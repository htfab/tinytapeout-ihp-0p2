module tt_um_no_time_for_squares_tommythorn (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire clknet_leaf_0_clk;
 wire \clock_inst.frameno[0] ;
 wire \clock_inst.frameno[1] ;
 wire \clock_inst.frameno[2] ;
 wire \clock_inst.frameno[3] ;
 wire \clock_inst.frameno[4] ;
 wire \clock_inst.frameno[5] ;
 wire \clock_inst.frameno[6] ;
 wire \clock_inst.hour[0] ;
 wire \clock_inst.hour[1] ;
 wire \clock_inst.hour[2] ;
 wire \clock_inst.hour[3] ;
 wire \clock_inst.hour_a[0] ;
 wire \clock_inst.hour_a[10] ;
 wire \clock_inst.hour_a[18] ;
 wire \clock_inst.hour_a[19] ;
 wire \clock_inst.hour_a[1] ;
 wire \clock_inst.hour_a[20] ;
 wire \clock_inst.hour_a[21] ;
 wire \clock_inst.hour_a[22] ;
 wire \clock_inst.hour_a[23] ;
 wire \clock_inst.hour_a[24] ;
 wire \clock_inst.hour_a[2] ;
 wire \clock_inst.hour_a[36] ;
 wire \clock_inst.hour_a[37] ;
 wire \clock_inst.hour_a[38] ;
 wire \clock_inst.hour_a[39] ;
 wire \clock_inst.hour_a[3] ;
 wire \clock_inst.hour_a[40] ;
 wire \clock_inst.hour_a[41] ;
 wire \clock_inst.hour_a[42] ;
 wire \clock_inst.hour_a[43] ;
 wire \clock_inst.hour_a[44] ;
 wire \clock_inst.hour_a[4] ;
 wire \clock_inst.hour_a[5] ;
 wire \clock_inst.hour_a[6] ;
 wire \clock_inst.hour_a[7] ;
 wire \clock_inst.hour_b[0] ;
 wire \clock_inst.hour_b[10] ;
 wire \clock_inst.hour_b[19] ;
 wire \clock_inst.hour_b[1] ;
 wire \clock_inst.hour_b[20] ;
 wire \clock_inst.hour_b[21] ;
 wire \clock_inst.hour_b[22] ;
 wire \clock_inst.hour_b[23] ;
 wire \clock_inst.hour_b[2] ;
 wire \clock_inst.hour_b[36] ;
 wire \clock_inst.hour_b[37] ;
 wire \clock_inst.hour_b[38] ;
 wire \clock_inst.hour_b[39] ;
 wire \clock_inst.hour_b[40] ;
 wire \clock_inst.hour_b[41] ;
 wire \clock_inst.hour_b[42] ;
 wire \clock_inst.hour_b[4] ;
 wire \clock_inst.hour_b[5] ;
 wire \clock_inst.hour_c[0] ;
 wire \clock_inst.hour_c[10] ;
 wire \clock_inst.hour_c[11] ;
 wire \clock_inst.hour_c[12] ;
 wire \clock_inst.hour_c[13] ;
 wire \clock_inst.hour_c[14] ;
 wire \clock_inst.hour_c[15] ;
 wire \clock_inst.hour_c[16] ;
 wire \clock_inst.hour_c[17] ;
 wire \clock_inst.hour_c[19] ;
 wire \clock_inst.hour_c[1] ;
 wire \clock_inst.hour_c[21] ;
 wire \clock_inst.hour_c[23] ;
 wire \clock_inst.hour_c[24] ;
 wire \clock_inst.hour_c[25] ;
 wire \clock_inst.hour_c[26] ;
 wire \clock_inst.hour_c[27] ;
 wire \clock_inst.hour_c[28] ;
 wire \clock_inst.hour_c[29] ;
 wire \clock_inst.hour_c[2] ;
 wire \clock_inst.hour_c[30] ;
 wire \clock_inst.hour_c[32] ;
 wire \clock_inst.hour_c[33] ;
 wire \clock_inst.hour_c[37] ;
 wire \clock_inst.hour_c[40] ;
 wire \clock_inst.hour_c[41] ;
 wire \clock_inst.hour_c[42] ;
 wire \clock_inst.hour_c[43] ;
 wire \clock_inst.hour_c[44] ;
 wire \clock_inst.hour_c[45] ;
 wire \clock_inst.hour_c[46] ;
 wire \clock_inst.hour_c[49] ;
 wire \clock_inst.hour_c[50] ;
 wire \clock_inst.hour_c[51] ;
 wire \clock_inst.hour_c[52] ;
 wire \clock_inst.hour_c[5] ;
 wire \clock_inst.hour_c[6] ;
 wire \clock_inst.hour_c[7] ;
 wire \clock_inst.hour_c[8] ;
 wire \clock_inst.hour_c[9] ;
 wire \clock_inst.hour_tile.e0[0] ;
 wire \clock_inst.hour_tile.e0[10] ;
 wire \clock_inst.hour_tile.e0[11] ;
 wire \clock_inst.hour_tile.e0[12] ;
 wire \clock_inst.hour_tile.e0[13] ;
 wire \clock_inst.hour_tile.e0[14] ;
 wire \clock_inst.hour_tile.e0[15] ;
 wire \clock_inst.hour_tile.e0[16] ;
 wire \clock_inst.hour_tile.e0[17] ;
 wire \clock_inst.hour_tile.e0[18] ;
 wire \clock_inst.hour_tile.e0[19] ;
 wire \clock_inst.hour_tile.e0[1] ;
 wire \clock_inst.hour_tile.e0[20] ;
 wire \clock_inst.hour_tile.e0[21] ;
 wire \clock_inst.hour_tile.e0[22] ;
 wire \clock_inst.hour_tile.e0[23] ;
 wire \clock_inst.hour_tile.e0[24] ;
 wire \clock_inst.hour_tile.e0[25] ;
 wire \clock_inst.hour_tile.e0[26] ;
 wire \clock_inst.hour_tile.e0[27] ;
 wire \clock_inst.hour_tile.e0[28] ;
 wire \clock_inst.hour_tile.e0[29] ;
 wire \clock_inst.hour_tile.e0[2] ;
 wire \clock_inst.hour_tile.e0[30] ;
 wire \clock_inst.hour_tile.e0[31] ;
 wire \clock_inst.hour_tile.e0[32] ;
 wire \clock_inst.hour_tile.e0[33] ;
 wire \clock_inst.hour_tile.e0[34] ;
 wire \clock_inst.hour_tile.e0[35] ;
 wire \clock_inst.hour_tile.e0[36] ;
 wire \clock_inst.hour_tile.e0[37] ;
 wire \clock_inst.hour_tile.e0[38] ;
 wire \clock_inst.hour_tile.e0[39] ;
 wire \clock_inst.hour_tile.e0[3] ;
 wire \clock_inst.hour_tile.e0[40] ;
 wire \clock_inst.hour_tile.e0[41] ;
 wire \clock_inst.hour_tile.e0[42] ;
 wire \clock_inst.hour_tile.e0[43] ;
 wire \clock_inst.hour_tile.e0[44] ;
 wire \clock_inst.hour_tile.e0[45] ;
 wire \clock_inst.hour_tile.e0[46] ;
 wire \clock_inst.hour_tile.e0[47] ;
 wire \clock_inst.hour_tile.e0[48] ;
 wire \clock_inst.hour_tile.e0[49] ;
 wire \clock_inst.hour_tile.e0[4] ;
 wire \clock_inst.hour_tile.e0[50] ;
 wire \clock_inst.hour_tile.e0[51] ;
 wire \clock_inst.hour_tile.e0[52] ;
 wire \clock_inst.hour_tile.e0[53] ;
 wire \clock_inst.hour_tile.e0[5] ;
 wire \clock_inst.hour_tile.e0[6] ;
 wire \clock_inst.hour_tile.e0[7] ;
 wire \clock_inst.hour_tile.e0[8] ;
 wire \clock_inst.hour_tile.e0[9] ;
 wire \clock_inst.hour_tile.e[0] ;
 wire \clock_inst.hour_tile.e[10] ;
 wire \clock_inst.hour_tile.e[11] ;
 wire \clock_inst.hour_tile.e[12] ;
 wire \clock_inst.hour_tile.e[13] ;
 wire \clock_inst.hour_tile.e[14] ;
 wire \clock_inst.hour_tile.e[15] ;
 wire \clock_inst.hour_tile.e[16] ;
 wire \clock_inst.hour_tile.e[17] ;
 wire \clock_inst.hour_tile.e[18] ;
 wire \clock_inst.hour_tile.e[19] ;
 wire \clock_inst.hour_tile.e[1] ;
 wire \clock_inst.hour_tile.e[20] ;
 wire \clock_inst.hour_tile.e[21] ;
 wire \clock_inst.hour_tile.e[22] ;
 wire \clock_inst.hour_tile.e[23] ;
 wire \clock_inst.hour_tile.e[24] ;
 wire \clock_inst.hour_tile.e[25] ;
 wire \clock_inst.hour_tile.e[26] ;
 wire \clock_inst.hour_tile.e[27] ;
 wire \clock_inst.hour_tile.e[28] ;
 wire \clock_inst.hour_tile.e[29] ;
 wire \clock_inst.hour_tile.e[2] ;
 wire \clock_inst.hour_tile.e[30] ;
 wire \clock_inst.hour_tile.e[31] ;
 wire \clock_inst.hour_tile.e[32] ;
 wire \clock_inst.hour_tile.e[33] ;
 wire \clock_inst.hour_tile.e[34] ;
 wire \clock_inst.hour_tile.e[35] ;
 wire \clock_inst.hour_tile.e[36] ;
 wire \clock_inst.hour_tile.e[37] ;
 wire \clock_inst.hour_tile.e[38] ;
 wire \clock_inst.hour_tile.e[39] ;
 wire \clock_inst.hour_tile.e[3] ;
 wire \clock_inst.hour_tile.e[40] ;
 wire \clock_inst.hour_tile.e[41] ;
 wire \clock_inst.hour_tile.e[42] ;
 wire \clock_inst.hour_tile.e[43] ;
 wire \clock_inst.hour_tile.e[44] ;
 wire \clock_inst.hour_tile.e[45] ;
 wire \clock_inst.hour_tile.e[46] ;
 wire \clock_inst.hour_tile.e[47] ;
 wire \clock_inst.hour_tile.e[48] ;
 wire \clock_inst.hour_tile.e[49] ;
 wire \clock_inst.hour_tile.e[4] ;
 wire \clock_inst.hour_tile.e[50] ;
 wire \clock_inst.hour_tile.e[51] ;
 wire \clock_inst.hour_tile.e[52] ;
 wire \clock_inst.hour_tile.e[53] ;
 wire \clock_inst.hour_tile.e[5] ;
 wire \clock_inst.hour_tile.e[6] ;
 wire \clock_inst.hour_tile.e[7] ;
 wire \clock_inst.hour_tile.e[8] ;
 wire \clock_inst.hour_tile.e[9] ;
 wire \clock_inst.min_a[0] ;
 wire \clock_inst.min_a[10] ;
 wire \clock_inst.min_a[18] ;
 wire \clock_inst.min_a[19] ;
 wire \clock_inst.min_a[1] ;
 wire \clock_inst.min_a[20] ;
 wire \clock_inst.min_a[21] ;
 wire \clock_inst.min_a[22] ;
 wire \clock_inst.min_a[23] ;
 wire \clock_inst.min_a[24] ;
 wire \clock_inst.min_a[2] ;
 wire \clock_inst.min_a[36] ;
 wire \clock_inst.min_a[37] ;
 wire \clock_inst.min_a[38] ;
 wire \clock_inst.min_a[39] ;
 wire \clock_inst.min_a[3] ;
 wire \clock_inst.min_a[40] ;
 wire \clock_inst.min_a[41] ;
 wire \clock_inst.min_a[42] ;
 wire \clock_inst.min_a[43] ;
 wire \clock_inst.min_a[44] ;
 wire \clock_inst.min_a[45] ;
 wire \clock_inst.min_a[4] ;
 wire \clock_inst.min_a[5] ;
 wire \clock_inst.min_a[6] ;
 wire \clock_inst.min_a[7] ;
 wire \clock_inst.min_a[8] ;
 wire \clock_inst.min_b[0] ;
 wire \clock_inst.min_b[10] ;
 wire \clock_inst.min_b[19] ;
 wire \clock_inst.min_b[1] ;
 wire \clock_inst.min_b[20] ;
 wire \clock_inst.min_b[21] ;
 wire \clock_inst.min_b[22] ;
 wire \clock_inst.min_b[23] ;
 wire \clock_inst.min_b[24] ;
 wire \clock_inst.min_b[2] ;
 wire \clock_inst.min_b[36] ;
 wire \clock_inst.min_b[37] ;
 wire \clock_inst.min_b[38] ;
 wire \clock_inst.min_b[39] ;
 wire \clock_inst.min_b[3] ;
 wire \clock_inst.min_b[40] ;
 wire \clock_inst.min_b[41] ;
 wire \clock_inst.min_b[42] ;
 wire \clock_inst.min_b[43] ;
 wire \clock_inst.min_b[44] ;
 wire \clock_inst.min_b[4] ;
 wire \clock_inst.min_b[5] ;
 wire \clock_inst.min_b[6] ;
 wire \clock_inst.min_b[7] ;
 wire \clock_inst.min_b[8] ;
 wire \clock_inst.min_c[0] ;
 wire \clock_inst.min_c[10] ;
 wire \clock_inst.min_c[11] ;
 wire \clock_inst.min_c[12] ;
 wire \clock_inst.min_c[13] ;
 wire \clock_inst.min_c[14] ;
 wire \clock_inst.min_c[15] ;
 wire \clock_inst.min_c[16] ;
 wire \clock_inst.min_c[17] ;
 wire \clock_inst.min_c[19] ;
 wire \clock_inst.min_c[1] ;
 wire \clock_inst.min_c[21] ;
 wire \clock_inst.min_c[22] ;
 wire \clock_inst.min_c[23] ;
 wire \clock_inst.min_c[24] ;
 wire \clock_inst.min_c[25] ;
 wire \clock_inst.min_c[26] ;
 wire \clock_inst.min_c[27] ;
 wire \clock_inst.min_c[28] ;
 wire \clock_inst.min_c[29] ;
 wire \clock_inst.min_c[2] ;
 wire \clock_inst.min_c[30] ;
 wire \clock_inst.min_c[31] ;
 wire \clock_inst.min_c[32] ;
 wire \clock_inst.min_c[33] ;
 wire \clock_inst.min_c[36] ;
 wire \clock_inst.min_c[37] ;
 wire \clock_inst.min_c[38] ;
 wire \clock_inst.min_c[39] ;
 wire \clock_inst.min_c[3] ;
 wire \clock_inst.min_c[40] ;
 wire \clock_inst.min_c[41] ;
 wire \clock_inst.min_c[42] ;
 wire \clock_inst.min_c[43] ;
 wire \clock_inst.min_c[44] ;
 wire \clock_inst.min_c[45] ;
 wire \clock_inst.min_c[46] ;
 wire \clock_inst.min_c[47] ;
 wire \clock_inst.min_c[48] ;
 wire \clock_inst.min_c[49] ;
 wire \clock_inst.min_c[4] ;
 wire \clock_inst.min_c[50] ;
 wire \clock_inst.min_c[51] ;
 wire \clock_inst.min_c[52] ;
 wire \clock_inst.min_c[53] ;
 wire \clock_inst.min_c[5] ;
 wire \clock_inst.min_c[6] ;
 wire \clock_inst.min_c[7] ;
 wire \clock_inst.min_c[8] ;
 wire \clock_inst.min_c[9] ;
 wire \clock_inst.min_tile.e0[0] ;
 wire \clock_inst.min_tile.e0[10] ;
 wire \clock_inst.min_tile.e0[11] ;
 wire \clock_inst.min_tile.e0[12] ;
 wire \clock_inst.min_tile.e0[13] ;
 wire \clock_inst.min_tile.e0[14] ;
 wire \clock_inst.min_tile.e0[15] ;
 wire \clock_inst.min_tile.e0[16] ;
 wire \clock_inst.min_tile.e0[17] ;
 wire \clock_inst.min_tile.e0[18] ;
 wire \clock_inst.min_tile.e0[19] ;
 wire \clock_inst.min_tile.e0[1] ;
 wire \clock_inst.min_tile.e0[20] ;
 wire \clock_inst.min_tile.e0[21] ;
 wire \clock_inst.min_tile.e0[22] ;
 wire \clock_inst.min_tile.e0[23] ;
 wire \clock_inst.min_tile.e0[24] ;
 wire \clock_inst.min_tile.e0[25] ;
 wire \clock_inst.min_tile.e0[26] ;
 wire \clock_inst.min_tile.e0[27] ;
 wire \clock_inst.min_tile.e0[28] ;
 wire \clock_inst.min_tile.e0[29] ;
 wire \clock_inst.min_tile.e0[2] ;
 wire \clock_inst.min_tile.e0[30] ;
 wire \clock_inst.min_tile.e0[31] ;
 wire \clock_inst.min_tile.e0[32] ;
 wire \clock_inst.min_tile.e0[33] ;
 wire \clock_inst.min_tile.e0[34] ;
 wire \clock_inst.min_tile.e0[35] ;
 wire \clock_inst.min_tile.e0[36] ;
 wire \clock_inst.min_tile.e0[37] ;
 wire \clock_inst.min_tile.e0[38] ;
 wire \clock_inst.min_tile.e0[39] ;
 wire \clock_inst.min_tile.e0[3] ;
 wire \clock_inst.min_tile.e0[40] ;
 wire \clock_inst.min_tile.e0[41] ;
 wire \clock_inst.min_tile.e0[42] ;
 wire \clock_inst.min_tile.e0[43] ;
 wire \clock_inst.min_tile.e0[44] ;
 wire \clock_inst.min_tile.e0[45] ;
 wire \clock_inst.min_tile.e0[46] ;
 wire \clock_inst.min_tile.e0[47] ;
 wire \clock_inst.min_tile.e0[48] ;
 wire \clock_inst.min_tile.e0[49] ;
 wire \clock_inst.min_tile.e0[4] ;
 wire \clock_inst.min_tile.e0[50] ;
 wire \clock_inst.min_tile.e0[51] ;
 wire \clock_inst.min_tile.e0[52] ;
 wire \clock_inst.min_tile.e0[53] ;
 wire \clock_inst.min_tile.e0[5] ;
 wire \clock_inst.min_tile.e0[6] ;
 wire \clock_inst.min_tile.e0[7] ;
 wire \clock_inst.min_tile.e0[8] ;
 wire \clock_inst.min_tile.e0[9] ;
 wire \clock_inst.min_tile.e[0] ;
 wire \clock_inst.min_tile.e[10] ;
 wire \clock_inst.min_tile.e[11] ;
 wire \clock_inst.min_tile.e[12] ;
 wire \clock_inst.min_tile.e[13] ;
 wire \clock_inst.min_tile.e[14] ;
 wire \clock_inst.min_tile.e[15] ;
 wire \clock_inst.min_tile.e[16] ;
 wire \clock_inst.min_tile.e[17] ;
 wire \clock_inst.min_tile.e[18] ;
 wire \clock_inst.min_tile.e[19] ;
 wire \clock_inst.min_tile.e[1] ;
 wire \clock_inst.min_tile.e[20] ;
 wire \clock_inst.min_tile.e[21] ;
 wire \clock_inst.min_tile.e[22] ;
 wire \clock_inst.min_tile.e[23] ;
 wire \clock_inst.min_tile.e[24] ;
 wire \clock_inst.min_tile.e[25] ;
 wire \clock_inst.min_tile.e[26] ;
 wire \clock_inst.min_tile.e[27] ;
 wire \clock_inst.min_tile.e[28] ;
 wire \clock_inst.min_tile.e[29] ;
 wire \clock_inst.min_tile.e[2] ;
 wire \clock_inst.min_tile.e[30] ;
 wire \clock_inst.min_tile.e[31] ;
 wire \clock_inst.min_tile.e[32] ;
 wire \clock_inst.min_tile.e[33] ;
 wire \clock_inst.min_tile.e[34] ;
 wire \clock_inst.min_tile.e[35] ;
 wire \clock_inst.min_tile.e[36] ;
 wire \clock_inst.min_tile.e[37] ;
 wire \clock_inst.min_tile.e[38] ;
 wire \clock_inst.min_tile.e[39] ;
 wire \clock_inst.min_tile.e[3] ;
 wire \clock_inst.min_tile.e[40] ;
 wire \clock_inst.min_tile.e[41] ;
 wire \clock_inst.min_tile.e[42] ;
 wire \clock_inst.min_tile.e[43] ;
 wire \clock_inst.min_tile.e[44] ;
 wire \clock_inst.min_tile.e[45] ;
 wire \clock_inst.min_tile.e[46] ;
 wire \clock_inst.min_tile.e[47] ;
 wire \clock_inst.min_tile.e[48] ;
 wire \clock_inst.min_tile.e[49] ;
 wire \clock_inst.min_tile.e[4] ;
 wire \clock_inst.min_tile.e[50] ;
 wire \clock_inst.min_tile.e[51] ;
 wire \clock_inst.min_tile.e[52] ;
 wire \clock_inst.min_tile.e[53] ;
 wire \clock_inst.min_tile.e[5] ;
 wire \clock_inst.min_tile.e[6] ;
 wire \clock_inst.min_tile.e[7] ;
 wire \clock_inst.min_tile.e[8] ;
 wire \clock_inst.min_tile.e[9] ;
 wire \clock_inst.minute[0] ;
 wire \clock_inst.minute[1] ;
 wire \clock_inst.minute[2] ;
 wire \clock_inst.minute[3] ;
 wire \clock_inst.minute[4] ;
 wire \clock_inst.minute[5] ;
 wire \clock_inst.sec_a[0] ;
 wire \clock_inst.sec_a[10] ;
 wire \clock_inst.sec_a[18] ;
 wire \clock_inst.sec_a[19] ;
 wire \clock_inst.sec_a[1] ;
 wire \clock_inst.sec_a[20] ;
 wire \clock_inst.sec_a[21] ;
 wire \clock_inst.sec_a[2] ;
 wire \clock_inst.sec_a[36] ;
 wire \clock_inst.sec_a[37] ;
 wire \clock_inst.sec_a[38] ;
 wire \clock_inst.sec_a[39] ;
 wire \clock_inst.sec_a[3] ;
 wire \clock_inst.sec_a[40] ;
 wire \clock_inst.sec_a[41] ;
 wire \clock_inst.sec_a[42] ;
 wire \clock_inst.sec_a[43] ;
 wire \clock_inst.sec_a[44] ;
 wire \clock_inst.sec_a[4] ;
 wire \clock_inst.sec_a[5] ;
 wire \clock_inst.sec_a[6] ;
 wire \clock_inst.sec_a[7] ;
 wire \clock_inst.sec_b[0] ;
 wire \clock_inst.sec_b[10] ;
 wire \clock_inst.sec_b[19] ;
 wire \clock_inst.sec_b[1] ;
 wire \clock_inst.sec_b[20] ;
 wire \clock_inst.sec_b[21] ;
 wire \clock_inst.sec_b[2] ;
 wire \clock_inst.sec_b[36] ;
 wire \clock_inst.sec_b[37] ;
 wire \clock_inst.sec_b[38] ;
 wire \clock_inst.sec_b[39] ;
 wire \clock_inst.sec_b[3] ;
 wire \clock_inst.sec_b[40] ;
 wire \clock_inst.sec_b[41] ;
 wire \clock_inst.sec_b[42] ;
 wire \clock_inst.sec_b[43] ;
 wire \clock_inst.sec_b[4] ;
 wire \clock_inst.sec_b[5] ;
 wire \clock_inst.sec_b[6] ;
 wire \clock_inst.sec_b[7] ;
 wire \clock_inst.sec_c[0] ;
 wire \clock_inst.sec_c[10] ;
 wire \clock_inst.sec_c[11] ;
 wire \clock_inst.sec_c[12] ;
 wire \clock_inst.sec_c[13] ;
 wire \clock_inst.sec_c[14] ;
 wire \clock_inst.sec_c[15] ;
 wire \clock_inst.sec_c[16] ;
 wire \clock_inst.sec_c[17] ;
 wire \clock_inst.sec_c[19] ;
 wire \clock_inst.sec_c[1] ;
 wire \clock_inst.sec_c[20] ;
 wire \clock_inst.sec_c[21] ;
 wire \clock_inst.sec_c[22] ;
 wire \clock_inst.sec_c[23] ;
 wire \clock_inst.sec_c[24] ;
 wire \clock_inst.sec_c[25] ;
 wire \clock_inst.sec_c[26] ;
 wire \clock_inst.sec_c[27] ;
 wire \clock_inst.sec_c[28] ;
 wire \clock_inst.sec_c[29] ;
 wire \clock_inst.sec_c[2] ;
 wire \clock_inst.sec_c[30] ;
 wire \clock_inst.sec_c[36] ;
 wire \clock_inst.sec_c[37] ;
 wire \clock_inst.sec_c[38] ;
 wire \clock_inst.sec_c[39] ;
 wire \clock_inst.sec_c[3] ;
 wire \clock_inst.sec_c[40] ;
 wire \clock_inst.sec_c[41] ;
 wire \clock_inst.sec_c[42] ;
 wire \clock_inst.sec_c[43] ;
 wire \clock_inst.sec_c[44] ;
 wire \clock_inst.sec_c[45] ;
 wire \clock_inst.sec_c[46] ;
 wire \clock_inst.sec_c[47] ;
 wire \clock_inst.sec_c[48] ;
 wire \clock_inst.sec_c[49] ;
 wire \clock_inst.sec_c[4] ;
 wire \clock_inst.sec_c[50] ;
 wire \clock_inst.sec_c[51] ;
 wire \clock_inst.sec_c[52] ;
 wire \clock_inst.sec_c[53] ;
 wire \clock_inst.sec_c[5] ;
 wire \clock_inst.sec_c[6] ;
 wire \clock_inst.sec_c[7] ;
 wire \clock_inst.sec_c[8] ;
 wire \clock_inst.sec_c[9] ;
 wire \clock_inst.sec_tile.e0[0] ;
 wire \clock_inst.sec_tile.e0[10] ;
 wire \clock_inst.sec_tile.e0[11] ;
 wire \clock_inst.sec_tile.e0[12] ;
 wire \clock_inst.sec_tile.e0[13] ;
 wire \clock_inst.sec_tile.e0[14] ;
 wire \clock_inst.sec_tile.e0[15] ;
 wire \clock_inst.sec_tile.e0[16] ;
 wire \clock_inst.sec_tile.e0[17] ;
 wire \clock_inst.sec_tile.e0[18] ;
 wire \clock_inst.sec_tile.e0[19] ;
 wire \clock_inst.sec_tile.e0[1] ;
 wire \clock_inst.sec_tile.e0[20] ;
 wire \clock_inst.sec_tile.e0[21] ;
 wire \clock_inst.sec_tile.e0[22] ;
 wire \clock_inst.sec_tile.e0[23] ;
 wire \clock_inst.sec_tile.e0[24] ;
 wire \clock_inst.sec_tile.e0[25] ;
 wire \clock_inst.sec_tile.e0[26] ;
 wire \clock_inst.sec_tile.e0[27] ;
 wire \clock_inst.sec_tile.e0[28] ;
 wire \clock_inst.sec_tile.e0[29] ;
 wire \clock_inst.sec_tile.e0[2] ;
 wire \clock_inst.sec_tile.e0[30] ;
 wire \clock_inst.sec_tile.e0[31] ;
 wire \clock_inst.sec_tile.e0[32] ;
 wire \clock_inst.sec_tile.e0[33] ;
 wire \clock_inst.sec_tile.e0[34] ;
 wire \clock_inst.sec_tile.e0[35] ;
 wire \clock_inst.sec_tile.e0[36] ;
 wire \clock_inst.sec_tile.e0[37] ;
 wire \clock_inst.sec_tile.e0[38] ;
 wire \clock_inst.sec_tile.e0[39] ;
 wire \clock_inst.sec_tile.e0[3] ;
 wire \clock_inst.sec_tile.e0[40] ;
 wire \clock_inst.sec_tile.e0[41] ;
 wire \clock_inst.sec_tile.e0[42] ;
 wire \clock_inst.sec_tile.e0[43] ;
 wire \clock_inst.sec_tile.e0[44] ;
 wire \clock_inst.sec_tile.e0[45] ;
 wire \clock_inst.sec_tile.e0[46] ;
 wire \clock_inst.sec_tile.e0[47] ;
 wire \clock_inst.sec_tile.e0[48] ;
 wire \clock_inst.sec_tile.e0[49] ;
 wire \clock_inst.sec_tile.e0[4] ;
 wire \clock_inst.sec_tile.e0[50] ;
 wire \clock_inst.sec_tile.e0[51] ;
 wire \clock_inst.sec_tile.e0[52] ;
 wire \clock_inst.sec_tile.e0[53] ;
 wire \clock_inst.sec_tile.e0[5] ;
 wire \clock_inst.sec_tile.e0[6] ;
 wire \clock_inst.sec_tile.e0[7] ;
 wire \clock_inst.sec_tile.e0[8] ;
 wire \clock_inst.sec_tile.e0[9] ;
 wire \clock_inst.sec_tile.e[0] ;
 wire \clock_inst.sec_tile.e[10] ;
 wire \clock_inst.sec_tile.e[11] ;
 wire \clock_inst.sec_tile.e[12] ;
 wire \clock_inst.sec_tile.e[13] ;
 wire \clock_inst.sec_tile.e[14] ;
 wire \clock_inst.sec_tile.e[15] ;
 wire \clock_inst.sec_tile.e[16] ;
 wire \clock_inst.sec_tile.e[17] ;
 wire \clock_inst.sec_tile.e[18] ;
 wire \clock_inst.sec_tile.e[19] ;
 wire \clock_inst.sec_tile.e[1] ;
 wire \clock_inst.sec_tile.e[20] ;
 wire \clock_inst.sec_tile.e[21] ;
 wire \clock_inst.sec_tile.e[22] ;
 wire \clock_inst.sec_tile.e[23] ;
 wire \clock_inst.sec_tile.e[24] ;
 wire \clock_inst.sec_tile.e[25] ;
 wire \clock_inst.sec_tile.e[26] ;
 wire \clock_inst.sec_tile.e[27] ;
 wire \clock_inst.sec_tile.e[28] ;
 wire \clock_inst.sec_tile.e[29] ;
 wire \clock_inst.sec_tile.e[2] ;
 wire \clock_inst.sec_tile.e[30] ;
 wire \clock_inst.sec_tile.e[31] ;
 wire \clock_inst.sec_tile.e[32] ;
 wire \clock_inst.sec_tile.e[33] ;
 wire \clock_inst.sec_tile.e[34] ;
 wire \clock_inst.sec_tile.e[35] ;
 wire \clock_inst.sec_tile.e[36] ;
 wire \clock_inst.sec_tile.e[37] ;
 wire \clock_inst.sec_tile.e[38] ;
 wire \clock_inst.sec_tile.e[39] ;
 wire \clock_inst.sec_tile.e[3] ;
 wire \clock_inst.sec_tile.e[40] ;
 wire \clock_inst.sec_tile.e[41] ;
 wire \clock_inst.sec_tile.e[42] ;
 wire \clock_inst.sec_tile.e[43] ;
 wire \clock_inst.sec_tile.e[44] ;
 wire \clock_inst.sec_tile.e[45] ;
 wire \clock_inst.sec_tile.e[46] ;
 wire \clock_inst.sec_tile.e[47] ;
 wire \clock_inst.sec_tile.e[48] ;
 wire \clock_inst.sec_tile.e[49] ;
 wire \clock_inst.sec_tile.e[4] ;
 wire \clock_inst.sec_tile.e[50] ;
 wire \clock_inst.sec_tile.e[51] ;
 wire \clock_inst.sec_tile.e[52] ;
 wire \clock_inst.sec_tile.e[53] ;
 wire \clock_inst.sec_tile.e[5] ;
 wire \clock_inst.sec_tile.e[6] ;
 wire \clock_inst.sec_tile.e[7] ;
 wire \clock_inst.sec_tile.e[8] ;
 wire \clock_inst.sec_tile.e[9] ;
 wire \clock_inst.second[0] ;
 wire \clock_inst.second[1] ;
 wire \clock_inst.second[2] ;
 wire \clock_inst.second[3] ;
 wire \clock_inst.second[4] ;
 wire \clock_inst.second[5] ;
 wire \clock_inst.vga_horizontal_blank_strobe ;
 wire \clock_inst.vga_hs ;
 wire \clock_inst.vga_inst.vga_horizontal_visible ;
 wire \clock_inst.vga_inst.vga_vertical_blank_strobe ;
 wire \clock_inst.vga_inst.vga_vertical_visible ;
 wire \clock_inst.vga_inst.vga_vs ;
 wire \clock_inst.vga_inst.vga_x[0] ;
 wire \clock_inst.vga_inst.vga_x[1] ;
 wire \clock_inst.vga_inst.vga_x[2] ;
 wire \clock_inst.vga_inst.vga_x[3] ;
 wire \clock_inst.vga_inst.vga_x[4] ;
 wire \clock_inst.vga_inst.vga_x[5] ;
 wire \clock_inst.vga_inst.vga_x[6] ;
 wire \clock_inst.vga_inst.vga_x[7] ;
 wire \clock_inst.vga_inst.vga_x[8] ;
 wire \clock_inst.vga_inst.vga_x[9] ;
 wire \clock_inst.vga_inst.vga_y[0] ;
 wire \clock_inst.vga_inst.vga_y[1] ;
 wire \clock_inst.vga_inst.vga_y[2] ;
 wire \clock_inst.vga_inst.vga_y[3] ;
 wire \clock_inst.vga_inst.vga_y[4] ;
 wire \clock_inst.vga_inst.vga_y[5] ;
 wire \clock_inst.vga_inst.vga_y[6] ;
 wire \clock_inst.vga_inst.vga_y[7] ;
 wire \clock_inst.vga_inst.vga_y[8] ;
 wire \clock_inst.vga_inst.vga_y[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_97_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;

 sg13g2_inv_1 _08018_ (.Y(_00655_),
    .A(\clock_inst.hour_a[0] ));
 sg13g2_buf_1 _08019_ (.A(\clock_inst.vga_inst.vga_vertical_blank_strobe ),
    .X(_00656_));
 sg13g2_buf_1 _08020_ (.A(\clock_inst.hour[2] ),
    .X(_00657_));
 sg13g2_buf_2 _08021_ (.A(\clock_inst.hour[3] ),
    .X(_00658_));
 sg13g2_nand2_2 _08022_ (.Y(_00659_),
    .A(net582),
    .B(_00658_));
 sg13g2_nand2_1 _08023_ (.Y(_00660_),
    .A(net583),
    .B(_00659_));
 sg13g2_buf_1 _08024_ (.A(_00660_),
    .X(_00661_));
 sg13g2_buf_1 _08025_ (.A(_00661_),
    .X(_00662_));
 sg13g2_buf_1 _08026_ (.A(net365),
    .X(_00663_));
 sg13g2_buf_1 _08027_ (.A(\clock_inst.hour[0] ),
    .X(_00664_));
 sg13g2_inv_1 _08028_ (.Y(_00665_),
    .A(net581));
 sg13g2_buf_1 _08029_ (.A(_00665_),
    .X(_00666_));
 sg13g2_inv_1 _08030_ (.Y(_00667_),
    .A(net582));
 sg13g2_buf_1 _08031_ (.A(_00667_),
    .X(_00668_));
 sg13g2_nor2_1 _08032_ (.A(_00666_),
    .B(net516),
    .Y(_00669_));
 sg13g2_buf_1 _08033_ (.A(\clock_inst.hour[1] ),
    .X(_00670_));
 sg13g2_inv_1 _08034_ (.Y(_00671_),
    .A(_00658_));
 sg13g2_buf_2 _08035_ (.A(_00671_),
    .X(_00672_));
 sg13g2_nand2_1 _08036_ (.Y(_00673_),
    .A(net580),
    .B(net515));
 sg13g2_buf_1 _08037_ (.A(_00673_),
    .X(_00674_));
 sg13g2_buf_2 _08038_ (.A(net517),
    .X(_00675_));
 sg13g2_inv_2 _08039_ (.Y(_00676_),
    .A(net580));
 sg13g2_buf_1 _08040_ (.A(_00658_),
    .X(_00677_));
 sg13g2_nand2_2 _08041_ (.Y(_00678_),
    .A(_00676_),
    .B(net550));
 sg13g2_inv_1 _08042_ (.Y(_00679_),
    .A(_00678_));
 sg13g2_buf_2 _08043_ (.A(net516),
    .X(_00680_));
 sg13g2_o21ai_1 _08044_ (.B1(net453),
    .Y(_00681_),
    .A1(net454),
    .A2(_00679_));
 sg13g2_o21ai_1 _08045_ (.B1(_00681_),
    .Y(_00682_),
    .A1(_00669_),
    .A2(net364));
 sg13g2_buf_1 _08046_ (.A(net583),
    .X(_00683_));
 sg13g2_buf_1 _08047_ (.A(net549),
    .X(_00684_));
 sg13g2_buf_1 _08048_ (.A(net514),
    .X(_00685_));
 sg13g2_a22oi_1 _08049_ (.Y(_00015_),
    .B1(_00682_),
    .B2(net452),
    .A2(net245),
    .A1(_00655_));
 sg13g2_buf_1 _08050_ (.A(\clock_inst.hour_a[10] ),
    .X(_00686_));
 sg13g2_buf_1 _08051_ (.A(_00661_),
    .X(_00687_));
 sg13g2_inv_1 _08052_ (.Y(_00688_),
    .A(net583));
 sg13g2_buf_1 _08053_ (.A(_00688_),
    .X(_00689_));
 sg13g2_nor2_1 _08054_ (.A(net513),
    .B(net582),
    .Y(_00690_));
 sg13g2_buf_1 _08055_ (.A(_00690_),
    .X(_00691_));
 sg13g2_a22oi_1 _08056_ (.Y(_00692_),
    .B1(_00678_),
    .B2(_00691_),
    .A2(net363),
    .A1(_00686_));
 sg13g2_inv_1 _08057_ (.Y(_00016_),
    .A(_00692_));
 sg13g2_inv_1 _08058_ (.Y(_00693_),
    .A(\clock_inst.hour_a[19] ));
 sg13g2_buf_1 _08059_ (.A(net580),
    .X(_00694_));
 sg13g2_buf_1 _08060_ (.A(net548),
    .X(_00695_));
 sg13g2_nor2_2 _08061_ (.A(net582),
    .B(_00658_),
    .Y(_00696_));
 sg13g2_inv_1 _08062_ (.Y(_00697_),
    .A(_00696_));
 sg13g2_buf_1 _08063_ (.A(_00664_),
    .X(_00698_));
 sg13g2_nand2_1 _08064_ (.Y(_00699_),
    .A(net547),
    .B(_00659_));
 sg13g2_o21ai_1 _08065_ (.B1(_00699_),
    .Y(_00700_),
    .A1(net512),
    .A2(_00697_));
 sg13g2_a22oi_1 _08066_ (.Y(_00017_),
    .B1(_00700_),
    .B2(net452),
    .A2(net245),
    .A1(_00693_));
 sg13g2_inv_1 _08067_ (.Y(_00701_),
    .A(\clock_inst.hour_a[1] ));
 sg13g2_and2_1 _08068_ (.A(net583),
    .B(_00659_),
    .X(_00702_));
 sg13g2_buf_1 _08069_ (.A(_00702_),
    .X(_00703_));
 sg13g2_nand2_1 _08070_ (.Y(_00704_),
    .A(_00657_),
    .B(_00671_));
 sg13g2_buf_2 _08071_ (.A(_00704_),
    .X(_00705_));
 sg13g2_nor2_1 _08072_ (.A(net517),
    .B(_00705_),
    .Y(_00706_));
 sg13g2_nand2_2 _08073_ (.Y(_00707_),
    .A(net517),
    .B(_00667_));
 sg13g2_a21oi_1 _08074_ (.A1(_00678_),
    .A2(net364),
    .Y(_00708_),
    .B1(_00707_));
 sg13g2_buf_1 _08075_ (.A(net549),
    .X(_00709_));
 sg13g2_o21ai_1 _08076_ (.B1(_00709_),
    .Y(_00710_),
    .A1(_00706_),
    .A2(_00708_));
 sg13g2_o21ai_1 _08077_ (.B1(_00710_),
    .Y(_00018_),
    .A1(_00701_),
    .A2(net451));
 sg13g2_inv_1 _08078_ (.Y(_00711_),
    .A(\clock_inst.hour_a[20] ));
 sg13g2_nor2_2 _08079_ (.A(net581),
    .B(net550),
    .Y(_00712_));
 sg13g2_nor2_1 _08080_ (.A(_00657_),
    .B(_00671_),
    .Y(_00713_));
 sg13g2_buf_2 _08081_ (.A(_00713_),
    .X(_00714_));
 sg13g2_nand2_1 _08082_ (.Y(_00715_),
    .A(net581),
    .B(_00714_));
 sg13g2_inv_1 _08083_ (.Y(_00716_),
    .A(_00715_));
 sg13g2_nor2_1 _08084_ (.A(_00712_),
    .B(_00716_),
    .Y(_00717_));
 sg13g2_buf_1 _08085_ (.A(_00694_),
    .X(_00718_));
 sg13g2_nand2_1 _08086_ (.Y(_00719_),
    .A(net510),
    .B(_00696_));
 sg13g2_o21ai_1 _08087_ (.B1(_00719_),
    .Y(_00720_),
    .A1(net512),
    .A2(_00717_));
 sg13g2_a22oi_1 _08088_ (.Y(_00019_),
    .B1(_00720_),
    .B2(net452),
    .A2(net245),
    .A1(_00711_));
 sg13g2_inv_1 _08089_ (.Y(_00721_),
    .A(\clock_inst.hour_a[21] ));
 sg13g2_nor2_2 _08090_ (.A(net513),
    .B(net550),
    .Y(_00722_));
 sg13g2_nand2_1 _08091_ (.Y(_00723_),
    .A(net548),
    .B(_00707_));
 sg13g2_a22oi_1 _08092_ (.Y(_00020_),
    .B1(_00722_),
    .B2(_00723_),
    .A2(_00663_),
    .A1(_00721_));
 sg13g2_buf_2 _08093_ (.A(\clock_inst.hour_a[22] ),
    .X(_00724_));
 sg13g2_inv_2 _08094_ (.Y(_00725_),
    .A(_00724_));
 sg13g2_nand2_1 _08095_ (.Y(_00726_),
    .A(_00699_),
    .B(_00697_));
 sg13g2_nand2_1 _08096_ (.Y(_00727_),
    .A(_00676_),
    .B(_00671_));
 sg13g2_nor2_1 _08097_ (.A(net581),
    .B(_00727_),
    .Y(_00728_));
 sg13g2_buf_2 _08098_ (.A(_00728_),
    .X(_00729_));
 sg13g2_a21o_1 _08099_ (.A2(_00726_),
    .A1(net512),
    .B1(_00729_),
    .X(_00730_));
 sg13g2_a22oi_1 _08100_ (.Y(_00021_),
    .B1(_00730_),
    .B2(net452),
    .A2(net245),
    .A1(_00725_));
 sg13g2_buf_8 _08101_ (.A(\clock_inst.hour_a[23] ),
    .X(_00731_));
 sg13g2_buf_1 _08102_ (.A(_00731_),
    .X(_00732_));
 sg13g2_nand2_1 _08103_ (.Y(_00733_),
    .A(net516),
    .B(_00658_));
 sg13g2_nor2_1 _08104_ (.A(_00698_),
    .B(_00733_),
    .Y(_00734_));
 sg13g2_buf_1 _08105_ (.A(net582),
    .X(_00735_));
 sg13g2_nand2_2 _08106_ (.Y(_00736_),
    .A(net581),
    .B(_00671_));
 sg13g2_buf_1 _08107_ (.A(net548),
    .X(_00737_));
 sg13g2_a21oi_1 _08108_ (.A1(net545),
    .A2(_00736_),
    .Y(_00738_),
    .B1(net509));
 sg13g2_o21ai_1 _08109_ (.B1(net514),
    .Y(_00739_),
    .A1(_00734_),
    .A2(_00738_));
 sg13g2_o21ai_1 _08110_ (.B1(_00739_),
    .Y(_00740_),
    .A1(_00732_),
    .A2(net451));
 sg13g2_inv_1 _08111_ (.Y(_00022_),
    .A(_00740_));
 sg13g2_buf_1 _08112_ (.A(\clock_inst.hour_a[2] ),
    .X(_00741_));
 sg13g2_buf_1 _08113_ (.A(net545),
    .X(_00742_));
 sg13g2_nand2_1 _08114_ (.Y(_00743_),
    .A(net517),
    .B(_00658_));
 sg13g2_nand2_1 _08115_ (.Y(_00744_),
    .A(_00736_),
    .B(_00743_));
 sg13g2_o21ai_1 _08116_ (.B1(net364),
    .Y(_00745_),
    .A1(net508),
    .A2(_00744_));
 sg13g2_buf_1 _08117_ (.A(net549),
    .X(_00746_));
 sg13g2_a22oi_1 _08118_ (.Y(_00747_),
    .B1(_00745_),
    .B2(_00746_),
    .A2(net363),
    .A1(_00741_));
 sg13g2_inv_1 _08119_ (.Y(_00023_),
    .A(_00747_));
 sg13g2_buf_1 _08120_ (.A(net513),
    .X(_00748_));
 sg13g2_nor2_1 _08121_ (.A(_00667_),
    .B(_00658_),
    .Y(_00749_));
 sg13g2_buf_2 _08122_ (.A(_00749_),
    .X(_00750_));
 sg13g2_a21oi_1 _08123_ (.A1(net548),
    .A2(_00750_),
    .Y(_00751_),
    .B1(_00714_));
 sg13g2_buf_1 _08124_ (.A(\clock_inst.hour_a[24] ),
    .X(_00752_));
 sg13g2_nand2_1 _08125_ (.Y(_00753_),
    .A(net583),
    .B(net515));
 sg13g2_buf_2 _08126_ (.A(_00753_),
    .X(_00754_));
 sg13g2_nand2_1 _08127_ (.Y(_00755_),
    .A(net579),
    .B(_00754_));
 sg13g2_o21ai_1 _08128_ (.B1(_00755_),
    .Y(_00024_),
    .A1(net450),
    .A2(_00751_));
 sg13g2_nand2_1 _08129_ (.Y(_00756_),
    .A(_00656_),
    .B(net516));
 sg13g2_buf_2 _08130_ (.A(_00756_),
    .X(_00757_));
 sg13g2_nor2_2 _08131_ (.A(net580),
    .B(net550),
    .Y(_00758_));
 sg13g2_a21oi_1 _08132_ (.A1(net509),
    .A2(_00714_),
    .Y(_00759_),
    .B1(_00758_));
 sg13g2_o21ai_1 _08133_ (.B1(_00705_),
    .Y(_00760_),
    .A1(net454),
    .A2(_00759_));
 sg13g2_a22oi_1 _08134_ (.Y(_00761_),
    .B1(_00760_),
    .B2(net507),
    .A2(_00757_),
    .A1(\clock_inst.hour_a[36] ));
 sg13g2_inv_1 _08135_ (.Y(_00025_),
    .A(_00761_));
 sg13g2_buf_1 _08136_ (.A(\clock_inst.hour_a[37] ),
    .X(_00762_));
 sg13g2_buf_1 _08137_ (.A(_00661_),
    .X(_00763_));
 sg13g2_nor2_2 _08138_ (.A(net517),
    .B(_00658_),
    .Y(_00764_));
 sg13g2_nand2_1 _08139_ (.Y(_00765_),
    .A(_00676_),
    .B(_00764_));
 sg13g2_buf_2 _08140_ (.A(_00765_),
    .X(_00766_));
 sg13g2_buf_1 _08141_ (.A(net550),
    .X(_00767_));
 sg13g2_nand2_1 _08142_ (.Y(_00768_),
    .A(_00718_),
    .B(net506));
 sg13g2_a21oi_1 _08143_ (.A1(_00766_),
    .A2(_00768_),
    .Y(_00769_),
    .B1(_00757_));
 sg13g2_a21o_1 _08144_ (.A2(net361),
    .A1(_00762_),
    .B1(_00769_),
    .X(_00026_));
 sg13g2_inv_1 _08145_ (.Y(_00770_),
    .A(\clock_inst.hour_a[38] ));
 sg13g2_o21ai_1 _08146_ (.B1(_00766_),
    .Y(_00771_),
    .A1(_00707_),
    .A2(_00758_));
 sg13g2_a22oi_1 _08147_ (.Y(_00027_),
    .B1(_00771_),
    .B2(net452),
    .A2(net245),
    .A1(_00770_));
 sg13g2_inv_1 _08148_ (.Y(_00772_),
    .A(\clock_inst.hour_a[39] ));
 sg13g2_nand2_1 _08149_ (.Y(_00773_),
    .A(_00694_),
    .B(_00764_));
 sg13g2_a22oi_1 _08150_ (.Y(_00028_),
    .B1(_00773_),
    .B2(net362),
    .A2(_00754_),
    .A1(_00772_));
 sg13g2_buf_1 _08151_ (.A(\clock_inst.hour_a[3] ),
    .X(_00774_));
 sg13g2_nand2_2 _08152_ (.Y(_00775_),
    .A(net580),
    .B(net547));
 sg13g2_a21oi_2 _08153_ (.B1(net545),
    .Y(_00776_),
    .A2(_00775_),
    .A1(_00677_));
 sg13g2_buf_1 _08154_ (.A(net549),
    .X(_00777_));
 sg13g2_a22oi_1 _08155_ (.Y(_00778_),
    .B1(_00776_),
    .B2(net505),
    .A2(net363),
    .A1(_00774_));
 sg13g2_inv_1 _08156_ (.Y(_00029_),
    .A(_00778_));
 sg13g2_inv_1 _08157_ (.Y(_00779_),
    .A(\clock_inst.hour_a[40] ));
 sg13g2_nor2_2 _08158_ (.A(net517),
    .B(net515),
    .Y(_00780_));
 sg13g2_o21ai_1 _08159_ (.B1(_00766_),
    .Y(_00781_),
    .A1(net508),
    .A2(_00780_));
 sg13g2_a22oi_1 _08160_ (.Y(_00030_),
    .B1(_00781_),
    .B2(_00685_),
    .A2(_00663_),
    .A1(_00779_));
 sg13g2_buf_1 _08161_ (.A(\clock_inst.hour_a[41] ),
    .X(_00782_));
 sg13g2_nor2_1 _08162_ (.A(_00670_),
    .B(_00707_),
    .Y(_00783_));
 sg13g2_nor2_1 _08163_ (.A(_00669_),
    .B(_00783_),
    .Y(_00784_));
 sg13g2_o21ai_1 _08164_ (.B1(_00718_),
    .Y(_00785_),
    .A1(_00734_),
    .A2(_00764_));
 sg13g2_o21ai_1 _08165_ (.B1(_00785_),
    .Y(_00786_),
    .A1(_00767_),
    .A2(_00784_));
 sg13g2_a22oi_1 _08166_ (.Y(_00787_),
    .B1(_00786_),
    .B2(net505),
    .A2(net363),
    .A1(_00782_));
 sg13g2_inv_1 _08167_ (.Y(_00031_),
    .A(_00787_));
 sg13g2_inv_1 _08168_ (.Y(_00788_),
    .A(\clock_inst.hour_a[42] ));
 sg13g2_nor2_1 _08169_ (.A(net517),
    .B(net582),
    .Y(_00789_));
 sg13g2_buf_2 _08170_ (.A(_00676_),
    .X(_00790_));
 sg13g2_o21ai_1 _08171_ (.B1(net504),
    .Y(_00791_),
    .A1(_00712_),
    .A2(_00789_));
 sg13g2_nand2_1 _08172_ (.Y(_00792_),
    .A(_00715_),
    .B(_00791_));
 sg13g2_a22oi_1 _08173_ (.Y(_00032_),
    .B1(_00792_),
    .B2(_00685_),
    .A2(net245),
    .A1(_00788_));
 sg13g2_buf_1 _08174_ (.A(\clock_inst.hour_a[43] ),
    .X(_00793_));
 sg13g2_nand2_2 _08175_ (.Y(_00794_),
    .A(net581),
    .B(net516));
 sg13g2_nor2_1 _08176_ (.A(_00676_),
    .B(_00794_),
    .Y(_00795_));
 sg13g2_a21oi_1 _08177_ (.A1(net454),
    .A2(_00659_),
    .Y(_00796_),
    .B1(_00696_));
 sg13g2_nor2_1 _08178_ (.A(_00737_),
    .B(_00796_),
    .Y(_00797_));
 sg13g2_or2_1 _08179_ (.X(_00798_),
    .B(_00797_),
    .A(_00795_));
 sg13g2_a22oi_1 _08180_ (.Y(_00799_),
    .B1(_00798_),
    .B2(net505),
    .A2(net363),
    .A1(_00793_));
 sg13g2_inv_1 _08181_ (.Y(_00033_),
    .A(_00799_));
 sg13g2_buf_1 _08182_ (.A(\clock_inst.hour_a[44] ),
    .X(_00800_));
 sg13g2_nor2_1 _08183_ (.A(net580),
    .B(_00664_),
    .Y(_00801_));
 sg13g2_nand2_1 _08184_ (.Y(_00802_),
    .A(_00714_),
    .B(_00801_));
 sg13g2_a21oi_1 _08185_ (.A1(_00773_),
    .A2(_00802_),
    .Y(_00803_),
    .B1(_00689_));
 sg13g2_a21oi_1 _08186_ (.A1(net450),
    .A2(_00800_),
    .Y(_00804_),
    .B1(_00803_));
 sg13g2_o21ai_1 _08187_ (.B1(net508),
    .Y(_00805_),
    .A1(_00800_),
    .A2(_00722_));
 sg13g2_nand2_1 _08188_ (.Y(_00034_),
    .A(_00804_),
    .B(_00805_));
 sg13g2_buf_2 _08189_ (.A(\clock_inst.hour_a[5] ),
    .X(_00806_));
 sg13g2_nor2_1 _08190_ (.A(net581),
    .B(_00705_),
    .Y(_00807_));
 sg13g2_o21ai_1 _08191_ (.B1(net509),
    .Y(_00808_),
    .A1(_00789_),
    .A2(_00807_));
 sg13g2_nor2_1 _08192_ (.A(net548),
    .B(_00743_),
    .Y(_00809_));
 sg13g2_o21ai_1 _08193_ (.B1(net453),
    .Y(_00810_),
    .A1(_00764_),
    .A2(_00809_));
 sg13g2_nand2_1 _08194_ (.Y(_00811_),
    .A(_00808_),
    .B(_00810_));
 sg13g2_a22oi_1 _08195_ (.Y(_00812_),
    .B1(_00811_),
    .B2(net505),
    .A2(net363),
    .A1(_00806_));
 sg13g2_inv_1 _08196_ (.Y(_00035_),
    .A(_00812_));
 sg13g2_buf_2 _08197_ (.A(\clock_inst.hour_a[6] ),
    .X(_00813_));
 sg13g2_inv_1 _08198_ (.Y(_00814_),
    .A(_00813_));
 sg13g2_nor2_1 _08199_ (.A(net580),
    .B(_00733_),
    .Y(_00815_));
 sg13g2_o21ai_1 _08200_ (.B1(net547),
    .Y(_00816_),
    .A1(_00750_),
    .A2(_00815_));
 sg13g2_nand2_1 _08201_ (.Y(_00817_),
    .A(net512),
    .B(_00712_));
 sg13g2_nand2_1 _08202_ (.Y(_00818_),
    .A(_00816_),
    .B(_00817_));
 sg13g2_a22oi_1 _08203_ (.Y(_00036_),
    .B1(_00818_),
    .B2(net452),
    .A2(net245),
    .A1(_00814_));
 sg13g2_buf_1 _08204_ (.A(\clock_inst.hour_a[7] ),
    .X(_00819_));
 sg13g2_inv_1 _08205_ (.Y(_00820_),
    .A(_00819_));
 sg13g2_o21ai_1 _08206_ (.B1(net504),
    .Y(_00821_),
    .A1(net516),
    .A2(_00712_));
 sg13g2_nand2_1 _08207_ (.Y(_00822_),
    .A(_00715_),
    .B(_00821_));
 sg13g2_a22oi_1 _08208_ (.Y(_00037_),
    .B1(_00822_),
    .B2(net452),
    .A2(net245),
    .A1(_00820_));
 sg13g2_buf_2 _08209_ (.A(\clock_inst.hour_b[0] ),
    .X(_00823_));
 sg13g2_inv_1 _08210_ (.Y(_00824_),
    .A(_00823_));
 sg13g2_buf_1 _08211_ (.A(_00661_),
    .X(_00825_));
 sg13g2_xnor2_1 _08212_ (.Y(_00826_),
    .A(net454),
    .B(_00758_));
 sg13g2_a22oi_1 _08213_ (.Y(_00038_),
    .B1(net362),
    .B2(_00826_),
    .A2(net360),
    .A1(_00824_));
 sg13g2_buf_1 _08214_ (.A(\clock_inst.hour_b[10] ),
    .X(_00827_));
 sg13g2_inv_1 _08215_ (.Y(_00828_),
    .A(net577));
 sg13g2_o21ai_1 _08216_ (.B1(net453),
    .Y(_00829_),
    .A1(net506),
    .A2(_00801_));
 sg13g2_o21ai_1 _08217_ (.B1(_00829_),
    .Y(_00830_),
    .A1(_00705_),
    .A2(_00775_));
 sg13g2_a22oi_1 _08218_ (.Y(_00039_),
    .B1(_00830_),
    .B2(net452),
    .A2(_00754_),
    .A1(_00828_));
 sg13g2_buf_2 _08219_ (.A(\clock_inst.hour_b[19] ),
    .X(_00831_));
 sg13g2_o21ai_1 _08220_ (.B1(net510),
    .Y(_00832_),
    .A1(_00750_),
    .A2(_00716_));
 sg13g2_nand2_1 _08221_ (.Y(_00833_),
    .A(_00766_),
    .B(_00832_));
 sg13g2_a22oi_1 _08222_ (.Y(_00834_),
    .B1(_00833_),
    .B2(net505),
    .A2(net363),
    .A1(_00831_));
 sg13g2_inv_1 _08223_ (.Y(_00040_),
    .A(_00834_));
 sg13g2_buf_2 _08224_ (.A(\clock_inst.hour_b[1] ),
    .X(_00835_));
 sg13g2_nor2_1 _08225_ (.A(_00670_),
    .B(_00666_),
    .Y(_00836_));
 sg13g2_buf_1 _08226_ (.A(_00836_),
    .X(_00837_));
 sg13g2_xnor2_1 _08227_ (.Y(_00838_),
    .A(_00672_),
    .B(net359));
 sg13g2_a22oi_1 _08228_ (.Y(_00839_),
    .B1(net362),
    .B2(_00838_),
    .A2(_00687_),
    .A1(_00835_));
 sg13g2_inv_1 _08229_ (.Y(_00041_),
    .A(_00839_));
 sg13g2_inv_1 _08230_ (.Y(_00840_),
    .A(\clock_inst.hour_b[20] ));
 sg13g2_nor2_2 _08231_ (.A(net580),
    .B(net582),
    .Y(_00841_));
 sg13g2_inv_1 _08232_ (.Y(_00842_),
    .A(_00744_));
 sg13g2_nand3_1 _08233_ (.B(net453),
    .C(_00842_),
    .A(net504),
    .Y(_00843_));
 sg13g2_o21ai_1 _08234_ (.B1(_00843_),
    .Y(_00844_),
    .A1(_00736_),
    .A2(_00841_));
 sg13g2_buf_1 _08235_ (.A(net514),
    .X(_00845_));
 sg13g2_a22oi_1 _08236_ (.Y(_00042_),
    .B1(_00844_),
    .B2(net449),
    .A2(_00825_),
    .A1(_00840_));
 sg13g2_inv_1 _08237_ (.Y(_00846_),
    .A(\clock_inst.hour_b[22] ));
 sg13g2_nor2_2 _08238_ (.A(net581),
    .B(net582),
    .Y(_00847_));
 sg13g2_o21ai_1 _08239_ (.B1(_00737_),
    .Y(_00848_),
    .A1(net515),
    .A2(_00847_));
 sg13g2_nand2_1 _08240_ (.Y(_00849_),
    .A(_00816_),
    .B(_00848_));
 sg13g2_a22oi_1 _08241_ (.Y(_00043_),
    .B1(_00849_),
    .B2(net449),
    .A2(net360),
    .A1(_00846_));
 sg13g2_inv_1 _08242_ (.Y(_00850_),
    .A(\clock_inst.hour_b[23] ));
 sg13g2_nand2_1 _08243_ (.Y(_00851_),
    .A(_00794_),
    .B(_00821_));
 sg13g2_a22oi_1 _08244_ (.Y(_00044_),
    .B1(_00851_),
    .B2(net449),
    .A2(net360),
    .A1(_00850_));
 sg13g2_buf_1 _08245_ (.A(\clock_inst.hour_b[2] ),
    .X(_00852_));
 sg13g2_inv_1 _08246_ (.Y(_00853_),
    .A(_00852_));
 sg13g2_nor2_2 _08247_ (.A(_00676_),
    .B(_00698_),
    .Y(_00854_));
 sg13g2_nor2_1 _08248_ (.A(_00837_),
    .B(_00854_),
    .Y(_00855_));
 sg13g2_a21oi_1 _08249_ (.A1(_00705_),
    .A2(_00733_),
    .Y(_00856_),
    .B1(_00689_));
 sg13g2_a22oi_1 _08250_ (.Y(_00045_),
    .B1(_00855_),
    .B2(_00856_),
    .A2(net360),
    .A1(_00853_));
 sg13g2_buf_1 _08251_ (.A(\clock_inst.hour_b[21] ),
    .X(_00857_));
 sg13g2_buf_1 _08252_ (.A(net576),
    .X(_00858_));
 sg13g2_nand2_1 _08253_ (.Y(_00859_),
    .A(net450),
    .B(net544));
 sg13g2_nand3b_1 _08254_ (.B(_00773_),
    .C(net514),
    .Y(_00860_),
    .A_N(_00815_));
 sg13g2_nand2_1 _08255_ (.Y(_00861_),
    .A(net544),
    .B(_00754_));
 sg13g2_a22oi_1 _08256_ (.Y(_00046_),
    .B1(_00861_),
    .B2(net508),
    .A2(_00860_),
    .A1(_00859_));
 sg13g2_buf_8 _08257_ (.A(\clock_inst.hour_b[36] ),
    .X(_00862_));
 sg13g2_inv_1 _08258_ (.Y(_00863_),
    .A(_00862_));
 sg13g2_o21ai_1 _08259_ (.B1(net453),
    .Y(_00864_),
    .A1(_00729_),
    .A2(_00780_));
 sg13g2_nand2_1 _08260_ (.Y(_00865_),
    .A(_00808_),
    .B(_00864_));
 sg13g2_a22oi_1 _08261_ (.Y(_00047_),
    .B1(_00865_),
    .B2(net449),
    .A2(net360),
    .A1(_00863_));
 sg13g2_buf_1 _08262_ (.A(\clock_inst.hour_b[37] ),
    .X(_00866_));
 sg13g2_and2_1 _08263_ (.A(_00723_),
    .B(_00784_),
    .X(_00867_));
 sg13g2_a22oi_1 _08264_ (.Y(_00868_),
    .B1(_00722_),
    .B2(_00867_),
    .A2(_00687_),
    .A1(_00866_));
 sg13g2_inv_1 _08265_ (.Y(_00048_),
    .A(_00868_));
 sg13g2_buf_8 _08266_ (.A(\clock_inst.hour_b[38] ),
    .X(_00869_));
 sg13g2_a21oi_1 _08267_ (.A1(net504),
    .A2(_00780_),
    .Y(_00870_),
    .B1(_00712_));
 sg13g2_o21ai_1 _08268_ (.B1(_00848_),
    .Y(_00871_),
    .A1(net508),
    .A2(_00870_));
 sg13g2_a22oi_1 _08269_ (.Y(_00872_),
    .B1(_00871_),
    .B2(net505),
    .A2(net363),
    .A1(_00869_));
 sg13g2_inv_1 _08270_ (.Y(_00049_),
    .A(_00872_));
 sg13g2_buf_8 _08271_ (.A(\clock_inst.hour_b[39] ),
    .X(_00873_));
 sg13g2_o21ai_1 _08272_ (.B1(_00684_),
    .Y(_00874_),
    .A1(_00758_),
    .A2(_00776_));
 sg13g2_o21ai_1 _08273_ (.B1(_00874_),
    .Y(_00875_),
    .A1(_00873_),
    .A2(_00703_));
 sg13g2_inv_1 _08274_ (.Y(_00050_),
    .A(_00875_));
 sg13g2_buf_2 _08275_ (.A(\clock_inst.hour_b[40] ),
    .X(_00876_));
 sg13g2_o21ai_1 _08276_ (.B1(net548),
    .Y(_00877_),
    .A1(_00706_),
    .A2(_00847_));
 sg13g2_o21ai_1 _08277_ (.B1(_00877_),
    .Y(_00878_),
    .A1(net508),
    .A2(_00870_));
 sg13g2_a22oi_1 _08278_ (.Y(_00879_),
    .B1(_00878_),
    .B2(net505),
    .A2(net365),
    .A1(_00876_));
 sg13g2_inv_1 _08279_ (.Y(_00051_),
    .A(_00879_));
 sg13g2_buf_8 _08280_ (.A(\clock_inst.hour_b[41] ),
    .X(_00880_));
 sg13g2_buf_1 _08281_ (.A(net547),
    .X(_00881_));
 sg13g2_nand2_1 _08282_ (.Y(_00882_),
    .A(net503),
    .B(_00696_));
 sg13g2_o21ai_1 _08283_ (.B1(_00882_),
    .Y(_00883_),
    .A1(net503),
    .A2(_00751_));
 sg13g2_a22oi_1 _08284_ (.Y(_00884_),
    .B1(_00883_),
    .B2(_00777_),
    .A2(net365),
    .A1(_00880_));
 sg13g2_inv_1 _08285_ (.Y(_00052_),
    .A(_00884_));
 sg13g2_nor2_1 _08286_ (.A(net547),
    .B(net516),
    .Y(_00885_));
 sg13g2_a21oi_1 _08287_ (.A1(net512),
    .A2(_00885_),
    .Y(_00886_),
    .B1(net359));
 sg13g2_buf_1 _08288_ (.A(\clock_inst.hour_b[42] ),
    .X(_00887_));
 sg13g2_a21oi_1 _08289_ (.A1(net511),
    .A2(_00659_),
    .Y(_00888_),
    .B1(_00887_));
 sg13g2_a21oi_1 _08290_ (.A1(_00722_),
    .A2(_00886_),
    .Y(_00053_),
    .B1(_00888_));
 sg13g2_buf_2 _08291_ (.A(\clock_inst.hour_b[4] ),
    .X(_00889_));
 sg13g2_o21ai_1 _08292_ (.B1(net453),
    .Y(_00890_),
    .A1(net515),
    .A2(_00854_));
 sg13g2_nand2_1 _08293_ (.Y(_00891_),
    .A(_00766_),
    .B(_00890_));
 sg13g2_a22oi_1 _08294_ (.Y(_00892_),
    .B1(_00891_),
    .B2(_00777_),
    .A2(_00662_),
    .A1(_00889_));
 sg13g2_inv_1 _08295_ (.Y(_00054_),
    .A(_00892_));
 sg13g2_inv_1 _08296_ (.Y(_00893_),
    .A(\clock_inst.hour_b[5] ));
 sg13g2_nor2_1 _08297_ (.A(_00754_),
    .B(_00841_),
    .Y(_00894_));
 sg13g2_a21oi_1 _08298_ (.A1(_00735_),
    .A2(_00893_),
    .Y(_00895_),
    .B1(_00894_));
 sg13g2_a221oi_1 _08299_ (.B2(net362),
    .C1(net503),
    .B1(_00674_),
    .A1(net550),
    .Y(_00896_),
    .A2(_00893_));
 sg13g2_a21oi_1 _08300_ (.A1(net503),
    .A2(_00895_),
    .Y(_00897_),
    .B1(_00896_));
 sg13g2_a21oi_1 _08301_ (.A1(_00748_),
    .A2(_00893_),
    .Y(_00055_),
    .B1(_00897_));
 sg13g2_inv_1 _08302_ (.Y(_00898_),
    .A(\clock_inst.hour_c[10] ));
 sg13g2_nand2_1 _08303_ (.Y(_00899_),
    .A(net517),
    .B(net545));
 sg13g2_nand2_1 _08304_ (.Y(_00900_),
    .A(_00794_),
    .B(_00899_));
 sg13g2_o21ai_1 _08305_ (.B1(_00715_),
    .Y(_00901_),
    .A1(net364),
    .A2(_00900_));
 sg13g2_a22oi_1 _08306_ (.Y(_00056_),
    .B1(_00901_),
    .B2(net449),
    .A2(net360),
    .A1(_00898_));
 sg13g2_inv_1 _08307_ (.Y(_00902_),
    .A(\clock_inst.hour_c[11] ));
 sg13g2_nand2_1 _08308_ (.Y(_00903_),
    .A(net504),
    .B(_00780_));
 sg13g2_nand2_1 _08309_ (.Y(_00904_),
    .A(net548),
    .B(_00744_));
 sg13g2_a21oi_1 _08310_ (.A1(_00903_),
    .A2(_00904_),
    .Y(_00905_),
    .B1(net545));
 sg13g2_and2_1 _08311_ (.A(_00750_),
    .B(_00854_),
    .X(_00906_));
 sg13g2_o21ai_1 _08312_ (.B1(net511),
    .Y(_00907_),
    .A1(_00905_),
    .A2(_00906_));
 sg13g2_o21ai_1 _08313_ (.B1(_00907_),
    .Y(_00057_),
    .A1(_00902_),
    .A2(net451));
 sg13g2_nand2_1 _08314_ (.Y(_00908_),
    .A(net548),
    .B(_00668_));
 sg13g2_a21oi_1 _08315_ (.A1(_00677_),
    .A2(_00908_),
    .Y(_00909_),
    .B1(net547));
 sg13g2_o21ai_1 _08316_ (.B1(net514),
    .Y(_00910_),
    .A1(_00758_),
    .A2(_00909_));
 sg13g2_o21ai_1 _08317_ (.B1(_00910_),
    .Y(_00911_),
    .A1(\clock_inst.hour_c[12] ),
    .A2(net451));
 sg13g2_inv_1 _08318_ (.Y(_00058_),
    .A(_00911_));
 sg13g2_nor3_1 _08319_ (.A(net506),
    .B(_00757_),
    .C(_00775_),
    .Y(_00912_));
 sg13g2_a21o_1 _08320_ (.A2(net361),
    .A1(\clock_inst.hour_c[13] ),
    .B1(_00912_),
    .X(_00059_));
 sg13g2_inv_1 _08321_ (.Y(_00913_),
    .A(\clock_inst.hour_c[14] ));
 sg13g2_a21oi_1 _08322_ (.A1(net510),
    .A2(_00899_),
    .Y(_00914_),
    .B1(_00789_));
 sg13g2_o21ai_1 _08323_ (.B1(_00802_),
    .Y(_00915_),
    .A1(net506),
    .A2(_00914_));
 sg13g2_a22oi_1 _08324_ (.Y(_00060_),
    .B1(_00915_),
    .B2(_00845_),
    .A2(net360),
    .A1(_00913_));
 sg13g2_a21oi_1 _08325_ (.A1(net509),
    .A2(_00744_),
    .Y(_00916_),
    .B1(_00729_));
 sg13g2_nand2_1 _08326_ (.Y(_00917_),
    .A(_00750_),
    .B(net359));
 sg13g2_o21ai_1 _08327_ (.B1(_00917_),
    .Y(_00918_),
    .A1(net545),
    .A2(_00916_));
 sg13g2_a22oi_1 _08328_ (.Y(_00919_),
    .B1(_00918_),
    .B2(net505),
    .A2(net365),
    .A1(\clock_inst.hour_c[15] ));
 sg13g2_inv_1 _08329_ (.Y(_00061_),
    .A(_00919_));
 sg13g2_o21ai_1 _08330_ (.B1(net514),
    .Y(_00920_),
    .A1(_00729_),
    .A2(_00795_));
 sg13g2_o21ai_1 _08331_ (.B1(_00920_),
    .Y(_00921_),
    .A1(\clock_inst.hour_c[16] ),
    .A2(net451));
 sg13g2_inv_1 _08332_ (.Y(_00062_),
    .A(_00921_));
 sg13g2_o21ai_1 _08333_ (.B1(net549),
    .Y(_00922_),
    .A1(_00729_),
    .A2(_00776_));
 sg13g2_o21ai_1 _08334_ (.B1(_00922_),
    .Y(_00923_),
    .A1(\clock_inst.hour_c[17] ),
    .A2(net451));
 sg13g2_inv_1 _08335_ (.Y(_00063_),
    .A(_00923_));
 sg13g2_nand2_1 _08336_ (.Y(_00924_),
    .A(net514),
    .B(_00854_));
 sg13g2_buf_8 _08337_ (.A(\clock_inst.hour_a[18] ),
    .X(_00925_));
 sg13g2_nand2_1 _08338_ (.Y(_00926_),
    .A(_00925_),
    .B(net361));
 sg13g2_o21ai_1 _08339_ (.B1(_00926_),
    .Y(_00064_),
    .A1(_00705_),
    .A2(_00924_));
 sg13g2_inv_1 _08340_ (.Y(_00927_),
    .A(\clock_inst.hour_c[19] ));
 sg13g2_a21oi_1 _08341_ (.A1(net510),
    .A2(_00900_),
    .Y(_00928_),
    .B1(_00783_));
 sg13g2_nand2_1 _08342_ (.Y(_00929_),
    .A(_00714_),
    .B(net359));
 sg13g2_o21ai_1 _08343_ (.B1(_00929_),
    .Y(_00930_),
    .A1(net506),
    .A2(_00928_));
 sg13g2_a22oi_1 _08344_ (.Y(_00065_),
    .B1(_00930_),
    .B2(_00845_),
    .A2(_00825_),
    .A1(_00927_));
 sg13g2_a21oi_1 _08345_ (.A1(_00695_),
    .A2(_00842_),
    .Y(_00931_),
    .B1(_00809_));
 sg13g2_nand2_1 _08346_ (.Y(_00932_),
    .A(\clock_inst.hour_c[1] ),
    .B(_00763_));
 sg13g2_o21ai_1 _08347_ (.B1(_00932_),
    .Y(_00066_),
    .A1(_00757_),
    .A2(_00931_));
 sg13g2_inv_1 _08348_ (.Y(_00933_),
    .A(\clock_inst.hour_c[21] ));
 sg13g2_nor2_1 _08349_ (.A(net547),
    .B(net515),
    .Y(_00934_));
 sg13g2_a21oi_1 _08350_ (.A1(net509),
    .A2(_00736_),
    .Y(_00935_),
    .B1(_00934_));
 sg13g2_and2_1 _08351_ (.A(_00766_),
    .B(_00935_),
    .X(_00936_));
 sg13g2_a22oi_1 _08352_ (.Y(_00067_),
    .B1(net362),
    .B2(_00936_),
    .A2(net360),
    .A1(_00933_));
 sg13g2_inv_1 _08353_ (.Y(_00937_),
    .A(\clock_inst.hour_c[23] ));
 sg13g2_a22oi_1 _08354_ (.Y(_00938_),
    .B1(_00729_),
    .B2(net549),
    .A2(_00937_),
    .A1(_00767_));
 sg13g2_inv_1 _08355_ (.Y(_00939_),
    .A(_00938_));
 sg13g2_nand3_1 _08356_ (.B(_00847_),
    .C(_00727_),
    .A(_00683_),
    .Y(_00940_));
 sg13g2_o21ai_1 _08357_ (.B1(_00940_),
    .Y(_00941_),
    .A1(net514),
    .A2(\clock_inst.hour_c[23] ));
 sg13g2_a21oi_1 _08358_ (.A1(net508),
    .A2(_00939_),
    .Y(_00068_),
    .B1(_00941_));
 sg13g2_inv_1 _08359_ (.Y(_00942_),
    .A(\clock_inst.hour_c[24] ));
 sg13g2_buf_1 _08360_ (.A(_00661_),
    .X(_00943_));
 sg13g2_o21ai_1 _08361_ (.B1(_00929_),
    .Y(_00944_),
    .A1(net506),
    .A2(_00867_));
 sg13g2_a22oi_1 _08362_ (.Y(_00069_),
    .B1(_00944_),
    .B2(net449),
    .A2(net358),
    .A1(_00942_));
 sg13g2_inv_1 _08363_ (.Y(_00945_),
    .A(\clock_inst.hour_c[25] ));
 sg13g2_o21ai_1 _08364_ (.B1(net512),
    .Y(_00946_),
    .A1(_00847_),
    .A2(_00764_));
 sg13g2_nand2_1 _08365_ (.Y(_00947_),
    .A(_00816_),
    .B(_00946_));
 sg13g2_a22oi_1 _08366_ (.Y(_00070_),
    .B1(_00947_),
    .B2(net449),
    .A2(net358),
    .A1(_00945_));
 sg13g2_a21oi_1 _08367_ (.A1(net508),
    .A2(\clock_inst.hour_c[26] ),
    .Y(_00948_),
    .B1(_00894_));
 sg13g2_a21o_1 _08368_ (.A2(\clock_inst.hour_c[26] ),
    .A1(net550),
    .B1(net362),
    .X(_00949_));
 sg13g2_a22oi_1 _08369_ (.Y(_00950_),
    .B1(_00949_),
    .B2(net503),
    .A2(\clock_inst.hour_c[26] ),
    .A1(_00748_));
 sg13g2_o21ai_1 _08370_ (.B1(_00950_),
    .Y(_00071_),
    .A1(net503),
    .A2(_00948_));
 sg13g2_a21o_1 _08371_ (.A2(_00934_),
    .A1(net510),
    .B1(net359),
    .X(_00951_));
 sg13g2_o21ai_1 _08372_ (.B1(_00754_),
    .Y(_00952_),
    .A1(_00680_),
    .A2(\clock_inst.hour_c[27] ));
 sg13g2_o21ai_1 _08373_ (.B1(net506),
    .Y(_00953_),
    .A1(_00837_),
    .A2(_00854_));
 sg13g2_a21oi_1 _08374_ (.A1(_00684_),
    .A2(_00953_),
    .Y(_00954_),
    .B1(\clock_inst.hour_c[27] ));
 sg13g2_a221oi_1 _08375_ (.B2(_00855_),
    .C1(_00954_),
    .B1(_00952_),
    .A1(net362),
    .Y(_00072_),
    .A2(_00951_));
 sg13g2_o21ai_1 _08376_ (.B1(_00766_),
    .Y(_00955_),
    .A1(_00742_),
    .A2(net359));
 sg13g2_nand2_1 _08377_ (.Y(_00956_),
    .A(net516),
    .B(_00836_));
 sg13g2_o21ai_1 _08378_ (.B1(_00956_),
    .Y(_00957_),
    .A1(net550),
    .A2(net359));
 sg13g2_a21oi_1 _08379_ (.A1(_00709_),
    .A2(_00957_),
    .Y(_00958_),
    .B1(\clock_inst.hour_c[28] ));
 sg13g2_a21oi_1 _08380_ (.A1(net507),
    .A2(_00955_),
    .Y(_00073_),
    .B1(_00958_));
 sg13g2_inv_1 _08381_ (.Y(_00959_),
    .A(\clock_inst.hour_c[29] ));
 sg13g2_a21o_1 _08382_ (.A2(_00801_),
    .A1(_00750_),
    .B1(_00905_),
    .X(_00960_));
 sg13g2_a22oi_1 _08383_ (.Y(_00074_),
    .B1(_00960_),
    .B2(net449),
    .A2(net358),
    .A1(_00959_));
 sg13g2_inv_1 _08384_ (.Y(_00961_),
    .A(\clock_inst.hour_c[30] ));
 sg13g2_nand2_1 _08385_ (.Y(_00962_),
    .A(net509),
    .B(_00847_));
 sg13g2_nand2_1 _08386_ (.Y(_00963_),
    .A(_00727_),
    .B(_00962_));
 sg13g2_a22oi_1 _08387_ (.Y(_00075_),
    .B1(_00963_),
    .B2(net507),
    .A2(net358),
    .A1(_00961_));
 sg13g2_buf_2 _08388_ (.A(\clock_inst.hour_a[4] ),
    .X(_00964_));
 sg13g2_nor2_1 _08389_ (.A(net503),
    .B(_00696_),
    .Y(_00965_));
 sg13g2_a21oi_1 _08390_ (.A1(net503),
    .A2(_00751_),
    .Y(_00966_),
    .B1(_00965_));
 sg13g2_a22oi_1 _08391_ (.Y(_00967_),
    .B1(_00966_),
    .B2(net511),
    .A2(net365),
    .A1(_00964_));
 sg13g2_inv_1 _08392_ (.Y(_00076_),
    .A(_00967_));
 sg13g2_inv_1 _08393_ (.Y(_00968_),
    .A(\clock_inst.hour_c[32] ));
 sg13g2_o21ai_1 _08394_ (.B1(net512),
    .Y(_00969_),
    .A1(net454),
    .A2(net515));
 sg13g2_a22oi_1 _08395_ (.Y(_00077_),
    .B1(net362),
    .B2(_00969_),
    .A2(net358),
    .A1(_00968_));
 sg13g2_a21o_1 _08396_ (.A2(_00757_),
    .A1(\clock_inst.hour_c[33] ),
    .B1(_00894_),
    .X(_00078_));
 sg13g2_nand2_1 _08397_ (.Y(_00970_),
    .A(\clock_inst.hour_c[0] ),
    .B(net361));
 sg13g2_o21ai_1 _08398_ (.B1(_00970_),
    .Y(_00079_),
    .A1(_00757_),
    .A2(_00935_));
 sg13g2_nand2_1 _08399_ (.Y(_00971_),
    .A(\clock_inst.hour_c[37] ),
    .B(_00763_));
 sg13g2_o21ai_1 _08400_ (.B1(_00971_),
    .Y(_00080_),
    .A1(_00733_),
    .A2(_00924_));
 sg13g2_a21o_1 _08401_ (.A2(_00707_),
    .A1(net504),
    .B1(_00669_),
    .X(_00972_));
 sg13g2_a22oi_1 _08402_ (.Y(_00973_),
    .B1(_00722_),
    .B2(_00972_),
    .A2(net365),
    .A1(\clock_inst.hour_c[2] ));
 sg13g2_inv_1 _08403_ (.Y(_00081_),
    .A(_00973_));
 sg13g2_inv_1 _08404_ (.Y(_00974_),
    .A(\clock_inst.hour_c[40] ));
 sg13g2_o21ai_1 _08405_ (.B1(_00940_),
    .Y(_00082_),
    .A1(_00974_),
    .A2(_00703_));
 sg13g2_o21ai_1 _08406_ (.B1(net510),
    .Y(_00975_),
    .A1(_00714_),
    .A2(_00706_));
 sg13g2_nand2b_1 _08407_ (.Y(_00976_),
    .B(_00975_),
    .A_N(_00734_));
 sg13g2_a22oi_1 _08408_ (.Y(_00977_),
    .B1(_00976_),
    .B2(net511),
    .A2(net365),
    .A1(\clock_inst.hour_c[41] ));
 sg13g2_inv_1 _08409_ (.Y(_00083_),
    .A(_00977_));
 sg13g2_inv_1 _08410_ (.Y(_00978_),
    .A(\clock_inst.hour_c[42] ));
 sg13g2_a21oi_1 _08411_ (.A1(_00735_),
    .A2(net364),
    .Y(_00979_),
    .B1(net454));
 sg13g2_or2_1 _08412_ (.X(_00980_),
    .B(_00979_),
    .A(_00729_));
 sg13g2_a22oi_1 _08413_ (.Y(_00084_),
    .B1(_00980_),
    .B2(net507),
    .A2(net358),
    .A1(_00978_));
 sg13g2_inv_1 _08414_ (.Y(_00981_),
    .A(\clock_inst.hour_c[43] ));
 sg13g2_o21ai_1 _08415_ (.B1(_00908_),
    .Y(_00982_),
    .A1(net509),
    .A2(_00705_));
 sg13g2_a21o_1 _08416_ (.A2(_00982_),
    .A1(_00675_),
    .B1(_00714_),
    .X(_00983_));
 sg13g2_a22oi_1 _08417_ (.Y(_00085_),
    .B1(_00983_),
    .B2(net507),
    .A2(_00754_),
    .A1(_00981_));
 sg13g2_inv_1 _08418_ (.Y(_00984_),
    .A(\clock_inst.hour_c[44] ));
 sg13g2_o21ai_1 _08419_ (.B1(net504),
    .Y(_00985_),
    .A1(_00750_),
    .A2(_00714_));
 sg13g2_nand2_1 _08420_ (.Y(_00986_),
    .A(_00794_),
    .B(_00985_));
 sg13g2_a22oi_1 _08421_ (.Y(_00086_),
    .B1(_00986_),
    .B2(net507),
    .A2(net358),
    .A1(_00984_));
 sg13g2_nand3_1 _08422_ (.B(_00678_),
    .C(net364),
    .A(_00668_),
    .Y(_00987_));
 sg13g2_nand2_1 _08423_ (.Y(_00988_),
    .A(_00736_),
    .B(_00987_));
 sg13g2_a22oi_1 _08424_ (.Y(_00989_),
    .B1(_00988_),
    .B2(net511),
    .A2(_00662_),
    .A1(\clock_inst.hour_c[45] ));
 sg13g2_inv_1 _08425_ (.Y(_00087_),
    .A(_00989_));
 sg13g2_nor2_1 _08426_ (.A(_00716_),
    .B(_00807_),
    .Y(_00990_));
 sg13g2_nand2_1 _08427_ (.Y(_00991_),
    .A(_00696_),
    .B(_00854_));
 sg13g2_o21ai_1 _08428_ (.B1(_00991_),
    .Y(_00992_),
    .A1(net510),
    .A2(_00990_));
 sg13g2_a22oi_1 _08429_ (.Y(_00993_),
    .B1(_00992_),
    .B2(net511),
    .A2(net365),
    .A1(\clock_inst.hour_c[46] ));
 sg13g2_inv_1 _08430_ (.Y(_00088_),
    .A(_00993_));
 sg13g2_inv_1 _08431_ (.Y(_00994_),
    .A(_00841_));
 sg13g2_nand2_1 _08432_ (.Y(_00995_),
    .A(_00683_),
    .B(net454));
 sg13g2_a21oi_1 _08433_ (.A1(net364),
    .A2(_00994_),
    .Y(_00996_),
    .B1(_00995_));
 sg13g2_a21o_1 _08434_ (.A2(net361),
    .A1(\clock_inst.hour_c[49] ),
    .B1(_00996_),
    .X(_00089_));
 sg13g2_a21oi_1 _08435_ (.A1(net512),
    .A2(_00750_),
    .Y(_00997_),
    .B1(_00815_));
 sg13g2_nand2_1 _08436_ (.Y(_00998_),
    .A(\clock_inst.hour_c[50] ),
    .B(net361));
 sg13g2_o21ai_1 _08437_ (.B1(_00998_),
    .Y(_00090_),
    .A1(_00995_),
    .A2(_00997_));
 sg13g2_inv_1 _08438_ (.Y(_00999_),
    .A(\clock_inst.hour_c[51] ));
 sg13g2_o21ai_1 _08439_ (.B1(_00877_),
    .Y(_01000_),
    .A1(_00669_),
    .A2(_00727_));
 sg13g2_a22oi_1 _08440_ (.Y(_00091_),
    .B1(_01000_),
    .B2(net507),
    .A2(_00943_),
    .A1(_00999_));
 sg13g2_inv_1 _08441_ (.Y(_01001_),
    .A(\clock_inst.hour_c[52] ));
 sg13g2_a22oi_1 _08442_ (.Y(_00092_),
    .B1(_00775_),
    .B2(_00856_),
    .A2(_00943_),
    .A1(_01001_));
 sg13g2_nor2b_1 _08443_ (.A(net359),
    .B_N(_00962_),
    .Y(_01002_));
 sg13g2_nand2_1 _08444_ (.Y(_01003_),
    .A(\clock_inst.hour_c[5] ),
    .B(net361));
 sg13g2_o21ai_1 _08445_ (.B1(_01003_),
    .Y(_00093_),
    .A1(_00754_),
    .A2(_01002_));
 sg13g2_inv_1 _08446_ (.Y(_01004_),
    .A(\clock_inst.hour_c[6] ));
 sg13g2_xnor2_1 _08447_ (.Y(_01005_),
    .A(_00790_),
    .B(_00885_));
 sg13g2_o21ai_1 _08448_ (.B1(_00794_),
    .Y(_01006_),
    .A1(net506),
    .A2(_01005_));
 sg13g2_a22oi_1 _08449_ (.Y(_00094_),
    .B1(_01006_),
    .B2(net507),
    .A2(net358),
    .A1(_01004_));
 sg13g2_inv_1 _08450_ (.Y(_01007_),
    .A(\clock_inst.hour_c[7] ));
 sg13g2_o21ai_1 _08451_ (.B1(net511),
    .Y(_01008_),
    .A1(_00841_),
    .A2(_00906_));
 sg13g2_o21ai_1 _08452_ (.B1(_01008_),
    .Y(_00095_),
    .A1(_01007_),
    .A2(net451));
 sg13g2_inv_1 _08453_ (.Y(_01009_),
    .A(\clock_inst.hour_c[8] ));
 sg13g2_o21ai_1 _08454_ (.B1(_00719_),
    .Y(_01010_),
    .A1(_00695_),
    .A2(_00699_));
 sg13g2_a22oi_1 _08455_ (.Y(_00096_),
    .B1(_01010_),
    .B2(_00746_),
    .A2(net361),
    .A1(_01009_));
 sg13g2_inv_1 _08456_ (.Y(_01011_),
    .A(\clock_inst.hour_c[9] ));
 sg13g2_o21ai_1 _08457_ (.B1(net511),
    .Y(_01012_),
    .A1(_00807_),
    .A2(_00795_));
 sg13g2_o21ai_1 _08458_ (.B1(_01012_),
    .Y(_00097_),
    .A1(_01011_),
    .A2(net451));
 sg13g2_buf_2 _08459_ (.A(\clock_inst.hour_tile.e0[0] ),
    .X(_01013_));
 sg13g2_buf_1 _08460_ (.A(\clock_inst.vga_inst.vga_x[3] ),
    .X(_01014_));
 sg13g2_buf_2 _08461_ (.A(\clock_inst.vga_inst.vga_x[7] ),
    .X(_01015_));
 sg13g2_nor2_1 _08462_ (.A(_01014_),
    .B(_01015_),
    .Y(_01016_));
 sg13g2_buf_2 _08463_ (.A(\clock_inst.vga_inst.vga_x[1] ),
    .X(_01017_));
 sg13g2_buf_2 _08464_ (.A(\clock_inst.vga_inst.vga_x[0] ),
    .X(_01018_));
 sg13g2_buf_1 _08465_ (.A(\clock_inst.vga_inst.vga_x[2] ),
    .X(_01019_));
 sg13g2_nor3_1 _08466_ (.A(_01017_),
    .B(_01018_),
    .C(_01019_),
    .Y(_01020_));
 sg13g2_nand2_2 _08467_ (.Y(_01021_),
    .A(_01016_),
    .B(_01020_));
 sg13g2_inv_1 _08468_ (.Y(_01022_),
    .A(\clock_inst.vga_inst.vga_x[4] ));
 sg13g2_buf_2 _08469_ (.A(\clock_inst.vga_inst.vga_x[8] ),
    .X(_01023_));
 sg13g2_buf_2 _08470_ (.A(\clock_inst.vga_inst.vga_x[9] ),
    .X(_01024_));
 sg13g2_nand3_1 _08471_ (.B(_01023_),
    .C(_01024_),
    .A(_01022_),
    .Y(_01025_));
 sg13g2_buf_1 _08472_ (.A(_01025_),
    .X(_01026_));
 sg13g2_buf_1 _08473_ (.A(\clock_inst.vga_inst.vga_x[6] ),
    .X(_01027_));
 sg13g2_buf_2 _08474_ (.A(\clock_inst.vga_inst.vga_x[5] ),
    .X(_01028_));
 sg13g2_nand2b_1 _08475_ (.Y(_01029_),
    .B(_01028_),
    .A_N(net574));
 sg13g2_or3_1 _08476_ (.A(_01021_),
    .B(_01026_),
    .C(_01029_),
    .X(_01030_));
 sg13g2_buf_2 _08477_ (.A(_01030_),
    .X(_01031_));
 sg13g2_buf_1 _08478_ (.A(_01031_),
    .X(_01032_));
 sg13g2_buf_1 _08479_ (.A(net244),
    .X(_01033_));
 sg13g2_buf_1 _08480_ (.A(_01033_),
    .X(_01034_));
 sg13g2_xnor2_1 _08481_ (.Y(_01035_),
    .A(_00823_),
    .B(_01013_));
 sg13g2_buf_1 _08482_ (.A(\clock_inst.vga_inst.vga_y[4] ),
    .X(_01036_));
 sg13g2_buf_1 _08483_ (.A(\clock_inst.vga_inst.vga_y[5] ),
    .X(_01037_));
 sg13g2_buf_1 _08484_ (.A(_01037_),
    .X(_01038_));
 sg13g2_buf_2 _08485_ (.A(\clock_inst.vga_inst.vga_y[9] ),
    .X(_01039_));
 sg13g2_buf_2 _08486_ (.A(\clock_inst.vga_inst.vga_y[6] ),
    .X(_01040_));
 sg13g2_buf_1 _08487_ (.A(\clock_inst.vga_inst.vga_y[7] ),
    .X(_01041_));
 sg13g2_buf_2 _08488_ (.A(\clock_inst.vga_inst.vga_y[8] ),
    .X(_01042_));
 sg13g2_nand3_1 _08489_ (.B(_01041_),
    .C(_01042_),
    .A(_01040_),
    .Y(_01043_));
 sg13g2_nor2_1 _08490_ (.A(_01039_),
    .B(_01043_),
    .Y(_01044_));
 sg13g2_buf_1 _08491_ (.A(\clock_inst.vga_inst.vga_y[1] ),
    .X(_01045_));
 sg13g2_nand2_2 _08492_ (.Y(_01046_),
    .A(_01045_),
    .B(\clock_inst.vga_inst.vga_y[0] ));
 sg13g2_buf_1 _08493_ (.A(\clock_inst.vga_inst.vga_y[3] ),
    .X(_01047_));
 sg13g2_buf_2 _08494_ (.A(\clock_inst.vga_inst.vga_y[2] ),
    .X(_01048_));
 sg13g2_nor2_1 _08495_ (.A(_01047_),
    .B(_01048_),
    .Y(_01049_));
 sg13g2_nor2b_1 _08496_ (.A(_01046_),
    .B_N(_01049_),
    .Y(_01050_));
 sg13g2_nand4_1 _08497_ (.B(net543),
    .C(_01044_),
    .A(net573),
    .Y(_01051_),
    .D(_01050_));
 sg13g2_buf_1 _08498_ (.A(_01051_),
    .X(_01052_));
 sg13g2_nand4_1 _08499_ (.B(_01037_),
    .C(_01044_),
    .A(_01036_),
    .Y(_01053_),
    .D(_01050_));
 sg13g2_buf_1 _08500_ (.A(_01053_),
    .X(_01054_));
 sg13g2_buf_1 _08501_ (.A(_01054_),
    .X(_01055_));
 sg13g2_nor3_1 _08502_ (.A(_01021_),
    .B(_01026_),
    .C(_01029_),
    .Y(_01056_));
 sg13g2_buf_2 _08503_ (.A(_01056_),
    .X(_01057_));
 sg13g2_o21ai_1 _08504_ (.B1(_01057_),
    .Y(_01058_),
    .A1(\clock_inst.hour_c[0] ),
    .A2(net243));
 sg13g2_a21oi_1 _08505_ (.A1(_01035_),
    .A2(_01052_),
    .Y(_01059_),
    .B1(_01058_));
 sg13g2_a21o_1 _08506_ (.A2(net112),
    .A1(_01013_),
    .B1(_01059_),
    .X(_00098_));
 sg13g2_inv_1 _08507_ (.Y(_01060_),
    .A(\clock_inst.hour_tile.e0[10] ));
 sg13g2_buf_1 _08508_ (.A(net244),
    .X(_01061_));
 sg13g2_buf_1 _08509_ (.A(net161),
    .X(_01062_));
 sg13g2_buf_1 _08510_ (.A(_01031_),
    .X(_01063_));
 sg13g2_buf_1 _08511_ (.A(net242),
    .X(_01064_));
 sg13g2_nand2_1 _08512_ (.Y(_01065_),
    .A(net573),
    .B(_01037_));
 sg13g2_or2_1 _08513_ (.X(_01066_),
    .B(_01043_),
    .A(_01039_));
 sg13g2_buf_2 _08514_ (.A(_01066_),
    .X(_01067_));
 sg13g2_nand2b_1 _08515_ (.Y(_01068_),
    .B(_01049_),
    .A_N(_01046_));
 sg13g2_nor3_1 _08516_ (.A(_01065_),
    .B(_01067_),
    .C(_01068_),
    .Y(_01069_));
 sg13g2_buf_1 _08517_ (.A(_01069_),
    .X(_01070_));
 sg13g2_buf_1 _08518_ (.A(net241),
    .X(_01071_));
 sg13g2_buf_1 _08519_ (.A(net159),
    .X(_01072_));
 sg13g2_buf_2 _08520_ (.A(\clock_inst.hour_tile.e0[8] ),
    .X(_01073_));
 sg13g2_inv_1 _08521_ (.Y(_01074_),
    .A(_01073_));
 sg13g2_buf_1 _08522_ (.A(\clock_inst.hour_tile.e0[6] ),
    .X(_01075_));
 sg13g2_inv_1 _08523_ (.Y(_01076_),
    .A(\clock_inst.hour_tile.e0[7] ));
 sg13g2_nor2_2 _08524_ (.A(_00725_),
    .B(_01076_),
    .Y(_01077_));
 sg13g2_buf_1 _08525_ (.A(\clock_inst.hour_tile.e0[3] ),
    .X(_01078_));
 sg13g2_inv_1 _08526_ (.Y(_01079_),
    .A(_01078_));
 sg13g2_buf_1 _08527_ (.A(\clock_inst.hour_tile.e0[2] ),
    .X(_01080_));
 sg13g2_nand2_1 _08528_ (.Y(_01081_),
    .A(_00852_),
    .B(_01080_));
 sg13g2_nor2_1 _08529_ (.A(_00852_),
    .B(_01080_),
    .Y(_01082_));
 sg13g2_buf_2 _08530_ (.A(\clock_inst.hour_tile.e0[1] ),
    .X(_01083_));
 sg13g2_nor2_1 _08531_ (.A(_00835_),
    .B(_01083_),
    .Y(_01084_));
 sg13g2_a22oi_1 _08532_ (.Y(_01085_),
    .B1(_00835_),
    .B2(_01083_),
    .A2(_01013_),
    .A1(_00823_));
 sg13g2_or3_1 _08533_ (.A(_01082_),
    .B(_01084_),
    .C(_01085_),
    .X(_01086_));
 sg13g2_xnor2_1 _08534_ (.Y(_01087_),
    .A(\clock_inst.hour_b[5] ),
    .B(\clock_inst.hour_tile.e0[5] ));
 sg13g2_buf_2 _08535_ (.A(\clock_inst.hour_tile.e0[4] ),
    .X(_01088_));
 sg13g2_xor2_1 _08536_ (.B(_01088_),
    .A(_00889_),
    .X(_01089_));
 sg13g2_nand2b_1 _08537_ (.Y(_01090_),
    .B(_01089_),
    .A_N(_01087_));
 sg13g2_a221oi_1 _08538_ (.B2(_01086_),
    .C1(_01090_),
    .B1(_01081_),
    .A1(_00828_),
    .Y(_01091_),
    .A2(_01079_));
 sg13g2_buf_2 _08539_ (.A(_01091_),
    .X(_01092_));
 sg13g2_nand2_1 _08540_ (.Y(_01093_),
    .A(net577),
    .B(_01078_));
 sg13g2_inv_1 _08541_ (.Y(_01094_),
    .A(\clock_inst.hour_tile.e0[5] ));
 sg13g2_a22oi_1 _08542_ (.Y(_01095_),
    .B1(\clock_inst.hour_b[5] ),
    .B2(\clock_inst.hour_tile.e0[5] ),
    .A2(_01088_),
    .A1(_00889_));
 sg13g2_a21o_1 _08543_ (.A2(_01094_),
    .A1(_00893_),
    .B1(_01095_),
    .X(_01096_));
 sg13g2_o21ai_1 _08544_ (.B1(_01096_),
    .Y(_01097_),
    .A1(_01090_),
    .A2(_01093_));
 sg13g2_buf_2 _08545_ (.A(_01097_),
    .X(_01098_));
 sg13g2_nor4_2 _08546_ (.A(_01075_),
    .B(_01077_),
    .C(_01092_),
    .Y(_01099_),
    .D(_01098_));
 sg13g2_nor4_2 _08547_ (.A(net546),
    .B(_01077_),
    .C(_01092_),
    .Y(_01100_),
    .D(_01098_));
 sg13g2_nand2_1 _08548_ (.Y(_01101_),
    .A(_00725_),
    .B(_01076_));
 sg13g2_nor2_1 _08549_ (.A(_00731_),
    .B(_01075_),
    .Y(_01102_));
 sg13g2_o21ai_1 _08550_ (.B1(_01102_),
    .Y(_01103_),
    .A1(_00725_),
    .A2(_01076_));
 sg13g2_nand2_1 _08551_ (.Y(_01104_),
    .A(_01101_),
    .B(_01103_));
 sg13g2_nor4_2 _08552_ (.A(_01074_),
    .B(_01099_),
    .C(_01100_),
    .Y(_01105_),
    .D(_01104_));
 sg13g2_buf_1 _08553_ (.A(\clock_inst.hour_tile.e0[9] ),
    .X(_01106_));
 sg13g2_nor2b_1 _08554_ (.A(net577),
    .B_N(_01106_),
    .Y(_01107_));
 sg13g2_inv_1 _08555_ (.Y(_01108_),
    .A(_01075_));
 sg13g2_nand2_1 _08556_ (.Y(_01109_),
    .A(_01108_),
    .B(_01074_));
 sg13g2_nor4_1 _08557_ (.A(_01077_),
    .B(_01092_),
    .C(_01098_),
    .D(_01109_),
    .Y(_01110_));
 sg13g2_or2_1 _08558_ (.X(_01111_),
    .B(_01073_),
    .A(net546));
 sg13g2_nor4_1 _08559_ (.A(_01077_),
    .B(_01092_),
    .C(_01098_),
    .D(_01111_),
    .Y(_01112_));
 sg13g2_a21oi_1 _08560_ (.A1(_01101_),
    .A2(_01103_),
    .Y(_01113_),
    .B1(_01073_));
 sg13g2_or3_1 _08561_ (.A(_01110_),
    .B(_01112_),
    .C(_01113_),
    .X(_01114_));
 sg13g2_buf_2 _08562_ (.A(_01114_),
    .X(_01115_));
 sg13g2_nor2b_1 _08563_ (.A(_01106_),
    .B_N(net577),
    .Y(_01116_));
 sg13g2_a22oi_1 _08564_ (.Y(_01117_),
    .B1(_01115_),
    .B2(_01116_),
    .A2(_01107_),
    .A1(_01105_));
 sg13g2_xnor2_1 _08565_ (.Y(_01118_),
    .A(_01060_),
    .B(_01117_));
 sg13g2_buf_1 _08566_ (.A(net241),
    .X(_01119_));
 sg13g2_buf_1 _08567_ (.A(net158),
    .X(_01120_));
 sg13g2_nand2_1 _08568_ (.Y(_01121_),
    .A(\clock_inst.hour_c[10] ),
    .B(_01120_));
 sg13g2_o21ai_1 _08569_ (.B1(_01121_),
    .Y(_01122_),
    .A1(net110),
    .A2(_01118_));
 sg13g2_nor2_1 _08570_ (.A(net160),
    .B(_01122_),
    .Y(_01123_));
 sg13g2_a21oi_1 _08571_ (.A1(_01060_),
    .A2(net111),
    .Y(_00099_),
    .B1(_01123_));
 sg13g2_inv_1 _08572_ (.Y(_01124_),
    .A(\clock_inst.hour_tile.e0[11] ));
 sg13g2_and2_1 _08573_ (.A(_01060_),
    .B(_01116_),
    .X(_01125_));
 sg13g2_and4_1 _08574_ (.A(_00828_),
    .B(_01073_),
    .C(_01106_),
    .D(\clock_inst.hour_tile.e0[10] ),
    .X(_01126_));
 sg13g2_nor3_2 _08575_ (.A(_01099_),
    .B(_01100_),
    .C(_01104_),
    .Y(_01127_));
 sg13g2_a22oi_1 _08576_ (.Y(_01128_),
    .B1(_01126_),
    .B2(_01127_),
    .A2(_01125_),
    .A1(_01115_));
 sg13g2_xnor2_1 _08577_ (.Y(_01129_),
    .A(\clock_inst.hour_tile.e0[11] ),
    .B(_01128_));
 sg13g2_buf_1 _08578_ (.A(net243),
    .X(_01130_));
 sg13g2_mux2_1 _08579_ (.A0(\clock_inst.hour_c[11] ),
    .A1(_01129_),
    .S(net157),
    .X(_01131_));
 sg13g2_nor2_1 _08580_ (.A(net160),
    .B(_01131_),
    .Y(_01132_));
 sg13g2_a21oi_1 _08581_ (.A1(_01124_),
    .A2(net111),
    .Y(_00100_),
    .B1(_01132_));
 sg13g2_buf_1 _08582_ (.A(\clock_inst.hour_tile.e0[12] ),
    .X(_01133_));
 sg13g2_inv_1 _08583_ (.Y(_01134_),
    .A(_01133_));
 sg13g2_buf_1 _08584_ (.A(_01057_),
    .X(_01135_));
 sg13g2_buf_1 _08585_ (.A(_01135_),
    .X(_01136_));
 sg13g2_buf_2 _08586_ (.A(_01136_),
    .X(_01137_));
 sg13g2_buf_1 _08587_ (.A(net240),
    .X(_01138_));
 sg13g2_and3_1 _08588_ (.X(_01139_),
    .A(\clock_inst.hour_tile.e0[10] ),
    .B(\clock_inst.hour_tile.e0[11] ),
    .C(_01107_));
 sg13g2_buf_1 _08589_ (.A(_01139_),
    .X(_01140_));
 sg13g2_nand3_1 _08590_ (.B(_01124_),
    .C(_01116_),
    .A(_01060_),
    .Y(_01141_));
 sg13g2_inv_1 _08591_ (.Y(_01142_),
    .A(_01141_));
 sg13g2_a22oi_1 _08592_ (.Y(_01143_),
    .B1(_01142_),
    .B2(_01115_),
    .A2(_01140_),
    .A1(_01105_));
 sg13g2_xnor2_1 _08593_ (.Y(_01144_),
    .A(_01134_),
    .B(_01143_));
 sg13g2_nor3_2 _08594_ (.A(_01065_),
    .B(_01067_),
    .C(_01068_),
    .Y(_01145_));
 sg13g2_nand2_1 _08595_ (.Y(_01146_),
    .A(\clock_inst.hour_c[12] ),
    .B(_01145_));
 sg13g2_o21ai_1 _08596_ (.B1(_01146_),
    .Y(_01147_),
    .A1(net110),
    .A2(_01144_));
 sg13g2_nand2_1 _08597_ (.Y(_01148_),
    .A(_01138_),
    .B(_01147_));
 sg13g2_o21ai_1 _08598_ (.B1(_01148_),
    .Y(_00101_),
    .A1(_01134_),
    .A2(_01137_));
 sg13g2_buf_1 _08599_ (.A(\clock_inst.hour_tile.e0[13] ),
    .X(_01149_));
 sg13g2_inv_1 _08600_ (.Y(_01150_),
    .A(_01149_));
 sg13g2_buf_2 _08601_ (.A(_01031_),
    .X(_01151_));
 sg13g2_buf_1 _08602_ (.A(net239),
    .X(_01152_));
 sg13g2_nor2_1 _08603_ (.A(_01150_),
    .B(_01119_),
    .Y(_01153_));
 sg13g2_nor2_1 _08604_ (.A(_01149_),
    .B(_01119_),
    .Y(_01154_));
 sg13g2_nand2_1 _08605_ (.Y(_01155_),
    .A(_01133_),
    .B(_01140_));
 sg13g2_nor3_1 _08606_ (.A(_01110_),
    .B(_01112_),
    .C(_01113_),
    .Y(_01156_));
 sg13g2_o21ai_1 _08607_ (.B1(_01156_),
    .Y(_01157_),
    .A1(net577),
    .A2(_01105_));
 sg13g2_buf_2 _08608_ (.A(_01157_),
    .X(_01158_));
 sg13g2_nand3_1 _08609_ (.B(_01115_),
    .C(_01142_),
    .A(_01134_),
    .Y(_01159_));
 sg13g2_o21ai_1 _08610_ (.B1(_01159_),
    .Y(_01160_),
    .A1(_01155_),
    .A2(_01158_));
 sg13g2_mux2_1 _08611_ (.A0(_01153_),
    .A1(_01154_),
    .S(_01160_),
    .X(_01161_));
 sg13g2_buf_1 _08612_ (.A(net158),
    .X(_01162_));
 sg13g2_and2_1 _08613_ (.A(\clock_inst.hour_c[13] ),
    .B(_01162_),
    .X(_01163_));
 sg13g2_nor3_1 _08614_ (.A(net154),
    .B(_01161_),
    .C(_01163_),
    .Y(_01164_));
 sg13g2_a21oi_1 _08615_ (.A1(_01150_),
    .A2(net111),
    .Y(_00102_),
    .B1(_01164_));
 sg13g2_inv_1 _08616_ (.Y(_01165_),
    .A(\clock_inst.hour_tile.e0[14] ));
 sg13g2_buf_2 _08617_ (.A(net156),
    .X(_01166_));
 sg13g2_o21ai_1 _08618_ (.B1(_01149_),
    .Y(_01167_),
    .A1(net577),
    .A2(_01073_));
 sg13g2_nor2_1 _08619_ (.A(_01155_),
    .B(_01167_),
    .Y(_01168_));
 sg13g2_nor3_1 _08620_ (.A(_01133_),
    .B(_01149_),
    .C(_01141_),
    .Y(_01169_));
 sg13g2_a22oi_1 _08621_ (.Y(_01170_),
    .B1(_01169_),
    .B2(_01115_),
    .A2(_01168_),
    .A1(_01127_));
 sg13g2_xnor2_1 _08622_ (.Y(_01171_),
    .A(_01165_),
    .B(_01170_));
 sg13g2_nand2_1 _08623_ (.Y(_01172_),
    .A(\clock_inst.hour_c[14] ),
    .B(_01120_));
 sg13g2_o21ai_1 _08624_ (.B1(_01172_),
    .Y(_01173_),
    .A1(net110),
    .A2(_01171_));
 sg13g2_nand2_1 _08625_ (.Y(_01174_),
    .A(net155),
    .B(_01173_));
 sg13g2_o21ai_1 _08626_ (.B1(_01174_),
    .Y(_00103_),
    .A1(_01165_),
    .A2(net106));
 sg13g2_inv_1 _08627_ (.Y(_01175_),
    .A(\clock_inst.hour_tile.e0[15] ));
 sg13g2_buf_1 _08628_ (.A(_01151_),
    .X(_01176_));
 sg13g2_buf_1 _08629_ (.A(net153),
    .X(_01177_));
 sg13g2_buf_1 _08630_ (.A(_01052_),
    .X(_01178_));
 sg13g2_buf_1 _08631_ (.A(_01178_),
    .X(_01179_));
 sg13g2_nor3_1 _08632_ (.A(_01150_),
    .B(_01165_),
    .C(_01155_),
    .Y(_01180_));
 sg13g2_and2_1 _08633_ (.A(_01165_),
    .B(_01169_),
    .X(_01181_));
 sg13g2_buf_1 _08634_ (.A(_01181_),
    .X(_01182_));
 sg13g2_mux2_1 _08635_ (.A0(_01180_),
    .A1(_01182_),
    .S(_01158_),
    .X(_01183_));
 sg13g2_xnor2_1 _08636_ (.Y(_01184_),
    .A(_01175_),
    .B(_01183_));
 sg13g2_nand2_1 _08637_ (.Y(_01185_),
    .A(_01179_),
    .B(_01184_));
 sg13g2_buf_2 _08638_ (.A(net109),
    .X(_01186_));
 sg13g2_a21oi_1 _08639_ (.A1(\clock_inst.hour_c[15] ),
    .A2(_01186_),
    .Y(_01187_),
    .B1(net162));
 sg13g2_a22oi_1 _08640_ (.Y(_00104_),
    .B1(_01185_),
    .B2(_01187_),
    .A2(_01177_),
    .A1(_01175_));
 sg13g2_inv_1 _08641_ (.Y(_01188_),
    .A(\clock_inst.hour_tile.e0[16] ));
 sg13g2_nand3_1 _08642_ (.B(_01175_),
    .C(_01182_),
    .A(_01074_),
    .Y(_01189_));
 sg13g2_nor2_1 _08643_ (.A(net577),
    .B(_01175_),
    .Y(_01190_));
 sg13g2_nand4_1 _08644_ (.B(_01149_),
    .C(\clock_inst.hour_tile.e0[14] ),
    .A(_01133_),
    .Y(_01191_),
    .D(_01190_));
 sg13g2_nor2_1 _08645_ (.A(_01073_),
    .B(_01141_),
    .Y(_01192_));
 sg13g2_a21oi_1 _08646_ (.A1(_01073_),
    .A2(_01140_),
    .Y(_01193_),
    .B1(_01192_));
 sg13g2_nor4_1 _08647_ (.A(_01099_),
    .B(_01100_),
    .C(_01104_),
    .D(_01193_),
    .Y(_01194_));
 sg13g2_mux2_1 _08648_ (.A0(_01189_),
    .A1(_01191_),
    .S(_01194_),
    .X(_01195_));
 sg13g2_xnor2_1 _08649_ (.Y(_01196_),
    .A(_01188_),
    .B(_01195_));
 sg13g2_nand2_1 _08650_ (.Y(_01197_),
    .A(\clock_inst.hour_c[16] ),
    .B(net109));
 sg13g2_o21ai_1 _08651_ (.B1(_01197_),
    .Y(_01198_),
    .A1(net110),
    .A2(_01196_));
 sg13g2_nor2_1 _08652_ (.A(net160),
    .B(_01198_),
    .Y(_01199_));
 sg13g2_a21oi_1 _08653_ (.A1(_01188_),
    .A2(_01062_),
    .Y(_00105_),
    .B1(_01199_));
 sg13g2_inv_1 _08654_ (.Y(_01200_),
    .A(\clock_inst.hour_tile.e0[17] ));
 sg13g2_buf_1 _08655_ (.A(net243),
    .X(_01201_));
 sg13g2_buf_1 _08656_ (.A(net151),
    .X(_01202_));
 sg13g2_buf_2 _08657_ (.A(_01202_),
    .X(_01203_));
 sg13g2_and3_1 _08658_ (.X(_01204_),
    .A(\clock_inst.hour_tile.e0[16] ),
    .B(_01180_),
    .C(_01190_));
 sg13g2_nand2_1 _08659_ (.Y(_01205_),
    .A(_01175_),
    .B(_01182_));
 sg13g2_nor2_1 _08660_ (.A(\clock_inst.hour_tile.e0[16] ),
    .B(_01205_),
    .Y(_01206_));
 sg13g2_a22oi_1 _08661_ (.Y(_01207_),
    .B1(_01206_),
    .B2(_01158_),
    .A2(_01204_),
    .A1(_01105_));
 sg13g2_xnor2_1 _08662_ (.Y(_01208_),
    .A(\clock_inst.hour_tile.e0[17] ),
    .B(_01207_));
 sg13g2_nand2_1 _08663_ (.Y(_01209_),
    .A(_01203_),
    .B(_01208_));
 sg13g2_buf_1 _08664_ (.A(_01145_),
    .X(_01210_));
 sg13g2_a21oi_1 _08665_ (.A1(\clock_inst.hour_c[17] ),
    .A2(_01210_),
    .Y(_01211_),
    .B1(net162));
 sg13g2_a22oi_1 _08666_ (.Y(_00106_),
    .B1(_01209_),
    .B2(_01211_),
    .A2(net105),
    .A1(_01200_));
 sg13g2_buf_2 _08667_ (.A(net156),
    .X(_01212_));
 sg13g2_buf_1 _08668_ (.A(net104),
    .X(_01213_));
 sg13g2_buf_2 _08669_ (.A(\clock_inst.hour_tile.e0[18] ),
    .X(_01214_));
 sg13g2_buf_1 _08670_ (.A(net243),
    .X(_01215_));
 sg13g2_buf_1 _08671_ (.A(net150),
    .X(_01216_));
 sg13g2_nand3_1 _08672_ (.B(net575),
    .C(_01216_),
    .A(_01214_),
    .Y(_01217_));
 sg13g2_o21ai_1 _08673_ (.B1(_01217_),
    .Y(_01218_),
    .A1(net575),
    .A2(net50));
 sg13g2_a21oi_1 _08674_ (.A1(net575),
    .A2(net155),
    .Y(_01219_),
    .B1(_01214_));
 sg13g2_a21oi_1 _08675_ (.A1(net103),
    .A2(_01218_),
    .Y(_00107_),
    .B1(_01219_));
 sg13g2_buf_2 _08676_ (.A(\clock_inst.hour_tile.e0[19] ),
    .X(_01220_));
 sg13g2_inv_1 _08677_ (.Y(_01221_),
    .A(_01220_));
 sg13g2_buf_1 _08678_ (.A(net151),
    .X(_01222_));
 sg13g2_nand2_1 _08679_ (.Y(_01223_),
    .A(_01214_),
    .B(net575));
 sg13g2_xor2_1 _08680_ (.B(_01220_),
    .A(_00831_),
    .X(_01224_));
 sg13g2_xnor2_1 _08681_ (.Y(_01225_),
    .A(_01223_),
    .B(_01224_));
 sg13g2_nand2_1 _08682_ (.Y(_01226_),
    .A(_01130_),
    .B(_01225_));
 sg13g2_o21ai_1 _08683_ (.B1(_01226_),
    .Y(_01227_),
    .A1(_00927_),
    .A2(net101));
 sg13g2_nor2_1 _08684_ (.A(net160),
    .B(_01227_),
    .Y(_01228_));
 sg13g2_a21oi_1 _08685_ (.A1(_01221_),
    .A2(net111),
    .Y(_00108_),
    .B1(_01228_));
 sg13g2_inv_1 _08686_ (.Y(_01229_),
    .A(_01083_));
 sg13g2_buf_1 _08687_ (.A(net161),
    .X(_01230_));
 sg13g2_nand2_1 _08688_ (.Y(_01231_),
    .A(_00823_),
    .B(_01013_));
 sg13g2_xnor2_1 _08689_ (.Y(_01232_),
    .A(_00835_),
    .B(_01083_));
 sg13g2_xnor2_1 _08690_ (.Y(_01233_),
    .A(_01231_),
    .B(_01232_));
 sg13g2_nand2_1 _08691_ (.Y(_01234_),
    .A(\clock_inst.hour_c[1] ),
    .B(net109));
 sg13g2_o21ai_1 _08692_ (.B1(_01234_),
    .Y(_01235_),
    .A1(net110),
    .A2(_01233_));
 sg13g2_nor2_1 _08693_ (.A(net160),
    .B(_01235_),
    .Y(_01236_));
 sg13g2_a21oi_1 _08694_ (.A1(_01229_),
    .A2(_01230_),
    .Y(_00109_),
    .B1(_01236_));
 sg13g2_buf_1 _08695_ (.A(\clock_inst.hour_tile.e0[20] ),
    .X(_01237_));
 sg13g2_nor2_1 _08696_ (.A(_01031_),
    .B(net241),
    .Y(_01238_));
 sg13g2_buf_1 _08697_ (.A(_01238_),
    .X(_01239_));
 sg13g2_buf_1 _08698_ (.A(net99),
    .X(_01240_));
 sg13g2_buf_1 _08699_ (.A(net49),
    .X(_01241_));
 sg13g2_a22oi_1 _08700_ (.Y(_01242_),
    .B1(_01214_),
    .B2(net575),
    .A2(_01220_),
    .A1(_00831_));
 sg13g2_nor2_1 _08701_ (.A(_00831_),
    .B(_01220_),
    .Y(_01243_));
 sg13g2_nor2_1 _08702_ (.A(_01242_),
    .B(_01243_),
    .Y(_01244_));
 sg13g2_xnor2_1 _08703_ (.Y(_01245_),
    .A(_00840_),
    .B(_01244_));
 sg13g2_nand2_1 _08704_ (.Y(_01246_),
    .A(_01241_),
    .B(_01245_));
 sg13g2_buf_1 _08705_ (.A(net159),
    .X(_01247_));
 sg13g2_buf_1 _08706_ (.A(_01057_),
    .X(_01248_));
 sg13g2_o21ai_1 _08707_ (.B1(net236),
    .Y(_01249_),
    .A1(_01247_),
    .A2(_01245_));
 sg13g2_nand2_1 _08708_ (.Y(_01250_),
    .A(_01237_),
    .B(_01249_));
 sg13g2_o21ai_1 _08709_ (.B1(_01250_),
    .Y(_00110_),
    .A1(_01237_),
    .A2(_01246_));
 sg13g2_inv_1 _08710_ (.Y(_01251_),
    .A(\clock_inst.hour_tile.e0[21] ));
 sg13g2_buf_1 _08711_ (.A(net159),
    .X(_01252_));
 sg13g2_nand2_1 _08712_ (.Y(_01253_),
    .A(\clock_inst.hour_c[21] ),
    .B(_01252_));
 sg13g2_and2_1 _08713_ (.A(\clock_inst.hour_b[20] ),
    .B(_01237_),
    .X(_01254_));
 sg13g2_nor2_1 _08714_ (.A(\clock_inst.hour_b[20] ),
    .B(_01237_),
    .Y(_01255_));
 sg13g2_nor3_1 _08715_ (.A(_01242_),
    .B(_01243_),
    .C(_01255_),
    .Y(_01256_));
 sg13g2_nor2_1 _08716_ (.A(_01254_),
    .B(_01256_),
    .Y(_01257_));
 sg13g2_xor2_1 _08717_ (.B(\clock_inst.hour_tile.e0[21] ),
    .A(net544),
    .X(_01258_));
 sg13g2_xnor2_1 _08718_ (.Y(_01259_),
    .A(_01257_),
    .B(_01258_));
 sg13g2_nand2_1 _08719_ (.Y(_01260_),
    .A(_01222_),
    .B(_01259_));
 sg13g2_and3_1 _08720_ (.X(_01261_),
    .A(net236),
    .B(_01253_),
    .C(_01260_));
 sg13g2_a21oi_1 _08721_ (.A1(_01251_),
    .A2(net100),
    .Y(_00111_),
    .B1(_01261_));
 sg13g2_buf_2 _08722_ (.A(\clock_inst.hour_tile.e0[22] ),
    .X(_01262_));
 sg13g2_buf_2 _08723_ (.A(net159),
    .X(_01263_));
 sg13g2_nor2_1 _08724_ (.A(net576),
    .B(\clock_inst.hour_tile.e0[21] ),
    .Y(_01264_));
 sg13g2_inv_1 _08725_ (.Y(_01265_),
    .A(_01264_));
 sg13g2_inv_1 _08726_ (.Y(_01266_),
    .A(net576));
 sg13g2_nor2_1 _08727_ (.A(_01266_),
    .B(_01251_),
    .Y(_01267_));
 sg13g2_or3_1 _08728_ (.A(_01254_),
    .B(_01256_),
    .C(_01267_),
    .X(_01268_));
 sg13g2_and2_1 _08729_ (.A(_01265_),
    .B(_01268_),
    .X(_01269_));
 sg13g2_buf_1 _08730_ (.A(_01269_),
    .X(_01270_));
 sg13g2_xnor2_1 _08731_ (.Y(_01271_),
    .A(_00846_),
    .B(_01270_));
 sg13g2_o21ai_1 _08732_ (.B1(net236),
    .Y(_01272_),
    .A1(net96),
    .A2(_01271_));
 sg13g2_nand2_1 _08733_ (.Y(_01273_),
    .A(_01057_),
    .B(_01054_));
 sg13g2_buf_2 _08734_ (.A(_01273_),
    .X(_01274_));
 sg13g2_buf_8 _08735_ (.A(_01274_),
    .X(_01275_));
 sg13g2_nor2_1 _08736_ (.A(_01262_),
    .B(net95),
    .Y(_01276_));
 sg13g2_a22oi_1 _08737_ (.Y(_01277_),
    .B1(_01276_),
    .B2(_01271_),
    .A2(_01272_),
    .A1(_01262_));
 sg13g2_inv_1 _08738_ (.Y(_00112_),
    .A(_01277_));
 sg13g2_inv_1 _08739_ (.Y(_01278_),
    .A(\clock_inst.hour_tile.e0[23] ));
 sg13g2_buf_1 _08740_ (.A(net150),
    .X(_01279_));
 sg13g2_a21o_1 _08741_ (.A2(_01270_),
    .A1(_01262_),
    .B1(\clock_inst.hour_b[22] ),
    .X(_01280_));
 sg13g2_o21ai_1 _08742_ (.B1(_01280_),
    .Y(_01281_),
    .A1(_01262_),
    .A2(_01270_));
 sg13g2_xnor2_1 _08743_ (.Y(_01282_),
    .A(\clock_inst.hour_b[23] ),
    .B(\clock_inst.hour_tile.e0[23] ));
 sg13g2_xnor2_1 _08744_ (.Y(_01283_),
    .A(_01281_),
    .B(_01282_));
 sg13g2_buf_1 _08745_ (.A(_01052_),
    .X(_01284_));
 sg13g2_nor2_1 _08746_ (.A(\clock_inst.hour_c[23] ),
    .B(net235),
    .Y(_01285_));
 sg13g2_a21oi_1 _08747_ (.A1(net94),
    .A2(_01283_),
    .Y(_01286_),
    .B1(_01285_));
 sg13g2_nor2_1 _08748_ (.A(_01064_),
    .B(_01286_),
    .Y(_01287_));
 sg13g2_a21oi_1 _08749_ (.A1(_01278_),
    .A2(net100),
    .Y(_00113_),
    .B1(_01287_));
 sg13g2_buf_1 _08750_ (.A(\clock_inst.hour_tile.e0[24] ),
    .X(_01288_));
 sg13g2_inv_2 _08751_ (.Y(_01289_),
    .A(_01288_));
 sg13g2_nor2_1 _08752_ (.A(_00850_),
    .B(_01278_),
    .Y(_01290_));
 sg13g2_a221oi_1 _08753_ (.B2(_01268_),
    .C1(_01290_),
    .B1(_01265_),
    .A1(\clock_inst.hour_b[22] ),
    .Y(_01291_),
    .A2(_01262_));
 sg13g2_buf_1 _08754_ (.A(_01291_),
    .X(_01292_));
 sg13g2_buf_8 _08755_ (.A(_01292_),
    .X(_01293_));
 sg13g2_or3_1 _08756_ (.A(\clock_inst.hour_b[22] ),
    .B(_01262_),
    .C(_01290_),
    .X(_01294_));
 sg13g2_o21ai_1 _08757_ (.B1(_01294_),
    .Y(_01295_),
    .A1(\clock_inst.hour_b[23] ),
    .A2(\clock_inst.hour_tile.e0[23] ));
 sg13g2_buf_1 _08758_ (.A(_01295_),
    .X(_01296_));
 sg13g2_buf_1 _08759_ (.A(_01296_),
    .X(_01297_));
 sg13g2_or2_1 _08760_ (.X(_01298_),
    .B(net234),
    .A(net149));
 sg13g2_buf_1 _08761_ (.A(_01298_),
    .X(_01299_));
 sg13g2_nand2_1 _08762_ (.Y(_01300_),
    .A(net576),
    .B(_01289_));
 sg13g2_inv_1 _08763_ (.Y(_01301_),
    .A(_01300_));
 sg13g2_nor2_1 _08764_ (.A(_00858_),
    .B(_01289_),
    .Y(_01302_));
 sg13g2_nor2_1 _08765_ (.A(_01301_),
    .B(_01302_),
    .Y(_01303_));
 sg13g2_xnor2_1 _08766_ (.Y(_01304_),
    .A(_01299_),
    .B(_01303_));
 sg13g2_nand2_1 _08767_ (.Y(_01305_),
    .A(\clock_inst.hour_c[24] ),
    .B(net109));
 sg13g2_o21ai_1 _08768_ (.B1(_01305_),
    .Y(_01306_),
    .A1(net110),
    .A2(_01304_));
 sg13g2_nor2_1 _08769_ (.A(_01064_),
    .B(_01306_),
    .Y(_01307_));
 sg13g2_a21oi_1 _08770_ (.A1(_01289_),
    .A2(net100),
    .Y(_00114_),
    .B1(_01307_));
 sg13g2_buf_2 _08771_ (.A(\clock_inst.hour_tile.e0[25] ),
    .X(_01308_));
 sg13g2_inv_1 _08772_ (.Y(_01309_),
    .A(_01308_));
 sg13g2_buf_1 _08773_ (.A(net242),
    .X(_01310_));
 sg13g2_o21ai_1 _08774_ (.B1(_01289_),
    .Y(_01311_),
    .A1(net149),
    .A2(net234));
 sg13g2_or4_1 _08775_ (.A(net576),
    .B(_01289_),
    .C(net149),
    .D(_01297_),
    .X(_01312_));
 sg13g2_o21ai_1 _08776_ (.B1(_01312_),
    .Y(_01313_),
    .A1(_01266_),
    .A2(_01311_));
 sg13g2_xnor2_1 _08777_ (.Y(_01314_),
    .A(_01308_),
    .B(_01313_));
 sg13g2_nand2_1 _08778_ (.Y(_01315_),
    .A(\clock_inst.hour_c[25] ),
    .B(net109));
 sg13g2_o21ai_1 _08779_ (.B1(_01315_),
    .Y(_01316_),
    .A1(net110),
    .A2(_01314_));
 sg13g2_nor2_1 _08780_ (.A(net148),
    .B(_01316_),
    .Y(_01317_));
 sg13g2_a21oi_1 _08781_ (.A1(_01309_),
    .A2(net100),
    .Y(_00115_),
    .B1(_01317_));
 sg13g2_buf_2 _08782_ (.A(\clock_inst.hour_tile.e0[26] ),
    .X(_01318_));
 sg13g2_inv_1 _08783_ (.Y(_01319_),
    .A(_01318_));
 sg13g2_nand2_1 _08784_ (.Y(_01320_),
    .A(_01266_),
    .B(_01288_));
 sg13g2_or4_1 _08785_ (.A(_01309_),
    .B(_01292_),
    .C(_01296_),
    .D(_01320_),
    .X(_01321_));
 sg13g2_buf_1 _08786_ (.A(_01321_),
    .X(_01322_));
 sg13g2_nor2_1 _08787_ (.A(_01308_),
    .B(_01300_),
    .Y(_01323_));
 sg13g2_o21ai_1 _08788_ (.B1(_01323_),
    .Y(_01324_),
    .A1(net149),
    .A2(net234));
 sg13g2_buf_1 _08789_ (.A(_01324_),
    .X(_01325_));
 sg13g2_nand2_1 _08790_ (.Y(_01326_),
    .A(_01322_),
    .B(_01325_));
 sg13g2_xnor2_1 _08791_ (.Y(_01327_),
    .A(_01318_),
    .B(_01326_));
 sg13g2_nand2_1 _08792_ (.Y(_01328_),
    .A(\clock_inst.hour_c[26] ),
    .B(net109));
 sg13g2_o21ai_1 _08793_ (.B1(_01328_),
    .Y(_01329_),
    .A1(net110),
    .A2(_01327_));
 sg13g2_nor2_1 _08794_ (.A(net148),
    .B(_01329_),
    .Y(_01330_));
 sg13g2_a21oi_1 _08795_ (.A1(_01319_),
    .A2(net100),
    .Y(_00116_),
    .B1(_01330_));
 sg13g2_buf_2 _08796_ (.A(\clock_inst.hour_tile.e0[27] ),
    .X(_01331_));
 sg13g2_inv_1 _08797_ (.Y(_01332_),
    .A(_01331_));
 sg13g2_mux2_1 _08798_ (.A0(_01322_),
    .A1(_01325_),
    .S(_01319_),
    .X(_01333_));
 sg13g2_xnor2_1 _08799_ (.Y(_01334_),
    .A(_01332_),
    .B(_01333_));
 sg13g2_nand2_1 _08800_ (.Y(_01335_),
    .A(\clock_inst.hour_c[27] ),
    .B(net109));
 sg13g2_o21ai_1 _08801_ (.B1(_01335_),
    .Y(_01336_),
    .A1(_01072_),
    .A2(_01334_));
 sg13g2_nor2_1 _08802_ (.A(net148),
    .B(_01336_),
    .Y(_01337_));
 sg13g2_a21oi_1 _08803_ (.A1(_01332_),
    .A2(net100),
    .Y(_00117_),
    .B1(_01337_));
 sg13g2_buf_1 _08804_ (.A(\clock_inst.hour_tile.e0[28] ),
    .X(_01338_));
 sg13g2_inv_1 _08805_ (.Y(_01339_),
    .A(_01338_));
 sg13g2_nand2_1 _08806_ (.Y(_01340_),
    .A(_01318_),
    .B(_01331_));
 sg13g2_nor2_1 _08807_ (.A(_01322_),
    .B(_01340_),
    .Y(_01341_));
 sg13g2_nor3_1 _08808_ (.A(_01318_),
    .B(_01331_),
    .C(_01325_),
    .Y(_01342_));
 sg13g2_o21ai_1 _08809_ (.B1(_01338_),
    .Y(_01343_),
    .A1(_01341_),
    .A2(_01342_));
 sg13g2_or3_1 _08810_ (.A(_01338_),
    .B(_01341_),
    .C(_01342_),
    .X(_01344_));
 sg13g2_a21o_1 _08811_ (.A2(_01344_),
    .A1(_01343_),
    .B1(_01210_),
    .X(_01345_));
 sg13g2_nand2b_1 _08812_ (.Y(_01346_),
    .B(_01252_),
    .A_N(\clock_inst.hour_c[28] ));
 sg13g2_buf_1 _08813_ (.A(net244),
    .X(_01347_));
 sg13g2_a21oi_1 _08814_ (.A1(_01345_),
    .A2(_01346_),
    .Y(_01348_),
    .B1(_01347_));
 sg13g2_a21oi_1 _08815_ (.A1(_01339_),
    .A2(net100),
    .Y(_00118_),
    .B1(_01348_));
 sg13g2_buf_1 _08816_ (.A(\clock_inst.hour_tile.e0[29] ),
    .X(_01349_));
 sg13g2_buf_2 _08817_ (.A(net150),
    .X(_01350_));
 sg13g2_nor4_1 _08818_ (.A(_01309_),
    .B(_01339_),
    .C(_01299_),
    .D(_01340_),
    .Y(_01351_));
 sg13g2_o21ai_1 _08819_ (.B1(_01309_),
    .Y(_01352_),
    .A1(_01293_),
    .A2(net234));
 sg13g2_nor4_1 _08820_ (.A(_01318_),
    .B(_01331_),
    .C(_01338_),
    .D(_01352_),
    .Y(_01353_));
 sg13g2_a22oi_1 _08821_ (.Y(_01354_),
    .B1(_01353_),
    .B2(_01301_),
    .A2(_01351_),
    .A1(_01302_));
 sg13g2_xor2_1 _08822_ (.B(_01354_),
    .A(_01349_),
    .X(_01355_));
 sg13g2_buf_1 _08823_ (.A(net151),
    .X(_01356_));
 sg13g2_o21ai_1 _08824_ (.B1(_01135_),
    .Y(_01357_),
    .A1(\clock_inst.hour_c[29] ),
    .A2(_01356_));
 sg13g2_a21oi_1 _08825_ (.A1(net93),
    .A2(_01355_),
    .Y(_01358_),
    .B1(_01357_));
 sg13g2_a21o_1 _08826_ (.A2(net112),
    .A1(_01349_),
    .B1(_01358_),
    .X(_00119_));
 sg13g2_inv_1 _08827_ (.Y(_01359_),
    .A(_01080_));
 sg13g2_buf_1 _08828_ (.A(_01130_),
    .X(_01360_));
 sg13g2_nor2_1 _08829_ (.A(_01084_),
    .B(_01085_),
    .Y(_01361_));
 sg13g2_xnor2_1 _08830_ (.Y(_01362_),
    .A(_00852_),
    .B(_01080_));
 sg13g2_xnor2_1 _08831_ (.Y(_01363_),
    .A(_01361_),
    .B(_01362_));
 sg13g2_a21o_1 _08832_ (.A2(net159),
    .A1(\clock_inst.hour_c[2] ),
    .B1(net239),
    .X(_01364_));
 sg13g2_a21oi_1 _08833_ (.A1(net91),
    .A2(_01363_),
    .Y(_01365_),
    .B1(_01364_));
 sg13g2_a21oi_1 _08834_ (.A1(_01359_),
    .A2(_01230_),
    .Y(_00120_),
    .B1(_01365_));
 sg13g2_buf_2 _08835_ (.A(\clock_inst.hour_tile.e0[30] ),
    .X(_01366_));
 sg13g2_or4_1 _08836_ (.A(_01318_),
    .B(_01331_),
    .C(_01338_),
    .D(_01349_),
    .X(_01367_));
 sg13g2_buf_1 _08837_ (.A(_01367_),
    .X(_01368_));
 sg13g2_o21ai_1 _08838_ (.B1(_00858_),
    .Y(_01369_),
    .A1(_01352_),
    .A2(_01368_));
 sg13g2_nand4_1 _08839_ (.B(_01331_),
    .C(_01338_),
    .A(_01318_),
    .Y(_01370_),
    .D(_01349_));
 sg13g2_buf_1 _08840_ (.A(_01370_),
    .X(_01371_));
 sg13g2_nor4_1 _08841_ (.A(_01309_),
    .B(_01293_),
    .C(_01297_),
    .D(_01371_),
    .Y(_01372_));
 sg13g2_o21ai_1 _08842_ (.B1(_01288_),
    .Y(_01373_),
    .A1(net544),
    .A2(_01372_));
 sg13g2_nand2_1 _08843_ (.Y(_01374_),
    .A(_01369_),
    .B(_01373_));
 sg13g2_xor2_1 _08844_ (.B(_01366_),
    .A(net544),
    .X(_01375_));
 sg13g2_xnor2_1 _08845_ (.Y(_01376_),
    .A(_01374_),
    .B(_01375_));
 sg13g2_buf_1 _08846_ (.A(net158),
    .X(_01377_));
 sg13g2_nand2_1 _08847_ (.Y(_01378_),
    .A(\clock_inst.hour_c[30] ),
    .B(_01377_));
 sg13g2_o21ai_1 _08848_ (.B1(_01378_),
    .Y(_01379_),
    .A1(net98),
    .A2(_01376_));
 sg13g2_buf_1 _08849_ (.A(_01057_),
    .X(_01380_));
 sg13g2_buf_1 _08850_ (.A(net233),
    .X(_01381_));
 sg13g2_mux2_1 _08851_ (.A0(_01366_),
    .A1(_01379_),
    .S(net146),
    .X(_00121_));
 sg13g2_nor3_1 _08852_ (.A(_01366_),
    .B(_01325_),
    .C(_01368_),
    .Y(_01382_));
 sg13g2_inv_1 _08853_ (.Y(_01383_),
    .A(_01366_));
 sg13g2_nor3_1 _08854_ (.A(_01383_),
    .B(_01322_),
    .C(_01371_),
    .Y(_01384_));
 sg13g2_nor2_1 _08855_ (.A(_01382_),
    .B(_01384_),
    .Y(_01385_));
 sg13g2_buf_2 _08856_ (.A(\clock_inst.hour_tile.e0[31] ),
    .X(_01386_));
 sg13g2_nand3b_1 _08857_ (.B(_01386_),
    .C(net235),
    .Y(_01387_),
    .A_N(_01385_));
 sg13g2_o21ai_1 _08858_ (.B1(_01387_),
    .Y(_01388_),
    .A1(_00964_),
    .A2(net152));
 sg13g2_a21oi_1 _08859_ (.A1(net93),
    .A2(_01385_),
    .Y(_01389_),
    .B1(net154));
 sg13g2_nor2_1 _08860_ (.A(_01386_),
    .B(_01389_),
    .Y(_01390_));
 sg13g2_a21oi_1 _08861_ (.A1(net103),
    .A2(_01388_),
    .Y(_00122_),
    .B1(_01390_));
 sg13g2_buf_2 _08862_ (.A(\clock_inst.hour_tile.e0[32] ),
    .X(_01391_));
 sg13g2_inv_1 _08863_ (.Y(_01392_),
    .A(_01391_));
 sg13g2_buf_2 _08864_ (.A(_01162_),
    .X(_01393_));
 sg13g2_mux2_1 _08865_ (.A0(_01382_),
    .A1(_01384_),
    .S(_01386_),
    .X(_01394_));
 sg13g2_o21ai_1 _08866_ (.B1(net155),
    .Y(_01395_),
    .A1(net48),
    .A2(_01394_));
 sg13g2_nand3_1 _08867_ (.B(net152),
    .C(_01394_),
    .A(_01391_),
    .Y(_01396_));
 sg13g2_o21ai_1 _08868_ (.B1(_01396_),
    .Y(_01397_),
    .A1(\clock_inst.hour_c[32] ),
    .A2(net152));
 sg13g2_a22oi_1 _08869_ (.Y(_00123_),
    .B1(_01397_),
    .B2(net103),
    .A2(_01395_),
    .A1(_01392_));
 sg13g2_inv_1 _08870_ (.Y(_01398_),
    .A(\clock_inst.hour_tile.e0[33] ));
 sg13g2_nor2_1 _08871_ (.A(_01386_),
    .B(_01391_),
    .Y(_01399_));
 sg13g2_nor4_1 _08872_ (.A(_00857_),
    .B(_01309_),
    .C(_01383_),
    .D(_01371_),
    .Y(_01400_));
 sg13g2_nand3_1 _08873_ (.B(_01391_),
    .C(_01400_),
    .A(_01386_),
    .Y(_01401_));
 sg13g2_nor3_1 _08874_ (.A(_01289_),
    .B(_01299_),
    .C(_01401_),
    .Y(_01402_));
 sg13g2_a21oi_1 _08875_ (.A1(_01382_),
    .A2(_01399_),
    .Y(_01403_),
    .B1(_01402_));
 sg13g2_xnor2_1 _08876_ (.Y(_01404_),
    .A(\clock_inst.hour_tile.e0[33] ),
    .B(_01403_));
 sg13g2_nand2_1 _08877_ (.Y(_01405_),
    .A(\clock_inst.hour_c[33] ),
    .B(_01070_));
 sg13g2_nand2_1 _08878_ (.Y(_01406_),
    .A(_01380_),
    .B(_01405_));
 sg13g2_a21oi_1 _08879_ (.A1(net91),
    .A2(_01404_),
    .Y(_01407_),
    .B1(_01406_));
 sg13g2_a21oi_1 _08880_ (.A1(_01398_),
    .A2(net100),
    .Y(_00124_),
    .B1(_01407_));
 sg13g2_buf_1 _08881_ (.A(\clock_inst.hour_tile.e0[34] ),
    .X(_01408_));
 sg13g2_buf_8 _08882_ (.A(net242),
    .X(_01409_));
 sg13g2_nor4_2 _08883_ (.A(_01366_),
    .B(_01386_),
    .C(_01391_),
    .Y(_01410_),
    .D(_01368_));
 sg13g2_nand2_1 _08884_ (.Y(_01411_),
    .A(_01398_),
    .B(_01410_));
 sg13g2_nand4_1 _08885_ (.B(_01408_),
    .C(_01055_),
    .A(net544),
    .Y(_01412_),
    .D(_01411_));
 sg13g2_a21oi_1 _08886_ (.A1(_01405_),
    .A2(_01412_),
    .Y(_01413_),
    .B1(_01031_));
 sg13g2_a21oi_1 _08887_ (.A1(_01408_),
    .A2(net145),
    .Y(_01414_),
    .B1(_01413_));
 sg13g2_inv_1 _08888_ (.Y(_01415_),
    .A(_01408_));
 sg13g2_nand3_1 _08889_ (.B(_01415_),
    .C(net99),
    .A(_01266_),
    .Y(_01416_));
 sg13g2_nand3_1 _08890_ (.B(_01408_),
    .C(_01239_),
    .A(net544),
    .Y(_01417_));
 sg13g2_nand4_1 _08891_ (.B(_01288_),
    .C(_01398_),
    .A(net576),
    .Y(_01418_),
    .D(_01410_));
 sg13g2_nand4_1 _08892_ (.B(_01308_),
    .C(_01398_),
    .A(net576),
    .Y(_01419_),
    .D(_01410_));
 sg13g2_or4_1 _08893_ (.A(_01266_),
    .B(net149),
    .C(net234),
    .D(_01411_),
    .X(_01420_));
 sg13g2_nand3_1 _08894_ (.B(_01386_),
    .C(_01391_),
    .A(_01366_),
    .Y(_01421_));
 sg13g2_nor4_1 _08895_ (.A(net576),
    .B(_01398_),
    .C(_01371_),
    .D(_01421_),
    .Y(_01422_));
 sg13g2_nand3_1 _08896_ (.B(_01308_),
    .C(_01422_),
    .A(_01288_),
    .Y(_01423_));
 sg13g2_or3_1 _08897_ (.A(net149),
    .B(net234),
    .C(_01423_),
    .X(_01424_));
 sg13g2_and4_1 _08898_ (.A(_01418_),
    .B(_01419_),
    .C(_01420_),
    .D(_01424_),
    .X(_01425_));
 sg13g2_a21o_1 _08899_ (.A2(_01417_),
    .A1(_01416_),
    .B1(_01425_),
    .X(_01426_));
 sg13g2_nor4_1 _08900_ (.A(_01266_),
    .B(_01408_),
    .C(_01274_),
    .D(_01411_),
    .Y(_01427_));
 sg13g2_nor3_1 _08901_ (.A(net544),
    .B(_01415_),
    .C(_01274_),
    .Y(_01428_));
 sg13g2_o21ai_1 _08902_ (.B1(_01425_),
    .Y(_01429_),
    .A1(_01427_),
    .A2(_01428_));
 sg13g2_nand3_1 _08903_ (.B(_01426_),
    .C(_01429_),
    .A(_01414_),
    .Y(_00125_));
 sg13g2_nor4_1 _08904_ (.A(_01308_),
    .B(_01408_),
    .C(_01300_),
    .D(_01411_),
    .Y(_01430_));
 sg13g2_o21ai_1 _08905_ (.B1(_01430_),
    .Y(_01431_),
    .A1(net149),
    .A2(net234));
 sg13g2_or4_1 _08906_ (.A(_01289_),
    .B(_01398_),
    .C(_01415_),
    .D(_01401_),
    .X(_01432_));
 sg13g2_or3_1 _08907_ (.A(net149),
    .B(net234),
    .C(_01432_),
    .X(_01433_));
 sg13g2_a21oi_1 _08908_ (.A1(_01431_),
    .A2(_01433_),
    .Y(_01434_),
    .B1(\clock_inst.hour_tile.e0[35] ));
 sg13g2_and3_1 _08909_ (.X(_01435_),
    .A(\clock_inst.hour_tile.e0[35] ),
    .B(_01431_),
    .C(_01433_));
 sg13g2_o21ai_1 _08910_ (.B1(_01055_),
    .Y(_01436_),
    .A1(_01434_),
    .A2(_01435_));
 sg13g2_a21oi_1 _08911_ (.A1(_01405_),
    .A2(_01436_),
    .Y(_01437_),
    .B1(_01032_));
 sg13g2_a21o_1 _08912_ (.A2(net112),
    .A1(\clock_inst.hour_tile.e0[35] ),
    .B1(_01437_),
    .X(_00126_));
 sg13g2_buf_8 _08913_ (.A(\clock_inst.hour_tile.e0[36] ),
    .X(_01438_));
 sg13g2_xnor2_1 _08914_ (.Y(_01439_),
    .A(_00862_),
    .B(_01438_));
 sg13g2_a21oi_1 _08915_ (.A1(_01178_),
    .A2(_01439_),
    .Y(_01440_),
    .B1(_01058_));
 sg13g2_a21o_1 _08916_ (.A2(net112),
    .A1(_01438_),
    .B1(_01440_),
    .X(_00127_));
 sg13g2_buf_8 _08917_ (.A(\clock_inst.hour_tile.e0[37] ),
    .X(_01441_));
 sg13g2_inv_1 _08918_ (.Y(_01442_),
    .A(_01441_));
 sg13g2_buf_1 _08919_ (.A(_01061_),
    .X(_01443_));
 sg13g2_nand2_1 _08920_ (.Y(_01444_),
    .A(_00862_),
    .B(_01438_));
 sg13g2_xnor2_1 _08921_ (.Y(_01445_),
    .A(_00866_),
    .B(_01441_));
 sg13g2_xnor2_1 _08922_ (.Y(_01446_),
    .A(_01444_),
    .B(_01445_));
 sg13g2_nand2_1 _08923_ (.Y(_01447_),
    .A(\clock_inst.hour_c[37] ),
    .B(net109));
 sg13g2_o21ai_1 _08924_ (.B1(_01447_),
    .Y(_01448_),
    .A1(_01072_),
    .A2(_01446_));
 sg13g2_nor2_1 _08925_ (.A(net148),
    .B(_01448_),
    .Y(_01449_));
 sg13g2_a21oi_1 _08926_ (.A1(_01442_),
    .A2(net89),
    .Y(_00128_),
    .B1(_01449_));
 sg13g2_buf_8 _08927_ (.A(\clock_inst.hour_tile.e0[38] ),
    .X(_01450_));
 sg13g2_inv_1 _08928_ (.Y(_01451_),
    .A(_01450_));
 sg13g2_a21o_1 _08929_ (.A2(_01438_),
    .A1(_00862_),
    .B1(_01441_),
    .X(_01452_));
 sg13g2_and3_1 _08930_ (.X(_01453_),
    .A(_01441_),
    .B(_00862_),
    .C(_01438_));
 sg13g2_a21oi_1 _08931_ (.A1(_00866_),
    .A2(_01452_),
    .Y(_01454_),
    .B1(_01453_));
 sg13g2_xor2_1 _08932_ (.B(_01450_),
    .A(_00869_),
    .X(_01455_));
 sg13g2_xnor2_1 _08933_ (.Y(_01456_),
    .A(_01454_),
    .B(_01455_));
 sg13g2_a21oi_1 _08934_ (.A1(net91),
    .A2(_01456_),
    .Y(_01457_),
    .B1(_01364_));
 sg13g2_a21oi_1 _08935_ (.A1(_01451_),
    .A2(net89),
    .Y(_00129_),
    .B1(_01457_));
 sg13g2_buf_2 _08936_ (.A(net156),
    .X(_01458_));
 sg13g2_buf_1 _08937_ (.A(\clock_inst.hour_tile.e0[39] ),
    .X(_01459_));
 sg13g2_buf_1 _08938_ (.A(net150),
    .X(_01460_));
 sg13g2_inv_1 _08939_ (.Y(_01461_),
    .A(_00873_));
 sg13g2_nand2_1 _08940_ (.Y(_01462_),
    .A(_00869_),
    .B(_01450_));
 sg13g2_or2_1 _08941_ (.X(_01463_),
    .B(_01450_),
    .A(_00869_));
 sg13g2_nand2_1 _08942_ (.Y(_01464_),
    .A(_01453_),
    .B(_01463_));
 sg13g2_nand3_1 _08943_ (.B(_01452_),
    .C(_01463_),
    .A(_00866_),
    .Y(_01465_));
 sg13g2_nand3_1 _08944_ (.B(_01464_),
    .C(_01465_),
    .A(_01462_),
    .Y(_01466_));
 sg13g2_buf_1 _08945_ (.A(_01466_),
    .X(_01467_));
 sg13g2_xnor2_1 _08946_ (.Y(_01468_),
    .A(_01461_),
    .B(_01467_));
 sg13g2_nand3_1 _08947_ (.B(net87),
    .C(_01468_),
    .A(_01459_),
    .Y(_01469_));
 sg13g2_o21ai_1 _08948_ (.B1(_01469_),
    .Y(_01470_),
    .A1(\clock_inst.hour_c[2] ),
    .A2(_01213_));
 sg13g2_buf_2 _08949_ (.A(net90),
    .X(_01471_));
 sg13g2_buf_1 _08950_ (.A(net233),
    .X(_01472_));
 sg13g2_o21ai_1 _08951_ (.B1(_01472_),
    .Y(_01473_),
    .A1(_01471_),
    .A2(_01468_));
 sg13g2_inv_1 _08952_ (.Y(_01474_),
    .A(_01459_));
 sg13g2_a22oi_1 _08953_ (.Y(_00130_),
    .B1(_01473_),
    .B2(_01474_),
    .A2(_01470_),
    .A1(_01458_));
 sg13g2_nor2_1 _08954_ (.A(_00853_),
    .B(_01359_),
    .Y(_01475_));
 sg13g2_nor3_1 _08955_ (.A(_01082_),
    .B(_01084_),
    .C(_01085_),
    .Y(_01476_));
 sg13g2_nor2_1 _08956_ (.A(_01475_),
    .B(_01476_),
    .Y(_01477_));
 sg13g2_xor2_1 _08957_ (.B(_01078_),
    .A(_00827_),
    .X(_01478_));
 sg13g2_xnor2_1 _08958_ (.Y(_01479_),
    .A(_01477_),
    .B(_01478_));
 sg13g2_a21oi_1 _08959_ (.A1(net91),
    .A2(_01479_),
    .Y(_01480_),
    .B1(_01364_));
 sg13g2_a21oi_1 _08960_ (.A1(_01079_),
    .A2(net89),
    .Y(_00131_),
    .B1(_01480_));
 sg13g2_buf_2 _08961_ (.A(\clock_inst.hour_tile.e0[40] ),
    .X(_01481_));
 sg13g2_inv_1 _08962_ (.Y(_01482_),
    .A(_01481_));
 sg13g2_xor2_1 _08963_ (.B(_01481_),
    .A(_00876_),
    .X(_01483_));
 sg13g2_a21o_1 _08964_ (.A2(_01467_),
    .A1(_00873_),
    .B1(_01459_),
    .X(_01484_));
 sg13g2_o21ai_1 _08965_ (.B1(_01484_),
    .Y(_01485_),
    .A1(_00873_),
    .A2(_01467_));
 sg13g2_xnor2_1 _08966_ (.Y(_01486_),
    .A(_01483_),
    .B(_01485_));
 sg13g2_a21oi_1 _08967_ (.A1(\clock_inst.hour_c[40] ),
    .A2(_01071_),
    .Y(_01487_),
    .B1(_01151_));
 sg13g2_inv_1 _08968_ (.Y(_01488_),
    .A(_01487_));
 sg13g2_a21oi_1 _08969_ (.A1(_01360_),
    .A2(_01486_),
    .Y(_01489_),
    .B1(_01488_));
 sg13g2_a21oi_1 _08970_ (.A1(_01482_),
    .A2(_01443_),
    .Y(_00132_),
    .B1(_01489_));
 sg13g2_buf_8 _08971_ (.A(\clock_inst.hour_tile.e0[41] ),
    .X(_01490_));
 sg13g2_inv_1 _08972_ (.Y(_01491_),
    .A(_01490_));
 sg13g2_buf_2 _08973_ (.A(net158),
    .X(_01492_));
 sg13g2_nand2_1 _08974_ (.Y(_01493_),
    .A(_00876_),
    .B(_01481_));
 sg13g2_and2_1 _08975_ (.A(_01462_),
    .B(_01493_),
    .X(_01494_));
 sg13g2_nand4_1 _08976_ (.B(_01464_),
    .C(_01465_),
    .A(_01474_),
    .Y(_01495_),
    .D(_01494_));
 sg13g2_nand4_1 _08977_ (.B(_01464_),
    .C(_01465_),
    .A(_01461_),
    .Y(_01496_),
    .D(_01494_));
 sg13g2_nor2_1 _08978_ (.A(_00873_),
    .B(_01459_),
    .Y(_01497_));
 sg13g2_nor2_1 _08979_ (.A(_00876_),
    .B(_01481_),
    .Y(_01498_));
 sg13g2_a21oi_1 _08980_ (.A1(_01493_),
    .A2(_01497_),
    .Y(_01499_),
    .B1(_01498_));
 sg13g2_nand3_1 _08981_ (.B(_01496_),
    .C(_01499_),
    .A(_01495_),
    .Y(_01500_));
 sg13g2_buf_1 _08982_ (.A(_01500_),
    .X(_01501_));
 sg13g2_xnor2_1 _08983_ (.Y(_01502_),
    .A(_00880_),
    .B(_01490_));
 sg13g2_xnor2_1 _08984_ (.Y(_01503_),
    .A(_01501_),
    .B(_01502_));
 sg13g2_buf_2 _08985_ (.A(net158),
    .X(_01504_));
 sg13g2_nand2_1 _08986_ (.Y(_01505_),
    .A(\clock_inst.hour_c[41] ),
    .B(net85));
 sg13g2_o21ai_1 _08987_ (.B1(_01505_),
    .Y(_01506_),
    .A1(net86),
    .A2(_01503_));
 sg13g2_nor2_1 _08988_ (.A(net148),
    .B(_01506_),
    .Y(_01507_));
 sg13g2_a21oi_1 _08989_ (.A1(_01491_),
    .A2(net89),
    .Y(_00133_),
    .B1(_01507_));
 sg13g2_buf_1 _08990_ (.A(\clock_inst.hour_tile.e0[42] ),
    .X(_01508_));
 sg13g2_inv_1 _08991_ (.Y(_01509_),
    .A(_01508_));
 sg13g2_nand2_1 _08992_ (.Y(_01510_),
    .A(_00880_),
    .B(_01490_));
 sg13g2_nor2_1 _08993_ (.A(_00880_),
    .B(_01490_),
    .Y(_01511_));
 sg13g2_a21oi_1 _08994_ (.A1(_01501_),
    .A2(_01510_),
    .Y(_01512_),
    .B1(_01511_));
 sg13g2_xor2_1 _08995_ (.B(_01508_),
    .A(_00887_),
    .X(_01513_));
 sg13g2_xnor2_1 _08996_ (.Y(_01514_),
    .A(_01512_),
    .B(_01513_));
 sg13g2_nand2_1 _08997_ (.Y(_01515_),
    .A(\clock_inst.hour_c[42] ),
    .B(_01504_));
 sg13g2_o21ai_1 _08998_ (.B1(_01515_),
    .Y(_01516_),
    .A1(_01492_),
    .A2(_01514_));
 sg13g2_nor2_1 _08999_ (.A(net148),
    .B(_01516_),
    .Y(_01517_));
 sg13g2_a21oi_1 _09000_ (.A1(_01509_),
    .A2(net89),
    .Y(_00134_),
    .B1(_01517_));
 sg13g2_inv_1 _09001_ (.Y(_01518_),
    .A(\clock_inst.hour_tile.e0[43] ));
 sg13g2_buf_2 _09002_ (.A(net150),
    .X(_01519_));
 sg13g2_xnor2_1 _09003_ (.Y(_01520_),
    .A(\clock_inst.hour_tile.e0[43] ),
    .B(net546));
 sg13g2_and2_1 _09004_ (.A(_00887_),
    .B(_01508_),
    .X(_01521_));
 sg13g2_buf_1 _09005_ (.A(_01521_),
    .X(_01522_));
 sg13g2_or2_1 _09006_ (.X(_01523_),
    .B(_01508_),
    .A(_00887_));
 sg13g2_buf_1 _09007_ (.A(_01523_),
    .X(_01524_));
 sg13g2_o21ai_1 _09008_ (.B1(_01524_),
    .Y(_01525_),
    .A1(_01512_),
    .A2(_01522_));
 sg13g2_xnor2_1 _09009_ (.Y(_01526_),
    .A(_01520_),
    .B(_01525_));
 sg13g2_buf_1 _09010_ (.A(_01052_),
    .X(_01527_));
 sg13g2_nor2_1 _09011_ (.A(\clock_inst.hour_c[43] ),
    .B(_01527_),
    .Y(_01528_));
 sg13g2_a21oi_1 _09012_ (.A1(_01519_),
    .A2(_01526_),
    .Y(_01529_),
    .B1(_01528_));
 sg13g2_nor2_1 _09013_ (.A(_01310_),
    .B(_01529_),
    .Y(_01530_));
 sg13g2_a21oi_1 _09014_ (.A1(_01518_),
    .A2(net89),
    .Y(_00135_),
    .B1(_01530_));
 sg13g2_buf_1 _09015_ (.A(\clock_inst.hour_tile.e0[44] ),
    .X(_01531_));
 sg13g2_inv_1 _09016_ (.Y(_01532_),
    .A(_01531_));
 sg13g2_nor3_1 _09017_ (.A(_00731_),
    .B(_01490_),
    .C(_01522_),
    .Y(_01533_));
 sg13g2_nor3_1 _09018_ (.A(_00731_),
    .B(_00880_),
    .C(_01522_),
    .Y(_01534_));
 sg13g2_o21ai_1 _09019_ (.B1(_01501_),
    .Y(_01535_),
    .A1(_01533_),
    .A2(_01534_));
 sg13g2_nor2_1 _09020_ (.A(net546),
    .B(_01524_),
    .Y(_01536_));
 sg13g2_a21oi_1 _09021_ (.A1(_01491_),
    .A2(_01534_),
    .Y(_01537_),
    .B1(_01536_));
 sg13g2_and3_1 _09022_ (.X(_01538_),
    .A(_00731_),
    .B(_01490_),
    .C(_01524_));
 sg13g2_nand4_1 _09023_ (.B(_01496_),
    .C(_01499_),
    .A(_01495_),
    .Y(_01539_),
    .D(_01538_));
 sg13g2_and3_1 _09024_ (.X(_01540_),
    .A(_00731_),
    .B(_00880_),
    .C(_01524_));
 sg13g2_nand4_1 _09025_ (.B(_01496_),
    .C(_01499_),
    .A(_01495_),
    .Y(_01541_),
    .D(_01540_));
 sg13g2_a22oi_1 _09026_ (.Y(_01542_),
    .B1(_01540_),
    .B2(_01490_),
    .A2(_01522_),
    .A1(_00731_));
 sg13g2_nand4_1 _09027_ (.B(_01539_),
    .C(_01541_),
    .A(_01518_),
    .Y(_01543_),
    .D(_01542_));
 sg13g2_and3_1 _09028_ (.X(_01544_),
    .A(_01535_),
    .B(_01537_),
    .C(_01543_));
 sg13g2_buf_1 _09029_ (.A(_01544_),
    .X(_01545_));
 sg13g2_inv_1 _09030_ (.Y(_01546_),
    .A(\clock_inst.hour_a[24] ));
 sg13g2_nand2_1 _09031_ (.Y(_01547_),
    .A(_01546_),
    .B(_01531_));
 sg13g2_nand2_1 _09032_ (.Y(_01548_),
    .A(_00752_),
    .B(_01532_));
 sg13g2_buf_8 _09033_ (.A(_01548_),
    .X(_01549_));
 sg13g2_nand2_1 _09034_ (.Y(_01550_),
    .A(_01547_),
    .B(_01549_));
 sg13g2_xnor2_1 _09035_ (.Y(_01551_),
    .A(net46),
    .B(_01550_));
 sg13g2_nand2_1 _09036_ (.Y(_01552_),
    .A(\clock_inst.hour_c[44] ),
    .B(_01504_));
 sg13g2_o21ai_1 _09037_ (.B1(_01552_),
    .Y(_01553_),
    .A1(_01492_),
    .A2(_01551_));
 sg13g2_nor2_1 _09038_ (.A(_01310_),
    .B(_01553_),
    .Y(_01554_));
 sg13g2_a21oi_1 _09039_ (.A1(_01532_),
    .A2(net89),
    .Y(_00136_),
    .B1(_01554_));
 sg13g2_mux2_1 _09040_ (.A0(_01549_),
    .A1(_01547_),
    .S(net46),
    .X(_01555_));
 sg13g2_buf_2 _09041_ (.A(\clock_inst.hour_tile.e0[45] ),
    .X(_01556_));
 sg13g2_nand3b_1 _09042_ (.B(_01556_),
    .C(net94),
    .Y(_01557_),
    .A_N(_01555_));
 sg13g2_o21ai_1 _09043_ (.B1(_01557_),
    .Y(_01558_),
    .A1(\clock_inst.hour_c[45] ),
    .A2(net50));
 sg13g2_buf_2 _09044_ (.A(net239),
    .X(_01559_));
 sg13g2_a21oi_1 _09045_ (.A1(net93),
    .A2(_01555_),
    .Y(_01560_),
    .B1(net143));
 sg13g2_nor2_1 _09046_ (.A(_01556_),
    .B(_01560_),
    .Y(_01561_));
 sg13g2_a21oi_1 _09047_ (.A1(net103),
    .A2(_01558_),
    .Y(_00137_),
    .B1(_01561_));
 sg13g2_buf_2 _09048_ (.A(\clock_inst.hour_tile.e0[46] ),
    .X(_01562_));
 sg13g2_inv_1 _09049_ (.Y(_01563_),
    .A(_01562_));
 sg13g2_and3_1 _09050_ (.X(_01564_),
    .A(_01546_),
    .B(_01556_),
    .C(_01531_));
 sg13g2_nand2b_1 _09051_ (.Y(_01565_),
    .B(_00752_),
    .A_N(_01556_));
 sg13g2_nor2_1 _09052_ (.A(_01531_),
    .B(_01565_),
    .Y(_01566_));
 sg13g2_nand2_1 _09053_ (.Y(_01567_),
    .A(_01535_),
    .B(_01537_));
 sg13g2_nand3_1 _09054_ (.B(_01541_),
    .C(_01542_),
    .A(_01539_),
    .Y(_01568_));
 sg13g2_nor4_1 _09055_ (.A(_01531_),
    .B(\clock_inst.hour_tile.e0[43] ),
    .C(_01568_),
    .D(_01565_),
    .Y(_01569_));
 sg13g2_a221oi_1 _09056_ (.B2(_01567_),
    .C1(_01569_),
    .B1(_01566_),
    .A1(_01545_),
    .Y(_01570_),
    .A2(_01564_));
 sg13g2_buf_1 _09057_ (.A(_01570_),
    .X(_01571_));
 sg13g2_a21o_1 _09058_ (.A2(_01571_),
    .A1(_01350_),
    .B1(_01176_),
    .X(_01572_));
 sg13g2_buf_1 _09059_ (.A(_01222_),
    .X(_01573_));
 sg13g2_nand3b_1 _09060_ (.B(_01562_),
    .C(net87),
    .Y(_01574_),
    .A_N(_01571_));
 sg13g2_o21ai_1 _09061_ (.B1(_01574_),
    .Y(_01575_),
    .A1(\clock_inst.hour_c[46] ),
    .A2(net45));
 sg13g2_a22oi_1 _09062_ (.Y(_00138_),
    .B1(_01575_),
    .B2(net103),
    .A2(_01572_),
    .A1(_01563_));
 sg13g2_buf_1 _09063_ (.A(\clock_inst.hour_tile.e0[47] ),
    .X(_01576_));
 sg13g2_inv_1 _09064_ (.Y(_01577_),
    .A(_01576_));
 sg13g2_nor3_1 _09065_ (.A(_01562_),
    .B(_01556_),
    .C(_01549_),
    .Y(_01578_));
 sg13g2_and2_1 _09066_ (.A(_01562_),
    .B(_01564_),
    .X(_01579_));
 sg13g2_mux2_1 _09067_ (.A0(_01578_),
    .A1(_01579_),
    .S(net46),
    .X(_01580_));
 sg13g2_xnor2_1 _09068_ (.Y(_01581_),
    .A(_01577_),
    .B(_01580_));
 sg13g2_nor2_1 _09069_ (.A(net95),
    .B(_01581_),
    .Y(_01582_));
 sg13g2_a21oi_1 _09070_ (.A1(_01577_),
    .A2(net89),
    .Y(_00139_),
    .B1(_01582_));
 sg13g2_buf_8 _09071_ (.A(_01275_),
    .X(_01583_));
 sg13g2_buf_8 _09072_ (.A(\clock_inst.hour_tile.e0[48] ),
    .X(_01584_));
 sg13g2_nor2_1 _09073_ (.A(net46),
    .B(_01549_),
    .Y(_01585_));
 sg13g2_nor3_1 _09074_ (.A(_01576_),
    .B(_01562_),
    .C(_01556_),
    .Y(_01586_));
 sg13g2_and2_1 _09075_ (.A(_01576_),
    .B(_01579_),
    .X(_01587_));
 sg13g2_a22oi_1 _09076_ (.Y(_01588_),
    .B1(_01587_),
    .B2(net46),
    .A2(_01586_),
    .A1(_01585_));
 sg13g2_xor2_1 _09077_ (.B(_01588_),
    .A(_01584_),
    .X(_01589_));
 sg13g2_buf_8 _09078_ (.A(net143),
    .X(_01590_));
 sg13g2_nand2_1 _09079_ (.Y(_01591_),
    .A(_01584_),
    .B(net83));
 sg13g2_o21ai_1 _09080_ (.B1(_01591_),
    .Y(_00140_),
    .A1(net44),
    .A2(_01589_));
 sg13g2_buf_8 _09081_ (.A(\clock_inst.hour_tile.e0[49] ),
    .X(_01592_));
 sg13g2_inv_1 _09082_ (.Y(_01593_),
    .A(_01592_));
 sg13g2_and3_1 _09083_ (.X(_01594_),
    .A(_01584_),
    .B(net46),
    .C(_01587_));
 sg13g2_buf_2 _09084_ (.A(_01594_),
    .X(_01595_));
 sg13g2_nand2b_1 _09085_ (.Y(_01596_),
    .B(_01586_),
    .A_N(_01584_));
 sg13g2_nor3_2 _09086_ (.A(net46),
    .B(_01549_),
    .C(_01596_),
    .Y(_01597_));
 sg13g2_or3_1 _09087_ (.A(_01592_),
    .B(_01595_),
    .C(_01597_),
    .X(_01598_));
 sg13g2_o21ai_1 _09088_ (.B1(_01592_),
    .Y(_01599_),
    .A1(_01595_),
    .A2(_01597_));
 sg13g2_nand3_1 _09089_ (.B(_01598_),
    .C(_01599_),
    .A(_01350_),
    .Y(_01600_));
 sg13g2_a21oi_1 _09090_ (.A1(\clock_inst.hour_c[49] ),
    .A2(net237),
    .Y(_01601_),
    .B1(_01033_));
 sg13g2_a22oi_1 _09091_ (.Y(_00141_),
    .B1(_01600_),
    .B2(_01601_),
    .A2(_01177_),
    .A1(_01593_));
 sg13g2_inv_1 _09092_ (.Y(_01602_),
    .A(_01088_));
 sg13g2_o21ai_1 _09093_ (.B1(_01078_),
    .Y(_01603_),
    .A1(_01475_),
    .A2(_01476_));
 sg13g2_nor3_1 _09094_ (.A(_01078_),
    .B(_01475_),
    .C(_01476_),
    .Y(_01604_));
 sg13g2_a21oi_2 _09095_ (.B1(_01604_),
    .Y(_01605_),
    .A2(_01603_),
    .A1(_00828_));
 sg13g2_xor2_1 _09096_ (.B(_01605_),
    .A(_01089_),
    .X(_01606_));
 sg13g2_a21oi_1 _09097_ (.A1(_01360_),
    .A2(_01606_),
    .Y(_01607_),
    .B1(_01488_));
 sg13g2_a21oi_1 _09098_ (.A1(_01602_),
    .A2(_01443_),
    .Y(_00142_),
    .B1(_01607_));
 sg13g2_inv_2 _09099_ (.Y(_01608_),
    .A(\clock_inst.hour_tile.e0[50] ));
 sg13g2_nor2_1 _09100_ (.A(_01031_),
    .B(_01054_),
    .Y(_01609_));
 sg13g2_buf_2 _09101_ (.A(_01609_),
    .X(_01610_));
 sg13g2_buf_8 _09102_ (.A(_01610_),
    .X(_01611_));
 sg13g2_nand2_1 _09103_ (.Y(_01612_),
    .A(\clock_inst.hour_c[50] ),
    .B(net82));
 sg13g2_or4_1 _09104_ (.A(_01592_),
    .B(_01608_),
    .C(_01275_),
    .D(_01597_),
    .X(_01613_));
 sg13g2_nor2_1 _09105_ (.A(_01592_),
    .B(\clock_inst.hour_tile.e0[50] ),
    .Y(_01614_));
 sg13g2_nand3_1 _09106_ (.B(_01597_),
    .C(_01614_),
    .A(net49),
    .Y(_01615_));
 sg13g2_nor2_2 _09107_ (.A(_01593_),
    .B(_01608_),
    .Y(_01616_));
 sg13g2_nand2_1 _09108_ (.Y(_01617_),
    .A(net49),
    .B(_01616_));
 sg13g2_nand3_1 _09109_ (.B(_01608_),
    .C(net49),
    .A(_01592_),
    .Y(_01618_));
 sg13g2_mux2_1 _09110_ (.A0(_01617_),
    .A1(_01618_),
    .S(_01595_),
    .X(_01619_));
 sg13g2_and4_1 _09111_ (.A(_01612_),
    .B(_01613_),
    .C(_01615_),
    .D(_01619_),
    .X(_01620_));
 sg13g2_o21ai_1 _09112_ (.B1(_01620_),
    .Y(_00143_),
    .A1(_01608_),
    .A2(net106));
 sg13g2_buf_8 _09113_ (.A(\clock_inst.hour_tile.e0[51] ),
    .X(_01621_));
 sg13g2_a22oi_1 _09114_ (.Y(_01622_),
    .B1(_01616_),
    .B2(_01595_),
    .A2(_01614_),
    .A1(_01597_));
 sg13g2_xor2_1 _09115_ (.B(_01622_),
    .A(_01621_),
    .X(_01623_));
 sg13g2_a22oi_1 _09116_ (.Y(_01624_),
    .B1(net82),
    .B2(\clock_inst.hour_c[51] ),
    .A2(net145),
    .A1(_01621_));
 sg13g2_o21ai_1 _09117_ (.B1(_01624_),
    .Y(_00144_),
    .A1(net44),
    .A2(_01623_));
 sg13g2_buf_8 _09118_ (.A(\clock_inst.hour_tile.e0[52] ),
    .X(_01625_));
 sg13g2_nor3_1 _09119_ (.A(_01592_),
    .B(\clock_inst.hour_tile.e0[50] ),
    .C(_01621_),
    .Y(_01626_));
 sg13g2_and2_1 _09120_ (.A(_01621_),
    .B(_01616_),
    .X(_01627_));
 sg13g2_a22oi_1 _09121_ (.Y(_01628_),
    .B1(_01627_),
    .B2(_01595_),
    .A2(_01626_),
    .A1(_01597_));
 sg13g2_xor2_1 _09122_ (.B(_01628_),
    .A(_01625_),
    .X(_01629_));
 sg13g2_a22oi_1 _09123_ (.Y(_01630_),
    .B1(net82),
    .B2(\clock_inst.hour_c[52] ),
    .A2(net145),
    .A1(_01625_));
 sg13g2_o21ai_1 _09124_ (.B1(_01630_),
    .Y(_00145_),
    .A1(net44),
    .A2(_01629_));
 sg13g2_inv_1 _09125_ (.Y(_01631_),
    .A(\clock_inst.hour_tile.e0[53] ));
 sg13g2_and4_1 _09126_ (.A(_01546_),
    .B(_01621_),
    .C(_01625_),
    .D(_01616_),
    .X(_01632_));
 sg13g2_nand2b_1 _09127_ (.Y(_01633_),
    .B(_01626_),
    .A_N(_01625_));
 sg13g2_nor4_1 _09128_ (.A(net46),
    .B(_01549_),
    .C(_01596_),
    .D(_01633_),
    .Y(_01634_));
 sg13g2_a21o_1 _09129_ (.A2(_01632_),
    .A1(_01595_),
    .B1(_01634_),
    .X(_01635_));
 sg13g2_buf_1 _09130_ (.A(_01635_),
    .X(_01636_));
 sg13g2_o21ai_1 _09131_ (.B1(net155),
    .Y(_01637_),
    .A1(_01393_),
    .A2(_01636_));
 sg13g2_nor2_1 _09132_ (.A(_01631_),
    .B(_01263_),
    .Y(_01638_));
 sg13g2_nor2_1 _09133_ (.A(_00774_),
    .B(_01460_),
    .Y(_01639_));
 sg13g2_a21o_1 _09134_ (.A2(_01638_),
    .A1(_01636_),
    .B1(_01639_),
    .X(_01640_));
 sg13g2_a22oi_1 _09135_ (.Y(_00146_),
    .B1(_01640_),
    .B2(_01212_),
    .A2(_01637_),
    .A1(_01631_));
 sg13g2_buf_1 _09136_ (.A(net240),
    .X(_01641_));
 sg13g2_a21o_1 _09137_ (.A2(_01605_),
    .A1(_01088_),
    .B1(_00889_),
    .X(_01642_));
 sg13g2_o21ai_1 _09138_ (.B1(_01642_),
    .Y(_01643_),
    .A1(_01088_),
    .A2(_01605_));
 sg13g2_xnor2_1 _09139_ (.Y(_01644_),
    .A(_01087_),
    .B(_01643_));
 sg13g2_nor2_1 _09140_ (.A(\clock_inst.hour_c[5] ),
    .B(net235),
    .Y(_01645_));
 sg13g2_a21oi_1 _09141_ (.A1(_01279_),
    .A2(_01644_),
    .Y(_01646_),
    .B1(_01645_));
 sg13g2_nand2_1 _09142_ (.Y(_01647_),
    .A(net142),
    .B(_01646_));
 sg13g2_o21ai_1 _09143_ (.B1(_01647_),
    .Y(_00147_),
    .A1(_01094_),
    .A2(net106));
 sg13g2_nor2_1 _09144_ (.A(_01092_),
    .B(_01098_),
    .Y(_01648_));
 sg13g2_xnor2_1 _09145_ (.Y(_01649_),
    .A(net546),
    .B(_01075_));
 sg13g2_xnor2_1 _09146_ (.Y(_01650_),
    .A(_01648_),
    .B(_01649_));
 sg13g2_nor2_1 _09147_ (.A(\clock_inst.hour_c[6] ),
    .B(_01284_),
    .Y(_01651_));
 sg13g2_a21oi_1 _09148_ (.A1(_01279_),
    .A2(_01650_),
    .Y(_01652_),
    .B1(_01651_));
 sg13g2_nand2_1 _09149_ (.Y(_01653_),
    .A(net142),
    .B(_01652_));
 sg13g2_o21ai_1 _09150_ (.B1(_01653_),
    .Y(_00148_),
    .A1(_01108_),
    .A2(_01166_));
 sg13g2_buf_1 _09151_ (.A(net161),
    .X(_01654_));
 sg13g2_buf_1 _09152_ (.A(net241),
    .X(_01655_));
 sg13g2_nand2_1 _09153_ (.Y(_01656_),
    .A(net546),
    .B(_01075_));
 sg13g2_a21oi_1 _09154_ (.A1(_01648_),
    .A2(_01656_),
    .Y(_01657_),
    .B1(_01102_));
 sg13g2_xor2_1 _09155_ (.B(\clock_inst.hour_tile.e0[7] ),
    .A(_00724_),
    .X(_01658_));
 sg13g2_xnor2_1 _09156_ (.Y(_01659_),
    .A(_01657_),
    .B(_01658_));
 sg13g2_nand2_1 _09157_ (.Y(_01660_),
    .A(\clock_inst.hour_c[7] ),
    .B(_01071_));
 sg13g2_o21ai_1 _09158_ (.B1(_01660_),
    .Y(_01661_),
    .A1(_01655_),
    .A2(_01659_));
 sg13g2_nor2_1 _09159_ (.A(net143),
    .B(_01661_),
    .Y(_01662_));
 sg13g2_a21oi_1 _09160_ (.A1(_01076_),
    .A2(_01654_),
    .Y(_00149_),
    .B1(_01662_));
 sg13g2_xor2_1 _09161_ (.B(_01073_),
    .A(net577),
    .X(_01663_));
 sg13g2_xnor2_1 _09162_ (.Y(_01664_),
    .A(_01127_),
    .B(_01663_));
 sg13g2_nor2_1 _09163_ (.A(\clock_inst.hour_c[8] ),
    .B(_01527_),
    .Y(_01665_));
 sg13g2_a21oi_1 _09164_ (.A1(_01284_),
    .A2(_01664_),
    .Y(_01666_),
    .B1(_01665_));
 sg13g2_nor2_1 _09165_ (.A(net148),
    .B(_01666_),
    .Y(_01667_));
 sg13g2_a21oi_1 _09166_ (.A1(_01074_),
    .A2(net81),
    .Y(_00150_),
    .B1(_01667_));
 sg13g2_nor2_1 _09167_ (.A(_01106_),
    .B(net146),
    .Y(_01668_));
 sg13g2_or2_1 _09168_ (.X(_01669_),
    .B(_01116_),
    .A(_01107_));
 sg13g2_xnor2_1 _09169_ (.Y(_01670_),
    .A(_01158_),
    .B(_01669_));
 sg13g2_nand2_1 _09170_ (.Y(_01671_),
    .A(_01202_),
    .B(_01670_));
 sg13g2_nand2_1 _09171_ (.Y(_01672_),
    .A(\clock_inst.hour_c[9] ),
    .B(net107));
 sg13g2_nand3_1 _09172_ (.B(_01671_),
    .C(_01672_),
    .A(net236),
    .Y(_01673_));
 sg13g2_nor2b_1 _09173_ (.A(_01668_),
    .B_N(_01673_),
    .Y(_00151_));
 sg13g2_inv_1 _09174_ (.Y(_01674_),
    .A(\clock_inst.hour_tile.e[0] ));
 sg13g2_nand2_2 _09175_ (.Y(_01675_),
    .A(\clock_inst.vga_inst.vga_horizontal_visible ),
    .B(\clock_inst.vga_inst.vga_vertical_visible ));
 sg13g2_buf_1 _09176_ (.A(_01675_),
    .X(_01676_));
 sg13g2_buf_1 _09177_ (.A(net542),
    .X(_01677_));
 sg13g2_nand2_1 _09178_ (.Y(_01678_),
    .A(net239),
    .B(net502));
 sg13g2_buf_1 _09179_ (.A(_01678_),
    .X(_01679_));
 sg13g2_o21ai_1 _09180_ (.B1(_01679_),
    .Y(_01680_),
    .A1(\clock_inst.hour_a[0] ),
    .A2(_01059_));
 sg13g2_buf_1 _09181_ (.A(_01676_),
    .X(_01681_));
 sg13g2_buf_1 _09182_ (.A(net501),
    .X(_01682_));
 sg13g2_nand2_1 _09183_ (.Y(_01683_),
    .A(\clock_inst.hour_a[0] ),
    .B(\clock_inst.hour_tile.e[0] ));
 sg13g2_o21ai_1 _09184_ (.B1(_01559_),
    .Y(_01684_),
    .A1(net448),
    .A2(_01683_));
 sg13g2_nor2b_1 _09185_ (.A(_01059_),
    .B_N(_01684_),
    .Y(_01685_));
 sg13g2_a21oi_1 _09186_ (.A1(_01674_),
    .A2(_01680_),
    .Y(_00152_),
    .B1(_01685_));
 sg13g2_buf_1 _09187_ (.A(_01032_),
    .X(_01686_));
 sg13g2_buf_1 _09188_ (.A(net140),
    .X(_01687_));
 sg13g2_buf_2 _09189_ (.A(\clock_inst.hour_tile.e[10] ),
    .X(_01688_));
 sg13g2_buf_1 _09190_ (.A(\clock_inst.hour_tile.e[7] ),
    .X(_01689_));
 sg13g2_nand2_1 _09191_ (.Y(_01690_),
    .A(_00819_),
    .B(_01689_));
 sg13g2_inv_1 _09192_ (.Y(_01691_),
    .A(\clock_inst.hour_tile.e[4] ));
 sg13g2_inv_1 _09193_ (.Y(_01692_),
    .A(_00964_));
 sg13g2_buf_1 _09194_ (.A(\clock_inst.hour_tile.e[2] ),
    .X(_01693_));
 sg13g2_or2_1 _09195_ (.X(_01694_),
    .B(_01693_),
    .A(_00741_));
 sg13g2_nor2_1 _09196_ (.A(\clock_inst.hour_a[1] ),
    .B(\clock_inst.hour_tile.e[1] ),
    .Y(_01695_));
 sg13g2_nand2_1 _09197_ (.Y(_01696_),
    .A(\clock_inst.hour_a[1] ),
    .B(\clock_inst.hour_tile.e[1] ));
 sg13g2_o21ai_1 _09198_ (.B1(_01696_),
    .Y(_01697_),
    .A1(_01683_),
    .A2(_01695_));
 sg13g2_buf_1 _09199_ (.A(_01697_),
    .X(_01698_));
 sg13g2_and2_1 _09200_ (.A(_00741_),
    .B(_01693_),
    .X(_01699_));
 sg13g2_a21oi_2 _09201_ (.B1(_01699_),
    .Y(_01700_),
    .A2(_01698_),
    .A1(_01694_));
 sg13g2_inv_1 _09202_ (.Y(_01701_),
    .A(_00774_));
 sg13g2_o21ai_1 _09203_ (.B1(_00774_),
    .Y(_01702_),
    .A1(_00741_),
    .A2(_01693_));
 sg13g2_inv_1 _09204_ (.Y(_01703_),
    .A(_01702_));
 sg13g2_a221oi_1 _09205_ (.B2(_01698_),
    .C1(\clock_inst.hour_tile.e[3] ),
    .B1(_01703_),
    .A1(_00774_),
    .Y(_01704_),
    .A2(_01699_));
 sg13g2_a221oi_1 _09206_ (.B2(_01701_),
    .C1(_01704_),
    .B1(_01700_),
    .A1(_01691_),
    .Y(_01705_),
    .A2(_01692_));
 sg13g2_buf_2 _09207_ (.A(_01705_),
    .X(_01706_));
 sg13g2_nor2_2 _09208_ (.A(_01691_),
    .B(_01692_),
    .Y(_01707_));
 sg13g2_buf_1 _09209_ (.A(\clock_inst.hour_tile.e[6] ),
    .X(_01708_));
 sg13g2_inv_1 _09210_ (.Y(_01709_),
    .A(_01708_));
 sg13g2_nor2_1 _09211_ (.A(_00819_),
    .B(_01689_),
    .Y(_01710_));
 sg13g2_buf_1 _09212_ (.A(\clock_inst.hour_tile.e[5] ),
    .X(_01711_));
 sg13g2_nor2_2 _09213_ (.A(_00806_),
    .B(_01711_),
    .Y(_01712_));
 sg13g2_nor3_1 _09214_ (.A(_01709_),
    .B(_01710_),
    .C(_01712_),
    .Y(_01713_));
 sg13g2_o21ai_1 _09215_ (.B1(_01713_),
    .Y(_01714_),
    .A1(_01706_),
    .A2(_01707_));
 sg13g2_nor3_1 _09216_ (.A(_00814_),
    .B(_01710_),
    .C(_01712_),
    .Y(_01715_));
 sg13g2_o21ai_1 _09217_ (.B1(_01715_),
    .Y(_01716_),
    .A1(_01706_),
    .A2(_01707_));
 sg13g2_nand2_1 _09218_ (.Y(_01717_),
    .A(_00813_),
    .B(_01708_));
 sg13g2_nor2_1 _09219_ (.A(_01710_),
    .B(_01717_),
    .Y(_01718_));
 sg13g2_or2_1 _09220_ (.X(_01719_),
    .B(_01689_),
    .A(_00819_));
 sg13g2_and3_1 _09221_ (.X(_01720_),
    .A(_00806_),
    .B(_01711_),
    .C(_01719_));
 sg13g2_o21ai_1 _09222_ (.B1(_01720_),
    .Y(_01721_),
    .A1(_00813_),
    .A2(_01708_));
 sg13g2_nor2b_1 _09223_ (.A(_01718_),
    .B_N(_01721_),
    .Y(_01722_));
 sg13g2_and4_1 _09224_ (.A(_01690_),
    .B(_01714_),
    .C(_01716_),
    .D(_01722_),
    .X(_01723_));
 sg13g2_buf_2 _09225_ (.A(_01723_),
    .X(_01724_));
 sg13g2_buf_1 _09226_ (.A(\clock_inst.hour_tile.e[9] ),
    .X(_01725_));
 sg13g2_and2_1 _09227_ (.A(\clock_inst.vga_inst.vga_horizontal_visible ),
    .B(\clock_inst.vga_inst.vga_vertical_visible ),
    .X(_01726_));
 sg13g2_buf_1 _09228_ (.A(_01726_),
    .X(_01727_));
 sg13g2_buf_1 _09229_ (.A(_01727_),
    .X(_01728_));
 sg13g2_buf_1 _09230_ (.A(\clock_inst.hour_tile.e[8] ),
    .X(_01729_));
 sg13g2_nor2b_1 _09231_ (.A(_00686_),
    .B_N(_01729_),
    .Y(_01730_));
 sg13g2_and2_1 _09232_ (.A(net500),
    .B(_01730_),
    .X(_01731_));
 sg13g2_nand2_1 _09233_ (.Y(_01732_),
    .A(_01725_),
    .B(_01731_));
 sg13g2_nand2b_1 _09234_ (.Y(_01733_),
    .B(_00686_),
    .A_N(_01729_));
 sg13g2_nor2_1 _09235_ (.A(net542),
    .B(_01733_),
    .Y(_01734_));
 sg13g2_nand3b_1 _09236_ (.B(_01724_),
    .C(_01734_),
    .Y(_01735_),
    .A_N(net572));
 sg13g2_o21ai_1 _09237_ (.B1(_01735_),
    .Y(_01736_),
    .A1(_01724_),
    .A2(_01732_));
 sg13g2_xnor2_1 _09238_ (.Y(_01737_),
    .A(_01688_),
    .B(_01736_));
 sg13g2_a21oi_1 _09239_ (.A1(net79),
    .A2(_01737_),
    .Y(_00153_),
    .B1(_01123_));
 sg13g2_buf_1 _09240_ (.A(\clock_inst.hour_tile.e[11] ),
    .X(_01738_));
 sg13g2_nand4_1 _09241_ (.B(_01714_),
    .C(_01716_),
    .A(_01690_),
    .Y(_01739_),
    .D(_01722_));
 sg13g2_buf_2 _09242_ (.A(_01739_),
    .X(_01740_));
 sg13g2_or4_1 _09243_ (.A(net572),
    .B(_01688_),
    .C(_01740_),
    .D(_01733_),
    .X(_01741_));
 sg13g2_nand4_1 _09244_ (.B(_01688_),
    .C(_01740_),
    .A(net572),
    .Y(_01742_),
    .D(_01730_));
 sg13g2_buf_1 _09245_ (.A(net502),
    .X(_01743_));
 sg13g2_a21oi_1 _09246_ (.A1(_01741_),
    .A2(_01742_),
    .Y(_01744_),
    .B1(_01743_));
 sg13g2_xnor2_1 _09247_ (.Y(_01745_),
    .A(_01738_),
    .B(_01744_));
 sg13g2_a21oi_1 _09248_ (.A1(net79),
    .A2(_01745_),
    .Y(_00154_),
    .B1(_01132_));
 sg13g2_buf_1 _09249_ (.A(net236),
    .X(_01746_));
 sg13g2_buf_1 _09250_ (.A(\clock_inst.hour_tile.e[12] ),
    .X(_01747_));
 sg13g2_or4_1 _09251_ (.A(net572),
    .B(_01688_),
    .C(_01738_),
    .D(_01733_),
    .X(_01748_));
 sg13g2_buf_1 _09252_ (.A(_01748_),
    .X(_01749_));
 sg13g2_nor3_2 _09253_ (.A(net542),
    .B(_01740_),
    .C(_01749_),
    .Y(_01750_));
 sg13g2_and4_1 _09254_ (.A(net572),
    .B(_01688_),
    .C(_01738_),
    .D(_01730_),
    .X(_01751_));
 sg13g2_nand2_1 _09255_ (.Y(_01752_),
    .A(net500),
    .B(_01751_));
 sg13g2_nor2_1 _09256_ (.A(_01724_),
    .B(_01752_),
    .Y(_01753_));
 sg13g2_nor2_1 _09257_ (.A(_01750_),
    .B(_01753_),
    .Y(_01754_));
 sg13g2_xor2_1 _09258_ (.B(_01754_),
    .A(_01747_),
    .X(_01755_));
 sg13g2_o21ai_1 _09259_ (.B1(_01148_),
    .Y(_00155_),
    .A1(_01746_),
    .A2(_01755_));
 sg13g2_buf_1 _09260_ (.A(\clock_inst.hour_tile.e[13] ),
    .X(_01756_));
 sg13g2_mux2_1 _09261_ (.A0(_01750_),
    .A1(_01753_),
    .S(_01747_),
    .X(_01757_));
 sg13g2_xnor2_1 _09262_ (.Y(_01758_),
    .A(_01756_),
    .B(_01757_));
 sg13g2_a21oi_1 _09263_ (.A1(net79),
    .A2(_01758_),
    .Y(_00156_),
    .B1(_01164_));
 sg13g2_buf_1 _09264_ (.A(\clock_inst.hour_tile.e[14] ),
    .X(_01759_));
 sg13g2_inv_1 _09265_ (.Y(_01760_),
    .A(_00686_));
 sg13g2_a221oi_1 _09266_ (.B2(_01711_),
    .C1(_01706_),
    .B1(_00806_),
    .A1(\clock_inst.hour_tile.e[4] ),
    .Y(_01761_),
    .A2(_00964_));
 sg13g2_buf_1 _09267_ (.A(_01761_),
    .X(_01762_));
 sg13g2_nand4_1 _09268_ (.B(_01688_),
    .C(_01738_),
    .A(net572),
    .Y(_01763_),
    .D(_01730_));
 sg13g2_nand2_1 _09269_ (.Y(_01764_),
    .A(_01749_),
    .B(_01763_));
 sg13g2_xor2_1 _09270_ (.B(_01708_),
    .A(_00813_),
    .X(_01765_));
 sg13g2_nand4_1 _09271_ (.B(_01719_),
    .C(_01764_),
    .A(_01690_),
    .Y(_01766_),
    .D(_01765_));
 sg13g2_nor3_1 _09272_ (.A(_01712_),
    .B(_01762_),
    .C(_01766_),
    .Y(_01767_));
 sg13g2_a21oi_1 _09273_ (.A1(_01690_),
    .A2(_01717_),
    .Y(_01768_),
    .B1(_01710_));
 sg13g2_nand4_1 _09274_ (.B(_01688_),
    .C(_01738_),
    .A(net572),
    .Y(_01769_),
    .D(_01768_));
 sg13g2_or4_1 _09275_ (.A(net572),
    .B(_01688_),
    .C(_01738_),
    .D(_01768_),
    .X(_01770_));
 sg13g2_a21oi_1 _09276_ (.A1(_00686_),
    .A2(_01770_),
    .Y(_01771_),
    .B1(_01729_));
 sg13g2_a21oi_1 _09277_ (.A1(_01760_),
    .A2(_01769_),
    .Y(_01772_),
    .B1(_01771_));
 sg13g2_or2_1 _09278_ (.X(_01773_),
    .B(_01756_),
    .A(_01747_));
 sg13g2_buf_1 _09279_ (.A(_01773_),
    .X(_01774_));
 sg13g2_or4_1 _09280_ (.A(_01760_),
    .B(_01767_),
    .C(_01772_),
    .D(_01774_),
    .X(_01775_));
 sg13g2_and3_1 _09281_ (.X(_01776_),
    .A(_01760_),
    .B(_01747_),
    .C(_01756_));
 sg13g2_o21ai_1 _09282_ (.B1(_01776_),
    .Y(_01777_),
    .A1(_01767_),
    .A2(_01772_));
 sg13g2_buf_1 _09283_ (.A(net502),
    .X(_01778_));
 sg13g2_a21oi_1 _09284_ (.A1(_01775_),
    .A2(_01777_),
    .Y(_01779_),
    .B1(_01778_));
 sg13g2_xnor2_1 _09285_ (.Y(_01780_),
    .A(_01759_),
    .B(_01779_));
 sg13g2_o21ai_1 _09286_ (.B1(_01174_),
    .Y(_00157_),
    .A1(_01746_),
    .A2(_01780_));
 sg13g2_inv_1 _09287_ (.Y(_01781_),
    .A(\clock_inst.hour_tile.e[15] ));
 sg13g2_nor2_1 _09288_ (.A(_01759_),
    .B(_01774_),
    .Y(_01782_));
 sg13g2_nand3_1 _09289_ (.B(_01756_),
    .C(_01759_),
    .A(_01747_),
    .Y(_01783_));
 sg13g2_nor2_1 _09290_ (.A(_01752_),
    .B(_01783_),
    .Y(_01784_));
 sg13g2_a22oi_1 _09291_ (.Y(_01785_),
    .B1(_01784_),
    .B2(_01740_),
    .A2(_01782_),
    .A1(_01750_));
 sg13g2_xnor2_1 _09292_ (.Y(_01786_),
    .A(_01781_),
    .B(_01785_));
 sg13g2_buf_1 _09293_ (.A(_01409_),
    .X(_01787_));
 sg13g2_a22oi_1 _09294_ (.Y(_00158_),
    .B1(_01786_),
    .B2(_01787_),
    .A2(_01187_),
    .A1(_01185_));
 sg13g2_nor3_1 _09295_ (.A(_01781_),
    .B(_01752_),
    .C(_01783_),
    .Y(_01788_));
 sg13g2_nor3_1 _09296_ (.A(_01759_),
    .B(\clock_inst.hour_tile.e[15] ),
    .C(_01774_),
    .Y(_01789_));
 sg13g2_a22oi_1 _09297_ (.Y(_01790_),
    .B1(_01789_),
    .B2(_01750_),
    .A2(_01788_),
    .A1(_01740_));
 sg13g2_xor2_1 _09298_ (.B(_01790_),
    .A(\clock_inst.hour_tile.e[16] ),
    .X(_01791_));
 sg13g2_a21oi_1 _09299_ (.A1(net79),
    .A2(_01791_),
    .Y(_00159_),
    .B1(_01199_));
 sg13g2_nand2b_1 _09300_ (.Y(_01792_),
    .B(_01782_),
    .A_N(\clock_inst.hour_tile.e[16] ));
 sg13g2_nor4_1 _09301_ (.A(\clock_inst.hour_tile.e[15] ),
    .B(_01740_),
    .C(_01749_),
    .D(_01792_),
    .Y(_01793_));
 sg13g2_nand2_1 _09302_ (.Y(_01794_),
    .A(\clock_inst.hour_tile.e[16] ),
    .B(_01751_));
 sg13g2_nor4_1 _09303_ (.A(_01781_),
    .B(_01724_),
    .C(_01783_),
    .D(_01794_),
    .Y(_01795_));
 sg13g2_buf_1 _09304_ (.A(net500),
    .X(_01796_));
 sg13g2_buf_1 _09305_ (.A(net445),
    .X(_01797_));
 sg13g2_o21ai_1 _09306_ (.B1(_01797_),
    .Y(_01798_),
    .A1(_01793_),
    .A2(_01795_));
 sg13g2_xor2_1 _09307_ (.B(_01798_),
    .A(\clock_inst.hour_tile.e[17] ),
    .X(_01799_));
 sg13g2_a22oi_1 _09308_ (.Y(_00160_),
    .B1(_01799_),
    .B2(net78),
    .A2(_01211_),
    .A1(_01209_));
 sg13g2_buf_2 _09309_ (.A(\clock_inst.hour_tile.e[18] ),
    .X(_01800_));
 sg13g2_nor2_1 _09310_ (.A(_01800_),
    .B(net80),
    .Y(_01801_));
 sg13g2_nor2_2 _09311_ (.A(_01057_),
    .B(net502),
    .Y(_01802_));
 sg13g2_a22oi_1 _09312_ (.Y(_01803_),
    .B1(_01802_),
    .B2(_01800_),
    .A2(net49),
    .A1(_01214_));
 sg13g2_nor2b_1 _09313_ (.A(_01803_),
    .B_N(net575),
    .Y(_01804_));
 sg13g2_nor2_1 _09314_ (.A(net239),
    .B(net237),
    .Y(_01805_));
 sg13g2_a221oi_1 _09315_ (.B2(_01214_),
    .C1(net575),
    .B1(_01805_),
    .A1(_01800_),
    .Y(_01806_),
    .A2(_01152_));
 sg13g2_nor3_1 _09316_ (.A(_01801_),
    .B(_01804_),
    .C(_01806_),
    .Y(_00161_));
 sg13g2_nand2_1 _09317_ (.Y(_01807_),
    .A(_00925_),
    .B(_01800_));
 sg13g2_xnor2_1 _09318_ (.Y(_01808_),
    .A(_00693_),
    .B(_01807_));
 sg13g2_nor2_1 _09319_ (.A(net448),
    .B(_01808_),
    .Y(_01809_));
 sg13g2_xnor2_1 _09320_ (.Y(_01810_),
    .A(\clock_inst.hour_tile.e[19] ),
    .B(_01809_));
 sg13g2_a21oi_1 _09321_ (.A1(_01687_),
    .A2(_01810_),
    .Y(_00162_),
    .B1(_01228_));
 sg13g2_buf_1 _09322_ (.A(net501),
    .X(_01811_));
 sg13g2_xnor2_1 _09323_ (.Y(_01812_),
    .A(_00701_),
    .B(_01683_));
 sg13g2_nor2_1 _09324_ (.A(net444),
    .B(_01812_),
    .Y(_01813_));
 sg13g2_xnor2_1 _09325_ (.Y(_01814_),
    .A(\clock_inst.hour_tile.e[1] ),
    .B(_01813_));
 sg13g2_a21oi_1 _09326_ (.A1(_01687_),
    .A2(_01814_),
    .Y(_00163_),
    .B1(_01236_));
 sg13g2_buf_1 _09327_ (.A(_01727_),
    .X(_01815_));
 sg13g2_buf_1 _09328_ (.A(net499),
    .X(_01816_));
 sg13g2_nor2_1 _09329_ (.A(\clock_inst.hour_a[19] ),
    .B(\clock_inst.hour_tile.e[19] ),
    .Y(_01817_));
 sg13g2_a22oi_1 _09330_ (.Y(_01818_),
    .B1(_01800_),
    .B2(net575),
    .A2(\clock_inst.hour_tile.e[19] ),
    .A1(\clock_inst.hour_a[19] ));
 sg13g2_nor2_1 _09331_ (.A(_01817_),
    .B(_01818_),
    .Y(_01819_));
 sg13g2_xnor2_1 _09332_ (.Y(_01820_),
    .A(_00711_),
    .B(_01819_));
 sg13g2_nand2_1 _09333_ (.Y(_01821_),
    .A(net443),
    .B(_01820_));
 sg13g2_xnor2_1 _09334_ (.Y(_01822_),
    .A(\clock_inst.hour_tile.e[20] ),
    .B(_01821_));
 sg13g2_xor2_1 _09335_ (.B(_01245_),
    .A(_01237_),
    .X(_01823_));
 sg13g2_a22oi_1 _09336_ (.Y(_01824_),
    .B1(_01823_),
    .B2(net23),
    .A2(_01822_),
    .A1(net83));
 sg13g2_inv_1 _09337_ (.Y(_00164_),
    .A(_01824_));
 sg13g2_and2_1 _09338_ (.A(\clock_inst.hour_a[20] ),
    .B(\clock_inst.hour_tile.e[20] ),
    .X(_01825_));
 sg13g2_buf_1 _09339_ (.A(_01825_),
    .X(_01826_));
 sg13g2_nor2_1 _09340_ (.A(\clock_inst.hour_a[20] ),
    .B(\clock_inst.hour_tile.e[20] ),
    .Y(_01827_));
 sg13g2_nor3_2 _09341_ (.A(_01817_),
    .B(_01818_),
    .C(_01827_),
    .Y(_01828_));
 sg13g2_o21ai_1 _09342_ (.B1(\clock_inst.hour_a[21] ),
    .Y(_01829_),
    .A1(_01826_),
    .A2(_01828_));
 sg13g2_or3_1 _09343_ (.A(\clock_inst.hour_a[21] ),
    .B(_01826_),
    .C(_01828_),
    .X(_01830_));
 sg13g2_and3_1 _09344_ (.X(_01831_),
    .A(net443),
    .B(_01829_),
    .C(_01830_));
 sg13g2_xnor2_1 _09345_ (.Y(_01832_),
    .A(\clock_inst.hour_tile.e[21] ),
    .B(_01831_));
 sg13g2_a21oi_1 _09346_ (.A1(net79),
    .A2(_01832_),
    .Y(_00165_),
    .B1(_01261_));
 sg13g2_inv_1 _09347_ (.Y(_01833_),
    .A(\clock_inst.hour_tile.e[22] ));
 sg13g2_inv_1 _09348_ (.Y(_01834_),
    .A(\clock_inst.hour_tile.e[21] ));
 sg13g2_nand2_1 _09349_ (.Y(_01835_),
    .A(_00721_),
    .B(_01834_));
 sg13g2_o21ai_1 _09350_ (.B1(_01835_),
    .Y(_01836_),
    .A1(_01826_),
    .A2(_01828_));
 sg13g2_buf_2 _09351_ (.A(_01836_),
    .X(_01837_));
 sg13g2_o21ai_1 _09352_ (.B1(_01837_),
    .Y(_01838_),
    .A1(_00721_),
    .A2(_01834_));
 sg13g2_xnor2_1 _09353_ (.Y(_01839_),
    .A(_00724_),
    .B(_01838_));
 sg13g2_nor2_1 _09354_ (.A(_01778_),
    .B(_01839_),
    .Y(_01840_));
 sg13g2_xnor2_1 _09355_ (.Y(_01841_),
    .A(_01833_),
    .B(_01840_));
 sg13g2_xnor2_1 _09356_ (.Y(_01842_),
    .A(_01262_),
    .B(_01271_));
 sg13g2_nor2_1 _09357_ (.A(net44),
    .B(_01842_),
    .Y(_01843_));
 sg13g2_a21o_1 _09358_ (.A2(_01841_),
    .A1(net112),
    .B1(_01843_),
    .X(_00166_));
 sg13g2_buf_1 _09359_ (.A(net140),
    .X(_01844_));
 sg13g2_buf_1 _09360_ (.A(\clock_inst.hour_tile.e[23] ),
    .X(_01845_));
 sg13g2_a22oi_1 _09361_ (.Y(_01846_),
    .B1(\clock_inst.hour_a[21] ),
    .B2(\clock_inst.hour_tile.e[21] ),
    .A2(_00724_),
    .A1(\clock_inst.hour_tile.e[22] ));
 sg13g2_buf_1 _09362_ (.A(_01846_),
    .X(_01847_));
 sg13g2_a22oi_1 _09363_ (.Y(_01848_),
    .B1(_01837_),
    .B2(_01847_),
    .A2(_00725_),
    .A1(_01833_));
 sg13g2_xnor2_1 _09364_ (.Y(_01849_),
    .A(net546),
    .B(_01848_));
 sg13g2_nor2_1 _09365_ (.A(net444),
    .B(_01849_),
    .Y(_01850_));
 sg13g2_xnor2_1 _09366_ (.Y(_01851_),
    .A(_01845_),
    .B(_01850_));
 sg13g2_a21oi_1 _09367_ (.A1(net77),
    .A2(_01851_),
    .Y(_00167_),
    .B1(_01287_));
 sg13g2_buf_1 _09368_ (.A(\clock_inst.hour_tile.e[24] ),
    .X(_01852_));
 sg13g2_nand2_1 _09369_ (.Y(_01853_),
    .A(_01833_),
    .B(_00725_));
 sg13g2_nand2_1 _09370_ (.Y(_01854_),
    .A(_01845_),
    .B(_01853_));
 sg13g2_a21oi_1 _09371_ (.A1(_01837_),
    .A2(_01847_),
    .Y(_01855_),
    .B1(_01854_));
 sg13g2_nand2_1 _09372_ (.Y(_01856_),
    .A(_00732_),
    .B(_01853_));
 sg13g2_a21oi_1 _09373_ (.A1(_01837_),
    .A2(_01847_),
    .Y(_01857_),
    .B1(_01856_));
 sg13g2_and2_1 _09374_ (.A(_00731_),
    .B(_01845_),
    .X(_01858_));
 sg13g2_buf_1 _09375_ (.A(_01858_),
    .X(_01859_));
 sg13g2_or3_1 _09376_ (.A(_01855_),
    .B(_01857_),
    .C(_01859_),
    .X(_01860_));
 sg13g2_buf_2 _09377_ (.A(_01860_),
    .X(_01861_));
 sg13g2_xnor2_1 _09378_ (.Y(_01862_),
    .A(net579),
    .B(_01861_));
 sg13g2_nor2_1 _09379_ (.A(net444),
    .B(_01862_),
    .Y(_01863_));
 sg13g2_xnor2_1 _09380_ (.Y(_01864_),
    .A(_01852_),
    .B(_01863_));
 sg13g2_a21oi_1 _09381_ (.A1(net77),
    .A2(_01864_),
    .Y(_00168_),
    .B1(_01307_));
 sg13g2_buf_2 _09382_ (.A(\clock_inst.hour_tile.e[25] ),
    .X(_01865_));
 sg13g2_nor2b_1 _09383_ (.A(net579),
    .B_N(_01852_),
    .Y(_01866_));
 sg13g2_nand2b_1 _09384_ (.Y(_01867_),
    .B(net579),
    .A_N(_01852_));
 sg13g2_nor2_1 _09385_ (.A(_01861_),
    .B(_01867_),
    .Y(_01868_));
 sg13g2_a21oi_1 _09386_ (.A1(_01861_),
    .A2(_01866_),
    .Y(_01869_),
    .B1(_01868_));
 sg13g2_nor2_1 _09387_ (.A(net444),
    .B(_01869_),
    .Y(_01870_));
 sg13g2_xnor2_1 _09388_ (.Y(_01871_),
    .A(_01865_),
    .B(_01870_));
 sg13g2_a21oi_1 _09389_ (.A1(net77),
    .A2(_01871_),
    .Y(_00169_),
    .B1(_01317_));
 sg13g2_buf_2 _09390_ (.A(\clock_inst.hour_tile.e[26] ),
    .X(_01872_));
 sg13g2_or3_1 _09391_ (.A(_01865_),
    .B(_01861_),
    .C(_01867_),
    .X(_01873_));
 sg13g2_nand3_1 _09392_ (.B(_01861_),
    .C(_01866_),
    .A(_01865_),
    .Y(_01874_));
 sg13g2_a21oi_1 _09393_ (.A1(_01873_),
    .A2(_01874_),
    .Y(_01875_),
    .B1(net447));
 sg13g2_xnor2_1 _09394_ (.Y(_01876_),
    .A(_01872_),
    .B(_01875_));
 sg13g2_a21oi_1 _09395_ (.A1(net77),
    .A2(_01876_),
    .Y(_00170_),
    .B1(_01330_));
 sg13g2_buf_1 _09396_ (.A(\clock_inst.hour_tile.e[27] ),
    .X(_01877_));
 sg13g2_nand4_1 _09397_ (.B(_01865_),
    .C(_01872_),
    .A(_01845_),
    .Y(_01878_),
    .D(_01853_));
 sg13g2_nand4_1 _09398_ (.B(_01865_),
    .C(_01872_),
    .A(net546),
    .Y(_01879_),
    .D(_01853_));
 sg13g2_a22oi_1 _09399_ (.Y(_01880_),
    .B1(_01878_),
    .B2(_01879_),
    .A2(_01847_),
    .A1(_01837_));
 sg13g2_nand3_1 _09400_ (.B(_01872_),
    .C(_01859_),
    .A(_01865_),
    .Y(_01881_));
 sg13g2_nand2b_1 _09401_ (.Y(_01882_),
    .B(_01881_),
    .A_N(_01880_));
 sg13g2_buf_2 _09402_ (.A(_01882_),
    .X(_01883_));
 sg13g2_nor4_2 _09403_ (.A(_01865_),
    .B(_01872_),
    .C(_01861_),
    .Y(_01884_),
    .D(_01867_));
 sg13g2_a21oi_1 _09404_ (.A1(_01866_),
    .A2(_01883_),
    .Y(_01885_),
    .B1(_01884_));
 sg13g2_nor2_1 _09405_ (.A(net444),
    .B(_01885_),
    .Y(_01886_));
 sg13g2_xnor2_1 _09406_ (.Y(_01887_),
    .A(_01877_),
    .B(_01886_));
 sg13g2_a21oi_1 _09407_ (.A1(net77),
    .A2(_01887_),
    .Y(_00171_),
    .B1(_01337_));
 sg13g2_buf_1 _09408_ (.A(\clock_inst.hour_tile.e[28] ),
    .X(_01888_));
 sg13g2_inv_1 _09409_ (.Y(_01889_),
    .A(_01877_));
 sg13g2_nand2_1 _09410_ (.Y(_01890_),
    .A(_01546_),
    .B(_01852_));
 sg13g2_nor2_1 _09411_ (.A(_01889_),
    .B(_01890_),
    .Y(_01891_));
 sg13g2_a22oi_1 _09412_ (.Y(_01892_),
    .B1(_01883_),
    .B2(_01891_),
    .A2(_01884_),
    .A1(_01889_));
 sg13g2_nor2_1 _09413_ (.A(net444),
    .B(_01892_),
    .Y(_01893_));
 sg13g2_xnor2_1 _09414_ (.Y(_01894_),
    .A(_01888_),
    .B(_01893_));
 sg13g2_a21oi_1 _09415_ (.A1(net77),
    .A2(_01894_),
    .Y(_00172_),
    .B1(_01348_));
 sg13g2_buf_1 _09416_ (.A(\clock_inst.hour_tile.e[29] ),
    .X(_01895_));
 sg13g2_nor4_1 _09417_ (.A(_01852_),
    .B(_01865_),
    .C(_01872_),
    .D(_01877_),
    .Y(_01896_));
 sg13g2_nand2b_1 _09418_ (.Y(_01897_),
    .B(_01896_),
    .A_N(_01888_));
 sg13g2_nor4_2 _09419_ (.A(_01855_),
    .B(_01857_),
    .C(_01859_),
    .Y(_01898_),
    .D(_01897_));
 sg13g2_and3_1 _09420_ (.X(_01899_),
    .A(_01852_),
    .B(_01877_),
    .C(_01888_));
 sg13g2_buf_1 _09421_ (.A(_01899_),
    .X(_01900_));
 sg13g2_and2_1 _09422_ (.A(_01546_),
    .B(_01900_),
    .X(_01901_));
 sg13g2_a22oi_1 _09423_ (.Y(_01902_),
    .B1(_01901_),
    .B2(_01883_),
    .A2(_01898_),
    .A1(net579));
 sg13g2_nor2_1 _09424_ (.A(net501),
    .B(_01902_),
    .Y(_01903_));
 sg13g2_xor2_1 _09425_ (.B(_01903_),
    .A(_01895_),
    .X(_01904_));
 sg13g2_a21o_1 _09426_ (.A2(_01904_),
    .A1(_01034_),
    .B1(_01358_),
    .X(_00173_));
 sg13g2_xnor2_1 _09427_ (.Y(_01905_),
    .A(_00741_),
    .B(_01698_));
 sg13g2_nor2_1 _09428_ (.A(net444),
    .B(_01905_),
    .Y(_01906_));
 sg13g2_xnor2_1 _09429_ (.Y(_01907_),
    .A(_01693_),
    .B(_01906_));
 sg13g2_a21oi_1 _09430_ (.A1(net77),
    .A2(_01907_),
    .Y(_00174_),
    .B1(_01365_));
 sg13g2_buf_1 _09431_ (.A(\clock_inst.hour_tile.e[30] ),
    .X(_01908_));
 sg13g2_nand4_1 _09432_ (.B(_01895_),
    .C(_01883_),
    .A(_01546_),
    .Y(_01909_),
    .D(_01900_));
 sg13g2_nand3b_1 _09433_ (.B(_01898_),
    .C(net579),
    .Y(_01910_),
    .A_N(_01895_));
 sg13g2_a21oi_1 _09434_ (.A1(_01909_),
    .A2(_01910_),
    .Y(_01911_),
    .B1(net446));
 sg13g2_xor2_1 _09435_ (.B(_01911_),
    .A(_01908_),
    .X(_01912_));
 sg13g2_buf_1 _09436_ (.A(net143),
    .X(_01913_));
 sg13g2_mux2_1 _09437_ (.A0(_01379_),
    .A1(_01912_),
    .S(net76),
    .X(_00175_));
 sg13g2_buf_1 _09438_ (.A(_01061_),
    .X(_01914_));
 sg13g2_buf_2 _09439_ (.A(\clock_inst.hour_tile.e[31] ),
    .X(_01915_));
 sg13g2_nor2b_1 _09440_ (.A(net579),
    .B_N(_01908_),
    .Y(_01916_));
 sg13g2_nand4_1 _09441_ (.B(_01883_),
    .C(_01900_),
    .A(_01895_),
    .Y(_01917_),
    .D(_01916_));
 sg13g2_nor2_1 _09442_ (.A(_01877_),
    .B(_01888_),
    .Y(_01918_));
 sg13g2_nor2_1 _09443_ (.A(_01895_),
    .B(_01908_),
    .Y(_01919_));
 sg13g2_nand3_1 _09444_ (.B(_01918_),
    .C(_01919_),
    .A(_01884_),
    .Y(_01920_));
 sg13g2_a21oi_1 _09445_ (.A1(_01917_),
    .A2(_01920_),
    .Y(_01921_),
    .B1(net447));
 sg13g2_xnor2_1 _09446_ (.Y(_01922_),
    .A(_01915_),
    .B(_01921_));
 sg13g2_xnor2_1 _09447_ (.Y(_01923_),
    .A(_01386_),
    .B(_01385_));
 sg13g2_nand2_1 _09448_ (.Y(_01924_),
    .A(net45),
    .B(_01923_));
 sg13g2_buf_1 _09449_ (.A(net96),
    .X(_01925_));
 sg13g2_buf_1 _09450_ (.A(net242),
    .X(_01926_));
 sg13g2_a21oi_1 _09451_ (.A1(_00964_),
    .A2(net43),
    .Y(_01927_),
    .B1(net138));
 sg13g2_a22oi_1 _09452_ (.Y(_00176_),
    .B1(_01924_),
    .B2(_01927_),
    .A2(_01922_),
    .A1(net75));
 sg13g2_buf_1 _09453_ (.A(\clock_inst.hour_tile.e[32] ),
    .X(_01928_));
 sg13g2_nor2_1 _09454_ (.A(_01677_),
    .B(_01917_),
    .Y(_01929_));
 sg13g2_nand4_1 _09455_ (.B(net500),
    .C(_01898_),
    .A(net579),
    .Y(_01930_),
    .D(_01919_));
 sg13g2_nor2_1 _09456_ (.A(_01915_),
    .B(_01930_),
    .Y(_01931_));
 sg13g2_a21oi_1 _09457_ (.A1(_01915_),
    .A2(_01929_),
    .Y(_01932_),
    .B1(_01931_));
 sg13g2_xor2_1 _09458_ (.B(_01932_),
    .A(_01928_),
    .X(_01933_));
 sg13g2_xnor2_1 _09459_ (.Y(_01934_),
    .A(_01392_),
    .B(_01394_));
 sg13g2_nand2_1 _09460_ (.Y(_01935_),
    .A(net152),
    .B(_01934_));
 sg13g2_a21oi_1 _09461_ (.A1(\clock_inst.hour_c[32] ),
    .A2(net43),
    .Y(_01936_),
    .B1(net138));
 sg13g2_a22oi_1 _09462_ (.Y(_00177_),
    .B1(_01935_),
    .B2(_01936_),
    .A2(_01933_),
    .A1(net75));
 sg13g2_nand2_1 _09463_ (.Y(_01937_),
    .A(_01915_),
    .B(_01928_));
 sg13g2_nor2_1 _09464_ (.A(_01898_),
    .B(_01937_),
    .Y(_01938_));
 sg13g2_nor3_1 _09465_ (.A(_01915_),
    .B(_01928_),
    .C(_01930_),
    .Y(_01939_));
 sg13g2_a21oi_1 _09466_ (.A1(_01929_),
    .A2(_01938_),
    .Y(_01940_),
    .B1(_01939_));
 sg13g2_xor2_1 _09467_ (.B(_01940_),
    .A(\clock_inst.hour_tile.e[33] ),
    .X(_01941_));
 sg13g2_a21oi_1 _09468_ (.A1(net77),
    .A2(_01941_),
    .Y(_00178_),
    .B1(_01407_));
 sg13g2_buf_1 _09469_ (.A(\clock_inst.hour_tile.e[34] ),
    .X(_01942_));
 sg13g2_nor2_1 _09470_ (.A(_01942_),
    .B(_01679_),
    .Y(_01943_));
 sg13g2_nand2_1 _09471_ (.Y(_01944_),
    .A(_01426_),
    .B(_01429_));
 sg13g2_nor3_1 _09472_ (.A(_01908_),
    .B(_01915_),
    .C(_01928_),
    .Y(_01945_));
 sg13g2_nor3_1 _09473_ (.A(_01888_),
    .B(_01895_),
    .C(\clock_inst.hour_tile.e[33] ),
    .Y(_01946_));
 sg13g2_and4_1 _09474_ (.A(_01889_),
    .B(_01884_),
    .C(_01945_),
    .D(_01946_),
    .X(_01947_));
 sg13g2_nand3_1 _09475_ (.B(_01928_),
    .C(\clock_inst.hour_tile.e[33] ),
    .A(_01915_),
    .Y(_01948_));
 sg13g2_nor2_1 _09476_ (.A(_01917_),
    .B(_01948_),
    .Y(_01949_));
 sg13g2_nor4_1 _09477_ (.A(_01942_),
    .B(_01413_),
    .C(_01947_),
    .D(_01949_),
    .Y(_01950_));
 sg13g2_nor2b_1 _09478_ (.A(_01944_),
    .B_N(_01950_),
    .Y(_01951_));
 sg13g2_and2_1 _09479_ (.A(_01942_),
    .B(net500),
    .X(_01952_));
 sg13g2_and4_1 _09480_ (.A(_01889_),
    .B(_01945_),
    .C(_01946_),
    .D(_01952_),
    .X(_01953_));
 sg13g2_a221oi_1 _09481_ (.B2(_01884_),
    .C1(net240),
    .B1(_01953_),
    .A1(_01949_),
    .Y(_01954_),
    .A2(_01952_));
 sg13g2_nor3_1 _09482_ (.A(_01413_),
    .B(_01944_),
    .C(_01954_),
    .Y(_01955_));
 sg13g2_nor3_1 _09483_ (.A(_01943_),
    .B(_01951_),
    .C(_01955_),
    .Y(_00179_));
 sg13g2_inv_1 _09484_ (.Y(_01956_),
    .A(\clock_inst.hour_tile.e[35] ));
 sg13g2_mux2_1 _09485_ (.A0(_01947_),
    .A1(_01949_),
    .S(_01942_),
    .X(_01957_));
 sg13g2_o21ai_1 _09486_ (.B1(net80),
    .Y(_01958_),
    .A1(_01437_),
    .A2(_01957_));
 sg13g2_nor2_1 _09487_ (.A(_01956_),
    .B(_01682_),
    .Y(_01959_));
 sg13g2_a21o_1 _09488_ (.A2(_01959_),
    .A1(_01957_),
    .B1(_01641_),
    .X(_01960_));
 sg13g2_a21o_1 _09489_ (.A2(_01436_),
    .A1(_01405_),
    .B1(net160),
    .X(_01961_));
 sg13g2_a22oi_1 _09490_ (.Y(_00180_),
    .B1(_01960_),
    .B2(_01961_),
    .A2(_01958_),
    .A1(_01956_));
 sg13g2_inv_1 _09491_ (.Y(_01962_),
    .A(\clock_inst.hour_tile.e[36] ));
 sg13g2_o21ai_1 _09492_ (.B1(net80),
    .Y(_01963_),
    .A1(\clock_inst.hour_a[36] ),
    .A2(_01440_));
 sg13g2_buf_1 _09493_ (.A(net499),
    .X(_01964_));
 sg13g2_buf_1 _09494_ (.A(_01964_),
    .X(_01965_));
 sg13g2_and2_1 _09495_ (.A(\clock_inst.hour_a[36] ),
    .B(\clock_inst.hour_tile.e[36] ),
    .X(_01966_));
 sg13g2_buf_1 _09496_ (.A(_01966_),
    .X(_01967_));
 sg13g2_a21oi_1 _09497_ (.A1(net356),
    .A2(_01967_),
    .Y(_01968_),
    .B1(_01248_));
 sg13g2_nor2_1 _09498_ (.A(_01440_),
    .B(_01968_),
    .Y(_01969_));
 sg13g2_a21oi_1 _09499_ (.A1(_01962_),
    .A2(_01963_),
    .Y(_00181_),
    .B1(_01969_));
 sg13g2_xnor2_1 _09500_ (.Y(_01970_),
    .A(_00762_),
    .B(_01967_));
 sg13g2_nor2_1 _09501_ (.A(_01811_),
    .B(_01970_),
    .Y(_01971_));
 sg13g2_xnor2_1 _09502_ (.Y(_01972_),
    .A(\clock_inst.hour_tile.e[37] ),
    .B(_01971_));
 sg13g2_a21oi_1 _09503_ (.A1(_01844_),
    .A2(_01972_),
    .Y(_00182_),
    .B1(_01449_));
 sg13g2_or2_1 _09504_ (.X(_01973_),
    .B(\clock_inst.hour_tile.e[37] ),
    .A(_00762_));
 sg13g2_and2_1 _09505_ (.A(_00762_),
    .B(\clock_inst.hour_tile.e[37] ),
    .X(_01974_));
 sg13g2_a21oi_1 _09506_ (.A1(_01967_),
    .A2(_01973_),
    .Y(_01975_),
    .B1(_01974_));
 sg13g2_xnor2_1 _09507_ (.Y(_01976_),
    .A(_00770_),
    .B(_01975_));
 sg13g2_nor2_1 _09508_ (.A(_01811_),
    .B(_01976_),
    .Y(_01977_));
 sg13g2_xnor2_1 _09509_ (.Y(_01978_),
    .A(\clock_inst.hour_tile.e[38] ),
    .B(_01977_));
 sg13g2_a21oi_1 _09510_ (.A1(_01844_),
    .A2(_01978_),
    .Y(_00183_),
    .B1(_01457_));
 sg13g2_xnor2_1 _09511_ (.Y(_01979_),
    .A(_01459_),
    .B(_01468_));
 sg13g2_nor2_1 _09512_ (.A(_01247_),
    .B(_01979_),
    .Y(_01980_));
 sg13g2_a21oi_1 _09513_ (.A1(\clock_inst.hour_c[2] ),
    .A2(_01393_),
    .Y(_01981_),
    .B1(_01980_));
 sg13g2_a221oi_1 _09514_ (.B2(_01973_),
    .C1(_01974_),
    .B1(_01967_),
    .A1(\clock_inst.hour_a[38] ),
    .Y(_01982_),
    .A2(\clock_inst.hour_tile.e[38] ));
 sg13g2_buf_1 _09515_ (.A(_01982_),
    .X(_01983_));
 sg13g2_nor2_2 _09516_ (.A(\clock_inst.hour_a[38] ),
    .B(\clock_inst.hour_tile.e[38] ),
    .Y(_01984_));
 sg13g2_nor2_1 _09517_ (.A(_01983_),
    .B(_01984_),
    .Y(_01985_));
 sg13g2_xnor2_1 _09518_ (.Y(_01986_),
    .A(_00772_),
    .B(_01985_));
 sg13g2_nand2_1 _09519_ (.Y(_01987_),
    .A(net443),
    .B(_01986_));
 sg13g2_xnor2_1 _09520_ (.Y(_01988_),
    .A(\clock_inst.hour_tile.e[39] ),
    .B(_01987_));
 sg13g2_nor2_1 _09521_ (.A(_01472_),
    .B(_01988_),
    .Y(_01989_));
 sg13g2_a21oi_1 _09522_ (.A1(_01212_),
    .A2(_01981_),
    .Y(_00184_),
    .B1(_01989_));
 sg13g2_buf_1 _09523_ (.A(net140),
    .X(_01990_));
 sg13g2_o21ai_1 _09524_ (.B1(net442),
    .Y(_01991_),
    .A1(_01701_),
    .A2(_01700_));
 sg13g2_a21oi_1 _09525_ (.A1(_01701_),
    .A2(_01700_),
    .Y(_01992_),
    .B1(_01991_));
 sg13g2_xnor2_1 _09526_ (.Y(_01993_),
    .A(\clock_inst.hour_tile.e[3] ),
    .B(_01992_));
 sg13g2_a21oi_1 _09527_ (.A1(net74),
    .A2(_01993_),
    .Y(_00185_),
    .B1(_01480_));
 sg13g2_buf_1 _09528_ (.A(\clock_inst.hour_tile.e[40] ),
    .X(_01994_));
 sg13g2_nand2_1 _09529_ (.Y(_01995_),
    .A(\clock_inst.hour_a[39] ),
    .B(\clock_inst.hour_tile.e[39] ));
 sg13g2_o21ai_1 _09530_ (.B1(_01995_),
    .Y(_01996_),
    .A1(_01983_),
    .A2(_01984_));
 sg13g2_or2_1 _09531_ (.X(_01997_),
    .B(\clock_inst.hour_tile.e[39] ),
    .A(\clock_inst.hour_a[39] ));
 sg13g2_nand2_1 _09532_ (.Y(_01998_),
    .A(_01996_),
    .B(_01997_));
 sg13g2_xnor2_1 _09533_ (.Y(_01999_),
    .A(_00779_),
    .B(_01998_));
 sg13g2_nor2_1 _09534_ (.A(net444),
    .B(_01999_),
    .Y(_02000_));
 sg13g2_xnor2_1 _09535_ (.Y(_02001_),
    .A(_01994_),
    .B(_02000_));
 sg13g2_a21oi_1 _09536_ (.A1(net74),
    .A2(_02001_),
    .Y(_00186_),
    .B1(_01489_));
 sg13g2_buf_1 _09537_ (.A(\clock_inst.hour_tile.e[41] ),
    .X(_02002_));
 sg13g2_buf_1 _09538_ (.A(net501),
    .X(_02003_));
 sg13g2_inv_1 _09539_ (.Y(_02004_),
    .A(_01994_));
 sg13g2_a21o_1 _09540_ (.A2(_01998_),
    .A1(_00779_),
    .B1(_02004_),
    .X(_02005_));
 sg13g2_o21ai_1 _09541_ (.B1(_02005_),
    .Y(_02006_),
    .A1(_00779_),
    .A2(_01998_));
 sg13g2_xnor2_1 _09542_ (.Y(_02007_),
    .A(_00782_),
    .B(_02006_));
 sg13g2_nor2_1 _09543_ (.A(net441),
    .B(_02007_),
    .Y(_02008_));
 sg13g2_xnor2_1 _09544_ (.Y(_02009_),
    .A(_02002_),
    .B(_02008_));
 sg13g2_a21oi_1 _09545_ (.A1(net74),
    .A2(_02009_),
    .Y(_00187_),
    .B1(_01507_));
 sg13g2_buf_1 _09546_ (.A(\clock_inst.hour_tile.e[42] ),
    .X(_02010_));
 sg13g2_nand2_1 _09547_ (.Y(_02011_),
    .A(_00782_),
    .B(_02002_));
 sg13g2_and3_1 _09548_ (.X(_02012_),
    .A(_02004_),
    .B(_01995_),
    .C(_02011_));
 sg13g2_o21ai_1 _09549_ (.B1(_02012_),
    .Y(_02013_),
    .A1(_01983_),
    .A2(_01984_));
 sg13g2_and3_1 _09550_ (.X(_02014_),
    .A(_00779_),
    .B(_01995_),
    .C(_02011_));
 sg13g2_o21ai_1 _09551_ (.B1(_02014_),
    .Y(_02015_),
    .A1(_01983_),
    .A2(_01984_));
 sg13g2_nor2_1 _09552_ (.A(\clock_inst.hour_a[40] ),
    .B(_01994_),
    .Y(_02016_));
 sg13g2_a221oi_1 _09553_ (.B2(_01994_),
    .C1(_01997_),
    .B1(\clock_inst.hour_a[40] ),
    .A1(_00782_),
    .Y(_02017_),
    .A2(_02002_));
 sg13g2_a21oi_1 _09554_ (.A1(_02011_),
    .A2(_02016_),
    .Y(_02018_),
    .B1(_02017_));
 sg13g2_nand3_1 _09555_ (.B(_02015_),
    .C(_02018_),
    .A(_02013_),
    .Y(_02019_));
 sg13g2_nor2_1 _09556_ (.A(_00782_),
    .B(_02002_),
    .Y(_02020_));
 sg13g2_or2_1 _09557_ (.X(_02021_),
    .B(_02020_),
    .A(_02019_));
 sg13g2_xnor2_1 _09558_ (.Y(_02022_),
    .A(_00788_),
    .B(_02021_));
 sg13g2_nor2_1 _09559_ (.A(net441),
    .B(_02022_),
    .Y(_02023_));
 sg13g2_xnor2_1 _09560_ (.Y(_02024_),
    .A(_02010_),
    .B(_02023_));
 sg13g2_a21oi_1 _09561_ (.A1(net74),
    .A2(_02024_),
    .Y(_00188_),
    .B1(_01517_));
 sg13g2_nor2_1 _09562_ (.A(\clock_inst.hour_a[42] ),
    .B(_02010_),
    .Y(_02025_));
 sg13g2_nand2_1 _09563_ (.Y(_02026_),
    .A(\clock_inst.hour_a[42] ),
    .B(_02010_));
 sg13g2_o21ai_1 _09564_ (.B1(_02026_),
    .Y(_02027_),
    .A1(_02021_),
    .A2(_02025_));
 sg13g2_xnor2_1 _09565_ (.Y(_02028_),
    .A(_00793_),
    .B(_02027_));
 sg13g2_nor2_1 _09566_ (.A(net441),
    .B(_02028_),
    .Y(_02029_));
 sg13g2_xnor2_1 _09567_ (.Y(_02030_),
    .A(\clock_inst.hour_tile.e[43] ),
    .B(_02029_));
 sg13g2_a21oi_1 _09568_ (.A1(net74),
    .A2(_02030_),
    .Y(_00189_),
    .B1(_01530_));
 sg13g2_buf_2 _09569_ (.A(\clock_inst.hour_tile.e[44] ),
    .X(_02031_));
 sg13g2_inv_1 _09570_ (.Y(_02032_),
    .A(_02010_));
 sg13g2_nor2_1 _09571_ (.A(_00793_),
    .B(\clock_inst.hour_tile.e[43] ),
    .Y(_02033_));
 sg13g2_nor3_1 _09572_ (.A(_02032_),
    .B(_02020_),
    .C(_02033_),
    .Y(_02034_));
 sg13g2_nand4_1 _09573_ (.B(_02015_),
    .C(_02018_),
    .A(_02013_),
    .Y(_02035_),
    .D(_02034_));
 sg13g2_nor3_1 _09574_ (.A(_00788_),
    .B(_02020_),
    .C(_02033_),
    .Y(_02036_));
 sg13g2_nand4_1 _09575_ (.B(_02015_),
    .C(_02018_),
    .A(_02013_),
    .Y(_02037_),
    .D(_02036_));
 sg13g2_nor2_1 _09576_ (.A(_02026_),
    .B(_02033_),
    .Y(_02038_));
 sg13g2_a21oi_1 _09577_ (.A1(_00793_),
    .A2(\clock_inst.hour_tile.e[43] ),
    .Y(_02039_),
    .B1(_02038_));
 sg13g2_nand3_1 _09578_ (.B(_02037_),
    .C(_02039_),
    .A(_02035_),
    .Y(_02040_));
 sg13g2_buf_1 _09579_ (.A(_02040_),
    .X(_02041_));
 sg13g2_buf_1 _09580_ (.A(_02041_),
    .X(_02042_));
 sg13g2_xnor2_1 _09581_ (.Y(_02043_),
    .A(net578),
    .B(net42));
 sg13g2_nor2_1 _09582_ (.A(_02003_),
    .B(_02043_),
    .Y(_02044_));
 sg13g2_xnor2_1 _09583_ (.Y(_02045_),
    .A(_02031_),
    .B(_02044_));
 sg13g2_a21oi_1 _09584_ (.A1(_01990_),
    .A2(_02045_),
    .Y(_00190_),
    .B1(_01554_));
 sg13g2_nor2_1 _09585_ (.A(_02031_),
    .B(_02041_),
    .Y(_02046_));
 sg13g2_nand2_1 _09586_ (.Y(_02047_),
    .A(net578),
    .B(_02046_));
 sg13g2_nand3b_1 _09587_ (.B(_02031_),
    .C(net42),
    .Y(_02048_),
    .A_N(net578));
 sg13g2_a21oi_1 _09588_ (.A1(_02047_),
    .A2(_02048_),
    .Y(_02049_),
    .B1(net447));
 sg13g2_xnor2_1 _09589_ (.Y(_02050_),
    .A(\clock_inst.hour_tile.e[45] ),
    .B(_02049_));
 sg13g2_xnor2_1 _09590_ (.Y(_02051_),
    .A(_01556_),
    .B(_01555_));
 sg13g2_nand2_1 _09591_ (.Y(_02052_),
    .A(_01573_),
    .B(_02051_));
 sg13g2_a21oi_1 _09592_ (.A1(\clock_inst.hour_c[45] ),
    .A2(_01925_),
    .Y(_02053_),
    .B1(_01926_));
 sg13g2_a22oi_1 _09593_ (.Y(_00191_),
    .B1(_02052_),
    .B2(_02053_),
    .A2(_02050_),
    .A1(net75));
 sg13g2_buf_1 _09594_ (.A(\clock_inst.hour_tile.e[46] ),
    .X(_02054_));
 sg13g2_inv_1 _09595_ (.Y(_02055_),
    .A(\clock_inst.hour_tile.e[45] ));
 sg13g2_inv_1 _09596_ (.Y(_02056_),
    .A(_02031_));
 sg13g2_nor3_1 _09597_ (.A(net578),
    .B(_02055_),
    .C(_02056_),
    .Y(_02057_));
 sg13g2_and2_1 _09598_ (.A(_02041_),
    .B(_02057_),
    .X(_02058_));
 sg13g2_nand2_1 _09599_ (.Y(_02059_),
    .A(net578),
    .B(_02055_));
 sg13g2_nor3_1 _09600_ (.A(_02031_),
    .B(net42),
    .C(_02059_),
    .Y(_02060_));
 sg13g2_buf_1 _09601_ (.A(_01796_),
    .X(_02061_));
 sg13g2_o21ai_1 _09602_ (.B1(_02061_),
    .Y(_02062_),
    .A1(_02058_),
    .A2(_02060_));
 sg13g2_xor2_1 _09603_ (.B(_02062_),
    .A(_02054_),
    .X(_02063_));
 sg13g2_xnor2_1 _09604_ (.Y(_02064_),
    .A(_01562_),
    .B(_01571_));
 sg13g2_nand2_1 _09605_ (.Y(_02065_),
    .A(net152),
    .B(_02064_));
 sg13g2_a21oi_1 _09606_ (.A1(\clock_inst.hour_c[46] ),
    .A2(net43),
    .Y(_02066_),
    .B1(net138));
 sg13g2_a22oi_1 _09607_ (.Y(_00192_),
    .B1(_02065_),
    .B2(_02066_),
    .A2(_02063_),
    .A1(net75));
 sg13g2_buf_1 _09608_ (.A(\clock_inst.hour_tile.e[47] ),
    .X(_02067_));
 sg13g2_nor2_1 _09609_ (.A(_02054_),
    .B(_02059_),
    .Y(_02068_));
 sg13g2_a22oi_1 _09610_ (.Y(_02069_),
    .B1(_02068_),
    .B2(_02046_),
    .A2(_02058_),
    .A1(_02054_));
 sg13g2_nor3_1 _09611_ (.A(_02067_),
    .B(_01682_),
    .C(_02069_),
    .Y(_02070_));
 sg13g2_nor2_1 _09612_ (.A(_01138_),
    .B(_02070_),
    .Y(_02071_));
 sg13g2_nor2_1 _09613_ (.A(_01057_),
    .B(net499),
    .Y(_02072_));
 sg13g2_buf_1 _09614_ (.A(_02072_),
    .X(_02073_));
 sg13g2_and2_1 _09615_ (.A(_02067_),
    .B(_02069_),
    .X(_02074_));
 sg13g2_nand2_1 _09616_ (.Y(_02075_),
    .A(_01577_),
    .B(_01240_));
 sg13g2_nand2_1 _09617_ (.Y(_02076_),
    .A(_01576_),
    .B(_01240_));
 sg13g2_mux2_1 _09618_ (.A0(_02075_),
    .A1(_02076_),
    .S(_01580_),
    .X(_02077_));
 sg13g2_a22oi_1 _09619_ (.Y(_02078_),
    .B1(_02074_),
    .B2(_02077_),
    .A2(net137),
    .A1(_02067_));
 sg13g2_o21ai_1 _09620_ (.B1(_02078_),
    .Y(_00193_),
    .A1(_01582_),
    .A2(_02071_));
 sg13g2_buf_2 _09621_ (.A(\clock_inst.hour_tile.e[48] ),
    .X(_02079_));
 sg13g2_nor3_1 _09622_ (.A(_02067_),
    .B(_02054_),
    .C(_02059_),
    .Y(_02080_));
 sg13g2_nand2_1 _09623_ (.Y(_02081_),
    .A(_02056_),
    .B(_02080_));
 sg13g2_or2_1 _09624_ (.X(_02082_),
    .B(_02081_),
    .A(net42));
 sg13g2_and2_1 _09625_ (.A(_02067_),
    .B(_02054_),
    .X(_02083_));
 sg13g2_nand3_1 _09626_ (.B(_02057_),
    .C(_02083_),
    .A(_02042_),
    .Y(_02084_));
 sg13g2_a21oi_1 _09627_ (.A1(_02082_),
    .A2(_02084_),
    .Y(_02085_),
    .B1(net501));
 sg13g2_xor2_1 _09628_ (.B(_02085_),
    .A(_02079_),
    .X(_02086_));
 sg13g2_nand2_1 _09629_ (.Y(_02087_),
    .A(net83),
    .B(_02086_));
 sg13g2_o21ai_1 _09630_ (.B1(_02087_),
    .Y(_00194_),
    .A1(net44),
    .A2(_01589_));
 sg13g2_buf_2 _09631_ (.A(\clock_inst.hour_tile.e[49] ),
    .X(_02088_));
 sg13g2_nand4_1 _09632_ (.B(_02031_),
    .C(_02079_),
    .A(\clock_inst.hour_tile.e[45] ),
    .Y(_02089_),
    .D(_02083_));
 sg13g2_nor2_1 _09633_ (.A(net578),
    .B(_02089_),
    .Y(_02090_));
 sg13g2_and2_1 _09634_ (.A(_02041_),
    .B(_02090_),
    .X(_02091_));
 sg13g2_nor2_1 _09635_ (.A(_02079_),
    .B(_02082_),
    .Y(_02092_));
 sg13g2_o21ai_1 _09636_ (.B1(_01797_),
    .Y(_02093_),
    .A1(_02091_),
    .A2(_02092_));
 sg13g2_xor2_1 _09637_ (.B(_02093_),
    .A(_02088_),
    .X(_02094_));
 sg13g2_a22oi_1 _09638_ (.Y(_00195_),
    .B1(_02094_),
    .B2(_01787_),
    .A2(_01601_),
    .A1(_01600_));
 sg13g2_a21oi_1 _09639_ (.A1(_01701_),
    .A2(_01700_),
    .Y(_02095_),
    .B1(_01704_));
 sg13g2_xnor2_1 _09640_ (.Y(_02096_),
    .A(_00964_),
    .B(_02095_));
 sg13g2_nor2_1 _09641_ (.A(_02003_),
    .B(_02096_),
    .Y(_02097_));
 sg13g2_xnor2_1 _09642_ (.Y(_02098_),
    .A(\clock_inst.hour_tile.e[4] ),
    .B(_02097_));
 sg13g2_a21oi_1 _09643_ (.A1(_01990_),
    .A2(_02098_),
    .Y(_00196_),
    .B1(_01607_));
 sg13g2_buf_1 _09644_ (.A(\clock_inst.hour_tile.e[50] ),
    .X(_02099_));
 sg13g2_inv_1 _09645_ (.Y(_02100_),
    .A(_02099_));
 sg13g2_buf_1 _09646_ (.A(net242),
    .X(_02101_));
 sg13g2_inv_1 _09647_ (.Y(_02102_),
    .A(_02080_));
 sg13g2_nor3_1 _09648_ (.A(_02079_),
    .B(_02088_),
    .C(_02102_),
    .Y(_02103_));
 sg13g2_a22oi_1 _09649_ (.Y(_02104_),
    .B1(_02103_),
    .B2(_02046_),
    .A2(_02091_),
    .A1(_02088_));
 sg13g2_nand2_1 _09650_ (.Y(_02105_),
    .A(_02100_),
    .B(_02104_));
 sg13g2_nand3b_1 _09651_ (.B(net356),
    .C(_02099_),
    .Y(_02106_),
    .A_N(_02104_));
 sg13g2_nand3_1 _09652_ (.B(_02105_),
    .C(_02106_),
    .A(_02101_),
    .Y(_02107_));
 sg13g2_a22oi_1 _09653_ (.Y(_00197_),
    .B1(_02107_),
    .B2(_01620_),
    .A2(net137),
    .A1(_02100_));
 sg13g2_a21oi_1 _09654_ (.A1(net578),
    .A2(_02031_),
    .Y(_02108_),
    .B1(_02099_));
 sg13g2_nand3b_1 _09655_ (.B(_02103_),
    .C(_02108_),
    .Y(_02109_),
    .A_N(net42));
 sg13g2_nand4_1 _09656_ (.B(_02099_),
    .C(net42),
    .A(_02088_),
    .Y(_02110_),
    .D(_02090_));
 sg13g2_a21oi_1 _09657_ (.A1(_02109_),
    .A2(_02110_),
    .Y(_02111_),
    .B1(_01681_));
 sg13g2_xor2_1 _09658_ (.B(_02111_),
    .A(\clock_inst.hour_tile.e[51] ),
    .X(_02112_));
 sg13g2_a22oi_1 _09659_ (.Y(_02113_),
    .B1(_02112_),
    .B2(_01590_),
    .A2(net82),
    .A1(\clock_inst.hour_c[51] ));
 sg13g2_o21ai_1 _09660_ (.B1(_02113_),
    .Y(_00198_),
    .A1(net44),
    .A2(_01623_));
 sg13g2_nand3_1 _09661_ (.B(_02099_),
    .C(\clock_inst.hour_tile.e[51] ),
    .A(_02088_),
    .Y(_02114_));
 sg13g2_o21ai_1 _09662_ (.B1(_02042_),
    .Y(_02115_),
    .A1(_02089_),
    .A2(_02114_));
 sg13g2_nor4_1 _09663_ (.A(_02088_),
    .B(_02099_),
    .C(\clock_inst.hour_tile.e[51] ),
    .D(_02081_),
    .Y(_02116_));
 sg13g2_or2_1 _09664_ (.X(_02117_),
    .B(_02116_),
    .A(net42));
 sg13g2_a21oi_1 _09665_ (.A1(net578),
    .A2(_02079_),
    .Y(_02118_),
    .B1(_01676_));
 sg13g2_nand3_1 _09666_ (.B(_02117_),
    .C(_02118_),
    .A(_02115_),
    .Y(_02119_));
 sg13g2_xnor2_1 _09667_ (.Y(_02120_),
    .A(\clock_inst.hour_tile.e[52] ),
    .B(_02119_));
 sg13g2_a22oi_1 _09668_ (.Y(_02121_),
    .B1(_02120_),
    .B2(_01590_),
    .A2(_01611_),
    .A1(\clock_inst.hour_c[52] ));
 sg13g2_o21ai_1 _09669_ (.B1(_02121_),
    .Y(_00199_),
    .A1(_01583_),
    .A2(_01629_));
 sg13g2_xnor2_1 _09670_ (.Y(_02122_),
    .A(\clock_inst.hour_tile.e0[53] ),
    .B(_01636_));
 sg13g2_nor2_1 _09671_ (.A(_02079_),
    .B(\clock_inst.hour_tile.e[52] ),
    .Y(_02123_));
 sg13g2_nand3_1 _09672_ (.B(_02116_),
    .C(_02123_),
    .A(net500),
    .Y(_02124_));
 sg13g2_inv_1 _09673_ (.Y(_02125_),
    .A(_02114_));
 sg13g2_nand4_1 _09674_ (.B(net500),
    .C(_02090_),
    .A(\clock_inst.hour_tile.e[52] ),
    .Y(_02126_),
    .D(_02125_));
 sg13g2_mux2_1 _09675_ (.A0(_02124_),
    .A1(_02126_),
    .S(net42),
    .X(_02127_));
 sg13g2_xnor2_1 _09676_ (.Y(_02128_),
    .A(\clock_inst.hour_tile.e[53] ),
    .B(_02127_));
 sg13g2_nor3_1 _09677_ (.A(_01701_),
    .B(_01559_),
    .C(net87),
    .Y(_02129_));
 sg13g2_a21oi_1 _09678_ (.A1(net145),
    .A2(_02128_),
    .Y(_02130_),
    .B1(_02129_));
 sg13g2_o21ai_1 _09679_ (.B1(_02130_),
    .Y(_00200_),
    .A1(_01583_),
    .A2(_02122_));
 sg13g2_buf_1 _09680_ (.A(net236),
    .X(_02131_));
 sg13g2_or3_1 _09681_ (.A(_00806_),
    .B(_01706_),
    .C(_01707_),
    .X(_02132_));
 sg13g2_o21ai_1 _09682_ (.B1(_00806_),
    .Y(_02133_),
    .A1(_01706_),
    .A2(_01707_));
 sg13g2_nand3_1 _09683_ (.B(_02132_),
    .C(_02133_),
    .A(net443),
    .Y(_02134_));
 sg13g2_xor2_1 _09684_ (.B(_02134_),
    .A(_01711_),
    .X(_02135_));
 sg13g2_o21ai_1 _09685_ (.B1(_01647_),
    .Y(_00201_),
    .A1(net135),
    .A2(_02135_));
 sg13g2_nor2_1 _09686_ (.A(_01712_),
    .B(_01762_),
    .Y(_02136_));
 sg13g2_xnor2_1 _09687_ (.Y(_02137_),
    .A(_00813_),
    .B(_02136_));
 sg13g2_nor2_1 _09688_ (.A(net447),
    .B(_02137_),
    .Y(_02138_));
 sg13g2_xnor2_1 _09689_ (.Y(_02139_),
    .A(_01708_),
    .B(_02138_));
 sg13g2_o21ai_1 _09690_ (.B1(_01653_),
    .Y(_00202_),
    .A1(net135),
    .A2(_02139_));
 sg13g2_nor3_1 _09691_ (.A(_01709_),
    .B(_01712_),
    .C(_01762_),
    .Y(_02140_));
 sg13g2_o21ai_1 _09692_ (.B1(_01709_),
    .Y(_02141_),
    .A1(_01712_),
    .A2(_01762_));
 sg13g2_o21ai_1 _09693_ (.B1(_02141_),
    .Y(_02142_),
    .A1(_00813_),
    .A2(_02140_));
 sg13g2_xnor2_1 _09694_ (.Y(_02143_),
    .A(_00819_),
    .B(_02142_));
 sg13g2_nor3_1 _09695_ (.A(_01689_),
    .B(_01248_),
    .C(_02143_),
    .Y(_02144_));
 sg13g2_and4_1 _09696_ (.A(_01689_),
    .B(net143),
    .C(_01965_),
    .D(_02143_),
    .X(_02145_));
 sg13g2_nor3_1 _09697_ (.A(_01689_),
    .B(net156),
    .C(_01965_),
    .Y(_02146_));
 sg13g2_nor4_1 _09698_ (.A(_01662_),
    .B(_02144_),
    .C(_02145_),
    .D(_02146_),
    .Y(_00203_));
 sg13g2_xnor2_1 _09699_ (.Y(_02147_),
    .A(_01760_),
    .B(_01724_));
 sg13g2_nor2_1 _09700_ (.A(net441),
    .B(_02147_),
    .Y(_02148_));
 sg13g2_xnor2_1 _09701_ (.Y(_02149_),
    .A(_01729_),
    .B(_02148_));
 sg13g2_a21oi_1 _09702_ (.A1(net74),
    .A2(_02149_),
    .Y(_00204_),
    .B1(_01667_));
 sg13g2_mux2_1 _09703_ (.A0(_01731_),
    .A1(_01734_),
    .S(_01724_),
    .X(_02150_));
 sg13g2_xnor2_1 _09704_ (.Y(_02151_),
    .A(_01725_),
    .B(_02150_));
 sg13g2_nand2_1 _09705_ (.Y(_02152_),
    .A(net136),
    .B(_02151_));
 sg13g2_and2_1 _09706_ (.A(_01673_),
    .B(_02152_),
    .X(_00205_));
 sg13g2_buf_1 _09707_ (.A(\clock_inst.minute[4] ),
    .X(_02153_));
 sg13g2_buf_1 _09708_ (.A(\clock_inst.minute[0] ),
    .X(_02154_));
 sg13g2_inv_1 _09709_ (.Y(_02155_),
    .A(_02154_));
 sg13g2_buf_1 _09710_ (.A(\clock_inst.minute[1] ),
    .X(_02156_));
 sg13g2_inv_1 _09711_ (.Y(_02157_),
    .A(_02156_));
 sg13g2_nor2_1 _09712_ (.A(_02155_),
    .B(_02157_),
    .Y(_02158_));
 sg13g2_buf_2 _09713_ (.A(_02158_),
    .X(_02159_));
 sg13g2_nor2_1 _09714_ (.A(net571),
    .B(_02159_),
    .Y(_02160_));
 sg13g2_buf_1 _09715_ (.A(\clock_inst.minute[5] ),
    .X(_02161_));
 sg13g2_buf_2 _09716_ (.A(\clock_inst.minute[3] ),
    .X(_02162_));
 sg13g2_inv_1 _09717_ (.Y(_02163_),
    .A(_02162_));
 sg13g2_buf_1 _09718_ (.A(\clock_inst.minute[2] ),
    .X(_02164_));
 sg13g2_inv_1 _09719_ (.Y(_02165_),
    .A(_02164_));
 sg13g2_nor2_1 _09720_ (.A(_02163_),
    .B(_02165_),
    .Y(_02166_));
 sg13g2_buf_1 _09721_ (.A(_02166_),
    .X(_02167_));
 sg13g2_nand2_1 _09722_ (.Y(_02168_),
    .A(_02161_),
    .B(_02167_));
 sg13g2_o21ai_1 _09723_ (.B1(net583),
    .Y(_02169_),
    .A1(_02160_),
    .A2(_02168_));
 sg13g2_buf_1 _09724_ (.A(_02169_),
    .X(_02170_));
 sg13g2_buf_1 _09725_ (.A(_02170_),
    .X(_02171_));
 sg13g2_buf_1 _09726_ (.A(net73),
    .X(_02172_));
 sg13g2_buf_1 _09727_ (.A(_02156_),
    .X(_02173_));
 sg13g2_nor2_1 _09728_ (.A(_02154_),
    .B(net541),
    .Y(_02174_));
 sg13g2_buf_2 _09729_ (.A(_02174_),
    .X(_02175_));
 sg13g2_buf_1 _09730_ (.A(_02164_),
    .X(_02176_));
 sg13g2_buf_1 _09731_ (.A(net540),
    .X(_02177_));
 sg13g2_inv_2 _09732_ (.Y(_02178_),
    .A(net570));
 sg13g2_nand2_1 _09733_ (.Y(_02179_),
    .A(net571),
    .B(_02178_));
 sg13g2_buf_2 _09734_ (.A(_02179_),
    .X(_02180_));
 sg13g2_nor2_2 _09735_ (.A(net498),
    .B(_02180_),
    .Y(_02181_));
 sg13g2_buf_1 _09736_ (.A(_02162_),
    .X(_02182_));
 sg13g2_buf_1 _09737_ (.A(net539),
    .X(_02183_));
 sg13g2_buf_1 _09738_ (.A(net497),
    .X(_02184_));
 sg13g2_buf_1 _09739_ (.A(net440),
    .X(_02185_));
 sg13g2_buf_1 _09740_ (.A(net541),
    .X(_02186_));
 sg13g2_buf_1 _09741_ (.A(net496),
    .X(_02187_));
 sg13g2_buf_1 _09742_ (.A(net439),
    .X(_02188_));
 sg13g2_buf_1 _09743_ (.A(_02165_),
    .X(_02189_));
 sg13g2_nor2_1 _09744_ (.A(net495),
    .B(_02178_),
    .Y(_02190_));
 sg13g2_buf_1 _09745_ (.A(_02190_),
    .X(_02191_));
 sg13g2_buf_1 _09746_ (.A(_02155_),
    .X(_02192_));
 sg13g2_inv_1 _09747_ (.Y(_02193_),
    .A(net571));
 sg13g2_buf_1 _09748_ (.A(_02193_),
    .X(_02194_));
 sg13g2_buf_1 _09749_ (.A(net493),
    .X(_02195_));
 sg13g2_nor2_1 _09750_ (.A(net494),
    .B(net438),
    .Y(_02196_));
 sg13g2_buf_1 _09751_ (.A(net541),
    .X(_02197_));
 sg13g2_buf_1 _09752_ (.A(net492),
    .X(_02198_));
 sg13g2_nor2_1 _09753_ (.A(_02164_),
    .B(net570),
    .Y(_02199_));
 sg13g2_buf_1 _09754_ (.A(_02199_),
    .X(_02200_));
 sg13g2_buf_1 _09755_ (.A(_02200_),
    .X(_02201_));
 sg13g2_nand2_1 _09756_ (.Y(_02202_),
    .A(_02198_),
    .B(net436));
 sg13g2_buf_1 _09757_ (.A(_02157_),
    .X(_02203_));
 sg13g2_nand2_2 _09758_ (.Y(_02204_),
    .A(_02203_),
    .B(net570));
 sg13g2_nand2_1 _09759_ (.Y(_02205_),
    .A(_02202_),
    .B(_02204_));
 sg13g2_buf_2 _09760_ (.A(net498),
    .X(_02206_));
 sg13g2_nor2_1 _09761_ (.A(net571),
    .B(\clock_inst.minute[5] ),
    .Y(_02207_));
 sg13g2_buf_2 _09762_ (.A(_02207_),
    .X(_02208_));
 sg13g2_buf_1 _09763_ (.A(net492),
    .X(_02209_));
 sg13g2_o21ai_1 _09764_ (.B1(net434),
    .Y(_02210_),
    .A1(net435),
    .A2(_02208_));
 sg13g2_buf_2 _09765_ (.A(net498),
    .X(_02211_));
 sg13g2_buf_1 _09766_ (.A(net571),
    .X(_02212_));
 sg13g2_nor2_2 _09767_ (.A(net492),
    .B(net538),
    .Y(_02213_));
 sg13g2_buf_1 _09768_ (.A(net570),
    .X(_02214_));
 sg13g2_buf_1 _09769_ (.A(net537),
    .X(_02215_));
 sg13g2_o21ai_1 _09770_ (.B1(net490),
    .Y(_02216_),
    .A1(net433),
    .A2(_02213_));
 sg13g2_buf_1 _09771_ (.A(_02154_),
    .X(_02217_));
 sg13g2_buf_1 _09772_ (.A(net536),
    .X(_02218_));
 sg13g2_buf_1 _09773_ (.A(net489),
    .X(_02219_));
 sg13g2_a21oi_1 _09774_ (.A1(_02210_),
    .A2(_02216_),
    .Y(_02220_),
    .B1(net432));
 sg13g2_a221oi_1 _09775_ (.B2(_02205_),
    .C1(_02220_),
    .B1(_02196_),
    .A1(net353),
    .Y(_02221_),
    .A2(net352));
 sg13g2_buf_1 _09776_ (.A(net538),
    .X(_02222_));
 sg13g2_buf_1 _09777_ (.A(net488),
    .X(_02223_));
 sg13g2_buf_1 _09778_ (.A(net495),
    .X(_02224_));
 sg13g2_buf_1 _09779_ (.A(net430),
    .X(_02225_));
 sg13g2_buf_1 _09780_ (.A(_02178_),
    .X(_02226_));
 sg13g2_nor2_1 _09781_ (.A(net491),
    .B(net487),
    .Y(_02227_));
 sg13g2_buf_2 _09782_ (.A(_02227_),
    .X(_02228_));
 sg13g2_nor2_2 _09783_ (.A(net540),
    .B(net487),
    .Y(_02229_));
 sg13g2_nand2_2 _09784_ (.Y(_02230_),
    .A(net496),
    .B(_02229_));
 sg13g2_o21ai_1 _09785_ (.B1(_02230_),
    .Y(_02231_),
    .A1(net351),
    .A2(_02228_));
 sg13g2_buf_1 _09786_ (.A(net437),
    .X(_02232_));
 sg13g2_nand2_2 _09787_ (.Y(_02233_),
    .A(net495),
    .B(net487));
 sg13g2_buf_1 _09788_ (.A(_02233_),
    .X(_02234_));
 sg13g2_buf_1 _09789_ (.A(net438),
    .X(_02235_));
 sg13g2_buf_1 _09790_ (.A(net348),
    .X(_02236_));
 sg13g2_o21ai_1 _09791_ (.B1(net231),
    .Y(_02237_),
    .A1(net350),
    .A2(net349));
 sg13g2_buf_1 _09792_ (.A(net494),
    .X(_02238_));
 sg13g2_buf_1 _09793_ (.A(_02238_),
    .X(_02239_));
 sg13g2_buf_1 _09794_ (.A(net539),
    .X(_02240_));
 sg13g2_buf_1 _09795_ (.A(net486),
    .X(_02241_));
 sg13g2_buf_1 _09796_ (.A(net428),
    .X(_02242_));
 sg13g2_a221oi_1 _09797_ (.B2(net347),
    .C1(net346),
    .B1(_02237_),
    .A1(_02223_),
    .Y(_02243_),
    .A2(_02231_));
 sg13g2_a21oi_1 _09798_ (.A1(net354),
    .A2(_02221_),
    .Y(_02244_),
    .B1(_02243_));
 sg13g2_a21oi_1 _09799_ (.A1(_02175_),
    .A2(_02181_),
    .Y(_02245_),
    .B1(_02244_));
 sg13g2_buf_1 _09800_ (.A(_02170_),
    .X(_02246_));
 sg13g2_buf_1 _09801_ (.A(net72),
    .X(_02247_));
 sg13g2_nand2_1 _09802_ (.Y(_02248_),
    .A(\clock_inst.min_a[0] ),
    .B(net40));
 sg13g2_o21ai_1 _09803_ (.B1(_02248_),
    .Y(_00206_),
    .A1(net41),
    .A2(_02245_));
 sg13g2_buf_1 _09804_ (.A(\clock_inst.min_a[10] ),
    .X(_02249_));
 sg13g2_inv_1 _09805_ (.Y(_02250_),
    .A(net569));
 sg13g2_buf_1 _09806_ (.A(net73),
    .X(_02251_));
 sg13g2_nor2_1 _09807_ (.A(_02160_),
    .B(_02168_),
    .Y(_02252_));
 sg13g2_nand2_1 _09808_ (.Y(_02253_),
    .A(_02165_),
    .B(_02208_));
 sg13g2_nand2_1 _09809_ (.Y(_02254_),
    .A(_02157_),
    .B(_02163_));
 sg13g2_buf_2 _09810_ (.A(_02254_),
    .X(_02255_));
 sg13g2_nor3_1 _09811_ (.A(_02154_),
    .B(_02253_),
    .C(_02255_),
    .Y(_02256_));
 sg13g2_or3_1 _09812_ (.A(net513),
    .B(_02252_),
    .C(_02256_),
    .X(_02257_));
 sg13g2_buf_1 _09813_ (.A(_02257_),
    .X(_02258_));
 sg13g2_nand2_1 _09814_ (.Y(_02259_),
    .A(net493),
    .B(_02178_));
 sg13g2_buf_2 _09815_ (.A(_02259_),
    .X(_02260_));
 sg13g2_nand2_1 _09816_ (.Y(_02261_),
    .A(_02159_),
    .B(_02167_));
 sg13g2_nor2_1 _09817_ (.A(_02260_),
    .B(_02261_),
    .Y(_02262_));
 sg13g2_nor2_1 _09818_ (.A(_02258_),
    .B(_02262_),
    .Y(_02263_));
 sg13g2_buf_1 _09819_ (.A(_02180_),
    .X(_02264_));
 sg13g2_buf_1 _09820_ (.A(net488),
    .X(_02265_));
 sg13g2_buf_1 _09821_ (.A(net427),
    .X(_02266_));
 sg13g2_buf_1 _09822_ (.A(_02159_),
    .X(_02267_));
 sg13g2_buf_1 _09823_ (.A(_02267_),
    .X(_02268_));
 sg13g2_buf_1 _09824_ (.A(_02167_),
    .X(_02269_));
 sg13g2_buf_1 _09825_ (.A(net342),
    .X(_02270_));
 sg13g2_o21ai_1 _09826_ (.B1(net229),
    .Y(_02271_),
    .A1(net344),
    .A2(net230));
 sg13g2_buf_1 _09827_ (.A(net231),
    .X(_02272_));
 sg13g2_buf_1 _09828_ (.A(net487),
    .X(_02273_));
 sg13g2_buf_1 _09829_ (.A(net426),
    .X(_02274_));
 sg13g2_nor2_1 _09830_ (.A(_02274_),
    .B(net342),
    .Y(_02275_));
 sg13g2_nand2_1 _09831_ (.Y(_02276_),
    .A(net134),
    .B(_02275_));
 sg13g2_buf_1 _09832_ (.A(net437),
    .X(_02277_));
 sg13g2_buf_1 _09833_ (.A(net340),
    .X(_02278_));
 sg13g2_nor2_1 _09834_ (.A(net540),
    .B(_02153_),
    .Y(_02279_));
 sg13g2_buf_1 _09835_ (.A(_02279_),
    .X(_02280_));
 sg13g2_buf_1 _09836_ (.A(_02280_),
    .X(_02281_));
 sg13g2_buf_1 _09837_ (.A(_02162_),
    .X(_02282_));
 sg13g2_nor2_1 _09838_ (.A(_02154_),
    .B(net534),
    .Y(_02283_));
 sg13g2_buf_2 _09839_ (.A(_02283_),
    .X(_02284_));
 sg13g2_nand2_1 _09840_ (.Y(_02285_),
    .A(_02162_),
    .B(_02164_));
 sg13g2_buf_1 _09841_ (.A(_02285_),
    .X(_02286_));
 sg13g2_nor2_2 _09842_ (.A(net426),
    .B(net485),
    .Y(_02287_));
 sg13g2_a21oi_1 _09843_ (.A1(net339),
    .A2(_02284_),
    .Y(_02288_),
    .B1(_02287_));
 sg13g2_or2_1 _09844_ (.X(_02289_),
    .B(_02288_),
    .A(_02278_));
 sg13g2_nand4_1 _09845_ (.B(_02271_),
    .C(_02276_),
    .A(_02264_),
    .Y(_02290_),
    .D(_02289_));
 sg13g2_a22oi_1 _09846_ (.Y(_00207_),
    .B1(_02263_),
    .B2(_02290_),
    .A2(net39),
    .A1(_02250_));
 sg13g2_nor2_1 _09847_ (.A(net433),
    .B(_02260_),
    .Y(_02291_));
 sg13g2_buf_1 _09848_ (.A(_02163_),
    .X(_02292_));
 sg13g2_nor2_1 _09849_ (.A(net541),
    .B(net484),
    .Y(_02293_));
 sg13g2_buf_2 _09850_ (.A(_02293_),
    .X(_02294_));
 sg13g2_buf_1 _09851_ (.A(_02294_),
    .X(_02295_));
 sg13g2_nand2_1 _09852_ (.Y(_02296_),
    .A(_02153_),
    .B(net570));
 sg13g2_buf_2 _09853_ (.A(_02296_),
    .X(_02297_));
 sg13g2_nand2_1 _09854_ (.Y(_02298_),
    .A(net540),
    .B(_02297_));
 sg13g2_inv_1 _09855_ (.Y(_02299_),
    .A(_02298_));
 sg13g2_nor2_1 _09856_ (.A(net491),
    .B(net534),
    .Y(_02300_));
 sg13g2_buf_2 _09857_ (.A(_02300_),
    .X(_02301_));
 sg13g2_buf_1 _09858_ (.A(net536),
    .X(_02302_));
 sg13g2_buf_1 _09859_ (.A(net483),
    .X(_02303_));
 sg13g2_buf_1 _09860_ (.A(net425),
    .X(_02304_));
 sg13g2_nand2_1 _09861_ (.Y(_02305_),
    .A(_02156_),
    .B(_02178_));
 sg13g2_buf_2 _09862_ (.A(_02305_),
    .X(_02306_));
 sg13g2_nand2_1 _09863_ (.Y(_02307_),
    .A(_02204_),
    .B(_02306_));
 sg13g2_buf_2 _09864_ (.A(_02307_),
    .X(_02308_));
 sg13g2_nand2_1 _09865_ (.Y(_02309_),
    .A(_02163_),
    .B(_02193_));
 sg13g2_buf_2 _09866_ (.A(_02309_),
    .X(_02310_));
 sg13g2_nor2_1 _09867_ (.A(net540),
    .B(net493),
    .Y(_02311_));
 sg13g2_nand2_2 _09868_ (.Y(_02312_),
    .A(_02182_),
    .B(_02311_));
 sg13g2_nand2_1 _09869_ (.Y(_02313_),
    .A(_02310_),
    .B(_02312_));
 sg13g2_nor2_1 _09870_ (.A(_02162_),
    .B(net493),
    .Y(_02314_));
 sg13g2_buf_1 _09871_ (.A(_02314_),
    .X(_02315_));
 sg13g2_nand2_1 _09872_ (.Y(_02316_),
    .A(net491),
    .B(net540));
 sg13g2_buf_2 _09873_ (.A(_02316_),
    .X(_02317_));
 sg13g2_nand2_1 _09874_ (.Y(_02318_),
    .A(_02230_),
    .B(_02317_));
 sg13g2_a22oi_1 _09875_ (.Y(_02319_),
    .B1(_02315_),
    .B2(_02318_),
    .A2(_02313_),
    .A1(_02308_));
 sg13g2_buf_1 _09876_ (.A(net536),
    .X(_02320_));
 sg13g2_buf_1 _09877_ (.A(net482),
    .X(_02321_));
 sg13g2_buf_1 _09878_ (.A(net424),
    .X(_02322_));
 sg13g2_buf_1 _09879_ (.A(net484),
    .X(_02323_));
 sg13g2_nor2_1 _09880_ (.A(net423),
    .B(_02177_),
    .Y(_02324_));
 sg13g2_nor2_1 _09881_ (.A(net571),
    .B(_02178_),
    .Y(_02325_));
 sg13g2_buf_2 _09882_ (.A(_02325_),
    .X(_02326_));
 sg13g2_nor2_1 _09883_ (.A(net539),
    .B(_02180_),
    .Y(_02327_));
 sg13g2_a21oi_1 _09884_ (.A1(_02324_),
    .A2(_02326_),
    .Y(_02328_),
    .B1(_02327_));
 sg13g2_buf_1 _09885_ (.A(_02214_),
    .X(_02329_));
 sg13g2_nor2_2 _09886_ (.A(net495),
    .B(net493),
    .Y(_02330_));
 sg13g2_nor2_1 _09887_ (.A(net537),
    .B(_02330_),
    .Y(_02331_));
 sg13g2_a221oi_1 _09888_ (.B2(net486),
    .C1(net434),
    .B1(_02331_),
    .A1(net481),
    .Y(_02332_),
    .A2(net337));
 sg13g2_a21oi_1 _09889_ (.A1(net340),
    .A2(_02328_),
    .Y(_02333_),
    .B1(_02332_));
 sg13g2_buf_1 _09890_ (.A(net492),
    .X(_02334_));
 sg13g2_nor2_1 _09891_ (.A(_02194_),
    .B(net570),
    .Y(_02335_));
 sg13g2_buf_2 _09892_ (.A(_02335_),
    .X(_02336_));
 sg13g2_nand2_1 _09893_ (.Y(_02337_),
    .A(net422),
    .B(_02336_));
 sg13g2_nand2_1 _09894_ (.Y(_02338_),
    .A(net484),
    .B(_02161_));
 sg13g2_buf_1 _09895_ (.A(_02338_),
    .X(_02339_));
 sg13g2_buf_1 _09896_ (.A(net351),
    .X(_02340_));
 sg13g2_a21oi_1 _09897_ (.A1(_02337_),
    .A2(net335),
    .Y(_02341_),
    .B1(net226));
 sg13g2_nor3_1 _09898_ (.A(net336),
    .B(_02333_),
    .C(_02341_),
    .Y(_02342_));
 sg13g2_a21oi_1 _09899_ (.A1(_02304_),
    .A2(_02319_),
    .Y(_02343_),
    .B1(_02342_));
 sg13g2_a221oi_1 _09900_ (.B2(_02301_),
    .C1(_02343_),
    .B1(_02299_),
    .A1(_02291_),
    .Y(_02344_),
    .A2(net227));
 sg13g2_buf_8 _09901_ (.A(\clock_inst.min_a[18] ),
    .X(_02345_));
 sg13g2_nand2_1 _09902_ (.Y(_02346_),
    .A(_02345_),
    .B(_02247_));
 sg13g2_o21ai_1 _09903_ (.B1(_02346_),
    .Y(_00208_),
    .A1(_02172_),
    .A2(_02344_));
 sg13g2_buf_1 _09904_ (.A(\clock_inst.min_a[19] ),
    .X(_02347_));
 sg13g2_inv_1 _09905_ (.Y(_02348_),
    .A(_02347_));
 sg13g2_nor2_1 _09906_ (.A(net513),
    .B(_02252_),
    .Y(_02349_));
 sg13g2_buf_1 _09907_ (.A(_02349_),
    .X(_02350_));
 sg13g2_buf_1 _09908_ (.A(_02350_),
    .X(_02351_));
 sg13g2_nand2_1 _09909_ (.Y(_02352_),
    .A(net495),
    .B(net570));
 sg13g2_buf_2 _09910_ (.A(_02352_),
    .X(_02353_));
 sg13g2_nor2_2 _09911_ (.A(net539),
    .B(_02353_),
    .Y(_02354_));
 sg13g2_buf_1 _09912_ (.A(_02282_),
    .X(_02355_));
 sg13g2_buf_1 _09913_ (.A(net480),
    .X(_02356_));
 sg13g2_a21oi_1 _09914_ (.A1(net421),
    .A2(net349),
    .Y(_02357_),
    .B1(_02277_));
 sg13g2_o21ai_1 _09915_ (.B1(net344),
    .Y(_02358_),
    .A1(_02354_),
    .A2(_02357_));
 sg13g2_buf_1 _09916_ (.A(net439),
    .X(_02359_));
 sg13g2_nand2_1 _09917_ (.Y(_02360_),
    .A(_02176_),
    .B(_02178_));
 sg13g2_buf_2 _09918_ (.A(_02360_),
    .X(_02361_));
 sg13g2_nand2_1 _09919_ (.Y(_02362_),
    .A(net488),
    .B(_02361_));
 sg13g2_nor2_1 _09920_ (.A(net495),
    .B(net538),
    .Y(_02363_));
 sg13g2_buf_1 _09921_ (.A(_02363_),
    .X(_02364_));
 sg13g2_buf_1 _09922_ (.A(net333),
    .X(_02365_));
 sg13g2_a21o_1 _09923_ (.A2(_02362_),
    .A1(_02183_),
    .B1(net225),
    .X(_02366_));
 sg13g2_nand2_1 _09924_ (.Y(_02367_),
    .A(_02194_),
    .B(net570));
 sg13g2_buf_1 _09925_ (.A(_02367_),
    .X(_02368_));
 sg13g2_nor2_2 _09926_ (.A(net423),
    .B(_02368_),
    .Y(_02369_));
 sg13g2_a21oi_1 _09927_ (.A1(_02359_),
    .A2(_02366_),
    .Y(_02370_),
    .B1(_02369_));
 sg13g2_buf_1 _09928_ (.A(net336),
    .X(_02371_));
 sg13g2_a21oi_1 _09929_ (.A1(_02358_),
    .A2(_02370_),
    .Y(_02372_),
    .B1(net224));
 sg13g2_buf_1 _09930_ (.A(_02359_),
    .X(_02373_));
 sg13g2_buf_1 _09931_ (.A(_02324_),
    .X(_02374_));
 sg13g2_buf_1 _09932_ (.A(_02326_),
    .X(_02375_));
 sg13g2_buf_1 _09933_ (.A(net332),
    .X(_02376_));
 sg13g2_nor2_1 _09934_ (.A(_02189_),
    .B(net537),
    .Y(_02377_));
 sg13g2_buf_2 _09935_ (.A(_02377_),
    .X(_02378_));
 sg13g2_buf_1 _09936_ (.A(_02378_),
    .X(_02379_));
 sg13g2_nor2_2 _09937_ (.A(net494),
    .B(_02355_),
    .Y(_02380_));
 sg13g2_a22oi_1 _09938_ (.Y(_02381_),
    .B1(net220),
    .B2(_02380_),
    .A2(net221),
    .A1(net222));
 sg13g2_buf_1 _09939_ (.A(net340),
    .X(_02382_));
 sg13g2_nor2_1 _09940_ (.A(net534),
    .B(net540),
    .Y(_02383_));
 sg13g2_buf_1 _09941_ (.A(_02383_),
    .X(_02384_));
 sg13g2_nand2_2 _09942_ (.Y(_02385_),
    .A(_02326_),
    .B(net420));
 sg13g2_nor2_1 _09943_ (.A(_02193_),
    .B(_02178_),
    .Y(_02386_));
 sg13g2_buf_1 _09944_ (.A(_02386_),
    .X(_02387_));
 sg13g2_nand2_1 _09945_ (.Y(_02388_),
    .A(net495),
    .B(_02387_));
 sg13g2_nand2_1 _09946_ (.Y(_02389_),
    .A(_02260_),
    .B(_02388_));
 sg13g2_nand2_1 _09947_ (.Y(_02390_),
    .A(net497),
    .B(_02389_));
 sg13g2_buf_1 _09948_ (.A(net429),
    .X(_02391_));
 sg13g2_a21oi_1 _09949_ (.A1(_02385_),
    .A2(_02390_),
    .Y(_02392_),
    .B1(net331));
 sg13g2_nor3_1 _09950_ (.A(net219),
    .B(_02327_),
    .C(_02392_),
    .Y(_02393_));
 sg13g2_a21oi_1 _09951_ (.A1(net223),
    .A2(_02381_),
    .Y(_02394_),
    .B1(_02393_));
 sg13g2_o21ai_1 _09952_ (.B1(net71),
    .Y(_02395_),
    .A1(_02372_),
    .A2(_02394_));
 sg13g2_o21ai_1 _09953_ (.B1(_02395_),
    .Y(_00209_),
    .A1(_02348_),
    .A2(net38));
 sg13g2_buf_1 _09954_ (.A(\clock_inst.min_a[1] ),
    .X(_02396_));
 sg13g2_inv_1 _09955_ (.Y(_02397_),
    .A(_02396_));
 sg13g2_buf_1 _09956_ (.A(_02361_),
    .X(_02398_));
 sg13g2_nand2_1 _09957_ (.Y(_02399_),
    .A(_02182_),
    .B(net537));
 sg13g2_buf_2 _09958_ (.A(_02399_),
    .X(_02400_));
 sg13g2_buf_1 _09959_ (.A(net491),
    .X(_02401_));
 sg13g2_buf_1 _09960_ (.A(net419),
    .X(_02402_));
 sg13g2_buf_1 _09961_ (.A(net329),
    .X(_02403_));
 sg13g2_a21oi_1 _09962_ (.A1(net330),
    .A2(_02400_),
    .Y(_02404_),
    .B1(net218));
 sg13g2_buf_1 _09963_ (.A(net489),
    .X(_02405_));
 sg13g2_buf_1 _09964_ (.A(net418),
    .X(_02406_));
 sg13g2_buf_1 _09965_ (.A(net328),
    .X(_02407_));
 sg13g2_o21ai_1 _09966_ (.B1(net217),
    .Y(_02408_),
    .A1(net229),
    .A2(_02404_));
 sg13g2_buf_1 _09967_ (.A(net481),
    .X(_02409_));
 sg13g2_buf_1 _09968_ (.A(net417),
    .X(_02410_));
 sg13g2_buf_1 _09969_ (.A(net490),
    .X(_02411_));
 sg13g2_nand2_2 _09970_ (.Y(_02412_),
    .A(net482),
    .B(net539));
 sg13g2_nand2_2 _09971_ (.Y(_02413_),
    .A(_02334_),
    .B(_02206_));
 sg13g2_o21ai_1 _09972_ (.B1(_02413_),
    .Y(_02414_),
    .A1(net416),
    .A2(_02412_));
 sg13g2_buf_1 _09973_ (.A(net431),
    .X(_02415_));
 sg13g2_buf_1 _09974_ (.A(_02356_),
    .X(_02416_));
 sg13g2_nand2_2 _09975_ (.Y(_02417_),
    .A(_02192_),
    .B(net433));
 sg13g2_buf_1 _09976_ (.A(net419),
    .X(_02418_));
 sg13g2_nor2_1 _09977_ (.A(net324),
    .B(_02353_),
    .Y(_02419_));
 sg13g2_a21oi_1 _09978_ (.A1(_02213_),
    .A2(_02417_),
    .Y(_02420_),
    .B1(_02419_));
 sg13g2_a22oi_1 _09979_ (.Y(_02421_),
    .B1(_02375_),
    .B2(_02294_),
    .A2(net337),
    .A1(net422));
 sg13g2_or2_1 _09980_ (.X(_02422_),
    .B(_02421_),
    .A(net418));
 sg13g2_o21ai_1 _09981_ (.B1(_02422_),
    .Y(_02423_),
    .A1(net325),
    .A2(_02420_));
 sg13g2_a221oi_1 _09982_ (.B2(net326),
    .C1(_02423_),
    .B1(_02414_),
    .A1(_02410_),
    .Y(_02424_),
    .A2(net229));
 sg13g2_nor3_2 _09983_ (.A(net513),
    .B(_02252_),
    .C(_02256_),
    .Y(_02425_));
 sg13g2_o21ai_1 _09984_ (.B1(_02425_),
    .Y(_02426_),
    .A1(net343),
    .A2(_02385_));
 sg13g2_buf_1 _09985_ (.A(_02426_),
    .X(_02427_));
 sg13g2_a21oi_1 _09986_ (.A1(_02408_),
    .A2(_02424_),
    .Y(_02428_),
    .B1(_02427_));
 sg13g2_a21oi_1 _09987_ (.A1(_02397_),
    .A2(net39),
    .Y(_00210_),
    .B1(_02428_));
 sg13g2_buf_1 _09988_ (.A(net73),
    .X(_02429_));
 sg13g2_buf_1 _09989_ (.A(net228),
    .X(_02430_));
 sg13g2_buf_1 _09990_ (.A(net489),
    .X(_02431_));
 sg13g2_buf_1 _09991_ (.A(net415),
    .X(_02432_));
 sg13g2_nand2_1 _09992_ (.Y(_02433_),
    .A(_02323_),
    .B(_02212_));
 sg13g2_buf_1 _09993_ (.A(_02433_),
    .X(_02434_));
 sg13g2_nor2_1 _09994_ (.A(net424),
    .B(net216),
    .Y(_02435_));
 sg13g2_buf_1 _09995_ (.A(net494),
    .X(_02436_));
 sg13g2_buf_1 _09996_ (.A(net414),
    .X(_02437_));
 sg13g2_nand2_1 _09997_ (.Y(_02438_),
    .A(net534),
    .B(net438));
 sg13g2_buf_2 _09998_ (.A(_02438_),
    .X(_02439_));
 sg13g2_nand2_2 _09999_ (.Y(_02440_),
    .A(_02433_),
    .B(_02439_));
 sg13g2_nor2_1 _10000_ (.A(_02437_),
    .B(_02440_),
    .Y(_02441_));
 sg13g2_buf_1 _10001_ (.A(net351),
    .X(_02442_));
 sg13g2_o21ai_1 _10002_ (.B1(net215),
    .Y(_02443_),
    .A1(_02435_),
    .A2(_02441_));
 sg13g2_o21ai_1 _10003_ (.B1(_02443_),
    .Y(_02444_),
    .A1(net323),
    .A2(net330));
 sg13g2_nor2_1 _10004_ (.A(net488),
    .B(net352),
    .Y(_02445_));
 sg13g2_a21oi_1 _10005_ (.A1(net325),
    .A2(_02445_),
    .Y(_02446_),
    .B1(_02181_));
 sg13g2_nand2_1 _10006_ (.Y(_02447_),
    .A(net495),
    .B(net493));
 sg13g2_buf_1 _10007_ (.A(_02447_),
    .X(_02448_));
 sg13g2_nand2_1 _10008_ (.Y(_02449_),
    .A(net324),
    .B(net321));
 sg13g2_nand2_1 _10009_ (.Y(_02450_),
    .A(net433),
    .B(_02387_));
 sg13g2_a21oi_1 _10010_ (.A1(_02449_),
    .A2(_02450_),
    .Y(_02451_),
    .B1(net428));
 sg13g2_buf_2 _10011_ (.A(net433),
    .X(_02452_));
 sg13g2_nand2_2 _10012_ (.Y(_02453_),
    .A(net534),
    .B(net538));
 sg13g2_buf_1 _10013_ (.A(net490),
    .X(_02454_));
 sg13g2_a21oi_1 _10014_ (.A1(net320),
    .A2(_02453_),
    .Y(_02455_),
    .B1(net413));
 sg13g2_buf_1 _10015_ (.A(net432),
    .X(_02456_));
 sg13g2_o21ai_1 _10016_ (.B1(net319),
    .Y(_02457_),
    .A1(_02451_),
    .A2(_02455_));
 sg13g2_o21ai_1 _10017_ (.B1(_02457_),
    .Y(_02458_),
    .A1(net223),
    .A2(_02446_));
 sg13g2_a21oi_1 _10018_ (.A1(net133),
    .A2(_02444_),
    .Y(_02459_),
    .B1(_02458_));
 sg13g2_buf_1 _10019_ (.A(\clock_inst.min_a[20] ),
    .X(_02460_));
 sg13g2_nand2_1 _10020_ (.Y(_02461_),
    .A(_02460_),
    .B(net40));
 sg13g2_o21ai_1 _10021_ (.B1(_02461_),
    .Y(_00211_),
    .A1(net37),
    .A2(_02459_));
 sg13g2_buf_1 _10022_ (.A(net428),
    .X(_02462_));
 sg13g2_buf_1 _10023_ (.A(net318),
    .X(_02463_));
 sg13g2_nand2_1 _10024_ (.Y(_02464_),
    .A(net340),
    .B(net332));
 sg13g2_buf_1 _10025_ (.A(_02330_),
    .X(_02465_));
 sg13g2_nand2_1 _10026_ (.Y(_02466_),
    .A(net329),
    .B(net317));
 sg13g2_a21oi_1 _10027_ (.A1(_02464_),
    .A2(_02466_),
    .Y(_02467_),
    .B1(_02303_));
 sg13g2_nand2_1 _10028_ (.Y(_02468_),
    .A(net498),
    .B(net537));
 sg13g2_buf_1 _10029_ (.A(_02468_),
    .X(_02469_));
 sg13g2_nand2_1 _10030_ (.Y(_02470_),
    .A(net424),
    .B(net329));
 sg13g2_a21oi_1 _10031_ (.A1(net431),
    .A2(net316),
    .Y(_02471_),
    .B1(_02470_));
 sg13g2_nand2_1 _10032_ (.Y(_02472_),
    .A(net491),
    .B(net487));
 sg13g2_buf_1 _10033_ (.A(_02472_),
    .X(_02473_));
 sg13g2_nand2_1 _10034_ (.Y(_02474_),
    .A(net427),
    .B(_02159_));
 sg13g2_buf_1 _10035_ (.A(net320),
    .X(_02475_));
 sg13g2_a21oi_1 _10036_ (.A1(net315),
    .A2(_02474_),
    .Y(_02476_),
    .B1(net213));
 sg13g2_nor3_1 _10037_ (.A(_02467_),
    .B(_02471_),
    .C(_02476_),
    .Y(_02477_));
 sg13g2_buf_1 _10038_ (.A(net320),
    .X(_02478_));
 sg13g2_nor2_1 _10039_ (.A(net324),
    .B(_02260_),
    .Y(_02479_));
 sg13g2_nor2_2 _10040_ (.A(net437),
    .B(net438),
    .Y(_02480_));
 sg13g2_buf_1 _10041_ (.A(net486),
    .X(_02481_));
 sg13g2_o21ai_1 _10042_ (.B1(net412),
    .Y(_02482_),
    .A1(_02479_),
    .A2(_02480_));
 sg13g2_buf_1 _10043_ (.A(_02336_),
    .X(_02483_));
 sg13g2_nand2_1 _10044_ (.Y(_02484_),
    .A(net322),
    .B(net211));
 sg13g2_nand2_1 _10045_ (.Y(_02485_),
    .A(_02482_),
    .B(_02484_));
 sg13g2_buf_1 _10046_ (.A(net429),
    .X(_02486_));
 sg13g2_nand2_1 _10047_ (.Y(_02487_),
    .A(_02162_),
    .B(_02226_));
 sg13g2_buf_1 _10048_ (.A(_02487_),
    .X(_02488_));
 sg13g2_nor2_1 _10049_ (.A(net496),
    .B(net313),
    .Y(_02489_));
 sg13g2_a21oi_1 _10050_ (.A1(net340),
    .A2(net332),
    .Y(_02490_),
    .B1(_02489_));
 sg13g2_buf_1 _10051_ (.A(_02208_),
    .X(_02491_));
 sg13g2_buf_1 _10052_ (.A(_02387_),
    .X(_02492_));
 sg13g2_a221oi_1 _10053_ (.B2(net421),
    .C1(net226),
    .B1(net312),
    .A1(net322),
    .Y(_02493_),
    .A2(net411));
 sg13g2_o21ai_1 _10054_ (.B1(_02493_),
    .Y(_02494_),
    .A1(net314),
    .A2(_02490_));
 sg13g2_o21ai_1 _10055_ (.B1(_02494_),
    .Y(_02495_),
    .A1(net212),
    .A2(_02485_));
 sg13g2_o21ai_1 _10056_ (.B1(_02495_),
    .Y(_02496_),
    .A1(net214),
    .A2(_02477_));
 sg13g2_buf_2 _10057_ (.A(\clock_inst.min_a[21] ),
    .X(_02497_));
 sg13g2_nand2_1 _10058_ (.Y(_02498_),
    .A(_02497_),
    .B(net40));
 sg13g2_o21ai_1 _10059_ (.B1(_02498_),
    .Y(_00212_),
    .A1(net37),
    .A2(_02496_));
 sg13g2_buf_1 _10060_ (.A(\clock_inst.min_a[22] ),
    .X(_02499_));
 sg13g2_nor2_1 _10061_ (.A(net484),
    .B(net487),
    .Y(_02500_));
 sg13g2_buf_1 _10062_ (.A(_02500_),
    .X(_02501_));
 sg13g2_nand2_1 _10063_ (.Y(_02502_),
    .A(net536),
    .B(net430));
 sg13g2_buf_1 _10064_ (.A(_02502_),
    .X(_02503_));
 sg13g2_nand2_2 _10065_ (.Y(_02504_),
    .A(net486),
    .B(_02208_));
 sg13g2_o21ai_1 _10066_ (.B1(_02504_),
    .Y(_02505_),
    .A1(net311),
    .A2(net210));
 sg13g2_nor2_1 _10067_ (.A(net484),
    .B(_02214_),
    .Y(_02506_));
 sg13g2_buf_2 _10068_ (.A(_02506_),
    .X(_02507_));
 sg13g2_nor2_1 _10069_ (.A(net536),
    .B(net438),
    .Y(_02508_));
 sg13g2_buf_1 _10070_ (.A(net324),
    .X(_02509_));
 sg13g2_o21ai_1 _10071_ (.B1(net209),
    .Y(_02510_),
    .A1(_02507_),
    .A2(_02508_));
 sg13g2_nand2_1 _10072_ (.Y(_02511_),
    .A(net416),
    .B(_02439_));
 sg13g2_nor2_1 _10073_ (.A(_02292_),
    .B(net571),
    .Y(_02512_));
 sg13g2_buf_2 _10074_ (.A(_02512_),
    .X(_02513_));
 sg13g2_nand2_1 _10075_ (.Y(_02514_),
    .A(net230),
    .B(_02513_));
 sg13g2_nand3_1 _10076_ (.B(_02511_),
    .C(_02514_),
    .A(_02510_),
    .Y(_02515_));
 sg13g2_buf_1 _10077_ (.A(net435),
    .X(_02516_));
 sg13g2_buf_1 _10078_ (.A(net310),
    .X(_02517_));
 sg13g2_nor2_2 _10079_ (.A(net480),
    .B(_02233_),
    .Y(_02518_));
 sg13g2_a221oi_1 _10080_ (.B2(net208),
    .C1(_02518_),
    .B1(_02515_),
    .A1(net133),
    .Y(_02519_),
    .A2(_02505_));
 sg13g2_mux2_1 _10081_ (.A0(_02499_),
    .A1(_02519_),
    .S(net38),
    .X(_00213_));
 sg13g2_buf_1 _10082_ (.A(net72),
    .X(_02520_));
 sg13g2_nor2_1 _10083_ (.A(_02321_),
    .B(_02317_),
    .Y(_02521_));
 sg13g2_nand2_1 _10084_ (.Y(_02522_),
    .A(_02154_),
    .B(net541));
 sg13g2_buf_1 _10085_ (.A(_02522_),
    .X(_02523_));
 sg13g2_a21oi_1 _10086_ (.A1(net416),
    .A2(net410),
    .Y(_02524_),
    .B1(net213));
 sg13g2_o21ai_1 _10087_ (.B1(net337),
    .Y(_02525_),
    .A1(_02521_),
    .A2(_02524_));
 sg13g2_nand2_1 _10088_ (.Y(_02526_),
    .A(net430),
    .B(net538));
 sg13g2_buf_1 _10089_ (.A(_02526_),
    .X(_02527_));
 sg13g2_nand2_2 _10090_ (.Y(_02528_),
    .A(net437),
    .B(_02507_));
 sg13g2_nand2_1 _10091_ (.Y(_02529_),
    .A(_02339_),
    .B(_02528_));
 sg13g2_nor2_2 _10092_ (.A(net498),
    .B(_02297_),
    .Y(_02530_));
 sg13g2_nor2_1 _10093_ (.A(net430),
    .B(_02260_),
    .Y(_02531_));
 sg13g2_buf_2 _10094_ (.A(_02531_),
    .X(_02532_));
 sg13g2_or2_1 _10095_ (.X(_02533_),
    .B(_02532_),
    .A(_02530_));
 sg13g2_a22oi_1 _10096_ (.Y(_02534_),
    .B1(_02533_),
    .B2(net354),
    .A2(_02529_),
    .A1(net207));
 sg13g2_buf_1 _10097_ (.A(_02170_),
    .X(_02535_));
 sg13g2_a21oi_1 _10098_ (.A1(_02525_),
    .A2(_02534_),
    .Y(_02536_),
    .B1(net70));
 sg13g2_a21o_1 _10099_ (.A2(net36),
    .A1(\clock_inst.min_a[23] ),
    .B1(_02536_),
    .X(_00214_));
 sg13g2_inv_1 _10100_ (.Y(_02537_),
    .A(\clock_inst.min_a[2] ));
 sg13g2_buf_1 _10101_ (.A(net73),
    .X(_02538_));
 sg13g2_buf_1 _10102_ (.A(_02260_),
    .X(_02539_));
 sg13g2_nor2_2 _10103_ (.A(net534),
    .B(net430),
    .Y(_02540_));
 sg13g2_a22oi_1 _10104_ (.Y(_02541_),
    .B1(_02540_),
    .B2(_02159_),
    .A2(_02324_),
    .A1(net414));
 sg13g2_nor2_1 _10105_ (.A(net206),
    .B(_02541_),
    .Y(_02542_));
 sg13g2_nor2_1 _10106_ (.A(_02258_),
    .B(_02542_),
    .Y(_02543_));
 sg13g2_buf_1 _10107_ (.A(_02432_),
    .X(_02544_));
 sg13g2_buf_1 _10108_ (.A(_02184_),
    .X(_02545_));
 sg13g2_nand2_1 _10109_ (.Y(_02546_),
    .A(net541),
    .B(net538));
 sg13g2_nand2_1 _10110_ (.Y(_02547_),
    .A(net481),
    .B(_02546_));
 sg13g2_buf_1 _10111_ (.A(net211),
    .X(_02548_));
 sg13g2_a21oi_1 _10112_ (.A1(net213),
    .A2(_02547_),
    .Y(_02549_),
    .B1(net132));
 sg13g2_buf_1 _10113_ (.A(_02509_),
    .X(_02550_));
 sg13g2_o21ai_1 _10114_ (.B1(net497),
    .Y(_02551_),
    .A1(net333),
    .A2(_02530_));
 sg13g2_nand3_1 _10115_ (.B(_02385_),
    .C(_02551_),
    .A(_02398_),
    .Y(_02552_));
 sg13g2_nand2_1 _10116_ (.Y(_02553_),
    .A(net131),
    .B(_02552_));
 sg13g2_o21ai_1 _10117_ (.B1(_02553_),
    .Y(_02554_),
    .A1(net309),
    .A2(_02549_));
 sg13g2_nor2_1 _10118_ (.A(net534),
    .B(_02226_),
    .Y(_02555_));
 sg13g2_buf_2 _10119_ (.A(_02555_),
    .X(_02556_));
 sg13g2_buf_1 _10120_ (.A(_02368_),
    .X(_02557_));
 sg13g2_buf_1 _10121_ (.A(net434),
    .X(_02558_));
 sg13g2_a21oi_1 _10122_ (.A1(_02434_),
    .A2(net204),
    .Y(_02559_),
    .B1(net308));
 sg13g2_o21ai_1 _10123_ (.B1(_02478_),
    .Y(_02560_),
    .A1(_02556_),
    .A2(_02559_));
 sg13g2_buf_1 _10124_ (.A(_02311_),
    .X(_02561_));
 sg13g2_o21ai_1 _10125_ (.B1(net497),
    .Y(_02562_),
    .A1(net307),
    .A2(net411));
 sg13g2_nand2_1 _10126_ (.Y(_02563_),
    .A(net349),
    .B(_02562_));
 sg13g2_a22oi_1 _10127_ (.Y(_02564_),
    .B1(_02563_),
    .B2(net228),
    .A2(net227),
    .A1(net132));
 sg13g2_nand3_1 _10128_ (.B(_02560_),
    .C(_02564_),
    .A(_02407_),
    .Y(_02565_));
 sg13g2_o21ai_1 _10129_ (.B1(_02565_),
    .Y(_02566_),
    .A1(net205),
    .A2(_02554_));
 sg13g2_a22oi_1 _10130_ (.Y(_00215_),
    .B1(_02543_),
    .B2(_02566_),
    .A2(net35),
    .A1(_02537_));
 sg13g2_buf_1 _10131_ (.A(\clock_inst.min_a[24] ),
    .X(_02567_));
 sg13g2_inv_1 _10132_ (.Y(_02568_),
    .A(net568));
 sg13g2_buf_1 _10133_ (.A(_02568_),
    .X(_02569_));
 sg13g2_buf_1 _10134_ (.A(net416),
    .X(_02570_));
 sg13g2_nor2_1 _10135_ (.A(net450),
    .B(net306),
    .Y(_02571_));
 sg13g2_nor2_1 _10136_ (.A(net419),
    .B(net438),
    .Y(_02572_));
 sg13g2_buf_2 _10137_ (.A(_02572_),
    .X(_02573_));
 sg13g2_nand2_1 _10138_ (.Y(_02574_),
    .A(net229),
    .B(_02573_));
 sg13g2_a22oi_1 _10139_ (.Y(_00216_),
    .B1(_02571_),
    .B2(_02574_),
    .A2(net35),
    .A1(_02569_));
 sg13g2_nand2_1 _10140_ (.Y(_02575_),
    .A(net329),
    .B(net348));
 sg13g2_buf_1 _10141_ (.A(net483),
    .X(_02576_));
 sg13g2_a22oi_1 _10142_ (.Y(_02577_),
    .B1(_02308_),
    .B2(net409),
    .A2(net310),
    .A1(net353));
 sg13g2_nor3_1 _10143_ (.A(net439),
    .B(net490),
    .C(net333),
    .Y(_02578_));
 sg13g2_nand2_1 _10144_ (.Y(_02579_),
    .A(net541),
    .B(net430));
 sg13g2_buf_1 _10145_ (.A(_02297_),
    .X(_02580_));
 sg13g2_nor2_1 _10146_ (.A(_02579_),
    .B(net408),
    .Y(_02581_));
 sg13g2_o21ai_1 _10147_ (.B1(net347),
    .Y(_02582_),
    .A1(_02578_),
    .A2(_02581_));
 sg13g2_o21ai_1 _10148_ (.B1(_02582_),
    .Y(_02583_),
    .A1(net344),
    .A2(_02577_));
 sg13g2_buf_1 _10149_ (.A(net423),
    .X(_02584_));
 sg13g2_buf_1 _10150_ (.A(net305),
    .X(_02585_));
 sg13g2_buf_2 _10151_ (.A(net203),
    .X(_02586_));
 sg13g2_o21ai_1 _10152_ (.B1(net414),
    .Y(_02587_),
    .A1(net539),
    .A2(net352));
 sg13g2_nand2_1 _10153_ (.Y(_02588_),
    .A(_02200_),
    .B(_02294_));
 sg13g2_buf_1 _10154_ (.A(_02266_),
    .X(_02589_));
 sg13g2_a21oi_1 _10155_ (.A1(_02587_),
    .A2(_02588_),
    .Y(_02590_),
    .B1(net202));
 sg13g2_a221oi_1 _10156_ (.B2(net130),
    .C1(_02590_),
    .B1(_02583_),
    .A1(_02287_),
    .Y(_02591_),
    .A2(_02575_));
 sg13g2_nand2_1 _10157_ (.Y(_02592_),
    .A(\clock_inst.min_a[36] ),
    .B(net40));
 sg13g2_o21ai_1 _10158_ (.B1(_02592_),
    .Y(_00217_),
    .A1(net37),
    .A2(_02591_));
 sg13g2_inv_1 _10159_ (.Y(_02593_),
    .A(\clock_inst.min_a[37] ));
 sg13g2_o21ai_1 _10160_ (.B1(net229),
    .Y(_02594_),
    .A1(net306),
    .A2(_02573_));
 sg13g2_nor2_1 _10161_ (.A(net480),
    .B(net352),
    .Y(_02595_));
 sg13g2_nand2_1 _10162_ (.Y(_02596_),
    .A(net491),
    .B(_02208_));
 sg13g2_nand2_1 _10163_ (.Y(_02597_),
    .A(_02387_),
    .B(_02301_));
 sg13g2_a21o_1 _10164_ (.A2(_02597_),
    .A1(_02596_),
    .B1(net320),
    .X(_02598_));
 sg13g2_o21ai_1 _10165_ (.B1(_02598_),
    .Y(_02599_),
    .A1(_02575_),
    .A2(_02595_));
 sg13g2_nor2_1 _10166_ (.A(net484),
    .B(net493),
    .Y(_02600_));
 sg13g2_buf_1 _10167_ (.A(_02600_),
    .X(_02601_));
 sg13g2_nor2_1 _10168_ (.A(_02383_),
    .B(net304),
    .Y(_02602_));
 sg13g2_o21ai_1 _10169_ (.B1(_02310_),
    .Y(_02603_),
    .A1(net439),
    .A2(_02602_));
 sg13g2_nand2_1 _10170_ (.Y(_02604_),
    .A(net341),
    .B(_02603_));
 sg13g2_nor2_1 _10171_ (.A(net534),
    .B(net538),
    .Y(_02605_));
 sg13g2_buf_1 _10172_ (.A(_02605_),
    .X(_02606_));
 sg13g2_nor2_1 _10173_ (.A(net305),
    .B(_02297_),
    .Y(_02607_));
 sg13g2_buf_1 _10174_ (.A(net434),
    .X(_02608_));
 sg13g2_o21ai_1 _10175_ (.B1(net303),
    .Y(_02609_),
    .A1(net407),
    .A2(_02607_));
 sg13g2_buf_1 _10176_ (.A(net435),
    .X(_02610_));
 sg13g2_o21ai_1 _10177_ (.B1(net302),
    .Y(_02611_),
    .A1(net340),
    .A2(net312));
 sg13g2_nand4_1 _10178_ (.B(_02604_),
    .C(_02609_),
    .A(net319),
    .Y(_02612_),
    .D(_02611_));
 sg13g2_o21ai_1 _10179_ (.B1(_02612_),
    .Y(_02613_),
    .A1(net338),
    .A2(_02599_));
 sg13g2_nand3_1 _10180_ (.B(_02594_),
    .C(_02613_),
    .A(net71),
    .Y(_02614_));
 sg13g2_o21ai_1 _10181_ (.B1(_02614_),
    .Y(_00218_),
    .A1(_02593_),
    .A2(net38));
 sg13g2_nand2_1 _10182_ (.Y(_02615_),
    .A(net434),
    .B(net490));
 sg13g2_o21ai_1 _10183_ (.B1(_02615_),
    .Y(_02616_),
    .A1(net308),
    .A2(net313));
 sg13g2_nor2_1 _10184_ (.A(net336),
    .B(_02453_),
    .Y(_02617_));
 sg13g2_a221oi_1 _10185_ (.B2(net323),
    .C1(_02617_),
    .B1(_02616_),
    .A1(net228),
    .Y(_02618_),
    .A2(net407));
 sg13g2_nor2_2 _10186_ (.A(net492),
    .B(net481),
    .Y(_02619_));
 sg13g2_nor3_1 _10187_ (.A(net322),
    .B(net311),
    .C(_02619_),
    .Y(_02620_));
 sg13g2_a21oi_1 _10188_ (.A1(net314),
    .A2(net335),
    .Y(_02621_),
    .B1(_02620_));
 sg13g2_nor2_1 _10189_ (.A(net541),
    .B(net498),
    .Y(_02622_));
 sg13g2_nand2_1 _10190_ (.Y(_02623_),
    .A(net490),
    .B(_02622_));
 sg13g2_a21oi_1 _10191_ (.A1(net434),
    .A2(net321),
    .Y(_02624_),
    .B1(_02400_));
 sg13g2_a21oi_1 _10192_ (.A1(net435),
    .A2(net206),
    .Y(_02625_),
    .B1(_02255_));
 sg13g2_o21ai_1 _10193_ (.B1(net347),
    .Y(_02626_),
    .A1(_02624_),
    .A2(_02625_));
 sg13g2_nand2_1 _10194_ (.Y(_02627_),
    .A(_02623_),
    .B(_02626_));
 sg13g2_a21oi_1 _10195_ (.A1(net202),
    .A2(_02621_),
    .Y(_02628_),
    .B1(_02627_));
 sg13g2_o21ai_1 _10196_ (.B1(_02628_),
    .Y(_02629_),
    .A1(net215),
    .A2(_02618_));
 sg13g2_buf_2 _10197_ (.A(\clock_inst.min_a[38] ),
    .X(_02630_));
 sg13g2_nand2_1 _10198_ (.Y(_02631_),
    .A(_02630_),
    .B(net40));
 sg13g2_o21ai_1 _10199_ (.B1(_02631_),
    .Y(_00219_),
    .A1(_02429_),
    .A2(_02629_));
 sg13g2_nand2_1 _10200_ (.Y(_02632_),
    .A(net484),
    .B(_02189_));
 sg13g2_buf_2 _10201_ (.A(_02632_),
    .X(_02633_));
 sg13g2_nor2_1 _10202_ (.A(net494),
    .B(_02173_),
    .Y(_02634_));
 sg13g2_buf_2 _10203_ (.A(_02634_),
    .X(_02635_));
 sg13g2_a21o_1 _10204_ (.A2(_02635_),
    .A1(_02633_),
    .B1(_02284_),
    .X(_02636_));
 sg13g2_nor2b_1 _10205_ (.A(_02413_),
    .B_N(_02412_),
    .Y(_02637_));
 sg13g2_a21oi_1 _10206_ (.A1(net134),
    .A2(_02636_),
    .Y(_02638_),
    .B1(_02637_));
 sg13g2_buf_1 _10207_ (.A(net419),
    .X(_02639_));
 sg13g2_o21ai_1 _10208_ (.B1(net427),
    .Y(_02640_),
    .A1(net301),
    .A2(_02556_));
 sg13g2_nor2_1 _10209_ (.A(net418),
    .B(_02369_),
    .Y(_02641_));
 sg13g2_nor2_2 _10210_ (.A(net437),
    .B(net480),
    .Y(_02642_));
 sg13g2_nand2_1 _10211_ (.Y(_02643_),
    .A(net348),
    .B(net313));
 sg13g2_a22oi_1 _10212_ (.Y(_02644_),
    .B1(_02643_),
    .B2(net303),
    .A2(net332),
    .A1(_02642_));
 sg13g2_a22oi_1 _10213_ (.Y(_02645_),
    .B1(_02644_),
    .B2(net328),
    .A2(_02641_),
    .A1(_02640_));
 sg13g2_nor2_1 _10214_ (.A(net414),
    .B(_02273_),
    .Y(_02646_));
 sg13g2_o21ai_1 _10215_ (.B1(net412),
    .Y(_02647_),
    .A1(net427),
    .A2(_02646_));
 sg13g2_nor2_1 _10216_ (.A(net536),
    .B(net419),
    .Y(_02648_));
 sg13g2_buf_1 _10217_ (.A(_02648_),
    .X(_02649_));
 sg13g2_nand2_1 _10218_ (.Y(_02650_),
    .A(net407),
    .B(net201));
 sg13g2_nand3_1 _10219_ (.B(_02647_),
    .C(_02650_),
    .A(net212),
    .Y(_02651_));
 sg13g2_o21ai_1 _10220_ (.B1(_02651_),
    .Y(_02652_),
    .A1(_02478_),
    .A2(_02645_));
 sg13g2_o21ai_1 _10221_ (.B1(_02652_),
    .Y(_02653_),
    .A1(_02570_),
    .A2(_02638_));
 sg13g2_buf_2 _10222_ (.A(\clock_inst.min_a[39] ),
    .X(_02654_));
 sg13g2_nand2_1 _10223_ (.Y(_02655_),
    .A(_02654_),
    .B(net40));
 sg13g2_o21ai_1 _10224_ (.B1(_02655_),
    .Y(_00220_),
    .A1(_02429_),
    .A2(_02653_));
 sg13g2_inv_1 _10225_ (.Y(_02656_),
    .A(\clock_inst.min_a[3] ));
 sg13g2_nand2_1 _10226_ (.Y(_02657_),
    .A(net482),
    .B(_02211_));
 sg13g2_nor2_1 _10227_ (.A(net419),
    .B(net498),
    .Y(_02658_));
 sg13g2_buf_2 _10228_ (.A(_02658_),
    .X(_02659_));
 sg13g2_nor2_2 _10229_ (.A(_02192_),
    .B(net488),
    .Y(_02660_));
 sg13g2_nor2_2 _10230_ (.A(_02508_),
    .B(_02660_),
    .Y(_02661_));
 sg13g2_nand2_1 _10231_ (.Y(_02662_),
    .A(_02659_),
    .B(_02661_));
 sg13g2_o21ai_1 _10232_ (.B1(_02662_),
    .Y(_02663_),
    .A1(_02573_),
    .A2(_02657_));
 sg13g2_buf_2 _10233_ (.A(net341),
    .X(_02664_));
 sg13g2_nand2_1 _10234_ (.Y(_02665_),
    .A(net324),
    .B(net333));
 sg13g2_a21oi_1 _10235_ (.A1(_02388_),
    .A2(_02665_),
    .Y(_02666_),
    .B1(net328));
 sg13g2_a221oi_1 _10236_ (.B2(net200),
    .C1(_02666_),
    .B1(_02663_),
    .A1(net339),
    .Y(_02667_),
    .A2(_02635_));
 sg13g2_nand2b_1 _10237_ (.Y(_02668_),
    .B(net214),
    .A_N(_02667_));
 sg13g2_nand2_2 _10238_ (.Y(_02669_),
    .A(net430),
    .B(_02336_));
 sg13g2_nand2_2 _10239_ (.Y(_02670_),
    .A(net492),
    .B(net423));
 sg13g2_nor3_2 _10240_ (.A(net482),
    .B(_02669_),
    .C(_02670_),
    .Y(_02671_));
 sg13g2_a21oi_1 _10241_ (.A1(net321),
    .A2(net216),
    .Y(_02672_),
    .B1(net331));
 sg13g2_nor2_2 _10242_ (.A(_02173_),
    .B(_02310_),
    .Y(_02673_));
 sg13g2_a21oi_1 _10243_ (.A1(net427),
    .A2(_02670_),
    .Y(_02674_),
    .B1(_02417_));
 sg13g2_nor3_1 _10244_ (.A(_02672_),
    .B(_02673_),
    .C(_02674_),
    .Y(_02675_));
 sg13g2_nand2_1 _10245_ (.Y(_02676_),
    .A(_02292_),
    .B(_02176_));
 sg13g2_buf_1 _10246_ (.A(_02676_),
    .X(_02677_));
 sg13g2_nor2_1 _10247_ (.A(net491),
    .B(_02212_),
    .Y(_02678_));
 sg13g2_buf_2 _10248_ (.A(_02678_),
    .X(_02679_));
 sg13g2_nor4_1 _10249_ (.A(net417),
    .B(_02196_),
    .C(net300),
    .D(_02679_),
    .Y(_02680_));
 sg13g2_nor2_1 _10250_ (.A(_02258_),
    .B(_02680_),
    .Y(_02681_));
 sg13g2_o21ai_1 _10251_ (.B1(_02681_),
    .Y(_02682_),
    .A1(net200),
    .A2(_02675_));
 sg13g2_nor2_1 _10252_ (.A(_02671_),
    .B(_02682_),
    .Y(_02683_));
 sg13g2_a22oi_1 _10253_ (.Y(_00221_),
    .B1(_02668_),
    .B2(_02683_),
    .A2(_02538_),
    .A1(_02656_));
 sg13g2_o21ai_1 _10254_ (.B1(net413),
    .Y(_02684_),
    .A1(net227),
    .A2(_02573_));
 sg13g2_nand2_1 _10255_ (.Y(_02685_),
    .A(_02197_),
    .B(_02513_));
 sg13g2_nor2_1 _10256_ (.A(net347),
    .B(_02480_),
    .Y(_02686_));
 sg13g2_a22oi_1 _10257_ (.Y(_02687_),
    .B1(_02685_),
    .B2(_02686_),
    .A2(_02684_),
    .A1(net314));
 sg13g2_a21oi_1 _10258_ (.A1(net353),
    .A2(_02298_),
    .Y(_02688_),
    .B1(_02181_));
 sg13g2_nand2_2 _10259_ (.Y(_02689_),
    .A(net414),
    .B(_02191_));
 sg13g2_nand2_1 _10260_ (.Y(_02690_),
    .A(net210),
    .B(_02689_));
 sg13g2_nand2_1 _10261_ (.Y(_02691_),
    .A(net437),
    .B(_02195_));
 sg13g2_a21oi_1 _10262_ (.A1(net417),
    .A2(_02691_),
    .Y(_02692_),
    .B1(net351));
 sg13g2_a22oi_1 _10263_ (.Y(_02693_),
    .B1(_02692_),
    .B2(net425),
    .A2(_02690_),
    .A1(net209));
 sg13g2_o21ai_1 _10264_ (.B1(_02693_),
    .Y(_02694_),
    .A1(net323),
    .A2(_02688_));
 sg13g2_nand2_1 _10265_ (.Y(_02695_),
    .A(net412),
    .B(_02213_));
 sg13g2_a21oi_1 _10266_ (.A1(net338),
    .A2(net316),
    .Y(_02696_),
    .B1(_02695_));
 sg13g2_a221oi_1 _10267_ (.B2(net130),
    .C1(_02696_),
    .B1(_02694_),
    .A1(net215),
    .Y(_02697_),
    .A2(_02687_));
 sg13g2_buf_2 _10268_ (.A(\clock_inst.min_a[40] ),
    .X(_02698_));
 sg13g2_nand2_1 _10269_ (.Y(_02699_),
    .A(_02698_),
    .B(net40));
 sg13g2_o21ai_1 _10270_ (.B1(_02699_),
    .Y(_00222_),
    .A1(net37),
    .A2(_02697_));
 sg13g2_nor2_2 _10271_ (.A(net329),
    .B(net349),
    .Y(_02700_));
 sg13g2_o21ai_1 _10272_ (.B1(net202),
    .Y(_02701_),
    .A1(net229),
    .A2(_02700_));
 sg13g2_nor2_1 _10273_ (.A(net433),
    .B(_02326_),
    .Y(_02702_));
 sg13g2_o21ai_1 _10274_ (.B1(_02468_),
    .Y(_02703_),
    .A1(net421),
    .A2(_02702_));
 sg13g2_nand2_1 _10275_ (.Y(_02704_),
    .A(net349),
    .B(_02615_));
 sg13g2_a22oi_1 _10276_ (.Y(_02705_),
    .B1(_02704_),
    .B2(net325),
    .A2(_02703_),
    .A1(net218));
 sg13g2_nand2b_1 _10277_ (.Y(_02706_),
    .B(net224),
    .A_N(_02705_));
 sg13g2_nor2_2 _10278_ (.A(net539),
    .B(net537),
    .Y(_02707_));
 sg13g2_o21ai_1 _10279_ (.B1(net301),
    .Y(_02708_),
    .A1(_02235_),
    .A2(_02707_));
 sg13g2_a21oi_1 _10280_ (.A1(net204),
    .A2(_02708_),
    .Y(_02709_),
    .B1(_02475_));
 sg13g2_a21oi_1 _10281_ (.A1(net216),
    .A2(net330),
    .Y(_02710_),
    .B1(_02403_));
 sg13g2_buf_1 _10282_ (.A(net331),
    .X(_02711_));
 sg13g2_o21ai_1 _10283_ (.B1(net199),
    .Y(_02712_),
    .A1(_02709_),
    .A2(_02710_));
 sg13g2_nand3_1 _10284_ (.B(_02706_),
    .C(_02712_),
    .A(_02701_),
    .Y(_02713_));
 sg13g2_buf_1 _10285_ (.A(\clock_inst.min_a[41] ),
    .X(_02714_));
 sg13g2_nand2_1 _10286_ (.Y(_02715_),
    .A(_02714_),
    .B(net40));
 sg13g2_o21ai_1 _10287_ (.B1(_02715_),
    .Y(_00223_),
    .A1(net37),
    .A2(_02713_));
 sg13g2_buf_1 _10288_ (.A(net411),
    .X(_02716_));
 sg13g2_nor2_2 _10289_ (.A(_02401_),
    .B(net423),
    .Y(_02717_));
 sg13g2_nor2_1 _10290_ (.A(net428),
    .B(net316),
    .Y(_02718_));
 sg13g2_a21o_1 _10291_ (.A2(_02717_),
    .A1(net299),
    .B1(_02718_),
    .X(_02719_));
 sg13g2_nand2_1 _10292_ (.Y(_02720_),
    .A(net438),
    .B(net335));
 sg13g2_nor2_1 _10293_ (.A(net302),
    .B(_02720_),
    .Y(_02721_));
 sg13g2_nand2_1 _10294_ (.Y(_02722_),
    .A(net486),
    .B(_02229_));
 sg13g2_a21oi_1 _10295_ (.A1(net300),
    .A2(_02722_),
    .Y(_02723_),
    .B1(net415));
 sg13g2_nor3_1 _10296_ (.A(net218),
    .B(_02721_),
    .C(_02723_),
    .Y(_02724_));
 sg13g2_nor2_1 _10297_ (.A(_02217_),
    .B(net484),
    .Y(_02725_));
 sg13g2_buf_2 _10298_ (.A(_02725_),
    .X(_02726_));
 sg13g2_a21oi_1 _10299_ (.A1(net333),
    .A2(_02726_),
    .Y(_02727_),
    .B1(net307));
 sg13g2_nor2_1 _10300_ (.A(net341),
    .B(_02727_),
    .Y(_02728_));
 sg13g2_nor2_1 _10301_ (.A(net498),
    .B(_02208_),
    .Y(_02729_));
 sg13g2_mux2_1 _10302_ (.A0(_02526_),
    .A1(_02729_),
    .S(net482),
    .X(_02730_));
 sg13g2_nor2_1 _10303_ (.A(net428),
    .B(_02730_),
    .Y(_02731_));
 sg13g2_nor3_1 _10304_ (.A(net334),
    .B(_02728_),
    .C(_02731_),
    .Y(_02732_));
 sg13g2_nor2_1 _10305_ (.A(_02724_),
    .B(_02732_),
    .Y(_02733_));
 sg13g2_a221oi_1 _10306_ (.B2(net217),
    .C1(_02733_),
    .B1(_02719_),
    .A1(_02284_),
    .Y(_02734_),
    .A2(net220));
 sg13g2_buf_2 _10307_ (.A(\clock_inst.min_a[42] ),
    .X(_02735_));
 sg13g2_buf_1 _10308_ (.A(net72),
    .X(_02736_));
 sg13g2_nand2_1 _10309_ (.Y(_02737_),
    .A(_02735_),
    .B(net34));
 sg13g2_o21ai_1 _10310_ (.B1(_02737_),
    .Y(_00224_),
    .A1(net37),
    .A2(_02734_));
 sg13g2_buf_1 _10311_ (.A(\clock_inst.min_a[43] ),
    .X(_02738_));
 sg13g2_nand2_1 _10312_ (.Y(_02739_),
    .A(_02164_),
    .B(net571));
 sg13g2_buf_1 _10313_ (.A(_02739_),
    .X(_02740_));
 sg13g2_nor2_2 _10314_ (.A(net481),
    .B(net478),
    .Y(_02741_));
 sg13g2_o21ai_1 _10315_ (.B1(net429),
    .Y(_02742_),
    .A1(_02225_),
    .A2(_02213_));
 sg13g2_o21ai_1 _10316_ (.B1(_02742_),
    .Y(_02743_),
    .A1(net302),
    .A2(_02573_));
 sg13g2_nand2_2 _10317_ (.Y(_02744_),
    .A(net419),
    .B(net430));
 sg13g2_o21ai_1 _10318_ (.B1(_02744_),
    .Y(_02745_),
    .A1(_02523_),
    .A2(net330));
 sg13g2_buf_1 _10319_ (.A(net305),
    .X(_02746_));
 sg13g2_buf_1 _10320_ (.A(net198),
    .X(_02747_));
 sg13g2_a221oi_1 _10321_ (.B2(net231),
    .C1(net129),
    .B1(_02745_),
    .A1(net327),
    .Y(_02748_),
    .A2(_02743_));
 sg13g2_nor2_1 _10322_ (.A(net536),
    .B(net538),
    .Y(_02749_));
 sg13g2_buf_2 _10323_ (.A(_02749_),
    .X(_02750_));
 sg13g2_buf_1 _10324_ (.A(_02622_),
    .X(_02751_));
 sg13g2_o21ai_1 _10325_ (.B1(net298),
    .Y(_02752_),
    .A1(net413),
    .A2(_02750_));
 sg13g2_a21oi_1 _10326_ (.A1(_02557_),
    .A2(_02752_),
    .Y(_02753_),
    .B1(net309));
 sg13g2_nor4_1 _10327_ (.A(net72),
    .B(_02741_),
    .C(_02748_),
    .D(_02753_),
    .Y(_02754_));
 sg13g2_a21o_1 _10328_ (.A2(net36),
    .A1(_02738_),
    .B1(_02754_),
    .X(_00225_));
 sg13g2_nand2_1 _10329_ (.Y(_02755_),
    .A(net494),
    .B(_02203_));
 sg13g2_buf_2 _10330_ (.A(_02755_),
    .X(_02756_));
 sg13g2_nor2_1 _10331_ (.A(net426),
    .B(_02756_),
    .Y(_02757_));
 sg13g2_o21ai_1 _10332_ (.B1(_02516_),
    .Y(_02758_),
    .A1(net431),
    .A2(_02757_));
 sg13g2_o21ai_1 _10333_ (.B1(_02758_),
    .Y(_02759_),
    .A1(net410),
    .A2(net339));
 sg13g2_a21oi_1 _10334_ (.A1(_02239_),
    .A2(net298),
    .Y(_02760_),
    .B1(net416));
 sg13g2_o21ai_1 _10335_ (.B1(_02353_),
    .Y(_02761_),
    .A1(_02462_),
    .A2(_02760_));
 sg13g2_a221oi_1 _10336_ (.B2(_02272_),
    .C1(net132),
    .B1(_02761_),
    .A1(net214),
    .Y(_02762_),
    .A2(_02759_));
 sg13g2_buf_1 _10337_ (.A(\clock_inst.min_a[44] ),
    .X(_02763_));
 sg13g2_nand2_1 _10338_ (.Y(_02764_),
    .A(_02763_),
    .B(net34));
 sg13g2_o21ai_1 _10339_ (.B1(_02764_),
    .Y(_00226_),
    .A1(net37),
    .A2(_02762_));
 sg13g2_buf_1 _10340_ (.A(\clock_inst.min_a[4] ),
    .X(_02765_));
 sg13g2_inv_1 _10341_ (.Y(_02766_),
    .A(_02765_));
 sg13g2_buf_1 _10342_ (.A(net307),
    .X(_02767_));
 sg13g2_a21oi_1 _10343_ (.A1(net336),
    .A2(net220),
    .Y(_02768_),
    .B1(net197));
 sg13g2_nand2_2 _10344_ (.Y(_02769_),
    .A(net486),
    .B(net333));
 sg13g2_a21o_1 _10345_ (.A2(_02769_),
    .A1(net216),
    .B1(_02322_),
    .X(_02770_));
 sg13g2_o21ai_1 _10346_ (.B1(_02770_),
    .Y(_02771_),
    .A1(_02545_),
    .A2(_02768_));
 sg13g2_buf_1 _10347_ (.A(_02229_),
    .X(_02772_));
 sg13g2_buf_1 _10348_ (.A(net297),
    .X(_02773_));
 sg13g2_nor2_1 _10349_ (.A(_02436_),
    .B(_02330_),
    .Y(_02774_));
 sg13g2_o21ai_1 _10350_ (.B1(_02242_),
    .Y(_02775_),
    .A1(_02773_),
    .A2(_02774_));
 sg13g2_o21ai_1 _10351_ (.B1(_02379_),
    .Y(_02776_),
    .A1(_02416_),
    .A2(_02660_));
 sg13g2_a21oi_1 _10352_ (.A1(_02775_),
    .A2(_02776_),
    .Y(_02777_),
    .B1(net223));
 sg13g2_a21oi_1 _10353_ (.A1(_02430_),
    .A2(_02771_),
    .Y(_02778_),
    .B1(_02777_));
 sg13g2_and2_1 _10354_ (.A(_02284_),
    .B(_02326_),
    .X(_02779_));
 sg13g2_a21oi_1 _10355_ (.A1(net208),
    .A2(_02779_),
    .Y(_02780_),
    .B1(_02427_));
 sg13g2_a22oi_1 _10356_ (.Y(_00227_),
    .B1(_02778_),
    .B2(_02780_),
    .A2(_02538_),
    .A1(_02766_));
 sg13g2_buf_1 _10357_ (.A(\clock_inst.min_a[45] ),
    .X(_02781_));
 sg13g2_inv_1 _10358_ (.Y(_02782_),
    .A(_02781_));
 sg13g2_buf_1 _10359_ (.A(net72),
    .X(_02783_));
 sg13g2_a21oi_1 _10360_ (.A1(net230),
    .A2(net342),
    .Y(_02784_),
    .B1(_02266_));
 sg13g2_o21ai_1 _10361_ (.B1(net221),
    .Y(_02785_),
    .A1(_02286_),
    .A2(_02175_));
 sg13g2_o21ai_1 _10362_ (.B1(_02785_),
    .Y(_02786_),
    .A1(_02570_),
    .A2(_02784_));
 sg13g2_nor2_1 _10363_ (.A(net33),
    .B(_02786_),
    .Y(_02787_));
 sg13g2_a21oi_1 _10364_ (.A1(net533),
    .A2(net39),
    .Y(_00228_),
    .B1(_02787_));
 sg13g2_buf_1 _10365_ (.A(\clock_inst.min_a[5] ),
    .X(_02788_));
 sg13g2_inv_1 _10366_ (.Y(_02789_),
    .A(_02788_));
 sg13g2_nand2_1 _10367_ (.Y(_02790_),
    .A(_02162_),
    .B(_02165_));
 sg13g2_buf_2 _10368_ (.A(_02790_),
    .X(_02791_));
 sg13g2_nand2_1 _10369_ (.Y(_02792_),
    .A(_02186_),
    .B(_02540_));
 sg13g2_o21ai_1 _10370_ (.B1(_02792_),
    .Y(_02793_),
    .A1(_02334_),
    .A2(_02791_));
 sg13g2_a22oi_1 _10371_ (.Y(_02794_),
    .B1(_02793_),
    .B2(net432),
    .A2(net201),
    .A1(net222));
 sg13g2_nor2_2 _10372_ (.A(_02323_),
    .B(_02361_),
    .Y(_02795_));
 sg13g2_nand2_1 _10373_ (.Y(_02796_),
    .A(_02635_),
    .B(_02795_));
 sg13g2_o21ai_1 _10374_ (.B1(_02796_),
    .Y(_02797_),
    .A1(net200),
    .A2(_02794_));
 sg13g2_nor2_1 _10375_ (.A(net345),
    .B(net300),
    .Y(_02798_));
 sg13g2_a221oi_1 _10376_ (.B2(_02175_),
    .C1(_02258_),
    .B1(_02798_),
    .A1(net134),
    .Y(_02799_),
    .A2(_02797_));
 sg13g2_nand2_2 _10377_ (.Y(_02800_),
    .A(net540),
    .B(net493));
 sg13g2_nand2_2 _10378_ (.Y(_02801_),
    .A(net480),
    .B(_02200_));
 sg13g2_o21ai_1 _10379_ (.B1(_02801_),
    .Y(_02802_),
    .A1(net497),
    .A2(_02800_));
 sg13g2_a22oi_1 _10380_ (.Y(_02803_),
    .B1(_02802_),
    .B2(net353),
    .A2(net221),
    .A1(net342));
 sg13g2_or2_1 _10381_ (.X(_02804_),
    .B(_02803_),
    .A(net319));
 sg13g2_nor2_1 _10382_ (.A(net206),
    .B(_02413_),
    .Y(_02805_));
 sg13g2_o21ai_1 _10383_ (.B1(net323),
    .Y(_02806_),
    .A1(_02354_),
    .A2(_02805_));
 sg13g2_nand2_1 _10384_ (.Y(_02807_),
    .A(_02320_),
    .B(net305));
 sg13g2_a22oi_1 _10385_ (.Y(_02808_),
    .B1(_02659_),
    .B2(_02807_),
    .A2(net342),
    .A1(net329));
 sg13g2_nor2_1 _10386_ (.A(net413),
    .B(_02808_),
    .Y(_02809_));
 sg13g2_nand3_1 _10387_ (.B(_02579_),
    .C(_02317_),
    .A(_02320_),
    .Y(_02810_));
 sg13g2_a21oi_1 _10388_ (.A1(_02689_),
    .A2(_02810_),
    .Y(_02811_),
    .B1(net412));
 sg13g2_o21ai_1 _10389_ (.B1(net326),
    .Y(_02812_),
    .A1(_02809_),
    .A2(_02811_));
 sg13g2_and4_1 _10390_ (.A(_02385_),
    .B(_02804_),
    .C(_02806_),
    .D(_02812_),
    .X(_02813_));
 sg13g2_a22oi_1 _10391_ (.Y(_00229_),
    .B1(_02799_),
    .B2(_02813_),
    .A2(net35),
    .A1(_02789_));
 sg13g2_buf_1 _10392_ (.A(\clock_inst.min_a[6] ),
    .X(_02814_));
 sg13g2_inv_1 _10393_ (.Y(_02815_),
    .A(_02814_));
 sg13g2_buf_1 _10394_ (.A(net218),
    .X(_02816_));
 sg13g2_nand2_1 _10395_ (.Y(_02817_),
    .A(net536),
    .B(_02195_));
 sg13g2_nand2_1 _10396_ (.Y(_02818_),
    .A(net417),
    .B(_02817_));
 sg13g2_nand2_1 _10397_ (.Y(_02819_),
    .A(net488),
    .B(_02234_));
 sg13g2_o21ai_1 _10398_ (.B1(_02469_),
    .Y(_02820_),
    .A1(net409),
    .A2(_02819_));
 sg13g2_a22oi_1 _10399_ (.Y(_02821_),
    .B1(_02820_),
    .B2(net129),
    .A2(_02818_),
    .A1(net222));
 sg13g2_nor2_1 _10400_ (.A(net328),
    .B(_02439_),
    .Y(_02822_));
 sg13g2_a21oi_1 _10401_ (.A1(_02434_),
    .A2(_02557_),
    .Y(_02823_),
    .B1(net210));
 sg13g2_nor3_1 _10402_ (.A(net131),
    .B(_02822_),
    .C(_02823_),
    .Y(_02824_));
 sg13g2_a21o_1 _10403_ (.A2(_02821_),
    .A1(net128),
    .B1(_02824_),
    .X(_02825_));
 sg13g2_nand2_1 _10404_ (.Y(_02826_),
    .A(net436),
    .B(_02726_));
 sg13g2_nand2b_1 _10405_ (.Y(_02827_),
    .B(_02425_),
    .A_N(_02262_));
 sg13g2_nand2_2 _10406_ (.Y(_02828_),
    .A(net539),
    .B(_02336_));
 sg13g2_nor2_1 _10407_ (.A(net410),
    .B(_02828_),
    .Y(_02829_));
 sg13g2_nor2_1 _10408_ (.A(_02779_),
    .B(_02829_),
    .Y(_02830_));
 sg13g2_nor2_1 _10409_ (.A(net310),
    .B(_02830_),
    .Y(_02831_));
 sg13g2_nand2_1 _10410_ (.Y(_02832_),
    .A(net342),
    .B(_02336_));
 sg13g2_buf_1 _10411_ (.A(net439),
    .X(_02833_));
 sg13g2_a21oi_1 _10412_ (.A1(_02385_),
    .A2(_02832_),
    .Y(_02834_),
    .B1(net296));
 sg13g2_nor3_1 _10413_ (.A(_02827_),
    .B(_02831_),
    .C(_02834_),
    .Y(_02835_));
 sg13g2_and2_1 _10414_ (.A(_02826_),
    .B(_02835_),
    .X(_02836_));
 sg13g2_a22oi_1 _10415_ (.Y(_00230_),
    .B1(_02825_),
    .B2(_02836_),
    .A2(net35),
    .A1(_02815_));
 sg13g2_buf_1 _10416_ (.A(\clock_inst.min_a[7] ),
    .X(_02837_));
 sg13g2_inv_1 _10417_ (.Y(_02838_),
    .A(_02837_));
 sg13g2_nor2_1 _10418_ (.A(net480),
    .B(_02361_),
    .Y(_02839_));
 sg13g2_nand2_1 _10419_ (.Y(_02840_),
    .A(net335),
    .B(_02487_));
 sg13g2_nor2_1 _10420_ (.A(net212),
    .B(net230),
    .Y(_02841_));
 sg13g2_a22oi_1 _10421_ (.Y(_02842_),
    .B1(_02840_),
    .B2(_02841_),
    .A2(_02839_),
    .A1(_02756_));
 sg13g2_nor2_1 _10422_ (.A(net429),
    .B(_02556_),
    .Y(_02843_));
 sg13g2_a22oi_1 _10423_ (.Y(_02844_),
    .B1(_02801_),
    .B2(_02843_),
    .A2(net485),
    .A1(net331));
 sg13g2_nand2_1 _10424_ (.Y(_02845_),
    .A(net429),
    .B(_02772_));
 sg13g2_nand2_1 _10425_ (.Y(_02846_),
    .A(net330),
    .B(_02845_));
 sg13g2_a221oi_1 _10426_ (.B2(_02295_),
    .C1(_02718_),
    .B1(_02846_),
    .A1(_02278_),
    .Y(_02847_),
    .A2(_02844_));
 sg13g2_mux2_1 _10427_ (.A0(_02842_),
    .A1(_02847_),
    .S(net134),
    .X(_02848_));
 sg13g2_a22oi_1 _10428_ (.Y(_00231_),
    .B1(_02835_),
    .B2(_02848_),
    .A2(net35),
    .A1(_02838_));
 sg13g2_nor2_1 _10429_ (.A(_02273_),
    .B(_02750_),
    .Y(_02849_));
 sg13g2_o21ai_1 _10430_ (.B1(net206),
    .Y(_02850_),
    .A1(net485),
    .A2(_02849_));
 sg13g2_a21oi_1 _10431_ (.A1(_02442_),
    .A2(_02284_),
    .Y(_02851_),
    .B1(net206));
 sg13g2_a221oi_1 _10432_ (.B2(net133),
    .C1(_02851_),
    .B1(_02850_),
    .A1(_02589_),
    .Y(_02852_),
    .A2(_02275_));
 sg13g2_buf_1 _10433_ (.A(\clock_inst.min_a[8] ),
    .X(_02853_));
 sg13g2_nand2_1 _10434_ (.Y(_02854_),
    .A(net567),
    .B(net34));
 sg13g2_o21ai_1 _10435_ (.B1(_02854_),
    .Y(_00232_),
    .A1(net37),
    .A2(_02852_));
 sg13g2_buf_1 _10436_ (.A(\clock_inst.min_b[0] ),
    .X(_02855_));
 sg13g2_nand2_2 _10437_ (.Y(_02856_),
    .A(net433),
    .B(_02326_));
 sg13g2_nand2_1 _10438_ (.Y(_02857_),
    .A(_02230_),
    .B(net315));
 sg13g2_nand2_1 _10439_ (.Y(_02858_),
    .A(net437),
    .B(_02330_));
 sg13g2_a21oi_1 _10440_ (.A1(_02810_),
    .A2(_02858_),
    .Y(_02859_),
    .B1(net417));
 sg13g2_a21oi_1 _10441_ (.A1(_02661_),
    .A2(_02857_),
    .Y(_02860_),
    .B1(_02859_));
 sg13g2_o21ai_1 _10442_ (.B1(_02265_),
    .Y(_02861_),
    .A1(net329),
    .A2(_02468_));
 sg13g2_a221oi_1 _10443_ (.B2(net415),
    .C1(net440),
    .B1(_02861_),
    .A1(net225),
    .Y(_02862_),
    .A2(net315));
 sg13g2_a21o_1 _10444_ (.A2(_02860_),
    .A1(net318),
    .B1(_02862_),
    .X(_02863_));
 sg13g2_o21ai_1 _10445_ (.B1(_02863_),
    .Y(_02864_),
    .A1(_02470_),
    .A2(_02856_));
 sg13g2_mux2_1 _10446_ (.A0(_02855_),
    .A1(_02864_),
    .S(net38),
    .X(_00233_));
 sg13g2_buf_1 _10447_ (.A(\clock_inst.min_b[10] ),
    .X(_02865_));
 sg13g2_buf_1 _10448_ (.A(_02865_),
    .X(_02866_));
 sg13g2_nand2_1 _10449_ (.Y(_02867_),
    .A(_02584_),
    .B(_02280_));
 sg13g2_nand3_1 _10450_ (.B(_02268_),
    .C(_02465_),
    .A(net346),
    .Y(_02868_));
 sg13g2_o21ai_1 _10451_ (.B1(_02868_),
    .Y(_02869_),
    .A1(_02756_),
    .A2(_02867_));
 sg13g2_nor3_1 _10452_ (.A(net450),
    .B(net306),
    .C(_02869_),
    .Y(_02870_));
 sg13g2_a21o_1 _10453_ (.A2(net36),
    .A1(net532),
    .B1(_02870_),
    .X(_00234_));
 sg13g2_buf_1 _10454_ (.A(_02171_),
    .X(_02871_));
 sg13g2_a21oi_1 _10455_ (.A1(net336),
    .A2(_02204_),
    .Y(_02872_),
    .B1(_02700_));
 sg13g2_inv_1 _10456_ (.Y(_02873_),
    .A(_02872_));
 sg13g2_buf_1 _10457_ (.A(_02558_),
    .X(_02874_));
 sg13g2_nand2_1 _10458_ (.Y(_02875_),
    .A(_02791_),
    .B(_02676_));
 sg13g2_inv_1 _10459_ (.Y(_02876_),
    .A(_02875_));
 sg13g2_o21ai_1 _10460_ (.B1(net313),
    .Y(_02877_),
    .A1(_02238_),
    .A2(_02876_));
 sg13g2_or2_1 _10461_ (.X(_02878_),
    .B(_02795_),
    .A(_02354_));
 sg13g2_a22oi_1 _10462_ (.Y(_02879_),
    .B1(_02878_),
    .B2(net347),
    .A2(_02877_),
    .A1(net431));
 sg13g2_o21ai_1 _10463_ (.B1(_02828_),
    .Y(_02880_),
    .A1(net410),
    .A2(net335));
 sg13g2_nand2_2 _10464_ (.Y(_02881_),
    .A(net423),
    .B(_02326_));
 sg13g2_a21oi_1 _10465_ (.A1(_02337_),
    .A2(_02881_),
    .Y(_02882_),
    .B1(net432));
 sg13g2_o21ai_1 _10466_ (.B1(net213),
    .Y(_02883_),
    .A1(_02880_),
    .A2(_02882_));
 sg13g2_o21ai_1 _10467_ (.B1(_02883_),
    .Y(_02884_),
    .A1(net195),
    .A2(_02879_));
 sg13g2_a221oi_1 _10468_ (.B2(net407),
    .C1(_02884_),
    .B1(_02873_),
    .A1(_02530_),
    .Y(_02885_),
    .A2(_02717_));
 sg13g2_buf_2 _10469_ (.A(\clock_inst.min_b[19] ),
    .X(_02886_));
 sg13g2_nand2_1 _10470_ (.Y(_02887_),
    .A(_02886_),
    .B(_02736_));
 sg13g2_o21ai_1 _10471_ (.B1(_02887_),
    .Y(_00235_),
    .A1(_02871_),
    .A2(_02885_));
 sg13g2_nand2_1 _10472_ (.Y(_02888_),
    .A(net421),
    .B(net349));
 sg13g2_nand2_1 _10473_ (.Y(_02889_),
    .A(net305),
    .B(_02200_));
 sg13g2_a21oi_1 _10474_ (.A1(net478),
    .A2(_02889_),
    .Y(_02890_),
    .B1(_02406_));
 sg13g2_a21oi_1 _10475_ (.A1(_02888_),
    .A2(_02660_),
    .Y(_02891_),
    .B1(_02890_));
 sg13g2_nand2_2 _10476_ (.Y(_02892_),
    .A(net414),
    .B(net438));
 sg13g2_nand2_1 _10477_ (.Y(_02893_),
    .A(net215),
    .B(_02892_));
 sg13g2_o21ai_1 _10478_ (.B1(net412),
    .Y(_02894_),
    .A1(net312),
    .A2(_02750_));
 sg13g2_nand2_1 _10479_ (.Y(_02895_),
    .A(net331),
    .B(_02299_));
 sg13g2_buf_1 _10480_ (.A(net312),
    .X(_02896_));
 sg13g2_nand3_1 _10481_ (.B(_02417_),
    .C(net210),
    .A(_02896_),
    .Y(_02897_));
 sg13g2_nand3_1 _10482_ (.B(_02895_),
    .C(_02897_),
    .A(_02894_),
    .Y(_02898_));
 sg13g2_a22oi_1 _10483_ (.Y(_02899_),
    .B1(_02898_),
    .B2(_02373_),
    .A2(_02893_),
    .A1(net311));
 sg13g2_o21ai_1 _10484_ (.B1(_02899_),
    .Y(_02900_),
    .A1(net133),
    .A2(_02891_));
 sg13g2_buf_2 _10485_ (.A(\clock_inst.min_b[1] ),
    .X(_02901_));
 sg13g2_nand2_1 _10486_ (.Y(_02902_),
    .A(_02901_),
    .B(net34));
 sg13g2_o21ai_1 _10487_ (.B1(_02902_),
    .Y(_00236_),
    .A1(net32),
    .A2(_02900_));
 sg13g2_buf_2 _10488_ (.A(\clock_inst.min_b[20] ),
    .X(_02903_));
 sg13g2_o21ai_1 _10489_ (.B1(_02716_),
    .Y(_02904_),
    .A1(net230),
    .A2(_02384_));
 sg13g2_o21ai_1 _10490_ (.B1(_02904_),
    .Y(_02905_),
    .A1(_02362_),
    .A2(_02470_));
 sg13g2_nand2_1 _10491_ (.Y(_02906_),
    .A(net408),
    .B(_02596_));
 sg13g2_a221oi_1 _10492_ (.B2(net310),
    .C1(_02660_),
    .B1(_02906_),
    .A1(_02188_),
    .Y(_02907_),
    .A2(net194));
 sg13g2_nand2_1 _10493_ (.Y(_02908_),
    .A(_02417_),
    .B(net210));
 sg13g2_a221oi_1 _10494_ (.B2(net296),
    .C1(net325),
    .B1(_02908_),
    .A1(net194),
    .Y(_02909_),
    .A2(net298));
 sg13g2_a21oi_1 _10495_ (.A1(net309),
    .A2(_02907_),
    .Y(_02910_),
    .B1(_02909_));
 sg13g2_nor3_1 _10496_ (.A(net70),
    .B(_02905_),
    .C(_02910_),
    .Y(_02911_));
 sg13g2_a21o_1 _10497_ (.A2(net36),
    .A1(_02903_),
    .B1(_02911_),
    .X(_00237_));
 sg13g2_nor2_2 _10498_ (.A(net494),
    .B(net537),
    .Y(_02912_));
 sg13g2_nand2_1 _10499_ (.Y(_02913_),
    .A(_02676_),
    .B(_02912_));
 sg13g2_and2_1 _10500_ (.A(_02587_),
    .B(_02913_),
    .X(_02914_));
 sg13g2_o21ai_1 _10501_ (.B1(_02400_),
    .Y(_02915_),
    .A1(_02595_),
    .A2(_02892_));
 sg13g2_a21oi_1 _10502_ (.A1(net431),
    .A2(_02914_),
    .Y(_02916_),
    .B1(_02915_));
 sg13g2_nand2_1 _10503_ (.Y(_02917_),
    .A(net195),
    .B(_02916_));
 sg13g2_o21ai_1 _10504_ (.B1(_02912_),
    .Y(_02918_),
    .A1(net231),
    .A2(net420));
 sg13g2_a22oi_1 _10505_ (.Y(_02919_),
    .B1(_02726_),
    .B2(net197),
    .A2(net225),
    .A1(net198));
 sg13g2_nand3_1 _10506_ (.B(_02918_),
    .C(_02919_),
    .A(net131),
    .Y(_02920_));
 sg13g2_a221oi_1 _10507_ (.B2(_02920_),
    .C1(_02607_),
    .B1(_02917_),
    .A1(net299),
    .Y(_02921_),
    .A2(net420));
 sg13g2_buf_1 _10508_ (.A(\clock_inst.min_b[21] ),
    .X(_02922_));
 sg13g2_nand2_1 _10509_ (.Y(_02923_),
    .A(_02922_),
    .B(net34));
 sg13g2_o21ai_1 _10510_ (.B1(_02923_),
    .Y(_00238_),
    .A1(net32),
    .A2(_02921_));
 sg13g2_buf_1 _10511_ (.A(\clock_inst.min_b[22] ),
    .X(_02924_));
 sg13g2_inv_1 _10512_ (.Y(_02925_),
    .A(_02924_));
 sg13g2_o21ai_1 _10513_ (.B1(_02315_),
    .Y(_02926_),
    .A1(net341),
    .A2(net343));
 sg13g2_o21ai_1 _10514_ (.B1(_02926_),
    .Y(_02927_),
    .A1(_02575_),
    .A2(net311));
 sg13g2_o21ai_1 _10515_ (.B1(_02310_),
    .Y(_02928_),
    .A1(net410),
    .A2(net304));
 sg13g2_o21ai_1 _10516_ (.B1(net311),
    .Y(_02929_),
    .A1(net344),
    .A2(net298));
 sg13g2_nand2_1 _10517_ (.Y(_02930_),
    .A(net422),
    .B(net333));
 sg13g2_o21ai_1 _10518_ (.B1(_02930_),
    .Y(_02931_),
    .A1(net303),
    .A2(net207));
 sg13g2_o21ai_1 _10519_ (.B1(_02931_),
    .Y(_02932_),
    .A1(net327),
    .A2(_02726_));
 sg13g2_nand3_1 _10520_ (.B(_02929_),
    .C(_02932_),
    .A(net71),
    .Y(_02933_));
 sg13g2_a221oi_1 _10521_ (.B2(net436),
    .C1(_02933_),
    .B1(_02928_),
    .A1(net208),
    .Y(_02934_),
    .A2(_02927_));
 sg13g2_a21oi_1 _10522_ (.A1(_02925_),
    .A2(net39),
    .Y(_00239_),
    .B1(_02934_));
 sg13g2_buf_1 _10523_ (.A(\clock_inst.min_b[23] ),
    .X(_02935_));
 sg13g2_a22oi_1 _10524_ (.Y(_02936_),
    .B1(_02440_),
    .B2(_02268_),
    .A2(net407),
    .A1(_02306_));
 sg13g2_inv_1 _10525_ (.Y(_02937_),
    .A(_02936_));
 sg13g2_a21oi_1 _10526_ (.A1(net331),
    .A2(net197),
    .Y(_02938_),
    .B1(_02454_));
 sg13g2_nand2_1 _10527_ (.Y(_02939_),
    .A(net481),
    .B(_02800_));
 sg13g2_o21ai_1 _10528_ (.B1(_02939_),
    .Y(_02940_),
    .A1(net228),
    .A2(_02938_));
 sg13g2_nor3_1 _10529_ (.A(_02183_),
    .B(net417),
    .C(net333),
    .Y(_02941_));
 sg13g2_a221oi_1 _10530_ (.B2(net354),
    .C1(_02941_),
    .B1(_02940_),
    .A1(_02517_),
    .Y(_02942_),
    .A2(_02937_));
 sg13g2_mux2_1 _10531_ (.A0(_02935_),
    .A1(_02942_),
    .S(net38),
    .X(_00240_));
 sg13g2_buf_2 _10532_ (.A(\clock_inst.min_b[2] ),
    .X(_02943_));
 sg13g2_inv_1 _10533_ (.Y(_02944_),
    .A(_02943_));
 sg13g2_nor2_1 _10534_ (.A(_02827_),
    .B(_02671_),
    .Y(_02945_));
 sg13g2_o21ai_1 _10535_ (.B1(net219),
    .Y(_02946_),
    .A1(net132),
    .A2(net222));
 sg13g2_nor2_2 _10536_ (.A(net496),
    .B(_02368_),
    .Y(_02947_));
 sg13g2_o21ai_1 _10537_ (.B1(_02585_),
    .Y(_02948_),
    .A1(_02741_),
    .A2(_02947_));
 sg13g2_nand3_1 _10538_ (.B(_02946_),
    .C(_02948_),
    .A(_02801_),
    .Y(_02949_));
 sg13g2_nor2_1 _10539_ (.A(net492),
    .B(net487),
    .Y(_02950_));
 sg13g2_buf_2 _10540_ (.A(_02950_),
    .X(_02951_));
 sg13g2_nand2_1 _10541_ (.Y(_02952_),
    .A(net321),
    .B(_02306_));
 sg13g2_a22oi_1 _10542_ (.Y(_02953_),
    .B1(_02952_),
    .B2(net346),
    .A2(_02602_),
    .A1(_02951_));
 sg13g2_nor2_2 _10543_ (.A(_02282_),
    .B(net478),
    .Y(_02954_));
 sg13g2_o21ai_1 _10544_ (.B1(net228),
    .Y(_02955_),
    .A1(net339),
    .A2(_02954_));
 sg13g2_a21oi_1 _10545_ (.A1(_02953_),
    .A2(_02955_),
    .Y(_02956_),
    .B1(net224));
 sg13g2_a221oi_1 _10546_ (.B2(net205),
    .C1(_02956_),
    .B1(_02949_),
    .A1(_02659_),
    .Y(_02957_),
    .A2(_02376_));
 sg13g2_a22oi_1 _10547_ (.Y(_00241_),
    .B1(_02945_),
    .B2(_02957_),
    .A2(net35),
    .A1(_02944_));
 sg13g2_buf_1 _10548_ (.A(\clock_inst.min_b[24] ),
    .X(_02958_));
 sg13g2_inv_2 _10549_ (.Y(_02959_),
    .A(net566));
 sg13g2_a22oi_1 _10550_ (.Y(_00242_),
    .B1(_02425_),
    .B2(_02290_),
    .A2(net35),
    .A1(_02959_));
 sg13g2_nand2_2 _10551_ (.Y(_02960_),
    .A(net423),
    .B(net487));
 sg13g2_a21oi_1 _10552_ (.A1(_02168_),
    .A2(_02960_),
    .Y(_02961_),
    .B1(net431));
 sg13g2_mux2_1 _10553_ (.A0(_02878_),
    .A1(_02961_),
    .S(net218),
    .X(_02962_));
 sg13g2_nor2_1 _10554_ (.A(net437),
    .B(_02233_),
    .Y(_02963_));
 sg13g2_a21oi_1 _10555_ (.A1(net425),
    .A2(net316),
    .Y(_02964_),
    .B1(_02963_));
 sg13g2_a221oi_1 _10556_ (.B2(_02239_),
    .C1(net325),
    .B1(_02308_),
    .A1(_02516_),
    .Y(_02965_),
    .A2(_02756_));
 sg13g2_a21oi_1 _10557_ (.A1(net309),
    .A2(_02964_),
    .Y(_02966_),
    .B1(_02965_));
 sg13g2_a22oi_1 _10558_ (.Y(_02967_),
    .B1(_02966_),
    .B2(net202),
    .A2(_02962_),
    .A1(net205));
 sg13g2_buf_1 _10559_ (.A(\clock_inst.min_b[36] ),
    .X(_02968_));
 sg13g2_nand2_1 _10560_ (.Y(_02969_),
    .A(_02968_),
    .B(net34));
 sg13g2_o21ai_1 _10561_ (.B1(_02969_),
    .Y(_00243_),
    .A1(net32),
    .A2(_02967_));
 sg13g2_buf_1 _10562_ (.A(\clock_inst.min_b[37] ),
    .X(_02970_));
 sg13g2_buf_1 _10563_ (.A(_02246_),
    .X(_02971_));
 sg13g2_a21oi_1 _10564_ (.A1(_02528_),
    .A2(_02744_),
    .Y(_02972_),
    .B1(net418));
 sg13g2_a221oi_1 _10565_ (.B2(_02707_),
    .C1(_02972_),
    .B1(_02635_),
    .A1(net308),
    .Y(_02973_),
    .A2(_02269_));
 sg13g2_a22oi_1 _10566_ (.Y(_02974_),
    .B1(_02941_),
    .B2(net314),
    .A2(_02817_),
    .A1(_02287_));
 sg13g2_o21ai_1 _10567_ (.B1(_02974_),
    .Y(_02975_),
    .A1(net326),
    .A2(_02973_));
 sg13g2_nor2_1 _10568_ (.A(net482),
    .B(_02224_),
    .Y(_02976_));
 sg13g2_a21oi_1 _10569_ (.A1(net426),
    .A2(_02791_),
    .Y(_02977_),
    .B1(net429));
 sg13g2_a21o_1 _10570_ (.A2(net210),
    .A1(net198),
    .B1(_02977_),
    .X(_02978_));
 sg13g2_a22oi_1 _10571_ (.Y(_02979_),
    .B1(_02978_),
    .B2(net344),
    .A2(_02960_),
    .A1(_02976_));
 sg13g2_nor2_1 _10572_ (.A(net128),
    .B(_02979_),
    .Y(_02980_));
 sg13g2_nor3_1 _10573_ (.A(net73),
    .B(_02975_),
    .C(_02980_),
    .Y(_02981_));
 sg13g2_a21o_1 _10574_ (.A2(net31),
    .A1(_02970_),
    .B1(_02981_),
    .X(_00244_));
 sg13g2_buf_1 _10575_ (.A(\clock_inst.min_b[38] ),
    .X(_02982_));
 sg13g2_inv_1 _10576_ (.Y(_02983_),
    .A(_02982_));
 sg13g2_nor2_1 _10577_ (.A(_02180_),
    .B(_02791_),
    .Y(_02984_));
 sg13g2_a21oi_1 _10578_ (.A1(_02828_),
    .A2(_02856_),
    .Y(_02985_),
    .B1(_02470_));
 sg13g2_nor2_1 _10579_ (.A(_02306_),
    .B(net478),
    .Y(_02986_));
 sg13g2_o21ai_1 _10580_ (.B1(net336),
    .Y(_02987_),
    .A1(_02751_),
    .A2(_02986_));
 sg13g2_a21oi_1 _10581_ (.A1(_02230_),
    .A2(_02987_),
    .Y(_02988_),
    .B1(_02185_));
 sg13g2_o21ai_1 _10582_ (.B1(_02801_),
    .Y(_02989_),
    .A1(net408),
    .A2(net300));
 sg13g2_nand3_1 _10583_ (.B(net348),
    .C(net313),
    .A(net435),
    .Y(_02990_));
 sg13g2_o21ai_1 _10584_ (.B1(net488),
    .Y(_02991_),
    .A1(net351),
    .A2(_02507_));
 sg13g2_nand3_1 _10585_ (.B(_02990_),
    .C(_02991_),
    .A(net303),
    .Y(_02992_));
 sg13g2_o21ai_1 _10586_ (.B1(_02992_),
    .Y(_02993_),
    .A1(net334),
    .A2(_02989_));
 sg13g2_a21oi_1 _10587_ (.A1(_02669_),
    .A2(_02993_),
    .Y(_02994_),
    .B1(net224));
 sg13g2_nor4_1 _10588_ (.A(_02984_),
    .B(_02985_),
    .C(_02988_),
    .D(_02994_),
    .Y(_02995_));
 sg13g2_a22oi_1 _10589_ (.Y(_00245_),
    .B1(_02799_),
    .B2(_02995_),
    .A2(net35),
    .A1(_02983_));
 sg13g2_nor2_1 _10590_ (.A(net488),
    .B(_02200_),
    .Y(_02996_));
 sg13g2_nand2_1 _10591_ (.Y(_02997_),
    .A(_02198_),
    .B(_02378_));
 sg13g2_nor2_2 _10592_ (.A(_02336_),
    .B(_02326_),
    .Y(_02998_));
 sg13g2_nand2_1 _10593_ (.Y(_02999_),
    .A(net298),
    .B(_02998_));
 sg13g2_nand3_1 _10594_ (.B(_02997_),
    .C(_02999_),
    .A(_02585_),
    .Y(_03000_));
 sg13g2_nand3_1 _10595_ (.B(net316),
    .C(_02669_),
    .A(net325),
    .Y(_03001_));
 sg13g2_a22oi_1 _10596_ (.Y(_03002_),
    .B1(_03000_),
    .B2(_03001_),
    .A2(_02996_),
    .A1(net195));
 sg13g2_nor2_2 _10597_ (.A(_02186_),
    .B(_02224_),
    .Y(_03003_));
 sg13g2_a221oi_1 _10598_ (.B2(net341),
    .C1(net352),
    .B1(net420),
    .A1(net497),
    .Y(_03004_),
    .A2(net207));
 sg13g2_o21ai_1 _10599_ (.B1(net198),
    .Y(_03005_),
    .A1(net320),
    .A2(net211));
 sg13g2_nor2_1 _10600_ (.A(net308),
    .B(_02607_),
    .Y(_03006_));
 sg13g2_a22oi_1 _10601_ (.Y(_03007_),
    .B1(_03005_),
    .B2(_03006_),
    .A2(_03004_),
    .A1(net219));
 sg13g2_a22oi_1 _10602_ (.Y(_03008_),
    .B1(_03007_),
    .B2(net224),
    .A2(_03003_),
    .A1(net132));
 sg13g2_o21ai_1 _10603_ (.B1(_03008_),
    .Y(_03009_),
    .A1(net205),
    .A2(_03002_));
 sg13g2_buf_1 _10604_ (.A(\clock_inst.min_b[39] ),
    .X(_03010_));
 sg13g2_nand2_1 _10605_ (.Y(_03011_),
    .A(_03010_),
    .B(net34));
 sg13g2_o21ai_1 _10606_ (.B1(_03011_),
    .Y(_00246_),
    .A1(net32),
    .A2(_03009_));
 sg13g2_buf_1 _10607_ (.A(\clock_inst.min_b[3] ),
    .X(_03012_));
 sg13g2_o21ai_1 _10608_ (.B1(net428),
    .Y(_03013_),
    .A1(net211),
    .A2(_02947_));
 sg13g2_o21ai_1 _10609_ (.B1(_03013_),
    .Y(_03014_),
    .A1(_02255_),
    .A2(net221));
 sg13g2_a22oi_1 _10610_ (.Y(_03015_),
    .B1(_03014_),
    .B2(net212),
    .A2(_02301_),
    .A1(net299));
 sg13g2_a21oi_1 _10611_ (.A1(net350),
    .A2(_02720_),
    .Y(_03016_),
    .B1(_02673_));
 sg13g2_nand2_1 _10612_ (.Y(_03017_),
    .A(net408),
    .B(_02685_));
 sg13g2_a21oi_1 _10613_ (.A1(net322),
    .A2(_03017_),
    .Y(_03018_),
    .B1(_02489_));
 sg13g2_o21ai_1 _10614_ (.B1(_03018_),
    .Y(_03019_),
    .A1(net347),
    .A2(_03016_));
 sg13g2_o21ai_1 _10615_ (.B1(_02504_),
    .Y(_03020_),
    .A1(net316),
    .A2(_02255_));
 sg13g2_a22oi_1 _10616_ (.Y(_03021_),
    .B1(_03020_),
    .B2(net338),
    .A2(_03019_),
    .A1(net215));
 sg13g2_o21ai_1 _10617_ (.B1(_03021_),
    .Y(_03022_),
    .A1(net217),
    .A2(_03015_));
 sg13g2_buf_1 _10618_ (.A(_02350_),
    .X(_03023_));
 sg13g2_mux2_1 _10619_ (.A0(_03012_),
    .A1(_03022_),
    .S(net30),
    .X(_00247_));
 sg13g2_buf_1 _10620_ (.A(\clock_inst.min_b[40] ),
    .X(_03024_));
 sg13g2_inv_1 _10621_ (.Y(_03025_),
    .A(_03024_));
 sg13g2_nor2_1 _10622_ (.A(net494),
    .B(_02229_),
    .Y(_03026_));
 sg13g2_nor2_1 _10623_ (.A(_02378_),
    .B(_03026_),
    .Y(_03027_));
 sg13g2_nand3_1 _10624_ (.B(net413),
    .C(net485),
    .A(net322),
    .Y(_03028_));
 sg13g2_o21ai_1 _10625_ (.B1(_03028_),
    .Y(_03029_),
    .A1(net203),
    .A2(_03027_));
 sg13g2_a22oi_1 _10626_ (.Y(_03030_),
    .B1(_03029_),
    .B2(net134),
    .A2(_02729_),
    .A1(net129));
 sg13g2_o21ai_1 _10627_ (.B1(net432),
    .Y(_03031_),
    .A1(net312),
    .A2(net220));
 sg13g2_nand3_1 _10628_ (.B(_02689_),
    .C(_03031_),
    .A(net203),
    .Y(_03032_));
 sg13g2_buf_1 _10629_ (.A(_02800_),
    .X(_03033_));
 sg13g2_nand3_1 _10630_ (.B(_02274_),
    .C(net295),
    .A(net432),
    .Y(_03034_));
 sg13g2_nand3_1 _10631_ (.B(_02527_),
    .C(_03034_),
    .A(net325),
    .Y(_03035_));
 sg13g2_a21oi_1 _10632_ (.A1(_03032_),
    .A2(_03035_),
    .Y(_03036_),
    .B1(net128));
 sg13g2_a21o_1 _10633_ (.A2(_03030_),
    .A1(net128),
    .B1(_03036_),
    .X(_03037_));
 sg13g2_a22oi_1 _10634_ (.Y(_00248_),
    .B1(_02681_),
    .B2(_03037_),
    .A2(net41),
    .A1(_03025_));
 sg13g2_buf_2 _10635_ (.A(\clock_inst.min_b[41] ),
    .X(_03038_));
 sg13g2_o21ai_1 _10636_ (.B1(net348),
    .Y(_03039_),
    .A1(_02354_),
    .A2(net220));
 sg13g2_o21ai_1 _10637_ (.B1(net428),
    .Y(_03040_),
    .A1(_02378_),
    .A2(_02530_));
 sg13g2_nand2_1 _10638_ (.Y(_03041_),
    .A(_03039_),
    .B(_03040_));
 sg13g2_a21oi_1 _10639_ (.A1(net198),
    .A2(net321),
    .Y(_03042_),
    .B1(_02741_));
 sg13g2_nand2_1 _10640_ (.Y(_03043_),
    .A(net219),
    .B(_03042_));
 sg13g2_o21ai_1 _10641_ (.B1(_03043_),
    .Y(_03044_),
    .A1(net195),
    .A2(_03041_));
 sg13g2_nand2_1 _10642_ (.Y(_03045_),
    .A(net216),
    .B(_02685_));
 sg13g2_nand2_1 _10643_ (.Y(_03046_),
    .A(net207),
    .B(_02310_));
 sg13g2_a22oi_1 _10644_ (.Y(_03047_),
    .B1(_03046_),
    .B2(net308),
    .A2(_02439_),
    .A1(net436));
 sg13g2_nor2_1 _10645_ (.A(net480),
    .B(_02297_),
    .Y(_03048_));
 sg13g2_o21ai_1 _10646_ (.B1(_03003_),
    .Y(_03049_),
    .A1(_03048_),
    .A2(_02513_));
 sg13g2_nand2_1 _10647_ (.Y(_03050_),
    .A(_03047_),
    .B(_03049_));
 sg13g2_a22oi_1 _10648_ (.Y(_03051_),
    .B1(_03050_),
    .B2(net338),
    .A2(_03045_),
    .A1(net436));
 sg13g2_o21ai_1 _10649_ (.B1(_03051_),
    .Y(_03052_),
    .A1(net217),
    .A2(_03044_));
 sg13g2_mux2_1 _10650_ (.A0(_03038_),
    .A1(_03052_),
    .S(net30),
    .X(_00249_));
 sg13g2_buf_1 _10651_ (.A(\clock_inst.min_b[42] ),
    .X(_03053_));
 sg13g2_inv_1 _10652_ (.Y(_03054_),
    .A(_03053_));
 sg13g2_a21oi_1 _10653_ (.A1(net489),
    .A2(_02306_),
    .Y(_03055_),
    .B1(_02648_));
 sg13g2_o21ai_1 _10654_ (.B1(_02997_),
    .Y(_03056_),
    .A1(net320),
    .A2(_03055_));
 sg13g2_a21oi_1 _10655_ (.A1(_02409_),
    .A2(_02657_),
    .Y(_03057_),
    .B1(net427));
 sg13g2_a22oi_1 _10656_ (.Y(_03058_),
    .B1(_03057_),
    .B2(_02403_),
    .A2(_03056_),
    .A1(net344));
 sg13g2_nand2_1 _10657_ (.Y(_03059_),
    .A(net354),
    .B(_03058_));
 sg13g2_a21oi_1 _10658_ (.A1(_02232_),
    .A2(net408),
    .Y(_03060_),
    .B1(net418));
 sg13g2_o21ai_1 _10659_ (.B1(net213),
    .Y(_03061_),
    .A1(_02951_),
    .A2(_03060_));
 sg13g2_nor2_2 _10660_ (.A(_02197_),
    .B(_02180_),
    .Y(_03062_));
 sg13g2_a21oi_1 _10661_ (.A1(_02659_),
    .A2(_02818_),
    .Y(_03063_),
    .B1(_03062_));
 sg13g2_nand3_1 _10662_ (.B(_03061_),
    .C(_03063_),
    .A(_02747_),
    .Y(_03064_));
 sg13g2_a221oi_1 _10663_ (.B2(_03064_),
    .C1(net70),
    .B1(_03059_),
    .A1(net299),
    .Y(_03065_),
    .A2(_02659_));
 sg13g2_a21oi_1 _10664_ (.A1(_03054_),
    .A2(net39),
    .Y(_00250_),
    .B1(_03065_));
 sg13g2_buf_1 _10665_ (.A(\clock_inst.min_b[43] ),
    .X(_03066_));
 sg13g2_inv_1 _10666_ (.Y(_03067_),
    .A(_03066_));
 sg13g2_nor2_2 _10667_ (.A(net491),
    .B(net537),
    .Y(_03068_));
 sg13g2_a21oi_1 _10668_ (.A1(net424),
    .A2(_02547_),
    .Y(_03069_),
    .B1(_03068_));
 sg13g2_o21ai_1 _10669_ (.B1(net345),
    .Y(_03070_),
    .A1(_02340_),
    .A2(_03069_));
 sg13g2_and2_1 _10670_ (.A(_02747_),
    .B(_03070_),
    .X(_03071_));
 sg13g2_nand2_1 _10671_ (.Y(_03072_),
    .A(_02418_),
    .B(net304));
 sg13g2_a21oi_1 _10672_ (.A1(_02881_),
    .A2(_03072_),
    .Y(_03073_),
    .B1(_02219_));
 sg13g2_a221oi_1 _10673_ (.B2(_02481_),
    .C1(_03073_),
    .B1(_02998_),
    .A1(_02642_),
    .Y(_03074_),
    .A2(net221));
 sg13g2_a21oi_1 _10674_ (.A1(net227),
    .A2(_03057_),
    .Y(_03075_),
    .B1(_02986_));
 sg13g2_o21ai_1 _10675_ (.B1(_03075_),
    .Y(_03076_),
    .A1(net208),
    .A2(_03074_));
 sg13g2_o21ai_1 _10676_ (.B1(net71),
    .Y(_03077_),
    .A1(_03071_),
    .A2(_03076_));
 sg13g2_o21ai_1 _10677_ (.B1(_03077_),
    .Y(_00251_),
    .A1(_03067_),
    .A2(_02351_));
 sg13g2_buf_1 _10678_ (.A(\clock_inst.min_b[44] ),
    .X(_03078_));
 sg13g2_nand2_2 _10679_ (.Y(_03079_),
    .A(_02167_),
    .B(_03068_));
 sg13g2_o21ai_1 _10680_ (.B1(net306),
    .Y(_03080_),
    .A1(net485),
    .A2(_02750_));
 sg13g2_a21oi_1 _10681_ (.A1(_03079_),
    .A2(_03080_),
    .Y(_03081_),
    .B1(_02535_));
 sg13g2_a21o_1 _10682_ (.A2(net31),
    .A1(_03078_),
    .B1(_03081_),
    .X(_00252_));
 sg13g2_o21ai_1 _10683_ (.B1(net478),
    .Y(_03082_),
    .A1(_02302_),
    .A2(net339));
 sg13g2_inv_1 _10684_ (.Y(_03083_),
    .A(_03082_));
 sg13g2_nand2_1 _10685_ (.Y(_03084_),
    .A(_02756_),
    .B(net478));
 sg13g2_a22oi_1 _10686_ (.Y(_03085_),
    .B1(_03084_),
    .B2(net416),
    .A2(_02819_),
    .A1(net343));
 sg13g2_o21ai_1 _10687_ (.B1(_03085_),
    .Y(_03086_),
    .A1(net228),
    .A2(_03083_));
 sg13g2_a21oi_1 _10688_ (.A1(net353),
    .A2(_02362_),
    .Y(_03087_),
    .B1(_02291_));
 sg13g2_o21ai_1 _10689_ (.B1(_02480_),
    .Y(_03088_),
    .A1(net297),
    .A2(net220));
 sg13g2_o21ai_1 _10690_ (.B1(_03088_),
    .Y(_03089_),
    .A1(net318),
    .A2(_03087_));
 sg13g2_buf_1 _10691_ (.A(_02486_),
    .X(_03090_));
 sg13g2_a21oi_1 _10692_ (.A1(_02213_),
    .A2(_02888_),
    .Y(_03091_),
    .B1(_03048_));
 sg13g2_nor2_1 _10693_ (.A(net199),
    .B(_03091_),
    .Y(_03092_));
 sg13g2_a221oi_1 _10694_ (.B2(net193),
    .C1(_03092_),
    .B1(_03089_),
    .A1(net214),
    .Y(_03093_),
    .A2(_03086_));
 sg13g2_buf_2 _10695_ (.A(\clock_inst.min_b[4] ),
    .X(_03094_));
 sg13g2_nand2_1 _10696_ (.Y(_03095_),
    .A(_03094_),
    .B(net34));
 sg13g2_o21ai_1 _10697_ (.B1(_03095_),
    .Y(_00253_),
    .A1(net32),
    .A2(_03093_));
 sg13g2_nor2_1 _10698_ (.A(_02452_),
    .B(_02513_),
    .Y(_03096_));
 sg13g2_nand3_1 _10699_ (.B(_02306_),
    .C(net216),
    .A(net226),
    .Y(_03097_));
 sg13g2_nor2_1 _10700_ (.A(net496),
    .B(_02433_),
    .Y(_03098_));
 sg13g2_o21ai_1 _10701_ (.B1(net213),
    .Y(_03099_),
    .A1(_02479_),
    .A2(_03098_));
 sg13g2_nand2_1 _10702_ (.Y(_03100_),
    .A(_03097_),
    .B(_03099_));
 sg13g2_o21ai_1 _10703_ (.B1(_02960_),
    .Y(_03101_),
    .A1(net439),
    .A2(_02400_));
 sg13g2_o21ai_1 _10704_ (.B1(net300),
    .Y(_03102_),
    .A1(net198),
    .A2(net321));
 sg13g2_a22oi_1 _10705_ (.Y(_03103_),
    .B1(_03102_),
    .B2(net219),
    .A2(_03101_),
    .A1(net225));
 sg13g2_nor2_1 _10706_ (.A(net301),
    .B(net335),
    .Y(_03104_));
 sg13g2_o21ai_1 _10707_ (.B1(net344),
    .Y(_03105_),
    .A1(_02795_),
    .A2(_03104_));
 sg13g2_a21oi_1 _10708_ (.A1(_03103_),
    .A2(_03105_),
    .Y(_03106_),
    .B1(net338));
 sg13g2_a221oi_1 _10709_ (.B2(net217),
    .C1(_03106_),
    .B1(_03100_),
    .A1(_02951_),
    .Y(_03107_),
    .A2(_03096_));
 sg13g2_buf_2 _10710_ (.A(\clock_inst.min_b[5] ),
    .X(_03108_));
 sg13g2_nand2_1 _10711_ (.Y(_03109_),
    .A(_03108_),
    .B(_02736_));
 sg13g2_o21ai_1 _10712_ (.B1(_03109_),
    .Y(_00254_),
    .A1(net32),
    .A2(_03107_));
 sg13g2_buf_2 _10713_ (.A(\clock_inst.min_b[6] ),
    .X(_03110_));
 sg13g2_a22oi_1 _10714_ (.Y(_03111_),
    .B1(_02440_),
    .B2(_02976_),
    .A2(net304),
    .A1(net425));
 sg13g2_a21oi_1 _10715_ (.A1(net417),
    .A2(_02453_),
    .Y(_03112_),
    .B1(_02417_));
 sg13g2_a21oi_1 _10716_ (.A1(net345),
    .A2(_02892_),
    .Y(_03113_),
    .B1(net421));
 sg13g2_a21oi_1 _10717_ (.A1(_02504_),
    .A2(net300),
    .Y(_03114_),
    .B1(net322));
 sg13g2_nor4_1 _10718_ (.A(net296),
    .B(_03112_),
    .C(_03113_),
    .D(_03114_),
    .Y(_03115_));
 sg13g2_a21oi_1 _10719_ (.A1(net223),
    .A2(_03111_),
    .Y(_03116_),
    .B1(_03115_));
 sg13g2_a21oi_1 _10720_ (.A1(net425),
    .A2(net352),
    .Y(_03117_),
    .B1(_02700_));
 sg13g2_nor2_1 _10721_ (.A(_02431_),
    .B(_02413_),
    .Y(_03118_));
 sg13g2_o21ai_1 _10722_ (.B1(net327),
    .Y(_03119_),
    .A1(_02673_),
    .A2(_03118_));
 sg13g2_o21ai_1 _10723_ (.B1(_03119_),
    .Y(_03120_),
    .A1(net407),
    .A2(_03117_));
 sg13g2_nor3_1 _10724_ (.A(net73),
    .B(_03116_),
    .C(_03120_),
    .Y(_03121_));
 sg13g2_a21o_1 _10725_ (.A2(net31),
    .A1(_03110_),
    .B1(_03121_),
    .X(_00255_));
 sg13g2_buf_1 _10726_ (.A(\clock_inst.min_b[7] ),
    .X(_03122_));
 sg13g2_o21ai_1 _10727_ (.B1(_02677_),
    .Y(_03123_),
    .A1(net415),
    .A2(_02400_));
 sg13g2_o21ai_1 _10728_ (.B1(_02255_),
    .Y(_03124_),
    .A1(net324),
    .A2(net485));
 sg13g2_nor2_1 _10729_ (.A(net324),
    .B(_02633_),
    .Y(_03125_));
 sg13g2_a21oi_1 _10730_ (.A1(net418),
    .A2(_03124_),
    .Y(_03126_),
    .B1(_03125_));
 sg13g2_nor2_1 _10731_ (.A(net416),
    .B(_03126_),
    .Y(_03127_));
 sg13g2_a221oi_1 _10732_ (.B2(_02550_),
    .C1(_03127_),
    .B1(_03123_),
    .A1(_02242_),
    .Y(_03128_),
    .A2(net196));
 sg13g2_a21oi_1 _10733_ (.A1(net350),
    .A2(_02657_),
    .Y(_03129_),
    .B1(_03003_));
 sg13g2_o21ai_1 _10734_ (.B1(net335),
    .Y(_03130_),
    .A1(_02488_),
    .A2(_03129_));
 sg13g2_a21oi_1 _10735_ (.A1(net326),
    .A2(_03130_),
    .Y(_03131_),
    .B1(_02718_));
 sg13g2_o21ai_1 _10736_ (.B1(_03131_),
    .Y(_03132_),
    .A1(net202),
    .A2(_03128_));
 sg13g2_mux2_1 _10737_ (.A0(_03122_),
    .A1(_03132_),
    .S(_03023_),
    .X(_00256_));
 sg13g2_buf_2 _10738_ (.A(\clock_inst.min_b[8] ),
    .X(_03133_));
 sg13g2_a22oi_1 _10739_ (.Y(_03134_),
    .B1(_02769_),
    .B2(net306),
    .A2(_02270_),
    .A1(net230));
 sg13g2_a21oi_1 _10740_ (.A1(net200),
    .A2(_02867_),
    .Y(_03135_),
    .B1(_02756_));
 sg13g2_nor2_1 _10741_ (.A(net72),
    .B(_03135_),
    .Y(_03136_));
 sg13g2_a22oi_1 _10742_ (.Y(_03137_),
    .B1(_03134_),
    .B2(_03136_),
    .A2(net70),
    .A1(_03133_));
 sg13g2_inv_1 _10743_ (.Y(_00257_),
    .A(_03137_));
 sg13g2_inv_1 _10744_ (.Y(_03138_),
    .A(\clock_inst.min_c[0] ));
 sg13g2_o21ai_1 _10745_ (.B1(_02633_),
    .Y(_03139_),
    .A1(_02269_),
    .A2(_02473_));
 sg13g2_o21ai_1 _10746_ (.B1(net422),
    .Y(_03140_),
    .A1(net480),
    .A2(_02378_));
 sg13g2_a22oi_1 _10747_ (.Y(_03141_),
    .B1(_02233_),
    .B2(net486),
    .A2(net352),
    .A1(net419));
 sg13g2_nand3_1 _10748_ (.B(_03140_),
    .C(_03141_),
    .A(net348),
    .Y(_03142_));
 sg13g2_o21ai_1 _10749_ (.B1(_03142_),
    .Y(_03143_),
    .A1(net231),
    .A2(_03139_));
 sg13g2_a21oi_1 _10750_ (.A1(_03079_),
    .A2(_03143_),
    .Y(_03144_),
    .B1(_02371_));
 sg13g2_o21ai_1 _10751_ (.B1(net321),
    .Y(_03145_),
    .A1(_02187_),
    .A2(net330));
 sg13g2_a22oi_1 _10752_ (.Y(_03146_),
    .B1(_03145_),
    .B2(_02576_),
    .A2(_02849_),
    .A1(net308));
 sg13g2_o21ai_1 _10753_ (.B1(_02225_),
    .Y(_03147_),
    .A1(_02222_),
    .A2(_02619_));
 sg13g2_a21o_1 _10754_ (.A2(_03147_),
    .A1(net345),
    .B1(_02412_),
    .X(_03148_));
 sg13g2_o21ai_1 _10755_ (.B1(_03148_),
    .Y(_03149_),
    .A1(net318),
    .A2(_03146_));
 sg13g2_o21ai_1 _10756_ (.B1(net71),
    .Y(_03150_),
    .A1(_03144_),
    .A2(_03149_));
 sg13g2_o21ai_1 _10757_ (.B1(_03150_),
    .Y(_00258_),
    .A1(_03138_),
    .A2(net38));
 sg13g2_nand2_1 _10758_ (.Y(_03151_),
    .A(_02180_),
    .B(_02800_));
 sg13g2_a22oi_1 _10759_ (.Y(_03152_),
    .B1(_03151_),
    .B2(net409),
    .A2(_02976_),
    .A1(net194));
 sg13g2_nor2_1 _10760_ (.A(_02217_),
    .B(net426),
    .Y(_03153_));
 sg13g2_nor3_1 _10761_ (.A(net435),
    .B(_03153_),
    .C(_02912_),
    .Y(_03154_));
 sg13g2_a21oi_1 _10762_ (.A1(net345),
    .A2(_02856_),
    .Y(_03155_),
    .B1(net483));
 sg13g2_o21ai_1 _10763_ (.B1(net296),
    .Y(_03156_),
    .A1(_03154_),
    .A2(_03155_));
 sg13g2_o21ai_1 _10764_ (.B1(_03156_),
    .Y(_03157_),
    .A1(net228),
    .A2(_03152_));
 sg13g2_a21oi_1 _10765_ (.A1(_02791_),
    .A2(net295),
    .Y(_03158_),
    .B1(_02306_));
 sg13g2_a21o_1 _10766_ (.A2(net227),
    .A1(net196),
    .B1(_03158_),
    .X(_03159_));
 sg13g2_o21ai_1 _10767_ (.B1(_02951_),
    .Y(_03160_),
    .A1(net226),
    .A2(_02726_));
 sg13g2_a21oi_1 _10768_ (.A1(_02528_),
    .A2(_03160_),
    .Y(_03161_),
    .B1(net202));
 sg13g2_a221oi_1 _10769_ (.B2(net217),
    .C1(_03161_),
    .B1(_03159_),
    .A1(net130),
    .Y(_03162_),
    .A2(_03157_));
 sg13g2_buf_1 _10770_ (.A(_02246_),
    .X(_03163_));
 sg13g2_nand2_1 _10771_ (.Y(_03164_),
    .A(\clock_inst.min_c[10] ),
    .B(net29));
 sg13g2_o21ai_1 _10772_ (.B1(_03164_),
    .Y(_00259_),
    .A1(net32),
    .A2(_03162_));
 sg13g2_o21ai_1 _10773_ (.B1(_02912_),
    .Y(_03165_),
    .A1(_02265_),
    .A2(net342));
 sg13g2_a21oi_1 _10774_ (.A1(_02740_),
    .A2(_03165_),
    .Y(_03166_),
    .B1(net195));
 sg13g2_nand2_1 _10775_ (.Y(_03167_),
    .A(_02639_),
    .B(net339));
 sg13g2_a21oi_1 _10776_ (.A1(_03079_),
    .A2(_03167_),
    .Y(_03168_),
    .B1(_02432_));
 sg13g2_nor2_1 _10777_ (.A(net481),
    .B(_02311_),
    .Y(_03169_));
 sg13g2_nand2_1 _10778_ (.Y(_03170_),
    .A(_02329_),
    .B(_02280_));
 sg13g2_o21ai_1 _10779_ (.B1(_03170_),
    .Y(_03171_),
    .A1(net329),
    .A2(_03169_));
 sg13g2_a22oi_1 _10780_ (.Y(_03172_),
    .B1(_03171_),
    .B2(net336),
    .A2(net194),
    .A1(net296));
 sg13g2_o21ai_1 _10781_ (.B1(net422),
    .Y(_03173_),
    .A1(_02280_),
    .A2(_02378_));
 sg13g2_nor2_1 _10782_ (.A(net297),
    .B(_02364_),
    .Y(_03174_));
 sg13g2_a22oi_1 _10783_ (.Y(_03175_),
    .B1(_03174_),
    .B2(_02391_),
    .A2(_03173_),
    .A1(_02774_));
 sg13g2_nor2_1 _10784_ (.A(net346),
    .B(_03175_),
    .Y(_03176_));
 sg13g2_a21oi_1 _10785_ (.A1(net309),
    .A2(_03172_),
    .Y(_03177_),
    .B1(_03176_));
 sg13g2_nor4_1 _10786_ (.A(net72),
    .B(_03166_),
    .C(_03168_),
    .D(_03177_),
    .Y(_03178_));
 sg13g2_a21o_1 _10787_ (.A2(net31),
    .A1(\clock_inst.min_c[11] ),
    .B1(_03178_),
    .X(_00260_));
 sg13g2_a21oi_1 _10788_ (.A1(net323),
    .A2(_02707_),
    .Y(_03179_),
    .B1(_02767_));
 sg13g2_nand2_1 _10789_ (.Y(_03180_),
    .A(net343),
    .B(_02954_));
 sg13g2_o21ai_1 _10790_ (.B1(_02391_),
    .Y(_03181_),
    .A1(net339),
    .A2(_03098_));
 sg13g2_nand2_1 _10791_ (.Y(_03182_),
    .A(_03180_),
    .B(_03181_));
 sg13g2_a21oi_1 _10792_ (.A1(_02405_),
    .A2(_02400_),
    .Y(_03183_),
    .B1(_02839_));
 sg13g2_a21oi_1 _10793_ (.A1(_02361_),
    .A2(net210),
    .Y(_03184_),
    .B1(_02584_));
 sg13g2_nand2_1 _10794_ (.Y(_03185_),
    .A(net308),
    .B(_03184_));
 sg13g2_o21ai_1 _10795_ (.B1(_03185_),
    .Y(_03186_),
    .A1(net334),
    .A2(_03183_));
 sg13g2_a22oi_1 _10796_ (.Y(_03187_),
    .B1(_03186_),
    .B2(net134),
    .A2(_03182_),
    .A1(net306));
 sg13g2_o21ai_1 _10797_ (.B1(_03187_),
    .Y(_03188_),
    .A1(net133),
    .A2(_03179_));
 sg13g2_mux2_1 _10798_ (.A0(\clock_inst.min_c[12] ),
    .A1(_03188_),
    .S(net30),
    .X(_00261_));
 sg13g2_a22oi_1 _10799_ (.Y(_03189_),
    .B1(_02875_),
    .B2(_02951_),
    .A2(_02717_),
    .A1(net436));
 sg13g2_o21ai_1 _10800_ (.B1(net350),
    .Y(_03190_),
    .A1(_02530_),
    .A2(_02839_));
 sg13g2_o21ai_1 _10801_ (.B1(_03190_),
    .Y(_03191_),
    .A1(net427),
    .A2(_03189_));
 sg13g2_or2_1 _10802_ (.X(_03192_),
    .B(_03191_),
    .A(_02798_));
 sg13g2_a21o_1 _10803_ (.A2(_02597_),
    .A1(_02439_),
    .B1(net226),
    .X(_03193_));
 sg13g2_o21ai_1 _10804_ (.B1(_02453_),
    .Y(_03194_),
    .A1(net492),
    .A2(_02605_));
 sg13g2_a22oi_1 _10805_ (.Y(_03195_),
    .B1(_03194_),
    .B2(net200),
    .A2(_02720_),
    .A1(net298));
 sg13g2_nor3_1 _10806_ (.A(net421),
    .B(net417),
    .C(net317),
    .Y(_03196_));
 sg13g2_o21ai_1 _10807_ (.B1(net219),
    .Y(_03197_),
    .A1(_02369_),
    .A2(_03196_));
 sg13g2_nand4_1 _10808_ (.B(_03193_),
    .C(_03195_),
    .A(net199),
    .Y(_03198_),
    .D(_03197_));
 sg13g2_o21ai_1 _10809_ (.B1(_03198_),
    .Y(_03199_),
    .A1(net193),
    .A2(_03192_));
 sg13g2_nand2_1 _10810_ (.Y(_03200_),
    .A(\clock_inst.min_c[13] ),
    .B(_03163_));
 sg13g2_o21ai_1 _10811_ (.B1(_03200_),
    .Y(_00262_),
    .A1(_02871_),
    .A2(_03199_));
 sg13g2_inv_1 _10812_ (.Y(_03201_),
    .A(\clock_inst.min_c[14] ));
 sg13g2_nor2_1 _10813_ (.A(_02291_),
    .B(_02492_),
    .Y(_03202_));
 sg13g2_o21ai_1 _10814_ (.B1(_02388_),
    .Y(_03203_),
    .A1(net409),
    .A2(_03202_));
 sg13g2_a22oi_1 _10815_ (.Y(_03204_),
    .B1(_03203_),
    .B2(net129),
    .A2(_02726_),
    .A1(_02181_));
 sg13g2_o21ai_1 _10816_ (.B1(_02769_),
    .Y(_03205_),
    .A1(_02481_),
    .A2(net207));
 sg13g2_a221oi_1 _10817_ (.B2(_02486_),
    .C1(net223),
    .B1(_03205_),
    .A1(net229),
    .Y(_03206_),
    .A2(net299));
 sg13g2_a21o_1 _10818_ (.A2(_03204_),
    .A1(net133),
    .B1(_03206_),
    .X(_03207_));
 sg13g2_a21oi_1 _10819_ (.A1(_02416_),
    .A2(_02281_),
    .Y(_03208_),
    .B1(_02741_));
 sg13g2_a21oi_1 _10820_ (.A1(_02312_),
    .A2(_02677_),
    .Y(_03209_),
    .B1(net341));
 sg13g2_nor3_1 _10821_ (.A(net219),
    .B(_02518_),
    .C(_03209_),
    .Y(_03210_));
 sg13g2_a21oi_1 _10822_ (.A1(net223),
    .A2(_03208_),
    .Y(_03211_),
    .B1(_03210_));
 sg13g2_nor3_1 _10823_ (.A(_02294_),
    .B(_02301_),
    .C(_02417_),
    .Y(_03212_));
 sg13g2_a21oi_1 _10824_ (.A1(net343),
    .A2(_02374_),
    .Y(_03213_),
    .B1(_03212_));
 sg13g2_o21ai_1 _10825_ (.B1(_02425_),
    .Y(_03214_),
    .A1(net345),
    .A2(_03213_));
 sg13g2_a21oi_1 _10826_ (.A1(_02544_),
    .A2(_03211_),
    .Y(_03215_),
    .B1(_03214_));
 sg13g2_a22oi_1 _10827_ (.Y(_00263_),
    .B1(_03207_),
    .B2(_03215_),
    .A2(net41),
    .A1(_03201_));
 sg13g2_o21ai_1 _10828_ (.B1(net228),
    .Y(_03216_),
    .A1(net420),
    .A2(_02795_));
 sg13g2_nand2b_1 _10829_ (.Y(_03217_),
    .B(_03216_),
    .A_N(_02963_));
 sg13g2_a221oi_1 _10830_ (.B2(net347),
    .C1(net196),
    .B1(_02875_),
    .A1(_02746_),
    .Y(_03218_),
    .A2(net220));
 sg13g2_o21ai_1 _10831_ (.B1(_02670_),
    .Y(_03219_),
    .A1(net340),
    .A2(net207));
 sg13g2_o21ai_1 _10832_ (.B1(_02791_),
    .Y(_03220_),
    .A1(net432),
    .A2(net204));
 sg13g2_a22oi_1 _10833_ (.Y(_03221_),
    .B1(_03220_),
    .B2(net131),
    .A2(_03219_),
    .A1(net328));
 sg13g2_o21ai_1 _10834_ (.B1(_03221_),
    .Y(_03222_),
    .A1(net326),
    .A2(_03218_));
 sg13g2_a21oi_1 _10835_ (.A1(net202),
    .A2(_03217_),
    .Y(_03223_),
    .B1(_03222_));
 sg13g2_nand2_1 _10836_ (.Y(_03224_),
    .A(\clock_inst.min_c[15] ),
    .B(_03163_));
 sg13g2_o21ai_1 _10837_ (.B1(_03224_),
    .Y(_00264_),
    .A1(net32),
    .A2(_03223_));
 sg13g2_buf_1 _10838_ (.A(_02171_),
    .X(_03225_));
 sg13g2_o21ai_1 _10839_ (.B1(net315),
    .Y(_03226_),
    .A1(net218),
    .A2(_02527_));
 sg13g2_a21oi_1 _10840_ (.A1(net353),
    .A2(_02707_),
    .Y(_03227_),
    .B1(net227));
 sg13g2_o21ai_1 _10841_ (.B1(_02184_),
    .Y(_03228_),
    .A1(_02228_),
    .A2(_02480_));
 sg13g2_o21ai_1 _10842_ (.B1(_03228_),
    .Y(_03229_),
    .A1(net314),
    .A2(_03227_));
 sg13g2_o21ai_1 _10843_ (.B1(_02539_),
    .Y(_03230_),
    .A1(net408),
    .A2(_02633_));
 sg13g2_a221oi_1 _10844_ (.B2(net208),
    .C1(_03230_),
    .B1(_03229_),
    .A1(net354),
    .Y(_03231_),
    .A2(_03226_));
 sg13g2_nand2_1 _10845_ (.Y(_03232_),
    .A(\clock_inst.min_c[16] ),
    .B(net29));
 sg13g2_o21ai_1 _10846_ (.B1(_03232_),
    .Y(_00265_),
    .A1(net28),
    .A2(_03231_));
 sg13g2_a21oi_1 _10847_ (.A1(_02523_),
    .A2(_02465_),
    .Y(_03233_),
    .B1(_02201_));
 sg13g2_o21ai_1 _10848_ (.B1(net408),
    .Y(_03234_),
    .A1(net410),
    .A2(net295));
 sg13g2_a221oi_1 _10849_ (.B2(net346),
    .C1(_02716_),
    .B1(_03234_),
    .A1(net213),
    .Y(_03235_),
    .A2(net194));
 sg13g2_o21ai_1 _10850_ (.B1(_03235_),
    .Y(_03236_),
    .A1(net214),
    .A2(_03233_));
 sg13g2_nand2_1 _10851_ (.Y(_03237_),
    .A(\clock_inst.min_c[17] ),
    .B(net29));
 sg13g2_o21ai_1 _10852_ (.B1(_03237_),
    .Y(_00266_),
    .A1(net28),
    .A2(_03236_));
 sg13g2_o21ai_1 _10853_ (.B1(_02619_),
    .Y(_03238_),
    .A1(net440),
    .A2(_02740_));
 sg13g2_o21ai_1 _10854_ (.B1(net305),
    .Y(_03239_),
    .A1(net426),
    .A2(_02561_));
 sg13g2_nand4_1 _10855_ (.B(_02234_),
    .C(_03033_),
    .A(_02833_),
    .Y(_03240_),
    .D(_03239_));
 sg13g2_nand2_1 _10856_ (.Y(_03241_),
    .A(_02469_),
    .B(_03167_));
 sg13g2_a22oi_1 _10857_ (.Y(_03242_),
    .B1(_03241_),
    .B2(net309),
    .A2(_03240_),
    .A1(_03238_));
 sg13g2_o21ai_1 _10858_ (.B1(net302),
    .Y(_03243_),
    .A1(net407),
    .A2(_02573_));
 sg13g2_a21o_1 _10859_ (.A2(_02312_),
    .A1(net206),
    .B1(_02277_),
    .X(_03244_));
 sg13g2_nor2_2 _10860_ (.A(_02211_),
    .B(net204),
    .Y(_03245_));
 sg13g2_o21ai_1 _10861_ (.B1(_02608_),
    .Y(_03246_),
    .A1(net211),
    .A2(_03245_));
 sg13g2_nand3_1 _10862_ (.B(_03244_),
    .C(_03246_),
    .A(_03243_),
    .Y(_03247_));
 sg13g2_a22oi_1 _10863_ (.Y(_03248_),
    .B1(_03247_),
    .B2(net193),
    .A2(net194),
    .A1(net131));
 sg13g2_o21ai_1 _10864_ (.B1(_03248_),
    .Y(_03249_),
    .A1(_03090_),
    .A2(_03242_));
 sg13g2_nand2_1 _10865_ (.Y(_03250_),
    .A(\clock_inst.min_c[19] ),
    .B(net29));
 sg13g2_o21ai_1 _10866_ (.B1(_03250_),
    .Y(_00267_),
    .A1(net28),
    .A2(_03249_));
 sg13g2_nand2_1 _10867_ (.Y(_03251_),
    .A(_02230_),
    .B(net330));
 sg13g2_a21oi_1 _10868_ (.A1(net422),
    .A2(_02960_),
    .Y(_03252_),
    .B1(net311));
 sg13g2_o21ai_1 _10869_ (.B1(_02588_),
    .Y(_03253_),
    .A1(net351),
    .A2(_03252_));
 sg13g2_nand2_1 _10870_ (.Y(_03254_),
    .A(net231),
    .B(_03253_));
 sg13g2_o21ai_1 _10871_ (.B1(_03254_),
    .Y(_03255_),
    .A1(_02669_),
    .A2(_02255_));
 sg13g2_a21oi_1 _10872_ (.A1(_02253_),
    .A2(_02450_),
    .Y(_03256_),
    .B1(net421));
 sg13g2_nor3_1 _10873_ (.A(net296),
    .B(_02795_),
    .C(_03256_),
    .Y(_03257_));
 sg13g2_a221oi_1 _10874_ (.B2(net412),
    .C1(net218),
    .B1(net196),
    .A1(net310),
    .Y(_03258_),
    .A2(net211));
 sg13g2_nor3_1 _10875_ (.A(net199),
    .B(_03257_),
    .C(_03258_),
    .Y(_03259_));
 sg13g2_a221oi_1 _10876_ (.B2(net193),
    .C1(_03259_),
    .B1(_03255_),
    .A1(net304),
    .Y(_03260_),
    .A2(_03251_));
 sg13g2_nand2_1 _10877_ (.Y(_03261_),
    .A(\clock_inst.min_c[1] ),
    .B(net29));
 sg13g2_o21ai_1 _10878_ (.B1(_03261_),
    .Y(_00268_),
    .A1(net28),
    .A2(_03260_));
 sg13g2_inv_1 _10879_ (.Y(_03262_),
    .A(\clock_inst.min_c[21] ));
 sg13g2_a22oi_1 _10880_ (.Y(_03263_),
    .B1(_02380_),
    .B2(net197),
    .A2(_02513_),
    .A1(_02175_));
 sg13g2_nor2_2 _10881_ (.A(net307),
    .B(_02363_),
    .Y(_03264_));
 sg13g2_nand3_1 _10882_ (.B(_02507_),
    .C(_03264_),
    .A(net319),
    .Y(_03265_));
 sg13g2_o21ai_1 _10883_ (.B1(_03265_),
    .Y(_03266_),
    .A1(net200),
    .A2(_03263_));
 sg13g2_a21oi_1 _10884_ (.A1(net351),
    .A2(_02817_),
    .Y(_03267_),
    .B1(net490));
 sg13g2_a21o_1 _10885_ (.A2(_03151_),
    .A1(net429),
    .B1(_03267_),
    .X(_03268_));
 sg13g2_a21oi_1 _10886_ (.A1(net489),
    .A2(_02387_),
    .Y(_03269_),
    .B1(_02750_));
 sg13g2_a22oi_1 _10887_ (.Y(_03270_),
    .B1(_03269_),
    .B2(net222),
    .A2(_03268_),
    .A1(net203));
 sg13g2_a21oi_1 _10888_ (.A1(_02240_),
    .A2(_02939_),
    .Y(_03271_),
    .B1(_02532_));
 sg13g2_nor2_1 _10889_ (.A(net432),
    .B(_03271_),
    .Y(_03272_));
 sg13g2_nor2_1 _10890_ (.A(_02580_),
    .B(net210),
    .Y(_03273_));
 sg13g2_o21ai_1 _10891_ (.B1(net483),
    .Y(_03274_),
    .A1(_02215_),
    .A2(net307));
 sg13g2_a21oi_1 _10892_ (.A1(_02939_),
    .A2(_03274_),
    .Y(_03275_),
    .B1(net412));
 sg13g2_nor4_1 _10893_ (.A(net218),
    .B(_03272_),
    .C(_03273_),
    .D(_03275_),
    .Y(_03276_));
 sg13g2_a21oi_1 _10894_ (.A1(net128),
    .A2(_03270_),
    .Y(_03277_),
    .B1(_03276_));
 sg13g2_nor3_1 _10895_ (.A(net70),
    .B(_03266_),
    .C(_03277_),
    .Y(_03278_));
 sg13g2_a21oi_1 _10896_ (.A1(_03262_),
    .A2(net39),
    .Y(_00269_),
    .B1(_03278_));
 sg13g2_nor2b_1 _10897_ (.A(_02331_),
    .B_N(_02450_),
    .Y(_03279_));
 sg13g2_nor3_1 _10898_ (.A(net350),
    .B(net307),
    .C(net332),
    .Y(_03280_));
 sg13g2_a21oi_1 _10899_ (.A1(net296),
    .A2(_03279_),
    .Y(_03281_),
    .B1(_03280_));
 sg13g2_nand3b_1 _10900_ (.B(net440),
    .C(net295),
    .Y(_03282_),
    .A_N(_03062_));
 sg13g2_o21ai_1 _10901_ (.B1(_03282_),
    .Y(_03283_),
    .A1(net318),
    .A2(_03281_));
 sg13g2_a21oi_1 _10902_ (.A1(_02353_),
    .A2(_02487_),
    .Y(_03284_),
    .B1(_02401_));
 sg13g2_a221oi_1 _10903_ (.B2(net324),
    .C1(_03284_),
    .B1(_02707_),
    .A1(net486),
    .Y(_03285_),
    .A2(net297));
 sg13g2_a21oi_1 _10904_ (.A1(_02633_),
    .A2(net313),
    .Y(_03286_),
    .B1(_02209_));
 sg13g2_nor3_1 _10905_ (.A(net427),
    .B(_02518_),
    .C(_03286_),
    .Y(_03287_));
 sg13g2_a21oi_1 _10906_ (.A1(net431),
    .A2(_03285_),
    .Y(_03288_),
    .B1(_03287_));
 sg13g2_nor2_1 _10907_ (.A(net410),
    .B(_02881_),
    .Y(_03289_));
 sg13g2_o21ai_1 _10908_ (.B1(net302),
    .Y(_03290_),
    .A1(_02489_),
    .A2(_03289_));
 sg13g2_inv_1 _10909_ (.Y(_03291_),
    .A(_03290_));
 sg13g2_a221oi_1 _10910_ (.B2(net323),
    .C1(_03291_),
    .B1(_03288_),
    .A1(net196),
    .Y(_03292_),
    .A2(_02717_));
 sg13g2_o21ai_1 _10911_ (.B1(_03292_),
    .Y(_03293_),
    .A1(net217),
    .A2(_03283_));
 sg13g2_mux2_1 _10912_ (.A0(\clock_inst.min_c[22] ),
    .A1(_03293_),
    .S(net30),
    .X(_00270_));
 sg13g2_inv_1 _10913_ (.Y(_03294_),
    .A(\clock_inst.min_c[23] ));
 sg13g2_o21ai_1 _10914_ (.B1(_02312_),
    .Y(_03295_),
    .A1(net490),
    .A2(_02540_));
 sg13g2_o21ai_1 _10915_ (.B1(net336),
    .Y(_03296_),
    .A1(net225),
    .A2(_03295_));
 sg13g2_nand3_1 _10916_ (.B(_02504_),
    .C(_03296_),
    .A(net131),
    .Y(_03297_));
 sg13g2_nand2_1 _10917_ (.Y(_03298_),
    .A(_02322_),
    .B(net196));
 sg13g2_nand3_1 _10918_ (.B(_02832_),
    .C(_03298_),
    .A(net195),
    .Y(_03299_));
 sg13g2_nor2_1 _10919_ (.A(_02405_),
    .B(net295),
    .Y(_03300_));
 sg13g2_a22oi_1 _10920_ (.Y(_03301_),
    .B1(_03300_),
    .B2(net200),
    .A2(_03264_),
    .A1(net409));
 sg13g2_nand3_1 _10921_ (.B(_02579_),
    .C(_03153_),
    .A(net344),
    .Y(_03302_));
 sg13g2_o21ai_1 _10922_ (.B1(_03302_),
    .Y(_03303_),
    .A1(net131),
    .A2(_03301_));
 sg13g2_a221oi_1 _10923_ (.B2(net130),
    .C1(_02827_),
    .B1(_03303_),
    .A1(_03297_),
    .Y(_03304_),
    .A2(_03299_));
 sg13g2_a21oi_1 _10924_ (.A1(_03294_),
    .A2(_02251_),
    .Y(_00271_),
    .B1(_03304_));
 sg13g2_o21ai_1 _10925_ (.B1(net303),
    .Y(_03305_),
    .A1(net222),
    .A2(_02954_));
 sg13g2_nand2_1 _10926_ (.Y(_03306_),
    .A(_02312_),
    .B(_03305_));
 sg13g2_a22oi_1 _10927_ (.Y(_03307_),
    .B1(_03306_),
    .B2(net327),
    .A2(_02518_),
    .A1(_02546_));
 sg13g2_nor2_1 _10928_ (.A(net482),
    .B(net433),
    .Y(_03308_));
 sg13g2_a21oi_1 _10929_ (.A1(_02353_),
    .A2(net330),
    .Y(_03309_),
    .B1(net418));
 sg13g2_or2_1 _10930_ (.X(_03310_),
    .B(_03309_),
    .A(_02532_));
 sg13g2_a22oi_1 _10931_ (.Y(_03311_),
    .B1(_03310_),
    .B2(net128),
    .A2(_03308_),
    .A1(_02529_));
 sg13g2_o21ai_1 _10932_ (.B1(_03311_),
    .Y(_03312_),
    .A1(net193),
    .A2(_03307_));
 sg13g2_mux2_1 _10933_ (.A0(\clock_inst.min_c[24] ),
    .A1(_03312_),
    .S(net30),
    .X(_00272_));
 sg13g2_a22oi_1 _10934_ (.Y(_03313_),
    .B1(_02440_),
    .B2(_02951_),
    .A2(_02310_),
    .A1(_03068_));
 sg13g2_nor2_1 _10935_ (.A(_02355_),
    .B(_02260_),
    .Y(_03314_));
 sg13g2_o21ai_1 _10936_ (.B1(net215),
    .Y(_03315_),
    .A1(_02573_),
    .A2(_03314_));
 sg13g2_nand2_1 _10937_ (.Y(_03316_),
    .A(_03313_),
    .B(_03315_));
 sg13g2_a22oi_1 _10938_ (.Y(_03317_),
    .B1(_02633_),
    .B2(_02679_),
    .A2(_02201_),
    .A1(net440));
 sg13g2_or2_1 _10939_ (.X(_03318_),
    .B(_03308_),
    .A(_02679_));
 sg13g2_a22oi_1 _10940_ (.Y(_03319_),
    .B1(_02556_),
    .B2(_03318_),
    .A2(net227),
    .A1(net132));
 sg13g2_o21ai_1 _10941_ (.B1(_03319_),
    .Y(_03320_),
    .A1(net323),
    .A2(_03317_));
 sg13g2_a21oi_1 _10942_ (.A1(net205),
    .A2(_03316_),
    .Y(_03321_),
    .B1(_03320_));
 sg13g2_mux2_1 _10943_ (.A0(\clock_inst.min_c[25] ),
    .A1(_03321_),
    .S(net30),
    .X(_00273_));
 sg13g2_a21oi_1 _10944_ (.A1(_02235_),
    .A2(_02488_),
    .Y(_03322_),
    .B1(net340));
 sg13g2_o21ai_1 _10945_ (.B1(net213),
    .Y(_03323_),
    .A1(_02601_),
    .A2(_03322_));
 sg13g2_a21oi_1 _10946_ (.A1(_02828_),
    .A2(_03323_),
    .Y(_03324_),
    .B1(net199));
 sg13g2_nand2_1 _10947_ (.Y(_03325_),
    .A(_02997_),
    .B(_03170_));
 sg13g2_a22oi_1 _10948_ (.Y(_03326_),
    .B1(_03325_),
    .B2(net328),
    .A2(_02649_),
    .A1(net436));
 sg13g2_o21ai_1 _10949_ (.B1(net429),
    .Y(_03327_),
    .A1(_02206_),
    .A2(_02294_));
 sg13g2_o21ai_1 _10950_ (.B1(_03327_),
    .Y(_03328_),
    .A1(net301),
    .A2(_02661_));
 sg13g2_a22oi_1 _10951_ (.Y(_03329_),
    .B1(_03328_),
    .B2(net327),
    .A2(net411),
    .A1(_02175_));
 sg13g2_o21ai_1 _10952_ (.B1(_03329_),
    .Y(_03330_),
    .A1(_02545_),
    .A2(_03326_));
 sg13g2_nor3_1 _10953_ (.A(net73),
    .B(_03324_),
    .C(_03330_),
    .Y(_03331_));
 sg13g2_a21o_1 _10954_ (.A2(net31),
    .A1(\clock_inst.min_c[26] ),
    .B1(_03331_),
    .X(_00274_));
 sg13g2_a21oi_1 _10955_ (.A1(net440),
    .A2(_03169_),
    .Y(_03332_),
    .B1(net225));
 sg13g2_o21ai_1 _10956_ (.B1(_02856_),
    .Y(_03333_),
    .A1(net131),
    .A2(_03332_));
 sg13g2_nand2_1 _10957_ (.Y(_03334_),
    .A(net216),
    .B(_02722_));
 sg13g2_a21oi_1 _10958_ (.A1(net348),
    .A2(net485),
    .Y(_03335_),
    .B1(net315));
 sg13g2_a221oi_1 _10959_ (.B2(net353),
    .C1(_03335_),
    .B1(_03334_),
    .A1(net198),
    .Y(_03336_),
    .A2(net197));
 sg13g2_a22oi_1 _10960_ (.Y(_03337_),
    .B1(_02726_),
    .B2(net332),
    .A2(net420),
    .A1(net211));
 sg13g2_or2_1 _10961_ (.X(_03338_),
    .B(_03337_),
    .A(net334));
 sg13g2_o21ai_1 _10962_ (.B1(_03338_),
    .Y(_03339_),
    .A1(net199),
    .A2(_03336_));
 sg13g2_a21oi_1 _10963_ (.A1(net193),
    .A2(_03333_),
    .Y(_03340_),
    .B1(_03339_));
 sg13g2_nand2_1 _10964_ (.Y(_03341_),
    .A(\clock_inst.min_c[27] ),
    .B(net29));
 sg13g2_o21ai_1 _10965_ (.B1(_03341_),
    .Y(_00275_),
    .A1(net28),
    .A2(_03340_));
 sg13g2_o21ai_1 _10966_ (.B1(net349),
    .Y(_03342_),
    .A1(_02746_),
    .A2(net478));
 sg13g2_a221oi_1 _10967_ (.B2(net323),
    .C1(_02718_),
    .B1(_03342_),
    .A1(net231),
    .Y(_03343_),
    .A2(net316));
 sg13g2_a21oi_1 _10968_ (.A1(net350),
    .A2(net307),
    .Y(_03344_),
    .B1(_02532_));
 sg13g2_nor2_1 _10969_ (.A(net423),
    .B(_02387_),
    .Y(_03345_));
 sg13g2_o21ai_1 _10970_ (.B1(net226),
    .Y(_03346_),
    .A1(net301),
    .A2(net411));
 sg13g2_a22oi_1 _10971_ (.Y(_03347_),
    .B1(_03345_),
    .B2(_03346_),
    .A2(_03344_),
    .A1(net203));
 sg13g2_o21ai_1 _10972_ (.B1(_02717_),
    .Y(_03348_),
    .A1(net413),
    .A2(net197));
 sg13g2_nand2_1 _10973_ (.Y(_03349_),
    .A(net310),
    .B(_03017_));
 sg13g2_nand3_1 _10974_ (.B(_03348_),
    .C(_03349_),
    .A(net319),
    .Y(_03350_));
 sg13g2_o21ai_1 _10975_ (.B1(_03350_),
    .Y(_03351_),
    .A1(net338),
    .A2(_03347_));
 sg13g2_o21ai_1 _10976_ (.B1(_03351_),
    .Y(_03352_),
    .A1(net133),
    .A2(_03343_));
 sg13g2_nand2_1 _10977_ (.Y(_03353_),
    .A(\clock_inst.min_c[28] ),
    .B(net29));
 sg13g2_o21ai_1 _10978_ (.B1(_03353_),
    .Y(_00276_),
    .A1(_03225_),
    .A2(_03352_));
 sg13g2_inv_1 _10979_ (.Y(_03354_),
    .A(\clock_inst.min_c[29] ));
 sg13g2_o21ai_1 _10980_ (.B1(_02939_),
    .Y(_03355_),
    .A1(_02329_),
    .A2(net307));
 sg13g2_nor4_1 _10981_ (.A(_02356_),
    .B(net343),
    .C(_02757_),
    .D(_03355_),
    .Y(_03356_));
 sg13g2_nor3_1 _10982_ (.A(_02258_),
    .B(_02542_),
    .C(_03356_),
    .Y(_03357_));
 sg13g2_a21oi_1 _10983_ (.A1(net334),
    .A2(_02548_),
    .Y(_03358_),
    .B1(_02947_));
 sg13g2_nand2_1 _10984_ (.Y(_03359_),
    .A(_02483_),
    .B(_02635_));
 sg13g2_o21ai_1 _10985_ (.B1(_03359_),
    .Y(_03360_),
    .A1(net338),
    .A2(_03358_));
 sg13g2_a22oi_1 _10986_ (.Y(_03361_),
    .B1(_02635_),
    .B2(net299),
    .A2(_02301_),
    .A1(net194));
 sg13g2_o21ai_1 _10987_ (.B1(net483),
    .Y(_03362_),
    .A1(_02209_),
    .A2(net337));
 sg13g2_nand2_1 _10988_ (.Y(_03363_),
    .A(_02756_),
    .B(_03362_));
 sg13g2_o21ai_1 _10989_ (.B1(_03072_),
    .Y(_03364_),
    .A1(net206),
    .A2(_02670_));
 sg13g2_a221oi_1 _10990_ (.B2(net314),
    .C1(net212),
    .B1(_03364_),
    .A1(_02411_),
    .Y(_03365_),
    .A2(_03363_));
 sg13g2_a21oi_1 _10991_ (.A1(net208),
    .A2(_03361_),
    .Y(_03366_),
    .B1(_03365_));
 sg13g2_a21oi_1 _10992_ (.A1(_02463_),
    .A2(_03360_),
    .Y(_03367_),
    .B1(_03366_));
 sg13g2_a22oi_1 _10993_ (.Y(_00277_),
    .B1(_03357_),
    .B2(_03367_),
    .A2(net41),
    .A1(_03354_));
 sg13g2_inv_1 _10994_ (.Y(_03368_),
    .A(\clock_inst.min_c[2] ));
 sg13g2_o21ai_1 _10995_ (.B1(_02845_),
    .Y(_03369_),
    .A1(_02874_),
    .A2(_02398_));
 sg13g2_nand2_1 _10996_ (.Y(_03370_),
    .A(_02402_),
    .B(_02996_));
 sg13g2_a21oi_1 _10997_ (.A1(_03173_),
    .A2(_03370_),
    .Y(_03371_),
    .B1(net409));
 sg13g2_a21oi_1 _10998_ (.A1(_03003_),
    .A2(_02376_),
    .Y(_03372_),
    .B1(_03371_));
 sg13g2_nor2_1 _10999_ (.A(net130),
    .B(_03372_),
    .Y(_03373_));
 sg13g2_a221oi_1 _11000_ (.B2(net337),
    .C1(_03373_),
    .B1(_03369_),
    .A1(_02532_),
    .Y(_03374_),
    .A2(_02649_));
 sg13g2_nor3_1 _11001_ (.A(net350),
    .B(_02378_),
    .C(_03245_),
    .Y(_03375_));
 sg13g2_a21o_1 _11002_ (.A2(_03202_),
    .A1(_02833_),
    .B1(_03375_),
    .X(_03376_));
 sg13g2_a21oi_1 _11003_ (.A1(_02610_),
    .A2(_02473_),
    .Y(_03377_),
    .B1(net231));
 sg13g2_nand2_1 _11004_ (.Y(_03378_),
    .A(net318),
    .B(_03377_));
 sg13g2_o21ai_1 _11005_ (.B1(_03378_),
    .Y(_03379_),
    .A1(net309),
    .A2(_03376_));
 sg13g2_a21oi_1 _11006_ (.A1(net425),
    .A2(_02659_),
    .Y(_03380_),
    .B1(_02521_));
 sg13g2_o21ai_1 _11007_ (.B1(_02945_),
    .Y(_03381_),
    .A1(_02881_),
    .A2(_03380_));
 sg13g2_a21oi_1 _11008_ (.A1(net205),
    .A2(_03379_),
    .Y(_03382_),
    .B1(_03381_));
 sg13g2_a22oi_1 _11009_ (.Y(_00278_),
    .B1(_03374_),
    .B2(_03382_),
    .A2(net41),
    .A1(_03368_));
 sg13g2_inv_1 _11010_ (.Y(_03383_),
    .A(\clock_inst.min_c[30] ));
 sg13g2_a21oi_1 _11011_ (.A1(_02202_),
    .A2(_02665_),
    .Y(_03384_),
    .B1(net328));
 sg13g2_nand2_1 _11012_ (.Y(_03385_),
    .A(net308),
    .B(_02281_));
 sg13g2_nand2_1 _11013_ (.Y(_03386_),
    .A(_02449_),
    .B(_02646_));
 sg13g2_o21ai_1 _11014_ (.B1(net317),
    .Y(_03387_),
    .A1(_02409_),
    .A2(_02267_));
 sg13g2_nand3_1 _11015_ (.B(_03386_),
    .C(_03387_),
    .A(_03385_),
    .Y(_03388_));
 sg13g2_o21ai_1 _11016_ (.B1(net354),
    .Y(_03389_),
    .A1(_03384_),
    .A2(_03388_));
 sg13g2_nand2_1 _11017_ (.Y(_03390_),
    .A(_02669_),
    .B(_02689_));
 sg13g2_nor2_1 _11018_ (.A(_02302_),
    .B(net321),
    .Y(_03391_));
 sg13g2_o21ai_1 _11019_ (.B1(net209),
    .Y(_03392_),
    .A1(_03026_),
    .A2(_03391_));
 sg13g2_o21ai_1 _11020_ (.B1(net201),
    .Y(_03393_),
    .A1(net197),
    .A2(net225));
 sg13g2_nand3_1 _11021_ (.B(_03392_),
    .C(_03393_),
    .A(net345),
    .Y(_03394_));
 sg13g2_a22oi_1 _11022_ (.Y(_03395_),
    .B1(_03394_),
    .B2(net130),
    .A2(_03390_),
    .A1(net128));
 sg13g2_nand3_1 _11023_ (.B(_03389_),
    .C(_03395_),
    .A(net71),
    .Y(_03396_));
 sg13g2_o21ai_1 _11024_ (.B1(_03396_),
    .Y(_00279_),
    .A1(_03383_),
    .A2(net38));
 sg13g2_inv_1 _11025_ (.Y(_03397_),
    .A(\clock_inst.min_c[31] ));
 sg13g2_nand2_1 _11026_ (.Y(_03398_),
    .A(_02175_),
    .B(_02353_));
 sg13g2_o21ai_1 _11027_ (.B1(net219),
    .Y(_03399_),
    .A1(_02340_),
    .A2(_03153_));
 sg13g2_a21oi_1 _11028_ (.A1(_03398_),
    .A2(_03399_),
    .Y(_03400_),
    .B1(_02589_));
 sg13g2_o21ai_1 _11029_ (.B1(_02456_),
    .Y(_03401_),
    .A1(_02947_),
    .A2(_02986_));
 sg13g2_nand2_1 _11030_ (.Y(_03402_),
    .A(_02230_),
    .B(_03401_));
 sg13g2_o21ai_1 _11031_ (.B1(net214),
    .Y(_03403_),
    .A1(_03400_),
    .A2(_03402_));
 sg13g2_nand2_1 _11032_ (.Y(_03404_),
    .A(_02744_),
    .B(_02792_));
 sg13g2_o21ai_1 _11033_ (.B1(_02580_),
    .Y(_03405_),
    .A1(_02711_),
    .A2(_02539_));
 sg13g2_a221oi_1 _11034_ (.B2(_03405_),
    .C1(_02427_),
    .B1(_03404_),
    .A1(net230),
    .Y(_03406_),
    .A2(net196));
 sg13g2_a22oi_1 _11035_ (.Y(_00280_),
    .B1(_03403_),
    .B2(_03406_),
    .A2(net41),
    .A1(_03397_));
 sg13g2_nand2_1 _11036_ (.Y(_03407_),
    .A(_02466_),
    .B(_03170_));
 sg13g2_a22oi_1 _11037_ (.Y(_03408_),
    .B1(_02379_),
    .B2(net319),
    .A2(_02284_),
    .A1(net197));
 sg13g2_nor2_1 _11038_ (.A(net128),
    .B(_03408_),
    .Y(_03409_));
 sg13g2_a221oi_1 _11039_ (.B2(_02586_),
    .C1(_03409_),
    .B1(_03407_),
    .A1(_02664_),
    .Y(_03410_),
    .A2(_02310_));
 sg13g2_nand2_1 _11040_ (.Y(_03411_),
    .A(\clock_inst.min_c[32] ),
    .B(net29));
 sg13g2_o21ai_1 _11041_ (.B1(_03411_),
    .Y(_00281_),
    .A1(_03225_),
    .A2(_03410_));
 sg13g2_nand2_1 _11042_ (.Y(_03412_),
    .A(net435),
    .B(_02159_));
 sg13g2_a21o_1 _11043_ (.A2(_03412_),
    .A1(_02606_),
    .B1(net327),
    .X(_03413_));
 sg13g2_a21oi_1 _11044_ (.A1(_02385_),
    .A2(_03413_),
    .Y(_03414_),
    .B1(_02535_));
 sg13g2_a21o_1 _11045_ (.A2(net31),
    .A1(\clock_inst.min_c[33] ),
    .B1(_03414_),
    .X(_00282_));
 sg13g2_inv_1 _11046_ (.Y(_03415_),
    .A(\clock_inst.min_c[36] ));
 sg13g2_nor2_1 _11047_ (.A(_02371_),
    .B(_03143_),
    .Y(_03416_));
 sg13g2_o21ai_1 _11048_ (.B1(net71),
    .Y(_03417_),
    .A1(_03149_),
    .A2(_03416_));
 sg13g2_o21ai_1 _11049_ (.B1(_03417_),
    .Y(_00283_),
    .A1(_03415_),
    .A2(net38));
 sg13g2_a21oi_1 _11050_ (.A1(_02215_),
    .A2(_02364_),
    .Y(_03418_),
    .B1(net436));
 sg13g2_nor2_1 _11051_ (.A(_02255_),
    .B(_03418_),
    .Y(_03419_));
 sg13g2_a22oi_1 _11052_ (.Y(_03420_),
    .B1(_02540_),
    .B2(net411),
    .A2(_02324_),
    .A1(net312));
 sg13g2_o21ai_1 _11053_ (.B1(_02832_),
    .Y(_03421_),
    .A1(net209),
    .A2(_03420_));
 sg13g2_or3_1 _11054_ (.A(net314),
    .B(_03419_),
    .C(_03421_),
    .X(_03422_));
 sg13g2_nand3_1 _11055_ (.B(net225),
    .C(net315),
    .A(net346),
    .Y(_03423_));
 sg13g2_nand3_1 _11056_ (.B(_02308_),
    .C(_03264_),
    .A(net129),
    .Y(_03424_));
 sg13g2_nand3_1 _11057_ (.B(_03423_),
    .C(_03424_),
    .A(net193),
    .Y(_03425_));
 sg13g2_a22oi_1 _11058_ (.Y(_03426_),
    .B1(_03422_),
    .B2(_03425_),
    .A2(_02642_),
    .A1(_02181_));
 sg13g2_nand2_1 _11059_ (.Y(_03427_),
    .A(\clock_inst.min_c[37] ),
    .B(net33));
 sg13g2_o21ai_1 _11060_ (.B1(_03427_),
    .Y(_00284_),
    .A1(net28),
    .A2(_03426_));
 sg13g2_inv_1 _11061_ (.Y(_03428_),
    .A(\clock_inst.min_c[38] ));
 sg13g2_a22oi_1 _11062_ (.Y(_03429_),
    .B1(_02840_),
    .B2(_02232_),
    .A2(_02375_),
    .A1(_02294_));
 sg13g2_inv_1 _11063_ (.Y(_03430_),
    .A(_03429_));
 sg13g2_a21oi_1 _11064_ (.A1(net497),
    .A2(_02702_),
    .Y(_03431_),
    .B1(_03314_));
 sg13g2_o21ai_1 _11065_ (.B1(_02867_),
    .Y(_03432_),
    .A1(_02558_),
    .A2(_03431_));
 sg13g2_a21oi_1 _11066_ (.A1(net212),
    .A2(_03430_),
    .Y(_03433_),
    .B1(_03432_));
 sg13g2_a21oi_1 _11067_ (.A1(net207),
    .A2(_02769_),
    .Y(_03434_),
    .B1(net315));
 sg13g2_a21oi_1 _11068_ (.A1(net439),
    .A2(_02361_),
    .Y(_03435_),
    .B1(net297));
 sg13g2_o21ai_1 _11069_ (.B1(net337),
    .Y(_03436_),
    .A1(net351),
    .A2(_02228_));
 sg13g2_o21ai_1 _11070_ (.B1(_03436_),
    .Y(_03437_),
    .A1(_02439_),
    .A2(_03435_));
 sg13g2_nor3_1 _11071_ (.A(net319),
    .B(_03434_),
    .C(_03437_),
    .Y(_03438_));
 sg13g2_a21oi_1 _11072_ (.A1(net217),
    .A2(_03433_),
    .Y(_03439_),
    .B1(_03438_));
 sg13g2_nor2_1 _11073_ (.A(_03214_),
    .B(_03439_),
    .Y(_03440_));
 sg13g2_a21oi_1 _11074_ (.A1(_03428_),
    .A2(net39),
    .Y(_00285_),
    .B1(_03440_));
 sg13g2_nor3_1 _11075_ (.A(net226),
    .B(_02228_),
    .C(_02619_),
    .Y(_03441_));
 sg13g2_o21ai_1 _11076_ (.B1(_02196_),
    .Y(_03442_),
    .A1(_03068_),
    .A2(_02751_));
 sg13g2_o21ai_1 _11077_ (.B1(_03442_),
    .Y(_03443_),
    .A1(_02892_),
    .A2(_03441_));
 sg13g2_nand2_1 _11078_ (.Y(_03444_),
    .A(_02218_),
    .B(_02492_));
 sg13g2_o21ai_1 _11079_ (.B1(_03444_),
    .Y(_03445_),
    .A1(net424),
    .A2(net295));
 sg13g2_nand2_1 _11080_ (.Y(_03446_),
    .A(_02218_),
    .B(_02222_));
 sg13g2_o21ai_1 _11081_ (.B1(_03446_),
    .Y(_03447_),
    .A1(net418),
    .A2(net204));
 sg13g2_nor3_1 _11082_ (.A(_02610_),
    .B(_02228_),
    .C(_02661_),
    .Y(_03448_));
 sg13g2_a221oi_1 _11083_ (.B2(net310),
    .C1(_03448_),
    .B1(_03447_),
    .A1(net334),
    .Y(_03449_),
    .A2(_03445_));
 sg13g2_nor2_1 _11084_ (.A(net354),
    .B(_03449_),
    .Y(_03450_));
 sg13g2_a21oi_1 _11085_ (.A1(net214),
    .A2(_03443_),
    .Y(_03451_),
    .B1(_03450_));
 sg13g2_nand2_1 _11086_ (.Y(_03452_),
    .A(\clock_inst.min_c[39] ),
    .B(net33));
 sg13g2_o21ai_1 _11087_ (.B1(_03452_),
    .Y(_00286_),
    .A1(net28),
    .A2(_03451_));
 sg13g2_a21o_1 _11088_ (.A2(_02313_),
    .A1(net328),
    .B1(_02435_),
    .X(_03453_));
 sg13g2_o21ai_1 _11089_ (.B1(_03359_),
    .Y(_03454_),
    .A1(_02228_),
    .A2(_02892_));
 sg13g2_a22oi_1 _11090_ (.Y(_03455_),
    .B1(_03454_),
    .B2(_02475_),
    .A2(_03245_),
    .A1(net201));
 sg13g2_inv_1 _11091_ (.Y(_03456_),
    .A(_03455_));
 sg13g2_a21oi_1 _11092_ (.A1(net300),
    .A2(_02588_),
    .Y(_03457_),
    .B1(_02661_));
 sg13g2_a221oi_1 _11093_ (.B2(_02463_),
    .C1(_03457_),
    .B1(_03456_),
    .A1(net315),
    .Y(_03458_),
    .A2(_03453_));
 sg13g2_nand2_1 _11094_ (.Y(_03459_),
    .A(\clock_inst.min_c[3] ),
    .B(_02783_));
 sg13g2_o21ai_1 _11095_ (.B1(_03459_),
    .Y(_00287_),
    .A1(net28),
    .A2(_03458_));
 sg13g2_a21oi_1 _11096_ (.A1(_02188_),
    .A2(_02707_),
    .Y(_03460_),
    .B1(_02480_));
 sg13g2_o21ai_1 _11097_ (.B1(net337),
    .Y(_03461_),
    .A1(_02419_),
    .A2(_02619_));
 sg13g2_o21ai_1 _11098_ (.B1(_03461_),
    .Y(_03462_),
    .A1(_02657_),
    .A2(_03460_));
 sg13g2_o21ai_1 _11099_ (.B1(_03412_),
    .Y(_03463_),
    .A1(_02321_),
    .A2(_02744_));
 sg13g2_or2_1 _11100_ (.X(_03464_),
    .B(_03308_),
    .A(_02380_));
 sg13g2_a22oi_1 _11101_ (.Y(_03465_),
    .B1(_03464_),
    .B2(_02308_),
    .A2(_03463_),
    .A1(net203));
 sg13g2_nor2_1 _11102_ (.A(net326),
    .B(_03465_),
    .Y(_03466_));
 sg13g2_a21o_1 _11103_ (.A2(_02596_),
    .A1(_02546_),
    .B1(net489),
    .X(_03467_));
 sg13g2_o21ai_1 _11104_ (.B1(_03467_),
    .Y(_03468_),
    .A1(net426),
    .A2(_02213_));
 sg13g2_a22oi_1 _11105_ (.Y(_03469_),
    .B1(net298),
    .B2(net411),
    .A2(net312),
    .A1(net434));
 sg13g2_nor2_1 _11106_ (.A(net322),
    .B(_03469_),
    .Y(_03470_));
 sg13g2_a221oi_1 _11107_ (.B2(net310),
    .C1(_03470_),
    .B1(_03468_),
    .A1(net339),
    .Y(_03471_),
    .A2(net201));
 sg13g2_nor2_1 _11108_ (.A(net130),
    .B(_03471_),
    .Y(_03472_));
 sg13g2_nor4_1 _11109_ (.A(net72),
    .B(_03462_),
    .C(_03466_),
    .D(_03472_),
    .Y(_03473_));
 sg13g2_a21o_1 _11110_ (.A2(_02971_),
    .A1(\clock_inst.min_c[40] ),
    .B1(_03473_),
    .X(_00288_));
 sg13g2_nand2_1 _11111_ (.Y(_03474_),
    .A(_02177_),
    .B(_02368_));
 sg13g2_o21ai_1 _11112_ (.B1(net322),
    .Y(_03475_),
    .A1(net211),
    .A2(net297));
 sg13g2_o21ai_1 _11113_ (.B1(_03475_),
    .Y(_03476_),
    .A1(net331),
    .A2(_03474_));
 sg13g2_o21ai_1 _11114_ (.B1(_02219_),
    .Y(_03477_),
    .A1(_02287_),
    .A2(net420));
 sg13g2_nand2_1 _11115_ (.Y(_03478_),
    .A(_02826_),
    .B(_03477_));
 sg13g2_a22oi_1 _11116_ (.Y(_03479_),
    .B1(_03478_),
    .B2(_02272_),
    .A2(_03476_),
    .A1(net129));
 sg13g2_nand3_1 _11117_ (.B(_02204_),
    .C(_02374_),
    .A(net415),
    .Y(_03480_));
 sg13g2_nand3_1 _11118_ (.B(net349),
    .C(_02301_),
    .A(_02437_),
    .Y(_03481_));
 sg13g2_nand2_1 _11119_ (.Y(_03482_),
    .A(_03480_),
    .B(_03481_));
 sg13g2_nand2_1 _11120_ (.Y(_03483_),
    .A(_02889_),
    .B(_02689_));
 sg13g2_a22oi_1 _11121_ (.Y(_03484_),
    .B1(_03483_),
    .B2(_02679_),
    .A2(_03482_),
    .A1(net326));
 sg13g2_o21ai_1 _11122_ (.B1(_03484_),
    .Y(_03485_),
    .A1(net133),
    .A2(_03479_));
 sg13g2_mux2_1 _11123_ (.A0(\clock_inst.min_c[41] ),
    .A1(_03485_),
    .S(net30),
    .X(_00289_));
 sg13g2_a21oi_1 _11124_ (.A1(net207),
    .A2(_02317_),
    .Y(_03486_),
    .B1(net416));
 sg13g2_a21oi_1 _11125_ (.A1(_02361_),
    .A2(_03170_),
    .Y(_03487_),
    .B1(_02402_));
 sg13g2_a21oi_1 _11126_ (.A1(_02639_),
    .A2(_02702_),
    .Y(_03488_),
    .B1(_03487_));
 sg13g2_nor2_1 _11127_ (.A(net346),
    .B(_03488_),
    .Y(_03489_));
 sg13g2_a21oi_1 _11128_ (.A1(net309),
    .A2(_03486_),
    .Y(_03490_),
    .B1(_03489_));
 sg13g2_o21ai_1 _11129_ (.B1(_02236_),
    .Y(_03491_),
    .A1(net209),
    .A2(net203));
 sg13g2_nor2_1 _11130_ (.A(_02501_),
    .B(_02532_),
    .Y(_03492_));
 sg13g2_a21oi_1 _11131_ (.A1(net335),
    .A2(_02439_),
    .Y(_03493_),
    .B1(net435));
 sg13g2_nor3_1 _11132_ (.A(net303),
    .B(net317),
    .C(_03493_),
    .Y(_03494_));
 sg13g2_a21oi_1 _11133_ (.A1(_02382_),
    .A2(_03492_),
    .Y(_03495_),
    .B1(_03494_));
 sg13g2_a22oi_1 _11134_ (.Y(_03496_),
    .B1(_03495_),
    .B2(net224),
    .A2(_03491_),
    .A1(net352));
 sg13g2_o21ai_1 _11135_ (.B1(_03496_),
    .Y(_03497_),
    .A1(net205),
    .A2(_03490_));
 sg13g2_nand2_1 _11136_ (.Y(_03498_),
    .A(\clock_inst.min_c[42] ),
    .B(net33));
 sg13g2_o21ai_1 _11137_ (.B1(_03498_),
    .Y(_00290_),
    .A1(net36),
    .A2(_03497_));
 sg13g2_nor2_1 _11138_ (.A(net334),
    .B(_02548_),
    .Y(_03499_));
 sg13g2_nor2_1 _11139_ (.A(_02241_),
    .B(_02362_),
    .Y(_03500_));
 sg13g2_nor2_1 _11140_ (.A(net299),
    .B(_03500_),
    .Y(_03501_));
 sg13g2_a22oi_1 _11141_ (.Y(_03502_),
    .B1(_03501_),
    .B2(_02373_),
    .A2(_03499_),
    .A1(_02867_));
 sg13g2_a21oi_1 _11142_ (.A1(net345),
    .A2(_02856_),
    .Y(_03503_),
    .B1(net301));
 sg13g2_a21oi_1 _11143_ (.A1(_02418_),
    .A2(_02556_),
    .Y(_03504_),
    .B1(_03345_));
 sg13g2_nor2_1 _11144_ (.A(net302),
    .B(_03504_),
    .Y(_03505_));
 sg13g2_nor3_1 _11145_ (.A(_02798_),
    .B(_03503_),
    .C(_03505_),
    .Y(_03506_));
 sg13g2_o21ai_1 _11146_ (.B1(_02270_),
    .Y(_03507_),
    .A1(_02896_),
    .A2(_02679_));
 sg13g2_o21ai_1 _11147_ (.B1(_03507_),
    .Y(_03508_),
    .A1(net199),
    .A2(_03506_));
 sg13g2_a21oi_1 _11148_ (.A1(_03090_),
    .A2(_03502_),
    .Y(_03509_),
    .B1(_03508_));
 sg13g2_nand2_1 _11149_ (.Y(_03510_),
    .A(\clock_inst.min_c[43] ),
    .B(_02783_));
 sg13g2_o21ai_1 _11150_ (.B1(_03510_),
    .Y(_00291_),
    .A1(_02520_),
    .A2(_03509_));
 sg13g2_nor3_1 _11151_ (.A(net209),
    .B(_02556_),
    .C(_02513_),
    .Y(_03511_));
 sg13g2_nand2_1 _11152_ (.Y(_03512_),
    .A(net414),
    .B(net481));
 sg13g2_a21oi_1 _11153_ (.A1(_02223_),
    .A2(_03512_),
    .Y(_03513_),
    .B1(net334));
 sg13g2_nor3_1 _11154_ (.A(net311),
    .B(_03511_),
    .C(_03513_),
    .Y(_03514_));
 sg13g2_a21oi_1 _11155_ (.A1(net411),
    .A2(net201),
    .Y(_03515_),
    .B1(_03098_));
 sg13g2_o21ai_1 _11156_ (.B1(net415),
    .Y(_03516_),
    .A1(net413),
    .A2(_02717_));
 sg13g2_nand2_1 _11157_ (.Y(_03517_),
    .A(_03515_),
    .B(_03516_));
 sg13g2_a22oi_1 _11158_ (.Y(_03518_),
    .B1(_03517_),
    .B2(net208),
    .A2(_02691_),
    .A1(net311));
 sg13g2_o21ai_1 _11159_ (.B1(_03518_),
    .Y(_03519_),
    .A1(net208),
    .A2(_03514_));
 sg13g2_nand2_1 _11160_ (.Y(_03520_),
    .A(\clock_inst.min_c[44] ),
    .B(net33));
 sg13g2_o21ai_1 _11161_ (.B1(_03520_),
    .Y(_00292_),
    .A1(net36),
    .A2(_03519_));
 sg13g2_inv_1 _11162_ (.Y(_03521_),
    .A(\clock_inst.min_c[45] ));
 sg13g2_a22oi_1 _11163_ (.Y(_03522_),
    .B1(_03245_),
    .B2(net343),
    .A2(_03003_),
    .A1(_02483_));
 sg13g2_nor2_1 _11164_ (.A(net203),
    .B(_03522_),
    .Y(_03523_));
 sg13g2_nor3_1 _11165_ (.A(_02827_),
    .B(_02671_),
    .C(_03523_),
    .Y(_03524_));
 sg13g2_o21ai_1 _11166_ (.B1(_03079_),
    .Y(_03525_),
    .A1(net350),
    .A2(_02876_));
 sg13g2_a21oi_1 _11167_ (.A1(_02241_),
    .A2(_02317_),
    .Y(_03526_),
    .B1(net204));
 sg13g2_a221oi_1 _11168_ (.B2(net431),
    .C1(_03526_),
    .B1(_03525_),
    .A1(_02700_),
    .Y(_03527_),
    .A2(_02453_));
 sg13g2_a221oi_1 _11169_ (.B2(_02295_),
    .C1(_02456_),
    .B1(_02819_),
    .A1(_02317_),
    .Y(_03528_),
    .A2(_03048_));
 sg13g2_a21oi_1 _11170_ (.A1(net224),
    .A2(_03527_),
    .Y(_03529_),
    .B1(_03528_));
 sg13g2_a21oi_1 _11171_ (.A1(_02301_),
    .A2(_02445_),
    .Y(_03530_),
    .B1(_03529_));
 sg13g2_a22oi_1 _11172_ (.Y(_00293_),
    .B1(_03524_),
    .B2(_03530_),
    .A2(net41),
    .A1(_03521_));
 sg13g2_o21ai_1 _11173_ (.B1(net496),
    .Y(_03531_),
    .A1(net337),
    .A2(_02369_));
 sg13g2_o21ai_1 _11174_ (.B1(net426),
    .Y(_03532_),
    .A1(net304),
    .A2(_02673_));
 sg13g2_nand2_1 _11175_ (.Y(_03533_),
    .A(_03531_),
    .B(_03532_));
 sg13g2_a21o_1 _11176_ (.A2(net407),
    .A1(net422),
    .B1(_03194_),
    .X(_03534_));
 sg13g2_a22oi_1 _11177_ (.Y(_03535_),
    .B1(_03534_),
    .B2(net297),
    .A2(_03533_),
    .A1(net302));
 sg13g2_or2_1 _11178_ (.X(_03536_),
    .B(_03535_),
    .A(_02406_));
 sg13g2_nand4_1 _11179_ (.B(_03033_),
    .C(_02400_),
    .A(_02264_),
    .Y(_03537_),
    .D(_02635_));
 sg13g2_nor2_1 _11180_ (.A(_02807_),
    .B(_03418_),
    .Y(_03538_));
 sg13g2_o21ai_1 _11181_ (.B1(net195),
    .Y(_03539_),
    .A1(_02741_),
    .A2(_03538_));
 sg13g2_nand4_1 _11182_ (.B(_03536_),
    .C(_03537_),
    .A(_03357_),
    .Y(_03540_),
    .D(_03539_));
 sg13g2_o21ai_1 _11183_ (.B1(_03540_),
    .Y(_03541_),
    .A1(\clock_inst.min_c[46] ),
    .A2(_03023_));
 sg13g2_inv_1 _11184_ (.Y(_00294_),
    .A(_03541_));
 sg13g2_inv_1 _11185_ (.Y(_03542_),
    .A(\clock_inst.min_c[47] ));
 sg13g2_o21ai_1 _11186_ (.B1(net425),
    .Y(_03543_),
    .A1(_02327_),
    .A2(_02947_));
 sg13g2_nand4_1 _11187_ (.B(_02597_),
    .C(_02695_),
    .A(net212),
    .Y(_03544_),
    .D(_03543_));
 sg13g2_nand2_1 _11188_ (.Y(_03545_),
    .A(_02507_),
    .B(_02635_));
 sg13g2_o21ai_1 _11189_ (.B1(_03545_),
    .Y(_03546_),
    .A1(net209),
    .A2(_03269_));
 sg13g2_nor3_1 _11190_ (.A(net483),
    .B(net332),
    .C(_03062_),
    .Y(_03547_));
 sg13g2_nor2_1 _11191_ (.A(_02436_),
    .B(_02998_),
    .Y(_03548_));
 sg13g2_nor3_1 _11192_ (.A(net412),
    .B(_03547_),
    .C(_03548_),
    .Y(_03549_));
 sg13g2_or3_1 _11193_ (.A(net212),
    .B(_03546_),
    .C(_03549_),
    .X(_03550_));
 sg13g2_nand2b_1 _11194_ (.Y(_03551_),
    .B(_02945_),
    .A_N(_03523_));
 sg13g2_a221oi_1 _11195_ (.B2(_03550_),
    .C1(_03551_),
    .B1(_03544_),
    .A1(net299),
    .Y(_03552_),
    .A2(_02726_));
 sg13g2_a21oi_1 _11196_ (.A1(_03542_),
    .A2(net39),
    .Y(_00295_),
    .B1(_03552_));
 sg13g2_inv_1 _11197_ (.Y(_03553_),
    .A(\clock_inst.min_c[48] ));
 sg13g2_o21ai_1 _11198_ (.B1(_02407_),
    .Y(_03554_),
    .A1(_02679_),
    .A2(_03062_));
 sg13g2_a221oi_1 _11199_ (.B2(net424),
    .C1(_02750_),
    .B1(net204),
    .A1(_02452_),
    .Y(_03555_),
    .A2(net341));
 sg13g2_a21oi_1 _11200_ (.A1(_02767_),
    .A2(net201),
    .Y(_03556_),
    .B1(_02532_));
 sg13g2_o21ai_1 _11201_ (.B1(_03556_),
    .Y(_03557_),
    .A1(_02382_),
    .A2(_03555_));
 sg13g2_o21ai_1 _11202_ (.B1(_02236_),
    .Y(_03558_),
    .A1(_02659_),
    .A2(_02646_));
 sg13g2_o21ai_1 _11203_ (.B1(net331),
    .Y(_03559_),
    .A1(_02963_),
    .A2(net317));
 sg13g2_nand4_1 _11204_ (.B(net316),
    .C(_03558_),
    .A(net318),
    .Y(_03560_),
    .D(_03559_));
 sg13g2_o21ai_1 _11205_ (.B1(_03560_),
    .Y(_03561_),
    .A1(net354),
    .A2(_03557_));
 sg13g2_nand2_1 _11206_ (.Y(_03562_),
    .A(_03554_),
    .B(_03561_));
 sg13g2_a22oi_1 _11207_ (.Y(_00296_),
    .B1(_02263_),
    .B2(_03562_),
    .A2(net41),
    .A1(_03553_));
 sg13g2_inv_1 _11208_ (.Y(_03563_),
    .A(\clock_inst.min_c[49] ));
 sg13g2_a21oi_1 _11209_ (.A1(_02204_),
    .A2(_02306_),
    .Y(_03564_),
    .B1(net224));
 sg13g2_a21oi_1 _11210_ (.A1(net302),
    .A2(_02670_),
    .Y(_03565_),
    .B1(_02431_));
 sg13g2_o21ai_1 _11211_ (.B1(net327),
    .Y(_03566_),
    .A1(_03125_),
    .A2(_03565_));
 sg13g2_o21ai_1 _11212_ (.B1(_03566_),
    .Y(_03567_),
    .A1(_02304_),
    .A2(net313));
 sg13g2_a22oi_1 _11213_ (.Y(_03568_),
    .B1(_03567_),
    .B2(net202),
    .A2(_03564_),
    .A1(net222));
 sg13g2_a21oi_1 _11214_ (.A1(_02286_),
    .A2(_02889_),
    .Y(_03569_),
    .B1(_02608_));
 sg13g2_a21oi_1 _11215_ (.A1(net325),
    .A2(_02773_),
    .Y(_03570_),
    .B1(_03569_));
 sg13g2_o21ai_1 _11216_ (.B1(net317),
    .Y(_03571_),
    .A1(_02642_),
    .A2(_03068_));
 sg13g2_o21ai_1 _11217_ (.B1(_03571_),
    .Y(_03572_),
    .A1(_02415_),
    .A2(_03570_));
 sg13g2_a21oi_1 _11218_ (.A1(_02544_),
    .A2(_03572_),
    .Y(_03573_),
    .B1(_03381_));
 sg13g2_a22oi_1 _11219_ (.Y(_00297_),
    .B1(_03568_),
    .B2(_03573_),
    .A2(_02172_),
    .A1(_03563_));
 sg13g2_a22oi_1 _11220_ (.Y(_03574_),
    .B1(_02472_),
    .B2(net414),
    .A2(net312),
    .A1(net422));
 sg13g2_nand3_1 _11221_ (.B(_02596_),
    .C(_03574_),
    .A(net320),
    .Y(_03575_));
 sg13g2_a21oi_1 _11222_ (.A1(net489),
    .A2(_02308_),
    .Y(_03576_),
    .B1(_02679_));
 sg13g2_nand2_1 _11223_ (.Y(_03577_),
    .A(net226),
    .B(_03576_));
 sg13g2_a22oi_1 _11224_ (.Y(_03578_),
    .B1(_03575_),
    .B2(_03577_),
    .A2(net221),
    .A1(net347));
 sg13g2_nor2_1 _11225_ (.A(net496),
    .B(_02998_),
    .Y(_03579_));
 sg13g2_a21oi_1 _11226_ (.A1(net434),
    .A2(_02389_),
    .Y(_03580_),
    .B1(_03579_));
 sg13g2_a21oi_1 _11227_ (.A1(_02526_),
    .A2(_02260_),
    .Y(_03581_),
    .B1(net496));
 sg13g2_nor3_1 _11228_ (.A(net483),
    .B(_02181_),
    .C(_03581_),
    .Y(_03582_));
 sg13g2_a21oi_1 _11229_ (.A1(net415),
    .A2(_03580_),
    .Y(_03583_),
    .B1(_03582_));
 sg13g2_nand2_1 _11230_ (.Y(_03584_),
    .A(net346),
    .B(_03583_));
 sg13g2_o21ai_1 _11231_ (.B1(_03584_),
    .Y(_03585_),
    .A1(net318),
    .A2(_03578_));
 sg13g2_a221oi_1 _11232_ (.B2(net221),
    .C1(_03585_),
    .B1(net201),
    .A1(net132),
    .Y(_03586_),
    .A2(net298));
 sg13g2_nand2_1 _11233_ (.Y(_03587_),
    .A(\clock_inst.min_c[4] ),
    .B(net33));
 sg13g2_o21ai_1 _11234_ (.B1(_03587_),
    .Y(_00298_),
    .A1(net36),
    .A2(_03586_));
 sg13g2_o21ai_1 _11235_ (.B1(net408),
    .Y(_03588_),
    .A1(_02576_),
    .A2(_02445_));
 sg13g2_o21ai_1 _11236_ (.B1(_02253_),
    .Y(_03589_),
    .A1(net440),
    .A2(_03027_));
 sg13g2_a21oi_1 _11237_ (.A1(_02462_),
    .A2(_03588_),
    .Y(_03590_),
    .B1(_03589_));
 sg13g2_nor2_1 _11238_ (.A(_02984_),
    .B(_02996_),
    .Y(_03591_));
 sg13g2_nor3_1 _11239_ (.A(net424),
    .B(_02491_),
    .C(_02384_),
    .Y(_03592_));
 sg13g2_a21oi_1 _11240_ (.A1(_02303_),
    .A2(_03591_),
    .Y(_03593_),
    .B1(_03592_));
 sg13g2_a221oi_1 _11241_ (.B2(_02874_),
    .C1(_02606_),
    .B1(_03593_),
    .A1(net229),
    .Y(_03594_),
    .A2(net194));
 sg13g2_o21ai_1 _11242_ (.B1(_03594_),
    .Y(_03595_),
    .A1(_02430_),
    .A2(_03590_));
 sg13g2_nand2_1 _11243_ (.Y(_03596_),
    .A(\clock_inst.min_c[50] ),
    .B(net33));
 sg13g2_o21ai_1 _11244_ (.B1(_03596_),
    .Y(_00299_),
    .A1(net36),
    .A2(_03595_));
 sg13g2_inv_1 _11245_ (.Y(_03597_),
    .A(\clock_inst.min_c[51] ));
 sg13g2_o21ai_1 _11246_ (.B1(net209),
    .Y(_03598_),
    .A1(_02454_),
    .A2(_02284_));
 sg13g2_o21ai_1 _11247_ (.B1(_03598_),
    .Y(_03599_),
    .A1(_02601_),
    .A2(_03512_));
 sg13g2_o21ai_1 _11248_ (.B1(net353),
    .Y(_03600_),
    .A1(net220),
    .A2(_03548_));
 sg13g2_nor2_1 _11249_ (.A(net317),
    .B(_02757_),
    .Y(_03601_));
 sg13g2_a21oi_1 _11250_ (.A1(_03600_),
    .A2(_03601_),
    .Y(_03602_),
    .B1(net129));
 sg13g2_a221oi_1 _11251_ (.B2(net215),
    .C1(_03602_),
    .B1(_03599_),
    .A1(_02204_),
    .Y(_03603_),
    .A2(net317));
 sg13g2_nor2_1 _11252_ (.A(_02427_),
    .B(_03603_),
    .Y(_03604_));
 sg13g2_a21oi_1 _11253_ (.A1(_03597_),
    .A2(_02251_),
    .Y(_00300_),
    .B1(_03604_));
 sg13g2_o21ai_1 _11254_ (.B1(net343),
    .Y(_03605_),
    .A1(net420),
    .A2(_02507_));
 sg13g2_o21ai_1 _11255_ (.B1(_03605_),
    .Y(_03606_),
    .A1(_02411_),
    .A2(_02875_));
 sg13g2_o21ai_1 _11256_ (.B1(net301),
    .Y(_03607_),
    .A1(net222),
    .A2(_02750_));
 sg13g2_nand3_1 _11257_ (.B(net300),
    .C(_03607_),
    .A(_02448_),
    .Y(_03608_));
 sg13g2_a22oi_1 _11258_ (.Y(_03609_),
    .B1(_03608_),
    .B2(net306),
    .A2(_03606_),
    .A1(net326));
 sg13g2_a21oi_1 _11259_ (.A1(_03079_),
    .A2(_03609_),
    .Y(_03610_),
    .B1(net70));
 sg13g2_a21o_1 _11260_ (.A2(net31),
    .A1(\clock_inst.min_c[52] ),
    .B1(_03610_),
    .X(_00301_));
 sg13g2_a21o_1 _11261_ (.A2(_02474_),
    .A1(_02410_),
    .B1(_02633_),
    .X(_03611_));
 sg13g2_a21oi_1 _11262_ (.A1(_03235_),
    .A2(_03611_),
    .Y(_03612_),
    .B1(net70));
 sg13g2_a21o_1 _11263_ (.A2(net31),
    .A1(\clock_inst.min_c[53] ),
    .B1(_03612_),
    .X(_00302_));
 sg13g2_o21ai_1 _11264_ (.B1(net485),
    .Y(_03613_),
    .A1(_02509_),
    .A2(_03096_));
 sg13g2_a22oi_1 _11265_ (.Y(_03614_),
    .B1(_03613_),
    .B2(net199),
    .A2(_02365_),
    .A1(net195));
 sg13g2_nor3_1 _11266_ (.A(net497),
    .B(net410),
    .C(_02561_),
    .Y(_03615_));
 sg13g2_o21ai_1 _11267_ (.B1(_02175_),
    .Y(_03616_),
    .A1(_02513_),
    .A2(_02954_));
 sg13g2_o21ai_1 _11268_ (.B1(_03616_),
    .Y(_03617_),
    .A1(_02175_),
    .A2(_02312_));
 sg13g2_or2_1 _11269_ (.X(_03618_),
    .B(_03617_),
    .A(_03615_));
 sg13g2_a21oi_1 _11270_ (.A1(net303),
    .A2(net304),
    .Y(_03619_),
    .B1(_02673_));
 sg13g2_nor2_1 _11271_ (.A(_02503_),
    .B(_03619_),
    .Y(_03620_));
 sg13g2_a221oi_1 _11272_ (.B2(net327),
    .C1(_03620_),
    .B1(_03618_),
    .A1(_02301_),
    .Y(_03621_),
    .A2(_02365_));
 sg13g2_o21ai_1 _11273_ (.B1(_03621_),
    .Y(_03622_),
    .A1(net306),
    .A2(_03614_));
 sg13g2_mux2_1 _11274_ (.A0(\clock_inst.min_c[5] ),
    .A1(_03622_),
    .S(net30),
    .X(_00303_));
 sg13g2_a22oi_1 _11275_ (.Y(_03623_),
    .B1(_03264_),
    .B2(net305),
    .A2(_02491_),
    .A1(net342));
 sg13g2_a221oi_1 _11276_ (.B2(net305),
    .C1(net424),
    .B1(_02702_),
    .A1(_02513_),
    .Y(_03624_),
    .A2(_02361_));
 sg13g2_a21o_1 _11277_ (.A2(_03623_),
    .A1(net409),
    .B1(_03624_),
    .X(_03625_));
 sg13g2_a21oi_1 _11278_ (.A1(net489),
    .A2(_02960_),
    .Y(_03626_),
    .B1(net304));
 sg13g2_nor2_1 _11279_ (.A(net320),
    .B(_03626_),
    .Y(_03627_));
 sg13g2_nor2_1 _11280_ (.A(net482),
    .B(_03474_),
    .Y(_03628_));
 sg13g2_a21oi_1 _11281_ (.A1(net483),
    .A2(net332),
    .Y(_03629_),
    .B1(_03628_));
 sg13g2_nor2_1 _11282_ (.A(net428),
    .B(_03629_),
    .Y(_03630_));
 sg13g2_nor4_1 _11283_ (.A(net296),
    .B(_02741_),
    .C(_03627_),
    .D(_03630_),
    .Y(_03631_));
 sg13g2_a21oi_1 _11284_ (.A1(net223),
    .A2(_03625_),
    .Y(_03632_),
    .B1(_03631_));
 sg13g2_a221oi_1 _11285_ (.B2(net132),
    .C1(_03632_),
    .B1(_02284_),
    .A1(_02185_),
    .Y(_03633_),
    .A2(net196));
 sg13g2_nand2_1 _11286_ (.Y(_03634_),
    .A(\clock_inst.min_c[6] ),
    .B(net33));
 sg13g2_o21ai_1 _11287_ (.B1(_03634_),
    .Y(_00304_),
    .A1(_02520_),
    .A2(_03633_));
 sg13g2_nand2_1 _11288_ (.Y(_03635_),
    .A(_02240_),
    .B(_02299_));
 sg13g2_a21oi_1 _11289_ (.A1(_02353_),
    .A2(_03635_),
    .Y(_03636_),
    .B1(net314));
 sg13g2_o21ai_1 _11290_ (.B1(_02484_),
    .Y(_03637_),
    .A1(net440),
    .A2(_03169_));
 sg13g2_o21ai_1 _11291_ (.B1(_02816_),
    .Y(_03638_),
    .A1(_03636_),
    .A2(_03637_));
 sg13g2_a21oi_1 _11292_ (.A1(net421),
    .A2(_02772_),
    .Y(_03639_),
    .B1(_02839_));
 sg13g2_o21ai_1 _11293_ (.B1(net216),
    .Y(_03640_),
    .A1(_02448_),
    .A2(_02412_));
 sg13g2_nand2_1 _11294_ (.Y(_03641_),
    .A(net341),
    .B(_03640_));
 sg13g2_o21ai_1 _11295_ (.B1(_03641_),
    .Y(_03642_),
    .A1(net425),
    .A2(_03639_));
 sg13g2_a22oi_1 _11296_ (.Y(_03643_),
    .B1(_03642_),
    .B2(net223),
    .A2(_02380_),
    .A1(net221));
 sg13g2_a21oi_1 _11297_ (.A1(_03638_),
    .A2(_03643_),
    .Y(_03644_),
    .B1(net70));
 sg13g2_a21o_1 _11298_ (.A2(_02971_),
    .A1(\clock_inst.min_c[7] ),
    .B1(_03644_),
    .X(_00305_));
 sg13g2_a21oi_1 _11299_ (.A1(_02528_),
    .A2(_03444_),
    .Y(_03645_),
    .B1(_02517_));
 sg13g2_o21ai_1 _11300_ (.B1(net478),
    .Y(_03646_),
    .A1(_02187_),
    .A2(_02998_));
 sg13g2_a21oi_1 _11301_ (.A1(net295),
    .A2(net313),
    .Y(_03647_),
    .B1(net301));
 sg13g2_a221oi_1 _11302_ (.B2(net198),
    .C1(_03647_),
    .B1(_03646_),
    .A1(net297),
    .Y(_03648_),
    .A2(net227));
 sg13g2_a21oi_1 _11303_ (.A1(net206),
    .A2(_03635_),
    .Y(_03649_),
    .B1(net303));
 sg13g2_o21ai_1 _11304_ (.B1(net319),
    .Y(_03650_),
    .A1(_02532_),
    .A2(_03649_));
 sg13g2_o21ai_1 _11305_ (.B1(_03650_),
    .Y(_03651_),
    .A1(net338),
    .A2(_03648_));
 sg13g2_nor3_1 _11306_ (.A(net73),
    .B(_03645_),
    .C(_03651_),
    .Y(_03652_));
 sg13g2_a21o_1 _11307_ (.A2(_02247_),
    .A1(\clock_inst.min_c[8] ),
    .B1(_03652_),
    .X(_00306_));
 sg13g2_inv_1 _11308_ (.Y(_03653_),
    .A(\clock_inst.min_c[9] ));
 sg13g2_nand2_1 _11309_ (.Y(_03654_),
    .A(net204),
    .B(_02858_));
 sg13g2_a21oi_1 _11310_ (.A1(net348),
    .A2(_02317_),
    .Y(_03655_),
    .B1(_03512_));
 sg13g2_a221oi_1 _11311_ (.B2(net409),
    .C1(_03655_),
    .B1(_03654_),
    .A1(_03446_),
    .Y(_03656_),
    .A2(_02659_));
 sg13g2_a21oi_1 _11312_ (.A1(_02623_),
    .A2(_02930_),
    .Y(_03657_),
    .B1(net415));
 sg13g2_nand2_1 _11313_ (.Y(_03658_),
    .A(net439),
    .B(net295));
 sg13g2_a21oi_1 _11314_ (.A1(_02665_),
    .A2(_03658_),
    .Y(_03659_),
    .B1(net413));
 sg13g2_nor3_1 _11315_ (.A(net129),
    .B(_03657_),
    .C(_03659_),
    .Y(_03660_));
 sg13g2_a21oi_1 _11316_ (.A1(net130),
    .A2(_03656_),
    .Y(_03661_),
    .B1(_03660_));
 sg13g2_o21ai_1 _11317_ (.B1(net71),
    .Y(_03662_),
    .A1(_03273_),
    .A2(_03661_));
 sg13g2_o21ai_1 _11318_ (.B1(_03662_),
    .Y(_00307_),
    .A1(_03653_),
    .A2(_02351_));
 sg13g2_buf_1 _11319_ (.A(\clock_inst.min_tile.e0[0] ),
    .X(_03663_));
 sg13g2_inv_1 _11320_ (.Y(_03664_),
    .A(_03663_));
 sg13g2_nor2_1 _11321_ (.A(_03138_),
    .B(net235),
    .Y(_03665_));
 sg13g2_xnor2_1 _11322_ (.Y(_03666_),
    .A(_02855_),
    .B(_03663_));
 sg13g2_nor2_1 _11323_ (.A(net237),
    .B(_03666_),
    .Y(_03667_));
 sg13g2_o21ai_1 _11324_ (.B1(net156),
    .Y(_03668_),
    .A1(_03665_),
    .A2(_03667_));
 sg13g2_o21ai_1 _11325_ (.B1(_03668_),
    .Y(_00308_),
    .A1(_03664_),
    .A2(net106));
 sg13g2_buf_2 _11326_ (.A(\clock_inst.min_tile.e0[10] ),
    .X(_03669_));
 sg13g2_inv_1 _11327_ (.Y(_03670_),
    .A(_03669_));
 sg13g2_buf_1 _11328_ (.A(net153),
    .X(_03671_));
 sg13g2_nand2_1 _11329_ (.Y(_03672_),
    .A(_03669_),
    .B(net104));
 sg13g2_nand2_1 _11330_ (.Y(_03673_),
    .A(_03670_),
    .B(net92));
 sg13g2_buf_1 _11331_ (.A(\clock_inst.min_tile.e0[9] ),
    .X(_03674_));
 sg13g2_nor2b_1 _11332_ (.A(_03674_),
    .B_N(net532),
    .Y(_03675_));
 sg13g2_buf_1 _11333_ (.A(_03675_),
    .X(_03676_));
 sg13g2_inv_1 _11334_ (.Y(_03677_),
    .A(_03674_));
 sg13g2_nor2_2 _11335_ (.A(net532),
    .B(_03677_),
    .Y(_03678_));
 sg13g2_buf_1 _11336_ (.A(\clock_inst.min_tile.e0[8] ),
    .X(_03679_));
 sg13g2_buf_1 _11337_ (.A(\clock_inst.min_tile.e0[7] ),
    .X(_03680_));
 sg13g2_xnor2_1 _11338_ (.Y(_03681_),
    .A(_03122_),
    .B(_03680_));
 sg13g2_buf_2 _11339_ (.A(\clock_inst.min_tile.e0[6] ),
    .X(_03682_));
 sg13g2_xor2_1 _11340_ (.B(_03682_),
    .A(_03110_),
    .X(_03683_));
 sg13g2_nor2b_1 _11341_ (.A(_03681_),
    .B_N(_03683_),
    .Y(_03684_));
 sg13g2_buf_2 _11342_ (.A(\clock_inst.min_tile.e0[1] ),
    .X(_03685_));
 sg13g2_a22oi_1 _11343_ (.Y(_03686_),
    .B1(_02901_),
    .B2(_03685_),
    .A2(_03663_),
    .A1(_02855_));
 sg13g2_nor2_1 _11344_ (.A(_02901_),
    .B(_03685_),
    .Y(_03687_));
 sg13g2_or2_1 _11345_ (.X(_03688_),
    .B(_03687_),
    .A(_03686_));
 sg13g2_buf_1 _11346_ (.A(_03688_),
    .X(_03689_));
 sg13g2_buf_1 _11347_ (.A(\clock_inst.min_tile.e0[3] ),
    .X(_03690_));
 sg13g2_inv_1 _11348_ (.Y(_03691_),
    .A(_03690_));
 sg13g2_buf_1 _11349_ (.A(\clock_inst.min_tile.e0[2] ),
    .X(_03692_));
 sg13g2_nand2_1 _11350_ (.Y(_03693_),
    .A(_02943_),
    .B(_03692_));
 sg13g2_buf_2 _11351_ (.A(\clock_inst.min_tile.e0[4] ),
    .X(_03694_));
 sg13g2_nand2_1 _11352_ (.Y(_03695_),
    .A(_03094_),
    .B(_03694_));
 sg13g2_and3_1 _11353_ (.X(_03696_),
    .A(_03691_),
    .B(_03693_),
    .C(_03695_));
 sg13g2_or2_1 _11354_ (.X(_03697_),
    .B(_03692_),
    .A(_02943_));
 sg13g2_buf_1 _11355_ (.A(_03697_),
    .X(_03698_));
 sg13g2_a221oi_1 _11356_ (.B2(_03694_),
    .C1(_03698_),
    .B1(_03094_),
    .A1(_03012_),
    .Y(_03699_),
    .A2(_03690_));
 sg13g2_a21oi_1 _11357_ (.A1(_03689_),
    .A2(_03696_),
    .Y(_03700_),
    .B1(_03699_));
 sg13g2_inv_1 _11358_ (.Y(_03701_),
    .A(_03012_));
 sg13g2_and3_1 _11359_ (.X(_03702_),
    .A(_03701_),
    .B(_03693_),
    .C(_03695_));
 sg13g2_nor2_1 _11360_ (.A(_03012_),
    .B(_03690_),
    .Y(_03703_));
 sg13g2_a22oi_1 _11361_ (.Y(_03704_),
    .B1(_03703_),
    .B2(_03695_),
    .A2(_03702_),
    .A1(_03689_));
 sg13g2_buf_1 _11362_ (.A(\clock_inst.min_tile.e0[5] ),
    .X(_03705_));
 sg13g2_or2_1 _11363_ (.X(_03706_),
    .B(_03694_),
    .A(_03094_));
 sg13g2_buf_1 _11364_ (.A(_03706_),
    .X(_03707_));
 sg13g2_and2_1 _11365_ (.A(_03705_),
    .B(_03707_),
    .X(_03708_));
 sg13g2_nand4_1 _11366_ (.B(_03700_),
    .C(_03704_),
    .A(_03684_),
    .Y(_03709_),
    .D(_03708_));
 sg13g2_and2_1 _11367_ (.A(_03108_),
    .B(_03707_),
    .X(_03710_));
 sg13g2_nand4_1 _11368_ (.B(_03700_),
    .C(_03704_),
    .A(_03684_),
    .Y(_03711_),
    .D(_03710_));
 sg13g2_inv_1 _11369_ (.Y(_03712_),
    .A(_03108_));
 sg13g2_inv_1 _11370_ (.Y(_03713_),
    .A(_03705_));
 sg13g2_nor2_1 _11371_ (.A(_03712_),
    .B(_03713_),
    .Y(_03714_));
 sg13g2_nor2_1 _11372_ (.A(_03122_),
    .B(_03680_),
    .Y(_03715_));
 sg13g2_a22oi_1 _11373_ (.Y(_03716_),
    .B1(_03122_),
    .B2(_03680_),
    .A2(_03682_),
    .A1(_03110_));
 sg13g2_nor2_1 _11374_ (.A(_03715_),
    .B(_03716_),
    .Y(_03717_));
 sg13g2_a21oi_1 _11375_ (.A1(_03684_),
    .A2(_03714_),
    .Y(_03718_),
    .B1(_03717_));
 sg13g2_nand3_1 _11376_ (.B(_03711_),
    .C(_03718_),
    .A(_03709_),
    .Y(_03719_));
 sg13g2_nand2_1 _11377_ (.Y(_03720_),
    .A(_03679_),
    .B(_03719_));
 sg13g2_o21ai_1 _11378_ (.B1(_03133_),
    .Y(_03721_),
    .A1(_03679_),
    .A2(_03719_));
 sg13g2_nand2_1 _11379_ (.Y(_03722_),
    .A(_03720_),
    .B(_03721_));
 sg13g2_mux2_1 _11380_ (.A0(_03676_),
    .A1(_03678_),
    .S(_03722_),
    .X(_03723_));
 sg13g2_mux2_1 _11381_ (.A0(_03672_),
    .A1(_03673_),
    .S(_03723_),
    .X(_03724_));
 sg13g2_a21oi_1 _11382_ (.A1(\clock_inst.min_c[10] ),
    .A2(net52),
    .Y(_03725_),
    .B1(net162));
 sg13g2_a22oi_1 _11383_ (.Y(_00309_),
    .B1(_03724_),
    .B2(_03725_),
    .A2(net69),
    .A1(_03670_));
 sg13g2_buf_1 _11384_ (.A(\clock_inst.min_tile.e0[11] ),
    .X(_03726_));
 sg13g2_inv_1 _11385_ (.Y(_03727_),
    .A(_03726_));
 sg13g2_nand2_1 _11386_ (.Y(_03728_),
    .A(_03727_),
    .B(net104));
 sg13g2_nand2_1 _11387_ (.Y(_03729_),
    .A(_03726_),
    .B(net92));
 sg13g2_nand2_1 _11388_ (.Y(_03730_),
    .A(_03669_),
    .B(_03678_));
 sg13g2_nand2_1 _11389_ (.Y(_03731_),
    .A(_03670_),
    .B(_03676_));
 sg13g2_and2_1 _11390_ (.A(_03720_),
    .B(_03721_),
    .X(_03732_));
 sg13g2_buf_1 _11391_ (.A(_03732_),
    .X(_03733_));
 sg13g2_mux2_1 _11392_ (.A0(_03730_),
    .A1(_03731_),
    .S(_03733_),
    .X(_03734_));
 sg13g2_mux2_1 _11393_ (.A0(_03728_),
    .A1(_03729_),
    .S(_03734_),
    .X(_03735_));
 sg13g2_a21oi_1 _11394_ (.A1(\clock_inst.min_c[11] ),
    .A2(net52),
    .Y(_03736_),
    .B1(net162));
 sg13g2_a22oi_1 _11395_ (.Y(_00310_),
    .B1(_03735_),
    .B2(_03736_),
    .A2(net69),
    .A1(_03727_));
 sg13g2_buf_2 _11396_ (.A(\clock_inst.min_tile.e0[12] ),
    .X(_03737_));
 sg13g2_xor2_1 _11397_ (.B(_03737_),
    .A(net532),
    .X(_03738_));
 sg13g2_nand2_1 _11398_ (.Y(_03739_),
    .A(net243),
    .B(_03738_));
 sg13g2_nand2b_1 _11399_ (.Y(_03740_),
    .B(net243),
    .A_N(_03738_));
 sg13g2_and3_1 _11400_ (.X(_03741_),
    .A(_03709_),
    .B(_03711_),
    .C(_03718_));
 sg13g2_xnor2_1 _11401_ (.Y(_03742_),
    .A(_03133_),
    .B(_03679_));
 sg13g2_nor4_1 _11402_ (.A(_02865_),
    .B(_03677_),
    .C(_03670_),
    .D(_03727_),
    .Y(_03743_));
 sg13g2_nand2b_1 _11403_ (.Y(_03744_),
    .B(_02865_),
    .A_N(_03674_));
 sg13g2_nor3_1 _11404_ (.A(_03669_),
    .B(_03726_),
    .C(_03744_),
    .Y(_03745_));
 sg13g2_nor2_1 _11405_ (.A(_03743_),
    .B(_03745_),
    .Y(_03746_));
 sg13g2_or2_1 _11406_ (.X(_03747_),
    .B(_03746_),
    .A(_03742_));
 sg13g2_nand3_1 _11407_ (.B(_03669_),
    .C(_03726_),
    .A(_03674_),
    .Y(_03748_));
 sg13g2_nor2b_1 _11408_ (.A(net532),
    .B_N(_03748_),
    .Y(_03749_));
 sg13g2_nand3_1 _11409_ (.B(_03670_),
    .C(_03727_),
    .A(_03677_),
    .Y(_03750_));
 sg13g2_a22oi_1 _11410_ (.Y(_03751_),
    .B1(net532),
    .B2(_03750_),
    .A2(_03679_),
    .A1(_03133_));
 sg13g2_or2_1 _11411_ (.X(_03752_),
    .B(_03751_),
    .A(_03749_));
 sg13g2_o21ai_1 _11412_ (.B1(_03752_),
    .Y(_03753_),
    .A1(_03741_),
    .A2(_03747_));
 sg13g2_mux2_1 _11413_ (.A0(_03739_),
    .A1(_03740_),
    .S(_03753_),
    .X(_03754_));
 sg13g2_nand2_1 _11414_ (.Y(_03755_),
    .A(\clock_inst.min_c[12] ),
    .B(_01145_));
 sg13g2_a21oi_1 _11415_ (.A1(_03754_),
    .A2(_03755_),
    .Y(_03756_),
    .B1(net239));
 sg13g2_a21o_1 _11416_ (.A2(net112),
    .A1(_03737_),
    .B1(_03756_),
    .X(_00311_));
 sg13g2_buf_1 _11417_ (.A(\clock_inst.min_tile.e0[13] ),
    .X(_03757_));
 sg13g2_inv_1 _11418_ (.Y(_03758_),
    .A(_03757_));
 sg13g2_nand2_1 _11419_ (.Y(_03759_),
    .A(_03758_),
    .B(net104));
 sg13g2_nand2_1 _11420_ (.Y(_03760_),
    .A(_03757_),
    .B(net92));
 sg13g2_nand2_1 _11421_ (.Y(_03761_),
    .A(_03737_),
    .B(_03743_));
 sg13g2_nand2b_1 _11422_ (.Y(_03762_),
    .B(_03745_),
    .A_N(_03737_));
 sg13g2_mux2_1 _11423_ (.A0(_03761_),
    .A1(_03762_),
    .S(_03733_),
    .X(_03763_));
 sg13g2_mux2_1 _11424_ (.A0(_03759_),
    .A1(_03760_),
    .S(_03763_),
    .X(_03764_));
 sg13g2_a21oi_1 _11425_ (.A1(\clock_inst.min_c[13] ),
    .A2(net52),
    .Y(_03765_),
    .B1(net162));
 sg13g2_a22oi_1 _11426_ (.Y(_00312_),
    .B1(_03764_),
    .B2(_03765_),
    .A2(net69),
    .A1(_03758_));
 sg13g2_inv_1 _11427_ (.Y(_03766_),
    .A(_03679_));
 sg13g2_or2_1 _11428_ (.X(_03767_),
    .B(_03716_),
    .A(_03715_));
 sg13g2_nand2_1 _11429_ (.Y(_03768_),
    .A(_03766_),
    .B(_03767_));
 sg13g2_nor2_1 _11430_ (.A(_03766_),
    .B(_03767_),
    .Y(_03769_));
 sg13g2_a21oi_1 _11431_ (.A1(_03133_),
    .A2(_03768_),
    .Y(_03770_),
    .B1(_03769_));
 sg13g2_and2_1 _11432_ (.A(_03737_),
    .B(_03757_),
    .X(_03771_));
 sg13g2_buf_1 _11433_ (.A(_03771_),
    .X(_03772_));
 sg13g2_nand3_1 _11434_ (.B(_03678_),
    .C(_03772_),
    .A(_03726_),
    .Y(_03773_));
 sg13g2_nor2_1 _11435_ (.A(_03737_),
    .B(_03757_),
    .Y(_03774_));
 sg13g2_nand2_1 _11436_ (.Y(_03775_),
    .A(net532),
    .B(_03774_));
 sg13g2_o21ai_1 _11437_ (.B1(_03775_),
    .Y(_03776_),
    .A1(_03770_),
    .A2(_03773_));
 sg13g2_nand2_1 _11438_ (.Y(_03777_),
    .A(_03669_),
    .B(_03776_));
 sg13g2_o21ai_1 _11439_ (.B1(_03693_),
    .Y(_03778_),
    .A1(_03686_),
    .A2(_03687_));
 sg13g2_nand3_1 _11440_ (.B(_03698_),
    .C(_03778_),
    .A(_03690_),
    .Y(_03779_));
 sg13g2_nand2_1 _11441_ (.Y(_03780_),
    .A(_03694_),
    .B(_03108_));
 sg13g2_nand2_1 _11442_ (.Y(_03781_),
    .A(_03094_),
    .B(_03108_));
 sg13g2_a21oi_1 _11443_ (.A1(_03698_),
    .A2(_03778_),
    .Y(_03782_),
    .B1(_03690_));
 sg13g2_a221oi_1 _11444_ (.B2(_03781_),
    .C1(_03782_),
    .B1(_03780_),
    .A1(_03701_),
    .Y(_03783_),
    .A2(_03779_));
 sg13g2_nand2_1 _11445_ (.Y(_03784_),
    .A(_03694_),
    .B(_03705_));
 sg13g2_nand2_1 _11446_ (.Y(_03785_),
    .A(_03094_),
    .B(_03705_));
 sg13g2_a221oi_1 _11447_ (.B2(_03785_),
    .C1(_03782_),
    .B1(_03784_),
    .A1(_03701_),
    .Y(_03786_),
    .A2(_03779_));
 sg13g2_a21oi_1 _11448_ (.A1(_03712_),
    .A2(_03713_),
    .Y(_03787_),
    .B1(_03695_));
 sg13g2_or4_1 _11449_ (.A(_03783_),
    .B(_03786_),
    .C(_03714_),
    .D(_03787_),
    .X(_03788_));
 sg13g2_buf_8 _11450_ (.A(_03788_),
    .X(_03789_));
 sg13g2_nand2b_1 _11451_ (.Y(_03790_),
    .B(_03683_),
    .A_N(_03681_));
 sg13g2_nor2_1 _11452_ (.A(_03790_),
    .B(_03747_),
    .Y(_03791_));
 sg13g2_nand3_1 _11453_ (.B(_03772_),
    .C(_03791_),
    .A(_03789_),
    .Y(_03792_));
 sg13g2_a21oi_2 _11454_ (.B1(net532),
    .Y(_03793_),
    .A2(_03792_),
    .A1(_03777_));
 sg13g2_nand4_1 _11455_ (.B(_03676_),
    .C(_03774_),
    .A(_03727_),
    .Y(_03794_),
    .D(_03770_));
 sg13g2_a221oi_1 _11456_ (.B2(_03789_),
    .C1(_03794_),
    .B1(_03791_),
    .A1(_03669_),
    .Y(_03795_),
    .A2(_03776_));
 sg13g2_buf_1 _11457_ (.A(_03795_),
    .X(_03796_));
 sg13g2_buf_2 _11458_ (.A(\clock_inst.min_tile.e0[14] ),
    .X(_03797_));
 sg13g2_nor2_1 _11459_ (.A(_03797_),
    .B(net107),
    .Y(_03798_));
 sg13g2_o21ai_1 _11460_ (.B1(_03798_),
    .Y(_03799_),
    .A1(_03793_),
    .A2(_03796_));
 sg13g2_nand2_1 _11461_ (.Y(_03800_),
    .A(\clock_inst.min_c[14] ),
    .B(net96));
 sg13g2_a21oi_1 _11462_ (.A1(_03799_),
    .A2(_03800_),
    .Y(_03801_),
    .B1(net136));
 sg13g2_nor3_1 _11463_ (.A(net96),
    .B(_03793_),
    .C(_03796_),
    .Y(_03802_));
 sg13g2_o21ai_1 _11464_ (.B1(_03797_),
    .Y(_03803_),
    .A1(net145),
    .A2(_03802_));
 sg13g2_nand2b_1 _11465_ (.Y(_00313_),
    .B(_03803_),
    .A_N(_03801_));
 sg13g2_buf_1 _11466_ (.A(\clock_inst.min_tile.e0[15] ),
    .X(_03804_));
 sg13g2_inv_1 _11467_ (.Y(_03805_),
    .A(_03804_));
 sg13g2_nand2_1 _11468_ (.Y(_03806_),
    .A(_03805_),
    .B(net92));
 sg13g2_nand2_1 _11469_ (.Y(_03807_),
    .A(_03804_),
    .B(net92));
 sg13g2_inv_1 _11470_ (.Y(_03808_),
    .A(_03745_));
 sg13g2_nor3_1 _11471_ (.A(_03737_),
    .B(_03757_),
    .C(_03797_),
    .Y(_03809_));
 sg13g2_inv_1 _11472_ (.Y(_03810_),
    .A(_03809_));
 sg13g2_nor2_1 _11473_ (.A(_03808_),
    .B(_03810_),
    .Y(_03811_));
 sg13g2_a22oi_1 _11474_ (.Y(_03812_),
    .B1(_03811_),
    .B2(_03733_),
    .A2(_03793_),
    .A1(_03797_));
 sg13g2_mux2_1 _11475_ (.A0(_03806_),
    .A1(_03807_),
    .S(_03812_),
    .X(_03813_));
 sg13g2_a21oi_1 _11476_ (.A1(\clock_inst.min_c[15] ),
    .A2(net52),
    .Y(_03814_),
    .B1(net162));
 sg13g2_a22oi_1 _11477_ (.Y(_00314_),
    .B1(_03813_),
    .B2(_03814_),
    .A2(net69),
    .A1(_03805_));
 sg13g2_buf_1 _11478_ (.A(\clock_inst.min_tile.e0[16] ),
    .X(_03815_));
 sg13g2_nand3_1 _11479_ (.B(_03805_),
    .C(_03809_),
    .A(_02866_),
    .Y(_03816_));
 sg13g2_nor2b_1 _11480_ (.A(_02866_),
    .B_N(_03797_),
    .Y(_03817_));
 sg13g2_nand3_1 _11481_ (.B(_03772_),
    .C(_03817_),
    .A(_03804_),
    .Y(_03818_));
 sg13g2_mux2_1 _11482_ (.A0(_03816_),
    .A1(_03818_),
    .S(_03753_),
    .X(_03819_));
 sg13g2_xor2_1 _11483_ (.B(_03819_),
    .A(_03815_),
    .X(_03820_));
 sg13g2_nand2_1 _11484_ (.Y(_03821_),
    .A(\clock_inst.min_c[16] ),
    .B(net237));
 sg13g2_o21ai_1 _11485_ (.B1(_03821_),
    .Y(_03822_),
    .A1(net98),
    .A2(_03820_));
 sg13g2_mux2_1 _11486_ (.A0(_03815_),
    .A1(_03822_),
    .S(net146),
    .X(_00315_));
 sg13g2_inv_1 _11487_ (.Y(_03823_),
    .A(\clock_inst.min_tile.e0[17] ));
 sg13g2_inv_1 _11488_ (.Y(_03824_),
    .A(\clock_inst.min_c[17] ));
 sg13g2_nor2_1 _11489_ (.A(_03823_),
    .B(net95),
    .Y(_03825_));
 sg13g2_nor2_1 _11490_ (.A(\clock_inst.min_tile.e0[17] ),
    .B(net95),
    .Y(_03826_));
 sg13g2_nor4_1 _11491_ (.A(_03804_),
    .B(_03815_),
    .C(_03808_),
    .D(_03810_),
    .Y(_03827_));
 sg13g2_and2_1 _11492_ (.A(_03815_),
    .B(_03772_),
    .X(_03828_));
 sg13g2_and3_1 _11493_ (.X(_03829_),
    .A(_03804_),
    .B(_03753_),
    .C(_03817_));
 sg13g2_a22oi_1 _11494_ (.Y(_03830_),
    .B1(_03828_),
    .B2(_03829_),
    .A2(_03827_),
    .A1(_03733_));
 sg13g2_mux2_1 _11495_ (.A0(_03825_),
    .A1(_03826_),
    .S(_03830_),
    .X(_03831_));
 sg13g2_a221oi_1 _11496_ (.B2(_03824_),
    .C1(_03831_),
    .B1(net82),
    .A1(_03823_),
    .Y(_00316_),
    .A2(net76));
 sg13g2_buf_1 _11497_ (.A(\clock_inst.min_tile.e0[18] ),
    .X(_03832_));
 sg13g2_nand3_1 _11498_ (.B(_02345_),
    .C(net102),
    .A(_03832_),
    .Y(_03833_));
 sg13g2_o21ai_1 _11499_ (.B1(_03833_),
    .Y(_03834_),
    .A1(_02345_),
    .A2(net50));
 sg13g2_a21oi_1 _11500_ (.A1(_02345_),
    .A2(net155),
    .Y(_03835_),
    .B1(_03832_));
 sg13g2_a21oi_1 _11501_ (.A1(net103),
    .A2(_03834_),
    .Y(_00317_),
    .B1(_03835_));
 sg13g2_buf_1 _11502_ (.A(\clock_inst.min_tile.e0[19] ),
    .X(_03836_));
 sg13g2_inv_1 _11503_ (.Y(_03837_),
    .A(_03836_));
 sg13g2_nand2_1 _11504_ (.Y(_03838_),
    .A(_03832_),
    .B(_02345_));
 sg13g2_xnor2_1 _11505_ (.Y(_03839_),
    .A(_02886_),
    .B(_03836_));
 sg13g2_xnor2_1 _11506_ (.Y(_03840_),
    .A(_03838_),
    .B(_03839_));
 sg13g2_nand2_1 _11507_ (.Y(_03841_),
    .A(\clock_inst.min_c[19] ),
    .B(net85));
 sg13g2_o21ai_1 _11508_ (.B1(_03841_),
    .Y(_03842_),
    .A1(net86),
    .A2(_03840_));
 sg13g2_nor2_1 _11509_ (.A(net148),
    .B(_03842_),
    .Y(_03843_));
 sg13g2_a21oi_1 _11510_ (.A1(_03837_),
    .A2(net81),
    .Y(_00318_),
    .B1(_03843_));
 sg13g2_inv_1 _11511_ (.Y(_03844_),
    .A(_03685_));
 sg13g2_buf_1 _11512_ (.A(net242),
    .X(_03845_));
 sg13g2_nand2_1 _11513_ (.Y(_03846_),
    .A(_02855_),
    .B(_03663_));
 sg13g2_xnor2_1 _11514_ (.Y(_03847_),
    .A(_02901_),
    .B(_03685_));
 sg13g2_xnor2_1 _11515_ (.Y(_03848_),
    .A(_03846_),
    .B(_03847_));
 sg13g2_nand2_1 _11516_ (.Y(_03849_),
    .A(\clock_inst.min_c[1] ),
    .B(net85));
 sg13g2_o21ai_1 _11517_ (.B1(_03849_),
    .Y(_03850_),
    .A1(net86),
    .A2(_03848_));
 sg13g2_nor2_1 _11518_ (.A(net127),
    .B(_03850_),
    .Y(_03851_));
 sg13g2_a21oi_1 _11519_ (.A1(_03844_),
    .A2(_01654_),
    .Y(_00319_),
    .B1(_03851_));
 sg13g2_buf_2 _11520_ (.A(\clock_inst.min_tile.e0[20] ),
    .X(_03852_));
 sg13g2_nand2_1 _11521_ (.Y(_03853_),
    .A(_02886_),
    .B(_03836_));
 sg13g2_nor2_1 _11522_ (.A(_02886_),
    .B(_03836_),
    .Y(_03854_));
 sg13g2_a21oi_2 _11523_ (.B1(_03854_),
    .Y(_03855_),
    .A2(_03853_),
    .A1(_03838_));
 sg13g2_xor2_1 _11524_ (.B(_03855_),
    .A(_02903_),
    .X(_03856_));
 sg13g2_nand2_1 _11525_ (.Y(_03857_),
    .A(net23),
    .B(_03856_));
 sg13g2_o21ai_1 _11526_ (.B1(net236),
    .Y(_03858_),
    .A1(net96),
    .A2(_03856_));
 sg13g2_nand2_1 _11527_ (.Y(_03859_),
    .A(_03852_),
    .B(_03858_));
 sg13g2_o21ai_1 _11528_ (.B1(_03859_),
    .Y(_00320_),
    .A1(_03852_),
    .A2(_03857_));
 sg13g2_buf_1 _11529_ (.A(\clock_inst.min_tile.e0[21] ),
    .X(_03860_));
 sg13g2_inv_1 _11530_ (.Y(_03861_),
    .A(_03860_));
 sg13g2_or2_1 _11531_ (.X(_03862_),
    .B(_03852_),
    .A(_02903_));
 sg13g2_and2_1 _11532_ (.A(_02903_),
    .B(_03852_),
    .X(_03863_));
 sg13g2_a21oi_1 _11533_ (.A1(_03855_),
    .A2(_03862_),
    .Y(_03864_),
    .B1(_03863_));
 sg13g2_xnor2_1 _11534_ (.Y(_03865_),
    .A(_02922_),
    .B(_03860_));
 sg13g2_xnor2_1 _11535_ (.Y(_03866_),
    .A(_03864_),
    .B(_03865_));
 sg13g2_nor2_1 _11536_ (.A(\clock_inst.min_c[21] ),
    .B(net232),
    .Y(_03867_));
 sg13g2_a21oi_1 _11537_ (.A1(_01519_),
    .A2(_03866_),
    .Y(_03868_),
    .B1(_03867_));
 sg13g2_nor2_1 _11538_ (.A(net127),
    .B(_03868_),
    .Y(_03869_));
 sg13g2_a21oi_1 _11539_ (.A1(_03861_),
    .A2(net81),
    .Y(_00321_),
    .B1(_03869_));
 sg13g2_inv_1 _11540_ (.Y(_03870_),
    .A(\clock_inst.min_tile.e0[22] ));
 sg13g2_nor2_1 _11541_ (.A(_02922_),
    .B(_03860_),
    .Y(_03871_));
 sg13g2_a221oi_1 _11542_ (.B2(_03862_),
    .C1(_03863_),
    .B1(_03855_),
    .A1(_02922_),
    .Y(_03872_),
    .A2(_03860_));
 sg13g2_nor2_1 _11543_ (.A(_03871_),
    .B(_03872_),
    .Y(_03873_));
 sg13g2_xor2_1 _11544_ (.B(\clock_inst.min_tile.e0[22] ),
    .A(_02924_),
    .X(_03874_));
 sg13g2_xnor2_1 _11545_ (.Y(_03875_),
    .A(_03873_),
    .B(_03874_));
 sg13g2_nor2_1 _11546_ (.A(\clock_inst.min_c[22] ),
    .B(net232),
    .Y(_03876_));
 sg13g2_a21oi_1 _11547_ (.A1(net84),
    .A2(_03875_),
    .Y(_03877_),
    .B1(_03876_));
 sg13g2_nor2_1 _11548_ (.A(net127),
    .B(_03877_),
    .Y(_03878_));
 sg13g2_a21oi_1 _11549_ (.A1(_03870_),
    .A2(net81),
    .Y(_00322_),
    .B1(_03878_));
 sg13g2_buf_1 _11550_ (.A(\clock_inst.min_tile.e0[23] ),
    .X(_03879_));
 sg13g2_inv_1 _11551_ (.Y(_03880_),
    .A(_03879_));
 sg13g2_o21ai_1 _11552_ (.B1(_03870_),
    .Y(_03881_),
    .A1(_03871_),
    .A2(_03872_));
 sg13g2_nor3_1 _11553_ (.A(_03870_),
    .B(_03871_),
    .C(_03872_),
    .Y(_03882_));
 sg13g2_a21oi_1 _11554_ (.A1(_02924_),
    .A2(_03881_),
    .Y(_03883_),
    .B1(_03882_));
 sg13g2_xnor2_1 _11555_ (.Y(_03884_),
    .A(_02935_),
    .B(_03879_));
 sg13g2_xnor2_1 _11556_ (.Y(_03885_),
    .A(_03883_),
    .B(_03884_));
 sg13g2_nor2_1 _11557_ (.A(\clock_inst.min_c[23] ),
    .B(net232),
    .Y(_03886_));
 sg13g2_a21oi_1 _11558_ (.A1(net84),
    .A2(_03885_),
    .Y(_03887_),
    .B1(_03886_));
 sg13g2_nor2_1 _11559_ (.A(_03845_),
    .B(_03887_),
    .Y(_03888_));
 sg13g2_a21oi_1 _11560_ (.A1(_03880_),
    .A2(net81),
    .Y(_00323_),
    .B1(_03888_));
 sg13g2_buf_2 _11561_ (.A(\clock_inst.min_tile.e0[24] ),
    .X(_03889_));
 sg13g2_inv_1 _11562_ (.Y(_03890_),
    .A(_03889_));
 sg13g2_nor2_1 _11563_ (.A(_02935_),
    .B(_03879_),
    .Y(_03891_));
 sg13g2_buf_1 _11564_ (.A(_03891_),
    .X(_03892_));
 sg13g2_a221oi_1 _11565_ (.B2(_02924_),
    .C1(_03882_),
    .B1(_03881_),
    .A1(_02935_),
    .Y(_03893_),
    .A2(_03879_));
 sg13g2_buf_8 _11566_ (.A(_03893_),
    .X(_03894_));
 sg13g2_or2_1 _11567_ (.X(_03895_),
    .B(net126),
    .A(net477));
 sg13g2_buf_2 _11568_ (.A(_03895_),
    .X(_03896_));
 sg13g2_nand2_1 _11569_ (.Y(_03897_),
    .A(_02959_),
    .B(_03889_));
 sg13g2_nand2_1 _11570_ (.Y(_03898_),
    .A(net566),
    .B(_03890_));
 sg13g2_nand2_1 _11571_ (.Y(_03899_),
    .A(_03897_),
    .B(_03898_));
 sg13g2_xnor2_1 _11572_ (.Y(_03900_),
    .A(_03896_),
    .B(_03899_));
 sg13g2_mux2_1 _11573_ (.A0(\clock_inst.min_c[24] ),
    .A1(_03900_),
    .S(net157),
    .X(_03901_));
 sg13g2_nor2_1 _11574_ (.A(_03845_),
    .B(_03901_),
    .Y(_03902_));
 sg13g2_a21oi_1 _11575_ (.A1(_03890_),
    .A2(net81),
    .Y(_00324_),
    .B1(_03902_));
 sg13g2_buf_2 _11576_ (.A(\clock_inst.min_tile.e0[25] ),
    .X(_03903_));
 sg13g2_inv_1 _11577_ (.Y(_03904_),
    .A(_03903_));
 sg13g2_nand2_1 _11578_ (.Y(_03905_),
    .A(_03903_),
    .B(net151));
 sg13g2_nand2_1 _11579_ (.Y(_03906_),
    .A(_03904_),
    .B(net151));
 sg13g2_mux2_1 _11580_ (.A0(_03897_),
    .A1(_03898_),
    .S(_03896_),
    .X(_03907_));
 sg13g2_mux2_1 _11581_ (.A0(_03905_),
    .A1(_03906_),
    .S(_03907_),
    .X(_03908_));
 sg13g2_nand2b_1 _11582_ (.Y(_03909_),
    .B(net97),
    .A_N(\clock_inst.min_c[25] ));
 sg13g2_a21oi_1 _11583_ (.A1(_03908_),
    .A2(_03909_),
    .Y(_03910_),
    .B1(net147));
 sg13g2_a21oi_1 _11584_ (.A1(_03904_),
    .A2(net81),
    .Y(_00325_),
    .B1(_03910_));
 sg13g2_buf_2 _11585_ (.A(\clock_inst.min_tile.e0[26] ),
    .X(_03911_));
 sg13g2_nor3_1 _11586_ (.A(_02959_),
    .B(_03889_),
    .C(_03903_),
    .Y(_03912_));
 sg13g2_nor2_1 _11587_ (.A(_03904_),
    .B(_03897_),
    .Y(_03913_));
 sg13g2_nor2_1 _11588_ (.A(net477),
    .B(net126),
    .Y(_03914_));
 sg13g2_mux2_1 _11589_ (.A0(_03912_),
    .A1(_03913_),
    .S(_03914_),
    .X(_03915_));
 sg13g2_nand3_1 _11590_ (.B(_01460_),
    .C(_03915_),
    .A(_03911_),
    .Y(_03916_));
 sg13g2_o21ai_1 _11591_ (.B1(_03916_),
    .Y(_03917_),
    .A1(\clock_inst.min_c[26] ),
    .A2(_01213_));
 sg13g2_buf_1 _11592_ (.A(_01380_),
    .X(_03918_));
 sg13g2_o21ai_1 _11593_ (.B1(_03918_),
    .Y(_03919_),
    .A1(_01471_),
    .A2(_03915_));
 sg13g2_inv_1 _11594_ (.Y(_03920_),
    .A(_03911_));
 sg13g2_a22oi_1 _11595_ (.Y(_00326_),
    .B1(_03919_),
    .B2(_03920_),
    .A2(_03917_),
    .A1(_01458_));
 sg13g2_buf_2 _11596_ (.A(\clock_inst.min_tile.e0[27] ),
    .X(_03921_));
 sg13g2_nor2_1 _11597_ (.A(_03903_),
    .B(_03911_),
    .Y(_03922_));
 sg13g2_o21ai_1 _11598_ (.B1(_03922_),
    .Y(_03923_),
    .A1(net477),
    .A2(net126));
 sg13g2_nand2_1 _11599_ (.Y(_03924_),
    .A(_03903_),
    .B(_03911_));
 sg13g2_or4_1 _11600_ (.A(net477),
    .B(net126),
    .C(_03897_),
    .D(_03924_),
    .X(_03925_));
 sg13g2_o21ai_1 _11601_ (.B1(_03925_),
    .Y(_03926_),
    .A1(_03898_),
    .A2(_03923_));
 sg13g2_xnor2_1 _11602_ (.Y(_03927_),
    .A(_03921_),
    .B(_03926_));
 sg13g2_nand2_1 _11603_ (.Y(_03928_),
    .A(\clock_inst.min_c[27] ),
    .B(net90));
 sg13g2_o21ai_1 _11604_ (.B1(_03928_),
    .Y(_03929_),
    .A1(net98),
    .A2(_03927_));
 sg13g2_mux2_1 _11605_ (.A0(_03921_),
    .A1(_03929_),
    .S(net146),
    .X(_00327_));
 sg13g2_buf_1 _11606_ (.A(\clock_inst.min_tile.e0[28] ),
    .X(_03930_));
 sg13g2_nor2_1 _11607_ (.A(_03930_),
    .B(_01136_),
    .Y(_03931_));
 sg13g2_o21ai_1 _11608_ (.B1(net566),
    .Y(_03932_),
    .A1(_03921_),
    .A2(_03923_));
 sg13g2_nand3_1 _11609_ (.B(_03911_),
    .C(_03921_),
    .A(_03903_),
    .Y(_03933_));
 sg13g2_nor3_1 _11610_ (.A(net477),
    .B(net126),
    .C(_03933_),
    .Y(_03934_));
 sg13g2_o21ai_1 _11611_ (.B1(_03889_),
    .Y(_03935_),
    .A1(net566),
    .A2(_03934_));
 sg13g2_nand2_1 _11612_ (.Y(_03936_),
    .A(_03932_),
    .B(_03935_));
 sg13g2_xor2_1 _11613_ (.B(_03930_),
    .A(net566),
    .X(_03937_));
 sg13g2_and3_1 _11614_ (.X(_03938_),
    .A(net23),
    .B(_03936_),
    .C(_03937_));
 sg13g2_nor3_1 _11615_ (.A(net95),
    .B(_03936_),
    .C(_03937_),
    .Y(_03939_));
 sg13g2_nor3_1 _11616_ (.A(\clock_inst.min_c[28] ),
    .B(net143),
    .C(net87),
    .Y(_03940_));
 sg13g2_nor4_1 _11617_ (.A(_03931_),
    .B(_03938_),
    .C(_03939_),
    .D(_03940_),
    .Y(_00328_));
 sg13g2_inv_1 _11618_ (.Y(_03941_),
    .A(\clock_inst.min_tile.e0[29] ));
 sg13g2_nor2_1 _11619_ (.A(_03941_),
    .B(net158),
    .Y(_03942_));
 sg13g2_nor2_1 _11620_ (.A(\clock_inst.min_tile.e0[29] ),
    .B(net158),
    .Y(_03943_));
 sg13g2_or3_1 _11621_ (.A(_03921_),
    .B(_03930_),
    .C(_03898_),
    .X(_03944_));
 sg13g2_nor2_1 _11622_ (.A(net566),
    .B(_03890_),
    .Y(_03945_));
 sg13g2_nand2_1 _11623_ (.Y(_03946_),
    .A(_03930_),
    .B(_03945_));
 sg13g2_or4_1 _11624_ (.A(net477),
    .B(net126),
    .C(_03933_),
    .D(_03946_),
    .X(_03947_));
 sg13g2_o21ai_1 _11625_ (.B1(_03947_),
    .Y(_03948_),
    .A1(_03923_),
    .A2(_03944_));
 sg13g2_mux2_1 _11626_ (.A0(_03942_),
    .A1(_03943_),
    .S(_03948_),
    .X(_03949_));
 sg13g2_nor2_1 _11627_ (.A(_03354_),
    .B(net101),
    .Y(_03950_));
 sg13g2_nor3_1 _11628_ (.A(_01152_),
    .B(_03949_),
    .C(_03950_),
    .Y(_03951_));
 sg13g2_a21oi_1 _11629_ (.A1(_03941_),
    .A2(net81),
    .Y(_00329_),
    .B1(_03951_));
 sg13g2_inv_1 _11630_ (.Y(_03952_),
    .A(_03692_));
 sg13g2_buf_1 _11631_ (.A(net161),
    .X(_03953_));
 sg13g2_xor2_1 _11632_ (.B(_03692_),
    .A(_02943_),
    .X(_03954_));
 sg13g2_xnor2_1 _11633_ (.Y(_03955_),
    .A(_03689_),
    .B(_03954_));
 sg13g2_nand2_1 _11634_ (.Y(_03956_),
    .A(net157),
    .B(_03955_));
 sg13g2_o21ai_1 _11635_ (.B1(_03956_),
    .Y(_03957_),
    .A1(_03368_),
    .A2(net101));
 sg13g2_nor2_1 _11636_ (.A(net127),
    .B(_03957_),
    .Y(_03958_));
 sg13g2_a21oi_1 _11637_ (.A1(_03952_),
    .A2(net68),
    .Y(_00330_),
    .B1(_03958_));
 sg13g2_buf_1 _11638_ (.A(\clock_inst.min_tile.e0[30] ),
    .X(_03959_));
 sg13g2_nor4_1 _11639_ (.A(_03911_),
    .B(_03921_),
    .C(_03930_),
    .D(\clock_inst.min_tile.e0[29] ),
    .Y(_03960_));
 sg13g2_nand4_1 _11640_ (.B(_03890_),
    .C(_03904_),
    .A(_02958_),
    .Y(_03961_),
    .D(_03960_));
 sg13g2_buf_1 _11641_ (.A(_03961_),
    .X(_03962_));
 sg13g2_inv_1 _11642_ (.Y(_03963_),
    .A(_03962_));
 sg13g2_o21ai_1 _11643_ (.B1(_03963_),
    .Y(_03964_),
    .A1(net477),
    .A2(net126));
 sg13g2_nand3_1 _11644_ (.B(_03930_),
    .C(\clock_inst.min_tile.e0[29] ),
    .A(_03921_),
    .Y(_03965_));
 sg13g2_nor2_1 _11645_ (.A(_03924_),
    .B(_03965_),
    .Y(_03966_));
 sg13g2_nand2_1 _11646_ (.Y(_03967_),
    .A(_03945_),
    .B(_03966_));
 sg13g2_or3_1 _11647_ (.A(net477),
    .B(net126),
    .C(_03967_),
    .X(_03968_));
 sg13g2_nand2_1 _11648_ (.Y(_03969_),
    .A(_03964_),
    .B(_03968_));
 sg13g2_nand3_1 _11649_ (.B(net87),
    .C(_03969_),
    .A(_03959_),
    .Y(_03970_));
 sg13g2_o21ai_1 _11650_ (.B1(_03970_),
    .Y(_03971_),
    .A1(\clock_inst.min_c[30] ),
    .A2(net50));
 sg13g2_o21ai_1 _11651_ (.B1(_03918_),
    .Y(_03972_),
    .A1(net47),
    .A2(_03969_));
 sg13g2_inv_1 _11652_ (.Y(_03973_),
    .A(_03959_));
 sg13g2_a22oi_1 _11653_ (.Y(_00331_),
    .B1(_03972_),
    .B2(_03973_),
    .A2(_03971_),
    .A1(_01137_));
 sg13g2_buf_1 _11654_ (.A(\clock_inst.min_tile.e0[31] ),
    .X(_03974_));
 sg13g2_inv_1 _11655_ (.Y(_03975_),
    .A(_03974_));
 sg13g2_nand2_1 _11656_ (.Y(_03976_),
    .A(_03974_),
    .B(net151));
 sg13g2_nand2_1 _11657_ (.Y(_03977_),
    .A(_03975_),
    .B(net151));
 sg13g2_mux2_1 _11658_ (.A0(_03964_),
    .A1(_03968_),
    .S(_03959_),
    .X(_03978_));
 sg13g2_mux2_1 _11659_ (.A0(_03976_),
    .A1(_03977_),
    .S(_03978_),
    .X(_03979_));
 sg13g2_nand2_1 _11660_ (.Y(_03980_),
    .A(_03397_),
    .B(net97));
 sg13g2_a21oi_1 _11661_ (.A1(_03979_),
    .A2(_03980_),
    .Y(_03981_),
    .B1(net140));
 sg13g2_a21oi_1 _11662_ (.A1(_03975_),
    .A2(_03953_),
    .Y(_00332_),
    .B1(_03981_));
 sg13g2_buf_2 _11663_ (.A(\clock_inst.min_tile.e0[32] ),
    .X(_03982_));
 sg13g2_nor3_1 _11664_ (.A(_03959_),
    .B(_03974_),
    .C(_03962_),
    .Y(_03983_));
 sg13g2_nor4_1 _11665_ (.A(_03973_),
    .B(_03975_),
    .C(_03924_),
    .D(_03965_),
    .Y(_03984_));
 sg13g2_and2_1 _11666_ (.A(_03945_),
    .B(_03984_),
    .X(_03985_));
 sg13g2_mux2_1 _11667_ (.A0(_03983_),
    .A1(_03985_),
    .S(_03914_),
    .X(_03986_));
 sg13g2_xnor2_1 _11668_ (.Y(_03987_),
    .A(_03982_),
    .B(_03986_));
 sg13g2_nand2_1 _11669_ (.Y(_03988_),
    .A(\clock_inst.min_c[32] ),
    .B(net90));
 sg13g2_o21ai_1 _11670_ (.B1(_03988_),
    .Y(_03989_),
    .A1(net98),
    .A2(_03987_));
 sg13g2_mux2_1 _11671_ (.A0(_03982_),
    .A1(_03989_),
    .S(net146),
    .X(_00333_));
 sg13g2_buf_1 _11672_ (.A(\clock_inst.min_tile.e0[33] ),
    .X(_03990_));
 sg13g2_and2_1 _11673_ (.A(_03990_),
    .B(net99),
    .X(_03991_));
 sg13g2_nor2_1 _11674_ (.A(_03990_),
    .B(_01274_),
    .Y(_03992_));
 sg13g2_nand2_1 _11675_ (.Y(_03993_),
    .A(_03982_),
    .B(_03985_));
 sg13g2_nor4_1 _11676_ (.A(_03959_),
    .B(_03974_),
    .C(_03982_),
    .D(_03962_),
    .Y(_03994_));
 sg13g2_o21ai_1 _11677_ (.B1(_03994_),
    .Y(_03995_),
    .A1(_03892_),
    .A2(_03894_));
 sg13g2_o21ai_1 _11678_ (.B1(_03995_),
    .Y(_03996_),
    .A1(_03896_),
    .A2(_03993_));
 sg13g2_mux2_1 _11679_ (.A0(_03991_),
    .A1(_03992_),
    .S(_03996_),
    .X(_03997_));
 sg13g2_and2_1 _11680_ (.A(\clock_inst.min_c[33] ),
    .B(_01610_),
    .X(_03998_));
 sg13g2_buf_1 _11681_ (.A(_03998_),
    .X(_03999_));
 sg13g2_a21oi_1 _11682_ (.A1(_03990_),
    .A2(_01409_),
    .Y(_04000_),
    .B1(_03999_));
 sg13g2_nand2b_1 _11683_ (.Y(_00334_),
    .B(_04000_),
    .A_N(_03997_));
 sg13g2_buf_1 _11684_ (.A(\clock_inst.min_tile.e0[34] ),
    .X(_04001_));
 sg13g2_inv_1 _11685_ (.Y(_04002_),
    .A(_04001_));
 sg13g2_nand2_1 _11686_ (.Y(_04003_),
    .A(_03982_),
    .B(_03990_));
 sg13g2_nor3_1 _11687_ (.A(_03973_),
    .B(_03975_),
    .C(_04003_),
    .Y(_04004_));
 sg13g2_nand4_1 _11688_ (.B(_03889_),
    .C(_03966_),
    .A(_02959_),
    .Y(_04005_),
    .D(_04004_));
 sg13g2_nor4_1 _11689_ (.A(_03959_),
    .B(_03974_),
    .C(_03982_),
    .D(_03990_),
    .Y(_04006_));
 sg13g2_nor2b_1 _11690_ (.A(_03962_),
    .B_N(_04006_),
    .Y(_04007_));
 sg13g2_o21ai_1 _11691_ (.B1(_04007_),
    .Y(_04008_),
    .A1(_03892_),
    .A2(_03894_));
 sg13g2_o21ai_1 _11692_ (.B1(_04008_),
    .Y(_04009_),
    .A1(_03896_),
    .A2(_04005_));
 sg13g2_xnor2_1 _11693_ (.Y(_04010_),
    .A(_04002_),
    .B(_04009_));
 sg13g2_a21oi_1 _11694_ (.A1(net23),
    .A2(_04010_),
    .Y(_04011_),
    .B1(_03999_));
 sg13g2_o21ai_1 _11695_ (.B1(_04011_),
    .Y(_00335_),
    .A1(_04002_),
    .A2(_01166_));
 sg13g2_buf_1 _11696_ (.A(\clock_inst.min_tile.e0[35] ),
    .X(_04012_));
 sg13g2_nor3_1 _11697_ (.A(_03982_),
    .B(_03990_),
    .C(_04001_),
    .Y(_04013_));
 sg13g2_nand2_1 _11698_ (.Y(_04014_),
    .A(_03983_),
    .B(_04013_));
 sg13g2_and4_1 _11699_ (.A(_04012_),
    .B(net99),
    .C(_03896_),
    .D(_04014_),
    .X(_04015_));
 sg13g2_nor4_1 _11700_ (.A(_04012_),
    .B(_01274_),
    .C(_03914_),
    .D(_04014_),
    .Y(_04016_));
 sg13g2_nor2_1 _11701_ (.A(net566),
    .B(_04003_),
    .Y(_04017_));
 sg13g2_nand4_1 _11702_ (.B(_04001_),
    .C(_03984_),
    .A(_03889_),
    .Y(_04018_),
    .D(_04017_));
 sg13g2_nand3_1 _11703_ (.B(net99),
    .C(_04018_),
    .A(_04012_),
    .Y(_04019_));
 sg13g2_or3_1 _11704_ (.A(_04012_),
    .B(_01274_),
    .C(_04018_),
    .X(_04020_));
 sg13g2_a21oi_1 _11705_ (.A1(_04019_),
    .A2(_04020_),
    .Y(_04021_),
    .B1(_03896_));
 sg13g2_or4_1 _11706_ (.A(_03999_),
    .B(_04015_),
    .C(_04016_),
    .D(_04021_),
    .X(_04022_));
 sg13g2_buf_1 _11707_ (.A(_04022_),
    .X(_04023_));
 sg13g2_a21o_1 _11708_ (.A2(_01034_),
    .A1(_04012_),
    .B1(_04023_),
    .X(_00336_));
 sg13g2_buf_1 _11709_ (.A(\clock_inst.min_tile.e0[36] ),
    .X(_04024_));
 sg13g2_inv_1 _11710_ (.Y(_04025_),
    .A(_04024_));
 sg13g2_nor2_1 _11711_ (.A(_03415_),
    .B(net235),
    .Y(_04026_));
 sg13g2_xnor2_1 _11712_ (.Y(_04027_),
    .A(_02968_),
    .B(_04024_));
 sg13g2_nor2_1 _11713_ (.A(net237),
    .B(_04027_),
    .Y(_04028_));
 sg13g2_o21ai_1 _11714_ (.B1(net156),
    .Y(_04029_),
    .A1(_04026_),
    .A2(_04028_));
 sg13g2_o21ai_1 _11715_ (.B1(_04029_),
    .Y(_00337_),
    .A1(_04025_),
    .A2(net106));
 sg13g2_buf_1 _11716_ (.A(\clock_inst.min_tile.e0[37] ),
    .X(_04030_));
 sg13g2_inv_1 _11717_ (.Y(_04031_),
    .A(_04030_));
 sg13g2_nand2_1 _11718_ (.Y(_04032_),
    .A(_02968_),
    .B(_04024_));
 sg13g2_xnor2_1 _11719_ (.Y(_04033_),
    .A(_02970_),
    .B(_04030_));
 sg13g2_xnor2_1 _11720_ (.Y(_04034_),
    .A(_04032_),
    .B(_04033_));
 sg13g2_nand2_1 _11721_ (.Y(_04035_),
    .A(\clock_inst.min_c[37] ),
    .B(net85));
 sg13g2_o21ai_1 _11722_ (.B1(_04035_),
    .Y(_04036_),
    .A1(net86),
    .A2(_04034_));
 sg13g2_nor2_1 _11723_ (.A(net127),
    .B(_04036_),
    .Y(_04037_));
 sg13g2_a21oi_1 _11724_ (.A1(_04031_),
    .A2(net68),
    .Y(_00338_),
    .B1(_04037_));
 sg13g2_buf_1 _11725_ (.A(\clock_inst.min_tile.e0[38] ),
    .X(_04038_));
 sg13g2_inv_1 _11726_ (.Y(_04039_),
    .A(_04038_));
 sg13g2_nor2_1 _11727_ (.A(_02970_),
    .B(_04030_),
    .Y(_04040_));
 sg13g2_a22oi_1 _11728_ (.Y(_04041_),
    .B1(_02970_),
    .B2(_04030_),
    .A2(_04024_),
    .A1(_02968_));
 sg13g2_nor2_1 _11729_ (.A(_04040_),
    .B(_04041_),
    .Y(_04042_));
 sg13g2_xnor2_1 _11730_ (.Y(_04043_),
    .A(_02982_),
    .B(_04038_));
 sg13g2_xnor2_1 _11731_ (.Y(_04044_),
    .A(_04042_),
    .B(_04043_));
 sg13g2_nor2_1 _11732_ (.A(net141),
    .B(_04044_),
    .Y(_04045_));
 sg13g2_a21oi_1 _11733_ (.A1(_03428_),
    .A2(net97),
    .Y(_04046_),
    .B1(_04045_));
 sg13g2_nor2_1 _11734_ (.A(net127),
    .B(_04046_),
    .Y(_04047_));
 sg13g2_a21oi_1 _11735_ (.A1(_04039_),
    .A2(net68),
    .Y(_00339_),
    .B1(_04047_));
 sg13g2_inv_1 _11736_ (.Y(_04048_),
    .A(\clock_inst.min_tile.e0[39] ));
 sg13g2_nor2_1 _11737_ (.A(_02983_),
    .B(_04039_),
    .Y(_04049_));
 sg13g2_nor2_1 _11738_ (.A(_02982_),
    .B(_04038_),
    .Y(_04050_));
 sg13g2_nor3_1 _11739_ (.A(_04040_),
    .B(_04041_),
    .C(_04050_),
    .Y(_04051_));
 sg13g2_nor2_1 _11740_ (.A(_04049_),
    .B(_04051_),
    .Y(_04052_));
 sg13g2_xnor2_1 _11741_ (.Y(_04053_),
    .A(_03010_),
    .B(\clock_inst.min_tile.e0[39] ));
 sg13g2_xnor2_1 _11742_ (.Y(_04054_),
    .A(_04052_),
    .B(_04053_));
 sg13g2_nor2_1 _11743_ (.A(\clock_inst.min_c[39] ),
    .B(net232),
    .Y(_04055_));
 sg13g2_a21oi_1 _11744_ (.A1(net84),
    .A2(_04054_),
    .Y(_04056_),
    .B1(_04055_));
 sg13g2_nor2_1 _11745_ (.A(net127),
    .B(_04056_),
    .Y(_04057_));
 sg13g2_a21oi_1 _11746_ (.A1(_04048_),
    .A2(net68),
    .Y(_00340_),
    .B1(_04057_));
 sg13g2_nand2_1 _11747_ (.Y(_04058_),
    .A(_03698_),
    .B(_03778_));
 sg13g2_xnor2_1 _11748_ (.Y(_04059_),
    .A(_03012_),
    .B(_03690_));
 sg13g2_xnor2_1 _11749_ (.Y(_04060_),
    .A(_04058_),
    .B(_04059_));
 sg13g2_nand2_1 _11750_ (.Y(_04061_),
    .A(\clock_inst.min_c[3] ),
    .B(net85));
 sg13g2_o21ai_1 _11751_ (.B1(_04061_),
    .Y(_04062_),
    .A1(net86),
    .A2(_04060_));
 sg13g2_nor2_1 _11752_ (.A(net127),
    .B(_04062_),
    .Y(_04063_));
 sg13g2_a21oi_1 _11753_ (.A1(_03691_),
    .A2(net68),
    .Y(_00341_),
    .B1(_04063_));
 sg13g2_buf_1 _11754_ (.A(\clock_inst.min_tile.e0[40] ),
    .X(_04064_));
 sg13g2_inv_1 _11755_ (.Y(_04065_),
    .A(_04064_));
 sg13g2_buf_1 _11756_ (.A(net244),
    .X(_04066_));
 sg13g2_inv_1 _11757_ (.Y(_04067_),
    .A(_03010_));
 sg13g2_nand2_1 _11758_ (.Y(_04068_),
    .A(_04067_),
    .B(_04048_));
 sg13g2_o21ai_1 _11759_ (.B1(_04068_),
    .Y(_04069_),
    .A1(_04049_),
    .A2(_04051_));
 sg13g2_nand2_1 _11760_ (.Y(_04070_),
    .A(_03010_),
    .B(\clock_inst.min_tile.e0[39] ));
 sg13g2_nand2_1 _11761_ (.Y(_04071_),
    .A(_04069_),
    .B(_04070_));
 sg13g2_xor2_1 _11762_ (.B(_04064_),
    .A(_03024_),
    .X(_04072_));
 sg13g2_xnor2_1 _11763_ (.Y(_04073_),
    .A(_04071_),
    .B(_04072_));
 sg13g2_nor2_1 _11764_ (.A(\clock_inst.min_c[40] ),
    .B(net232),
    .Y(_04074_));
 sg13g2_a21oi_1 _11765_ (.A1(net84),
    .A2(_04073_),
    .Y(_04075_),
    .B1(_04074_));
 sg13g2_nor2_1 _11766_ (.A(net124),
    .B(_04075_),
    .Y(_04076_));
 sg13g2_a21oi_1 _11767_ (.A1(_04065_),
    .A2(net68),
    .Y(_00342_),
    .B1(_04076_));
 sg13g2_buf_1 _11768_ (.A(\clock_inst.min_tile.e0[41] ),
    .X(_04077_));
 sg13g2_inv_1 _11769_ (.Y(_04078_),
    .A(_04077_));
 sg13g2_xor2_1 _11770_ (.B(_04077_),
    .A(_03038_),
    .X(_04079_));
 sg13g2_nor2_1 _11771_ (.A(_03024_),
    .B(_04064_),
    .Y(_04080_));
 sg13g2_nor3_1 _11772_ (.A(_04048_),
    .B(_04050_),
    .C(_04080_),
    .Y(_04081_));
 sg13g2_nand2_1 _11773_ (.Y(_04082_),
    .A(_02982_),
    .B(_04038_));
 sg13g2_a221oi_1 _11774_ (.B2(_04065_),
    .C1(_04082_),
    .B1(_03025_),
    .A1(_04067_),
    .Y(_04083_),
    .A2(_04048_));
 sg13g2_a21o_1 _11775_ (.A2(_04081_),
    .A1(_04042_),
    .B1(_04083_),
    .X(_04084_));
 sg13g2_buf_2 _11776_ (.A(_04084_),
    .X(_04085_));
 sg13g2_nor3_1 _11777_ (.A(_04067_),
    .B(_04050_),
    .C(_04080_),
    .Y(_04086_));
 sg13g2_nor2_1 _11778_ (.A(_04070_),
    .B(_04080_),
    .Y(_04087_));
 sg13g2_a21o_1 _11779_ (.A2(_04086_),
    .A1(_04042_),
    .B1(_04087_),
    .X(_04088_));
 sg13g2_buf_2 _11780_ (.A(_04088_),
    .X(_04089_));
 sg13g2_nor2_1 _11781_ (.A(_04085_),
    .B(_04089_),
    .Y(_04090_));
 sg13g2_o21ai_1 _11782_ (.B1(_04090_),
    .Y(_04091_),
    .A1(_03025_),
    .A2(_04065_));
 sg13g2_xnor2_1 _11783_ (.Y(_04092_),
    .A(_04079_),
    .B(_04091_));
 sg13g2_nor2_1 _11784_ (.A(\clock_inst.min_c[41] ),
    .B(net232),
    .Y(_04093_));
 sg13g2_a21oi_1 _11785_ (.A1(net84),
    .A2(_04092_),
    .Y(_04094_),
    .B1(_04093_));
 sg13g2_nor2_1 _11786_ (.A(net124),
    .B(_04094_),
    .Y(_04095_));
 sg13g2_a21oi_1 _11787_ (.A1(_04078_),
    .A2(net68),
    .Y(_00343_),
    .B1(_04095_));
 sg13g2_buf_1 _11788_ (.A(\clock_inst.min_tile.e0[42] ),
    .X(_04096_));
 sg13g2_inv_1 _11789_ (.Y(_04097_),
    .A(_04096_));
 sg13g2_a22oi_1 _11790_ (.Y(_04098_),
    .B1(_03038_),
    .B2(_04077_),
    .A2(_04064_),
    .A1(_03024_));
 sg13g2_nor2_1 _11791_ (.A(_03038_),
    .B(_04077_),
    .Y(_04099_));
 sg13g2_a21oi_1 _11792_ (.A1(_04090_),
    .A2(_04098_),
    .Y(_04100_),
    .B1(_04099_));
 sg13g2_xor2_1 _11793_ (.B(_04096_),
    .A(_03053_),
    .X(_04101_));
 sg13g2_xnor2_1 _11794_ (.Y(_04102_),
    .A(_04100_),
    .B(_04101_));
 sg13g2_nor2_1 _11795_ (.A(\clock_inst.min_c[42] ),
    .B(net232),
    .Y(_04103_));
 sg13g2_a21oi_1 _11796_ (.A1(net84),
    .A2(_04102_),
    .Y(_04104_),
    .B1(_04103_));
 sg13g2_nor2_1 _11797_ (.A(net124),
    .B(_04104_),
    .Y(_04105_));
 sg13g2_a21oi_1 _11798_ (.A1(_04097_),
    .A2(_03953_),
    .Y(_00344_),
    .B1(_04105_));
 sg13g2_buf_2 _11799_ (.A(\clock_inst.min_tile.e0[43] ),
    .X(_04106_));
 sg13g2_inv_1 _11800_ (.Y(_04107_),
    .A(_04106_));
 sg13g2_nor2_1 _11801_ (.A(_03053_),
    .B(_04096_),
    .Y(_04108_));
 sg13g2_inv_1 _11802_ (.Y(_04109_),
    .A(_04108_));
 sg13g2_nand2_1 _11803_ (.Y(_04110_),
    .A(_03053_),
    .B(_04096_));
 sg13g2_o21ai_1 _11804_ (.B1(_04110_),
    .Y(_04111_),
    .A1(_04099_),
    .A2(_04098_));
 sg13g2_and2_1 _11805_ (.A(_04109_),
    .B(_04111_),
    .X(_04112_));
 sg13g2_buf_2 _11806_ (.A(_04112_),
    .X(_04113_));
 sg13g2_or2_1 _11807_ (.X(_04114_),
    .B(_04077_),
    .A(_03038_));
 sg13g2_nand2_1 _11808_ (.Y(_04115_),
    .A(_04114_),
    .B(_04109_));
 sg13g2_a221oi_1 _11809_ (.B2(_04070_),
    .C1(_04115_),
    .B1(_04069_),
    .A1(_03025_),
    .Y(_04116_),
    .A2(_04065_));
 sg13g2_nor2_1 _11810_ (.A(_04113_),
    .B(_04116_),
    .Y(_04117_));
 sg13g2_xor2_1 _11811_ (.B(_04106_),
    .A(_03066_),
    .X(_04118_));
 sg13g2_xnor2_1 _11812_ (.Y(_04119_),
    .A(_04117_),
    .B(_04118_));
 sg13g2_nor2_1 _11813_ (.A(net107),
    .B(_04119_),
    .Y(_04120_));
 sg13g2_nor2_1 _11814_ (.A(\clock_inst.min_c[43] ),
    .B(net104),
    .Y(_04121_));
 sg13g2_or3_1 _11815_ (.A(net143),
    .B(_04120_),
    .C(_04121_),
    .X(_04122_));
 sg13g2_o21ai_1 _11816_ (.B1(_04122_),
    .Y(_00345_),
    .A1(_04107_),
    .A2(net106));
 sg13g2_buf_1 _11817_ (.A(\clock_inst.min_tile.e0[44] ),
    .X(_04123_));
 sg13g2_inv_1 _11818_ (.Y(_04124_),
    .A(_04123_));
 sg13g2_xor2_1 _11819_ (.B(_04123_),
    .A(_03078_),
    .X(_04125_));
 sg13g2_o21ai_1 _11820_ (.B1(_04106_),
    .Y(_04126_),
    .A1(_04113_),
    .A2(_04116_));
 sg13g2_nor3_1 _11821_ (.A(_04106_),
    .B(_04113_),
    .C(_04116_),
    .Y(_04127_));
 sg13g2_a21oi_1 _11822_ (.A1(_03067_),
    .A2(_04126_),
    .Y(_04128_),
    .B1(_04127_));
 sg13g2_xnor2_1 _11823_ (.Y(_04129_),
    .A(_04125_),
    .B(_04128_));
 sg13g2_nor2_1 _11824_ (.A(\clock_inst.min_c[44] ),
    .B(net232),
    .Y(_04130_));
 sg13g2_a21oi_1 _11825_ (.A1(net84),
    .A2(_04129_),
    .Y(_04131_),
    .B1(_04130_));
 sg13g2_nor2_1 _11826_ (.A(net124),
    .B(_04131_),
    .Y(_04132_));
 sg13g2_a21oi_1 _11827_ (.A1(_04124_),
    .A2(net68),
    .Y(_00346_),
    .B1(_04132_));
 sg13g2_inv_1 _11828_ (.Y(_04133_),
    .A(\clock_inst.min_tile.e0[45] ));
 sg13g2_buf_1 _11829_ (.A(net153),
    .X(_04134_));
 sg13g2_a22oi_1 _11830_ (.Y(_04135_),
    .B1(_03078_),
    .B2(_04123_),
    .A2(_04106_),
    .A1(_03066_));
 sg13g2_inv_1 _11831_ (.Y(_04136_),
    .A(_04135_));
 sg13g2_nor4_2 _11832_ (.A(_04085_),
    .B(_04089_),
    .C(_04113_),
    .Y(_04137_),
    .D(_04136_));
 sg13g2_nor2_1 _11833_ (.A(_03078_),
    .B(_04123_),
    .Y(_04138_));
 sg13g2_o21ai_1 _11834_ (.B1(_04110_),
    .Y(_04139_),
    .A1(_04099_),
    .A2(_04108_));
 sg13g2_a21o_1 _11835_ (.A2(_04139_),
    .A1(_04106_),
    .B1(_03066_),
    .X(_04140_));
 sg13g2_or2_1 _11836_ (.X(_04141_),
    .B(_04139_),
    .A(_04106_));
 sg13g2_nand2_1 _11837_ (.Y(_04142_),
    .A(_03078_),
    .B(_04123_));
 sg13g2_inv_1 _11838_ (.Y(_04143_),
    .A(_04142_));
 sg13g2_a21oi_1 _11839_ (.A1(_04140_),
    .A2(_04141_),
    .Y(_04144_),
    .B1(_04143_));
 sg13g2_or3_1 _11840_ (.A(_04137_),
    .B(_04138_),
    .C(_04144_),
    .X(_04145_));
 sg13g2_buf_1 _11841_ (.A(_04145_),
    .X(_04146_));
 sg13g2_nand2_2 _11842_ (.Y(_04147_),
    .A(net568),
    .B(_04133_));
 sg13g2_nand2_1 _11843_ (.Y(_04148_),
    .A(net479),
    .B(\clock_inst.min_tile.e0[45] ));
 sg13g2_nand2_1 _11844_ (.Y(_04149_),
    .A(_04147_),
    .B(_04148_));
 sg13g2_xor2_1 _11845_ (.B(_04149_),
    .A(net66),
    .X(_04150_));
 sg13g2_nand2_1 _11846_ (.Y(_04151_),
    .A(\clock_inst.min_c[45] ),
    .B(net241));
 sg13g2_o21ai_1 _11847_ (.B1(_04151_),
    .Y(_04152_),
    .A1(net158),
    .A2(_04150_));
 sg13g2_nor2_1 _11848_ (.A(net244),
    .B(_04152_),
    .Y(_04153_));
 sg13g2_a21oi_1 _11849_ (.A1(_04133_),
    .A2(net67),
    .Y(_00347_),
    .B1(_04153_));
 sg13g2_buf_1 _11850_ (.A(\clock_inst.min_tile.e0[46] ),
    .X(_04154_));
 sg13g2_inv_1 _11851_ (.Y(_04155_),
    .A(_04154_));
 sg13g2_mux2_1 _11852_ (.A0(_04148_),
    .A1(_04147_),
    .S(net66),
    .X(_04156_));
 sg13g2_xnor2_1 _11853_ (.Y(_04157_),
    .A(_04155_),
    .B(_04156_));
 sg13g2_nand2_1 _11854_ (.Y(_04158_),
    .A(\clock_inst.min_c[46] ),
    .B(net85));
 sg13g2_o21ai_1 _11855_ (.B1(_04158_),
    .Y(_04159_),
    .A1(net86),
    .A2(_04157_));
 sg13g2_nor2_1 _11856_ (.A(net124),
    .B(_04159_),
    .Y(_04160_));
 sg13g2_a21oi_1 _11857_ (.A1(_04155_),
    .A2(net67),
    .Y(_00348_),
    .B1(_04160_));
 sg13g2_buf_1 _11858_ (.A(\clock_inst.min_tile.e0[47] ),
    .X(_04161_));
 sg13g2_inv_1 _11859_ (.Y(_04162_),
    .A(_04161_));
 sg13g2_nor2_1 _11860_ (.A(net568),
    .B(_04133_),
    .Y(_04163_));
 sg13g2_nand2_1 _11861_ (.Y(_04164_),
    .A(_04154_),
    .B(_04163_));
 sg13g2_buf_1 _11862_ (.A(net568),
    .X(_04165_));
 sg13g2_nand4_1 _11863_ (.B(_04133_),
    .C(_04155_),
    .A(_04165_),
    .Y(_04166_),
    .D(net66));
 sg13g2_o21ai_1 _11864_ (.B1(_04166_),
    .Y(_04167_),
    .A1(net66),
    .A2(_04164_));
 sg13g2_xnor2_1 _11865_ (.Y(_04168_),
    .A(_04162_),
    .B(_04167_));
 sg13g2_o21ai_1 _11866_ (.B1(net240),
    .Y(_04169_),
    .A1(_03542_),
    .A2(net157));
 sg13g2_a21oi_1 _11867_ (.A1(net93),
    .A2(_04168_),
    .Y(_04170_),
    .B1(_04169_));
 sg13g2_a21oi_1 _11868_ (.A1(_04162_),
    .A2(_04134_),
    .Y(_00349_),
    .B1(_04170_));
 sg13g2_buf_1 _11869_ (.A(\clock_inst.min_tile.e0[48] ),
    .X(_04171_));
 sg13g2_nor4_1 _11870_ (.A(net568),
    .B(_04133_),
    .C(_04155_),
    .D(_04162_),
    .Y(_04172_));
 sg13g2_nor3_1 _11871_ (.A(_04154_),
    .B(_04161_),
    .C(_04147_),
    .Y(_04173_));
 sg13g2_mux2_1 _11872_ (.A0(_04172_),
    .A1(_04173_),
    .S(net66),
    .X(_04174_));
 sg13g2_nand3_1 _11873_ (.B(net87),
    .C(_04174_),
    .A(_04171_),
    .Y(_04175_));
 sg13g2_o21ai_1 _11874_ (.B1(_04175_),
    .Y(_04176_),
    .A1(\clock_inst.min_c[48] ),
    .A2(net51));
 sg13g2_o21ai_1 _11875_ (.B1(net125),
    .Y(_04177_),
    .A1(net47),
    .A2(_04174_));
 sg13g2_inv_1 _11876_ (.Y(_04178_),
    .A(_04171_));
 sg13g2_a22oi_1 _11877_ (.Y(_00350_),
    .B1(_04177_),
    .B2(_04178_),
    .A2(_04176_),
    .A1(net108));
 sg13g2_buf_1 _11878_ (.A(\clock_inst.min_tile.e0[49] ),
    .X(_04179_));
 sg13g2_and2_1 _11879_ (.A(_04171_),
    .B(_04172_),
    .X(_04180_));
 sg13g2_nor3_1 _11880_ (.A(_04154_),
    .B(_04161_),
    .C(_04171_),
    .Y(_04181_));
 sg13g2_nor2b_1 _11881_ (.A(_04147_),
    .B_N(_04181_),
    .Y(_04182_));
 sg13g2_mux2_1 _11882_ (.A0(_04180_),
    .A1(_04182_),
    .S(net66),
    .X(_04183_));
 sg13g2_nand3_1 _11883_ (.B(_01216_),
    .C(_04183_),
    .A(_04179_),
    .Y(_04184_));
 sg13g2_o21ai_1 _11884_ (.B1(_04184_),
    .Y(_04185_),
    .A1(\clock_inst.min_c[49] ),
    .A2(net51));
 sg13g2_o21ai_1 _11885_ (.B1(net125),
    .Y(_04186_),
    .A1(net47),
    .A2(_04183_));
 sg13g2_inv_1 _11886_ (.Y(_04187_),
    .A(_04179_));
 sg13g2_a22oi_1 _11887_ (.Y(_00351_),
    .B1(_04186_),
    .B2(_04187_),
    .A2(_04185_),
    .A1(net108));
 sg13g2_inv_1 _11888_ (.Y(_04188_),
    .A(_03694_));
 sg13g2_a21oi_1 _11889_ (.A1(_03701_),
    .A2(_03779_),
    .Y(_04189_),
    .B1(_03782_));
 sg13g2_xor2_1 _11890_ (.B(_03694_),
    .A(_03094_),
    .X(_04190_));
 sg13g2_xnor2_1 _11891_ (.Y(_04191_),
    .A(_04189_),
    .B(_04190_));
 sg13g2_nand2_1 _11892_ (.Y(_04192_),
    .A(\clock_inst.min_c[4] ),
    .B(net85));
 sg13g2_o21ai_1 _11893_ (.B1(_04192_),
    .Y(_04193_),
    .A1(net86),
    .A2(_04191_));
 sg13g2_nor2_1 _11894_ (.A(net124),
    .B(_04193_),
    .Y(_04194_));
 sg13g2_a21oi_1 _11895_ (.A1(_04188_),
    .A2(net67),
    .Y(_00352_),
    .B1(_04194_));
 sg13g2_buf_1 _11896_ (.A(\clock_inst.min_tile.e0[50] ),
    .X(_04195_));
 sg13g2_inv_1 _11897_ (.Y(_04196_),
    .A(_04195_));
 sg13g2_and2_1 _11898_ (.A(_04187_),
    .B(_04182_),
    .X(_04197_));
 sg13g2_buf_1 _11899_ (.A(_04197_),
    .X(_04198_));
 sg13g2_nor3_1 _11900_ (.A(_04155_),
    .B(_04187_),
    .C(_04138_),
    .Y(_04199_));
 sg13g2_and4_1 _11901_ (.A(_04161_),
    .B(_04171_),
    .C(_04163_),
    .D(_04199_),
    .X(_04200_));
 sg13g2_nand2_1 _11902_ (.Y(_04201_),
    .A(_04107_),
    .B(_04142_));
 sg13g2_nand2_1 _11903_ (.Y(_04202_),
    .A(_03067_),
    .B(_04142_));
 sg13g2_a221oi_1 _11904_ (.B2(_04202_),
    .C1(_04113_),
    .B1(_04201_),
    .A1(_04114_),
    .Y(_04203_),
    .A2(_04109_));
 sg13g2_nor4_1 _11905_ (.A(_04085_),
    .B(_04089_),
    .C(_04113_),
    .D(_04201_),
    .Y(_04204_));
 sg13g2_nor4_1 _11906_ (.A(_04085_),
    .B(_04089_),
    .C(_04113_),
    .D(_04202_),
    .Y(_04205_));
 sg13g2_nor3_1 _11907_ (.A(_03066_),
    .B(_04106_),
    .C(_04143_),
    .Y(_04206_));
 sg13g2_nor4_1 _11908_ (.A(_04203_),
    .B(_04204_),
    .C(_04205_),
    .D(_04206_),
    .Y(_04207_));
 sg13g2_nand2_1 _11909_ (.Y(_04208_),
    .A(_04195_),
    .B(net99));
 sg13g2_a221oi_1 _11910_ (.B2(_04207_),
    .C1(_04208_),
    .B1(_04200_),
    .A1(_04146_),
    .Y(_04209_),
    .A2(_04198_));
 sg13g2_nor2_1 _11911_ (.A(_04195_),
    .B(_01274_),
    .Y(_04210_));
 sg13g2_and3_1 _11912_ (.X(_04211_),
    .A(_04146_),
    .B(_04198_),
    .C(_04210_));
 sg13g2_nand2_1 _11913_ (.Y(_04212_),
    .A(_04179_),
    .B(_04180_));
 sg13g2_nor4_2 _11914_ (.A(_04137_),
    .B(_04138_),
    .C(_04144_),
    .Y(_04213_),
    .D(_04212_));
 sg13g2_and2_1 _11915_ (.A(_04213_),
    .B(_04210_),
    .X(_04214_));
 sg13g2_and2_1 _11916_ (.A(\clock_inst.min_c[50] ),
    .B(_01610_),
    .X(_04215_));
 sg13g2_nor4_2 _11917_ (.A(_04209_),
    .B(_04211_),
    .C(_04214_),
    .Y(_04216_),
    .D(_04215_));
 sg13g2_o21ai_1 _11918_ (.B1(_04216_),
    .Y(_00353_),
    .A1(_04196_),
    .A2(net106));
 sg13g2_inv_1 _11919_ (.Y(_04217_),
    .A(\clock_inst.min_tile.e0[51] ));
 sg13g2_and3_1 _11920_ (.X(_04218_),
    .A(_04196_),
    .B(net66),
    .C(_04198_));
 sg13g2_a21oi_1 _11921_ (.A1(_04195_),
    .A2(_04213_),
    .Y(_04219_),
    .B1(_04218_));
 sg13g2_a21o_1 _11922_ (.A2(_04219_),
    .A1(net93),
    .B1(net153),
    .X(_04220_));
 sg13g2_nand3b_1 _11923_ (.B(\clock_inst.min_tile.e0[51] ),
    .C(net152),
    .Y(_04221_),
    .A_N(_04219_));
 sg13g2_o21ai_1 _11924_ (.B1(_04221_),
    .Y(_04222_),
    .A1(\clock_inst.min_c[51] ),
    .A2(net152));
 sg13g2_a22oi_1 _11925_ (.Y(_00354_),
    .B1(_04222_),
    .B2(net103),
    .A2(_04220_),
    .A1(_04217_));
 sg13g2_inv_1 _11926_ (.Y(_04223_),
    .A(\clock_inst.min_tile.e0[52] ));
 sg13g2_nor2_1 _11927_ (.A(_04196_),
    .B(_04217_),
    .Y(_04224_));
 sg13g2_a22oi_1 _11928_ (.Y(_04225_),
    .B1(_04224_),
    .B2(_04213_),
    .A2(_04218_),
    .A1(_04217_));
 sg13g2_xnor2_1 _11929_ (.Y(_04226_),
    .A(\clock_inst.min_tile.e0[52] ),
    .B(_04225_));
 sg13g2_nand2_1 _11930_ (.Y(_04227_),
    .A(net152),
    .B(_04226_));
 sg13g2_a21oi_1 _11931_ (.A1(\clock_inst.min_c[52] ),
    .A2(_01186_),
    .Y(_04228_),
    .B1(net162));
 sg13g2_a22oi_1 _11932_ (.Y(_00355_),
    .B1(_04227_),
    .B2(_04228_),
    .A2(net69),
    .A1(_04223_));
 sg13g2_nor2_1 _11933_ (.A(\clock_inst.min_tile.e0[53] ),
    .B(_01274_),
    .Y(_04229_));
 sg13g2_and2_1 _11934_ (.A(\clock_inst.min_tile.e0[53] ),
    .B(net99),
    .X(_04230_));
 sg13g2_nor3_1 _11935_ (.A(_04179_),
    .B(_04195_),
    .C(_04147_),
    .Y(_04231_));
 sg13g2_and4_1 _11936_ (.A(_04217_),
    .B(_04223_),
    .C(_04181_),
    .D(_04231_),
    .X(_04232_));
 sg13g2_and2_1 _11937_ (.A(\clock_inst.min_tile.e0[52] ),
    .B(_04224_),
    .X(_04233_));
 sg13g2_a22oi_1 _11938_ (.Y(_04234_),
    .B1(_04233_),
    .B2(_04213_),
    .A2(_04232_),
    .A1(net66));
 sg13g2_mux2_1 _11939_ (.A0(_04229_),
    .A1(_04230_),
    .S(_04234_),
    .X(_04235_));
 sg13g2_a21o_1 _11940_ (.A2(_01610_),
    .A1(\clock_inst.min_c[53] ),
    .B1(_04235_),
    .X(_04236_));
 sg13g2_a21o_1 _11941_ (.A2(net76),
    .A1(\clock_inst.min_tile.e0[53] ),
    .B1(_04236_),
    .X(_00356_));
 sg13g2_nand3_1 _11942_ (.B(_03704_),
    .C(_03707_),
    .A(_03700_),
    .Y(_04237_));
 sg13g2_xnor2_1 _11943_ (.Y(_04238_),
    .A(_03108_),
    .B(_03705_));
 sg13g2_xnor2_1 _11944_ (.Y(_04239_),
    .A(_04237_),
    .B(_04238_));
 sg13g2_nand2_1 _11945_ (.Y(_04240_),
    .A(\clock_inst.min_c[5] ),
    .B(net85));
 sg13g2_o21ai_1 _11946_ (.B1(_04240_),
    .Y(_04241_),
    .A1(net86),
    .A2(_04239_));
 sg13g2_nor2_1 _11947_ (.A(net124),
    .B(_04241_),
    .Y(_04242_));
 sg13g2_a21oi_1 _11948_ (.A1(_03713_),
    .A2(net67),
    .Y(_00357_),
    .B1(_04242_));
 sg13g2_inv_1 _11949_ (.Y(_04243_),
    .A(_03682_));
 sg13g2_xnor2_1 _11950_ (.Y(_04244_),
    .A(_03683_),
    .B(_03789_));
 sg13g2_nand2_1 _11951_ (.Y(_04245_),
    .A(\clock_inst.min_c[6] ),
    .B(net141));
 sg13g2_o21ai_1 _11952_ (.B1(_04245_),
    .Y(_04246_),
    .A1(net90),
    .A2(_04244_));
 sg13g2_nor2_1 _11953_ (.A(net124),
    .B(_04246_),
    .Y(_04247_));
 sg13g2_a21oi_1 _11954_ (.A1(_04243_),
    .A2(net67),
    .Y(_00358_),
    .B1(_04247_));
 sg13g2_inv_1 _11955_ (.Y(_04248_),
    .A(_03680_));
 sg13g2_a21o_1 _11956_ (.A2(_03789_),
    .A1(_03682_),
    .B1(_03110_),
    .X(_04249_));
 sg13g2_o21ai_1 _11957_ (.B1(_04249_),
    .Y(_04250_),
    .A1(_03682_),
    .A2(_03789_));
 sg13g2_xnor2_1 _11958_ (.Y(_04251_),
    .A(_03681_),
    .B(_04250_));
 sg13g2_o21ai_1 _11959_ (.B1(net240),
    .Y(_04252_),
    .A1(\clock_inst.min_c[7] ),
    .A2(net104));
 sg13g2_a21o_1 _11960_ (.A2(_04251_),
    .A1(net91),
    .B1(_04252_),
    .X(_04253_));
 sg13g2_o21ai_1 _11961_ (.B1(_04253_),
    .Y(_00359_),
    .A1(_04248_),
    .A2(net106));
 sg13g2_xnor2_1 _11962_ (.Y(_04254_),
    .A(_03741_),
    .B(_03742_));
 sg13g2_nor2_1 _11963_ (.A(\clock_inst.min_c[8] ),
    .B(net150),
    .Y(_04255_));
 sg13g2_a21oi_1 _11964_ (.A1(net101),
    .A2(_04254_),
    .Y(_04256_),
    .B1(_04255_));
 sg13g2_nand2_1 _11965_ (.Y(_04257_),
    .A(net144),
    .B(_04256_));
 sg13g2_o21ai_1 _11966_ (.B1(_04257_),
    .Y(_00360_),
    .A1(_03766_),
    .A2(net139));
 sg13g2_nand2_1 _11967_ (.Y(_04258_),
    .A(\clock_inst.min_c[9] ),
    .B(net107));
 sg13g2_o21ai_1 _11968_ (.B1(net243),
    .Y(_04259_),
    .A1(_03676_),
    .A2(_03678_));
 sg13g2_or3_1 _11969_ (.A(net241),
    .B(_03676_),
    .C(_03678_),
    .X(_04260_));
 sg13g2_mux2_1 _11970_ (.A0(_04259_),
    .A1(_04260_),
    .S(_03722_),
    .X(_04261_));
 sg13g2_a21o_1 _11971_ (.A2(_04261_),
    .A1(_04258_),
    .B1(net154),
    .X(_04262_));
 sg13g2_o21ai_1 _11972_ (.B1(_04262_),
    .Y(_00361_),
    .A1(_03677_),
    .A2(net139));
 sg13g2_nand2_1 _11973_ (.Y(_04263_),
    .A(\clock_inst.min_a[0] ),
    .B(net355));
 sg13g2_xor2_1 _11974_ (.B(_04263_),
    .A(\clock_inst.min_tile.e[0] ),
    .X(_04264_));
 sg13g2_o21ai_1 _11975_ (.B1(_03668_),
    .Y(_00362_),
    .A1(net135),
    .A2(_04264_));
 sg13g2_buf_1 _11976_ (.A(\clock_inst.min_tile.e[10] ),
    .X(_04265_));
 sg13g2_buf_1 _11977_ (.A(\clock_inst.min_tile.e[9] ),
    .X(_04266_));
 sg13g2_nand3_1 _11978_ (.B(net565),
    .C(net499),
    .A(net535),
    .Y(_04267_));
 sg13g2_nand3b_1 _11979_ (.B(net499),
    .C(net569),
    .Y(_04268_),
    .A_N(_04266_));
 sg13g2_buf_2 _11980_ (.A(\clock_inst.min_tile.e[8] ),
    .X(_04269_));
 sg13g2_buf_1 _11981_ (.A(\clock_inst.min_tile.e[3] ),
    .X(_04270_));
 sg13g2_inv_1 _11982_ (.Y(_04271_),
    .A(_04270_));
 sg13g2_or2_1 _11983_ (.X(_04272_),
    .B(\clock_inst.min_tile.e[2] ),
    .A(\clock_inst.min_a[2] ));
 sg13g2_nand2_1 _11984_ (.Y(_04273_),
    .A(\clock_inst.min_a[0] ),
    .B(\clock_inst.min_tile.e[0] ));
 sg13g2_nor2_1 _11985_ (.A(_02396_),
    .B(\clock_inst.min_tile.e[1] ),
    .Y(_04274_));
 sg13g2_nand2_1 _11986_ (.Y(_04275_),
    .A(_02396_),
    .B(\clock_inst.min_tile.e[1] ));
 sg13g2_o21ai_1 _11987_ (.B1(_04275_),
    .Y(_04276_),
    .A1(_04273_),
    .A2(_04274_));
 sg13g2_buf_1 _11988_ (.A(_04276_),
    .X(_04277_));
 sg13g2_and2_1 _11989_ (.A(\clock_inst.min_a[2] ),
    .B(\clock_inst.min_tile.e[2] ),
    .X(_04278_));
 sg13g2_buf_1 _11990_ (.A(_04278_),
    .X(_04279_));
 sg13g2_a21oi_2 _11991_ (.B1(_04279_),
    .Y(_04280_),
    .A2(_04277_),
    .A1(_04272_));
 sg13g2_and2_1 _11992_ (.A(_04270_),
    .B(_04272_),
    .X(_04281_));
 sg13g2_a221oi_1 _11993_ (.B2(_04277_),
    .C1(\clock_inst.min_a[3] ),
    .B1(_04281_),
    .A1(_04270_),
    .Y(_04282_),
    .A2(_04279_));
 sg13g2_a21oi_2 _11994_ (.B1(_04282_),
    .Y(_04283_),
    .A2(_04280_),
    .A1(_04271_));
 sg13g2_buf_1 _11995_ (.A(\clock_inst.min_tile.e[4] ),
    .X(_04284_));
 sg13g2_inv_1 _11996_ (.Y(_04285_),
    .A(_04284_));
 sg13g2_nor2_1 _11997_ (.A(_02788_),
    .B(\clock_inst.min_tile.e[5] ),
    .Y(_04286_));
 sg13g2_a21oi_1 _11998_ (.A1(_02766_),
    .A2(_04285_),
    .Y(_04287_),
    .B1(_04286_));
 sg13g2_buf_2 _11999_ (.A(\clock_inst.min_tile.e[6] ),
    .X(_04288_));
 sg13g2_buf_1 _12000_ (.A(\clock_inst.min_tile.e[7] ),
    .X(_04289_));
 sg13g2_nand2_1 _12001_ (.Y(_04290_),
    .A(_02837_),
    .B(_04289_));
 sg13g2_nand2b_1 _12002_ (.Y(_04291_),
    .B(_04290_),
    .A_N(_04288_));
 sg13g2_nand2_1 _12003_ (.Y(_04292_),
    .A(_02815_),
    .B(_04290_));
 sg13g2_a22oi_1 _12004_ (.Y(_04293_),
    .B1(_02788_),
    .B2(\clock_inst.min_tile.e[5] ),
    .A2(_04284_),
    .A1(_02765_));
 sg13g2_nor2_1 _12005_ (.A(_04286_),
    .B(_04293_),
    .Y(_04294_));
 sg13g2_a221oi_1 _12006_ (.B2(_04292_),
    .C1(_04294_),
    .B1(_04291_),
    .A1(_04283_),
    .Y(_04295_),
    .A2(_04287_));
 sg13g2_nor2_1 _12007_ (.A(_02814_),
    .B(_04288_),
    .Y(_04296_));
 sg13g2_nor2_1 _12008_ (.A(_02837_),
    .B(_04289_),
    .Y(_04297_));
 sg13g2_a21o_1 _12009_ (.A2(_04296_),
    .A1(_04290_),
    .B1(_04297_),
    .X(_04298_));
 sg13g2_nor2_1 _12010_ (.A(_04295_),
    .B(_04298_),
    .Y(_04299_));
 sg13g2_nor2b_1 _12011_ (.A(_04297_),
    .B_N(net567),
    .Y(_04300_));
 sg13g2_nand2_1 _12012_ (.Y(_04301_),
    .A(\clock_inst.min_a[3] ),
    .B(_04287_));
 sg13g2_a21oi_2 _12013_ (.B1(_04301_),
    .Y(_04302_),
    .A2(_04280_),
    .A1(_04271_));
 sg13g2_and2_1 _12014_ (.A(_04270_),
    .B(_04279_),
    .X(_04303_));
 sg13g2_a21o_1 _12015_ (.A2(_04281_),
    .A1(_04277_),
    .B1(_04303_),
    .X(_04304_));
 sg13g2_a21o_1 _12016_ (.A2(_04287_),
    .A1(_04304_),
    .B1(_04294_),
    .X(_04305_));
 sg13g2_buf_1 _12017_ (.A(_04305_),
    .X(_04306_));
 sg13g2_nor3_1 _12018_ (.A(_04288_),
    .B(_04302_),
    .C(_04306_),
    .Y(_04307_));
 sg13g2_o21ai_1 _12019_ (.B1(_04288_),
    .Y(_04308_),
    .A1(_04302_),
    .A2(_04306_));
 sg13g2_o21ai_1 _12020_ (.B1(_04308_),
    .Y(_04309_),
    .A1(_02815_),
    .A2(_04307_));
 sg13g2_and2_1 _12021_ (.A(_02837_),
    .B(_04289_),
    .X(_04310_));
 sg13g2_o21ai_1 _12022_ (.B1(net567),
    .Y(_04311_),
    .A1(_04269_),
    .A2(_04310_));
 sg13g2_inv_1 _12023_ (.Y(_04312_),
    .A(_04311_));
 sg13g2_a221oi_1 _12024_ (.B2(_04309_),
    .C1(_04312_),
    .B1(_04300_),
    .A1(_04269_),
    .Y(_04313_),
    .A2(_04299_));
 sg13g2_buf_2 _12025_ (.A(_04313_),
    .X(_04314_));
 sg13g2_mux2_1 _12026_ (.A0(_04267_),
    .A1(_04268_),
    .S(_04314_),
    .X(_04315_));
 sg13g2_xor2_1 _12027_ (.B(_04315_),
    .A(_04265_),
    .X(_04316_));
 sg13g2_a22oi_1 _12028_ (.Y(_00363_),
    .B1(_04316_),
    .B2(net78),
    .A2(_03725_),
    .A1(_03724_));
 sg13g2_buf_1 _12029_ (.A(\clock_inst.min_tile.e[11] ),
    .X(_04317_));
 sg13g2_nand4_1 _12030_ (.B(net565),
    .C(_04265_),
    .A(net535),
    .Y(_04318_),
    .D(net499));
 sg13g2_nor2_1 _12031_ (.A(net565),
    .B(_04265_),
    .Y(_04319_));
 sg13g2_nand3_1 _12032_ (.B(net445),
    .C(_04319_),
    .A(net569),
    .Y(_04320_));
 sg13g2_mux2_1 _12033_ (.A0(_04318_),
    .A1(_04320_),
    .S(_04314_),
    .X(_04321_));
 sg13g2_xor2_1 _12034_ (.B(_04321_),
    .A(_04317_),
    .X(_04322_));
 sg13g2_a22oi_1 _12035_ (.Y(_00364_),
    .B1(_04322_),
    .B2(net78),
    .A2(_03736_),
    .A1(_03735_));
 sg13g2_nand2b_1 _12036_ (.Y(_04323_),
    .B(_04319_),
    .A_N(_04317_));
 sg13g2_a22oi_1 _12037_ (.Y(_04324_),
    .B1(net569),
    .B2(_04323_),
    .A2(_04269_),
    .A1(net567));
 sg13g2_buf_1 _12038_ (.A(_04324_),
    .X(_04325_));
 sg13g2_nand3_1 _12039_ (.B(_04265_),
    .C(_04317_),
    .A(net565),
    .Y(_04326_));
 sg13g2_nor2_1 _12040_ (.A(_04325_),
    .B(_04326_),
    .Y(_04327_));
 sg13g2_nor3_1 _12041_ (.A(net565),
    .B(_04265_),
    .C(_04317_),
    .Y(_04328_));
 sg13g2_and3_1 _12042_ (.X(_04329_),
    .A(net565),
    .B(_04265_),
    .C(_04317_));
 sg13g2_buf_1 _12043_ (.A(_04329_),
    .X(_04330_));
 sg13g2_a21oi_1 _12044_ (.A1(net569),
    .A2(_04328_),
    .Y(_04331_),
    .B1(_04330_));
 sg13g2_nor2_1 _12045_ (.A(net567),
    .B(_04269_),
    .Y(_04332_));
 sg13g2_nand3_1 _12046_ (.B(_04269_),
    .C(_04326_),
    .A(net567),
    .Y(_04333_));
 sg13g2_nand2b_1 _12047_ (.Y(_04334_),
    .B(_04333_),
    .A_N(_04332_));
 sg13g2_nor4_1 _12048_ (.A(_04295_),
    .B(_04298_),
    .C(_04331_),
    .D(_04334_),
    .Y(_04335_));
 sg13g2_o21ai_1 _12049_ (.B1(net535),
    .Y(_04336_),
    .A1(_04327_),
    .A2(_04335_));
 sg13g2_inv_1 _12050_ (.Y(_04337_),
    .A(_04298_));
 sg13g2_nand2_1 _12051_ (.Y(_04338_),
    .A(net569),
    .B(_04328_));
 sg13g2_nand2_1 _12052_ (.Y(_04339_),
    .A(net535),
    .B(_04330_));
 sg13g2_xnor2_1 _12053_ (.Y(_04340_),
    .A(net567),
    .B(_04269_));
 sg13g2_a21oi_1 _12054_ (.A1(_04338_),
    .A2(_04339_),
    .Y(_04341_),
    .B1(_04340_));
 sg13g2_nand3b_1 _12055_ (.B(_04337_),
    .C(_04341_),
    .Y(_04342_),
    .A_N(_04295_));
 sg13g2_nand3_1 _12056_ (.B(_04325_),
    .C(_04342_),
    .A(net569),
    .Y(_04343_));
 sg13g2_buf_2 _12057_ (.A(\clock_inst.min_tile.e[12] ),
    .X(_04344_));
 sg13g2_nand2_1 _12058_ (.Y(_04345_),
    .A(_04344_),
    .B(net442));
 sg13g2_a21o_1 _12059_ (.A2(_04343_),
    .A1(_04336_),
    .B1(_04345_),
    .X(_04346_));
 sg13g2_a21oi_1 _12060_ (.A1(net161),
    .A2(_04346_),
    .Y(_04347_),
    .B1(_03756_));
 sg13g2_nand3b_1 _12061_ (.B(_04336_),
    .C(_04343_),
    .Y(_04348_),
    .A_N(_04344_));
 sg13g2_nor2_1 _12062_ (.A(_03756_),
    .B(_04348_),
    .Y(_04349_));
 sg13g2_nor2_1 _12063_ (.A(_04344_),
    .B(net80),
    .Y(_04350_));
 sg13g2_nor3_1 _12064_ (.A(_04347_),
    .B(_04349_),
    .C(_04350_),
    .Y(_00365_));
 sg13g2_buf_1 _12065_ (.A(\clock_inst.min_tile.e[13] ),
    .X(_04351_));
 sg13g2_nand4_1 _12066_ (.B(_04344_),
    .C(net499),
    .A(net535),
    .Y(_04352_),
    .D(_04330_));
 sg13g2_nor3_1 _12067_ (.A(net535),
    .B(_04344_),
    .C(net542),
    .Y(_04353_));
 sg13g2_nand3_1 _12068_ (.B(_04342_),
    .C(_04353_),
    .A(_04325_),
    .Y(_04354_));
 sg13g2_o21ai_1 _12069_ (.B1(_04354_),
    .Y(_04355_),
    .A1(_04314_),
    .A2(_04352_));
 sg13g2_xnor2_1 _12070_ (.Y(_04356_),
    .A(_04351_),
    .B(_04355_));
 sg13g2_a22oi_1 _12071_ (.Y(_00366_),
    .B1(_04356_),
    .B2(net78),
    .A2(_03765_),
    .A1(_03764_));
 sg13g2_buf_1 _12072_ (.A(\clock_inst.min_tile.e[14] ),
    .X(_04357_));
 sg13g2_and2_1 _12073_ (.A(_02814_),
    .B(_04288_),
    .X(_04358_));
 sg13g2_nor4_1 _12074_ (.A(_04310_),
    .B(_04297_),
    .C(_04296_),
    .D(_04358_),
    .Y(_04359_));
 sg13g2_nand2_1 _12075_ (.Y(_04360_),
    .A(_04344_),
    .B(_04351_));
 sg13g2_or3_1 _12076_ (.A(_02250_),
    .B(_04344_),
    .C(_04351_),
    .X(_04361_));
 sg13g2_buf_1 _12077_ (.A(_04361_),
    .X(_04362_));
 sg13g2_o21ai_1 _12078_ (.B1(_04362_),
    .Y(_04363_),
    .A1(net569),
    .A2(_04360_));
 sg13g2_and3_1 _12079_ (.X(_04364_),
    .A(_04341_),
    .B(_04359_),
    .C(_04363_));
 sg13g2_o21ai_1 _12080_ (.B1(_04364_),
    .Y(_04365_),
    .A1(_04302_),
    .A2(_04306_));
 sg13g2_nand2_1 _12081_ (.Y(_04366_),
    .A(_02814_),
    .B(_04288_));
 sg13g2_a21oi_1 _12082_ (.A1(_04290_),
    .A2(_04366_),
    .Y(_04367_),
    .B1(_04297_));
 sg13g2_a21oi_1 _12083_ (.A1(net567),
    .A2(_04269_),
    .Y(_04368_),
    .B1(_04367_));
 sg13g2_nor2_1 _12084_ (.A(_04332_),
    .B(_04368_),
    .Y(_04369_));
 sg13g2_nand4_1 _12085_ (.B(_04351_),
    .C(_04330_),
    .A(_04344_),
    .Y(_04370_),
    .D(_04369_));
 sg13g2_a21o_1 _12086_ (.A2(_04370_),
    .A1(_04365_),
    .B1(_02249_),
    .X(_04371_));
 sg13g2_nor3_1 _12087_ (.A(_04323_),
    .B(_04362_),
    .C(_04369_),
    .Y(_04372_));
 sg13g2_nand2_1 _12088_ (.Y(_04373_),
    .A(_04365_),
    .B(_04372_));
 sg13g2_a21oi_1 _12089_ (.A1(_04371_),
    .A2(_04373_),
    .Y(_04374_),
    .B1(net502));
 sg13g2_xnor2_1 _12090_ (.Y(_04375_),
    .A(_04357_),
    .B(_04374_));
 sg13g2_nand3_1 _12091_ (.B(net150),
    .C(_03796_),
    .A(_03797_),
    .Y(_04376_));
 sg13g2_nand2_1 _12092_ (.Y(_04377_),
    .A(_03201_),
    .B(net141));
 sg13g2_nand3_1 _12093_ (.B(_04376_),
    .C(_04377_),
    .A(net233),
    .Y(_04378_));
 sg13g2_o21ai_1 _12094_ (.B1(_04378_),
    .Y(_04379_),
    .A1(net156),
    .A2(_04375_));
 sg13g2_and2_1 _12095_ (.A(_03797_),
    .B(_03793_),
    .X(_04380_));
 sg13g2_nor3_1 _12096_ (.A(_03797_),
    .B(_03793_),
    .C(_03796_),
    .Y(_04381_));
 sg13g2_a21oi_1 _12097_ (.A1(\clock_inst.min_c[14] ),
    .A2(net96),
    .Y(_04382_),
    .B1(net143));
 sg13g2_o21ai_1 _12098_ (.B1(_04382_),
    .Y(_04383_),
    .A1(_04380_),
    .A2(_04381_));
 sg13g2_and2_1 _12099_ (.A(_04379_),
    .B(_04383_),
    .X(_00367_));
 sg13g2_nand2_1 _12100_ (.Y(_04384_),
    .A(net535),
    .B(_04357_));
 sg13g2_nor4_1 _12101_ (.A(net542),
    .B(_04326_),
    .C(_04360_),
    .D(_04384_),
    .Y(_04385_));
 sg13g2_nor4_1 _12102_ (.A(_04357_),
    .B(net542),
    .C(_04323_),
    .D(_04362_),
    .Y(_04386_));
 sg13g2_mux2_1 _12103_ (.A0(_04385_),
    .A1(_04386_),
    .S(_04314_),
    .X(_04387_));
 sg13g2_xnor2_1 _12104_ (.Y(_04388_),
    .A(\clock_inst.min_tile.e[15] ),
    .B(_04387_));
 sg13g2_a22oi_1 _12105_ (.Y(_00368_),
    .B1(_04388_),
    .B2(net78),
    .A2(_03814_),
    .A1(_03813_));
 sg13g2_inv_1 _12106_ (.Y(_04389_),
    .A(\clock_inst.min_tile.e[15] ));
 sg13g2_nor4_1 _12107_ (.A(_04389_),
    .B(_01675_),
    .C(_04360_),
    .D(_04384_),
    .Y(_04390_));
 sg13g2_o21ai_1 _12108_ (.B1(_04390_),
    .Y(_04391_),
    .A1(_04327_),
    .A2(_04335_));
 sg13g2_nor4_1 _12109_ (.A(_04357_),
    .B(\clock_inst.min_tile.e[15] ),
    .C(_01675_),
    .D(_04362_),
    .Y(_04392_));
 sg13g2_nand3_1 _12110_ (.B(_04342_),
    .C(_04392_),
    .A(_04325_),
    .Y(_04393_));
 sg13g2_nand2_1 _12111_ (.Y(_04394_),
    .A(_04391_),
    .B(_04393_));
 sg13g2_xor2_1 _12112_ (.B(_04394_),
    .A(\clock_inst.min_tile.e[16] ),
    .X(_04395_));
 sg13g2_mux2_1 _12113_ (.A0(_03822_),
    .A1(_04395_),
    .S(net76),
    .X(_00369_));
 sg13g2_mux2_1 _12114_ (.A0(_04393_),
    .A1(_04391_),
    .S(\clock_inst.min_tile.e[16] ),
    .X(_04396_));
 sg13g2_xor2_1 _12115_ (.B(_04396_),
    .A(\clock_inst.min_tile.e[17] ),
    .X(_04397_));
 sg13g2_a221oi_1 _12116_ (.B2(net76),
    .C1(_03831_),
    .B1(_04397_),
    .A1(_03824_),
    .Y(_00370_),
    .A2(net82));
 sg13g2_buf_1 _12117_ (.A(\clock_inst.min_tile.e[18] ),
    .X(_04398_));
 sg13g2_inv_1 _12118_ (.Y(_04399_),
    .A(_04398_));
 sg13g2_a22oi_1 _12119_ (.Y(_04400_),
    .B1(_01802_),
    .B2(_04398_),
    .A2(net49),
    .A1(_03832_));
 sg13g2_nand3_1 _12120_ (.B(net240),
    .C(_01215_),
    .A(_03832_),
    .Y(_04401_));
 sg13g2_nand2_1 _12121_ (.Y(_04402_),
    .A(_04398_),
    .B(net239));
 sg13g2_a21oi_1 _12122_ (.A1(_04401_),
    .A2(_04402_),
    .Y(_04403_),
    .B1(_02345_));
 sg13g2_a21oi_1 _12123_ (.A1(_02345_),
    .A2(_04400_),
    .Y(_04404_),
    .B1(_04403_));
 sg13g2_a21oi_1 _12124_ (.A1(_04399_),
    .A2(net137),
    .Y(_00371_),
    .B1(_04404_));
 sg13g2_nand2_1 _12125_ (.Y(_04405_),
    .A(_02345_),
    .B(_04398_));
 sg13g2_xor2_1 _12126_ (.B(_04405_),
    .A(_02347_),
    .X(_04406_));
 sg13g2_nor2_1 _12127_ (.A(net441),
    .B(_04406_),
    .Y(_04407_));
 sg13g2_xnor2_1 _12128_ (.Y(_04408_),
    .A(\clock_inst.min_tile.e[19] ),
    .B(_04407_));
 sg13g2_a21oi_1 _12129_ (.A1(net74),
    .A2(_04408_),
    .Y(_00372_),
    .B1(_03843_));
 sg13g2_xnor2_1 _12130_ (.Y(_04409_),
    .A(_02396_),
    .B(_04273_));
 sg13g2_nand2_1 _12131_ (.Y(_04410_),
    .A(net357),
    .B(_04409_));
 sg13g2_xor2_1 _12132_ (.B(_04410_),
    .A(\clock_inst.min_tile.e[1] ),
    .X(_04411_));
 sg13g2_a21oi_1 _12133_ (.A1(net74),
    .A2(_04411_),
    .Y(_00373_),
    .B1(_03851_));
 sg13g2_nor2_1 _12134_ (.A(_02347_),
    .B(\clock_inst.min_tile.e[19] ),
    .Y(_04412_));
 sg13g2_nand2_1 _12135_ (.Y(_04413_),
    .A(_02347_),
    .B(\clock_inst.min_tile.e[19] ));
 sg13g2_o21ai_1 _12136_ (.B1(_04413_),
    .Y(_04414_),
    .A1(_04405_),
    .A2(_04412_));
 sg13g2_xor2_1 _12137_ (.B(_04414_),
    .A(_02460_),
    .X(_04415_));
 sg13g2_nand2_1 _12138_ (.Y(_04416_),
    .A(net442),
    .B(_04415_));
 sg13g2_xnor2_1 _12139_ (.Y(_04417_),
    .A(\clock_inst.min_tile.e[20] ),
    .B(_04416_));
 sg13g2_xor2_1 _12140_ (.B(_03856_),
    .A(_03852_),
    .X(_04418_));
 sg13g2_a22oi_1 _12141_ (.Y(_04419_),
    .B1(_04418_),
    .B2(net23),
    .A2(_04417_),
    .A1(net83));
 sg13g2_inv_1 _12142_ (.Y(_00374_),
    .A(_04419_));
 sg13g2_buf_1 _12143_ (.A(net140),
    .X(_04420_));
 sg13g2_buf_1 _12144_ (.A(\clock_inst.min_tile.e[21] ),
    .X(_04421_));
 sg13g2_or2_1 _12145_ (.X(_04422_),
    .B(\clock_inst.min_tile.e[20] ),
    .A(_02460_));
 sg13g2_and2_1 _12146_ (.A(_02460_),
    .B(\clock_inst.min_tile.e[20] ),
    .X(_04423_));
 sg13g2_a21o_1 _12147_ (.A2(_04422_),
    .A1(_04414_),
    .B1(_04423_),
    .X(_04424_));
 sg13g2_buf_1 _12148_ (.A(_04424_),
    .X(_04425_));
 sg13g2_xnor2_1 _12149_ (.Y(_04426_),
    .A(_02497_),
    .B(_04425_));
 sg13g2_nor2_1 _12150_ (.A(net441),
    .B(_04426_),
    .Y(_04427_));
 sg13g2_xnor2_1 _12151_ (.Y(_04428_),
    .A(_04421_),
    .B(_04427_));
 sg13g2_a21oi_1 _12152_ (.A1(net65),
    .A2(_04428_),
    .Y(_00375_),
    .B1(_03869_));
 sg13g2_a21o_1 _12153_ (.A2(_04425_),
    .A1(_04421_),
    .B1(_02497_),
    .X(_04429_));
 sg13g2_o21ai_1 _12154_ (.B1(_04429_),
    .Y(_04430_),
    .A1(_04421_),
    .A2(_04425_));
 sg13g2_xor2_1 _12155_ (.B(_04430_),
    .A(_02499_),
    .X(_04431_));
 sg13g2_nor2_1 _12156_ (.A(net441),
    .B(_04431_),
    .Y(_04432_));
 sg13g2_xnor2_1 _12157_ (.Y(_04433_),
    .A(\clock_inst.min_tile.e[22] ),
    .B(_04432_));
 sg13g2_a21oi_1 _12158_ (.A1(net65),
    .A2(_04433_),
    .Y(_00376_),
    .B1(_03878_));
 sg13g2_buf_1 _12159_ (.A(\clock_inst.min_tile.e[23] ),
    .X(_04434_));
 sg13g2_a221oi_1 _12160_ (.B2(_04422_),
    .C1(_04423_),
    .B1(_04414_),
    .A1(_02497_),
    .Y(_04435_),
    .A2(_04421_));
 sg13g2_or2_1 _12161_ (.X(_04436_),
    .B(\clock_inst.min_tile.e[22] ),
    .A(_02499_));
 sg13g2_o21ai_1 _12162_ (.B1(_04436_),
    .Y(_04437_),
    .A1(_02497_),
    .A2(_04421_));
 sg13g2_nand2_1 _12163_ (.Y(_04438_),
    .A(_02499_),
    .B(\clock_inst.min_tile.e[22] ));
 sg13g2_o21ai_1 _12164_ (.B1(_04438_),
    .Y(_04439_),
    .A1(_04435_),
    .A2(_04437_));
 sg13g2_buf_2 _12165_ (.A(_04439_),
    .X(_04440_));
 sg13g2_xnor2_1 _12166_ (.Y(_04441_),
    .A(\clock_inst.min_a[23] ),
    .B(_04440_));
 sg13g2_nor2_1 _12167_ (.A(net441),
    .B(_04441_),
    .Y(_04442_));
 sg13g2_xnor2_1 _12168_ (.Y(_04443_),
    .A(_04434_),
    .B(_04442_));
 sg13g2_a21oi_1 _12169_ (.A1(net65),
    .A2(_04443_),
    .Y(_00377_),
    .B1(_03888_));
 sg13g2_buf_1 _12170_ (.A(\clock_inst.min_tile.e[24] ),
    .X(_04444_));
 sg13g2_buf_1 _12171_ (.A(_01677_),
    .X(_04445_));
 sg13g2_nor2_1 _12172_ (.A(_04434_),
    .B(_04440_),
    .Y(_04446_));
 sg13g2_buf_2 _12173_ (.A(_04446_),
    .X(_04447_));
 sg13g2_a21oi_1 _12174_ (.A1(_04434_),
    .A2(_04440_),
    .Y(_04448_),
    .B1(\clock_inst.min_a[23] ));
 sg13g2_buf_2 _12175_ (.A(_04448_),
    .X(_04449_));
 sg13g2_nor2_2 _12176_ (.A(_04447_),
    .B(_04449_),
    .Y(_04450_));
 sg13g2_xnor2_1 _12177_ (.Y(_04451_),
    .A(net531),
    .B(_04450_));
 sg13g2_nor2_1 _12178_ (.A(_04445_),
    .B(_04451_),
    .Y(_04452_));
 sg13g2_xnor2_1 _12179_ (.Y(_04453_),
    .A(net564),
    .B(_04452_));
 sg13g2_a21oi_1 _12180_ (.A1(net65),
    .A2(_04453_),
    .Y(_00378_),
    .B1(_03902_));
 sg13g2_buf_2 _12181_ (.A(\clock_inst.min_tile.e[25] ),
    .X(_04454_));
 sg13g2_or2_1 _12182_ (.X(_04455_),
    .B(_04449_),
    .A(_04447_));
 sg13g2_buf_2 _12183_ (.A(_04455_),
    .X(_04456_));
 sg13g2_nor2_1 _12184_ (.A(net479),
    .B(net564),
    .Y(_04457_));
 sg13g2_nand2_1 _12185_ (.Y(_04458_),
    .A(_04456_),
    .B(_04457_));
 sg13g2_inv_1 _12186_ (.Y(_04459_),
    .A(net564));
 sg13g2_nor2_1 _12187_ (.A(net568),
    .B(_04459_),
    .Y(_04460_));
 sg13g2_nand2_1 _12188_ (.Y(_04461_),
    .A(_04450_),
    .B(_04460_));
 sg13g2_a21oi_1 _12189_ (.A1(_04458_),
    .A2(_04461_),
    .Y(_04462_),
    .B1(_01743_));
 sg13g2_xnor2_1 _12190_ (.Y(_04463_),
    .A(_04454_),
    .B(_04462_));
 sg13g2_a21oi_1 _12191_ (.A1(net65),
    .A2(_04463_),
    .Y(_00379_),
    .B1(_03910_));
 sg13g2_buf_1 _12192_ (.A(\clock_inst.min_tile.e[26] ),
    .X(_04464_));
 sg13g2_inv_1 _12193_ (.Y(_04465_),
    .A(_04454_));
 sg13g2_nor4_1 _12194_ (.A(net531),
    .B(_04459_),
    .C(_04465_),
    .D(_04456_),
    .Y(_04466_));
 sg13g2_o21ai_1 _12195_ (.B1(_04465_),
    .Y(_04467_),
    .A1(_04447_),
    .A2(_04449_));
 sg13g2_buf_2 _12196_ (.A(_04467_),
    .X(_04468_));
 sg13g2_nor3_1 _12197_ (.A(net479),
    .B(net564),
    .C(_04468_),
    .Y(_04469_));
 sg13g2_o21ai_1 _12198_ (.B1(_02061_),
    .Y(_04470_),
    .A1(_04466_),
    .A2(_04469_));
 sg13g2_xor2_1 _12199_ (.B(_04470_),
    .A(net563),
    .X(_04471_));
 sg13g2_xnor2_1 _12200_ (.Y(_04472_),
    .A(_03920_),
    .B(_03915_));
 sg13g2_nand2_1 _12201_ (.Y(_04473_),
    .A(_01573_),
    .B(_04472_));
 sg13g2_a21oi_1 _12202_ (.A1(\clock_inst.min_c[26] ),
    .A2(_01925_),
    .Y(_04474_),
    .B1(_01926_));
 sg13g2_a22oi_1 _12203_ (.Y(_00380_),
    .B1(_04473_),
    .B2(_04474_),
    .A2(_04471_),
    .A1(_01914_));
 sg13g2_buf_1 _12204_ (.A(\clock_inst.min_tile.e[27] ),
    .X(_04475_));
 sg13g2_nor3_1 _12205_ (.A(net564),
    .B(_04454_),
    .C(net563),
    .Y(_04476_));
 sg13g2_o21ai_1 _12206_ (.B1(_04476_),
    .Y(_04477_),
    .A1(_04447_),
    .A2(_04449_));
 sg13g2_buf_1 _12207_ (.A(_04477_),
    .X(_04478_));
 sg13g2_nand2_1 _12208_ (.Y(_04479_),
    .A(net531),
    .B(net445));
 sg13g2_nand2_2 _12209_ (.Y(_04480_),
    .A(_04454_),
    .B(net563));
 sg13g2_nor4_1 _12210_ (.A(_04459_),
    .B(_04447_),
    .C(_04449_),
    .D(_04480_),
    .Y(_04481_));
 sg13g2_nand3_1 _12211_ (.B(net445),
    .C(_04481_),
    .A(net479),
    .Y(_04482_));
 sg13g2_o21ai_1 _12212_ (.B1(_04482_),
    .Y(_04483_),
    .A1(_04478_),
    .A2(_04479_));
 sg13g2_xor2_1 _12213_ (.B(_04483_),
    .A(net562),
    .X(_04484_));
 sg13g2_mux2_1 _12214_ (.A0(_03929_),
    .A1(_04484_),
    .S(_01913_),
    .X(_00381_));
 sg13g2_buf_2 _12215_ (.A(\clock_inst.min_tile.e[28] ),
    .X(_04485_));
 sg13g2_nand3b_1 _12216_ (.B(net500),
    .C(net531),
    .Y(_04486_),
    .A_N(net562));
 sg13g2_nand4_1 _12217_ (.B(net564),
    .C(net562),
    .A(net479),
    .Y(_04487_),
    .D(_01727_));
 sg13g2_or4_1 _12218_ (.A(_04447_),
    .B(_04449_),
    .C(_04480_),
    .D(_04487_),
    .X(_04488_));
 sg13g2_o21ai_1 _12219_ (.B1(_04488_),
    .Y(_04489_),
    .A1(_04478_),
    .A2(_04486_));
 sg13g2_xor2_1 _12220_ (.B(_04489_),
    .A(_04485_),
    .X(_04490_));
 sg13g2_nor2_1 _12221_ (.A(_01641_),
    .B(_04490_),
    .Y(_04491_));
 sg13g2_nor4_1 _12222_ (.A(_03938_),
    .B(_03939_),
    .C(_03940_),
    .D(_04491_),
    .Y(_00382_));
 sg13g2_buf_2 _12223_ (.A(\clock_inst.min_tile.e[29] ),
    .X(_04492_));
 sg13g2_nand3_1 _12224_ (.B(_04485_),
    .C(_04460_),
    .A(net562),
    .Y(_04493_));
 sg13g2_nor3_1 _12225_ (.A(_04456_),
    .B(_04480_),
    .C(_04493_),
    .Y(_04494_));
 sg13g2_or4_1 _12226_ (.A(net564),
    .B(_04454_),
    .C(net563),
    .D(_04485_),
    .X(_04495_));
 sg13g2_nor4_1 _12227_ (.A(net479),
    .B(net562),
    .C(_04450_),
    .D(_04495_),
    .Y(_04496_));
 sg13g2_o21ai_1 _12228_ (.B1(net355),
    .Y(_04497_),
    .A1(_04494_),
    .A2(_04496_));
 sg13g2_xor2_1 _12229_ (.B(_04497_),
    .A(_04492_),
    .X(_04498_));
 sg13g2_a21oi_1 _12230_ (.A1(_04420_),
    .A2(_04498_),
    .Y(_00383_),
    .B1(_03951_));
 sg13g2_xnor2_1 _12231_ (.Y(_04499_),
    .A(_02537_),
    .B(_04277_));
 sg13g2_nand2_1 _12232_ (.Y(_04500_),
    .A(net357),
    .B(_04499_));
 sg13g2_xor2_1 _12233_ (.B(_04500_),
    .A(\clock_inst.min_tile.e[2] ),
    .X(_04501_));
 sg13g2_a21oi_1 _12234_ (.A1(net65),
    .A2(_04501_),
    .Y(_00384_),
    .B1(_03958_));
 sg13g2_buf_2 _12235_ (.A(\clock_inst.min_tile.e[30] ),
    .X(_04502_));
 sg13g2_nor4_1 _12236_ (.A(_04444_),
    .B(net563),
    .C(net562),
    .D(_04485_),
    .Y(_04503_));
 sg13g2_nand3b_1 _12237_ (.B(_04503_),
    .C(net568),
    .Y(_04504_),
    .A_N(_04492_));
 sg13g2_nor3_1 _12238_ (.A(_04454_),
    .B(net502),
    .C(_04504_),
    .Y(_04505_));
 sg13g2_and3_1 _12239_ (.X(_04506_),
    .A(net562),
    .B(_04485_),
    .C(_04460_));
 sg13g2_and4_1 _12240_ (.A(net563),
    .B(_04492_),
    .C(_04450_),
    .D(_04506_),
    .X(_04507_));
 sg13g2_nor2_1 _12241_ (.A(_04465_),
    .B(_01681_),
    .Y(_04508_));
 sg13g2_a22oi_1 _12242_ (.Y(_04509_),
    .B1(_04507_),
    .B2(_04508_),
    .A2(_04505_),
    .A1(_04456_));
 sg13g2_xor2_1 _12243_ (.B(_04509_),
    .A(_04502_),
    .X(_04510_));
 sg13g2_a21oi_1 _12244_ (.A1(\clock_inst.min_c[30] ),
    .A2(net47),
    .Y(_04511_),
    .B1(_02101_));
 sg13g2_xnor2_1 _12245_ (.Y(_04512_),
    .A(_03973_),
    .B(_03969_));
 sg13g2_nand2_1 _12246_ (.Y(_04513_),
    .A(net45),
    .B(_04512_));
 sg13g2_a22oi_1 _12247_ (.Y(_00385_),
    .B1(_04511_),
    .B2(_04513_),
    .A2(_04510_),
    .A1(_01914_));
 sg13g2_buf_2 _12248_ (.A(\clock_inst.min_tile.e[31] ),
    .X(_04514_));
 sg13g2_nand4_1 _12249_ (.B(_04485_),
    .C(_04492_),
    .A(net562),
    .Y(_04515_),
    .D(_04502_));
 sg13g2_nor2_1 _12250_ (.A(net568),
    .B(_04515_),
    .Y(_04516_));
 sg13g2_a221oi_1 _12251_ (.B2(_04476_),
    .C1(_04516_),
    .B1(_04456_),
    .A1(net479),
    .Y(_04517_),
    .A2(_04459_));
 sg13g2_nor2_1 _12252_ (.A(_04485_),
    .B(_04492_),
    .Y(_04518_));
 sg13g2_nor3_1 _12253_ (.A(_02568_),
    .B(\clock_inst.min_tile.e[27] ),
    .C(_04502_),
    .Y(_04519_));
 sg13g2_and2_1 _12254_ (.A(_04518_),
    .B(_04519_),
    .X(_04520_));
 sg13g2_buf_1 _12255_ (.A(_04520_),
    .X(_04521_));
 sg13g2_nor2_1 _12256_ (.A(_04478_),
    .B(_04521_),
    .Y(_04522_));
 sg13g2_o21ai_1 _12257_ (.B1(net445),
    .Y(_04523_),
    .A1(_04165_),
    .A2(_04481_));
 sg13g2_nor3_1 _12258_ (.A(_04517_),
    .B(_04522_),
    .C(_04523_),
    .Y(_04524_));
 sg13g2_xnor2_1 _12259_ (.Y(_04525_),
    .A(_04514_),
    .B(_04524_));
 sg13g2_a21oi_1 _12260_ (.A1(_04420_),
    .A2(_04525_),
    .Y(_00386_),
    .B1(_03981_));
 sg13g2_buf_1 _12261_ (.A(\clock_inst.min_tile.e[32] ),
    .X(_04526_));
 sg13g2_nand4_1 _12262_ (.B(_04502_),
    .C(_04514_),
    .A(_04492_),
    .Y(_04527_),
    .D(_04506_));
 sg13g2_nor3_1 _12263_ (.A(_04456_),
    .B(_04480_),
    .C(_04527_),
    .Y(_04528_));
 sg13g2_nor2_1 _12264_ (.A(net563),
    .B(_04475_),
    .Y(_04529_));
 sg13g2_nand3_1 _12265_ (.B(_04529_),
    .C(_04518_),
    .A(_04457_),
    .Y(_04530_));
 sg13g2_nor4_1 _12266_ (.A(_04502_),
    .B(_04514_),
    .C(_04468_),
    .D(_04530_),
    .Y(_04531_));
 sg13g2_o21ai_1 _12267_ (.B1(_01816_),
    .Y(_04532_),
    .A1(_04528_),
    .A2(_04531_));
 sg13g2_xnor2_1 _12268_ (.Y(_04533_),
    .A(_04526_),
    .B(_04532_));
 sg13g2_mux2_1 _12269_ (.A0(_03989_),
    .A1(_04533_),
    .S(_01913_),
    .X(_00387_));
 sg13g2_buf_1 _12270_ (.A(\clock_inst.min_tile.e[33] ),
    .X(_04534_));
 sg13g2_nor4_1 _12271_ (.A(_04492_),
    .B(_04502_),
    .C(_04514_),
    .D(_04526_),
    .Y(_04535_));
 sg13g2_nand2_1 _12272_ (.Y(_04536_),
    .A(net531),
    .B(_04535_));
 sg13g2_nor4_1 _12273_ (.A(_04475_),
    .B(_04450_),
    .C(_04495_),
    .D(_04536_),
    .Y(_04537_));
 sg13g2_nand4_1 _12274_ (.B(_04502_),
    .C(_04514_),
    .A(_04492_),
    .Y(_04538_),
    .D(_04526_));
 sg13g2_nor4_1 _12275_ (.A(_04456_),
    .B(_04480_),
    .C(_04493_),
    .D(_04538_),
    .Y(_04539_));
 sg13g2_or4_1 _12276_ (.A(_04534_),
    .B(_03999_),
    .C(_04537_),
    .D(_04539_),
    .X(_04540_));
 sg13g2_nand2b_1 _12277_ (.Y(_04541_),
    .B(_02073_),
    .A_N(_04534_));
 sg13g2_o21ai_1 _12278_ (.B1(_04541_),
    .Y(_04542_),
    .A1(_03997_),
    .A2(_04540_));
 sg13g2_and2_1 _12279_ (.A(_04534_),
    .B(net445),
    .X(_04543_));
 sg13g2_o21ai_1 _12280_ (.B1(_04543_),
    .Y(_04544_),
    .A1(_04537_),
    .A2(_04539_));
 sg13g2_a221oi_1 _12281_ (.B2(_01176_),
    .C1(_03997_),
    .B1(_04544_),
    .A1(\clock_inst.min_c[33] ),
    .Y(_04545_),
    .A2(_01611_));
 sg13g2_nor2_1 _12282_ (.A(_04542_),
    .B(_04545_),
    .Y(_00388_));
 sg13g2_buf_1 _12283_ (.A(\clock_inst.min_tile.e[34] ),
    .X(_04546_));
 sg13g2_and2_1 _12284_ (.A(_04546_),
    .B(_01816_),
    .X(_04547_));
 sg13g2_and3_1 _12285_ (.X(_04548_),
    .A(_04514_),
    .B(_04526_),
    .C(_04534_));
 sg13g2_nand3_1 _12286_ (.B(_04516_),
    .C(_04548_),
    .A(net563),
    .Y(_04549_));
 sg13g2_o21ai_1 _12287_ (.B1(_04454_),
    .Y(_04550_),
    .A1(_04434_),
    .A2(_04440_));
 sg13g2_o21ai_1 _12288_ (.B1(net479),
    .Y(_04551_),
    .A1(_04449_),
    .A2(_04550_));
 sg13g2_a22oi_1 _12289_ (.Y(_04552_),
    .B1(_04551_),
    .B2(net564),
    .A2(_04468_),
    .A1(net531));
 sg13g2_nor4_1 _12290_ (.A(_04502_),
    .B(_04514_),
    .C(_04526_),
    .D(_04534_),
    .Y(_04553_));
 sg13g2_nand2b_1 _12291_ (.Y(_04554_),
    .B(_04553_),
    .A_N(_04530_));
 sg13g2_a21o_1 _12292_ (.A2(_04468_),
    .A1(net531),
    .B1(_04554_),
    .X(_04555_));
 sg13g2_o21ai_1 _12293_ (.B1(_04555_),
    .Y(_04556_),
    .A1(_04549_),
    .A2(_04552_));
 sg13g2_a21o_1 _12294_ (.A2(_04556_),
    .A1(_04547_),
    .B1(net156),
    .X(_04557_));
 sg13g2_nor2_1 _12295_ (.A(_04002_),
    .B(net95),
    .Y(_04558_));
 sg13g2_nor2_1 _12296_ (.A(_04001_),
    .B(net95),
    .Y(_04559_));
 sg13g2_nand4_1 _12297_ (.B(_03889_),
    .C(_03903_),
    .A(_02959_),
    .Y(_04560_),
    .D(_04004_));
 sg13g2_nand2_1 _12298_ (.Y(_04561_),
    .A(_02959_),
    .B(_03911_));
 sg13g2_nand2_1 _12299_ (.Y(_04562_),
    .A(net566),
    .B(_03960_));
 sg13g2_o21ai_1 _12300_ (.B1(_04562_),
    .Y(_04563_),
    .A1(_03965_),
    .A2(_04561_));
 sg13g2_nand2b_1 _12301_ (.Y(_04564_),
    .B(_04563_),
    .A_N(_04560_));
 sg13g2_o21ai_1 _12302_ (.B1(_04008_),
    .Y(_04565_),
    .A1(_03896_),
    .A2(_04564_));
 sg13g2_mux2_1 _12303_ (.A0(_04558_),
    .A1(_04559_),
    .S(_04565_),
    .X(_04566_));
 sg13g2_nand2b_1 _12304_ (.Y(_04567_),
    .B(_04553_),
    .A_N(_04504_));
 sg13g2_a21oi_1 _12305_ (.A1(net531),
    .A2(_04468_),
    .Y(_04568_),
    .B1(_04567_));
 sg13g2_nor2_1 _12306_ (.A(_04459_),
    .B(_04549_),
    .Y(_04569_));
 sg13g2_and2_1 _12307_ (.A(_04551_),
    .B(_04569_),
    .X(_04570_));
 sg13g2_or4_1 _12308_ (.A(_04546_),
    .B(_03999_),
    .C(_04568_),
    .D(_04570_),
    .X(_04571_));
 sg13g2_nand2b_1 _12309_ (.Y(_04572_),
    .B(_02073_),
    .A_N(_04546_));
 sg13g2_o21ai_1 _12310_ (.B1(_04572_),
    .Y(_04573_),
    .A1(_04566_),
    .A2(_04571_));
 sg13g2_a21oi_1 _12311_ (.A1(_04011_),
    .A2(_04557_),
    .Y(_00389_),
    .B1(_04573_));
 sg13g2_nor4_1 _12312_ (.A(_04514_),
    .B(_04526_),
    .C(_04534_),
    .D(_04546_),
    .Y(_04574_));
 sg13g2_nand2_1 _12313_ (.Y(_04575_),
    .A(_02567_),
    .B(_04574_));
 sg13g2_nand4_1 _12314_ (.B(_04454_),
    .C(_04546_),
    .A(_02569_),
    .Y(_04576_),
    .D(_04548_));
 sg13g2_nor2_1 _12315_ (.A(_04516_),
    .B(_04521_),
    .Y(_04577_));
 sg13g2_a21oi_1 _12316_ (.A1(_04575_),
    .A2(_04576_),
    .Y(_04578_),
    .B1(_04577_));
 sg13g2_nand2_1 _12317_ (.Y(_04579_),
    .A(_04521_),
    .B(_04574_));
 sg13g2_a21oi_1 _12318_ (.A1(_04478_),
    .A2(_04578_),
    .Y(_04580_),
    .B1(_04579_));
 sg13g2_and4_1 _12319_ (.A(_04464_),
    .B(_04450_),
    .C(_04460_),
    .D(_04578_),
    .X(_04581_));
 sg13g2_or3_1 _12320_ (.A(\clock_inst.min_tile.e[35] ),
    .B(_04580_),
    .C(_04581_),
    .X(_04582_));
 sg13g2_nand2b_1 _12321_ (.Y(_04583_),
    .B(net137),
    .A_N(\clock_inst.min_tile.e[35] ));
 sg13g2_o21ai_1 _12322_ (.B1(_04583_),
    .Y(_04584_),
    .A1(_04023_),
    .A2(_04582_));
 sg13g2_and2_1 _12323_ (.A(\clock_inst.min_tile.e[35] ),
    .B(_01964_),
    .X(_04585_));
 sg13g2_o21ai_1 _12324_ (.B1(_04585_),
    .Y(_04586_),
    .A1(_04580_),
    .A2(_04581_));
 sg13g2_a21oi_1 _12325_ (.A1(net136),
    .A2(_04586_),
    .Y(_04587_),
    .B1(_04023_));
 sg13g2_nor2_1 _12326_ (.A(_04584_),
    .B(_04587_),
    .Y(_00390_));
 sg13g2_nand2_1 _12327_ (.Y(_04588_),
    .A(\clock_inst.min_a[36] ),
    .B(net355));
 sg13g2_xor2_1 _12328_ (.B(_04588_),
    .A(\clock_inst.min_tile.e[36] ),
    .X(_04589_));
 sg13g2_o21ai_1 _12329_ (.B1(_04029_),
    .Y(_00391_),
    .A1(net135),
    .A2(_04589_));
 sg13g2_buf_8 _12330_ (.A(\clock_inst.min_tile.e[37] ),
    .X(_04590_));
 sg13g2_nand2_1 _12331_ (.Y(_04591_),
    .A(\clock_inst.min_a[36] ),
    .B(\clock_inst.min_tile.e[36] ));
 sg13g2_xnor2_1 _12332_ (.Y(_04592_),
    .A(_02593_),
    .B(_04591_));
 sg13g2_nor2_1 _12333_ (.A(net406),
    .B(_04592_),
    .Y(_04593_));
 sg13g2_xnor2_1 _12334_ (.Y(_04594_),
    .A(_04590_),
    .B(_04593_));
 sg13g2_a21oi_1 _12335_ (.A1(net65),
    .A2(_04594_),
    .Y(_00392_),
    .B1(_04037_));
 sg13g2_buf_2 _12336_ (.A(\clock_inst.min_tile.e[38] ),
    .X(_04595_));
 sg13g2_nor2_1 _12337_ (.A(\clock_inst.min_a[37] ),
    .B(_04590_),
    .Y(_04596_));
 sg13g2_a22oi_1 _12338_ (.Y(_04597_),
    .B1(\clock_inst.min_a[37] ),
    .B2(_04590_),
    .A2(\clock_inst.min_tile.e[36] ),
    .A1(\clock_inst.min_a[36] ));
 sg13g2_nor2_1 _12339_ (.A(_04596_),
    .B(_04597_),
    .Y(_04598_));
 sg13g2_xnor2_1 _12340_ (.Y(_04599_),
    .A(_02630_),
    .B(_04598_));
 sg13g2_nor2_1 _12341_ (.A(net406),
    .B(_04599_),
    .Y(_04600_));
 sg13g2_xnor2_1 _12342_ (.Y(_04601_),
    .A(_04595_),
    .B(_04600_));
 sg13g2_a21oi_1 _12343_ (.A1(net65),
    .A2(_04601_),
    .Y(_00393_),
    .B1(_04047_));
 sg13g2_buf_1 _12344_ (.A(net140),
    .X(_04602_));
 sg13g2_or2_1 _12345_ (.X(_04603_),
    .B(_04595_),
    .A(_02630_));
 sg13g2_and2_1 _12346_ (.A(_02630_),
    .B(_04595_),
    .X(_04604_));
 sg13g2_a21oi_1 _12347_ (.A1(_04598_),
    .A2(_04603_),
    .Y(_04605_),
    .B1(_04604_));
 sg13g2_xnor2_1 _12348_ (.Y(_04606_),
    .A(_02654_),
    .B(_04605_));
 sg13g2_nand2_1 _12349_ (.Y(_04607_),
    .A(net357),
    .B(_04606_));
 sg13g2_xor2_1 _12350_ (.B(_04607_),
    .A(\clock_inst.min_tile.e[39] ),
    .X(_04608_));
 sg13g2_a21oi_1 _12351_ (.A1(net64),
    .A2(_04608_),
    .Y(_00394_),
    .B1(_04057_));
 sg13g2_xnor2_1 _12352_ (.Y(_04609_),
    .A(_02656_),
    .B(_04280_));
 sg13g2_nor2_1 _12353_ (.A(net406),
    .B(_04609_),
    .Y(_04610_));
 sg13g2_xnor2_1 _12354_ (.Y(_04611_),
    .A(_04270_),
    .B(_04610_));
 sg13g2_a21oi_1 _12355_ (.A1(net64),
    .A2(_04611_),
    .Y(_00395_),
    .B1(_04063_));
 sg13g2_a22oi_1 _12356_ (.Y(_04612_),
    .B1(_02630_),
    .B2(_04595_),
    .A2(_04590_),
    .A1(\clock_inst.min_a[37] ));
 sg13g2_o21ai_1 _12357_ (.B1(_04612_),
    .Y(_04613_),
    .A1(_04591_),
    .A2(_04596_));
 sg13g2_buf_1 _12358_ (.A(_04613_),
    .X(_04614_));
 sg13g2_and2_1 _12359_ (.A(\clock_inst.min_tile.e[39] ),
    .B(_04603_),
    .X(_04615_));
 sg13g2_buf_1 _12360_ (.A(_04615_),
    .X(_04616_));
 sg13g2_o21ai_1 _12361_ (.B1(_02654_),
    .Y(_04617_),
    .A1(_02630_),
    .A2(_04595_));
 sg13g2_nor3_1 _12362_ (.A(_04596_),
    .B(_04597_),
    .C(_04617_),
    .Y(_04618_));
 sg13g2_o21ai_1 _12363_ (.B1(_02654_),
    .Y(_04619_),
    .A1(\clock_inst.min_tile.e[39] ),
    .A2(_04604_));
 sg13g2_nand2b_1 _12364_ (.Y(_04620_),
    .B(_04619_),
    .A_N(_04618_));
 sg13g2_a21o_1 _12365_ (.A2(_04616_),
    .A1(_04614_),
    .B1(_04620_),
    .X(_04621_));
 sg13g2_xnor2_1 _12366_ (.Y(_04622_),
    .A(_02698_),
    .B(_04621_));
 sg13g2_nor2_1 _12367_ (.A(net406),
    .B(_04622_),
    .Y(_04623_));
 sg13g2_xnor2_1 _12368_ (.Y(_04624_),
    .A(\clock_inst.min_tile.e[40] ),
    .B(_04623_));
 sg13g2_a21oi_1 _12369_ (.A1(net64),
    .A2(_04624_),
    .Y(_00396_),
    .B1(_04076_));
 sg13g2_buf_1 _12370_ (.A(\clock_inst.min_tile.e[41] ),
    .X(_04625_));
 sg13g2_nand2_1 _12371_ (.Y(_04626_),
    .A(_02698_),
    .B(\clock_inst.min_tile.e[40] ));
 sg13g2_or2_1 _12372_ (.X(_04627_),
    .B(\clock_inst.min_tile.e[40] ),
    .A(_02698_));
 sg13g2_nand2_1 _12373_ (.Y(_04628_),
    .A(_04621_),
    .B(_04627_));
 sg13g2_and2_1 _12374_ (.A(_04626_),
    .B(_04628_),
    .X(_04629_));
 sg13g2_xor2_1 _12375_ (.B(_04629_),
    .A(_02714_),
    .X(_04630_));
 sg13g2_nor2_1 _12376_ (.A(net406),
    .B(_04630_),
    .Y(_04631_));
 sg13g2_xnor2_1 _12377_ (.Y(_04632_),
    .A(_04625_),
    .B(_04631_));
 sg13g2_a21oi_1 _12378_ (.A1(_04602_),
    .A2(_04632_),
    .Y(_00397_),
    .B1(_04095_));
 sg13g2_buf_2 _12379_ (.A(\clock_inst.min_tile.e[42] ),
    .X(_04633_));
 sg13g2_nand2b_1 _12380_ (.Y(_04634_),
    .B(_04626_),
    .A_N(_04625_));
 sg13g2_nand2b_1 _12381_ (.Y(_04635_),
    .B(_04626_),
    .A_N(_02714_));
 sg13g2_a221oi_1 _12382_ (.B2(_04635_),
    .C1(_04620_),
    .B1(_04634_),
    .A1(_04614_),
    .Y(_04636_),
    .A2(_04616_));
 sg13g2_buf_1 _12383_ (.A(_04636_),
    .X(_04637_));
 sg13g2_nor2_1 _12384_ (.A(_02714_),
    .B(_04625_),
    .Y(_04638_));
 sg13g2_a21oi_1 _12385_ (.A1(_02714_),
    .A2(_04625_),
    .Y(_04639_),
    .B1(_04627_));
 sg13g2_or2_1 _12386_ (.X(_04640_),
    .B(_04639_),
    .A(_04638_));
 sg13g2_buf_1 _12387_ (.A(_04640_),
    .X(_04641_));
 sg13g2_nor2_1 _12388_ (.A(_04637_),
    .B(_04641_),
    .Y(_04642_));
 sg13g2_xnor2_1 _12389_ (.Y(_04643_),
    .A(_02735_),
    .B(_04642_));
 sg13g2_nor2_1 _12390_ (.A(net406),
    .B(_04643_),
    .Y(_04644_));
 sg13g2_xnor2_1 _12391_ (.Y(_04645_),
    .A(_04633_),
    .B(_04644_));
 sg13g2_a21oi_1 _12392_ (.A1(net64),
    .A2(_04645_),
    .Y(_00398_),
    .B1(_04105_));
 sg13g2_buf_1 _12393_ (.A(\clock_inst.min_tile.e[43] ),
    .X(_04646_));
 sg13g2_nor2_1 _12394_ (.A(_04633_),
    .B(_04642_),
    .Y(_04647_));
 sg13g2_a21oi_1 _12395_ (.A1(_04633_),
    .A2(_04642_),
    .Y(_04648_),
    .B1(_02735_));
 sg13g2_o21ai_1 _12396_ (.B1(_02738_),
    .Y(_04649_),
    .A1(_04647_),
    .A2(_04648_));
 sg13g2_or3_1 _12397_ (.A(_02738_),
    .B(_04647_),
    .C(_04648_),
    .X(_04650_));
 sg13g2_a21oi_1 _12398_ (.A1(_04649_),
    .A2(_04650_),
    .Y(_04651_),
    .B1(net446));
 sg13g2_xnor2_1 _12399_ (.Y(_04652_),
    .A(_04646_),
    .B(_04651_));
 sg13g2_o21ai_1 _12400_ (.B1(_04122_),
    .Y(_00399_),
    .A1(_02131_),
    .A2(_04652_));
 sg13g2_buf_2 _12401_ (.A(\clock_inst.min_tile.e[44] ),
    .X(_04653_));
 sg13g2_inv_1 _12402_ (.Y(_04654_),
    .A(_02763_));
 sg13g2_nand2_1 _12403_ (.Y(_04655_),
    .A(_02738_),
    .B(_04646_));
 sg13g2_buf_2 _12404_ (.A(_04655_),
    .X(_04656_));
 sg13g2_or2_1 _12405_ (.X(_04657_),
    .B(_04646_),
    .A(_02738_));
 sg13g2_buf_1 _12406_ (.A(_04657_),
    .X(_04658_));
 sg13g2_nand3_1 _12407_ (.B(_04633_),
    .C(_04658_),
    .A(_02735_),
    .Y(_04659_));
 sg13g2_nand2_1 _12408_ (.Y(_04660_),
    .A(_04656_),
    .B(_04659_));
 sg13g2_nor2_1 _12409_ (.A(_02738_),
    .B(_04646_),
    .Y(_04661_));
 sg13g2_nor2_1 _12410_ (.A(_02735_),
    .B(_04633_),
    .Y(_04662_));
 sg13g2_nor4_1 _12411_ (.A(_04637_),
    .B(_04641_),
    .C(_04661_),
    .D(_04662_),
    .Y(_04663_));
 sg13g2_nor2_1 _12412_ (.A(_04660_),
    .B(_04663_),
    .Y(_04664_));
 sg13g2_xnor2_1 _12413_ (.Y(_04665_),
    .A(_04654_),
    .B(_04664_));
 sg13g2_nor2_1 _12414_ (.A(_04445_),
    .B(_04665_),
    .Y(_04666_));
 sg13g2_xnor2_1 _12415_ (.Y(_04667_),
    .A(_04653_),
    .B(_04666_));
 sg13g2_a21oi_1 _12416_ (.A1(net64),
    .A2(_04667_),
    .Y(_00400_),
    .B1(_04132_));
 sg13g2_buf_2 _12417_ (.A(\clock_inst.min_tile.e[45] ),
    .X(_04668_));
 sg13g2_o21ai_1 _12418_ (.B1(_04653_),
    .Y(_04669_),
    .A1(_04660_),
    .A2(_04663_));
 sg13g2_buf_2 _12419_ (.A(_04669_),
    .X(_04670_));
 sg13g2_a21oi_1 _12420_ (.A1(_04614_),
    .A2(_04616_),
    .Y(_04671_),
    .B1(_04634_));
 sg13g2_a21oi_1 _12421_ (.A1(_04614_),
    .A2(_04616_),
    .Y(_04672_),
    .B1(_04635_));
 sg13g2_nor2b_1 _12422_ (.A(_04618_),
    .B_N(_04619_),
    .Y(_04673_));
 sg13g2_o21ai_1 _12423_ (.B1(_04673_),
    .Y(_04674_),
    .A1(_04671_),
    .A2(_04672_));
 sg13g2_nor2_1 _12424_ (.A(_04638_),
    .B(_04639_),
    .Y(_04675_));
 sg13g2_inv_1 _12425_ (.Y(_04676_),
    .A(_04633_));
 sg13g2_inv_1 _12426_ (.Y(_04677_),
    .A(_04653_));
 sg13g2_nand3_1 _12427_ (.B(_04677_),
    .C(_04656_),
    .A(_04676_),
    .Y(_04678_));
 sg13g2_nand3b_1 _12428_ (.B(_04677_),
    .C(_04656_),
    .Y(_04679_),
    .A_N(_02735_));
 sg13g2_a22oi_1 _12429_ (.Y(_04680_),
    .B1(_04678_),
    .B2(_04679_),
    .A2(_04675_),
    .A1(_04674_));
 sg13g2_nand2_1 _12430_ (.Y(_04681_),
    .A(_04656_),
    .B(_04662_));
 sg13g2_a21oi_1 _12431_ (.A1(_04658_),
    .A2(_04681_),
    .Y(_04682_),
    .B1(_04653_));
 sg13g2_or3_1 _12432_ (.A(_04654_),
    .B(_04680_),
    .C(_04682_),
    .X(_04683_));
 sg13g2_buf_2 _12433_ (.A(_04683_),
    .X(_04684_));
 sg13g2_nand2_2 _12434_ (.Y(_04685_),
    .A(_04670_),
    .B(_04684_));
 sg13g2_xnor2_1 _12435_ (.Y(_04686_),
    .A(net533),
    .B(_04685_));
 sg13g2_or3_1 _12436_ (.A(_04668_),
    .B(net233),
    .C(_04686_),
    .X(_04687_));
 sg13g2_nand4_1 _12437_ (.B(net153),
    .C(net356),
    .A(_04668_),
    .Y(_04688_),
    .D(_04686_));
 sg13g2_nor3_1 _12438_ (.A(_04668_),
    .B(net240),
    .C(net356),
    .Y(_04689_));
 sg13g2_nor2_1 _12439_ (.A(_04153_),
    .B(_04689_),
    .Y(_04690_));
 sg13g2_and3_1 _12440_ (.X(_00401_),
    .A(_04687_),
    .B(_04688_),
    .C(_04690_));
 sg13g2_buf_1 _12441_ (.A(\clock_inst.min_tile.e[46] ),
    .X(_04691_));
 sg13g2_nor2_1 _12442_ (.A(net533),
    .B(_04668_),
    .Y(_04692_));
 sg13g2_nand2_1 _12443_ (.Y(_04693_),
    .A(net445),
    .B(_04692_));
 sg13g2_nand3_1 _12444_ (.B(_04668_),
    .C(net499),
    .A(net533),
    .Y(_04694_));
 sg13g2_mux2_1 _12445_ (.A0(_04693_),
    .A1(_04694_),
    .S(_04685_),
    .X(_04695_));
 sg13g2_xor2_1 _12446_ (.B(_04695_),
    .A(_04691_),
    .X(_04696_));
 sg13g2_a21oi_1 _12447_ (.A1(net64),
    .A2(_04696_),
    .Y(_00402_),
    .B1(_04160_));
 sg13g2_buf_1 _12448_ (.A(\clock_inst.min_tile.e[47] ),
    .X(_04697_));
 sg13g2_and3_1 _12449_ (.X(_04698_),
    .A(_04697_),
    .B(net239),
    .C(net443));
 sg13g2_nor2_1 _12450_ (.A(_04697_),
    .B(net240),
    .Y(_04699_));
 sg13g2_nand2b_1 _12451_ (.Y(_04700_),
    .B(_04692_),
    .A_N(_04691_));
 sg13g2_nand3_1 _12452_ (.B(_04668_),
    .C(_04691_),
    .A(net533),
    .Y(_04701_));
 sg13g2_mux2_1 _12453_ (.A0(_04700_),
    .A1(_04701_),
    .S(_04685_),
    .X(_04702_));
 sg13g2_mux2_1 _12454_ (.A0(_04698_),
    .A1(_04699_),
    .S(_04702_),
    .X(_04703_));
 sg13g2_nor3_1 _12455_ (.A(_04697_),
    .B(net142),
    .C(net356),
    .Y(_04704_));
 sg13g2_nor3_1 _12456_ (.A(_04170_),
    .B(_04703_),
    .C(_04704_),
    .Y(_00403_));
 sg13g2_buf_1 _12457_ (.A(\clock_inst.min_tile.e[48] ),
    .X(_04705_));
 sg13g2_nor2_1 _12458_ (.A(_04661_),
    .B(_04662_),
    .Y(_04706_));
 sg13g2_nor3_1 _12459_ (.A(_04668_),
    .B(_04691_),
    .C(_04697_),
    .Y(_04707_));
 sg13g2_nand2_1 _12460_ (.Y(_04708_),
    .A(_02781_),
    .B(_04707_));
 sg13g2_nand3_1 _12461_ (.B(_04691_),
    .C(_04697_),
    .A(_04668_),
    .Y(_04709_));
 sg13g2_nand2b_1 _12462_ (.Y(_04710_),
    .B(net533),
    .A_N(_04709_));
 sg13g2_xnor2_1 _12463_ (.Y(_04711_),
    .A(_02763_),
    .B(_04653_));
 sg13g2_a21oi_1 _12464_ (.A1(_04708_),
    .A2(_04710_),
    .Y(_04712_),
    .B1(_04711_));
 sg13g2_nand4_1 _12465_ (.B(_04675_),
    .C(_04706_),
    .A(_04674_),
    .Y(_04713_),
    .D(_04712_));
 sg13g2_nand2_1 _12466_ (.Y(_04714_),
    .A(net533),
    .B(_04709_));
 sg13g2_nand2_1 _12467_ (.Y(_04715_),
    .A(_02763_),
    .B(_04653_));
 sg13g2_o21ai_1 _12468_ (.B1(_04715_),
    .Y(_04716_),
    .A1(_02782_),
    .A2(_04707_));
 sg13g2_a22oi_1 _12469_ (.Y(_04717_),
    .B1(_04712_),
    .B2(_04660_),
    .A2(_04716_),
    .A1(_04714_));
 sg13g2_a21oi_2 _12470_ (.B1(_02781_),
    .Y(_04718_),
    .A2(_04717_),
    .A1(_04713_));
 sg13g2_and3_1 _12471_ (.X(_04719_),
    .A(_02781_),
    .B(_04713_),
    .C(_04717_));
 sg13g2_o21ai_1 _12472_ (.B1(net355),
    .Y(_04720_),
    .A1(_04718_),
    .A2(_04719_));
 sg13g2_xor2_1 _12473_ (.B(_04720_),
    .A(_04705_),
    .X(_04721_));
 sg13g2_xnor2_1 _12474_ (.Y(_04722_),
    .A(_04178_),
    .B(_04174_));
 sg13g2_nand2_1 _12475_ (.Y(_04723_),
    .A(net45),
    .B(_04722_));
 sg13g2_a21oi_1 _12476_ (.A1(\clock_inst.min_c[48] ),
    .A2(net43),
    .Y(_04724_),
    .B1(net138));
 sg13g2_a22oi_1 _12477_ (.Y(_00404_),
    .B1(_04723_),
    .B2(_04724_),
    .A2(_04721_),
    .A1(net75));
 sg13g2_buf_1 _12478_ (.A(\clock_inst.min_tile.e[49] ),
    .X(_04725_));
 sg13g2_nor2_1 _12479_ (.A(_04705_),
    .B(_04708_),
    .Y(_04726_));
 sg13g2_nand3_1 _12480_ (.B(_04684_),
    .C(_04726_),
    .A(_04670_),
    .Y(_04727_));
 sg13g2_nand2_1 _12481_ (.Y(_04728_),
    .A(_04705_),
    .B(_04718_));
 sg13g2_a21oi_1 _12482_ (.A1(_04727_),
    .A2(_04728_),
    .Y(_04729_),
    .B1(net447));
 sg13g2_xnor2_1 _12483_ (.Y(_04730_),
    .A(_04725_),
    .B(_04729_));
 sg13g2_xnor2_1 _12484_ (.Y(_04731_),
    .A(_04179_),
    .B(_04183_));
 sg13g2_nand2_1 _12485_ (.Y(_04732_),
    .A(\clock_inst.min_c[49] ),
    .B(net107));
 sg13g2_o21ai_1 _12486_ (.B1(_04732_),
    .Y(_04733_),
    .A1(net98),
    .A2(_04731_));
 sg13g2_nor2_1 _12487_ (.A(net83),
    .B(_04733_),
    .Y(_04734_));
 sg13g2_a21oi_1 _12488_ (.A1(_04602_),
    .A2(_04730_),
    .Y(_00405_),
    .B1(_04734_));
 sg13g2_xnor2_1 _12489_ (.Y(_04735_),
    .A(_02765_),
    .B(_04283_));
 sg13g2_nor2_1 _12490_ (.A(net406),
    .B(_04735_),
    .Y(_04736_));
 sg13g2_xnor2_1 _12491_ (.Y(_04737_),
    .A(_04284_),
    .B(_04736_));
 sg13g2_a21oi_1 _12492_ (.A1(net64),
    .A2(_04737_),
    .Y(_00406_),
    .B1(_04194_));
 sg13g2_nand3_1 _12493_ (.B(_04653_),
    .C(_04658_),
    .A(_04633_),
    .Y(_04738_));
 sg13g2_nor3_1 _12494_ (.A(_04637_),
    .B(_04641_),
    .C(_04738_),
    .Y(_04739_));
 sg13g2_nand3_1 _12495_ (.B(_04653_),
    .C(_04658_),
    .A(_02735_),
    .Y(_04740_));
 sg13g2_nor3_1 _12496_ (.A(_04637_),
    .B(_04641_),
    .C(_04740_),
    .Y(_04741_));
 sg13g2_a21oi_1 _12497_ (.A1(_04656_),
    .A2(_04659_),
    .Y(_04742_),
    .B1(_04677_));
 sg13g2_nand2b_1 _12498_ (.Y(_04743_),
    .B(_04726_),
    .A_N(_04725_));
 sg13g2_nor4_1 _12499_ (.A(_04739_),
    .B(_04741_),
    .C(_04742_),
    .D(_04743_),
    .Y(_04744_));
 sg13g2_nand2_1 _12500_ (.Y(_04745_),
    .A(_04705_),
    .B(_04725_));
 sg13g2_or2_1 _12501_ (.X(_04746_),
    .B(_04745_),
    .A(_04710_));
 sg13g2_nor2_1 _12502_ (.A(_04654_),
    .B(_04746_),
    .Y(_04747_));
 sg13g2_nor2_1 _12503_ (.A(_04680_),
    .B(_04682_),
    .Y(_04748_));
 sg13g2_nand2_1 _12504_ (.Y(_04749_),
    .A(_04676_),
    .B(_04656_));
 sg13g2_nand2b_1 _12505_ (.Y(_04750_),
    .B(_04656_),
    .A_N(_02735_));
 sg13g2_a22oi_1 _12506_ (.Y(_04751_),
    .B1(_04749_),
    .B2(_04750_),
    .A2(_04675_),
    .A1(_04674_));
 sg13g2_nand2_1 _12507_ (.Y(_04752_),
    .A(_04658_),
    .B(_04681_));
 sg13g2_nor4_1 _12508_ (.A(_04677_),
    .B(_04751_),
    .C(_04752_),
    .D(_04746_),
    .Y(_04753_));
 sg13g2_a221oi_1 _12509_ (.B2(_04748_),
    .C1(_04753_),
    .B1(_04747_),
    .A1(_04684_),
    .Y(_04754_),
    .A2(_04744_));
 sg13g2_buf_1 _12510_ (.A(\clock_inst.min_tile.e[50] ),
    .X(_04755_));
 sg13g2_nand2_1 _12511_ (.Y(_04756_),
    .A(_04755_),
    .B(net356));
 sg13g2_o21ai_1 _12512_ (.B1(net145),
    .Y(_04757_),
    .A1(_04754_),
    .A2(_04756_));
 sg13g2_a21oi_1 _12513_ (.A1(_04216_),
    .A2(_04754_),
    .Y(_04758_),
    .B1(net137));
 sg13g2_nor2_1 _12514_ (.A(_04755_),
    .B(_04758_),
    .Y(_04759_));
 sg13g2_a21oi_1 _12515_ (.A1(_04216_),
    .A2(_04757_),
    .Y(_00407_),
    .B1(_04759_));
 sg13g2_xnor2_1 _12516_ (.Y(_04760_),
    .A(_04217_),
    .B(_04219_));
 sg13g2_nand2_1 _12517_ (.Y(_04761_),
    .A(\clock_inst.min_c[51] ),
    .B(net96));
 sg13g2_o21ai_1 _12518_ (.B1(_04761_),
    .Y(_04762_),
    .A1(net48),
    .A2(_04760_));
 sg13g2_buf_1 _12519_ (.A(\clock_inst.min_tile.e[51] ),
    .X(_04763_));
 sg13g2_and3_1 _12520_ (.X(_04764_),
    .A(_04705_),
    .B(_04725_),
    .C(_04755_));
 sg13g2_buf_1 _12521_ (.A(_04764_),
    .X(_04765_));
 sg13g2_nand2_1 _12522_ (.Y(_04766_),
    .A(_04718_),
    .B(_04765_));
 sg13g2_nor2_1 _12523_ (.A(_04725_),
    .B(_04755_),
    .Y(_04767_));
 sg13g2_nand4_1 _12524_ (.B(_04684_),
    .C(_04726_),
    .A(_04670_),
    .Y(_04768_),
    .D(_04767_));
 sg13g2_a21oi_1 _12525_ (.A1(_04766_),
    .A2(_04768_),
    .Y(_04769_),
    .B1(net501));
 sg13g2_xor2_1 _12526_ (.B(_04769_),
    .A(_04763_),
    .X(_04770_));
 sg13g2_mux2_1 _12527_ (.A0(_04762_),
    .A1(_04770_),
    .S(net76),
    .X(_00408_));
 sg13g2_nor3_1 _12528_ (.A(_04725_),
    .B(_04755_),
    .C(_04763_),
    .Y(_04771_));
 sg13g2_nor2_1 _12529_ (.A(net533),
    .B(_04705_),
    .Y(_04772_));
 sg13g2_nand4_1 _12530_ (.B(_04717_),
    .C(_04771_),
    .A(_04713_),
    .Y(_04773_),
    .D(_04772_));
 sg13g2_nand3_1 _12531_ (.B(_04718_),
    .C(_04765_),
    .A(_04763_),
    .Y(_04774_));
 sg13g2_a21o_1 _12532_ (.A2(_04774_),
    .A1(_04773_),
    .B1(net446),
    .X(_04775_));
 sg13g2_xor2_1 _12533_ (.B(_04775_),
    .A(\clock_inst.min_tile.e[52] ),
    .X(_04776_));
 sg13g2_a22oi_1 _12534_ (.Y(_00409_),
    .B1(_04776_),
    .B2(net78),
    .A2(_04228_),
    .A1(_04227_));
 sg13g2_nor2b_1 _12535_ (.A(\clock_inst.min_tile.e[52] ),
    .B_N(_04771_),
    .Y(_04777_));
 sg13g2_nand4_1 _12536_ (.B(_04684_),
    .C(_04726_),
    .A(_04670_),
    .Y(_04778_),
    .D(_04777_));
 sg13g2_nand4_1 _12537_ (.B(\clock_inst.min_tile.e[52] ),
    .C(_04718_),
    .A(_04763_),
    .Y(_04779_),
    .D(_04765_));
 sg13g2_nand2_1 _12538_ (.Y(_04780_),
    .A(_04778_),
    .B(_04779_));
 sg13g2_nor3_1 _12539_ (.A(\clock_inst.min_tile.e[53] ),
    .B(_04236_),
    .C(_04780_),
    .Y(_04781_));
 sg13g2_nor2_1 _12540_ (.A(\clock_inst.min_tile.e[53] ),
    .B(net80),
    .Y(_04782_));
 sg13g2_nand2_1 _12541_ (.Y(_04783_),
    .A(\clock_inst.min_tile.e[53] ),
    .B(net442));
 sg13g2_a21o_1 _12542_ (.A2(_04779_),
    .A1(_04778_),
    .B1(_04783_),
    .X(_04784_));
 sg13g2_a21oi_1 _12543_ (.A1(net160),
    .A2(_04784_),
    .Y(_04785_),
    .B1(_04236_));
 sg13g2_nor3_1 _12544_ (.A(_04781_),
    .B(_04782_),
    .C(_04785_),
    .Y(_00410_));
 sg13g2_o21ai_1 _12545_ (.B1(_02765_),
    .Y(_04786_),
    .A1(_04284_),
    .A2(_04283_));
 sg13g2_nand2_1 _12546_ (.Y(_04787_),
    .A(_04284_),
    .B(_04283_));
 sg13g2_nand2_1 _12547_ (.Y(_04788_),
    .A(_04786_),
    .B(_04787_));
 sg13g2_xnor2_1 _12548_ (.Y(_04789_),
    .A(_02788_),
    .B(_04788_));
 sg13g2_nor2_1 _12549_ (.A(net406),
    .B(_04789_),
    .Y(_04790_));
 sg13g2_xnor2_1 _12550_ (.Y(_04791_),
    .A(\clock_inst.min_tile.e[5] ),
    .B(_04790_));
 sg13g2_a21oi_1 _12551_ (.A1(net64),
    .A2(_04791_),
    .Y(_00411_),
    .B1(_04242_));
 sg13g2_buf_1 _12552_ (.A(net140),
    .X(_04792_));
 sg13g2_buf_1 _12553_ (.A(net502),
    .X(_04793_));
 sg13g2_nor2_1 _12554_ (.A(_04302_),
    .B(_04306_),
    .Y(_04794_));
 sg13g2_xnor2_1 _12555_ (.Y(_04795_),
    .A(_02815_),
    .B(_04794_));
 sg13g2_nor2_1 _12556_ (.A(_04793_),
    .B(_04795_),
    .Y(_04796_));
 sg13g2_xnor2_1 _12557_ (.Y(_04797_),
    .A(_04288_),
    .B(_04796_));
 sg13g2_a21oi_1 _12558_ (.A1(net63),
    .A2(_04797_),
    .Y(_00412_),
    .B1(_04247_));
 sg13g2_xnor2_1 _12559_ (.Y(_04798_),
    .A(_02837_),
    .B(_04309_));
 sg13g2_nor2_1 _12560_ (.A(net446),
    .B(_04798_),
    .Y(_04799_));
 sg13g2_xnor2_1 _12561_ (.Y(_04800_),
    .A(_04289_),
    .B(_04799_));
 sg13g2_o21ai_1 _12562_ (.B1(_04253_),
    .Y(_00413_),
    .A1(net135),
    .A2(_04800_));
 sg13g2_xnor2_1 _12563_ (.Y(_04801_),
    .A(_02853_),
    .B(_04299_));
 sg13g2_nor2_1 _12564_ (.A(net405),
    .B(_04801_),
    .Y(_04802_));
 sg13g2_xnor2_1 _12565_ (.Y(_04803_),
    .A(_04269_),
    .B(_04802_));
 sg13g2_nor2_1 _12566_ (.A(net83),
    .B(_04256_),
    .Y(_04804_));
 sg13g2_a21oi_1 _12567_ (.A1(net63),
    .A2(_04803_),
    .Y(_00414_),
    .B1(_04804_));
 sg13g2_xnor2_1 _12568_ (.Y(_04805_),
    .A(net535),
    .B(_04314_));
 sg13g2_nand3_1 _12569_ (.B(net147),
    .C(_04805_),
    .A(net565),
    .Y(_04806_));
 sg13g2_or4_1 _12570_ (.A(net565),
    .B(net233),
    .C(net448),
    .D(_04805_),
    .X(_04807_));
 sg13g2_nand3_1 _12571_ (.B(net161),
    .C(net448),
    .A(_04266_),
    .Y(_04808_));
 sg13g2_nand4_1 _12572_ (.B(_04806_),
    .C(_04807_),
    .A(_04262_),
    .Y(_00415_),
    .D(_04808_));
 sg13g2_inv_1 _12573_ (.Y(_04809_),
    .A(\clock_inst.sec_a[0] ));
 sg13g2_buf_1 _12574_ (.A(\clock_inst.second[4] ),
    .X(_04810_));
 sg13g2_inv_1 _12575_ (.Y(_04811_),
    .A(net561));
 sg13g2_buf_2 _12576_ (.A(\clock_inst.second[5] ),
    .X(_04812_));
 sg13g2_inv_2 _12577_ (.Y(_04813_),
    .A(_04812_));
 sg13g2_nor2_1 _12578_ (.A(_04811_),
    .B(_04813_),
    .Y(_04814_));
 sg13g2_buf_2 _12579_ (.A(_04814_),
    .X(_04815_));
 sg13g2_buf_1 _12580_ (.A(\clock_inst.second[3] ),
    .X(_04816_));
 sg13g2_inv_1 _12581_ (.Y(_04817_),
    .A(net560));
 sg13g2_buf_1 _12582_ (.A(_04817_),
    .X(_04818_));
 sg13g2_buf_1 _12583_ (.A(\clock_inst.second[2] ),
    .X(_04819_));
 sg13g2_inv_1 _12584_ (.Y(_04820_),
    .A(_04819_));
 sg13g2_nor2_1 _12585_ (.A(net476),
    .B(_04820_),
    .Y(_04821_));
 sg13g2_buf_2 _12586_ (.A(_04821_),
    .X(_04822_));
 sg13g2_a21oi_1 _12587_ (.A1(_04815_),
    .A2(_04822_),
    .Y(_04823_),
    .B1(_00688_));
 sg13g2_buf_1 _12588_ (.A(_04823_),
    .X(_04824_));
 sg13g2_buf_1 _12589_ (.A(_04824_),
    .X(_04825_));
 sg13g2_buf_1 _12590_ (.A(\clock_inst.second[1] ),
    .X(_04826_));
 sg13g2_buf_1 _12591_ (.A(_04826_),
    .X(_04827_));
 sg13g2_buf_1 _12592_ (.A(net530),
    .X(_04828_));
 sg13g2_buf_1 _12593_ (.A(net475),
    .X(_04829_));
 sg13g2_buf_1 _12594_ (.A(_04829_),
    .X(_04830_));
 sg13g2_buf_1 _12595_ (.A(net294),
    .X(_04831_));
 sg13g2_buf_2 _12596_ (.A(\clock_inst.second[0] ),
    .X(_04832_));
 sg13g2_buf_1 _12597_ (.A(_04832_),
    .X(_04833_));
 sg13g2_buf_1 _12598_ (.A(_04811_),
    .X(_04834_));
 sg13g2_nor2_1 _12599_ (.A(net529),
    .B(_04834_),
    .Y(_04835_));
 sg13g2_buf_2 _12600_ (.A(_04835_),
    .X(_04836_));
 sg13g2_inv_2 _12601_ (.Y(_04837_),
    .A(_04832_));
 sg13g2_nor2_1 _12602_ (.A(_04837_),
    .B(net561),
    .Y(_04838_));
 sg13g2_buf_1 _12603_ (.A(_04838_),
    .X(_04839_));
 sg13g2_nor2_1 _12604_ (.A(_04836_),
    .B(net403),
    .Y(_04840_));
 sg13g2_buf_1 _12605_ (.A(_04820_),
    .X(_04841_));
 sg13g2_buf_1 _12606_ (.A(_04813_),
    .X(_04842_));
 sg13g2_nand2_1 _12607_ (.Y(_04843_),
    .A(net473),
    .B(net472));
 sg13g2_buf_1 _12608_ (.A(_04843_),
    .X(_04844_));
 sg13g2_nor3_1 _12609_ (.A(net192),
    .B(_04840_),
    .C(net293),
    .Y(_04845_));
 sg13g2_buf_1 _12610_ (.A(net560),
    .X(_04846_));
 sg13g2_buf_1 _12611_ (.A(net528),
    .X(_04847_));
 sg13g2_buf_1 _12612_ (.A(net471),
    .X(_04848_));
 sg13g2_buf_1 _12613_ (.A(net402),
    .X(_04849_));
 sg13g2_buf_1 _12614_ (.A(net561),
    .X(_04850_));
 sg13g2_nor2_1 _12615_ (.A(net529),
    .B(net527),
    .Y(_04851_));
 sg13g2_buf_2 _12616_ (.A(_04851_),
    .X(_04852_));
 sg13g2_buf_1 _12617_ (.A(net530),
    .X(_04853_));
 sg13g2_buf_1 _12618_ (.A(_04819_),
    .X(_04854_));
 sg13g2_buf_1 _12619_ (.A(_04812_),
    .X(_04855_));
 sg13g2_nor2_1 _12620_ (.A(net526),
    .B(net525),
    .Y(_04856_));
 sg13g2_buf_1 _12621_ (.A(_04856_),
    .X(_04857_));
 sg13g2_buf_1 _12622_ (.A(net473),
    .X(_04858_));
 sg13g2_nand2_2 _12623_ (.Y(_04859_),
    .A(net475),
    .B(net400));
 sg13g2_o21ai_1 _12624_ (.B1(_04859_),
    .Y(_04860_),
    .A1(net470),
    .A2(net401));
 sg13g2_buf_2 _12625_ (.A(net526),
    .X(_04861_));
 sg13g2_buf_1 _12626_ (.A(net469),
    .X(_04862_));
 sg13g2_nand2_2 _12627_ (.Y(_04863_),
    .A(net399),
    .B(_04815_));
 sg13g2_nor2_1 _12628_ (.A(_04841_),
    .B(net472),
    .Y(_04864_));
 sg13g2_nor2_1 _12629_ (.A(net526),
    .B(net474),
    .Y(_04865_));
 sg13g2_buf_1 _12630_ (.A(_04865_),
    .X(_04866_));
 sg13g2_buf_1 _12631_ (.A(net529),
    .X(_04867_));
 sg13g2_buf_1 _12632_ (.A(net468),
    .X(_04868_));
 sg13g2_o21ai_1 _12633_ (.B1(net398),
    .Y(_04869_),
    .A1(_04864_),
    .A2(net291));
 sg13g2_nand2_1 _12634_ (.Y(_04870_),
    .A(_04863_),
    .B(_04869_));
 sg13g2_buf_1 _12635_ (.A(net470),
    .X(_04871_));
 sg13g2_buf_1 _12636_ (.A(net525),
    .X(_04872_));
 sg13g2_buf_1 _12637_ (.A(net467),
    .X(_04873_));
 sg13g2_buf_1 _12638_ (.A(net530),
    .X(_04874_));
 sg13g2_buf_1 _12639_ (.A(_04837_),
    .X(_04875_));
 sg13g2_nor2_2 _12640_ (.A(net530),
    .B(net465),
    .Y(_04876_));
 sg13g2_nor2_1 _12641_ (.A(_04820_),
    .B(_04811_),
    .Y(_04877_));
 sg13g2_buf_1 _12642_ (.A(_04877_),
    .X(_04878_));
 sg13g2_a22oi_1 _12643_ (.Y(_04879_),
    .B1(_04876_),
    .B2(net395),
    .A2(_04852_),
    .A1(net466));
 sg13g2_nor2_1 _12644_ (.A(net465),
    .B(net526),
    .Y(_04880_));
 sg13g2_buf_2 _12645_ (.A(_04880_),
    .X(_04881_));
 sg13g2_nand2_1 _12646_ (.Y(_04882_),
    .A(_04815_),
    .B(_04881_));
 sg13g2_o21ai_1 _12647_ (.B1(_04882_),
    .Y(_04883_),
    .A1(net396),
    .A2(_04879_));
 sg13g2_a221oi_1 _12648_ (.B2(net397),
    .C1(_04883_),
    .B1(_04870_),
    .A1(_04852_),
    .Y(_04884_),
    .A2(_04860_));
 sg13g2_inv_1 _12649_ (.Y(_04885_),
    .A(_04826_));
 sg13g2_buf_1 _12650_ (.A(_04885_),
    .X(_04886_));
 sg13g2_buf_1 _12651_ (.A(net464),
    .X(_04887_));
 sg13g2_buf_1 _12652_ (.A(net394),
    .X(_04888_));
 sg13g2_nand2_1 _12653_ (.Y(_04889_),
    .A(net526),
    .B(net474));
 sg13g2_buf_1 _12654_ (.A(_04889_),
    .X(_04890_));
 sg13g2_nor2_1 _12655_ (.A(_04832_),
    .B(_04855_),
    .Y(_04891_));
 sg13g2_buf_2 _12656_ (.A(_04891_),
    .X(_04892_));
 sg13g2_nand2_1 _12657_ (.Y(_04893_),
    .A(_04811_),
    .B(_04812_));
 sg13g2_buf_1 _12658_ (.A(_04893_),
    .X(_04894_));
 sg13g2_nand2_1 _12659_ (.Y(_04895_),
    .A(net529),
    .B(_04813_));
 sg13g2_buf_2 _12660_ (.A(_04895_),
    .X(_04896_));
 sg13g2_o21ai_1 _12661_ (.B1(_04896_),
    .Y(_04897_),
    .A1(net468),
    .A2(net393));
 sg13g2_buf_1 _12662_ (.A(net469),
    .X(_04898_));
 sg13g2_a22oi_1 _12663_ (.Y(_04899_),
    .B1(_04897_),
    .B2(net392),
    .A2(_04892_),
    .A1(_04890_));
 sg13g2_nor2_1 _12664_ (.A(net290),
    .B(_04899_),
    .Y(_04900_));
 sg13g2_nand2_1 _12665_ (.Y(_04901_),
    .A(net464),
    .B(_04837_));
 sg13g2_buf_2 _12666_ (.A(_04901_),
    .X(_04902_));
 sg13g2_nand2_1 _12667_ (.Y(_04903_),
    .A(net473),
    .B(net525));
 sg13g2_buf_1 _12668_ (.A(_04903_),
    .X(_04904_));
 sg13g2_nor2_1 _12669_ (.A(net526),
    .B(net561),
    .Y(_04905_));
 sg13g2_buf_1 _12670_ (.A(_04905_),
    .X(_04906_));
 sg13g2_buf_1 _12671_ (.A(net527),
    .X(_04907_));
 sg13g2_a21oi_1 _12672_ (.A1(net463),
    .A2(_04843_),
    .Y(_04908_),
    .B1(net475));
 sg13g2_buf_1 _12673_ (.A(_04867_),
    .X(_04909_));
 sg13g2_o21ai_1 _12674_ (.B1(net390),
    .Y(_04910_),
    .A1(net391),
    .A2(_04908_));
 sg13g2_o21ai_1 _12675_ (.B1(_04910_),
    .Y(_04911_),
    .A1(_04902_),
    .A2(net289));
 sg13g2_buf_1 _12676_ (.A(net560),
    .X(_04912_));
 sg13g2_buf_1 _12677_ (.A(net524),
    .X(_04913_));
 sg13g2_buf_1 _12678_ (.A(net462),
    .X(_04914_));
 sg13g2_buf_1 _12679_ (.A(net389),
    .X(_04915_));
 sg13g2_o21ai_1 _12680_ (.B1(net288),
    .Y(_04916_),
    .A1(_04900_),
    .A2(_04911_));
 sg13g2_o21ai_1 _12681_ (.B1(_04916_),
    .Y(_04917_),
    .A1(net292),
    .A2(_04884_));
 sg13g2_nand2_1 _12682_ (.Y(_04918_),
    .A(net561),
    .B(_04812_));
 sg13g2_buf_1 _12683_ (.A(_04918_),
    .X(_04919_));
 sg13g2_nand2_1 _12684_ (.Y(_04920_),
    .A(net560),
    .B(_04819_));
 sg13g2_buf_1 _12685_ (.A(_04920_),
    .X(_04921_));
 sg13g2_o21ai_1 _12686_ (.B1(net583),
    .Y(_04922_),
    .A1(net461),
    .A2(net460));
 sg13g2_buf_1 _12687_ (.A(_04922_),
    .X(_04923_));
 sg13g2_nand2_1 _12688_ (.Y(_04924_),
    .A(net476),
    .B(_04820_));
 sg13g2_buf_2 _12689_ (.A(_04924_),
    .X(_04925_));
 sg13g2_nor2_1 _12690_ (.A(_04826_),
    .B(_04832_),
    .Y(_04926_));
 sg13g2_buf_2 _12691_ (.A(_04926_),
    .X(_04927_));
 sg13g2_nor2_1 _12692_ (.A(net561),
    .B(_04812_),
    .Y(_04928_));
 sg13g2_buf_1 _12693_ (.A(_04928_),
    .X(_04929_));
 sg13g2_nand2_1 _12694_ (.Y(_04930_),
    .A(_04927_),
    .B(_04929_));
 sg13g2_nor2_1 _12695_ (.A(_04925_),
    .B(_04930_),
    .Y(_04931_));
 sg13g2_nor2_1 _12696_ (.A(_04923_),
    .B(_04931_),
    .Y(_04932_));
 sg13g2_buf_1 _12697_ (.A(_04932_),
    .X(_04933_));
 sg13g2_o21ai_1 _12698_ (.B1(_04933_),
    .Y(_04934_),
    .A1(_04845_),
    .A2(_04917_));
 sg13g2_o21ai_1 _12699_ (.B1(_04934_),
    .Y(_00422_),
    .A1(_04809_),
    .A2(net62));
 sg13g2_buf_2 _12700_ (.A(\clock_inst.sec_a[10] ),
    .X(_04935_));
 sg13g2_buf_1 _12701_ (.A(_04923_),
    .X(_04936_));
 sg13g2_buf_1 _12702_ (.A(net191),
    .X(_04937_));
 sg13g2_buf_1 _12703_ (.A(net191),
    .X(_04938_));
 sg13g2_nor2_1 _12704_ (.A(_04811_),
    .B(_04812_),
    .Y(_04939_));
 sg13g2_buf_1 _12705_ (.A(_04939_),
    .X(_04940_));
 sg13g2_buf_1 _12706_ (.A(net388),
    .X(_04941_));
 sg13g2_buf_1 _12707_ (.A(net399),
    .X(_04942_));
 sg13g2_buf_1 _12708_ (.A(net286),
    .X(_04943_));
 sg13g2_buf_1 _12709_ (.A(net476),
    .X(_04944_));
 sg13g2_buf_1 _12710_ (.A(net387),
    .X(_04945_));
 sg13g2_nor2_2 _12711_ (.A(net394),
    .B(net285),
    .Y(_04946_));
 sg13g2_buf_1 _12712_ (.A(net393),
    .X(_04947_));
 sg13g2_a21oi_1 _12713_ (.A1(net190),
    .A2(_04946_),
    .Y(_04948_),
    .B1(net284));
 sg13g2_nor3_1 _12714_ (.A(net122),
    .B(_04941_),
    .C(_04948_),
    .Y(_04949_));
 sg13g2_a21o_1 _12715_ (.A2(net123),
    .A1(_04935_),
    .B1(_04949_),
    .X(_00423_));
 sg13g2_buf_1 _12716_ (.A(net191),
    .X(_04950_));
 sg13g2_buf_1 _12717_ (.A(net470),
    .X(_04951_));
 sg13g2_buf_1 _12718_ (.A(net386),
    .X(_04952_));
 sg13g2_buf_1 _12719_ (.A(net283),
    .X(_04953_));
 sg13g2_buf_1 _12720_ (.A(net463),
    .X(_04954_));
 sg13g2_buf_1 _12721_ (.A(net385),
    .X(_04955_));
 sg13g2_buf_1 _12722_ (.A(net465),
    .X(_04956_));
 sg13g2_buf_1 _12723_ (.A(net384),
    .X(_04957_));
 sg13g2_nand2_1 _12724_ (.Y(_04958_),
    .A(net387),
    .B(_04854_));
 sg13g2_buf_2 _12725_ (.A(_04958_),
    .X(_04959_));
 sg13g2_buf_1 _12726_ (.A(net472),
    .X(_04960_));
 sg13g2_buf_1 _12727_ (.A(_04960_),
    .X(_04961_));
 sg13g2_o21ai_1 _12728_ (.B1(net280),
    .Y(_04962_),
    .A1(_04957_),
    .A2(_04959_));
 sg13g2_nand2_1 _12729_ (.Y(_04963_),
    .A(net528),
    .B(net391));
 sg13g2_buf_2 _12730_ (.A(_04963_),
    .X(_04964_));
 sg13g2_nand2_1 _12731_ (.Y(_04965_),
    .A(net280),
    .B(_04964_));
 sg13g2_buf_1 _12732_ (.A(net398),
    .X(_04966_));
 sg13g2_buf_1 _12733_ (.A(_04966_),
    .X(_04967_));
 sg13g2_nand2_1 _12734_ (.Y(_04968_),
    .A(net474),
    .B(net472));
 sg13g2_buf_2 _12735_ (.A(_04968_),
    .X(_04969_));
 sg13g2_buf_1 _12736_ (.A(_04969_),
    .X(_04970_));
 sg13g2_nand2_1 _12737_ (.Y(_04971_),
    .A(net528),
    .B(_04865_));
 sg13g2_buf_1 _12738_ (.A(_04833_),
    .X(_04972_));
 sg13g2_buf_1 _12739_ (.A(net458),
    .X(_04973_));
 sg13g2_buf_1 _12740_ (.A(net382),
    .X(_04974_));
 sg13g2_a21oi_1 _12741_ (.A1(_04970_),
    .A2(_04971_),
    .Y(_04975_),
    .B1(net278));
 sg13g2_a221oi_1 _12742_ (.B2(net188),
    .C1(_04975_),
    .B1(_04965_),
    .A1(net282),
    .Y(_04976_),
    .A2(_04962_));
 sg13g2_nand2_1 _12743_ (.Y(_04977_),
    .A(net466),
    .B(net383));
 sg13g2_inv_1 _12744_ (.Y(_04978_),
    .A(_04977_));
 sg13g2_buf_1 _12745_ (.A(net392),
    .X(_04979_));
 sg13g2_nor2_1 _12746_ (.A(net277),
    .B(_04852_),
    .Y(_04980_));
 sg13g2_nand2_1 _12747_ (.Y(_04981_),
    .A(net473),
    .B(net474));
 sg13g2_buf_1 _12748_ (.A(_04981_),
    .X(_04982_));
 sg13g2_nand2_2 _12749_ (.Y(_04983_),
    .A(_04826_),
    .B(_04837_));
 sg13g2_nand2_1 _12750_ (.Y(_04984_),
    .A(net528),
    .B(net395));
 sg13g2_buf_1 _12751_ (.A(_04984_),
    .X(_04985_));
 sg13g2_o21ai_1 _12752_ (.B1(_04985_),
    .Y(_04986_),
    .A1(_04982_),
    .A2(_04983_));
 sg13g2_buf_1 _12753_ (.A(net396),
    .X(_04987_));
 sg13g2_nor2_1 _12754_ (.A(net473),
    .B(net527),
    .Y(_04988_));
 sg13g2_buf_1 _12755_ (.A(_04988_),
    .X(_04989_));
 sg13g2_nand2_1 _12756_ (.Y(_04990_),
    .A(net384),
    .B(_04989_));
 sg13g2_nand2_2 _12757_ (.Y(_04991_),
    .A(_04832_),
    .B(net561));
 sg13g2_and2_1 _12758_ (.A(net469),
    .B(_04991_),
    .X(_04992_));
 sg13g2_buf_1 _12759_ (.A(_04992_),
    .X(_04993_));
 sg13g2_nand2_1 _12760_ (.Y(_04994_),
    .A(net473),
    .B(net527));
 sg13g2_a21oi_1 _12761_ (.A1(net467),
    .A2(_04994_),
    .Y(_04995_),
    .B1(net384));
 sg13g2_buf_1 _12762_ (.A(net466),
    .X(_04996_));
 sg13g2_o21ai_1 _12763_ (.B1(net381),
    .Y(_04997_),
    .A1(_04993_),
    .A2(_04995_));
 sg13g2_a21oi_1 _12764_ (.A1(_04990_),
    .A2(_04997_),
    .Y(_04998_),
    .B1(net288));
 sg13g2_a221oi_1 _12765_ (.B2(_04987_),
    .C1(_04998_),
    .B1(_04986_),
    .A1(_04978_),
    .Y(_04999_),
    .A2(_04980_));
 sg13g2_o21ai_1 _12766_ (.B1(_04999_),
    .Y(_05000_),
    .A1(net189),
    .A2(_04976_));
 sg13g2_buf_1 _12767_ (.A(\clock_inst.sec_a[18] ),
    .X(_05001_));
 sg13g2_buf_1 _12768_ (.A(net191),
    .X(_05002_));
 sg13g2_nand2_1 _12769_ (.Y(_05003_),
    .A(net559),
    .B(net120));
 sg13g2_o21ai_1 _12770_ (.B1(_05003_),
    .Y(_00424_),
    .A1(net121),
    .A2(_05000_));
 sg13g2_nand2b_1 _12771_ (.Y(_05004_),
    .B(_04824_),
    .A_N(_04931_));
 sg13g2_buf_1 _12772_ (.A(_05004_),
    .X(_05005_));
 sg13g2_buf_1 _12773_ (.A(_05005_),
    .X(_05006_));
 sg13g2_nor2_1 _12774_ (.A(_04827_),
    .B(net524),
    .Y(_05007_));
 sg13g2_buf_1 _12775_ (.A(_05007_),
    .X(_05008_));
 sg13g2_nand2_2 _12776_ (.Y(_05009_),
    .A(net399),
    .B(net459));
 sg13g2_inv_1 _12777_ (.Y(_05010_),
    .A(_05009_));
 sg13g2_buf_1 _12778_ (.A(net290),
    .X(_05011_));
 sg13g2_nand2_1 _12779_ (.Y(_05012_),
    .A(_04810_),
    .B(_04813_));
 sg13g2_buf_2 _12780_ (.A(_05012_),
    .X(_05013_));
 sg13g2_buf_1 _12781_ (.A(_05013_),
    .X(_05014_));
 sg13g2_nor2_1 _12782_ (.A(net561),
    .B(net472),
    .Y(_05015_));
 sg13g2_buf_1 _12783_ (.A(_05015_),
    .X(_05016_));
 sg13g2_nand2_1 _12784_ (.Y(_05017_),
    .A(net392),
    .B(net273));
 sg13g2_o21ai_1 _12785_ (.B1(_05017_),
    .Y(_05018_),
    .A1(net186),
    .A2(net274));
 sg13g2_buf_1 _12786_ (.A(net462),
    .X(_05019_));
 sg13g2_buf_1 _12787_ (.A(net379),
    .X(_05020_));
 sg13g2_buf_1 _12788_ (.A(net272),
    .X(_05021_));
 sg13g2_buf_1 _12789_ (.A(net390),
    .X(_05022_));
 sg13g2_nor2_2 _12790_ (.A(net476),
    .B(net474),
    .Y(_05023_));
 sg13g2_nand2_1 _12791_ (.Y(_05024_),
    .A(net529),
    .B(net387));
 sg13g2_buf_2 _12792_ (.A(_05024_),
    .X(_05025_));
 sg13g2_nand2_1 _12793_ (.Y(_05026_),
    .A(net524),
    .B(net527));
 sg13g2_buf_2 _12794_ (.A(_05026_),
    .X(_05027_));
 sg13g2_o21ai_1 _12795_ (.B1(_05027_),
    .Y(_05028_),
    .A1(_04969_),
    .A2(_05025_));
 sg13g2_buf_1 _12796_ (.A(net475),
    .X(_05029_));
 sg13g2_buf_1 _12797_ (.A(net378),
    .X(_05030_));
 sg13g2_a22oi_1 _12798_ (.Y(_05031_),
    .B1(_05028_),
    .B2(net270),
    .A2(_05023_),
    .A1(net271));
 sg13g2_buf_1 _12799_ (.A(_04873_),
    .X(_05032_));
 sg13g2_nor2_2 _12800_ (.A(_04875_),
    .B(_04846_),
    .Y(_05033_));
 sg13g2_nor2_2 _12801_ (.A(net468),
    .B(net387),
    .Y(_05034_));
 sg13g2_o21ai_1 _12802_ (.B1(net381),
    .Y(_05035_),
    .A1(_05033_),
    .A2(_05034_));
 sg13g2_buf_1 _12803_ (.A(_04886_),
    .X(_05036_));
 sg13g2_nand2_1 _12804_ (.Y(_05037_),
    .A(net465),
    .B(net524));
 sg13g2_nand2_1 _12805_ (.Y(_05038_),
    .A(net476),
    .B(net474));
 sg13g2_buf_2 _12806_ (.A(_05038_),
    .X(_05039_));
 sg13g2_nand3_1 _12807_ (.B(_05037_),
    .C(_05039_),
    .A(_05036_),
    .Y(_05040_));
 sg13g2_nand3_1 _12808_ (.B(_05035_),
    .C(_05040_),
    .A(net269),
    .Y(_05041_));
 sg13g2_buf_1 _12809_ (.A(net392),
    .X(_05042_));
 sg13g2_buf_1 _12810_ (.A(net268),
    .X(_05043_));
 sg13g2_a21oi_1 _12811_ (.A1(_05031_),
    .A2(_05041_),
    .Y(_05044_),
    .B1(net184));
 sg13g2_a221oi_1 _12812_ (.B2(net185),
    .C1(_05044_),
    .B1(_05018_),
    .A1(net380),
    .Y(_05045_),
    .A2(_05010_));
 sg13g2_buf_1 _12813_ (.A(\clock_inst.sec_a[19] ),
    .X(_05046_));
 sg13g2_nand2_1 _12814_ (.Y(_05047_),
    .A(_05046_),
    .B(_05002_));
 sg13g2_o21ai_1 _12815_ (.B1(_05047_),
    .Y(_00425_),
    .A1(_05006_),
    .A2(_05045_));
 sg13g2_inv_1 _12816_ (.Y(_05048_),
    .A(\clock_inst.sec_a[1] ));
 sg13g2_buf_1 _12817_ (.A(net122),
    .X(_05049_));
 sg13g2_nand2_1 _12818_ (.Y(_05050_),
    .A(net560),
    .B(_04820_));
 sg13g2_buf_2 _12819_ (.A(_05050_),
    .X(_05051_));
 sg13g2_nand2_2 _12820_ (.Y(_05052_),
    .A(net464),
    .B(_04832_));
 sg13g2_nand2_1 _12821_ (.Y(_05053_),
    .A(_05052_),
    .B(_04983_));
 sg13g2_nor3_1 _12822_ (.A(net393),
    .B(_05051_),
    .C(_05053_),
    .Y(_05054_));
 sg13g2_nor2_1 _12823_ (.A(_05005_),
    .B(_05054_),
    .Y(_05055_));
 sg13g2_nor2_1 _12824_ (.A(net464),
    .B(net468),
    .Y(_05056_));
 sg13g2_buf_1 _12825_ (.A(_05056_),
    .X(_05057_));
 sg13g2_nor2_1 _12826_ (.A(net475),
    .B(_04896_),
    .Y(_05058_));
 sg13g2_nor2_1 _12827_ (.A(net524),
    .B(_04981_),
    .Y(_05059_));
 sg13g2_o21ai_1 _12828_ (.B1(_05059_),
    .Y(_05060_),
    .A1(net267),
    .A2(_05058_));
 sg13g2_and2_1 _12829_ (.A(_05055_),
    .B(_05060_),
    .X(_05061_));
 sg13g2_buf_1 _12830_ (.A(net395),
    .X(_05062_));
 sg13g2_nor2_1 _12831_ (.A(net392),
    .B(net273),
    .Y(_05063_));
 sg13g2_nand2_2 _12832_ (.Y(_05064_),
    .A(_04862_),
    .B(net463));
 sg13g2_a21oi_1 _12833_ (.A1(_05064_),
    .A2(_04896_),
    .Y(_05065_),
    .B1(net386));
 sg13g2_a221oi_1 _12834_ (.B2(_05063_),
    .C1(_05065_),
    .B1(net267),
    .A1(net271),
    .Y(_05066_),
    .A2(net266));
 sg13g2_buf_1 _12835_ (.A(net389),
    .X(_05067_));
 sg13g2_buf_1 _12836_ (.A(net459),
    .X(_05068_));
 sg13g2_nand2_1 _12837_ (.Y(_05069_),
    .A(net530),
    .B(net468));
 sg13g2_buf_2 _12838_ (.A(_05069_),
    .X(_05070_));
 sg13g2_a21oi_1 _12839_ (.A1(net385),
    .A2(_05070_),
    .Y(_05071_),
    .B1(net286));
 sg13g2_nand2_1 _12840_ (.Y(_05072_),
    .A(net398),
    .B(_04864_));
 sg13g2_buf_1 _12841_ (.A(net465),
    .X(_05073_));
 sg13g2_nand2_1 _12842_ (.Y(_05074_),
    .A(net375),
    .B(net401));
 sg13g2_a21oi_1 _12843_ (.A1(_05072_),
    .A2(_05074_),
    .Y(_05075_),
    .B1(net386));
 sg13g2_nor4_1 _12844_ (.A(net265),
    .B(net376),
    .C(_05071_),
    .D(_05075_),
    .Y(_05076_));
 sg13g2_a21oi_1 _12845_ (.A1(net292),
    .A2(_05066_),
    .Y(_05077_),
    .B1(_05076_));
 sg13g2_nor2_1 _12846_ (.A(net530),
    .B(net469),
    .Y(_05078_));
 sg13g2_buf_2 _12847_ (.A(_05078_),
    .X(_05079_));
 sg13g2_buf_1 _12848_ (.A(net273),
    .X(_05080_));
 sg13g2_nand2_2 _12849_ (.Y(_05081_),
    .A(net465),
    .B(_04861_));
 sg13g2_nand2_1 _12850_ (.Y(_05082_),
    .A(_04854_),
    .B(net472));
 sg13g2_buf_2 _12851_ (.A(_05082_),
    .X(_05083_));
 sg13g2_nand2_1 _12852_ (.Y(_05084_),
    .A(_05083_),
    .B(net289));
 sg13g2_nand2_1 _12853_ (.Y(_05085_),
    .A(net271),
    .B(_05084_));
 sg13g2_o21ai_1 _12854_ (.B1(_05085_),
    .Y(_05086_),
    .A1(net461),
    .A2(_05081_));
 sg13g2_buf_1 _12855_ (.A(_05030_),
    .X(_05087_));
 sg13g2_a22oi_1 _12856_ (.Y(_05088_),
    .B1(_05086_),
    .B2(net182),
    .A2(net183),
    .A1(_05079_));
 sg13g2_nand2b_1 _12857_ (.Y(_05089_),
    .B(_05088_),
    .A_N(_05077_));
 sg13g2_a22oi_1 _12858_ (.Y(_00426_),
    .B1(_05061_),
    .B2(_05089_),
    .A2(net60),
    .A1(_05048_));
 sg13g2_buf_2 _12859_ (.A(\clock_inst.sec_a[20] ),
    .X(_05090_));
 sg13g2_buf_1 _12860_ (.A(_04936_),
    .X(_05091_));
 sg13g2_buf_1 _12861_ (.A(net61),
    .X(_05092_));
 sg13g2_buf_1 _12862_ (.A(net265),
    .X(_05093_));
 sg13g2_buf_1 _12863_ (.A(_04815_),
    .X(_05094_));
 sg13g2_a21oi_1 _12864_ (.A1(net264),
    .A2(net267),
    .Y(_05095_),
    .B1(net459));
 sg13g2_nand2_1 _12865_ (.Y(_05096_),
    .A(net377),
    .B(net459));
 sg13g2_o21ai_1 _12866_ (.B1(_05096_),
    .Y(_05097_),
    .A1(net190),
    .A2(_05095_));
 sg13g2_buf_1 _12867_ (.A(net467),
    .X(_05098_));
 sg13g2_nor2_1 _12868_ (.A(_04827_),
    .B(net474),
    .Y(_05099_));
 sg13g2_buf_2 _12869_ (.A(_05099_),
    .X(_05100_));
 sg13g2_o21ai_1 _12870_ (.B1(net277),
    .Y(_05101_),
    .A1(net374),
    .A2(_05100_));
 sg13g2_buf_1 _12871_ (.A(net394),
    .X(_05102_));
 sg13g2_nand2_1 _12872_ (.Y(_05103_),
    .A(net468),
    .B(_04939_));
 sg13g2_o21ai_1 _12873_ (.B1(_05103_),
    .Y(_05104_),
    .A1(net458),
    .A2(net393));
 sg13g2_nand2_1 _12874_ (.Y(_05105_),
    .A(_04841_),
    .B(net388));
 sg13g2_buf_2 _12875_ (.A(_05105_),
    .X(_05106_));
 sg13g2_nand2_1 _12876_ (.Y(_05107_),
    .A(net458),
    .B(_05015_));
 sg13g2_a21oi_1 _12877_ (.A1(_05106_),
    .A2(_05107_),
    .Y(_05108_),
    .B1(net290));
 sg13g2_a21oi_1 _12878_ (.A1(net263),
    .A2(_05104_),
    .Y(_05109_),
    .B1(_05108_));
 sg13g2_nand3_1 _12879_ (.B(_05101_),
    .C(_05109_),
    .A(net272),
    .Y(_05110_));
 sg13g2_o21ai_1 _12880_ (.B1(_05110_),
    .Y(_05111_),
    .A1(net181),
    .A2(_05097_));
 sg13g2_a22oi_1 _12881_ (.Y(_05112_),
    .B1(net27),
    .B2(_05111_),
    .A2(net119),
    .A1(_05090_));
 sg13g2_inv_1 _12882_ (.Y(_00427_),
    .A(_05112_));
 sg13g2_buf_1 _12883_ (.A(\clock_inst.sec_a[2] ),
    .X(_05113_));
 sg13g2_inv_1 _12884_ (.Y(_05114_),
    .A(_05113_));
 sg13g2_nor2_1 _12885_ (.A(net289),
    .B(_05039_),
    .Y(_05115_));
 sg13g2_nand2_1 _12886_ (.Y(_05116_),
    .A(_04945_),
    .B(net395));
 sg13g2_nand2_1 _12887_ (.Y(_05117_),
    .A(_05096_),
    .B(_05116_));
 sg13g2_buf_1 _12888_ (.A(net278),
    .X(_05118_));
 sg13g2_nand3_1 _12889_ (.B(_04927_),
    .C(net388),
    .A(_04822_),
    .Y(_05119_));
 sg13g2_nand2_1 _12890_ (.Y(_05120_),
    .A(_04933_),
    .B(_05119_));
 sg13g2_a221oi_1 _12891_ (.B2(net180),
    .C1(_05120_),
    .B1(_05117_),
    .A1(_05052_),
    .Y(_05121_),
    .A2(_05115_));
 sg13g2_nor2_1 _12892_ (.A(net476),
    .B(_04812_),
    .Y(_05122_));
 sg13g2_buf_1 _12893_ (.A(_05122_),
    .X(_05123_));
 sg13g2_nand2_1 _12894_ (.Y(_05124_),
    .A(_04868_),
    .B(net262));
 sg13g2_nand2b_1 _12895_ (.Y(_05125_),
    .B(_05124_),
    .A_N(_04836_));
 sg13g2_nor2_1 _12896_ (.A(net285),
    .B(_04894_),
    .Y(_05126_));
 sg13g2_buf_1 _12897_ (.A(_04927_),
    .X(_05127_));
 sg13g2_nor2_2 _12898_ (.A(net462),
    .B(_05013_),
    .Y(_05128_));
 sg13g2_a221oi_1 _12899_ (.B2(_05127_),
    .C1(_05128_),
    .B1(_05126_),
    .A1(net283),
    .Y(_05129_),
    .A2(_05125_));
 sg13g2_nand2_1 _12900_ (.Y(_05130_),
    .A(net476),
    .B(net525));
 sg13g2_buf_1 _12901_ (.A(_05130_),
    .X(_05131_));
 sg13g2_nor2_1 _12902_ (.A(_04972_),
    .B(net261),
    .Y(_05132_));
 sg13g2_a21oi_1 _12903_ (.A1(net292),
    .A2(_05068_),
    .Y(_05133_),
    .B1(_05132_));
 sg13g2_buf_1 _12904_ (.A(_04943_),
    .X(_05134_));
 sg13g2_mux2_1 _12905_ (.A0(_05129_),
    .A1(_05133_),
    .S(_05134_),
    .X(_05135_));
 sg13g2_a22oi_1 _12906_ (.Y(_00428_),
    .B1(_05121_),
    .B2(_05135_),
    .A2(net60),
    .A1(_05114_));
 sg13g2_buf_1 _12907_ (.A(net269),
    .X(_05136_));
 sg13g2_nor2_1 _12908_ (.A(_04977_),
    .B(_04985_),
    .Y(_05137_));
 sg13g2_a21oi_1 _12909_ (.A1(net179),
    .A2(_04985_),
    .Y(_05138_),
    .B1(_05137_));
 sg13g2_buf_1 _12910_ (.A(\clock_inst.sec_a[21] ),
    .X(_05139_));
 sg13g2_buf_1 _12911_ (.A(_05139_),
    .X(_05140_));
 sg13g2_buf_1 _12912_ (.A(net523),
    .X(_05141_));
 sg13g2_buf_1 _12913_ (.A(_05141_),
    .X(_05142_));
 sg13g2_nand2_1 _12914_ (.Y(_05143_),
    .A(net372),
    .B(net120));
 sg13g2_o21ai_1 _12915_ (.B1(_05143_),
    .Y(_00429_),
    .A1(net22),
    .A2(_05138_));
 sg13g2_buf_2 _12916_ (.A(net463),
    .X(_05144_));
 sg13g2_buf_1 _12917_ (.A(net371),
    .X(_05145_));
 sg13g2_buf_1 _12918_ (.A(net286),
    .X(_05146_));
 sg13g2_nand2_2 _12919_ (.Y(_05147_),
    .A(net384),
    .B(net467));
 sg13g2_nand3_1 _12920_ (.B(_04896_),
    .C(_05147_),
    .A(net404),
    .Y(_05148_));
 sg13g2_o21ai_1 _12921_ (.B1(_05148_),
    .Y(_05149_),
    .A1(_04951_),
    .A2(_05147_));
 sg13g2_nor2_1 _12922_ (.A(_04956_),
    .B(_04945_),
    .Y(_05150_));
 sg13g2_nand2_2 _12923_ (.Y(_05151_),
    .A(net394),
    .B(net467));
 sg13g2_nand2_1 _12924_ (.Y(_05152_),
    .A(net293),
    .B(_05151_));
 sg13g2_a22oi_1 _12925_ (.Y(_05153_),
    .B1(_05150_),
    .B2(_05152_),
    .A2(_05149_),
    .A1(_05146_));
 sg13g2_buf_1 _12926_ (.A(net390),
    .X(_05154_));
 sg13g2_nor2_1 _12927_ (.A(net560),
    .B(_04813_),
    .Y(_05155_));
 sg13g2_buf_1 _12928_ (.A(_05155_),
    .X(_05156_));
 sg13g2_nor2_1 _12929_ (.A(net387),
    .B(net469),
    .Y(_05157_));
 sg13g2_buf_2 _12930_ (.A(_05157_),
    .X(_05158_));
 sg13g2_a21oi_1 _12931_ (.A1(net470),
    .A2(_05156_),
    .Y(_05159_),
    .B1(_05158_));
 sg13g2_nor2_2 _12932_ (.A(_04912_),
    .B(net469),
    .Y(_05160_));
 sg13g2_nand2_1 _12933_ (.Y(_05161_),
    .A(net398),
    .B(_05160_));
 sg13g2_o21ai_1 _12934_ (.B1(_05161_),
    .Y(_05162_),
    .A1(_05154_),
    .A2(_05159_));
 sg13g2_nor2_1 _12935_ (.A(_04820_),
    .B(_04812_),
    .Y(_05163_));
 sg13g2_buf_1 _12936_ (.A(_05163_),
    .X(_05164_));
 sg13g2_buf_1 _12937_ (.A(_05164_),
    .X(_05165_));
 sg13g2_nand2_1 _12938_ (.Y(_05166_),
    .A(net377),
    .B(net258));
 sg13g2_nor2_1 _12939_ (.A(net526),
    .B(_04813_),
    .Y(_05167_));
 sg13g2_buf_2 _12940_ (.A(_05167_),
    .X(_05168_));
 sg13g2_buf_1 _12941_ (.A(_05168_),
    .X(_05169_));
 sg13g2_nand2_1 _12942_ (.Y(_05170_),
    .A(net381),
    .B(_05169_));
 sg13g2_nor2_1 _12943_ (.A(_04818_),
    .B(_04850_),
    .Y(_05171_));
 sg13g2_buf_1 _12944_ (.A(_05171_),
    .X(_05172_));
 sg13g2_buf_1 _12945_ (.A(_05172_),
    .X(_05173_));
 sg13g2_a21oi_1 _12946_ (.A1(_05166_),
    .A2(_05170_),
    .Y(_05174_),
    .B1(_05173_));
 sg13g2_a21oi_1 _12947_ (.A1(_04955_),
    .A2(_05162_),
    .Y(_05175_),
    .B1(_05174_));
 sg13g2_o21ai_1 _12948_ (.B1(_05175_),
    .Y(_05176_),
    .A1(_05145_),
    .A2(_05153_));
 sg13g2_a22oi_1 _12949_ (.Y(_05177_),
    .B1(_05092_),
    .B2(_05176_),
    .A2(net119),
    .A1(\clock_inst.sec_a[36] ));
 sg13g2_inv_1 _12950_ (.Y(_00430_),
    .A(_05177_));
 sg13g2_inv_1 _12951_ (.Y(_05178_),
    .A(\clock_inst.sec_a[37] ));
 sg13g2_o21ai_1 _12952_ (.B1(_05161_),
    .Y(_05179_),
    .A1(net188),
    .A2(_04947_));
 sg13g2_nor2_2 _12953_ (.A(net387),
    .B(_04940_),
    .Y(_05180_));
 sg13g2_nor2_1 _12954_ (.A(net475),
    .B(net525),
    .Y(_05181_));
 sg13g2_buf_2 _12955_ (.A(_05181_),
    .X(_05182_));
 sg13g2_o21ai_1 _12956_ (.B1(_05067_),
    .Y(_05183_),
    .A1(net403),
    .A2(_05182_));
 sg13g2_o21ai_1 _12957_ (.B1(_05183_),
    .Y(_05184_),
    .A1(_04983_),
    .A2(_05180_));
 sg13g2_nor2_1 _12958_ (.A(net529),
    .B(net560),
    .Y(_05185_));
 sg13g2_buf_1 _12959_ (.A(_05185_),
    .X(_05186_));
 sg13g2_nand2_2 _12960_ (.Y(_05187_),
    .A(net463),
    .B(net369));
 sg13g2_nor2_1 _12961_ (.A(net258),
    .B(_05187_),
    .Y(_05188_));
 sg13g2_a21oi_1 _12962_ (.A1(_04881_),
    .A2(_05080_),
    .Y(_05189_),
    .B1(_05188_));
 sg13g2_nand2_1 _12963_ (.Y(_05190_),
    .A(net61),
    .B(_05189_));
 sg13g2_a221oi_1 _12964_ (.B2(net118),
    .C1(_05190_),
    .B1(_05184_),
    .A1(net189),
    .Y(_05191_),
    .A2(_05179_));
 sg13g2_nor2_2 _12965_ (.A(net468),
    .B(net469),
    .Y(_05192_));
 sg13g2_nand2_1 _12966_ (.Y(_05193_),
    .A(net269),
    .B(_05192_));
 sg13g2_a21oi_1 _12967_ (.A1(net260),
    .A2(_05193_),
    .Y(_05194_),
    .B1(net192));
 sg13g2_nor2_1 _12968_ (.A(net529),
    .B(_04981_),
    .Y(_05195_));
 sg13g2_o21ai_1 _12969_ (.B1(_05021_),
    .Y(_05196_),
    .A1(_05194_),
    .A2(_05195_));
 sg13g2_a22oi_1 _12970_ (.Y(_00431_),
    .B1(_05191_),
    .B2(_05196_),
    .A2(net60),
    .A1(_05178_));
 sg13g2_buf_2 _12971_ (.A(\clock_inst.sec_a[38] ),
    .X(_05197_));
 sg13g2_inv_1 _12972_ (.Y(_05198_),
    .A(_05197_));
 sg13g2_buf_1 _12973_ (.A(_04864_),
    .X(_05199_));
 sg13g2_nand2_1 _12974_ (.Y(_05200_),
    .A(net375),
    .B(net256));
 sg13g2_a21oi_1 _12975_ (.A1(_05106_),
    .A2(_05200_),
    .Y(_05201_),
    .B1(net181));
 sg13g2_buf_1 _12976_ (.A(net377),
    .X(_05202_));
 sg13g2_buf_1 _12977_ (.A(net255),
    .X(_05203_));
 sg13g2_nor2_1 _12978_ (.A(net524),
    .B(net527),
    .Y(_05204_));
 sg13g2_buf_1 _12979_ (.A(_05204_),
    .X(_05205_));
 sg13g2_o21ai_1 _12980_ (.B1(_04990_),
    .Y(_05206_),
    .A1(net375),
    .A2(net368));
 sg13g2_a21oi_1 _12981_ (.A1(_05039_),
    .A2(_05051_),
    .Y(_05207_),
    .B1(net398));
 sg13g2_nand2_1 _12982_ (.Y(_05208_),
    .A(net285),
    .B(_04989_));
 sg13g2_nand3b_1 _12983_ (.B(_05208_),
    .C(net374),
    .Y(_05209_),
    .A_N(_05207_));
 sg13g2_o21ai_1 _12984_ (.B1(_05209_),
    .Y(_05210_),
    .A1(net269),
    .A2(_05206_));
 sg13g2_nand2_1 _12985_ (.Y(_05211_),
    .A(net528),
    .B(_05164_));
 sg13g2_nand2_2 _12986_ (.Y(_05212_),
    .A(net400),
    .B(_04815_));
 sg13g2_a21oi_1 _12987_ (.A1(_05211_),
    .A2(_05212_),
    .Y(_05213_),
    .B1(net382));
 sg13g2_buf_1 _12988_ (.A(_04811_),
    .X(_05214_));
 sg13g2_nand2_1 _12989_ (.Y(_05215_),
    .A(_04868_),
    .B(net456));
 sg13g2_a21oi_1 _12990_ (.A1(net374),
    .A2(_04925_),
    .Y(_05216_),
    .B1(_05215_));
 sg13g2_a21oi_1 _12991_ (.A1(net293),
    .A2(_04863_),
    .Y(_05217_),
    .B1(net379));
 sg13g2_nor4_1 _12992_ (.A(net255),
    .B(_05213_),
    .C(_05216_),
    .D(_05217_),
    .Y(_05218_));
 sg13g2_a21oi_1 _12993_ (.A1(net176),
    .A2(_05210_),
    .Y(_05219_),
    .B1(_05218_));
 sg13g2_o21ai_1 _12994_ (.B1(net61),
    .Y(_05220_),
    .A1(_05201_),
    .A2(_05219_));
 sg13g2_o21ai_1 _12995_ (.B1(_05220_),
    .Y(_00432_),
    .A1(_05198_),
    .A2(net62));
 sg13g2_buf_2 _12996_ (.A(\clock_inst.sec_a[39] ),
    .X(_05221_));
 sg13g2_inv_1 _12997_ (.Y(_05222_),
    .A(_05221_));
 sg13g2_o21ai_1 _12998_ (.B1(net284),
    .Y(_05223_),
    .A1(_04859_),
    .A2(net274));
 sg13g2_nand2_1 _12999_ (.Y(_05224_),
    .A(net399),
    .B(net388));
 sg13g2_buf_1 _13000_ (.A(net285),
    .X(_05225_));
 sg13g2_o21ai_1 _13001_ (.B1(net175),
    .Y(_05226_),
    .A1(net395),
    .A2(net257));
 sg13g2_nand3_1 _13002_ (.B(_05224_),
    .C(_05226_),
    .A(_04964_),
    .Y(_05227_));
 sg13g2_nor2_1 _13003_ (.A(net469),
    .B(_04893_),
    .Y(_05228_));
 sg13g2_buf_2 _13004_ (.A(_05228_),
    .X(_05229_));
 sg13g2_a221oi_1 _13005_ (.B2(net186),
    .C1(_05229_),
    .B1(_05227_),
    .A1(net272),
    .Y(_05230_),
    .A2(_05223_));
 sg13g2_buf_1 _13006_ (.A(net175),
    .X(_05231_));
 sg13g2_nand2_1 _13007_ (.Y(_05232_),
    .A(net526),
    .B(net525));
 sg13g2_buf_1 _13008_ (.A(_05232_),
    .X(_05233_));
 sg13g2_buf_1 _13009_ (.A(_05233_),
    .X(_05234_));
 sg13g2_o21ai_1 _13010_ (.B1(net293),
    .Y(_05235_),
    .A1(net290),
    .A2(net254));
 sg13g2_buf_1 _13011_ (.A(_04890_),
    .X(_05236_));
 sg13g2_o21ai_1 _13012_ (.B1(net174),
    .Y(_05237_),
    .A1(net263),
    .A2(net291));
 sg13g2_nor2_1 _13013_ (.A(net461),
    .B(_04859_),
    .Y(_05238_));
 sg13g2_a221oi_1 _13014_ (.B2(net262),
    .C1(_05238_),
    .B1(_05237_),
    .A1(net117),
    .Y(_05239_),
    .A2(_05235_));
 sg13g2_mux2_1 _13015_ (.A0(_05230_),
    .A1(_05239_),
    .S(net180),
    .X(_05240_));
 sg13g2_buf_1 _13016_ (.A(net400),
    .X(_05241_));
 sg13g2_xnor2_1 _13017_ (.Y(_05242_),
    .A(_05241_),
    .B(_04927_));
 sg13g2_nor2_1 _13018_ (.A(net471),
    .B(_04969_),
    .Y(_05243_));
 sg13g2_a21oi_2 _13019_ (.B1(_04923_),
    .Y(_05244_),
    .A2(_05243_),
    .A1(_05242_));
 sg13g2_buf_1 _13020_ (.A(net264),
    .X(_05245_));
 sg13g2_nor2_1 _13021_ (.A(net464),
    .B(net560),
    .Y(_05246_));
 sg13g2_buf_1 _13022_ (.A(_05246_),
    .X(_05247_));
 sg13g2_nand3_1 _13023_ (.B(net173),
    .C(net252),
    .A(net184),
    .Y(_05248_));
 sg13g2_and2_1 _13024_ (.A(_05244_),
    .B(_05248_),
    .X(_05249_));
 sg13g2_a22oi_1 _13025_ (.Y(_00433_),
    .B1(_05240_),
    .B2(_05249_),
    .A2(net60),
    .A1(_05222_));
 sg13g2_buf_1 _13026_ (.A(net188),
    .X(_05250_));
 sg13g2_buf_1 _13027_ (.A(net470),
    .X(_05251_));
 sg13g2_nand2_2 _13028_ (.Y(_05252_),
    .A(_04959_),
    .B(_05051_));
 sg13g2_buf_1 _13029_ (.A(_04989_),
    .X(_05253_));
 sg13g2_o21ai_1 _13030_ (.B1(_05029_),
    .Y(_05254_),
    .A1(net291),
    .A2(net172));
 sg13g2_o21ai_1 _13031_ (.B1(_05254_),
    .Y(_05255_),
    .A1(net367),
    .A2(_05252_));
 sg13g2_buf_1 _13032_ (.A(net280),
    .X(_05256_));
 sg13g2_a221oi_1 _13033_ (.B2(net171),
    .C1(_05115_),
    .B1(_05255_),
    .A1(net186),
    .Y(_05257_),
    .A2(_05062_));
 sg13g2_nor2_1 _13034_ (.A(net262),
    .B(_05155_),
    .Y(_05258_));
 sg13g2_nand2_1 _13035_ (.Y(_05259_),
    .A(net456),
    .B(_05258_));
 sg13g2_nor2_2 _13036_ (.A(_04846_),
    .B(_04858_),
    .Y(_05260_));
 sg13g2_o21ai_1 _13037_ (.B1(_04888_),
    .Y(_05261_),
    .A1(net396),
    .A2(_05260_));
 sg13g2_buf_1 _13038_ (.A(net375),
    .X(_05262_));
 sg13g2_a21oi_1 _13039_ (.A1(_05259_),
    .A2(_05261_),
    .Y(_05263_),
    .B1(net251));
 sg13g2_a221oi_1 _13040_ (.B2(_05011_),
    .C1(_05263_),
    .B1(net391),
    .A1(net178),
    .Y(_05264_),
    .A2(net173));
 sg13g2_o21ai_1 _13041_ (.B1(_05264_),
    .Y(_05265_),
    .A1(net116),
    .A2(_05257_));
 sg13g2_nand2_1 _13042_ (.Y(_05266_),
    .A(\clock_inst.sec_a[3] ),
    .B(net120));
 sg13g2_o21ai_1 _13043_ (.B1(_05266_),
    .Y(_00434_),
    .A1(net121),
    .A2(_05265_));
 sg13g2_buf_2 _13044_ (.A(\clock_inst.sec_a[40] ),
    .X(_05267_));
 sg13g2_nor2_1 _13045_ (.A(_04833_),
    .B(net473),
    .Y(_05268_));
 sg13g2_buf_1 _13046_ (.A(_05268_),
    .X(_05269_));
 sg13g2_nand2_2 _13047_ (.Y(_05270_),
    .A(net529),
    .B(_04861_));
 sg13g2_o21ai_1 _13048_ (.B1(_05270_),
    .Y(_05271_),
    .A1(net458),
    .A2(net276));
 sg13g2_nor2_2 _13049_ (.A(net466),
    .B(net383),
    .Y(_05272_));
 sg13g2_a22oi_1 _13050_ (.Y(_05273_),
    .B1(_05271_),
    .B2(_05272_),
    .A2(net250),
    .A1(net376));
 sg13g2_nor2_1 _13051_ (.A(net400),
    .B(_04892_),
    .Y(_05274_));
 sg13g2_nor2_2 _13052_ (.A(net530),
    .B(_04944_),
    .Y(_05275_));
 sg13g2_o21ai_1 _13053_ (.B1(net458),
    .Y(_05276_),
    .A1(net252),
    .A2(_05275_));
 sg13g2_nand2_1 _13054_ (.Y(_05277_),
    .A(net460),
    .B(_05276_));
 sg13g2_a22oi_1 _13055_ (.Y(_05278_),
    .B1(_05275_),
    .B2(_05168_),
    .A2(net252),
    .A1(_05083_));
 sg13g2_nor2_1 _13056_ (.A(net390),
    .B(_05278_),
    .Y(_05279_));
 sg13g2_a221oi_1 _13057_ (.B2(net280),
    .C1(_05279_),
    .B1(_05277_),
    .A1(net380),
    .Y(_05280_),
    .A2(_05274_));
 sg13g2_o21ai_1 _13058_ (.B1(net285),
    .Y(_05281_),
    .A1(net375),
    .A2(_05164_));
 sg13g2_a221oi_1 _13059_ (.B2(net381),
    .C1(net385),
    .B1(_05281_),
    .A1(_04857_),
    .Y(_05282_),
    .A2(_05034_));
 sg13g2_a21o_1 _13060_ (.A2(_05280_),
    .A1(net282),
    .B1(_05282_),
    .X(_05283_));
 sg13g2_o21ai_1 _13061_ (.B1(_05283_),
    .Y(_05284_),
    .A1(net181),
    .A2(_05273_));
 sg13g2_a22oi_1 _13062_ (.Y(_05285_),
    .B1(net27),
    .B2(_05284_),
    .A2(_05091_),
    .A1(_05267_));
 sg13g2_inv_1 _13063_ (.Y(_00435_),
    .A(_05285_));
 sg13g2_inv_1 _13064_ (.Y(_05286_),
    .A(\clock_inst.sec_a[41] ));
 sg13g2_o21ai_1 _13065_ (.B1(net367),
    .Y(_05287_),
    .A1(net385),
    .A2(net401));
 sg13g2_a21oi_1 _13066_ (.A1(_05106_),
    .A2(_05287_),
    .Y(_05288_),
    .B1(_05025_));
 sg13g2_nor2_2 _13067_ (.A(net464),
    .B(net527),
    .Y(_05289_));
 sg13g2_o21ai_1 _13068_ (.B1(_05289_),
    .Y(_05290_),
    .A1(_04881_),
    .A2(net250));
 sg13g2_a21oi_1 _13069_ (.A1(_05224_),
    .A2(_05290_),
    .Y(_05291_),
    .B1(net117));
 sg13g2_nor2_2 _13070_ (.A(net399),
    .B(_04969_),
    .Y(_05292_));
 sg13g2_nor2_1 _13071_ (.A(net382),
    .B(net256),
    .Y(_05293_));
 sg13g2_o21ai_1 _13072_ (.B1(net402),
    .Y(_05294_),
    .A1(_05292_),
    .A2(_05293_));
 sg13g2_nor2_1 _13073_ (.A(net465),
    .B(net473),
    .Y(_05295_));
 sg13g2_o21ai_1 _13074_ (.B1(_04890_),
    .Y(_05296_),
    .A1(net390),
    .A2(net401));
 sg13g2_a22oi_1 _13075_ (.Y(_05297_),
    .B1(_05296_),
    .B2(net175),
    .A2(_05295_),
    .A1(net183));
 sg13g2_buf_2 _13076_ (.A(net367),
    .X(_05298_));
 sg13g2_a21oi_1 _13077_ (.A1(_05294_),
    .A2(_05297_),
    .Y(_05299_),
    .B1(net249));
 sg13g2_or4_1 _13078_ (.A(_04936_),
    .B(_05288_),
    .C(_05291_),
    .D(_05299_),
    .X(_05300_));
 sg13g2_o21ai_1 _13079_ (.B1(_05300_),
    .Y(_00436_),
    .A1(_05286_),
    .A2(net62));
 sg13g2_buf_1 _13080_ (.A(net253),
    .X(_05301_));
 sg13g2_nand2_1 _13081_ (.Y(_05302_),
    .A(net387),
    .B(net472));
 sg13g2_buf_1 _13082_ (.A(_05302_),
    .X(_05303_));
 sg13g2_nor2_1 _13083_ (.A(_04875_),
    .B(net525),
    .Y(_05304_));
 sg13g2_buf_2 _13084_ (.A(_05304_),
    .X(_05305_));
 sg13g2_o21ai_1 _13085_ (.B1(_05147_),
    .Y(_05306_),
    .A1(net470),
    .A2(_05305_));
 sg13g2_nand2_1 _13086_ (.Y(_05307_),
    .A(_04954_),
    .B(_05306_));
 sg13g2_o21ai_1 _13087_ (.B1(_05307_),
    .Y(_05308_),
    .A1(net283),
    .A2(net169));
 sg13g2_nand2_1 _13088_ (.Y(_05309_),
    .A(net276),
    .B(_05116_));
 sg13g2_o21ai_1 _13089_ (.B1(net471),
    .Y(_05310_),
    .A1(net459),
    .A2(_05168_));
 sg13g2_a21oi_1 _13090_ (.A1(_05116_),
    .A2(_05310_),
    .Y(_05311_),
    .B1(net251));
 sg13g2_a21o_1 _13091_ (.A2(_05309_),
    .A1(net280),
    .B1(_05311_),
    .X(_05312_));
 sg13g2_o21ai_1 _13092_ (.B1(net172),
    .Y(_05313_),
    .A1(_05127_),
    .A2(net370));
 sg13g2_o21ai_1 _13093_ (.B1(_05313_),
    .Y(_05314_),
    .A1(_05052_),
    .A2(net169));
 sg13g2_a221oi_1 _13094_ (.B2(_05087_),
    .C1(_05314_),
    .B1(_05312_),
    .A1(net170),
    .Y(_05315_),
    .A2(_05308_));
 sg13g2_buf_1 _13095_ (.A(\clock_inst.sec_a[42] ),
    .X(_05316_));
 sg13g2_nand2_1 _13096_ (.Y(_05317_),
    .A(_05316_),
    .B(net120));
 sg13g2_o21ai_1 _13097_ (.B1(_05317_),
    .Y(_00437_),
    .A1(_04950_),
    .A2(_05315_));
 sg13g2_inv_1 _13098_ (.Y(_05318_),
    .A(\clock_inst.sec_a[43] ));
 sg13g2_buf_1 _13099_ (.A(_04938_),
    .X(_05319_));
 sg13g2_buf_1 _13100_ (.A(net271),
    .X(_05320_));
 sg13g2_buf_1 _13101_ (.A(net175),
    .X(_05321_));
 sg13g2_nor2_1 _13102_ (.A(net476),
    .B(net472),
    .Y(_05322_));
 sg13g2_buf_1 _13103_ (.A(_05322_),
    .X(_05323_));
 sg13g2_a21oi_1 _13104_ (.A1(net115),
    .A2(net266),
    .Y(_05324_),
    .B1(net248));
 sg13g2_o21ai_1 _13105_ (.B1(_04964_),
    .Y(_05325_),
    .A1(net168),
    .A2(_05324_));
 sg13g2_a21oi_1 _13106_ (.A1(net176),
    .A2(_05325_),
    .Y(_05326_),
    .B1(net450));
 sg13g2_buf_1 _13107_ (.A(net115),
    .X(_05327_));
 sg13g2_nor2_1 _13108_ (.A(net464),
    .B(_04837_),
    .Y(_05328_));
 sg13g2_buf_1 _13109_ (.A(_05328_),
    .X(_05329_));
 sg13g2_buf_1 _13110_ (.A(_05329_),
    .X(_05330_));
 sg13g2_o21ai_1 _13111_ (.B1(net371),
    .Y(_05331_),
    .A1(net277),
    .A2(net167));
 sg13g2_a21oi_1 _13112_ (.A1(net58),
    .A2(_05331_),
    .Y(_05332_),
    .B1(net172));
 sg13g2_o21ai_1 _13113_ (.B1(net293),
    .Y(_05333_),
    .A1(_05236_),
    .A2(net167));
 sg13g2_nor2_2 _13114_ (.A(net400),
    .B(_05013_),
    .Y(_05334_));
 sg13g2_a21oi_1 _13115_ (.A1(_05093_),
    .A2(_05333_),
    .Y(_05335_),
    .B1(_05334_));
 sg13g2_o21ai_1 _13116_ (.B1(_05335_),
    .Y(_05336_),
    .A1(_05256_),
    .A2(_05332_));
 sg13g2_a22oi_1 _13117_ (.Y(_00438_),
    .B1(_05326_),
    .B2(_05336_),
    .A2(net59),
    .A1(_05318_));
 sg13g2_inv_1 _13118_ (.Y(_05337_),
    .A(\clock_inst.sec_a[4] ));
 sg13g2_nor2_2 _13119_ (.A(net394),
    .B(net456),
    .Y(_05338_));
 sg13g2_nand2_1 _13120_ (.Y(_05339_),
    .A(_04979_),
    .B(net261));
 sg13g2_a21oi_1 _13121_ (.A1(_04829_),
    .A2(_05131_),
    .Y(_05340_),
    .B1(net380));
 sg13g2_nand2_1 _13122_ (.Y(_05341_),
    .A(_04888_),
    .B(net370));
 sg13g2_o21ai_1 _13123_ (.B1(_05341_),
    .Y(_05342_),
    .A1(_05144_),
    .A2(_05340_));
 sg13g2_nor2_1 _13124_ (.A(_04969_),
    .B(_05051_),
    .Y(_05343_));
 sg13g2_a221oi_1 _13125_ (.B2(net184),
    .C1(_05343_),
    .B1(_05342_),
    .A1(_05338_),
    .Y(_05344_),
    .A2(_05339_));
 sg13g2_nand2b_1 _13126_ (.Y(_05345_),
    .B(net116),
    .A_N(_05344_));
 sg13g2_buf_1 _13127_ (.A(net291),
    .X(_05346_));
 sg13g2_a22oi_1 _13128_ (.Y(_05347_),
    .B1(net172),
    .B2(net373),
    .A2(_05346_),
    .A1(_04952_));
 sg13g2_inv_1 _13129_ (.Y(_05348_),
    .A(_05347_));
 sg13g2_nand2_1 _13130_ (.Y(_05349_),
    .A(_04887_),
    .B(_04858_));
 sg13g2_nand2_1 _13131_ (.Y(_05350_),
    .A(net285),
    .B(_05164_));
 sg13g2_o21ai_1 _13132_ (.B1(_05350_),
    .Y(_05351_),
    .A1(_05349_),
    .A2(net248));
 sg13g2_a22oi_1 _13133_ (.Y(_05352_),
    .B1(_05351_),
    .B2(net282),
    .A2(_05260_),
    .A1(net183));
 sg13g2_o21ai_1 _13134_ (.B1(_05061_),
    .Y(_05353_),
    .A1(net180),
    .A2(_05352_));
 sg13g2_a21oi_1 _13135_ (.A1(net185),
    .A2(_05348_),
    .Y(_05354_),
    .B1(_05353_));
 sg13g2_a22oi_1 _13136_ (.Y(_00439_),
    .B1(_05345_),
    .B2(_05354_),
    .A2(net59),
    .A1(_05337_));
 sg13g2_buf_1 _13137_ (.A(\clock_inst.sec_a[44] ),
    .X(_05355_));
 sg13g2_inv_1 _13138_ (.Y(_05356_),
    .A(net558));
 sg13g2_a21oi_1 _13139_ (.A1(_04822_),
    .A2(_05330_),
    .Y(_05357_),
    .B1(net371));
 sg13g2_nor2_1 _13140_ (.A(net275),
    .B(_05357_),
    .Y(_05358_));
 sg13g2_a21oi_1 _13141_ (.A1(_04822_),
    .A2(_04902_),
    .Y(_05359_),
    .B1(net284));
 sg13g2_buf_1 _13142_ (.A(_04824_),
    .X(_05360_));
 sg13g2_o21ai_1 _13143_ (.B1(net57),
    .Y(_05361_),
    .A1(_05358_),
    .A2(_05359_));
 sg13g2_o21ai_1 _13144_ (.B1(_05361_),
    .Y(_00440_),
    .A1(_05356_),
    .A2(net62));
 sg13g2_buf_2 _13145_ (.A(\clock_inst.sec_a[5] ),
    .X(_05362_));
 sg13g2_nor2_1 _13146_ (.A(net467),
    .B(_05172_),
    .Y(_05363_));
 sg13g2_nor2_1 _13147_ (.A(net268),
    .B(_05363_),
    .Y(_05364_));
 sg13g2_nand2_1 _13148_ (.Y(_05365_),
    .A(_04816_),
    .B(_04842_));
 sg13g2_buf_2 _13149_ (.A(_05365_),
    .X(_05366_));
 sg13g2_a21oi_1 _13150_ (.A1(_04959_),
    .A2(_05366_),
    .Y(_05367_),
    .B1(net259));
 sg13g2_nand2_1 _13151_ (.Y(_05368_),
    .A(_04909_),
    .B(net291));
 sg13g2_a21oi_1 _13152_ (.A1(net174),
    .A2(_05368_),
    .Y(_05369_),
    .B1(_04848_));
 sg13g2_nor3_1 _13153_ (.A(_05364_),
    .B(_05367_),
    .C(_05369_),
    .Y(_05370_));
 sg13g2_nand2_2 _13154_ (.Y(_05371_),
    .A(_04837_),
    .B(net474));
 sg13g2_nand2_1 _13155_ (.Y(_05372_),
    .A(_04855_),
    .B(_05371_));
 sg13g2_nand2_1 _13156_ (.Y(_05373_),
    .A(_04874_),
    .B(_05372_));
 sg13g2_nand2_1 _13157_ (.Y(_05374_),
    .A(_05014_),
    .B(_05373_));
 sg13g2_nor2_2 _13158_ (.A(net528),
    .B(net467),
    .Y(_05375_));
 sg13g2_a21oi_1 _13159_ (.A1(net404),
    .A2(_05375_),
    .Y(_05376_),
    .B1(net248));
 sg13g2_nand3_1 _13160_ (.B(net293),
    .C(net252),
    .A(net385),
    .Y(_05377_));
 sg13g2_o21ai_1 _13161_ (.B1(_05377_),
    .Y(_05378_),
    .A1(net276),
    .A2(_05376_));
 sg13g2_a22oi_1 _13162_ (.Y(_05379_),
    .B1(_05378_),
    .B2(net168),
    .A2(_05374_),
    .A1(_04822_));
 sg13g2_o21ai_1 _13163_ (.B1(_05379_),
    .Y(_05380_),
    .A1(net182),
    .A2(_05370_));
 sg13g2_a22oi_1 _13164_ (.Y(_05381_),
    .B1(net27),
    .B2(_05380_),
    .A2(net119),
    .A1(_05362_));
 sg13g2_inv_1 _13165_ (.Y(_00441_),
    .A(_05381_));
 sg13g2_nand2_1 _13166_ (.Y(_05382_),
    .A(_05169_),
    .B(net252));
 sg13g2_o21ai_1 _13167_ (.B1(_05382_),
    .Y(_05383_),
    .A1(net270),
    .A2(_05366_));
 sg13g2_nor2_1 _13168_ (.A(net383),
    .B(_05329_),
    .Y(_05384_));
 sg13g2_o21ai_1 _13169_ (.B1(net187),
    .Y(_05385_),
    .A1(_05225_),
    .A2(net264));
 sg13g2_nor2_2 _13170_ (.A(net399),
    .B(_05013_),
    .Y(_05386_));
 sg13g2_a21oi_1 _13171_ (.A1(net277),
    .A2(_05385_),
    .Y(_05387_),
    .B1(_05386_));
 sg13g2_a221oi_1 _13172_ (.B2(net250),
    .C1(net294),
    .B1(net287),
    .A1(net402),
    .Y(_05388_),
    .A2(net391));
 sg13g2_a21oi_1 _13173_ (.A1(net192),
    .A2(_05387_),
    .Y(_05389_),
    .B1(_05388_));
 sg13g2_a221oi_1 _13174_ (.B2(_05309_),
    .C1(_05389_),
    .B1(_05384_),
    .A1(net180),
    .Y(_05390_),
    .A2(_05383_));
 sg13g2_nand2_1 _13175_ (.Y(_05391_),
    .A(\clock_inst.sec_a[6] ),
    .B(net120));
 sg13g2_o21ai_1 _13176_ (.B1(_05391_),
    .Y(_00442_),
    .A1(net22),
    .A2(_05390_));
 sg13g2_buf_1 _13177_ (.A(\clock_inst.sec_a[7] ),
    .X(_05392_));
 sg13g2_buf_1 _13178_ (.A(net282),
    .X(_05393_));
 sg13g2_nor2_1 _13179_ (.A(net404),
    .B(_05081_),
    .Y(_05394_));
 sg13g2_a21oi_1 _13180_ (.A1(net386),
    .A2(_04881_),
    .Y(_05395_),
    .B1(_05394_));
 sg13g2_o21ai_1 _13181_ (.B1(_05234_),
    .Y(_05396_),
    .A1(_04915_),
    .A2(_05395_));
 sg13g2_o21ai_1 _13182_ (.B1(_05202_),
    .Y(_05397_),
    .A1(net374),
    .A2(net391));
 sg13g2_nand2_1 _13183_ (.Y(_05398_),
    .A(_04904_),
    .B(_05397_));
 sg13g2_nor2_1 _13184_ (.A(net266),
    .B(net169),
    .Y(_05399_));
 sg13g2_a221oi_1 _13185_ (.B2(net181),
    .C1(_05399_),
    .B1(_05398_),
    .A1(net165),
    .Y(_05400_),
    .A2(_05396_));
 sg13g2_mux2_1 _13186_ (.A0(_05392_),
    .A1(_05400_),
    .S(_04825_),
    .X(_00443_));
 sg13g2_nand2_1 _13187_ (.Y(_05401_),
    .A(_04818_),
    .B(_04810_));
 sg13g2_buf_1 _13188_ (.A(_05401_),
    .X(_05402_));
 sg13g2_nor2_1 _13189_ (.A(_05241_),
    .B(_05182_),
    .Y(_05403_));
 sg13g2_nand2_2 _13190_ (.Y(_05404_),
    .A(_04816_),
    .B(_04834_));
 sg13g2_a21oi_1 _13191_ (.A1(net396),
    .A2(_05404_),
    .Y(_05405_),
    .B1(net286));
 sg13g2_o21ai_1 _13192_ (.B1(net471),
    .Y(_05406_),
    .A1(net392),
    .A2(net459));
 sg13g2_nand3_1 _13193_ (.B(net254),
    .C(_05406_),
    .A(net386),
    .Y(_05407_));
 sg13g2_o21ai_1 _13194_ (.B1(_05407_),
    .Y(_05408_),
    .A1(net294),
    .A2(_05405_));
 sg13g2_o21ai_1 _13195_ (.B1(_05408_),
    .Y(_05409_),
    .A1(_05402_),
    .A2(_05403_));
 sg13g2_nand2_1 _13196_ (.Y(_05410_),
    .A(net524),
    .B(net525));
 sg13g2_buf_2 _13197_ (.A(_05410_),
    .X(_05411_));
 sg13g2_nand2_1 _13198_ (.Y(_05412_),
    .A(net387),
    .B(_05015_));
 sg13g2_nor2_1 _13199_ (.A(net394),
    .B(net262),
    .Y(_05413_));
 sg13g2_a22oi_1 _13200_ (.Y(_05414_),
    .B1(_05412_),
    .B2(_05413_),
    .A2(_05411_),
    .A1(net377));
 sg13g2_nand2_1 _13201_ (.Y(_05415_),
    .A(net466),
    .B(_04872_));
 sg13g2_nor2_1 _13202_ (.A(net462),
    .B(_04890_),
    .Y(_05416_));
 sg13g2_a221oi_1 _13203_ (.B2(_05416_),
    .C1(_05023_),
    .B1(_05415_),
    .A1(net253),
    .Y(_05417_),
    .A2(_05414_));
 sg13g2_o21ai_1 _13204_ (.B1(_05027_),
    .Y(_05418_),
    .A1(net290),
    .A2(net368));
 sg13g2_a22oi_1 _13205_ (.Y(_05419_),
    .B1(_05418_),
    .B2(net256),
    .A2(net380),
    .A1(_04857_));
 sg13g2_o21ai_1 _13206_ (.B1(_05419_),
    .Y(_05420_),
    .A1(net168),
    .A2(_05417_));
 sg13g2_a21oi_1 _13207_ (.A1(net116),
    .A2(_05409_),
    .Y(_05421_),
    .B1(_05420_));
 sg13g2_buf_1 _13208_ (.A(\clock_inst.sec_b[0] ),
    .X(_05422_));
 sg13g2_nand2_1 _13209_ (.Y(_05423_),
    .A(_05422_),
    .B(net120));
 sg13g2_o21ai_1 _13210_ (.B1(_05423_),
    .Y(_00444_),
    .A1(net121),
    .A2(_05421_));
 sg13g2_buf_1 _13211_ (.A(\clock_inst.sec_b[10] ),
    .X(_05424_));
 sg13g2_nand2_1 _13212_ (.Y(_05425_),
    .A(net373),
    .B(_05059_));
 sg13g2_o21ai_1 _13213_ (.B1(_05425_),
    .Y(_05426_),
    .A1(_04985_),
    .A2(_05070_));
 sg13g2_nor3_1 _13214_ (.A(net179),
    .B(net450),
    .C(_05426_),
    .Y(_05427_));
 sg13g2_a21o_1 _13215_ (.A2(net123),
    .A1(_05424_),
    .B1(_05427_),
    .X(_00445_));
 sg13g2_buf_1 _13216_ (.A(\clock_inst.sec_b[19] ),
    .X(_05428_));
 sg13g2_inv_1 _13217_ (.Y(_05429_),
    .A(_05428_));
 sg13g2_a22oi_1 _13218_ (.Y(_05430_),
    .B1(_05375_),
    .B2(net278),
    .A2(_05084_),
    .A1(_05067_));
 sg13g2_nor2_1 _13219_ (.A(_04912_),
    .B(net456),
    .Y(_05431_));
 sg13g2_buf_2 _13220_ (.A(_05431_),
    .X(_05432_));
 sg13g2_o21ai_1 _13221_ (.B1(net289),
    .Y(_05433_),
    .A1(net279),
    .A2(_05083_));
 sg13g2_nand2_1 _13222_ (.Y(_05434_),
    .A(_05432_),
    .B(_05433_));
 sg13g2_o21ai_1 _13223_ (.B1(_05434_),
    .Y(_05435_),
    .A1(net260),
    .A2(_05430_));
 sg13g2_nor2_1 _13224_ (.A(_04862_),
    .B(net403),
    .Y(_05436_));
 sg13g2_nor2_2 _13225_ (.A(net463),
    .B(_04921_),
    .Y(_05437_));
 sg13g2_a22oi_1 _13226_ (.Y(_05438_),
    .B1(_05437_),
    .B2(_04896_),
    .A2(_05436_),
    .A1(_05258_));
 sg13g2_nor2_1 _13227_ (.A(net461),
    .B(_04959_),
    .Y(_05439_));
 sg13g2_o21ai_1 _13228_ (.B1(net188),
    .Y(_05440_),
    .A1(_05343_),
    .A2(_05439_));
 sg13g2_nand3_1 _13229_ (.B(_05438_),
    .C(_05440_),
    .A(net182),
    .Y(_05441_));
 sg13g2_o21ai_1 _13230_ (.B1(_05441_),
    .Y(_05442_),
    .A1(net189),
    .A2(_05435_));
 sg13g2_a22oi_1 _13231_ (.Y(_00446_),
    .B1(net27),
    .B2(_05442_),
    .A2(net59),
    .A1(_05429_));
 sg13g2_buf_2 _13232_ (.A(\clock_inst.sec_b[1] ),
    .X(_05443_));
 sg13g2_inv_1 _13233_ (.Y(_05444_),
    .A(_05443_));
 sg13g2_nor2_1 _13234_ (.A(_04837_),
    .B(_04813_),
    .Y(_05445_));
 sg13g2_buf_2 _13235_ (.A(_05445_),
    .X(_05446_));
 sg13g2_o21ai_1 _13236_ (.B1(_05416_),
    .Y(_05447_),
    .A1(_04927_),
    .A2(_05446_));
 sg13g2_nand2_1 _13237_ (.Y(_05448_),
    .A(net61),
    .B(_05447_));
 sg13g2_a22oi_1 _13238_ (.Y(_05449_),
    .B1(net376),
    .B2(net249),
    .A2(_05245_),
    .A1(net188));
 sg13g2_nor2_1 _13239_ (.A(net118),
    .B(_05449_),
    .Y(_05450_));
 sg13g2_nor2_1 _13240_ (.A(_05448_),
    .B(_05450_),
    .Y(_05451_));
 sg13g2_a221oi_1 _13241_ (.B2(_04871_),
    .C1(_05446_),
    .B1(_05274_),
    .A1(_04961_),
    .Y(_05452_),
    .A2(_05079_));
 sg13g2_a221oi_1 _13242_ (.B2(_05102_),
    .C1(net282),
    .B1(net257),
    .A1(_05022_),
    .Y(_05453_),
    .A2(_05234_));
 sg13g2_a21oi_1 _13243_ (.A1(net260),
    .A2(_05452_),
    .Y(_05454_),
    .B1(_05453_));
 sg13g2_nand2_1 _13244_ (.Y(_05455_),
    .A(net384),
    .B(_04929_));
 sg13g2_nand2_1 _13245_ (.Y(_05456_),
    .A(net393),
    .B(_05013_));
 sg13g2_nand2_1 _13246_ (.Y(_05457_),
    .A(_04909_),
    .B(_05456_));
 sg13g2_nand2_1 _13247_ (.Y(_05458_),
    .A(_05455_),
    .B(_05457_));
 sg13g2_nor2_1 _13248_ (.A(net475),
    .B(net400),
    .Y(_05459_));
 sg13g2_buf_2 _13249_ (.A(_05459_),
    .X(_05460_));
 sg13g2_a22oi_1 _13250_ (.Y(_05461_),
    .B1(_05458_),
    .B2(_05460_),
    .A2(_05436_),
    .A1(net283));
 sg13g2_nand2_1 _13251_ (.Y(_05462_),
    .A(net185),
    .B(_05461_));
 sg13g2_o21ai_1 _13252_ (.B1(_05462_),
    .Y(_05463_),
    .A1(net185),
    .A2(_05454_));
 sg13g2_a22oi_1 _13253_ (.Y(_00447_),
    .B1(_05451_),
    .B2(_05463_),
    .A2(net59),
    .A1(_05444_));
 sg13g2_nand2_1 _13254_ (.Y(_05464_),
    .A(_04951_),
    .B(net174));
 sg13g2_o21ai_1 _13255_ (.B1(_05464_),
    .Y(_05465_),
    .A1(net294),
    .A2(net166));
 sg13g2_a22oi_1 _13256_ (.Y(_05466_),
    .B1(_05465_),
    .B2(net292),
    .A2(net167),
    .A1(_05062_));
 sg13g2_inv_1 _13257_ (.Y(_05467_),
    .A(_05436_));
 sg13g2_o21ai_1 _13258_ (.B1(_05467_),
    .Y(_05468_),
    .A1(net397),
    .A2(_04840_));
 sg13g2_a221oi_1 _13259_ (.B2(_05231_),
    .C1(net179),
    .B1(_05468_),
    .A1(net167),
    .Y(_05469_),
    .A2(_05437_));
 sg13g2_a21oi_1 _13260_ (.A1(net179),
    .A2(_05466_),
    .Y(_05470_),
    .B1(_05469_));
 sg13g2_nand2_1 _13261_ (.Y(_05471_),
    .A(\clock_inst.sec_b[20] ),
    .B(_05002_));
 sg13g2_o21ai_1 _13262_ (.B1(_05471_),
    .Y(_00448_),
    .A1(_05006_),
    .A2(_05470_));
 sg13g2_buf_2 _13263_ (.A(\clock_inst.sec_b[2] ),
    .X(_05472_));
 sg13g2_o21ai_1 _13264_ (.B1(_04853_),
    .Y(_05473_),
    .A1(net370),
    .A2(_05172_));
 sg13g2_nand2_1 _13265_ (.Y(_05474_),
    .A(_05366_),
    .B(_05473_));
 sg13g2_buf_1 _13266_ (.A(net253),
    .X(_05475_));
 sg13g2_nor2_1 _13267_ (.A(net466),
    .B(_05013_),
    .Y(_05476_));
 sg13g2_a221oi_1 _13268_ (.B2(net164),
    .C1(_05476_),
    .B1(_05474_),
    .A1(net115),
    .Y(_05477_),
    .A2(_05080_));
 sg13g2_nand2_1 _13269_ (.Y(_05478_),
    .A(net285),
    .B(_04815_));
 sg13g2_o21ai_1 _13270_ (.B1(_05079_),
    .Y(_05479_),
    .A1(_05156_),
    .A2(_05172_));
 sg13g2_o21ai_1 _13271_ (.B1(_05083_),
    .Y(_05480_),
    .A1(_04887_),
    .A2(net393));
 sg13g2_nand2_1 _13272_ (.Y(_05481_),
    .A(_04914_),
    .B(_05480_));
 sg13g2_nand4_1 _13273_ (.B(_05478_),
    .C(_05479_),
    .A(_05009_),
    .Y(_05482_),
    .D(_05481_));
 sg13g2_a22oi_1 _13274_ (.Y(_05483_),
    .B1(_05482_),
    .B2(_05320_),
    .A2(_04946_),
    .A1(_04941_));
 sg13g2_o21ai_1 _13275_ (.B1(_05483_),
    .Y(_05484_),
    .A1(net180),
    .A2(_05477_));
 sg13g2_a22oi_1 _13276_ (.Y(_05485_),
    .B1(net27),
    .B2(_05484_),
    .A2(net119),
    .A1(_05472_));
 sg13g2_inv_1 _13277_ (.Y(_00449_),
    .A(_05485_));
 sg13g2_buf_1 _13278_ (.A(\clock_inst.sec_b[21] ),
    .X(_05486_));
 sg13g2_inv_1 _13279_ (.Y(_05487_),
    .A(net557));
 sg13g2_or3_1 _13280_ (.A(net191),
    .B(_04948_),
    .C(_05358_),
    .X(_05488_));
 sg13g2_o21ai_1 _13281_ (.B1(_05488_),
    .Y(_00450_),
    .A1(net522),
    .A2(net62));
 sg13g2_buf_8 _13282_ (.A(\clock_inst.sec_b[36] ),
    .X(_05489_));
 sg13g2_inv_1 _13283_ (.Y(_05490_),
    .A(_05489_));
 sg13g2_nor2_1 _13284_ (.A(net375),
    .B(net177),
    .Y(_05491_));
 sg13g2_nand2_1 _13285_ (.Y(_05492_),
    .A(net528),
    .B(net388));
 sg13g2_nor2_1 _13286_ (.A(net271),
    .B(net368),
    .Y(_05493_));
 sg13g2_a221oi_1 _13287_ (.B2(_05493_),
    .C1(_05043_),
    .B1(_05492_),
    .A1(_05478_),
    .Y(_05494_),
    .A2(_05491_));
 sg13g2_nor2_1 _13288_ (.A(net273),
    .B(net388),
    .Y(_05495_));
 sg13g2_o21ai_1 _13289_ (.B1(net398),
    .Y(_05496_),
    .A1(_04865_),
    .A2(_05015_));
 sg13g2_a21oi_1 _13290_ (.A1(net289),
    .A2(_05496_),
    .Y(_05497_),
    .B1(net379));
 sg13g2_a221oi_1 _13291_ (.B2(net250),
    .C1(_05497_),
    .B1(_05495_),
    .A1(net173),
    .Y(_05498_),
    .A2(_05150_));
 sg13g2_o21ai_1 _13292_ (.B1(net390),
    .Y(_05499_),
    .A1(net383),
    .A2(_05023_));
 sg13g2_a21oi_1 _13293_ (.A1(net384),
    .A2(net248),
    .Y(_05500_),
    .B1(_05375_));
 sg13g2_a21oi_1 _13294_ (.A1(_05499_),
    .A2(_05500_),
    .Y(_05501_),
    .B1(net253));
 sg13g2_a21oi_1 _13295_ (.A1(_04971_),
    .A2(_05039_),
    .Y(_05502_),
    .B1(net259));
 sg13g2_nor3_1 _13296_ (.A(net270),
    .B(_05501_),
    .C(_05502_),
    .Y(_05503_));
 sg13g2_a21oi_1 _13297_ (.A1(net192),
    .A2(_05498_),
    .Y(_05504_),
    .B1(_05503_));
 sg13g2_o21ai_1 _13298_ (.B1(_04824_),
    .Y(_05505_),
    .A1(_05494_),
    .A2(_05504_));
 sg13g2_o21ai_1 _13299_ (.B1(_05505_),
    .Y(_00451_),
    .A1(_05490_),
    .A2(net62));
 sg13g2_buf_8 _13300_ (.A(\clock_inst.sec_b[37] ),
    .X(_05506_));
 sg13g2_inv_1 _13301_ (.Y(_05507_),
    .A(_05506_));
 sg13g2_nand2_1 _13302_ (.Y(_05508_),
    .A(net404),
    .B(net258));
 sg13g2_o21ai_1 _13303_ (.B1(_05508_),
    .Y(_05509_),
    .A1(net397),
    .A2(_05274_));
 sg13g2_nor2_2 _13304_ (.A(net458),
    .B(net289),
    .Y(_05510_));
 sg13g2_a21o_1 _13305_ (.A2(_05509_),
    .A1(net272),
    .B1(_05510_),
    .X(_05511_));
 sg13g2_nand2_1 _13306_ (.Y(_05512_),
    .A(net466),
    .B(net462));
 sg13g2_o21ai_1 _13307_ (.B1(_05116_),
    .Y(_05513_),
    .A1(net256),
    .A2(_05512_));
 sg13g2_o21ai_1 _13308_ (.B1(_04967_),
    .Y(_05514_),
    .A1(_05292_),
    .A2(_05513_));
 sg13g2_nand2_1 _13309_ (.Y(_05515_),
    .A(_04898_),
    .B(_05172_));
 sg13g2_a21oi_1 _13310_ (.A1(_05025_),
    .A2(_05515_),
    .Y(_05516_),
    .B1(_05151_));
 sg13g2_a21oi_1 _13311_ (.A1(_05160_),
    .A2(net267),
    .Y(_05517_),
    .B1(_05516_));
 sg13g2_nand3_1 _13312_ (.B(_05514_),
    .C(_05517_),
    .A(_05244_),
    .Y(_05518_));
 sg13g2_a21oi_1 _13313_ (.A1(net165),
    .A2(_05511_),
    .Y(_05519_),
    .B1(_05518_));
 sg13g2_a21oi_1 _13314_ (.A1(_05507_),
    .A2(net60),
    .Y(_00452_),
    .B1(_05519_));
 sg13g2_buf_2 _13315_ (.A(\clock_inst.sec_b[38] ),
    .X(_05520_));
 sg13g2_a22oi_1 _13316_ (.Y(_05521_),
    .B1(net287),
    .B2(_05033_),
    .A2(_04852_),
    .A1(net367));
 sg13g2_nand2_1 _13317_ (.Y(_05522_),
    .A(_04867_),
    .B(net528));
 sg13g2_nand2_1 _13318_ (.Y(_05523_),
    .A(net383),
    .B(_05522_));
 sg13g2_a221oi_1 _13319_ (.B2(_05100_),
    .C1(net268),
    .B1(_05523_),
    .A1(net279),
    .Y(_05524_),
    .A2(_05323_));
 sg13g2_a21oi_1 _13320_ (.A1(net178),
    .A2(_05521_),
    .Y(_05525_),
    .B1(_05524_));
 sg13g2_nand3_1 _13321_ (.B(net269),
    .C(_04925_),
    .A(net397),
    .Y(_05526_));
 sg13g2_nand2_1 _13322_ (.Y(_05527_),
    .A(_05027_),
    .B(_05182_));
 sg13g2_a21oi_1 _13323_ (.A1(_05526_),
    .A2(_05527_),
    .Y(_05528_),
    .B1(net168));
 sg13g2_nand2_2 _13324_ (.Y(_05529_),
    .A(net524),
    .B(_04815_));
 sg13g2_nand2_1 _13325_ (.Y(_05530_),
    .A(net61),
    .B(_05529_));
 sg13g2_nand2_1 _13326_ (.Y(_05531_),
    .A(_05161_),
    .B(_05211_));
 sg13g2_nand2_1 _13327_ (.Y(_05532_),
    .A(net293),
    .B(_05072_));
 sg13g2_a22oi_1 _13328_ (.Y(_05533_),
    .B1(_05532_),
    .B2(net115),
    .A2(_05531_),
    .A1(net294));
 sg13g2_nor2_1 _13329_ (.A(net260),
    .B(_05533_),
    .Y(_05534_));
 sg13g2_nor4_1 _13330_ (.A(_05525_),
    .B(_05528_),
    .C(_05530_),
    .D(_05534_),
    .Y(_05535_));
 sg13g2_a21o_1 _13331_ (.A2(net123),
    .A1(_05520_),
    .B1(_05535_),
    .X(_00453_));
 sg13g2_buf_2 _13332_ (.A(\clock_inst.sec_b[39] ),
    .X(_05536_));
 sg13g2_a21oi_1 _13333_ (.A1(net404),
    .A2(net368),
    .Y(_05537_),
    .B1(net248));
 sg13g2_o21ai_1 _13334_ (.B1(_05537_),
    .Y(_05538_),
    .A1(net386),
    .A2(_05456_));
 sg13g2_a22oi_1 _13335_ (.Y(_05539_),
    .B1(_05538_),
    .B2(net188),
    .A2(net369),
    .A1(net183));
 sg13g2_nand2_1 _13336_ (.Y(_05540_),
    .A(net393),
    .B(_05260_));
 sg13g2_o21ai_1 _13337_ (.B1(_04914_),
    .Y(_05541_),
    .A1(net172),
    .A2(_04892_));
 sg13g2_nand2_1 _13338_ (.Y(_05542_),
    .A(_05540_),
    .B(_05541_));
 sg13g2_o21ai_1 _13339_ (.B1(_04959_),
    .Y(_05543_),
    .A1(_05154_),
    .A2(_05158_));
 sg13g2_a22oi_1 _13340_ (.Y(_05544_),
    .B1(_05543_),
    .B2(net287),
    .A2(_05542_),
    .A1(net249));
 sg13g2_o21ai_1 _13341_ (.B1(_05544_),
    .Y(_05545_),
    .A1(_05134_),
    .A2(_05539_));
 sg13g2_a22oi_1 _13342_ (.Y(_05546_),
    .B1(_05092_),
    .B2(_05545_),
    .A2(_05091_),
    .A1(_05536_));
 sg13g2_inv_1 _13343_ (.Y(_00454_),
    .A(_05546_));
 sg13g2_o21ai_1 _13344_ (.B1(net169),
    .Y(_05547_),
    .A1(net378),
    .A2(_05027_));
 sg13g2_a21oi_1 _13345_ (.A1(net294),
    .A2(_05495_),
    .Y(_05548_),
    .B1(_05547_));
 sg13g2_o21ai_1 _13346_ (.B1(_05460_),
    .Y(_05549_),
    .A1(_05214_),
    .A2(net370));
 sg13g2_o21ai_1 _13347_ (.B1(_05549_),
    .Y(_05550_),
    .A1(net184),
    .A2(_05548_));
 sg13g2_a21oi_1 _13348_ (.A1(net284),
    .A2(_05224_),
    .Y(_05551_),
    .B1(net175));
 sg13g2_nor2_1 _13349_ (.A(_05229_),
    .B(_05551_),
    .Y(_05552_));
 sg13g2_a21oi_1 _13350_ (.A1(net174),
    .A2(_05492_),
    .Y(_05553_),
    .B1(_04966_));
 sg13g2_a21oi_1 _13351_ (.A1(net382),
    .A2(net174),
    .Y(_05554_),
    .B1(net261));
 sg13g2_o21ai_1 _13352_ (.B1(net283),
    .Y(_05555_),
    .A1(_05553_),
    .A2(_05554_));
 sg13g2_o21ai_1 _13353_ (.B1(_05555_),
    .Y(_05556_),
    .A1(net168),
    .A2(_05552_));
 sg13g2_a21oi_1 _13354_ (.A1(net116),
    .A2(_05550_),
    .Y(_05557_),
    .B1(_05556_));
 sg13g2_buf_1 _13355_ (.A(\clock_inst.sec_b[3] ),
    .X(_05558_));
 sg13g2_buf_1 _13356_ (.A(net191),
    .X(_05559_));
 sg13g2_nand2_1 _13357_ (.Y(_05560_),
    .A(_05558_),
    .B(net114));
 sg13g2_o21ai_1 _13358_ (.B1(_05560_),
    .Y(_00455_),
    .A1(net22),
    .A2(_05557_));
 sg13g2_buf_2 _13359_ (.A(\clock_inst.sec_b[40] ),
    .X(_05561_));
 sg13g2_a21oi_1 _13360_ (.A1(_05079_),
    .A2(_05016_),
    .Y(_05562_),
    .B1(_05338_));
 sg13g2_o21ai_1 _13361_ (.B1(_05247_),
    .Y(_05563_),
    .A1(net374),
    .A2(_04906_));
 sg13g2_o21ai_1 _13362_ (.B1(_05563_),
    .Y(_05564_),
    .A1(net117),
    .A2(_05562_));
 sg13g2_nand2_1 _13363_ (.Y(_05565_),
    .A(_04925_),
    .B(_05027_));
 sg13g2_a22oi_1 _13364_ (.Y(_05566_),
    .B1(_05565_),
    .B2(net263),
    .A2(_04946_),
    .A1(_04906_));
 sg13g2_nor2_1 _13365_ (.A(net285),
    .B(_05456_),
    .Y(_05567_));
 sg13g2_nor2_1 _13366_ (.A(net458),
    .B(_04842_),
    .Y(_05568_));
 sg13g2_nor3_1 _13367_ (.A(net471),
    .B(_05305_),
    .C(_05568_),
    .Y(_05569_));
 sg13g2_o21ai_1 _13368_ (.B1(net190),
    .Y(_05570_),
    .A1(_05567_),
    .A2(_05569_));
 sg13g2_o21ai_1 _13369_ (.B1(_05570_),
    .Y(_05571_),
    .A1(_04967_),
    .A2(_05566_));
 sg13g2_a221oi_1 _13370_ (.B2(net180),
    .C1(_05571_),
    .B1(_05564_),
    .A1(net166),
    .Y(_05572_),
    .A2(net380));
 sg13g2_mux2_1 _13371_ (.A0(_05561_),
    .A1(_05572_),
    .S(net62),
    .X(_00456_));
 sg13g2_buf_2 _13372_ (.A(\clock_inst.sec_b[41] ),
    .X(_05573_));
 sg13g2_nand3_1 _13373_ (.B(_05037_),
    .C(_05460_),
    .A(_05025_),
    .Y(_05574_));
 sg13g2_o21ai_1 _13374_ (.B1(_05574_),
    .Y(_05575_),
    .A1(_04844_),
    .A2(_05037_));
 sg13g2_o21ai_1 _13375_ (.B1(_04913_),
    .Y(_05576_),
    .A1(net383),
    .A2(_04836_));
 sg13g2_a21oi_1 _13376_ (.A1(_05014_),
    .A2(_05576_),
    .Y(_05577_),
    .B1(net286));
 sg13g2_a21oi_1 _13377_ (.A1(_05019_),
    .A2(net276),
    .Y(_05578_),
    .B1(net281));
 sg13g2_or3_1 _13378_ (.A(_05416_),
    .B(_05577_),
    .C(_05578_),
    .X(_05579_));
 sg13g2_a21oi_1 _13379_ (.A1(net397),
    .A2(_05205_),
    .Y(_05580_),
    .B1(_04822_));
 sg13g2_nor2_1 _13380_ (.A(_04850_),
    .B(_05446_),
    .Y(_05581_));
 sg13g2_nand3_1 _13381_ (.B(_05079_),
    .C(_05581_),
    .A(net115),
    .Y(_05582_));
 sg13g2_o21ai_1 _13382_ (.B1(_05582_),
    .Y(_05583_),
    .A1(net171),
    .A2(_05580_));
 sg13g2_a221oi_1 _13383_ (.B2(net182),
    .C1(_05583_),
    .B1(_05579_),
    .A1(net165),
    .Y(_05584_),
    .A2(_05575_));
 sg13g2_mux2_1 _13384_ (.A0(_05573_),
    .A1(_05584_),
    .S(net57),
    .X(_00457_));
 sg13g2_o21ai_1 _13385_ (.B1(net263),
    .Y(_05585_),
    .A1(_05042_),
    .A2(_04852_));
 sg13g2_nand2b_1 _13386_ (.Y(_05586_),
    .B(_05585_),
    .A_N(_04993_));
 sg13g2_a22oi_1 _13387_ (.Y(_05587_),
    .B1(net261),
    .B2(_05144_),
    .A2(net284),
    .A1(net259));
 sg13g2_o21ai_1 _13388_ (.B1(_05366_),
    .Y(_05588_),
    .A1(net178),
    .A2(_05587_));
 sg13g2_a21o_1 _13389_ (.A2(_05187_),
    .A1(net174),
    .B1(net397),
    .X(_05589_));
 sg13g2_a21oi_1 _13390_ (.A1(_05368_),
    .A2(_05589_),
    .Y(_05590_),
    .B1(_05136_));
 sg13g2_a221oi_1 _13391_ (.B2(net182),
    .C1(_05590_),
    .B1(_05588_),
    .A1(net370),
    .Y(_05591_),
    .A2(_05586_));
 sg13g2_nand2_1 _13392_ (.Y(_05592_),
    .A(\clock_inst.sec_b[42] ),
    .B(net114));
 sg13g2_o21ai_1 _13393_ (.B1(_05592_),
    .Y(_00458_),
    .A1(net22),
    .A2(_05591_));
 sg13g2_buf_1 _13394_ (.A(\clock_inst.sec_b[43] ),
    .X(_05593_));
 sg13g2_inv_1 _13395_ (.Y(_05594_),
    .A(_05593_));
 sg13g2_nand2_2 _13396_ (.Y(_05595_),
    .A(net383),
    .B(_04902_));
 sg13g2_a21oi_1 _13397_ (.A1(net166),
    .A2(_05595_),
    .Y(_05596_),
    .B1(net376));
 sg13g2_nor3_1 _13398_ (.A(_04915_),
    .B(net287),
    .C(_05229_),
    .Y(_05597_));
 sg13g2_a21oi_1 _13399_ (.A1(_04849_),
    .A2(_05596_),
    .Y(_05598_),
    .B1(_05597_));
 sg13g2_nand2_1 _13400_ (.Y(_05599_),
    .A(_04828_),
    .B(net399));
 sg13g2_a21oi_1 _13401_ (.A1(net278),
    .A2(_05432_),
    .Y(_05600_),
    .B1(net171));
 sg13g2_nor2_1 _13402_ (.A(_05599_),
    .B(_05600_),
    .Y(_05601_));
 sg13g2_o21ai_1 _13403_ (.B1(net61),
    .Y(_05602_),
    .A1(_05598_),
    .A2(_05601_));
 sg13g2_o21ai_1 _13404_ (.B1(_05602_),
    .Y(_00459_),
    .A1(_05594_),
    .A2(_04825_));
 sg13g2_o21ai_1 _13405_ (.B1(net279),
    .Y(_05603_),
    .A1(net385),
    .A2(net401));
 sg13g2_a21oi_1 _13406_ (.A1(_05081_),
    .A2(_05603_),
    .Y(_05604_),
    .B1(net117));
 sg13g2_o21ai_1 _13407_ (.B1(net176),
    .Y(_05605_),
    .A1(_05510_),
    .A2(_05604_));
 sg13g2_o21ai_1 _13408_ (.B1(_05200_),
    .Y(_05606_),
    .A1(net276),
    .A2(_05522_));
 sg13g2_nor2_1 _13409_ (.A(net530),
    .B(net527),
    .Y(_05607_));
 sg13g2_a22oi_1 _13410_ (.Y(_05608_),
    .B1(_05270_),
    .B2(_05607_),
    .A2(net258),
    .A1(net382));
 sg13g2_o21ai_1 _13411_ (.B1(_05338_),
    .Y(_05609_),
    .A1(_05305_),
    .A2(_05192_));
 sg13g2_a21oi_1 _13412_ (.A1(_05608_),
    .A2(_05609_),
    .Y(_05610_),
    .B1(net288));
 sg13g2_a221oi_1 _13413_ (.B2(net249),
    .C1(_05610_),
    .B1(_05606_),
    .A1(net272),
    .Y(_05611_),
    .A2(net256));
 sg13g2_nand2_1 _13414_ (.Y(_05612_),
    .A(_05605_),
    .B(_05611_));
 sg13g2_buf_1 _13415_ (.A(\clock_inst.sec_b[4] ),
    .X(_05613_));
 sg13g2_nand2_1 _13416_ (.Y(_05614_),
    .A(_05613_),
    .B(_05559_));
 sg13g2_o21ai_1 _13417_ (.B1(_05614_),
    .Y(_00460_),
    .A1(net121),
    .A2(_05612_));
 sg13g2_buf_1 _13418_ (.A(\clock_inst.sec_b[5] ),
    .X(_05615_));
 sg13g2_buf_1 _13419_ (.A(net281),
    .X(_05616_));
 sg13g2_a21oi_1 _13420_ (.A1(_05334_),
    .A2(_05275_),
    .Y(_05617_),
    .B1(net252));
 sg13g2_o21ai_1 _13421_ (.B1(_05039_),
    .Y(_05618_),
    .A1(_05013_),
    .A2(_05037_));
 sg13g2_nor3_1 _13422_ (.A(net471),
    .B(_04902_),
    .C(_05016_),
    .Y(_05619_));
 sg13g2_a221oi_1 _13423_ (.B2(_04996_),
    .C1(_05619_),
    .B1(_05618_),
    .A1(net177),
    .Y(_05620_),
    .A2(_05595_));
 sg13g2_nor2_1 _13424_ (.A(_05023_),
    .B(_05155_),
    .Y(_05621_));
 sg13g2_o21ai_1 _13425_ (.B1(_05529_),
    .Y(_05622_),
    .A1(_04874_),
    .A2(_05621_));
 sg13g2_o21ai_1 _13426_ (.B1(net458),
    .Y(_05623_),
    .A1(_04828_),
    .A2(_05204_));
 sg13g2_nand2_1 _13427_ (.Y(_05624_),
    .A(_05402_),
    .B(_05404_));
 sg13g2_nand2_1 _13428_ (.Y(_05625_),
    .A(net475),
    .B(_05624_));
 sg13g2_a21oi_1 _13429_ (.A1(_05623_),
    .A2(_05625_),
    .Y(_05626_),
    .B1(_04873_));
 sg13g2_a221oi_1 _13430_ (.B2(net281),
    .C1(_05626_),
    .B1(_05622_),
    .A1(net381),
    .Y(_05627_),
    .A2(_04839_));
 sg13g2_mux2_1 _13431_ (.A0(_05620_),
    .A1(_05627_),
    .S(net164),
    .X(_05628_));
 sg13g2_o21ai_1 _13432_ (.B1(_05628_),
    .Y(_05629_),
    .A1(_05616_),
    .A2(_05617_));
 sg13g2_a22oi_1 _13433_ (.Y(_05630_),
    .B1(net27),
    .B2(_05629_),
    .A2(net119),
    .A1(_05615_));
 sg13g2_inv_1 _13434_ (.Y(_00461_),
    .A(_05630_));
 sg13g2_buf_1 _13435_ (.A(\clock_inst.sec_b[6] ),
    .X(_05631_));
 sg13g2_inv_1 _13436_ (.Y(_05632_),
    .A(_05631_));
 sg13g2_nor2_1 _13437_ (.A(net400),
    .B(net388),
    .Y(_05633_));
 sg13g2_nor2_1 _13438_ (.A(net259),
    .B(_05039_),
    .Y(_05634_));
 sg13g2_nand2_1 _13439_ (.Y(_05635_),
    .A(net465),
    .B(_04944_));
 sg13g2_a21oi_1 _13440_ (.A1(_05635_),
    .A2(_05368_),
    .Y(_05636_),
    .B1(net275));
 sg13g2_nor4_1 _13441_ (.A(net249),
    .B(_05633_),
    .C(_05634_),
    .D(_05636_),
    .Y(_05637_));
 sg13g2_a21o_1 _13442_ (.A2(_04991_),
    .A1(net374),
    .B1(net402),
    .X(_05638_));
 sg13g2_a21oi_1 _13443_ (.A1(net251),
    .A2(net287),
    .Y(_05639_),
    .B1(net253));
 sg13g2_nand2_1 _13444_ (.Y(_05640_),
    .A(net274),
    .B(net369));
 sg13g2_a221oi_1 _13445_ (.B2(_05063_),
    .C1(_05203_),
    .B1(_05640_),
    .A1(_05638_),
    .Y(_05641_),
    .A2(_05639_));
 sg13g2_nor4_1 _13446_ (.A(net191),
    .B(_05126_),
    .C(_05637_),
    .D(_05641_),
    .Y(_05642_));
 sg13g2_a21oi_1 _13447_ (.A1(_05632_),
    .A2(net60),
    .Y(_00462_),
    .B1(_05642_));
 sg13g2_buf_1 _13448_ (.A(\clock_inst.sec_b[7] ),
    .X(_05643_));
 sg13g2_nand3_1 _13449_ (.B(_05402_),
    .C(_05404_),
    .A(net373),
    .Y(_05644_));
 sg13g2_a21oi_1 _13450_ (.A1(_05412_),
    .A2(_05644_),
    .Y(_05645_),
    .B1(net184));
 sg13g2_a21oi_1 _13451_ (.A1(_04991_),
    .A2(net169),
    .Y(_05646_),
    .B1(_05599_));
 sg13g2_nor4_1 _13452_ (.A(_05128_),
    .B(_05567_),
    .C(_05645_),
    .D(_05646_),
    .Y(_05647_));
 sg13g2_mux2_1 _13453_ (.A0(_05643_),
    .A1(_05647_),
    .S(net57),
    .X(_00463_));
 sg13g2_inv_1 _13454_ (.Y(_05648_),
    .A(\clock_inst.sec_c[0] ));
 sg13g2_nand2_1 _13455_ (.Y(_05649_),
    .A(net187),
    .B(_05529_));
 sg13g2_a22oi_1 _13456_ (.Y(_05650_),
    .B1(_05649_),
    .B2(net270),
    .A2(net380),
    .A1(net183));
 sg13g2_o21ai_1 _13457_ (.B1(_05182_),
    .Y(_05651_),
    .A1(_05432_),
    .A2(_05491_));
 sg13g2_o21ai_1 _13458_ (.B1(_05651_),
    .Y(_05652_),
    .A1(net168),
    .A2(_05650_));
 sg13g2_a22oi_1 _13459_ (.Y(_05653_),
    .B1(net370),
    .B2(net167),
    .A2(net262),
    .A1(net281));
 sg13g2_nor2_1 _13460_ (.A(net456),
    .B(_05653_),
    .Y(_05654_));
 sg13g2_a21oi_1 _13461_ (.A1(_04896_),
    .A2(net284),
    .Y(_05655_),
    .B1(net263));
 sg13g2_o21ai_1 _13462_ (.B1(net288),
    .Y(_05656_),
    .A1(net403),
    .A2(_05655_));
 sg13g2_nand3b_1 _13463_ (.B(net118),
    .C(_05656_),
    .Y(_05657_),
    .A_N(_05654_));
 sg13g2_o21ai_1 _13464_ (.B1(_05657_),
    .Y(_05658_),
    .A1(net118),
    .A2(_05652_));
 sg13g2_a22oi_1 _13465_ (.Y(_00464_),
    .B1(_05055_),
    .B2(_05658_),
    .A2(net59),
    .A1(_05648_));
 sg13g2_inv_1 _13466_ (.Y(_05659_),
    .A(\clock_inst.sec_c[10] ));
 sg13g2_nor3_1 _13467_ (.A(net279),
    .B(net286),
    .C(_05432_),
    .Y(_05660_));
 sg13g2_a21oi_1 _13468_ (.A1(net278),
    .A2(_05173_),
    .Y(_05661_),
    .B1(_05660_));
 sg13g2_nor2_1 _13469_ (.A(net171),
    .B(_05661_),
    .Y(_05662_));
 sg13g2_o21ai_1 _13470_ (.B1(net189),
    .Y(_05663_),
    .A1(_05128_),
    .A2(_05662_));
 sg13g2_a21oi_1 _13471_ (.A1(_05064_),
    .A2(_05123_),
    .Y(_05664_),
    .B1(_05432_));
 sg13g2_o21ai_1 _13472_ (.B1(_05540_),
    .Y(_05665_),
    .A1(_04831_),
    .A2(_05664_));
 sg13g2_a22oi_1 _13473_ (.Y(_05666_),
    .B1(net370),
    .B2(_05100_),
    .A2(net262),
    .A1(net250));
 sg13g2_nand2b_1 _13474_ (.Y(_05667_),
    .B(_05666_),
    .A_N(_05448_));
 sg13g2_a21oi_1 _13475_ (.A1(_05250_),
    .A2(_05665_),
    .Y(_05668_),
    .B1(_05667_));
 sg13g2_a22oi_1 _13476_ (.Y(_00465_),
    .B1(_05663_),
    .B2(_05668_),
    .A2(_05319_),
    .A1(_05659_));
 sg13g2_a21oi_1 _13477_ (.A1(net396),
    .A2(_04890_),
    .Y(_05669_),
    .B1(net378));
 sg13g2_o21ai_1 _13478_ (.B1(net115),
    .Y(_05670_),
    .A1(net258),
    .A2(_05669_));
 sg13g2_nand2_1 _13479_ (.Y(_05671_),
    .A(net266),
    .B(_05275_));
 sg13g2_a21oi_1 _13480_ (.A1(_05670_),
    .A2(_05671_),
    .Y(_05672_),
    .B1(net168));
 sg13g2_nand2_1 _13481_ (.Y(_05673_),
    .A(net378),
    .B(_04907_));
 sg13g2_nand2_1 _13482_ (.Y(_05674_),
    .A(_05215_),
    .B(_05415_));
 sg13g2_a22oi_1 _13483_ (.Y(_05675_),
    .B1(_05674_),
    .B2(net288),
    .A2(_05446_),
    .A1(_05673_));
 sg13g2_a21oi_1 _13484_ (.A1(_04972_),
    .A2(_04907_),
    .Y(_05676_),
    .B1(_04872_));
 sg13g2_o21ai_1 _13485_ (.B1(_05373_),
    .Y(_05677_),
    .A1(_04853_),
    .A2(_05676_));
 sg13g2_a21o_1 _13486_ (.A2(_05305_),
    .A1(net404),
    .B1(_05132_),
    .X(_05678_));
 sg13g2_a221oi_1 _13487_ (.B2(net371),
    .C1(net190),
    .B1(_05678_),
    .A1(net402),
    .Y(_05679_),
    .A2(_05677_));
 sg13g2_a21oi_1 _13488_ (.A1(net184),
    .A2(_05675_),
    .Y(_05680_),
    .B1(_05679_));
 sg13g2_nor3_1 _13489_ (.A(net122),
    .B(_05672_),
    .C(_05680_),
    .Y(_05681_));
 sg13g2_a21o_1 _13490_ (.A2(_04937_),
    .A1(\clock_inst.sec_c[11] ),
    .B1(_05681_),
    .X(_00466_));
 sg13g2_inv_1 _13491_ (.Y(_05682_),
    .A(\clock_inst.sec_c[12] ));
 sg13g2_nand2_1 _13492_ (.Y(_05683_),
    .A(net167),
    .B(_05633_));
 sg13g2_nor2_1 _13493_ (.A(net395),
    .B(_05168_),
    .Y(_05684_));
 sg13g2_nand2_1 _13494_ (.Y(_05685_),
    .A(net398),
    .B(_05684_));
 sg13g2_o21ai_1 _13495_ (.B1(_05685_),
    .Y(_05686_),
    .A1(net382),
    .A2(net291));
 sg13g2_a21o_1 _13496_ (.A2(_05295_),
    .A1(net394),
    .B1(_05195_),
    .X(_05687_));
 sg13g2_a22oi_1 _13497_ (.Y(_05688_),
    .B1(_05687_),
    .B2(net280),
    .A2(net267),
    .A1(net395));
 sg13g2_o21ai_1 _13498_ (.B1(_05688_),
    .Y(_05689_),
    .A1(net294),
    .A2(_05686_));
 sg13g2_o21ai_1 _13499_ (.B1(net286),
    .Y(_05690_),
    .A1(net396),
    .A2(_05329_));
 sg13g2_o21ai_1 _13500_ (.B1(net381),
    .Y(_05691_),
    .A1(net264),
    .A2(net403));
 sg13g2_nand4_1 _13501_ (.B(_05107_),
    .C(_05690_),
    .A(net288),
    .Y(_05692_),
    .D(_05691_));
 sg13g2_o21ai_1 _13502_ (.B1(_05692_),
    .Y(_05693_),
    .A1(net292),
    .A2(_05689_));
 sg13g2_nand4_1 _13503_ (.B(_04930_),
    .C(_05683_),
    .A(_04824_),
    .Y(_05694_),
    .D(_05693_));
 sg13g2_o21ai_1 _13504_ (.B1(_05694_),
    .Y(_00467_),
    .A1(_05682_),
    .A2(net62));
 sg13g2_inv_1 _13505_ (.Y(_05695_),
    .A(\clock_inst.sec_c[13] ));
 sg13g2_nand2_1 _13506_ (.Y(_05696_),
    .A(_05168_),
    .B(_05204_));
 sg13g2_o21ai_1 _13507_ (.B1(_05696_),
    .Y(_05697_),
    .A1(net460),
    .A2(net274));
 sg13g2_nand2b_1 _13508_ (.Y(_05698_),
    .B(_04932_),
    .A_N(_05054_));
 sg13g2_a21oi_1 _13509_ (.A1(_04876_),
    .A2(_05697_),
    .Y(_05699_),
    .B1(_05698_));
 sg13g2_o21ai_1 _13510_ (.B1(_05699_),
    .Y(_05700_),
    .A1(_05208_),
    .A2(_05384_));
 sg13g2_nor2_2 _13511_ (.A(net377),
    .B(net400),
    .Y(_05701_));
 sg13g2_o21ai_1 _13512_ (.B1(_05027_),
    .Y(_05702_),
    .A1(net378),
    .A2(_05039_));
 sg13g2_a22oi_1 _13513_ (.Y(_05703_),
    .B1(_05702_),
    .B2(_04881_),
    .A2(_05624_),
    .A1(_05701_));
 sg13g2_buf_1 _13514_ (.A(_04994_),
    .X(_05704_));
 sg13g2_nor2_1 _13515_ (.A(net379),
    .B(net247),
    .Y(_05705_));
 sg13g2_o21ai_1 _13516_ (.B1(_05446_),
    .Y(_05706_),
    .A1(_05437_),
    .A2(_05705_));
 sg13g2_o21ai_1 _13517_ (.B1(_05706_),
    .Y(_05707_),
    .A1(net275),
    .A2(_05703_));
 sg13g2_o21ai_1 _13518_ (.B1(_05083_),
    .Y(_05708_),
    .A1(net377),
    .A2(net257));
 sg13g2_a221oi_1 _13519_ (.B2(net371),
    .C1(net288),
    .B1(_05708_),
    .A1(_05079_),
    .Y(_05709_),
    .A2(net183));
 sg13g2_and3_1 _13520_ (.X(_05710_),
    .A(net265),
    .B(_05096_),
    .C(_05212_));
 sg13g2_nor3_1 _13521_ (.A(net180),
    .B(_05709_),
    .C(_05710_),
    .Y(_05711_));
 sg13g2_nor3_1 _13522_ (.A(_05700_),
    .B(_05707_),
    .C(_05711_),
    .Y(_05712_));
 sg13g2_a21oi_1 _13523_ (.A1(_05695_),
    .A2(net60),
    .Y(_00468_),
    .B1(_05712_));
 sg13g2_nor2_1 _13524_ (.A(_05029_),
    .B(_05303_),
    .Y(_05713_));
 sg13g2_a21oi_1 _13525_ (.A1(net397),
    .A2(_05252_),
    .Y(_05714_),
    .B1(_05713_));
 sg13g2_a22oi_1 _13526_ (.Y(_05715_),
    .B1(_05199_),
    .B2(net265),
    .A2(net373),
    .A1(_04925_));
 sg13g2_o21ai_1 _13527_ (.B1(_05715_),
    .Y(_05716_),
    .A1(net163),
    .A2(_05714_));
 sg13g2_nor3_1 _13528_ (.A(net389),
    .B(net392),
    .C(_04836_),
    .Y(_05717_));
 sg13g2_nor3_1 _13529_ (.A(_05568_),
    .B(_05437_),
    .C(_05717_),
    .Y(_05718_));
 sg13g2_o21ai_1 _13530_ (.B1(_05412_),
    .Y(_05719_),
    .A1(net192),
    .A2(_05718_));
 sg13g2_a21oi_1 _13531_ (.A1(net165),
    .A2(_05716_),
    .Y(_05720_),
    .B1(_05719_));
 sg13g2_mux2_1 _13532_ (.A0(\clock_inst.sec_c[14] ),
    .A1(_05720_),
    .S(net57),
    .X(_00469_));
 sg13g2_o21ai_1 _13533_ (.B1(_05032_),
    .Y(_05721_),
    .A1(net379),
    .A2(_04836_));
 sg13g2_o21ai_1 _13534_ (.B1(_05102_),
    .Y(_05722_),
    .A1(_05034_),
    .A2(_05432_));
 sg13g2_a21oi_1 _13535_ (.A1(_05721_),
    .A2(_05722_),
    .Y(_05723_),
    .B1(net170));
 sg13g2_o21ai_1 _13536_ (.B1(net396),
    .Y(_05724_),
    .A1(net375),
    .A2(_05027_));
 sg13g2_nand2_1 _13537_ (.Y(_05725_),
    .A(_05251_),
    .B(_05724_));
 sg13g2_a21oi_1 _13538_ (.A1(_05124_),
    .A2(_05725_),
    .Y(_05726_),
    .B1(_05146_));
 sg13g2_nor2_1 _13539_ (.A(net187),
    .B(_04946_),
    .Y(_05727_));
 sg13g2_nor4_1 _13540_ (.A(net191),
    .B(_05723_),
    .C(_05726_),
    .D(_05727_),
    .Y(_05728_));
 sg13g2_a21o_1 _13541_ (.A2(net123),
    .A1(\clock_inst.sec_c[15] ),
    .B1(_05728_),
    .X(_00470_));
 sg13g2_inv_1 _13542_ (.Y(_05729_),
    .A(\clock_inst.sec_c[16] ));
 sg13g2_and2_1 _13543_ (.A(net61),
    .B(_05119_),
    .X(_05730_));
 sg13g2_buf_1 _13544_ (.A(_05730_),
    .X(_05731_));
 sg13g2_o21ai_1 _13545_ (.B1(_05017_),
    .Y(_05732_),
    .A1(net247),
    .A2(_05070_));
 sg13g2_nor2b_1 _13546_ (.A(_05192_),
    .B_N(_05607_),
    .Y(_05733_));
 sg13g2_a21oi_1 _13547_ (.A1(net247),
    .A2(net252),
    .Y(_05734_),
    .B1(_05733_));
 sg13g2_a21oi_1 _13548_ (.A1(_05051_),
    .A2(_05734_),
    .Y(_05735_),
    .B1(net179));
 sg13g2_a221oi_1 _13549_ (.B2(_05021_),
    .C1(_05735_),
    .B1(_05732_),
    .A1(net173),
    .Y(_05736_),
    .A2(_05160_));
 sg13g2_a22oi_1 _13550_ (.Y(_00471_),
    .B1(_05731_),
    .B2(_05736_),
    .A2(_05319_),
    .A1(_05729_));
 sg13g2_inv_1 _13551_ (.Y(_05737_),
    .A(\clock_inst.sec_c[17] ));
 sg13g2_a21oi_1 _13552_ (.A1(net282),
    .A2(_04925_),
    .Y(_05738_),
    .B1(net280));
 sg13g2_nor2_1 _13553_ (.A(net513),
    .B(_05738_),
    .Y(_05739_));
 sg13g2_nor2_1 _13554_ (.A(net464),
    .B(_05083_),
    .Y(_05740_));
 sg13g2_nor2_1 _13555_ (.A(net115),
    .B(net257),
    .Y(_05741_));
 sg13g2_o21ai_1 _13556_ (.B1(net165),
    .Y(_05742_),
    .A1(_05740_),
    .A2(_05741_));
 sg13g2_a22oi_1 _13557_ (.Y(_00472_),
    .B1(_05739_),
    .B2(_05742_),
    .A2(net59),
    .A1(_05737_));
 sg13g2_inv_1 _13558_ (.Y(_05743_),
    .A(\clock_inst.sec_c[19] ));
 sg13g2_o21ai_1 _13559_ (.B1(net254),
    .Y(_05744_),
    .A1(_04979_),
    .A2(_05595_));
 sg13g2_nor2_1 _13560_ (.A(_04902_),
    .B(net169),
    .Y(_05745_));
 sg13g2_a221oi_1 _13561_ (.B2(net247),
    .C1(net513),
    .B1(_05745_),
    .A1(_05023_),
    .Y(_05746_),
    .A2(_05744_));
 sg13g2_a21oi_1 _13562_ (.A1(net278),
    .A2(net376),
    .Y(_05747_),
    .B1(net166));
 sg13g2_nand2_1 _13563_ (.Y(_05748_),
    .A(net468),
    .B(net467));
 sg13g2_a221oi_1 _13564_ (.B2(net164),
    .C1(net255),
    .B1(_05748_),
    .A1(net173),
    .Y(_05749_),
    .A2(_05295_));
 sg13g2_a21oi_1 _13565_ (.A1(net176),
    .A2(_05747_),
    .Y(_05750_),
    .B1(_05749_));
 sg13g2_nor2_1 _13566_ (.A(_05272_),
    .B(_05289_),
    .Y(_05751_));
 sg13g2_nand3_1 _13567_ (.B(net293),
    .C(_04863_),
    .A(net272),
    .Y(_05752_));
 sg13g2_o21ai_1 _13568_ (.B1(_05752_),
    .Y(_05753_),
    .A1(net184),
    .A2(_05751_));
 sg13g2_a21oi_1 _13569_ (.A1(net58),
    .A2(_05750_),
    .Y(_05754_),
    .B1(_05753_));
 sg13g2_a22oi_1 _13570_ (.Y(_00473_),
    .B1(_05746_),
    .B2(_05754_),
    .A2(net59),
    .A1(_05743_));
 sg13g2_inv_1 _13571_ (.Y(_05755_),
    .A(\clock_inst.sec_c[1] ));
 sg13g2_a21oi_1 _13572_ (.A1(net393),
    .A2(_05103_),
    .Y(_05756_),
    .B1(net470));
 sg13g2_a21oi_1 _13573_ (.A1(_04977_),
    .A2(_05151_),
    .Y(_05757_),
    .B1(net279));
 sg13g2_o21ai_1 _13574_ (.B1(net164),
    .Y(_05758_),
    .A1(_05756_),
    .A2(_05757_));
 sg13g2_a21o_1 _13575_ (.A2(_05166_),
    .A1(_04859_),
    .B1(_04840_),
    .X(_05759_));
 sg13g2_nand2_1 _13576_ (.Y(_05760_),
    .A(_05758_),
    .B(_05759_));
 sg13g2_nor2_1 _13577_ (.A(_04898_),
    .B(net461),
    .Y(_05761_));
 sg13g2_o21ai_1 _13578_ (.B1(net378),
    .Y(_05762_),
    .A1(net403),
    .A2(_04892_));
 sg13g2_nand2b_1 _13579_ (.Y(_05763_),
    .B(_05762_),
    .A_N(_05756_));
 sg13g2_a22oi_1 _13580_ (.Y(_05764_),
    .B1(_05763_),
    .B2(net178),
    .A2(_05761_),
    .A1(net167));
 sg13g2_nand2_1 _13581_ (.Y(_05765_),
    .A(net181),
    .B(_05764_));
 sg13g2_o21ai_1 _13582_ (.B1(_05765_),
    .Y(_05766_),
    .A1(net185),
    .A2(_05760_));
 sg13g2_a22oi_1 _13583_ (.Y(_00474_),
    .B1(net27),
    .B2(_05766_),
    .A2(net59),
    .A1(_05755_));
 sg13g2_inv_1 _13584_ (.Y(_05767_),
    .A(\clock_inst.sec_c[20] ));
 sg13g2_buf_1 _13585_ (.A(net122),
    .X(_05768_));
 sg13g2_a21oi_1 _13586_ (.A1(net456),
    .A2(net261),
    .Y(_05769_),
    .B1(net270));
 sg13g2_o21ai_1 _13587_ (.B1(_05147_),
    .Y(_05770_),
    .A1(net255),
    .A2(_05245_));
 sg13g2_o21ai_1 _13588_ (.B1(net118),
    .Y(_05771_),
    .A1(_05769_),
    .A2(_05770_));
 sg13g2_a21oi_1 _13589_ (.A1(net264),
    .A2(net167),
    .Y(_05772_),
    .B1(_05182_));
 sg13g2_nor2_1 _13590_ (.A(net178),
    .B(_05772_),
    .Y(_05773_));
 sg13g2_a21oi_1 _13591_ (.A1(_05415_),
    .A2(_05634_),
    .Y(_05774_),
    .B1(_05773_));
 sg13g2_nor2_1 _13592_ (.A(net255),
    .B(_05581_),
    .Y(_05775_));
 sg13g2_o21ai_1 _13593_ (.B1(net181),
    .Y(_05776_),
    .A1(_05058_),
    .A2(_05775_));
 sg13g2_nand3_1 _13594_ (.B(_05774_),
    .C(_05776_),
    .A(_05771_),
    .Y(_05777_));
 sg13g2_a22oi_1 _13595_ (.Y(_00475_),
    .B1(_05746_),
    .B2(_05777_),
    .A2(net56),
    .A1(_05767_));
 sg13g2_a21oi_1 _13596_ (.A1(_04971_),
    .A2(_05208_),
    .Y(_05778_),
    .B1(net281));
 sg13g2_nor4_1 _13597_ (.A(net382),
    .B(_04847_),
    .C(_04866_),
    .D(net172),
    .Y(_05779_));
 sg13g2_o21ai_1 _13598_ (.B1(net255),
    .Y(_05780_),
    .A1(_05778_),
    .A2(_05779_));
 sg13g2_o21ai_1 _13599_ (.B1(_05780_),
    .Y(_05781_),
    .A1(_04983_),
    .A2(_04964_));
 sg13g2_o21ai_1 _13600_ (.B1(net390),
    .Y(_05782_),
    .A1(net395),
    .A2(_05059_));
 sg13g2_o21ai_1 _13601_ (.B1(_05782_),
    .Y(_05783_),
    .A1(net247),
    .A2(_05635_));
 sg13g2_a21o_1 _13602_ (.A2(_05271_),
    .A1(net290),
    .B1(net266),
    .X(_05784_));
 sg13g2_a22oi_1 _13603_ (.Y(_05785_),
    .B1(_05784_),
    .B2(net272),
    .A2(_05783_),
    .A1(net270));
 sg13g2_nor2_1 _13604_ (.A(net171),
    .B(_05785_),
    .Y(_05786_));
 sg13g2_a21oi_1 _13605_ (.A1(net171),
    .A2(_05781_),
    .Y(_05787_),
    .B1(_05786_));
 sg13g2_nand2_1 _13606_ (.Y(_05788_),
    .A(\clock_inst.sec_c[21] ),
    .B(net114));
 sg13g2_o21ai_1 _13607_ (.B1(_05788_),
    .Y(_00476_),
    .A1(net121),
    .A2(_05787_));
 sg13g2_o21ai_1 _13608_ (.B1(_05131_),
    .Y(_05789_),
    .A1(_04844_),
    .A2(_04852_));
 sg13g2_a21oi_1 _13609_ (.A1(_04942_),
    .A2(_05455_),
    .Y(_05790_),
    .B1(net367));
 sg13g2_nor2_1 _13610_ (.A(_05195_),
    .B(_05790_),
    .Y(_05791_));
 sg13g2_a22oi_1 _13611_ (.Y(_05792_),
    .B1(_05791_),
    .B2(net181),
    .A2(_05372_),
    .A1(_05160_));
 sg13g2_a21oi_1 _13612_ (.A1(net189),
    .A2(_05789_),
    .Y(_05793_),
    .B1(_05792_));
 sg13g2_nand2_1 _13613_ (.Y(_05794_),
    .A(\clock_inst.sec_c[22] ),
    .B(net114));
 sg13g2_o21ai_1 _13614_ (.B1(_05794_),
    .Y(_00477_),
    .A1(net22),
    .A2(_05793_));
 sg13g2_o21ai_1 _13615_ (.B1(_04964_),
    .Y(_05795_),
    .A1(_05064_),
    .A2(_05070_));
 sg13g2_o21ai_1 _13616_ (.B1(net268),
    .Y(_05796_),
    .A1(net385),
    .A2(_04927_));
 sg13g2_nand3_1 _13617_ (.B(net247),
    .C(_05329_),
    .A(net254),
    .Y(_05797_));
 sg13g2_nand3_1 _13618_ (.B(_05796_),
    .C(_05797_),
    .A(net288),
    .Y(_05798_));
 sg13g2_nor2_1 _13619_ (.A(net398),
    .B(_05633_),
    .Y(_05799_));
 sg13g2_o21ai_1 _13620_ (.B1(_04994_),
    .Y(_05800_),
    .A1(_04969_),
    .A2(_05270_));
 sg13g2_o21ai_1 _13621_ (.B1(net263),
    .Y(_05801_),
    .A1(_05799_),
    .A2(_05800_));
 sg13g2_nand3_1 _13622_ (.B(_05106_),
    .C(_05801_),
    .A(net117),
    .Y(_05802_));
 sg13g2_a221oi_1 _13623_ (.B2(_05802_),
    .C1(_05005_),
    .B1(_05798_),
    .A1(net179),
    .Y(_05803_),
    .A2(_05795_));
 sg13g2_a21oi_1 _13624_ (.A1(\clock_inst.sec_c[23] ),
    .A2(net119),
    .Y(_05804_),
    .B1(_05803_));
 sg13g2_inv_1 _13625_ (.Y(_00478_),
    .A(_05804_));
 sg13g2_o21ai_1 _13626_ (.B1(net259),
    .Y(_05805_),
    .A1(net291),
    .A2(_05205_));
 sg13g2_a21o_1 _13627_ (.A2(_05805_),
    .A1(_05187_),
    .B1(net275),
    .X(_05806_));
 sg13g2_o21ai_1 _13628_ (.B1(net254),
    .Y(_05807_),
    .A1(net279),
    .A2(net401));
 sg13g2_a221oi_1 _13629_ (.B2(_05807_),
    .C1(net249),
    .B1(net177),
    .A1(_05231_),
    .Y(_05808_),
    .A2(net166));
 sg13g2_a21o_1 _13630_ (.A2(_05068_),
    .A1(_04848_),
    .B1(_05439_),
    .X(_05809_));
 sg13g2_nor2_1 _13631_ (.A(net384),
    .B(_05432_),
    .Y(_05810_));
 sg13g2_o21ai_1 _13632_ (.B1(net374),
    .Y(_05811_),
    .A1(_04836_),
    .A2(_05810_));
 sg13g2_a21oi_1 _13633_ (.A1(_05455_),
    .A2(_05811_),
    .Y(_05812_),
    .B1(net190));
 sg13g2_a21oi_1 _13634_ (.A1(_05320_),
    .A2(_05809_),
    .Y(_05813_),
    .B1(_05812_));
 sg13g2_a22oi_1 _13635_ (.Y(_05814_),
    .B1(_05813_),
    .B2(_04953_),
    .A2(_05808_),
    .A1(_05806_));
 sg13g2_mux2_1 _13636_ (.A0(\clock_inst.sec_c[24] ),
    .A1(_05814_),
    .S(net57),
    .X(_00479_));
 sg13g2_inv_1 _13637_ (.Y(_05815_),
    .A(\clock_inst.sec_c[25] ));
 sg13g2_a21oi_1 _13638_ (.A1(net275),
    .A2(_05270_),
    .Y(_05816_),
    .B1(net255));
 sg13g2_a21oi_1 _13639_ (.A1(net371),
    .A2(_04896_),
    .Y(_05817_),
    .B1(net164));
 sg13g2_nor3_1 _13640_ (.A(net376),
    .B(_05816_),
    .C(_05817_),
    .Y(_05818_));
 sg13g2_a21oi_1 _13641_ (.A1(net367),
    .A2(_05192_),
    .Y(_05819_),
    .B1(net374));
 sg13g2_nor2_1 _13642_ (.A(net282),
    .B(_05819_),
    .Y(_05820_));
 sg13g2_nor4_1 _13643_ (.A(net58),
    .B(net256),
    .C(_05100_),
    .D(_05820_),
    .Y(_05821_));
 sg13g2_a21oi_1 _13644_ (.A1(net58),
    .A2(_05818_),
    .Y(_05822_),
    .B1(_05821_));
 sg13g2_a22oi_1 _13645_ (.Y(_00480_),
    .B1(_05244_),
    .B2(_05822_),
    .A2(net56),
    .A1(_05815_));
 sg13g2_inv_1 _13646_ (.Y(_05823_),
    .A(\clock_inst.sec_c[26] ));
 sg13g2_nor2_1 _13647_ (.A(_04866_),
    .B(_04989_),
    .Y(_05824_));
 sg13g2_a22oi_1 _13648_ (.Y(_05825_),
    .B1(_05824_),
    .B2(_05022_),
    .A2(_05236_),
    .A1(_04871_));
 sg13g2_nand2_1 _13649_ (.Y(_05826_),
    .A(net373),
    .B(_05253_));
 sg13g2_o21ai_1 _13650_ (.B1(_05826_),
    .Y(_05827_),
    .A1(_04987_),
    .A2(_05825_));
 sg13g2_nor2_1 _13651_ (.A(_05160_),
    .B(net376),
    .Y(_05828_));
 sg13g2_o21ai_1 _13652_ (.B1(net260),
    .Y(_05829_),
    .A1(_05043_),
    .A2(_05272_));
 sg13g2_a221oi_1 _13653_ (.B2(_05829_),
    .C1(net22),
    .B1(_05828_),
    .A1(_05327_),
    .Y(_05830_),
    .A2(_05827_));
 sg13g2_a21oi_1 _13654_ (.A1(_05823_),
    .A2(net60),
    .Y(_00481_),
    .B1(_05830_));
 sg13g2_nand2_1 _13655_ (.Y(_05831_),
    .A(net375),
    .B(net248));
 sg13g2_o21ai_1 _13656_ (.B1(_05831_),
    .Y(_05832_),
    .A1(_05305_),
    .A2(_05252_));
 sg13g2_a22oi_1 _13657_ (.Y(_05833_),
    .B1(_05832_),
    .B2(_05298_),
    .A2(_04959_),
    .A1(_04876_));
 sg13g2_o21ai_1 _13658_ (.B1(_05165_),
    .Y(_05834_),
    .A1(_05100_),
    .A2(net252));
 sg13g2_o21ai_1 _13659_ (.B1(_05079_),
    .Y(_05835_),
    .A1(net379),
    .A2(_05094_));
 sg13g2_and2_1 _13660_ (.A(_05834_),
    .B(_05835_),
    .X(_05836_));
 sg13g2_o21ai_1 _13661_ (.B1(_05836_),
    .Y(_05837_),
    .A1(net260),
    .A2(_05833_));
 sg13g2_a22oi_1 _13662_ (.Y(_05838_),
    .B1(net27),
    .B2(_05837_),
    .A2(_04938_),
    .A1(\clock_inst.sec_c[27] ));
 sg13g2_inv_1 _13663_ (.Y(_00482_),
    .A(_05838_));
 sg13g2_nand3_1 _13664_ (.B(net261),
    .C(_05404_),
    .A(net367),
    .Y(_05839_));
 sg13g2_nand3b_1 _13665_ (.B(_05411_),
    .C(_05839_),
    .Y(_05840_),
    .A_N(_05128_));
 sg13g2_o21ai_1 _13666_ (.B1(net261),
    .Y(_05841_),
    .A1(net175),
    .A2(_05384_));
 sg13g2_nor2_1 _13667_ (.A(_04902_),
    .B(_05252_),
    .Y(_05842_));
 sg13g2_a21o_1 _13668_ (.A2(_05841_),
    .A1(_05475_),
    .B1(_05842_),
    .X(_05843_));
 sg13g2_o21ai_1 _13669_ (.B1(_05529_),
    .Y(_05844_),
    .A1(_05349_),
    .A2(_05621_));
 sg13g2_a221oi_1 _13670_ (.B2(net456),
    .C1(_05844_),
    .B1(_05843_),
    .A1(net118),
    .Y(_05845_),
    .A2(_05840_));
 sg13g2_nand2_1 _13671_ (.Y(_05846_),
    .A(\clock_inst.sec_c[28] ),
    .B(net114));
 sg13g2_o21ai_1 _13672_ (.B1(_05846_),
    .Y(_00483_),
    .A1(net121),
    .A2(_05845_));
 sg13g2_a21oi_1 _13673_ (.A1(net186),
    .A2(_05346_),
    .Y(_05847_),
    .B1(net275));
 sg13g2_a21oi_1 _13674_ (.A1(_05212_),
    .A2(_05208_),
    .Y(_05848_),
    .B1(net270));
 sg13g2_a221oi_1 _13675_ (.B2(_05375_),
    .C1(_05848_),
    .B1(_05824_),
    .A1(net178),
    .Y(_05849_),
    .A2(net183));
 sg13g2_o21ai_1 _13676_ (.B1(_05849_),
    .Y(_05850_),
    .A1(net58),
    .A2(_05847_));
 sg13g2_nand2_1 _13677_ (.Y(_05851_),
    .A(\clock_inst.sec_c[29] ),
    .B(net114));
 sg13g2_o21ai_1 _13678_ (.B1(_05851_),
    .Y(_00484_),
    .A1(net121),
    .A2(_05850_));
 sg13g2_inv_1 _13679_ (.Y(_05852_),
    .A(\clock_inst.sec_c[2] ));
 sg13g2_a22oi_1 _13680_ (.Y(_05853_),
    .B1(_05252_),
    .B2(net267),
    .A2(_05158_),
    .A1(_04876_));
 sg13g2_nand3_1 _13681_ (.B(_05371_),
    .C(_05460_),
    .A(_05321_),
    .Y(_05854_));
 sg13g2_o21ai_1 _13682_ (.B1(_05854_),
    .Y(_05855_),
    .A1(_04955_),
    .A2(_05853_));
 sg13g2_a21oi_1 _13683_ (.A1(_05256_),
    .A2(_05855_),
    .Y(_05856_),
    .B1(_05005_));
 sg13g2_a22oi_1 _13684_ (.Y(_05857_),
    .B1(_05460_),
    .B2(_05025_),
    .A2(_05158_),
    .A1(net251));
 sg13g2_nand2_1 _13685_ (.Y(_05858_),
    .A(_05371_),
    .B(_05247_));
 sg13g2_o21ai_1 _13686_ (.B1(_05858_),
    .Y(_05859_),
    .A1(_05145_),
    .A2(_05857_));
 sg13g2_a22oi_1 _13687_ (.Y(_05860_),
    .B1(_05081_),
    .B2(_05100_),
    .A2(_04993_),
    .A1(net378));
 sg13g2_or2_1 _13688_ (.X(_05861_),
    .B(_05860_),
    .A(net269));
 sg13g2_nand3_1 _13689_ (.B(_05368_),
    .C(_05861_),
    .A(_05826_),
    .Y(_05862_));
 sg13g2_a22oi_1 _13690_ (.Y(_05863_),
    .B1(_05862_),
    .B2(net185),
    .A2(_05859_),
    .A1(_05136_));
 sg13g2_a22oi_1 _13691_ (.Y(_00485_),
    .B1(_05856_),
    .B2(_05863_),
    .A2(_05768_),
    .A1(_05852_));
 sg13g2_buf_1 _13692_ (.A(\clock_inst.sec_c[30] ),
    .X(_05864_));
 sg13g2_o21ai_1 _13693_ (.B1(net171),
    .Y(_05865_),
    .A1(_05039_),
    .A2(_05701_));
 sg13g2_a21oi_1 _13694_ (.A1(_05696_),
    .A2(_05865_),
    .Y(_05866_),
    .B1(net122));
 sg13g2_a21o_1 _13695_ (.A2(net123),
    .A1(_05864_),
    .B1(_05866_),
    .X(_00486_));
 sg13g2_inv_1 _13696_ (.Y(_05867_),
    .A(\clock_inst.sec_c[36] ));
 sg13g2_a21oi_1 _13697_ (.A1(_05305_),
    .A2(_05402_),
    .Y(_05868_),
    .B1(_05126_));
 sg13g2_nand2_1 _13698_ (.Y(_05869_),
    .A(_04881_),
    .B(net287));
 sg13g2_o21ai_1 _13699_ (.B1(_04957_),
    .Y(_05870_),
    .A1(_05229_),
    .A2(_05334_));
 sg13g2_a21o_1 _13700_ (.A2(_05870_),
    .A1(_05869_),
    .B1(net265),
    .X(_05871_));
 sg13g2_o21ai_1 _13701_ (.B1(_05871_),
    .Y(_05872_),
    .A1(net170),
    .A2(_05868_));
 sg13g2_nand2_1 _13702_ (.Y(_05873_),
    .A(_04956_),
    .B(net383));
 sg13g2_o21ai_1 _13703_ (.B1(_05748_),
    .Y(_05874_),
    .A1(_05873_),
    .A2(_05158_));
 sg13g2_nand3_1 _13704_ (.B(_04959_),
    .C(_05874_),
    .A(_05214_),
    .Y(_05875_));
 sg13g2_o21ai_1 _13705_ (.B1(net257),
    .Y(_05876_),
    .A1(_04836_),
    .A2(_05150_));
 sg13g2_nand3_1 _13706_ (.B(_05875_),
    .C(_05876_),
    .A(_05087_),
    .Y(_05877_));
 sg13g2_o21ai_1 _13707_ (.B1(_05877_),
    .Y(_05878_),
    .A1(_04953_),
    .A2(_05872_));
 sg13g2_a22oi_1 _13708_ (.Y(_00487_),
    .B1(_05731_),
    .B2(_05878_),
    .A2(net56),
    .A1(_05867_));
 sg13g2_inv_1 _13709_ (.Y(_05879_),
    .A(\clock_inst.sec_c[37] ));
 sg13g2_a22oi_1 _13710_ (.Y(_05880_),
    .B1(_05180_),
    .B2(net283),
    .A2(net380),
    .A1(net287));
 sg13g2_o21ai_1 _13711_ (.B1(_04876_),
    .Y(_05881_),
    .A1(_05023_),
    .A2(_05243_));
 sg13g2_o21ai_1 _13712_ (.B1(_05881_),
    .Y(_05882_),
    .A1(_05118_),
    .A2(_05880_));
 sg13g2_nand2_1 _13713_ (.Y(_05883_),
    .A(net170),
    .B(_05882_));
 sg13g2_a21oi_1 _13714_ (.A1(_05032_),
    .A2(_05260_),
    .Y(_05884_),
    .B1(net262));
 sg13g2_nand2_1 _13715_ (.Y(_05885_),
    .A(_05272_),
    .B(_05437_));
 sg13g2_o21ai_1 _13716_ (.B1(_05885_),
    .Y(_05886_),
    .A1(_05673_),
    .A2(_05884_));
 sg13g2_xnor2_1 _13717_ (.Y(_05887_),
    .A(_04961_),
    .B(net267));
 sg13g2_o21ai_1 _13718_ (.B1(_05055_),
    .Y(_05888_),
    .A1(_05515_),
    .A2(_05887_));
 sg13g2_a221oi_1 _13719_ (.B2(_05250_),
    .C1(_05888_),
    .B1(_05886_),
    .A1(_05034_),
    .Y(_05889_),
    .A2(_05334_));
 sg13g2_a22oi_1 _13720_ (.Y(_00488_),
    .B1(_05883_),
    .B2(_05889_),
    .A2(net56),
    .A1(_05879_));
 sg13g2_inv_1 _13721_ (.Y(_05890_),
    .A(\clock_inst.sec_c[38] ));
 sg13g2_a22oi_1 _13722_ (.Y(_05891_),
    .B1(_05253_),
    .B2(net373),
    .A2(_05371_),
    .A1(_04830_));
 sg13g2_o21ai_1 _13723_ (.B1(_05475_),
    .Y(_05892_),
    .A1(_04836_),
    .A2(net403));
 sg13g2_o21ai_1 _13724_ (.B1(_05892_),
    .Y(_05893_),
    .A1(net171),
    .A2(_05891_));
 sg13g2_a22oi_1 _13725_ (.Y(_05894_),
    .B1(_05104_),
    .B2(net378),
    .A2(net273),
    .A1(_04876_));
 sg13g2_inv_1 _13726_ (.Y(_05895_),
    .A(_05894_));
 sg13g2_o21ai_1 _13727_ (.B1(net274),
    .Y(_05896_),
    .A1(_04973_),
    .A2(_04894_));
 sg13g2_a22oi_1 _13728_ (.Y(_05897_),
    .B1(_05896_),
    .B2(_05079_),
    .A2(_05895_),
    .A1(net178));
 sg13g2_nand2_1 _13729_ (.Y(_05898_),
    .A(_05093_),
    .B(_05897_));
 sg13g2_o21ai_1 _13730_ (.B1(_05898_),
    .Y(_05899_),
    .A1(net185),
    .A2(_05893_));
 sg13g2_a22oi_1 _13731_ (.Y(_00489_),
    .B1(_05856_),
    .B2(_05899_),
    .A2(_05768_),
    .A1(_05890_));
 sg13g2_a22oi_1 _13732_ (.Y(_05900_),
    .B1(_05411_),
    .B2(_04852_),
    .A2(_05033_),
    .A1(net287));
 sg13g2_nand2_1 _13733_ (.Y(_05901_),
    .A(_05073_),
    .B(net274));
 sg13g2_a221oi_1 _13734_ (.B2(_05901_),
    .C1(net253),
    .B1(_05457_),
    .A1(net379),
    .Y(_05902_),
    .A2(_05873_));
 sg13g2_a21oi_1 _13735_ (.A1(net170),
    .A2(_05900_),
    .Y(_05903_),
    .B1(_05902_));
 sg13g2_o21ai_1 _13736_ (.B1(net463),
    .Y(_05904_),
    .A1(net462),
    .A2(_05192_));
 sg13g2_o21ai_1 _13737_ (.B1(net390),
    .Y(_05905_),
    .A1(net462),
    .A2(net391));
 sg13g2_nand2_1 _13738_ (.Y(_05906_),
    .A(_05904_),
    .B(_05905_));
 sg13g2_nand2_1 _13739_ (.Y(_05907_),
    .A(_04940_),
    .B(_05033_));
 sg13g2_o21ai_1 _13740_ (.B1(_05907_),
    .Y(_05908_),
    .A1(_05371_),
    .A2(_05258_));
 sg13g2_a22oi_1 _13741_ (.Y(_05909_),
    .B1(_05908_),
    .B2(net190),
    .A2(_05906_),
    .A1(net269));
 sg13g2_nor2_1 _13742_ (.A(net186),
    .B(_05909_),
    .Y(_05910_));
 sg13g2_a221oi_1 _13743_ (.B2(net176),
    .C1(_05910_),
    .B1(_05903_),
    .A1(net369),
    .Y(_05911_),
    .A2(_05292_));
 sg13g2_mux2_1 _13744_ (.A0(\clock_inst.sec_c[39] ),
    .A1(_05911_),
    .S(_05360_),
    .X(_00490_));
 sg13g2_o21ai_1 _13745_ (.B1(net271),
    .Y(_05912_),
    .A1(_05063_),
    .A2(_05128_));
 sg13g2_a21oi_1 _13746_ (.A1(_04847_),
    .A2(net276),
    .Y(_05913_),
    .B1(net382));
 sg13g2_o21ai_1 _13747_ (.B1(net269),
    .Y(_05914_),
    .A1(net368),
    .A2(_05913_));
 sg13g2_nand3_1 _13748_ (.B(_05912_),
    .C(_05914_),
    .A(_05106_),
    .Y(_05915_));
 sg13g2_nor2_1 _13749_ (.A(net281),
    .B(_05363_),
    .Y(_05916_));
 sg13g2_o21ai_1 _13750_ (.B1(net164),
    .Y(_05917_),
    .A1(net173),
    .A2(_05916_));
 sg13g2_nand2_1 _13751_ (.Y(_05918_),
    .A(net462),
    .B(_04856_));
 sg13g2_nand2_1 _13752_ (.Y(_05919_),
    .A(net174),
    .B(_05918_));
 sg13g2_o21ai_1 _13753_ (.B1(net169),
    .Y(_05920_),
    .A1(_04991_),
    .A2(net248));
 sg13g2_a22oi_1 _13754_ (.Y(_05921_),
    .B1(_05920_),
    .B2(net277),
    .A2(_05919_),
    .A1(_05262_));
 sg13g2_a21oi_1 _13755_ (.A1(_05917_),
    .A2(_05921_),
    .Y(_05922_),
    .B1(net192));
 sg13g2_a221oi_1 _13756_ (.B2(net182),
    .C1(_05922_),
    .B1(_05915_),
    .A1(net376),
    .Y(_05923_),
    .A2(_05269_));
 sg13g2_nand2_1 _13757_ (.Y(_05924_),
    .A(\clock_inst.sec_c[3] ),
    .B(net114));
 sg13g2_o21ai_1 _13758_ (.B1(_05924_),
    .Y(_00491_),
    .A1(net22),
    .A2(_05923_));
 sg13g2_inv_1 _13759_ (.Y(_05925_),
    .A(\clock_inst.sec_c[40] ));
 sg13g2_o21ai_1 _13760_ (.B1(_05098_),
    .Y(_05926_),
    .A1(_04878_),
    .A2(net368));
 sg13g2_nand2_1 _13761_ (.Y(_05927_),
    .A(net251),
    .B(_05926_));
 sg13g2_nand3b_1 _13762_ (.B(_04974_),
    .C(_05017_),
    .Y(_05928_),
    .A_N(_05128_));
 sg13g2_o21ai_1 _13763_ (.B1(_05748_),
    .Y(_05929_),
    .A1(net187),
    .A2(_05081_));
 sg13g2_a221oi_1 _13764_ (.B2(_04849_),
    .C1(net176),
    .B1(_05929_),
    .A1(_05927_),
    .Y(_05930_),
    .A2(_05928_));
 sg13g2_a21oi_1 _13765_ (.A1(net279),
    .A2(net177),
    .Y(_05931_),
    .B1(_05207_));
 sg13g2_o21ai_1 _13766_ (.B1(net460),
    .Y(_05932_),
    .A1(_05164_),
    .A2(_05025_));
 sg13g2_a22oi_1 _13767_ (.Y(_05933_),
    .B1(_05932_),
    .B2(net371),
    .A2(net256),
    .A1(net379));
 sg13g2_o21ai_1 _13768_ (.B1(_05933_),
    .Y(_05934_),
    .A1(net275),
    .A2(_05931_));
 sg13g2_o21ai_1 _13769_ (.B1(_05731_),
    .Y(_05935_),
    .A1(net182),
    .A2(_05934_));
 sg13g2_nor2_1 _13770_ (.A(_05930_),
    .B(_05935_),
    .Y(_05936_));
 sg13g2_a21oi_1 _13771_ (.A1(_05925_),
    .A2(_05049_),
    .Y(_00492_),
    .B1(_05936_));
 sg13g2_inv_1 _13772_ (.Y(_05937_),
    .A(\clock_inst.sec_c[41] ));
 sg13g2_o21ai_1 _13773_ (.B1(net389),
    .Y(_05938_),
    .A1(net264),
    .A2(net172));
 sg13g2_a21oi_1 _13774_ (.A1(net187),
    .A2(_05938_),
    .Y(_05939_),
    .B1(_05030_));
 sg13g2_a221oi_1 _13775_ (.B2(net117),
    .C1(_05939_),
    .B1(net166),
    .A1(net249),
    .Y(_05940_),
    .A2(_05199_));
 sg13g2_nand2_1 _13776_ (.Y(_05941_),
    .A(net268),
    .B(net274));
 sg13g2_nor2_1 _13777_ (.A(net290),
    .B(net401),
    .Y(_05942_));
 sg13g2_o21ai_1 _13778_ (.B1(net279),
    .Y(_05943_),
    .A1(net258),
    .A2(net273));
 sg13g2_a22oi_1 _13779_ (.Y(_05944_),
    .B1(_05943_),
    .B2(net186),
    .A2(_05942_),
    .A1(_05941_));
 sg13g2_a21oi_1 _13780_ (.A1(net463),
    .A2(_05748_),
    .Y(_05945_),
    .B1(net377));
 sg13g2_o21ai_1 _13781_ (.B1(net253),
    .Y(_05946_),
    .A1(_05058_),
    .A2(_05945_));
 sg13g2_nand3_1 _13782_ (.B(_04863_),
    .C(_05946_),
    .A(net272),
    .Y(_05947_));
 sg13g2_o21ai_1 _13783_ (.B1(_05947_),
    .Y(_05948_),
    .A1(net292),
    .A2(_05944_));
 sg13g2_o21ai_1 _13784_ (.B1(_05948_),
    .Y(_05949_),
    .A1(net116),
    .A2(_05940_));
 sg13g2_a21oi_1 _13785_ (.A1(_05053_),
    .A2(_05343_),
    .Y(_05950_),
    .B1(net22));
 sg13g2_a22oi_1 _13786_ (.Y(_00493_),
    .B1(_05949_),
    .B2(_05950_),
    .A2(net56),
    .A1(_05937_));
 sg13g2_o21ai_1 _13787_ (.B1(_05366_),
    .Y(_05951_),
    .A1(net281),
    .A2(_05158_));
 sg13g2_or2_1 _13788_ (.X(_05952_),
    .B(_05182_),
    .A(_05158_));
 sg13g2_a21oi_1 _13789_ (.A1(_05411_),
    .A2(_05350_),
    .Y(_05953_),
    .B1(_04830_));
 sg13g2_a221oi_1 _13790_ (.B2(net163),
    .C1(_05953_),
    .B1(_05952_),
    .A1(net283),
    .Y(_05954_),
    .A2(_05951_));
 sg13g2_o21ai_1 _13791_ (.B1(_05508_),
    .Y(_05955_),
    .A1(_05251_),
    .A2(_05704_));
 sg13g2_nand3_1 _13792_ (.B(_04982_),
    .C(net370),
    .A(net381),
    .Y(_05956_));
 sg13g2_a21oi_1 _13793_ (.A1(_05166_),
    .A2(_05956_),
    .Y(_05957_),
    .B1(net278));
 sg13g2_a221oi_1 _13794_ (.B2(net188),
    .C1(_05957_),
    .B1(_05955_),
    .A1(net380),
    .Y(_05958_),
    .A2(_05761_));
 sg13g2_o21ai_1 _13795_ (.B1(_05958_),
    .Y(_05959_),
    .A1(net165),
    .A2(_05954_));
 sg13g2_mux2_1 _13796_ (.A0(\clock_inst.sec_c[42] ),
    .A1(_05959_),
    .S(net57),
    .X(_00494_));
 sg13g2_o21ai_1 _13797_ (.B1(net286),
    .Y(_05960_),
    .A1(_04852_),
    .A2(_05305_));
 sg13g2_nand2b_1 _13798_ (.Y(_05961_),
    .B(_05960_),
    .A_N(_05229_));
 sg13g2_a21oi_1 _13799_ (.A1(net247),
    .A2(_05151_),
    .Y(_05962_),
    .B1(net278));
 sg13g2_a221oi_1 _13800_ (.B2(net283),
    .C1(_05962_),
    .B1(_05961_),
    .A1(_05083_),
    .Y(_05963_),
    .A2(_05100_));
 sg13g2_nor2_1 _13801_ (.A(_04943_),
    .B(_04902_),
    .Y(_05964_));
 sg13g2_a22oi_1 _13802_ (.Y(_05965_),
    .B1(_04970_),
    .B2(net268),
    .A2(net264),
    .A1(net386));
 sg13g2_o21ai_1 _13803_ (.B1(net259),
    .Y(_05966_),
    .A1(_05292_),
    .A2(_05460_));
 sg13g2_nand2_1 _13804_ (.Y(_05967_),
    .A(_05965_),
    .B(_05966_));
 sg13g2_a22oi_1 _13805_ (.Y(_05968_),
    .B1(_05967_),
    .B2(net181),
    .A2(_05964_),
    .A1(net461));
 sg13g2_o21ai_1 _13806_ (.B1(_05968_),
    .Y(_05969_),
    .A1(net185),
    .A2(_05963_));
 sg13g2_nand2_1 _13807_ (.Y(_05970_),
    .A(\clock_inst.sec_c[43] ),
    .B(_05559_));
 sg13g2_o21ai_1 _13808_ (.B1(_05970_),
    .Y(_00495_),
    .A1(_04950_),
    .A2(_05969_));
 sg13g2_nor2_1 _13809_ (.A(\clock_inst.sec_c[44] ),
    .B(_05360_),
    .Y(_05971_));
 sg13g2_o21ai_1 _13810_ (.B1(net377),
    .Y(_05972_),
    .A1(net459),
    .A2(net256));
 sg13g2_a21oi_1 _13811_ (.A1(_05009_),
    .A2(_05972_),
    .Y(_05973_),
    .B1(net402));
 sg13g2_a22oi_1 _13812_ (.Y(_05974_),
    .B1(_05338_),
    .B2(_05366_),
    .A2(_05180_),
    .A1(net290));
 sg13g2_nor2_1 _13813_ (.A(net277),
    .B(_05974_),
    .Y(_05975_));
 sg13g2_nor3_1 _13814_ (.A(net163),
    .B(_05973_),
    .C(_05975_),
    .Y(_05976_));
 sg13g2_xnor2_1 _13815_ (.Y(_05977_),
    .A(_04913_),
    .B(net459));
 sg13g2_nor3_1 _13816_ (.A(net404),
    .B(net262),
    .C(_05432_),
    .Y(_05978_));
 sg13g2_a21oi_1 _13817_ (.A1(net397),
    .A2(_05977_),
    .Y(_05979_),
    .B1(_05978_));
 sg13g2_a221oi_1 _13818_ (.B2(net170),
    .C1(net168),
    .B1(_05979_),
    .A1(net177),
    .Y(_05980_),
    .A2(_05403_));
 sg13g2_a21oi_1 _13819_ (.A1(_05052_),
    .A2(_05115_),
    .Y(_05981_),
    .B1(_05120_));
 sg13g2_o21ai_1 _13820_ (.B1(_05981_),
    .Y(_05982_),
    .A1(_05976_),
    .A2(_05980_));
 sg13g2_nor2b_1 _13821_ (.A(_05971_),
    .B_N(_05982_),
    .Y(_00496_));
 sg13g2_inv_1 _13822_ (.Y(_05983_),
    .A(\clock_inst.sec_c[45] ));
 sg13g2_o21ai_1 _13823_ (.B1(net247),
    .Y(_05984_),
    .A1(net173),
    .A2(_05270_));
 sg13g2_a22oi_1 _13824_ (.Y(_05985_),
    .B1(_05984_),
    .B2(net58),
    .A2(_05034_),
    .A1(net257));
 sg13g2_a22oi_1 _13825_ (.Y(_05986_),
    .B1(net289),
    .B2(_05330_),
    .A2(_04896_),
    .A1(net266));
 sg13g2_nor2_1 _13826_ (.A(net117),
    .B(_05986_),
    .Y(_05987_));
 sg13g2_o21ai_1 _13827_ (.B1(_05701_),
    .Y(_05988_),
    .A1(net280),
    .A2(net369));
 sg13g2_a21oi_1 _13828_ (.A1(net257),
    .A2(_05033_),
    .Y(_05989_),
    .B1(_04892_));
 sg13g2_a21oi_1 _13829_ (.A1(_05988_),
    .A2(_05989_),
    .Y(_05990_),
    .B1(net282));
 sg13g2_nor2_1 _13830_ (.A(_05987_),
    .B(_05990_),
    .Y(_05991_));
 sg13g2_o21ai_1 _13831_ (.B1(_05991_),
    .Y(_05992_),
    .A1(net189),
    .A2(_05985_));
 sg13g2_a22oi_1 _13832_ (.Y(_00497_),
    .B1(_05244_),
    .B2(_05992_),
    .A2(net56),
    .A1(_05983_));
 sg13g2_a21o_1 _13833_ (.A2(net266),
    .A1(_04996_),
    .B1(_05229_),
    .X(_05993_));
 sg13g2_o21ai_1 _13834_ (.B1(_05704_),
    .Y(_05994_),
    .A1(_05019_),
    .A2(net172));
 sg13g2_a21oi_1 _13835_ (.A1(net164),
    .A2(_05402_),
    .Y(_05995_),
    .B1(_05415_));
 sg13g2_a221oi_1 _13836_ (.B2(_05182_),
    .C1(_05995_),
    .B1(_05994_),
    .A1(_05020_),
    .Y(_05996_),
    .A2(_05993_));
 sg13g2_nand2_1 _13837_ (.Y(_05997_),
    .A(net461),
    .B(_05096_));
 sg13g2_o21ai_1 _13838_ (.B1(net386),
    .Y(_05998_),
    .A1(net291),
    .A2(_05323_));
 sg13g2_o21ai_1 _13839_ (.B1(_04942_),
    .Y(_05999_),
    .A1(net177),
    .A2(_05476_));
 sg13g2_nand3_1 _13840_ (.B(_05998_),
    .C(_05999_),
    .A(_05212_),
    .Y(_06000_));
 sg13g2_a22oi_1 _13841_ (.Y(_06001_),
    .B1(_06000_),
    .B2(_05118_),
    .A2(_05997_),
    .A1(_04822_));
 sg13g2_o21ai_1 _13842_ (.B1(_06001_),
    .Y(_06002_),
    .A1(net116),
    .A2(_05996_));
 sg13g2_nand2_1 _13843_ (.Y(_06003_),
    .A(\clock_inst.sec_c[46] ),
    .B(net114));
 sg13g2_o21ai_1 _13844_ (.B1(_06003_),
    .Y(_00498_),
    .A1(net123),
    .A2(_06002_));
 sg13g2_a22oi_1 _13845_ (.Y(_06004_),
    .B1(_05446_),
    .B2(_05512_),
    .A2(_05411_),
    .A1(net373));
 sg13g2_o21ai_1 _13846_ (.B1(_05225_),
    .Y(_06005_),
    .A1(net250),
    .A2(_05386_));
 sg13g2_o21ai_1 _13847_ (.B1(_06005_),
    .Y(_06006_),
    .A1(_04919_),
    .A2(_05051_));
 sg13g2_o21ai_1 _13848_ (.B1(net389),
    .Y(_06007_),
    .A1(_05165_),
    .A2(_05510_));
 sg13g2_a21oi_1 _13849_ (.A1(_04959_),
    .A2(_05366_),
    .Y(_06008_),
    .B1(net384));
 sg13g2_nor2_1 _13850_ (.A(net392),
    .B(_05635_),
    .Y(_06009_));
 sg13g2_o21ai_1 _13851_ (.B1(net385),
    .Y(_06010_),
    .A1(_06008_),
    .A2(_06009_));
 sg13g2_nand4_1 _13852_ (.B(_05017_),
    .C(_06007_),
    .A(net270),
    .Y(_06011_),
    .D(_06010_));
 sg13g2_o21ai_1 _13853_ (.B1(_06011_),
    .Y(_06012_),
    .A1(net192),
    .A2(_06006_));
 sg13g2_o21ai_1 _13854_ (.B1(_06012_),
    .Y(_06013_),
    .A1(net165),
    .A2(_06004_));
 sg13g2_mux2_1 _13855_ (.A0(\clock_inst.sec_c[47] ),
    .A1(_06013_),
    .S(net57),
    .X(_00499_));
 sg13g2_inv_1 _13856_ (.Y(_06014_),
    .A(\clock_inst.sec_c[48] ));
 sg13g2_o21ai_1 _13857_ (.B1(net186),
    .Y(_06015_),
    .A1(net190),
    .A2(_05446_));
 sg13g2_nand2_1 _13858_ (.Y(_06016_),
    .A(net254),
    .B(_06015_));
 sg13g2_a21o_1 _13859_ (.A2(net391),
    .A1(net192),
    .B1(_05275_),
    .X(_06017_));
 sg13g2_a22oi_1 _13860_ (.Y(_06018_),
    .B1(_06017_),
    .B2(_04892_),
    .A2(_06016_),
    .A1(net177));
 sg13g2_o21ai_1 _13861_ (.B1(_05036_),
    .Y(_06019_),
    .A1(net396),
    .A2(net250));
 sg13g2_a21oi_1 _13862_ (.A1(_05200_),
    .A2(_06019_),
    .Y(_06020_),
    .B1(net265));
 sg13g2_a21oi_1 _13863_ (.A1(net389),
    .A2(_05233_),
    .Y(_06021_),
    .B1(net401));
 sg13g2_o21ai_1 _13864_ (.B1(_05918_),
    .Y(_06022_),
    .A1(_05070_),
    .A2(_06021_));
 sg13g2_o21ai_1 _13865_ (.B1(net260),
    .Y(_06023_),
    .A1(_06020_),
    .A2(_06022_));
 sg13g2_nor2b_1 _13866_ (.A(_05700_),
    .B_N(_06023_),
    .Y(_06024_));
 sg13g2_a22oi_1 _13867_ (.Y(_00500_),
    .B1(_06018_),
    .B2(_06024_),
    .A2(net56),
    .A1(_06014_));
 sg13g2_o21ai_1 _13868_ (.B1(_05106_),
    .Y(_06025_),
    .A1(net254),
    .A2(_05289_));
 sg13g2_a21oi_1 _13869_ (.A1(_05233_),
    .A2(_05607_),
    .Y(_06026_),
    .B1(_05740_));
 sg13g2_a21oi_1 _13870_ (.A1(_05212_),
    .A2(_06026_),
    .Y(_06027_),
    .B1(net115));
 sg13g2_a21oi_1 _13871_ (.A1(net117),
    .A2(_06025_),
    .Y(_06028_),
    .B1(_06027_));
 sg13g2_a21oi_1 _13872_ (.A1(net470),
    .A2(net388),
    .Y(_06029_),
    .B1(net273));
 sg13g2_o21ai_1 _13873_ (.B1(_05492_),
    .Y(_06030_),
    .A1(net253),
    .A2(_06029_));
 sg13g2_a22oi_1 _13874_ (.Y(_06031_),
    .B1(_05289_),
    .B2(_05522_),
    .A2(net369),
    .A1(net264));
 sg13g2_nor2_1 _13875_ (.A(net277),
    .B(_06031_),
    .Y(_06032_));
 sg13g2_a21oi_1 _13876_ (.A1(net163),
    .A2(_06030_),
    .Y(_06033_),
    .B1(_06032_));
 sg13g2_o21ai_1 _13877_ (.B1(_06033_),
    .Y(_06034_),
    .A1(net163),
    .A2(_06028_));
 sg13g2_a22oi_1 _13878_ (.Y(_06035_),
    .B1(net61),
    .B2(_06034_),
    .A2(net122),
    .A1(\clock_inst.sec_c[49] ));
 sg13g2_inv_1 _13879_ (.Y(_00501_),
    .A(_06035_));
 sg13g2_o21ai_1 _13880_ (.B1(net263),
    .Y(_06036_),
    .A1(net258),
    .A2(net177));
 sg13g2_nand3_1 _13881_ (.B(_05211_),
    .C(_06036_),
    .A(net276),
    .Y(_06037_));
 sg13g2_o21ai_1 _13882_ (.B1(_05193_),
    .Y(_06038_),
    .A1(_04921_),
    .A2(net187));
 sg13g2_a22oi_1 _13883_ (.Y(_06039_),
    .B1(net174),
    .B2(_05182_),
    .A2(net166),
    .A1(net271));
 sg13g2_nor2_1 _13884_ (.A(net466),
    .B(_05168_),
    .Y(_06040_));
 sg13g2_o21ai_1 _13885_ (.B1(_05233_),
    .Y(_06041_),
    .A1(net399),
    .A2(_04815_));
 sg13g2_inv_1 _13886_ (.Y(_06042_),
    .A(_06041_));
 sg13g2_a22oi_1 _13887_ (.Y(_06043_),
    .B1(_06042_),
    .B2(net381),
    .A2(_06040_),
    .A1(_05009_));
 sg13g2_a21oi_1 _13888_ (.A1(_05151_),
    .A2(_05599_),
    .Y(_06044_),
    .B1(_04991_));
 sg13g2_nor3_1 _13889_ (.A(net265),
    .B(_06043_),
    .C(_06044_),
    .Y(_06045_));
 sg13g2_a21oi_1 _13890_ (.A1(net292),
    .A2(_06039_),
    .Y(_06046_),
    .B1(_06045_));
 sg13g2_a221oi_1 _13891_ (.B2(net182),
    .C1(_06046_),
    .B1(_06038_),
    .A1(net163),
    .Y(_06047_),
    .A2(_06037_));
 sg13g2_nand2_1 _13892_ (.Y(_06048_),
    .A(\clock_inst.sec_c[4] ),
    .B(net119));
 sg13g2_o21ai_1 _13893_ (.B1(_06048_),
    .Y(_00502_),
    .A1(net123),
    .A2(_06047_));
 sg13g2_inv_1 _13894_ (.Y(_06049_),
    .A(\clock_inst.sec_c[50] ));
 sg13g2_a21oi_1 _13895_ (.A1(net284),
    .A2(_04946_),
    .Y(_06050_),
    .B1(_05008_));
 sg13g2_nand2_1 _13896_ (.Y(_06051_),
    .A(net373),
    .B(net187));
 sg13g2_o21ai_1 _13897_ (.B1(_06051_),
    .Y(_06052_),
    .A1(_05616_),
    .A2(_06050_));
 sg13g2_o21ai_1 _13898_ (.B1(net284),
    .Y(_06053_),
    .A1(_05064_),
    .A2(_05070_));
 sg13g2_a21oi_1 _13899_ (.A1(_05187_),
    .A2(_05515_),
    .Y(_06054_),
    .B1(_04831_));
 sg13g2_a221oi_1 _13900_ (.B2(_05327_),
    .C1(_06054_),
    .B1(_06053_),
    .A1(_05301_),
    .Y(_06055_),
    .A2(_06052_));
 sg13g2_a22oi_1 _13901_ (.Y(_00503_),
    .B1(_05731_),
    .B2(_06055_),
    .A2(net56),
    .A1(_06049_));
 sg13g2_a21oi_1 _13902_ (.A1(_05307_),
    .A2(_05411_),
    .Y(_06056_),
    .B1(net170));
 sg13g2_nor3_1 _13903_ (.A(_05726_),
    .B(_05727_),
    .C(_06056_),
    .Y(_06057_));
 sg13g2_nand2_1 _13904_ (.Y(_06058_),
    .A(\clock_inst.sec_c[51] ),
    .B(net119));
 sg13g2_o21ai_1 _13905_ (.B1(_06058_),
    .Y(_00504_),
    .A1(net123),
    .A2(_06057_));
 sg13g2_a21oi_1 _13906_ (.A1(net255),
    .A2(_04991_),
    .Y(_06059_),
    .B1(_05083_));
 sg13g2_o21ai_1 _13907_ (.B1(net292),
    .Y(_06060_),
    .A1(_05510_),
    .A2(_06059_));
 sg13g2_a22oi_1 _13908_ (.Y(_06061_),
    .B1(net369),
    .B2(net266),
    .A2(net257),
    .A1(net389));
 sg13g2_nor2_1 _13909_ (.A(net294),
    .B(_06061_),
    .Y(_06062_));
 sg13g2_a21oi_1 _13910_ (.A1(net254),
    .A2(_05106_),
    .Y(_06063_),
    .B1(net265));
 sg13g2_nor3_1 _13911_ (.A(_05229_),
    .B(_06062_),
    .C(_06063_),
    .Y(_06064_));
 sg13g2_a21oi_1 _13912_ (.A1(_06060_),
    .A2(_06064_),
    .Y(_06065_),
    .B1(_05005_));
 sg13g2_a21o_1 _13913_ (.A2(_04937_),
    .A1(\clock_inst.sec_c[52] ),
    .B1(_06065_),
    .X(_00505_));
 sg13g2_nor2_1 _13914_ (.A(_05301_),
    .B(_05595_),
    .Y(_06066_));
 sg13g2_o21ai_1 _13915_ (.B1(_05393_),
    .Y(_06067_),
    .A1(_05741_),
    .A2(_06066_));
 sg13g2_a22oi_1 _13916_ (.Y(_06068_),
    .B1(_05739_),
    .B2(_06067_),
    .A2(net122),
    .A1(\clock_inst.sec_c[53] ));
 sg13g2_inv_1 _13917_ (.Y(_00506_),
    .A(_06068_));
 sg13g2_inv_1 _13918_ (.Y(_06069_),
    .A(\clock_inst.sec_c[5] ));
 sg13g2_nand3_1 _13919_ (.B(net274),
    .C(net369),
    .A(net164),
    .Y(_06070_));
 sg13g2_o21ai_1 _13920_ (.B1(_06070_),
    .Y(_06071_),
    .A1(net460),
    .A2(_04947_));
 sg13g2_o21ai_1 _13921_ (.B1(_05051_),
    .Y(_06072_),
    .A1(_04973_),
    .A2(_05064_));
 sg13g2_a22oi_1 _13922_ (.Y(_06073_),
    .B1(_06072_),
    .B2(_05202_),
    .A2(_05034_),
    .A1(net166));
 sg13g2_o21ai_1 _13923_ (.B1(_05699_),
    .Y(_06074_),
    .A1(net275),
    .A2(_06073_));
 sg13g2_a221oi_1 _13924_ (.B2(net189),
    .C1(_06074_),
    .B1(_06071_),
    .A1(net183),
    .Y(_06075_),
    .A2(_05186_));
 sg13g2_a22oi_1 _13925_ (.Y(_06076_),
    .B1(net169),
    .B2(_05460_),
    .A2(_04978_),
    .A1(net460));
 sg13g2_a21oi_1 _13926_ (.A1(_04925_),
    .A2(_04985_),
    .Y(_06077_),
    .B1(_05098_));
 sg13g2_o21ai_1 _13927_ (.B1(_05298_),
    .Y(_06078_),
    .A1(_05761_),
    .A2(_06077_));
 sg13g2_o21ai_1 _13928_ (.B1(_06078_),
    .Y(_06079_),
    .A1(net260),
    .A2(_06076_));
 sg13g2_nand2_1 _13929_ (.Y(_06080_),
    .A(net116),
    .B(_06079_));
 sg13g2_a22oi_1 _13930_ (.Y(_00507_),
    .B1(_06075_),
    .B2(_06080_),
    .A2(net121),
    .A1(_06069_));
 sg13g2_inv_1 _13931_ (.Y(_06081_),
    .A(\clock_inst.sec_c[6] ));
 sg13g2_nor2_1 _13932_ (.A(net404),
    .B(_05581_),
    .Y(_06082_));
 sg13g2_a21oi_1 _13933_ (.A1(net259),
    .A2(_05094_),
    .Y(_06083_),
    .B1(_06082_));
 sg13g2_a21oi_1 _13934_ (.A1(net367),
    .A2(net403),
    .Y(_06084_),
    .B1(_05042_));
 sg13g2_o21ai_1 _13935_ (.B1(_05262_),
    .Y(_06085_),
    .A1(_04954_),
    .A2(_05272_));
 sg13g2_a221oi_1 _13936_ (.B2(_06085_),
    .C1(_05020_),
    .B1(_06084_),
    .A1(net178),
    .Y(_06086_),
    .A2(_06083_));
 sg13g2_o21ai_1 _13937_ (.B1(_05321_),
    .Y(_06087_),
    .A1(_04881_),
    .A2(net250));
 sg13g2_a21oi_1 _13938_ (.A1(_04964_),
    .A2(_06087_),
    .Y(_06088_),
    .B1(_04977_));
 sg13g2_nand2_1 _13939_ (.Y(_06089_),
    .A(_04904_),
    .B(_05124_));
 sg13g2_a22oi_1 _13940_ (.Y(_06090_),
    .B1(_06089_),
    .B2(_05011_),
    .A2(_05057_),
    .A1(net258));
 sg13g2_nor2_1 _13941_ (.A(net456),
    .B(_06090_),
    .Y(_06091_));
 sg13g2_nor4_1 _13942_ (.A(_05888_),
    .B(_06086_),
    .C(_06088_),
    .D(_06091_),
    .Y(_06092_));
 sg13g2_a21oi_1 _13943_ (.A1(_06081_),
    .A2(_05049_),
    .Y(_00508_),
    .B1(_06092_));
 sg13g2_a21oi_1 _13944_ (.A1(net259),
    .A2(net368),
    .Y(_06093_),
    .B1(net248));
 sg13g2_nor2_1 _13945_ (.A(net281),
    .B(net261),
    .Y(_06094_));
 sg13g2_a21oi_1 _13946_ (.A1(net251),
    .A2(_05621_),
    .Y(_06095_),
    .B1(_06094_));
 sg13g2_o21ai_1 _13947_ (.B1(_06095_),
    .Y(_06096_),
    .A1(net186),
    .A2(_06093_));
 sg13g2_nand2_1 _13948_ (.Y(_06097_),
    .A(_04969_),
    .B(_05411_));
 sg13g2_a22oi_1 _13949_ (.Y(_06098_),
    .B1(_06097_),
    .B2(net251),
    .A2(net391),
    .A1(net402));
 sg13g2_nor3_1 _13950_ (.A(net471),
    .B(_04843_),
    .C(_05070_),
    .Y(_06099_));
 sg13g2_o21ai_1 _13951_ (.B1(net371),
    .Y(_06100_),
    .A1(_05460_),
    .A2(_06099_));
 sg13g2_o21ai_1 _13952_ (.B1(_06100_),
    .Y(_06101_),
    .A1(net249),
    .A2(_06098_));
 sg13g2_a221oi_1 _13953_ (.B2(net118),
    .C1(_06101_),
    .B1(_06096_),
    .A1(net267),
    .Y(_06102_),
    .A2(_05229_));
 sg13g2_mux2_1 _13954_ (.A0(\clock_inst.sec_c[7] ),
    .A1(_06102_),
    .S(net57),
    .X(_00509_));
 sg13g2_o21ai_1 _13955_ (.B1(_04863_),
    .Y(_06103_),
    .A1(net471),
    .A2(net276));
 sg13g2_a221oi_1 _13956_ (.B2(net263),
    .C1(_05386_),
    .B1(_06103_),
    .A1(net268),
    .Y(_06104_),
    .A2(_06097_));
 sg13g2_a22oi_1 _13957_ (.Y(_06105_),
    .B1(_05289_),
    .B2(_05233_),
    .A2(_05100_),
    .A1(net289));
 sg13g2_nand2_1 _13958_ (.Y(_06106_),
    .A(net389),
    .B(_06105_));
 sg13g2_a21oi_1 _13959_ (.A1(net394),
    .A2(_04989_),
    .Y(_06107_),
    .B1(_05168_));
 sg13g2_nand2_1 _13960_ (.Y(_06108_),
    .A(net175),
    .B(_06107_));
 sg13g2_a221oi_1 _13961_ (.B2(_06108_),
    .C1(net251),
    .B1(_06106_),
    .A1(net173),
    .Y(_06109_),
    .A2(_05701_));
 sg13g2_a21oi_1 _13962_ (.A1(net163),
    .A2(_06104_),
    .Y(_06110_),
    .B1(_06109_));
 sg13g2_nor3_1 _13963_ (.A(_05005_),
    .B(_05115_),
    .C(_06110_),
    .Y(_06111_));
 sg13g2_a21o_1 _13964_ (.A2(net120),
    .A1(\clock_inst.sec_c[8] ),
    .B1(_06111_),
    .X(_00510_));
 sg13g2_a22oi_1 _13965_ (.Y(_06112_),
    .B1(_05684_),
    .B2(net402),
    .A2(net273),
    .A1(net268));
 sg13g2_nand2b_1 _13966_ (.Y(_06113_),
    .B(net188),
    .A_N(_06112_));
 sg13g2_a21oi_1 _13967_ (.A1(_05009_),
    .A2(_05402_),
    .Y(_06114_),
    .B1(net271));
 sg13g2_nor3_1 _13968_ (.A(_04952_),
    .B(_05386_),
    .C(_06114_),
    .Y(_06115_));
 sg13g2_o21ai_1 _13969_ (.B1(net175),
    .Y(_06116_),
    .A1(_04960_),
    .A2(_04878_));
 sg13g2_nand2_1 _13970_ (.Y(_06117_),
    .A(net187),
    .B(_06116_));
 sg13g2_o21ai_1 _13971_ (.B1(_05073_),
    .Y(_06118_),
    .A1(net368),
    .A2(_05123_));
 sg13g2_a21oi_1 _13972_ (.A1(_05529_),
    .A2(_06118_),
    .Y(_06119_),
    .B1(net277));
 sg13g2_a221oi_1 _13973_ (.B2(_04974_),
    .C1(_06119_),
    .B1(_06117_),
    .A1(net190),
    .Y(_06120_),
    .A2(_05896_));
 sg13g2_a221oi_1 _13974_ (.B2(net189),
    .C1(net122),
    .B1(_06120_),
    .A1(_06113_),
    .Y(_06121_),
    .A2(_06115_));
 sg13g2_a21o_1 _13975_ (.A2(net120),
    .A1(\clock_inst.sec_c[9] ),
    .B1(_06121_),
    .X(_00511_));
 sg13g2_buf_1 _13976_ (.A(\clock_inst.sec_tile.e0[0] ),
    .X(_06122_));
 sg13g2_inv_1 _13977_ (.Y(_06123_),
    .A(_06122_));
 sg13g2_xor2_1 _13978_ (.B(_06122_),
    .A(_05422_),
    .X(_06124_));
 sg13g2_nor2_1 _13979_ (.A(net141),
    .B(_06124_),
    .Y(_06125_));
 sg13g2_a21oi_1 _13980_ (.A1(_05648_),
    .A2(net97),
    .Y(_06126_),
    .B1(_06125_));
 sg13g2_nand2_1 _13981_ (.Y(_06127_),
    .A(net142),
    .B(_06126_));
 sg13g2_o21ai_1 _13982_ (.B1(_06127_),
    .Y(_00512_),
    .A1(_06123_),
    .A2(net139));
 sg13g2_buf_1 _13983_ (.A(\clock_inst.sec_tile.e0[10] ),
    .X(_06128_));
 sg13g2_inv_1 _13984_ (.Y(_06129_),
    .A(_06128_));
 sg13g2_inv_1 _13985_ (.Y(_06130_),
    .A(\clock_inst.sec_tile.e0[6] ));
 sg13g2_buf_1 _13986_ (.A(\clock_inst.sec_tile.e0[7] ),
    .X(_06131_));
 sg13g2_nor2_1 _13987_ (.A(_05643_),
    .B(_06131_),
    .Y(_06132_));
 sg13g2_buf_1 _13988_ (.A(\clock_inst.sec_tile.e0[2] ),
    .X(_06133_));
 sg13g2_buf_2 _13989_ (.A(\clock_inst.sec_tile.e0[1] ),
    .X(_06134_));
 sg13g2_or2_1 _13990_ (.X(_06135_),
    .B(_06134_),
    .A(_05443_));
 sg13g2_and2_1 _13991_ (.A(_05422_),
    .B(_06122_),
    .X(_06136_));
 sg13g2_and2_1 _13992_ (.A(_05443_),
    .B(_06134_),
    .X(_06137_));
 sg13g2_a221oi_1 _13993_ (.B2(_06136_),
    .C1(_06137_),
    .B1(_06135_),
    .A1(_05472_),
    .Y(_06138_),
    .A2(_06133_));
 sg13g2_inv_1 _13994_ (.Y(_06139_),
    .A(_06138_));
 sg13g2_buf_1 _13995_ (.A(\clock_inst.sec_tile.e0[3] ),
    .X(_06140_));
 sg13g2_or2_1 _13996_ (.X(_06141_),
    .B(_06133_),
    .A(_05472_));
 sg13g2_nand2_1 _13997_ (.Y(_06142_),
    .A(_06140_),
    .B(_06141_));
 sg13g2_inv_1 _13998_ (.Y(_06143_),
    .A(_06142_));
 sg13g2_buf_1 _13999_ (.A(\clock_inst.sec_tile.e0[4] ),
    .X(_06144_));
 sg13g2_inv_1 _14000_ (.Y(_06145_),
    .A(_06144_));
 sg13g2_buf_1 _14001_ (.A(\clock_inst.sec_tile.e0[5] ),
    .X(_06146_));
 sg13g2_nand2_1 _14002_ (.Y(_06147_),
    .A(_05615_),
    .B(_06146_));
 sg13g2_nand2_1 _14003_ (.Y(_06148_),
    .A(_06145_),
    .B(_06147_));
 sg13g2_nand2b_1 _14004_ (.Y(_06149_),
    .B(_06147_),
    .A_N(_05613_));
 sg13g2_nor2_1 _14005_ (.A(_05443_),
    .B(_06134_),
    .Y(_06150_));
 sg13g2_a22oi_1 _14006_ (.Y(_06151_),
    .B1(_05443_),
    .B2(_06134_),
    .A2(_06122_),
    .A1(_05422_));
 sg13g2_o21ai_1 _14007_ (.B1(_05558_),
    .Y(_06152_),
    .A1(_05472_),
    .A2(_06133_));
 sg13g2_nor3_1 _14008_ (.A(_06150_),
    .B(_06151_),
    .C(_06152_),
    .Y(_06153_));
 sg13g2_and2_1 _14009_ (.A(_05472_),
    .B(_06133_),
    .X(_06154_));
 sg13g2_o21ai_1 _14010_ (.B1(_05558_),
    .Y(_06155_),
    .A1(_06140_),
    .A2(_06154_));
 sg13g2_nand2b_1 _14011_ (.Y(_06156_),
    .B(_06155_),
    .A_N(_06153_));
 sg13g2_a221oi_1 _14012_ (.B2(_06149_),
    .C1(_06156_),
    .B1(_06148_),
    .A1(_06139_),
    .Y(_06157_),
    .A2(_06143_));
 sg13g2_buf_2 _14013_ (.A(_06157_),
    .X(_06158_));
 sg13g2_nand3b_1 _14014_ (.B(_06145_),
    .C(_06147_),
    .Y(_06159_),
    .A_N(_05613_));
 sg13g2_o21ai_1 _14015_ (.B1(_06159_),
    .Y(_06160_),
    .A1(_05615_),
    .A2(_06146_));
 sg13g2_buf_1 _14016_ (.A(_06160_),
    .X(_06161_));
 sg13g2_nor4_1 _14017_ (.A(_06130_),
    .B(_06132_),
    .C(_06158_),
    .D(_06161_),
    .Y(_06162_));
 sg13g2_nor4_1 _14018_ (.A(_05632_),
    .B(_06132_),
    .C(_06158_),
    .D(_06161_),
    .Y(_06163_));
 sg13g2_nand2_1 _14019_ (.Y(_06164_),
    .A(_05631_),
    .B(\clock_inst.sec_tile.e0[6] ));
 sg13g2_nand2_1 _14020_ (.Y(_06165_),
    .A(_05643_),
    .B(_06131_));
 sg13g2_o21ai_1 _14021_ (.B1(_06165_),
    .Y(_06166_),
    .A1(_06132_),
    .A2(_06164_));
 sg13g2_nor3_2 _14022_ (.A(_06162_),
    .B(_06163_),
    .C(_06166_),
    .Y(_06167_));
 sg13g2_nor2b_1 _14023_ (.A(\clock_inst.sec_tile.e0[8] ),
    .B_N(_05424_),
    .Y(_06168_));
 sg13g2_buf_1 _14024_ (.A(_06168_),
    .X(_06169_));
 sg13g2_and2_1 _14025_ (.A(_06167_),
    .B(_06169_),
    .X(_06170_));
 sg13g2_buf_1 _14026_ (.A(_06170_),
    .X(_06171_));
 sg13g2_inv_1 _14027_ (.Y(_06172_),
    .A(\clock_inst.sec_tile.e0[8] ));
 sg13g2_nor2_1 _14028_ (.A(_05424_),
    .B(_06172_),
    .Y(_06173_));
 sg13g2_nor2b_1 _14029_ (.A(_06167_),
    .B_N(_06173_),
    .Y(_06174_));
 sg13g2_buf_1 _14030_ (.A(_06174_),
    .X(_06175_));
 sg13g2_buf_2 _14031_ (.A(\clock_inst.sec_tile.e0[9] ),
    .X(_06176_));
 sg13g2_mux2_1 _14032_ (.A0(_06171_),
    .A1(_06175_),
    .S(_06176_),
    .X(_06177_));
 sg13g2_o21ai_1 _14033_ (.B1(net155),
    .Y(_06178_),
    .A1(net48),
    .A2(_06177_));
 sg13g2_nor2_1 _14034_ (.A(_06129_),
    .B(net96),
    .Y(_06179_));
 sg13g2_nor2_1 _14035_ (.A(\clock_inst.sec_c[10] ),
    .B(net87),
    .Y(_06180_));
 sg13g2_a21o_1 _14036_ (.A2(_06179_),
    .A1(_06177_),
    .B1(_06180_),
    .X(_06181_));
 sg13g2_a22oi_1 _14037_ (.Y(_00513_),
    .B1(_06181_),
    .B2(net103),
    .A2(_06178_),
    .A1(_06129_));
 sg13g2_and2_1 _14038_ (.A(_06176_),
    .B(_06128_),
    .X(_06182_));
 sg13g2_buf_1 _14039_ (.A(_06182_),
    .X(_06183_));
 sg13g2_buf_8 _14040_ (.A(_06167_),
    .X(_06184_));
 sg13g2_nor2_1 _14041_ (.A(_06176_),
    .B(_06128_),
    .Y(_06185_));
 sg13g2_and3_1 _14042_ (.X(_06186_),
    .A(net26),
    .B(_06169_),
    .C(_06185_));
 sg13g2_a21o_1 _14043_ (.A2(_06183_),
    .A1(_06175_),
    .B1(_06186_),
    .X(_06187_));
 sg13g2_buf_1 _14044_ (.A(\clock_inst.sec_tile.e0[11] ),
    .X(_06188_));
 sg13g2_nor2_1 _14045_ (.A(_06188_),
    .B(_01377_),
    .Y(_06189_));
 sg13g2_a22oi_1 _14046_ (.Y(_06190_),
    .B1(_06187_),
    .B2(_06189_),
    .A2(net48),
    .A1(\clock_inst.sec_c[11] ));
 sg13g2_a221oi_1 _14047_ (.B2(_06175_),
    .C1(_01263_),
    .B1(_06183_),
    .A1(_06171_),
    .Y(_06191_),
    .A2(_06185_));
 sg13g2_o21ai_1 _14048_ (.B1(_06188_),
    .Y(_06192_),
    .A1(net160),
    .A2(_06191_));
 sg13g2_o21ai_1 _14049_ (.B1(_06192_),
    .Y(_00514_),
    .A1(net112),
    .A2(_06190_));
 sg13g2_inv_1 _14050_ (.Y(_06193_),
    .A(\clock_inst.sec_tile.e0[12] ));
 sg13g2_nand2_1 _14051_ (.Y(_06194_),
    .A(\clock_inst.sec_tile.e0[12] ),
    .B(_01201_));
 sg13g2_nand2_1 _14052_ (.Y(_06195_),
    .A(_06193_),
    .B(_01201_));
 sg13g2_nand3_1 _14053_ (.B(_06173_),
    .C(_06183_),
    .A(_06188_),
    .Y(_06196_));
 sg13g2_nand3b_1 _14054_ (.B(_06169_),
    .C(_06185_),
    .Y(_06197_),
    .A_N(_06188_));
 sg13g2_mux2_1 _14055_ (.A0(_06196_),
    .A1(_06197_),
    .S(net26),
    .X(_06198_));
 sg13g2_mux2_1 _14056_ (.A0(_06194_),
    .A1(_06195_),
    .S(_06198_),
    .X(_06199_));
 sg13g2_nand2b_1 _14057_ (.Y(_06200_),
    .B(net237),
    .A_N(\clock_inst.sec_c[12] ));
 sg13g2_a21oi_1 _14058_ (.A1(_06199_),
    .A2(_06200_),
    .Y(_06201_),
    .B1(net140));
 sg13g2_a21oi_1 _14059_ (.A1(_06193_),
    .A2(_04134_),
    .Y(_00515_),
    .B1(_06201_));
 sg13g2_inv_1 _14060_ (.Y(_06202_),
    .A(\clock_inst.sec_tile.e0[13] ));
 sg13g2_nand2_1 _14061_ (.Y(_06203_),
    .A(_06202_),
    .B(net92));
 sg13g2_nand2_1 _14062_ (.Y(_06204_),
    .A(\clock_inst.sec_tile.e0[13] ),
    .B(_01356_));
 sg13g2_nor4_1 _14063_ (.A(_06176_),
    .B(_06128_),
    .C(_06188_),
    .D(\clock_inst.sec_tile.e0[12] ),
    .Y(_06205_));
 sg13g2_nand3_1 _14064_ (.B(\clock_inst.sec_tile.e0[12] ),
    .C(_06183_),
    .A(_06188_),
    .Y(_06206_));
 sg13g2_inv_1 _14065_ (.Y(_06207_),
    .A(_06206_));
 sg13g2_a22oi_1 _14066_ (.Y(_06208_),
    .B1(_06207_),
    .B2(_06175_),
    .A2(_06205_),
    .A1(_06171_));
 sg13g2_mux2_1 _14067_ (.A0(_06203_),
    .A1(_06204_),
    .S(_06208_),
    .X(_06209_));
 sg13g2_a21oi_1 _14068_ (.A1(\clock_inst.sec_c[13] ),
    .A2(net52),
    .Y(_06210_),
    .B1(net162));
 sg13g2_a22oi_1 _14069_ (.Y(_00516_),
    .B1(_06209_),
    .B2(_06210_),
    .A2(net69),
    .A1(_06202_));
 sg13g2_buf_1 _14070_ (.A(\clock_inst.sec_tile.e0[14] ),
    .X(_06211_));
 sg13g2_nor4_1 _14071_ (.A(_05424_),
    .B(_06172_),
    .C(_06202_),
    .D(_06206_),
    .Y(_06212_));
 sg13g2_and3_1 _14072_ (.X(_06213_),
    .A(_06202_),
    .B(_06169_),
    .C(_06205_));
 sg13g2_mux2_1 _14073_ (.A0(_06212_),
    .A1(_06213_),
    .S(_06184_),
    .X(_06214_));
 sg13g2_xnor2_1 _14074_ (.Y(_06215_),
    .A(_06211_),
    .B(_06214_));
 sg13g2_nand2_1 _14075_ (.Y(_06216_),
    .A(\clock_inst.sec_c[14] ),
    .B(net237));
 sg13g2_o21ai_1 _14076_ (.B1(_06216_),
    .Y(_06217_),
    .A1(net98),
    .A2(_06215_));
 sg13g2_mux2_1 _14077_ (.A0(_06211_),
    .A1(_06217_),
    .S(_01381_),
    .X(_00517_));
 sg13g2_inv_1 _14078_ (.Y(_06218_),
    .A(\clock_inst.sec_tile.e0[15] ));
 sg13g2_nand2_1 _14079_ (.Y(_06219_),
    .A(_06211_),
    .B(_06212_));
 sg13g2_nand2b_1 _14080_ (.Y(_06220_),
    .B(_06213_),
    .A_N(_06211_));
 sg13g2_mux2_1 _14081_ (.A0(_06219_),
    .A1(_06220_),
    .S(net26),
    .X(_06221_));
 sg13g2_xnor2_1 _14082_ (.Y(_06222_),
    .A(_06218_),
    .B(_06221_));
 sg13g2_nand2_1 _14083_ (.Y(_06223_),
    .A(\clock_inst.sec_c[15] ),
    .B(net237));
 sg13g2_o21ai_1 _14084_ (.B1(_06223_),
    .Y(_06224_),
    .A1(net98),
    .A2(_06222_));
 sg13g2_mux2_1 _14085_ (.A0(\clock_inst.sec_tile.e0[15] ),
    .A1(_06224_),
    .S(_01381_),
    .X(_00518_));
 sg13g2_inv_1 _14086_ (.Y(_06225_),
    .A(\clock_inst.sec_tile.e0[16] ));
 sg13g2_nand3b_1 _14087_ (.B(net26),
    .C(_06218_),
    .Y(_06226_),
    .A_N(_06220_));
 sg13g2_or3_1 _14088_ (.A(_06218_),
    .B(net26),
    .C(_06219_),
    .X(_06227_));
 sg13g2_and3_1 _14089_ (.X(_06228_),
    .A(\clock_inst.sec_tile.e0[16] ),
    .B(_06226_),
    .C(_06227_));
 sg13g2_a21oi_1 _14090_ (.A1(_06226_),
    .A2(_06227_),
    .Y(_06229_),
    .B1(\clock_inst.sec_tile.e0[16] ));
 sg13g2_o21ai_1 _14091_ (.B1(_01179_),
    .Y(_06230_),
    .A1(_06228_),
    .A2(_06229_));
 sg13g2_a21oi_1 _14092_ (.A1(\clock_inst.sec_c[16] ),
    .A2(net52),
    .Y(_06231_),
    .B1(net154));
 sg13g2_a22oi_1 _14093_ (.Y(_00519_),
    .B1(_06230_),
    .B2(_06231_),
    .A2(net69),
    .A1(_06225_));
 sg13g2_inv_1 _14094_ (.Y(_06232_),
    .A(\clock_inst.sec_tile.e0[17] ));
 sg13g2_nand2_1 _14095_ (.Y(_06233_),
    .A(_06232_),
    .B(net92));
 sg13g2_nand2_1 _14096_ (.Y(_06234_),
    .A(\clock_inst.sec_tile.e0[17] ),
    .B(net92));
 sg13g2_nor2b_1 _14097_ (.A(_06220_),
    .B_N(net26),
    .Y(_06235_));
 sg13g2_nor2_1 _14098_ (.A(\clock_inst.sec_tile.e0[15] ),
    .B(\clock_inst.sec_tile.e0[16] ),
    .Y(_06236_));
 sg13g2_nor4_1 _14099_ (.A(_06218_),
    .B(_06225_),
    .C(_06184_),
    .D(_06219_),
    .Y(_06237_));
 sg13g2_a21oi_1 _14100_ (.A1(_06235_),
    .A2(_06236_),
    .Y(_06238_),
    .B1(_06237_));
 sg13g2_mux2_1 _14101_ (.A0(_06233_),
    .A1(_06234_),
    .S(_06238_),
    .X(_06239_));
 sg13g2_a21oi_1 _14102_ (.A1(\clock_inst.sec_c[17] ),
    .A2(net52),
    .Y(_06240_),
    .B1(net154));
 sg13g2_a22oi_1 _14103_ (.Y(_00520_),
    .B1(_06239_),
    .B2(_06240_),
    .A2(net69),
    .A1(_06232_));
 sg13g2_buf_2 _14104_ (.A(\clock_inst.sec_tile.e0[18] ),
    .X(_06241_));
 sg13g2_nand3_1 _14105_ (.B(net559),
    .C(net102),
    .A(_06241_),
    .Y(_06242_));
 sg13g2_o21ai_1 _14106_ (.B1(_06242_),
    .Y(_06243_),
    .A1(net559),
    .A2(net50));
 sg13g2_a21oi_1 _14107_ (.A1(net559),
    .A2(net155),
    .Y(_06244_),
    .B1(_06241_));
 sg13g2_a21oi_1 _14108_ (.A1(net88),
    .A2(_06243_),
    .Y(_00521_),
    .B1(_06244_));
 sg13g2_buf_1 _14109_ (.A(\clock_inst.sec_tile.e0[19] ),
    .X(_06245_));
 sg13g2_inv_1 _14110_ (.Y(_06246_),
    .A(_06245_));
 sg13g2_nand2_1 _14111_ (.Y(_06247_),
    .A(_06241_),
    .B(net559));
 sg13g2_xor2_1 _14112_ (.B(_06245_),
    .A(_05428_),
    .X(_06248_));
 sg13g2_xnor2_1 _14113_ (.Y(_06249_),
    .A(_06247_),
    .B(_06248_));
 sg13g2_nand2_1 _14114_ (.Y(_06250_),
    .A(net157),
    .B(_06249_));
 sg13g2_o21ai_1 _14115_ (.B1(_06250_),
    .Y(_06251_),
    .A1(_05743_),
    .A2(net101));
 sg13g2_nor2_1 _14116_ (.A(_04066_),
    .B(_06251_),
    .Y(_06252_));
 sg13g2_a21oi_1 _14117_ (.A1(_06246_),
    .A2(net67),
    .Y(_00522_),
    .B1(_06252_));
 sg13g2_inv_1 _14118_ (.Y(_06253_),
    .A(_06134_));
 sg13g2_xnor2_1 _14119_ (.Y(_06254_),
    .A(_05443_),
    .B(_06134_));
 sg13g2_xnor2_1 _14120_ (.Y(_06255_),
    .A(_06136_),
    .B(_06254_));
 sg13g2_nand2_1 _14121_ (.Y(_06256_),
    .A(net157),
    .B(_06255_));
 sg13g2_o21ai_1 _14122_ (.B1(_06256_),
    .Y(_06257_),
    .A1(_05755_),
    .A2(net101));
 sg13g2_nor2_1 _14123_ (.A(_04066_),
    .B(_06257_),
    .Y(_06258_));
 sg13g2_a21oi_1 _14124_ (.A1(_06253_),
    .A2(net67),
    .Y(_00523_),
    .B1(_06258_));
 sg13g2_inv_1 _14125_ (.Y(_06259_),
    .A(\clock_inst.sec_tile.e0[20] ));
 sg13g2_buf_1 _14126_ (.A(net244),
    .X(_06260_));
 sg13g2_nor2_1 _14127_ (.A(_05428_),
    .B(_06245_),
    .Y(_06261_));
 sg13g2_a22oi_1 _14128_ (.Y(_06262_),
    .B1(_05428_),
    .B2(_06245_),
    .A2(net559),
    .A1(_06241_));
 sg13g2_nor2_1 _14129_ (.A(_06261_),
    .B(_06262_),
    .Y(_06263_));
 sg13g2_xnor2_1 _14130_ (.Y(_06264_),
    .A(\clock_inst.sec_b[20] ),
    .B(\clock_inst.sec_tile.e0[20] ));
 sg13g2_xnor2_1 _14131_ (.Y(_06265_),
    .A(_06263_),
    .B(_06264_));
 sg13g2_nor2_1 _14132_ (.A(net159),
    .B(_06265_),
    .Y(_06266_));
 sg13g2_a21oi_1 _14133_ (.A1(_05767_),
    .A2(net97),
    .Y(_06267_),
    .B1(_06266_));
 sg13g2_nor2_1 _14134_ (.A(net113),
    .B(_06267_),
    .Y(_06268_));
 sg13g2_a21oi_1 _14135_ (.A1(_06259_),
    .A2(net67),
    .Y(_00524_),
    .B1(_06268_));
 sg13g2_buf_1 _14136_ (.A(\clock_inst.sec_tile.e0[21] ),
    .X(_06269_));
 sg13g2_buf_1 _14137_ (.A(_06269_),
    .X(_06270_));
 sg13g2_inv_1 _14138_ (.Y(_06271_),
    .A(net521));
 sg13g2_buf_1 _14139_ (.A(net153),
    .X(_06272_));
 sg13g2_o21ai_1 _14140_ (.B1(_06259_),
    .Y(_06273_),
    .A1(_06261_),
    .A2(_06262_));
 sg13g2_nor3_1 _14141_ (.A(_06259_),
    .B(_06261_),
    .C(_06262_),
    .Y(_06274_));
 sg13g2_a21o_1 _14142_ (.A2(_06273_),
    .A1(\clock_inst.sec_b[20] ),
    .B1(_06274_),
    .X(_06275_));
 sg13g2_buf_1 _14143_ (.A(_06275_),
    .X(_06276_));
 sg13g2_buf_1 _14144_ (.A(net557),
    .X(_06277_));
 sg13g2_xor2_1 _14145_ (.B(net521),
    .A(net520),
    .X(_06278_));
 sg13g2_xnor2_1 _14146_ (.Y(_06279_),
    .A(net246),
    .B(_06278_));
 sg13g2_nor2_1 _14147_ (.A(\clock_inst.sec_c[21] ),
    .B(net238),
    .Y(_06280_));
 sg13g2_a21oi_1 _14148_ (.A1(net84),
    .A2(_06279_),
    .Y(_06281_),
    .B1(_06280_));
 sg13g2_nor2_1 _14149_ (.A(net113),
    .B(_06281_),
    .Y(_06282_));
 sg13g2_a21oi_1 _14150_ (.A1(_06271_),
    .A2(net55),
    .Y(_00525_),
    .B1(_06282_));
 sg13g2_buf_1 _14151_ (.A(\clock_inst.sec_tile.e0[22] ),
    .X(_06283_));
 sg13g2_inv_1 _14152_ (.Y(_06284_),
    .A(_06283_));
 sg13g2_and2_1 _14153_ (.A(_06269_),
    .B(net246),
    .X(_06285_));
 sg13g2_buf_1 _14154_ (.A(_06285_),
    .X(_06286_));
 sg13g2_nor3_1 _14155_ (.A(net522),
    .B(net521),
    .C(net246),
    .Y(_06287_));
 sg13g2_a21o_1 _14156_ (.A2(_06286_),
    .A1(net522),
    .B1(_06287_),
    .X(_06288_));
 sg13g2_xnor2_1 _14157_ (.Y(_06289_),
    .A(_06283_),
    .B(_06288_));
 sg13g2_nand2_1 _14158_ (.Y(_06290_),
    .A(\clock_inst.sec_c[22] ),
    .B(net141));
 sg13g2_o21ai_1 _14159_ (.B1(_06290_),
    .Y(_06291_),
    .A1(net90),
    .A2(_06289_));
 sg13g2_nor2_1 _14160_ (.A(net113),
    .B(_06291_),
    .Y(_06292_));
 sg13g2_a21oi_1 _14161_ (.A1(_06284_),
    .A2(net55),
    .Y(_00526_),
    .B1(_06292_));
 sg13g2_buf_1 _14162_ (.A(\clock_inst.sec_tile.e0[23] ),
    .X(_06293_));
 sg13g2_inv_1 _14163_ (.Y(_06294_),
    .A(_06293_));
 sg13g2_nor3_1 _14164_ (.A(net521),
    .B(_06283_),
    .C(net246),
    .Y(_06295_));
 sg13g2_nor2_1 _14165_ (.A(net520),
    .B(_06284_),
    .Y(_06296_));
 sg13g2_a22oi_1 _14166_ (.Y(_06297_),
    .B1(_06296_),
    .B2(_06286_),
    .A2(_06295_),
    .A1(net520));
 sg13g2_xnor2_1 _14167_ (.Y(_06298_),
    .A(_06294_),
    .B(_06297_));
 sg13g2_nand2_1 _14168_ (.Y(_06299_),
    .A(\clock_inst.sec_c[23] ),
    .B(net141));
 sg13g2_o21ai_1 _14169_ (.B1(_06299_),
    .Y(_06300_),
    .A1(net90),
    .A2(_06298_));
 sg13g2_nor2_1 _14170_ (.A(net113),
    .B(_06300_),
    .Y(_06301_));
 sg13g2_a21oi_1 _14171_ (.A1(_06294_),
    .A2(net55),
    .Y(_00527_),
    .B1(_06301_));
 sg13g2_buf_2 _14172_ (.A(\clock_inst.sec_tile.e0[24] ),
    .X(_06302_));
 sg13g2_inv_1 _14173_ (.Y(_06303_),
    .A(_06302_));
 sg13g2_buf_1 _14174_ (.A(net151),
    .X(_06304_));
 sg13g2_nor2_1 _14175_ (.A(_06284_),
    .B(_06294_),
    .Y(_06305_));
 sg13g2_a21o_1 _14176_ (.A2(_06305_),
    .A1(net246),
    .B1(net557),
    .X(_06306_));
 sg13g2_or3_1 _14177_ (.A(_06283_),
    .B(_06293_),
    .C(net246),
    .X(_06307_));
 sg13g2_a22oi_1 _14178_ (.Y(_06308_),
    .B1(_06307_),
    .B2(net557),
    .A2(_06306_),
    .A1(net521));
 sg13g2_xnor2_1 _14179_ (.Y(_06309_),
    .A(net520),
    .B(_06302_));
 sg13g2_xnor2_1 _14180_ (.Y(_06310_),
    .A(_06308_),
    .B(_06309_));
 sg13g2_nor2_1 _14181_ (.A(\clock_inst.sec_c[24] ),
    .B(net238),
    .Y(_06311_));
 sg13g2_a21oi_1 _14182_ (.A1(_06304_),
    .A2(_06310_),
    .Y(_06312_),
    .B1(_06311_));
 sg13g2_nor2_1 _14183_ (.A(_06260_),
    .B(_06312_),
    .Y(_06313_));
 sg13g2_a21oi_1 _14184_ (.A1(_06303_),
    .A2(net55),
    .Y(_00528_),
    .B1(_06313_));
 sg13g2_buf_1 _14185_ (.A(\clock_inst.sec_tile.e0[25] ),
    .X(_06314_));
 sg13g2_and2_1 _14186_ (.A(_06302_),
    .B(_06305_),
    .X(_06315_));
 sg13g2_a21o_1 _14187_ (.A2(_06315_),
    .A1(_06276_),
    .B1(net557),
    .X(_06316_));
 sg13g2_or4_1 _14188_ (.A(_06283_),
    .B(_06293_),
    .C(_06302_),
    .D(net246),
    .X(_06317_));
 sg13g2_buf_2 _14189_ (.A(_06317_),
    .X(_06318_));
 sg13g2_a22oi_1 _14190_ (.Y(_06319_),
    .B1(_06318_),
    .B2(net520),
    .A2(_06316_),
    .A1(net521));
 sg13g2_xnor2_1 _14191_ (.Y(_06320_),
    .A(net520),
    .B(_06319_));
 sg13g2_nand3_1 _14192_ (.B(net102),
    .C(_06320_),
    .A(_06314_),
    .Y(_06321_));
 sg13g2_o21ai_1 _14193_ (.B1(_06321_),
    .Y(_06322_),
    .A1(\clock_inst.sec_c[25] ),
    .A2(net51));
 sg13g2_o21ai_1 _14194_ (.B1(net125),
    .Y(_06323_),
    .A1(net47),
    .A2(_06320_));
 sg13g2_inv_1 _14195_ (.Y(_06324_),
    .A(_06314_));
 sg13g2_a22oi_1 _14196_ (.Y(_00529_),
    .B1(_06323_),
    .B2(_06324_),
    .A2(_06322_),
    .A1(net108));
 sg13g2_buf_1 _14197_ (.A(\clock_inst.sec_tile.e0[26] ),
    .X(_06325_));
 sg13g2_inv_1 _14198_ (.Y(_06326_),
    .A(_06325_));
 sg13g2_nand3b_1 _14199_ (.B(_06324_),
    .C(_06271_),
    .Y(_06327_),
    .A_N(_06318_));
 sg13g2_nand3_1 _14200_ (.B(_06293_),
    .C(net246),
    .A(net521),
    .Y(_06328_));
 sg13g2_nand3_1 _14201_ (.B(_06302_),
    .C(_06314_),
    .A(_06283_),
    .Y(_06329_));
 sg13g2_a21oi_1 _14202_ (.A1(net522),
    .A2(_06328_),
    .Y(_06330_),
    .B1(_06329_));
 sg13g2_a21o_1 _14203_ (.A2(_06327_),
    .A1(net557),
    .B1(_06330_),
    .X(_06331_));
 sg13g2_buf_1 _14204_ (.A(_06331_),
    .X(_06332_));
 sg13g2_xor2_1 _14205_ (.B(_06325_),
    .A(net520),
    .X(_06333_));
 sg13g2_xnor2_1 _14206_ (.Y(_06334_),
    .A(_06332_),
    .B(_06333_));
 sg13g2_nor2_1 _14207_ (.A(\clock_inst.sec_c[26] ),
    .B(_01215_),
    .Y(_06335_));
 sg13g2_a21oi_1 _14208_ (.A1(net94),
    .A2(_06334_),
    .Y(_06336_),
    .B1(_06335_));
 sg13g2_nand2_1 _14209_ (.Y(_06337_),
    .A(net142),
    .B(_06336_));
 sg13g2_o21ai_1 _14210_ (.B1(_06337_),
    .Y(_00530_),
    .A1(_06326_),
    .A2(net139));
 sg13g2_buf_1 _14211_ (.A(\clock_inst.sec_tile.e0[27] ),
    .X(_06338_));
 sg13g2_nor2_1 _14212_ (.A(_06324_),
    .B(_06326_),
    .Y(_06339_));
 sg13g2_nand2_1 _14213_ (.Y(_06340_),
    .A(net522),
    .B(_06339_));
 sg13g2_nand3_1 _14214_ (.B(_06324_),
    .C(_06326_),
    .A(net557),
    .Y(_06341_));
 sg13g2_or3_1 _14215_ (.A(net521),
    .B(_06318_),
    .C(_06341_),
    .X(_06342_));
 sg13g2_o21ai_1 _14216_ (.B1(_06342_),
    .Y(_06343_),
    .A1(_06319_),
    .A2(_06340_));
 sg13g2_nand3_1 _14217_ (.B(net102),
    .C(_06343_),
    .A(_06338_),
    .Y(_06344_));
 sg13g2_o21ai_1 _14218_ (.B1(_06344_),
    .Y(_06345_),
    .A1(\clock_inst.sec_c[27] ),
    .A2(net51));
 sg13g2_o21ai_1 _14219_ (.B1(net125),
    .Y(_06346_),
    .A1(net47),
    .A2(_06343_));
 sg13g2_inv_1 _14220_ (.Y(_06347_),
    .A(_06338_));
 sg13g2_a22oi_1 _14221_ (.Y(_00531_),
    .B1(_06346_),
    .B2(_06347_),
    .A2(_06345_),
    .A1(net108));
 sg13g2_buf_1 _14222_ (.A(\clock_inst.sec_tile.e0[28] ),
    .X(_06348_));
 sg13g2_inv_1 _14223_ (.Y(_06349_),
    .A(_06348_));
 sg13g2_nor2_1 _14224_ (.A(_06338_),
    .B(_06341_),
    .Y(_06350_));
 sg13g2_nand2_1 _14225_ (.Y(_06351_),
    .A(_06308_),
    .B(_06350_));
 sg13g2_and4_1 _14226_ (.A(_06338_),
    .B(_06286_),
    .C(_06305_),
    .D(_06339_),
    .X(_06352_));
 sg13g2_o21ai_1 _14227_ (.B1(_06302_),
    .Y(_06353_),
    .A1(net557),
    .A2(_06352_));
 sg13g2_mux2_1 _14228_ (.A0(_06277_),
    .A1(_06351_),
    .S(_06353_),
    .X(_06354_));
 sg13g2_xnor2_1 _14229_ (.Y(_06355_),
    .A(_06348_),
    .B(_06354_));
 sg13g2_a21o_1 _14230_ (.A2(net107),
    .A1(\clock_inst.sec_c[28] ),
    .B1(net244),
    .X(_06356_));
 sg13g2_a21oi_1 _14231_ (.A1(net91),
    .A2(_06355_),
    .Y(_06357_),
    .B1(_06356_));
 sg13g2_a21oi_1 _14232_ (.A1(_06349_),
    .A2(_06272_),
    .Y(_00532_),
    .B1(_06357_));
 sg13g2_buf_1 _14233_ (.A(\clock_inst.sec_tile.e0[29] ),
    .X(_06358_));
 sg13g2_inv_1 _14234_ (.Y(_06359_),
    .A(_06358_));
 sg13g2_or2_1 _14235_ (.X(_06360_),
    .B(_06348_),
    .A(_06338_));
 sg13g2_nor2_1 _14236_ (.A(\clock_inst.sec_b[21] ),
    .B(_06349_),
    .Y(_06361_));
 sg13g2_and2_1 _14237_ (.A(_06338_),
    .B(_06361_),
    .X(_06362_));
 sg13g2_buf_1 _14238_ (.A(_06362_),
    .X(_06363_));
 sg13g2_nand4_1 _14239_ (.B(_06316_),
    .C(_06339_),
    .A(_06270_),
    .Y(_06364_),
    .D(_06363_));
 sg13g2_o21ai_1 _14240_ (.B1(_06364_),
    .Y(_06365_),
    .A1(_06342_),
    .A2(_06360_));
 sg13g2_xnor2_1 _14241_ (.Y(_06366_),
    .A(_06358_),
    .B(_06365_));
 sg13g2_nand2_1 _14242_ (.Y(_06367_),
    .A(\clock_inst.sec_c[29] ),
    .B(net141));
 sg13g2_o21ai_1 _14243_ (.B1(_06367_),
    .Y(_06368_),
    .A1(net90),
    .A2(_06366_));
 sg13g2_nor2_1 _14244_ (.A(_06260_),
    .B(_06368_),
    .Y(_06369_));
 sg13g2_a21oi_1 _14245_ (.A1(_06359_),
    .A2(_06272_),
    .Y(_00533_),
    .B1(_06369_));
 sg13g2_inv_1 _14246_ (.Y(_06370_),
    .A(_06133_));
 sg13g2_nor2_1 _14247_ (.A(_06150_),
    .B(_06151_),
    .Y(_06371_));
 sg13g2_xnor2_1 _14248_ (.Y(_06372_),
    .A(_05472_),
    .B(_06133_));
 sg13g2_xnor2_1 _14249_ (.Y(_06373_),
    .A(_06371_),
    .B(_06372_));
 sg13g2_nor2_1 _14250_ (.A(net159),
    .B(_06373_),
    .Y(_06374_));
 sg13g2_a21oi_1 _14251_ (.A1(_05852_),
    .A2(net97),
    .Y(_06375_),
    .B1(_06374_));
 sg13g2_nor2_1 _14252_ (.A(net113),
    .B(_06375_),
    .Y(_06376_));
 sg13g2_a21oi_1 _14253_ (.A1(_06370_),
    .A2(net55),
    .Y(_00534_),
    .B1(_06376_));
 sg13g2_buf_2 _14254_ (.A(\clock_inst.sec_tile.e0[30] ),
    .X(_06377_));
 sg13g2_and2_1 _14255_ (.A(_05864_),
    .B(_01610_),
    .X(_06378_));
 sg13g2_buf_2 _14256_ (.A(_06378_),
    .X(_06379_));
 sg13g2_a21oi_1 _14257_ (.A1(_06377_),
    .A2(net136),
    .Y(_06380_),
    .B1(_06379_));
 sg13g2_nor2_1 _14258_ (.A(_06358_),
    .B(_06360_),
    .Y(_06381_));
 sg13g2_nand3_1 _14259_ (.B(_06326_),
    .C(_06381_),
    .A(_05486_),
    .Y(_06382_));
 sg13g2_nand4_1 _14260_ (.B(_06358_),
    .C(_06330_),
    .A(_06325_),
    .Y(_06383_),
    .D(_06363_));
 sg13g2_o21ai_1 _14261_ (.B1(_06383_),
    .Y(_06384_),
    .A1(_06332_),
    .A2(_06382_));
 sg13g2_xor2_1 _14262_ (.B(_06384_),
    .A(_06377_),
    .X(_06385_));
 sg13g2_nand2_1 _14263_ (.Y(_06386_),
    .A(net23),
    .B(_06385_));
 sg13g2_nand2_1 _14264_ (.Y(_00535_),
    .A(_06380_),
    .B(_06386_));
 sg13g2_buf_1 _14265_ (.A(\clock_inst.sec_tile.e0[31] ),
    .X(_06387_));
 sg13g2_and2_1 _14266_ (.A(_06358_),
    .B(_06377_),
    .X(_06388_));
 sg13g2_buf_1 _14267_ (.A(_06388_),
    .X(_06389_));
 sg13g2_nor2_1 _14268_ (.A(net522),
    .B(_06377_),
    .Y(_06390_));
 sg13g2_a22oi_1 _14269_ (.Y(_06391_),
    .B1(_06390_),
    .B2(_06381_),
    .A2(_06389_),
    .A1(_06363_));
 sg13g2_nor2_1 _14270_ (.A(_06377_),
    .B(net556),
    .Y(_06392_));
 sg13g2_nand2_1 _14271_ (.Y(_06393_),
    .A(_06381_),
    .B(_06392_));
 sg13g2_inv_1 _14272_ (.Y(_06394_),
    .A(_06393_));
 sg13g2_nand4_1 _14273_ (.B(_06325_),
    .C(_06276_),
    .A(_06269_),
    .Y(_06395_),
    .D(_06315_));
 sg13g2_a21o_1 _14274_ (.A2(_06395_),
    .A1(net522),
    .B1(_06324_),
    .X(_06396_));
 sg13g2_buf_1 _14275_ (.A(_06396_),
    .X(_06397_));
 sg13g2_nand2_1 _14276_ (.Y(_06398_),
    .A(_06271_),
    .B(_06326_));
 sg13g2_nor2_1 _14277_ (.A(_06318_),
    .B(_06398_),
    .Y(_06399_));
 sg13g2_and2_1 _14278_ (.A(_06397_),
    .B(_06399_),
    .X(_06400_));
 sg13g2_mux2_1 _14279_ (.A0(net556),
    .A1(_06394_),
    .S(_06400_),
    .X(_06401_));
 sg13g2_or3_1 _14280_ (.A(net556),
    .B(_06391_),
    .C(_06397_),
    .X(_06402_));
 sg13g2_nand2_1 _14281_ (.Y(_06403_),
    .A(net556),
    .B(_06397_));
 sg13g2_a21oi_1 _14282_ (.A1(_06402_),
    .A2(_06403_),
    .Y(_06404_),
    .B1(_06277_));
 sg13g2_a221oi_1 _14283_ (.B2(net520),
    .C1(_06404_),
    .B1(_06401_),
    .A1(net556),
    .Y(_06405_),
    .A2(_06391_));
 sg13g2_o21ai_1 _14284_ (.B1(net233),
    .Y(_06406_),
    .A1(_05864_),
    .A2(net94));
 sg13g2_a21oi_1 _14285_ (.A1(net45),
    .A2(_06405_),
    .Y(_06407_),
    .B1(_06406_));
 sg13g2_a21o_1 _14286_ (.A2(net76),
    .A1(_06387_),
    .B1(_06407_),
    .X(_00536_));
 sg13g2_buf_2 _14287_ (.A(\clock_inst.sec_tile.e0[32] ),
    .X(_06408_));
 sg13g2_a21oi_1 _14288_ (.A1(_06408_),
    .A2(net136),
    .Y(_06409_),
    .B1(_06379_));
 sg13g2_nand3_1 _14289_ (.B(_06361_),
    .C(_06389_),
    .A(net556),
    .Y(_06410_));
 sg13g2_nor4_1 _14290_ (.A(_06302_),
    .B(_06348_),
    .C(_06377_),
    .D(net556),
    .Y(_06411_));
 sg13g2_nand4_1 _14291_ (.B(_06308_),
    .C(_06350_),
    .A(_06359_),
    .Y(_06412_),
    .D(_06411_));
 sg13g2_o21ai_1 _14292_ (.B1(_06412_),
    .Y(_06413_),
    .A1(_06353_),
    .A2(_06410_));
 sg13g2_xor2_1 _14293_ (.B(_06413_),
    .A(_06408_),
    .X(_06414_));
 sg13g2_nand2_1 _14294_ (.Y(_06415_),
    .A(_01241_),
    .B(_06414_));
 sg13g2_nand2_1 _14295_ (.Y(_00537_),
    .A(_06409_),
    .B(_06415_));
 sg13g2_inv_1 _14296_ (.Y(_06416_),
    .A(\clock_inst.sec_tile.e0[33] ));
 sg13g2_nand3_1 _14297_ (.B(_06408_),
    .C(_06389_),
    .A(net556),
    .Y(_06417_));
 sg13g2_nor4_1 _14298_ (.A(_06270_),
    .B(_06408_),
    .C(_06341_),
    .D(_06393_),
    .Y(_06418_));
 sg13g2_nand2b_1 _14299_ (.Y(_06419_),
    .B(_06418_),
    .A_N(_06318_));
 sg13g2_o21ai_1 _14300_ (.B1(_06419_),
    .Y(_06420_),
    .A1(_06364_),
    .A2(_06417_));
 sg13g2_xnor2_1 _14301_ (.Y(_06421_),
    .A(_06416_),
    .B(_06420_));
 sg13g2_a21oi_1 _14302_ (.A1(net49),
    .A2(_06421_),
    .Y(_06422_),
    .B1(_06379_));
 sg13g2_o21ai_1 _14303_ (.B1(_06422_),
    .Y(_00538_),
    .A1(_06416_),
    .A2(net139));
 sg13g2_buf_1 _14304_ (.A(\clock_inst.sec_tile.e0[34] ),
    .X(_06423_));
 sg13g2_nor3_1 _14305_ (.A(net522),
    .B(_06408_),
    .C(\clock_inst.sec_tile.e0[33] ),
    .Y(_06424_));
 sg13g2_nor2b_1 _14306_ (.A(_06393_),
    .B_N(_06424_),
    .Y(_06425_));
 sg13g2_and2_1 _14307_ (.A(_06326_),
    .B(_06425_),
    .X(_06426_));
 sg13g2_nand3_1 _14308_ (.B(_06358_),
    .C(_06363_),
    .A(_06325_),
    .Y(_06427_));
 sg13g2_and4_1 _14309_ (.A(_05487_),
    .B(_06387_),
    .C(_06408_),
    .D(\clock_inst.sec_tile.e0[33] ),
    .X(_06428_));
 sg13g2_a22oi_1 _14310_ (.Y(_06429_),
    .B1(_06424_),
    .B2(_06392_),
    .A2(_06428_),
    .A1(_06377_));
 sg13g2_a21oi_1 _14311_ (.A1(_06382_),
    .A2(_06427_),
    .Y(_06430_),
    .B1(_06429_));
 sg13g2_nand2_1 _14312_ (.Y(_06431_),
    .A(_06332_),
    .B(_06430_));
 sg13g2_mux2_1 _14313_ (.A0(_05487_),
    .A1(_06426_),
    .S(_06431_),
    .X(_06432_));
 sg13g2_xnor2_1 _14314_ (.Y(_06433_),
    .A(_06423_),
    .B(_06432_));
 sg13g2_a21oi_1 _14315_ (.A1(_06423_),
    .A2(net145),
    .Y(_06434_),
    .B1(_06379_));
 sg13g2_o21ai_1 _14316_ (.B1(_06434_),
    .Y(_00539_),
    .A1(net44),
    .A2(_06433_));
 sg13g2_a21oi_1 _14317_ (.A1(\clock_inst.sec_tile.e0[35] ),
    .A2(net136),
    .Y(_06435_),
    .B1(_06379_));
 sg13g2_nand2b_1 _14318_ (.Y(_06436_),
    .B(_06425_),
    .A_N(_06423_));
 sg13g2_nand2_1 _14319_ (.Y(_06437_),
    .A(_06423_),
    .B(_06428_));
 sg13g2_o21ai_1 _14320_ (.B1(_05486_),
    .Y(_06438_),
    .A1(_06318_),
    .A2(_06398_));
 sg13g2_a21oi_1 _14321_ (.A1(_06397_),
    .A2(_06438_),
    .Y(_06439_),
    .B1(_06391_));
 sg13g2_mux2_1 _14322_ (.A0(_06436_),
    .A1(_06437_),
    .S(_06439_),
    .X(_06440_));
 sg13g2_xnor2_1 _14323_ (.Y(_06441_),
    .A(\clock_inst.sec_tile.e0[35] ),
    .B(_06440_));
 sg13g2_nand2_1 _14324_ (.Y(_06442_),
    .A(net23),
    .B(_06441_));
 sg13g2_nand2_1 _14325_ (.Y(_00540_),
    .A(_06435_),
    .B(_06442_));
 sg13g2_buf_8 _14326_ (.A(\clock_inst.sec_tile.e0[36] ),
    .X(_06443_));
 sg13g2_inv_1 _14327_ (.Y(_06444_),
    .A(_06443_));
 sg13g2_xor2_1 _14328_ (.B(_06443_),
    .A(_05489_),
    .X(_06445_));
 sg13g2_nor2_1 _14329_ (.A(_01655_),
    .B(_06445_),
    .Y(_06446_));
 sg13g2_a21oi_1 _14330_ (.A1(_05867_),
    .A2(net97),
    .Y(_06447_),
    .B1(_06446_));
 sg13g2_nand2_1 _14331_ (.Y(_06448_),
    .A(net142),
    .B(_06447_));
 sg13g2_o21ai_1 _14332_ (.B1(_06448_),
    .Y(_00541_),
    .A1(_06444_),
    .A2(net139));
 sg13g2_buf_8 _14333_ (.A(\clock_inst.sec_tile.e0[37] ),
    .X(_06449_));
 sg13g2_inv_1 _14334_ (.Y(_06450_),
    .A(_06449_));
 sg13g2_nand2_1 _14335_ (.Y(_06451_),
    .A(_05489_),
    .B(_06443_));
 sg13g2_xor2_1 _14336_ (.B(_06449_),
    .A(_05506_),
    .X(_06452_));
 sg13g2_xnor2_1 _14337_ (.Y(_06453_),
    .A(_06451_),
    .B(_06452_));
 sg13g2_nand2_1 _14338_ (.Y(_06454_),
    .A(net157),
    .B(_06453_));
 sg13g2_o21ai_1 _14339_ (.B1(_06454_),
    .Y(_06455_),
    .A1(_05879_),
    .A2(net101));
 sg13g2_nor2_1 _14340_ (.A(net113),
    .B(_06455_),
    .Y(_06456_));
 sg13g2_a21oi_1 _14341_ (.A1(_06450_),
    .A2(net55),
    .Y(_00542_),
    .B1(_06456_));
 sg13g2_buf_2 _14342_ (.A(\clock_inst.sec_tile.e0[38] ),
    .X(_06457_));
 sg13g2_inv_1 _14343_ (.Y(_06458_),
    .A(_06457_));
 sg13g2_nor2_1 _14344_ (.A(_05506_),
    .B(_06449_),
    .Y(_06459_));
 sg13g2_a22oi_1 _14345_ (.Y(_06460_),
    .B1(_05506_),
    .B2(_06449_),
    .A2(_06443_),
    .A1(_05489_));
 sg13g2_nor2_1 _14346_ (.A(_06459_),
    .B(_06460_),
    .Y(_06461_));
 sg13g2_xnor2_1 _14347_ (.Y(_06462_),
    .A(_05520_),
    .B(_06457_));
 sg13g2_xnor2_1 _14348_ (.Y(_06463_),
    .A(_06461_),
    .B(_06462_));
 sg13g2_nor2_1 _14349_ (.A(net159),
    .B(_06463_),
    .Y(_06464_));
 sg13g2_a21oi_1 _14350_ (.A1(_05890_),
    .A2(net97),
    .Y(_06465_),
    .B1(_06464_));
 sg13g2_nor2_1 _14351_ (.A(net113),
    .B(_06465_),
    .Y(_06466_));
 sg13g2_a21oi_1 _14352_ (.A1(_06458_),
    .A2(net55),
    .Y(_00543_),
    .B1(_06466_));
 sg13g2_buf_1 _14353_ (.A(\clock_inst.sec_tile.e0[39] ),
    .X(_06467_));
 sg13g2_inv_1 _14354_ (.Y(_06468_),
    .A(_06467_));
 sg13g2_or2_1 _14355_ (.X(_06469_),
    .B(_06457_),
    .A(_05520_));
 sg13g2_buf_1 _14356_ (.A(_06469_),
    .X(_06470_));
 sg13g2_and2_1 _14357_ (.A(_05520_),
    .B(_06457_),
    .X(_06471_));
 sg13g2_buf_1 _14358_ (.A(_06471_),
    .X(_06472_));
 sg13g2_a21oi_1 _14359_ (.A1(_06461_),
    .A2(_06470_),
    .Y(_06473_),
    .B1(_06472_));
 sg13g2_xnor2_1 _14360_ (.Y(_06474_),
    .A(_05536_),
    .B(_06467_));
 sg13g2_xnor2_1 _14361_ (.Y(_06475_),
    .A(_06473_),
    .B(_06474_));
 sg13g2_nor2_1 _14362_ (.A(\clock_inst.sec_c[39] ),
    .B(net238),
    .Y(_06476_));
 sg13g2_a21oi_1 _14363_ (.A1(net54),
    .A2(_06475_),
    .Y(_06477_),
    .B1(_06476_));
 sg13g2_nor2_1 _14364_ (.A(net113),
    .B(_06477_),
    .Y(_06478_));
 sg13g2_a21oi_1 _14365_ (.A1(_06468_),
    .A2(net55),
    .Y(_00544_),
    .B1(_06478_));
 sg13g2_inv_1 _14366_ (.Y(_06479_),
    .A(_06140_));
 sg13g2_a21oi_1 _14367_ (.A1(_06371_),
    .A2(_06141_),
    .Y(_06480_),
    .B1(_06154_));
 sg13g2_xnor2_1 _14368_ (.Y(_06481_),
    .A(_05558_),
    .B(_06140_));
 sg13g2_xnor2_1 _14369_ (.Y(_06482_),
    .A(_06480_),
    .B(_06481_));
 sg13g2_nor2_1 _14370_ (.A(\clock_inst.sec_c[3] ),
    .B(net238),
    .Y(_06483_));
 sg13g2_a21oi_1 _14371_ (.A1(net54),
    .A2(_06482_),
    .Y(_06484_),
    .B1(_06483_));
 sg13g2_nor2_1 _14372_ (.A(net147),
    .B(_06484_),
    .Y(_06485_));
 sg13g2_a21oi_1 _14373_ (.A1(_06479_),
    .A2(net105),
    .Y(_00545_),
    .B1(_06485_));
 sg13g2_buf_2 _14374_ (.A(\clock_inst.sec_tile.e0[40] ),
    .X(_06486_));
 sg13g2_inv_1 _14375_ (.Y(_06487_),
    .A(_06486_));
 sg13g2_a221oi_1 _14376_ (.B2(_06470_),
    .C1(_06472_),
    .B1(_06461_),
    .A1(_05536_),
    .Y(_06488_),
    .A2(_06467_));
 sg13g2_nor2_1 _14377_ (.A(_05536_),
    .B(_06467_),
    .Y(_06489_));
 sg13g2_nor2_1 _14378_ (.A(_06488_),
    .B(_06489_),
    .Y(_06490_));
 sg13g2_xor2_1 _14379_ (.B(_06486_),
    .A(_05561_),
    .X(_06491_));
 sg13g2_xnor2_1 _14380_ (.Y(_06492_),
    .A(_06490_),
    .B(_06491_));
 sg13g2_nor2_1 _14381_ (.A(\clock_inst.sec_c[40] ),
    .B(net238),
    .Y(_06493_));
 sg13g2_a21oi_1 _14382_ (.A1(net54),
    .A2(_06492_),
    .Y(_06494_),
    .B1(_06493_));
 sg13g2_nor2_1 _14383_ (.A(net147),
    .B(_06494_),
    .Y(_06495_));
 sg13g2_a21oi_1 _14384_ (.A1(_06487_),
    .A2(net105),
    .Y(_00546_),
    .B1(_06495_));
 sg13g2_buf_2 _14385_ (.A(\clock_inst.sec_tile.e0[41] ),
    .X(_06496_));
 sg13g2_xor2_1 _14386_ (.B(_06496_),
    .A(_05573_),
    .X(_06497_));
 sg13g2_a21o_1 _14387_ (.A2(_06490_),
    .A1(_06486_),
    .B1(_05561_),
    .X(_06498_));
 sg13g2_o21ai_1 _14388_ (.B1(_06498_),
    .Y(_06499_),
    .A1(_06486_),
    .A2(_06490_));
 sg13g2_xor2_1 _14389_ (.B(_06499_),
    .A(_06497_),
    .X(_06500_));
 sg13g2_nand2_1 _14390_ (.Y(_06501_),
    .A(net54),
    .B(_06500_));
 sg13g2_o21ai_1 _14391_ (.B1(_06501_),
    .Y(_06502_),
    .A1(\clock_inst.sec_c[41] ),
    .A2(net93));
 sg13g2_nor2_1 _14392_ (.A(_06496_),
    .B(net144),
    .Y(_06503_));
 sg13g2_a21oi_1 _14393_ (.A1(net88),
    .A2(_06502_),
    .Y(_00547_),
    .B1(_06503_));
 sg13g2_buf_1 _14394_ (.A(\clock_inst.sec_tile.e0[42] ),
    .X(_06504_));
 sg13g2_inv_1 _14395_ (.Y(_06505_),
    .A(_06504_));
 sg13g2_and2_1 _14396_ (.A(_06491_),
    .B(_06497_),
    .X(_06506_));
 sg13g2_nand2b_1 _14397_ (.Y(_06507_),
    .B(_06506_),
    .A_N(_06489_));
 sg13g2_nor2_1 _14398_ (.A(_05573_),
    .B(_06496_),
    .Y(_06508_));
 sg13g2_a22oi_1 _14399_ (.Y(_06509_),
    .B1(_05573_),
    .B2(_06496_),
    .A2(_06486_),
    .A1(_05561_));
 sg13g2_or2_1 _14400_ (.X(_06510_),
    .B(_06509_),
    .A(_06508_));
 sg13g2_o21ai_1 _14401_ (.B1(_06510_),
    .Y(_06511_),
    .A1(_06488_),
    .A2(_06507_));
 sg13g2_xor2_1 _14402_ (.B(_06504_),
    .A(\clock_inst.sec_b[42] ),
    .X(_06512_));
 sg13g2_xnor2_1 _14403_ (.Y(_06513_),
    .A(_06511_),
    .B(_06512_));
 sg13g2_nor2_1 _14404_ (.A(\clock_inst.sec_c[42] ),
    .B(net235),
    .Y(_06514_));
 sg13g2_a21oi_1 _14405_ (.A1(net94),
    .A2(_06513_),
    .Y(_06515_),
    .B1(_06514_));
 sg13g2_nand2_1 _14406_ (.Y(_06516_),
    .A(net142),
    .B(_06515_));
 sg13g2_o21ai_1 _14407_ (.B1(_06516_),
    .Y(_00548_),
    .A1(_06505_),
    .A2(net139));
 sg13g2_nor2b_1 _14408_ (.A(_06506_),
    .B_N(_06510_),
    .Y(_06517_));
 sg13g2_a22oi_1 _14409_ (.Y(_06518_),
    .B1(_05520_),
    .B2(_06457_),
    .A2(_06449_),
    .A1(_05506_));
 sg13g2_o21ai_1 _14410_ (.B1(_06518_),
    .Y(_06519_),
    .A1(_06451_),
    .A2(_06459_));
 sg13g2_and2_1 _14411_ (.A(_06467_),
    .B(_06470_),
    .X(_06520_));
 sg13g2_o21ai_1 _14412_ (.B1(_06505_),
    .Y(_06521_),
    .A1(_06508_),
    .A2(_06509_));
 sg13g2_a21oi_1 _14413_ (.A1(_06519_),
    .A2(_06520_),
    .Y(_06522_),
    .B1(_06521_));
 sg13g2_o21ai_1 _14414_ (.B1(_05536_),
    .Y(_06523_),
    .A1(_05520_),
    .A2(_06457_));
 sg13g2_nor3_1 _14415_ (.A(_06459_),
    .B(_06460_),
    .C(_06523_),
    .Y(_06524_));
 sg13g2_o21ai_1 _14416_ (.B1(_05536_),
    .Y(_06525_),
    .A1(_06467_),
    .A2(_06472_));
 sg13g2_nor2b_1 _14417_ (.A(_06524_),
    .B_N(_06525_),
    .Y(_06526_));
 sg13g2_inv_1 _14418_ (.Y(_06527_),
    .A(\clock_inst.sec_b[42] ));
 sg13g2_a221oi_1 _14419_ (.B2(_06526_),
    .C1(_06527_),
    .B1(_06522_),
    .A1(_06505_),
    .Y(_06528_),
    .A2(_06517_));
 sg13g2_a21o_1 _14420_ (.A2(_06511_),
    .A1(_06504_),
    .B1(_06528_),
    .X(_06529_));
 sg13g2_buf_1 _14421_ (.A(\clock_inst.sec_tile.e0[43] ),
    .X(_06530_));
 sg13g2_xor2_1 _14422_ (.B(_06530_),
    .A(_05593_),
    .X(_06531_));
 sg13g2_xnor2_1 _14423_ (.Y(_06532_),
    .A(_06529_),
    .B(_06531_));
 sg13g2_nand2_1 _14424_ (.Y(_06533_),
    .A(net54),
    .B(_06532_));
 sg13g2_o21ai_1 _14425_ (.B1(_06533_),
    .Y(_06534_),
    .A1(\clock_inst.sec_c[43] ),
    .A2(net93));
 sg13g2_nor2_1 _14426_ (.A(_06530_),
    .B(net144),
    .Y(_06535_));
 sg13g2_a21oi_1 _14427_ (.A1(net88),
    .A2(_06534_),
    .Y(_00549_),
    .B1(_06535_));
 sg13g2_buf_1 _14428_ (.A(\clock_inst.sec_tile.e0[44] ),
    .X(_06536_));
 sg13g2_inv_1 _14429_ (.Y(_06537_),
    .A(_06536_));
 sg13g2_nor2_1 _14430_ (.A(_05593_),
    .B(_06530_),
    .Y(_06538_));
 sg13g2_buf_2 _14431_ (.A(_06538_),
    .X(_06539_));
 sg13g2_a221oi_1 _14432_ (.B2(_06504_),
    .C1(_06528_),
    .B1(_06511_),
    .A1(_05593_),
    .Y(_06540_),
    .A2(_06530_));
 sg13g2_buf_2 _14433_ (.A(_06540_),
    .X(_06541_));
 sg13g2_or2_1 _14434_ (.X(_06542_),
    .B(_06541_),
    .A(_06539_));
 sg13g2_buf_2 _14435_ (.A(_06542_),
    .X(_06543_));
 sg13g2_inv_1 _14436_ (.Y(_06544_),
    .A(_05139_));
 sg13g2_buf_1 _14437_ (.A(_06544_),
    .X(_06545_));
 sg13g2_nor2_1 _14438_ (.A(net455),
    .B(_06536_),
    .Y(_06546_));
 sg13g2_nor2_1 _14439_ (.A(net457),
    .B(_06537_),
    .Y(_06547_));
 sg13g2_nor2_1 _14440_ (.A(_06546_),
    .B(_06547_),
    .Y(_06548_));
 sg13g2_xnor2_1 _14441_ (.Y(_06549_),
    .A(_06543_),
    .B(_06548_));
 sg13g2_nand2_1 _14442_ (.Y(_06550_),
    .A(\clock_inst.sec_c[44] ),
    .B(net141));
 sg13g2_o21ai_1 _14443_ (.B1(_06550_),
    .Y(_06551_),
    .A1(net90),
    .A2(_06549_));
 sg13g2_nor2_1 _14444_ (.A(net147),
    .B(_06551_),
    .Y(_06552_));
 sg13g2_a21oi_1 _14445_ (.A1(_06537_),
    .A2(net105),
    .Y(_00550_),
    .B1(_06552_));
 sg13g2_buf_1 _14446_ (.A(\clock_inst.sec_tile.e0[45] ),
    .X(_06553_));
 sg13g2_mux2_1 _14447_ (.A0(_06547_),
    .A1(_06546_),
    .S(_06543_),
    .X(_06554_));
 sg13g2_nand3_1 _14448_ (.B(net102),
    .C(_06554_),
    .A(_06553_),
    .Y(_06555_));
 sg13g2_o21ai_1 _14449_ (.B1(_06555_),
    .Y(_06556_),
    .A1(\clock_inst.sec_c[45] ),
    .A2(net51));
 sg13g2_o21ai_1 _14450_ (.B1(net125),
    .Y(_06557_),
    .A1(net47),
    .A2(_06554_));
 sg13g2_inv_1 _14451_ (.Y(_06558_),
    .A(_06553_));
 sg13g2_a22oi_1 _14452_ (.Y(_00551_),
    .B1(_06557_),
    .B2(_06558_),
    .A2(_06556_),
    .A1(net108));
 sg13g2_buf_1 _14453_ (.A(\clock_inst.sec_tile.e0[46] ),
    .X(_06559_));
 sg13g2_inv_1 _14454_ (.Y(_06560_),
    .A(_06559_));
 sg13g2_nand3_1 _14455_ (.B(_06536_),
    .C(_06553_),
    .A(net455),
    .Y(_06561_));
 sg13g2_nand3_1 _14456_ (.B(_06537_),
    .C(_06558_),
    .A(net457),
    .Y(_06562_));
 sg13g2_mux2_1 _14457_ (.A0(_06561_),
    .A1(_06562_),
    .S(_06543_),
    .X(_06563_));
 sg13g2_xnor2_1 _14458_ (.Y(_06564_),
    .A(_06559_),
    .B(_06563_));
 sg13g2_nand2_1 _14459_ (.Y(_06565_),
    .A(net51),
    .B(_06564_));
 sg13g2_a21oi_1 _14460_ (.A1(\clock_inst.sec_c[46] ),
    .A2(net52),
    .Y(_06566_),
    .B1(net154));
 sg13g2_a22oi_1 _14461_ (.Y(_00552_),
    .B1(_06565_),
    .B2(_06566_),
    .A2(_03671_),
    .A1(_06560_));
 sg13g2_buf_1 _14462_ (.A(\clock_inst.sec_tile.e0[47] ),
    .X(_06567_));
 sg13g2_nor3_1 _14463_ (.A(_06537_),
    .B(_06558_),
    .C(_06560_),
    .Y(_06568_));
 sg13g2_nand2_1 _14464_ (.Y(_06569_),
    .A(net455),
    .B(_06568_));
 sg13g2_nor4_1 _14465_ (.A(net455),
    .B(_06536_),
    .C(_06553_),
    .D(_06559_),
    .Y(_06570_));
 sg13g2_o21ai_1 _14466_ (.B1(_06570_),
    .Y(_06571_),
    .A1(_06539_),
    .A2(_06541_));
 sg13g2_o21ai_1 _14467_ (.B1(_06571_),
    .Y(_06572_),
    .A1(_06543_),
    .A2(_06569_));
 sg13g2_nand3_1 _14468_ (.B(net102),
    .C(_06572_),
    .A(_06567_),
    .Y(_06573_));
 sg13g2_o21ai_1 _14469_ (.B1(_06573_),
    .Y(_06574_),
    .A1(\clock_inst.sec_c[47] ),
    .A2(net51));
 sg13g2_o21ai_1 _14470_ (.B1(net125),
    .Y(_06575_),
    .A1(net48),
    .A2(_06572_));
 sg13g2_inv_1 _14471_ (.Y(_06576_),
    .A(_06567_));
 sg13g2_a22oi_1 _14472_ (.Y(_00553_),
    .B1(_06575_),
    .B2(_06576_),
    .A2(_06574_),
    .A1(net108));
 sg13g2_buf_1 _14473_ (.A(\clock_inst.sec_tile.e0[48] ),
    .X(_06577_));
 sg13g2_inv_1 _14474_ (.Y(_06578_),
    .A(_06577_));
 sg13g2_nand2_1 _14475_ (.Y(_06579_),
    .A(_06567_),
    .B(_06568_));
 sg13g2_or3_1 _14476_ (.A(_06539_),
    .B(_06541_),
    .C(_06579_),
    .X(_06580_));
 sg13g2_nor4_2 _14477_ (.A(_06536_),
    .B(_06553_),
    .C(_06559_),
    .Y(_06581_),
    .D(_06567_));
 sg13g2_a22oi_1 _14478_ (.Y(_06582_),
    .B1(_06581_),
    .B2(_06543_),
    .A2(_06580_),
    .A1(net455));
 sg13g2_xnor2_1 _14479_ (.Y(_06583_),
    .A(net372),
    .B(_06577_));
 sg13g2_xnor2_1 _14480_ (.Y(_06584_),
    .A(_06582_),
    .B(_06583_));
 sg13g2_nand2_1 _14481_ (.Y(_06585_),
    .A(net91),
    .B(_06584_));
 sg13g2_a21oi_1 _14482_ (.A1(\clock_inst.sec_c[48] ),
    .A2(net98),
    .Y(_06586_),
    .B1(net154));
 sg13g2_a22oi_1 _14483_ (.Y(_00554_),
    .B1(_06585_),
    .B2(_06586_),
    .A2(_03671_),
    .A1(_06578_));
 sg13g2_buf_2 _14484_ (.A(\clock_inst.sec_tile.e0[49] ),
    .X(_06587_));
 sg13g2_and2_1 _14485_ (.A(_06587_),
    .B(net99),
    .X(_06588_));
 sg13g2_nor2_1 _14486_ (.A(_06587_),
    .B(net95),
    .Y(_06589_));
 sg13g2_nor2_1 _14487_ (.A(_06544_),
    .B(_06577_),
    .Y(_06590_));
 sg13g2_and2_1 _14488_ (.A(_06581_),
    .B(_06590_),
    .X(_06591_));
 sg13g2_buf_1 _14489_ (.A(_06591_),
    .X(_06592_));
 sg13g2_o21ai_1 _14490_ (.B1(_06592_),
    .Y(_06593_),
    .A1(_06539_),
    .A2(_06541_));
 sg13g2_nand2_1 _14491_ (.Y(_06594_),
    .A(_06544_),
    .B(_06577_));
 sg13g2_or4_1 _14492_ (.A(_06539_),
    .B(_06541_),
    .C(_06579_),
    .D(_06594_),
    .X(_06595_));
 sg13g2_nand2_1 _14493_ (.Y(_06596_),
    .A(_06593_),
    .B(_06595_));
 sg13g2_mux2_1 _14494_ (.A0(_06588_),
    .A1(_06589_),
    .S(_06596_),
    .X(_06597_));
 sg13g2_a221oi_1 _14495_ (.B2(\clock_inst.sec_c[49] ),
    .C1(_06597_),
    .B1(net82),
    .A1(_06587_),
    .Y(_06598_),
    .A2(net147));
 sg13g2_inv_1 _14496_ (.Y(_00555_),
    .A(_06598_));
 sg13g2_a21o_1 _14497_ (.A2(_06143_),
    .A1(_06139_),
    .B1(_06156_),
    .X(_06599_));
 sg13g2_buf_1 _14498_ (.A(_06599_),
    .X(_06600_));
 sg13g2_xor2_1 _14499_ (.B(_06600_),
    .A(_05613_),
    .X(_06601_));
 sg13g2_nand3_1 _14500_ (.B(net102),
    .C(_06601_),
    .A(_06144_),
    .Y(_06602_));
 sg13g2_o21ai_1 _14501_ (.B1(_06602_),
    .Y(_06603_),
    .A1(\clock_inst.sec_c[4] ),
    .A2(net51));
 sg13g2_o21ai_1 _14502_ (.B1(net125),
    .Y(_06604_),
    .A1(net48),
    .A2(_06601_));
 sg13g2_a22oi_1 _14503_ (.Y(_00556_),
    .B1(_06604_),
    .B2(_06145_),
    .A2(_06603_),
    .A1(net108));
 sg13g2_buf_1 _14504_ (.A(\clock_inst.sec_tile.e0[50] ),
    .X(_06605_));
 sg13g2_inv_1 _14505_ (.Y(_06606_),
    .A(_06605_));
 sg13g2_nand2_1 _14506_ (.Y(_06607_),
    .A(_06606_),
    .B(net104));
 sg13g2_nand2_1 _14507_ (.Y(_06608_),
    .A(_06605_),
    .B(net104));
 sg13g2_mux2_1 _14508_ (.A0(_06593_),
    .A1(_06595_),
    .S(_06587_),
    .X(_06609_));
 sg13g2_mux2_1 _14509_ (.A0(_06607_),
    .A1(_06608_),
    .S(_06609_),
    .X(_06610_));
 sg13g2_a21oi_1 _14510_ (.A1(\clock_inst.sec_c[50] ),
    .A2(net48),
    .Y(_06611_),
    .B1(net153));
 sg13g2_a22oi_1 _14511_ (.Y(_00557_),
    .B1(_06610_),
    .B2(_06611_),
    .A2(net112),
    .A1(_06606_));
 sg13g2_buf_1 _14512_ (.A(\clock_inst.sec_tile.e0[51] ),
    .X(_06612_));
 sg13g2_inv_1 _14513_ (.Y(_06613_),
    .A(_06592_));
 sg13g2_nor3_1 _14514_ (.A(_06587_),
    .B(_06605_),
    .C(_06613_),
    .Y(_06614_));
 sg13g2_nand2_1 _14515_ (.Y(_06615_),
    .A(_06587_),
    .B(_06605_));
 sg13g2_nor3_1 _14516_ (.A(_06576_),
    .B(_06594_),
    .C(_06615_),
    .Y(_06616_));
 sg13g2_nor2_1 _14517_ (.A(net457),
    .B(_06568_),
    .Y(_06617_));
 sg13g2_nor3_1 _14518_ (.A(_06539_),
    .B(_06541_),
    .C(_06617_),
    .Y(_06618_));
 sg13g2_mux2_1 _14519_ (.A0(_06614_),
    .A1(_06616_),
    .S(_06618_),
    .X(_06619_));
 sg13g2_nand3_1 _14520_ (.B(net102),
    .C(_06619_),
    .A(_06612_),
    .Y(_06620_));
 sg13g2_o21ai_1 _14521_ (.B1(_06620_),
    .Y(_06621_),
    .A1(\clock_inst.sec_c[51] ),
    .A2(_01203_));
 sg13g2_o21ai_1 _14522_ (.B1(net125),
    .Y(_06622_),
    .A1(net48),
    .A2(_06619_));
 sg13g2_inv_1 _14523_ (.Y(_06623_),
    .A(_06612_));
 sg13g2_a22oi_1 _14524_ (.Y(_00558_),
    .B1(_06622_),
    .B2(_06623_),
    .A2(_06621_),
    .A1(net108));
 sg13g2_inv_1 _14525_ (.Y(_06624_),
    .A(\clock_inst.sec_tile.e0[52] ));
 sg13g2_nor3_1 _14526_ (.A(_06587_),
    .B(_06605_),
    .C(_06612_),
    .Y(_06625_));
 sg13g2_and2_1 _14527_ (.A(_06592_),
    .B(_06625_),
    .X(_06626_));
 sg13g2_nor2_1 _14528_ (.A(_06594_),
    .B(_06615_),
    .Y(_06627_));
 sg13g2_a22oi_1 _14529_ (.Y(_06628_),
    .B1(_06625_),
    .B2(_06590_),
    .A2(_06627_),
    .A1(_06612_));
 sg13g2_nor2_1 _14530_ (.A(net523),
    .B(_06579_),
    .Y(_06629_));
 sg13g2_a21oi_1 _14531_ (.A1(net523),
    .A2(_06581_),
    .Y(_06630_),
    .B1(_06629_));
 sg13g2_nor4_1 _14532_ (.A(_06539_),
    .B(_06541_),
    .C(_06628_),
    .D(_06630_),
    .Y(_06631_));
 sg13g2_mux2_1 _14533_ (.A0(_06626_),
    .A1(net455),
    .S(_06631_),
    .X(_06632_));
 sg13g2_xnor2_1 _14534_ (.Y(_06633_),
    .A(_06624_),
    .B(_06632_));
 sg13g2_a21o_1 _14535_ (.A2(net107),
    .A1(\clock_inst.sec_c[52] ),
    .B1(net244),
    .X(_06634_));
 sg13g2_a21oi_1 _14536_ (.A1(net91),
    .A2(_06633_),
    .Y(_06635_),
    .B1(_06634_));
 sg13g2_a21oi_1 _14537_ (.A1(_06624_),
    .A2(net105),
    .Y(_00559_),
    .B1(_06635_));
 sg13g2_nand4_1 _14538_ (.B(_06587_),
    .C(_06605_),
    .A(_06544_),
    .Y(_06636_),
    .D(_06612_));
 sg13g2_nor4_1 _14539_ (.A(_06624_),
    .B(_06579_),
    .C(_06594_),
    .D(_06636_),
    .Y(_06637_));
 sg13g2_nor3_1 _14540_ (.A(_06539_),
    .B(_06541_),
    .C(_06637_),
    .Y(_06638_));
 sg13g2_or2_1 _14541_ (.X(_06639_),
    .B(_06530_),
    .A(_05593_));
 sg13g2_and2_1 _14542_ (.A(_05593_),
    .B(_06530_),
    .X(_06640_));
 sg13g2_a221oi_1 _14543_ (.B2(_06624_),
    .C1(_06640_),
    .B1(_06626_),
    .A1(_06529_),
    .Y(_06641_),
    .A2(_06639_));
 sg13g2_nor2_1 _14544_ (.A(\clock_inst.sec_tile.e0[53] ),
    .B(net241),
    .Y(_06642_));
 sg13g2_o21ai_1 _14545_ (.B1(_06642_),
    .Y(_06643_),
    .A1(_06638_),
    .A2(_06641_));
 sg13g2_nand2_1 _14546_ (.Y(_06644_),
    .A(\clock_inst.sec_tile.e0[53] ),
    .B(net243));
 sg13g2_or3_1 _14547_ (.A(_06638_),
    .B(_06641_),
    .C(_06644_),
    .X(_06645_));
 sg13g2_nand2b_1 _14548_ (.Y(_06646_),
    .B(net241),
    .A_N(\clock_inst.sec_c[53] ));
 sg13g2_and4_1 _14549_ (.A(_01057_),
    .B(_06643_),
    .C(_06645_),
    .D(_06646_),
    .X(_06647_));
 sg13g2_buf_1 _14550_ (.A(_06647_),
    .X(_06648_));
 sg13g2_a21o_1 _14551_ (.A2(net76),
    .A1(\clock_inst.sec_tile.e0[53] ),
    .B1(_06648_),
    .X(_00560_));
 sg13g2_inv_1 _14552_ (.Y(_06649_),
    .A(_06146_));
 sg13g2_a21o_1 _14553_ (.A2(_06600_),
    .A1(_06144_),
    .B1(_05613_),
    .X(_06650_));
 sg13g2_o21ai_1 _14554_ (.B1(_06650_),
    .Y(_06651_),
    .A1(_06144_),
    .A2(_06600_));
 sg13g2_xnor2_1 _14555_ (.Y(_06652_),
    .A(_05615_),
    .B(_06146_));
 sg13g2_xnor2_1 _14556_ (.Y(_06653_),
    .A(_06651_),
    .B(_06652_));
 sg13g2_nor2_1 _14557_ (.A(\clock_inst.sec_c[5] ),
    .B(net238),
    .Y(_06654_));
 sg13g2_a21oi_1 _14558_ (.A1(net54),
    .A2(_06653_),
    .Y(_06655_),
    .B1(_06654_));
 sg13g2_nor2_1 _14559_ (.A(net147),
    .B(_06655_),
    .Y(_06656_));
 sg13g2_a21oi_1 _14560_ (.A1(_06649_),
    .A2(net105),
    .Y(_00561_),
    .B1(_06656_));
 sg13g2_nor2_1 _14561_ (.A(_06158_),
    .B(_06161_),
    .Y(_06657_));
 sg13g2_xor2_1 _14562_ (.B(\clock_inst.sec_tile.e0[6] ),
    .A(_05631_),
    .X(_06658_));
 sg13g2_xnor2_1 _14563_ (.Y(_06659_),
    .A(_06657_),
    .B(_06658_));
 sg13g2_nor2_1 _14564_ (.A(\clock_inst.sec_c[6] ),
    .B(net238),
    .Y(_06660_));
 sg13g2_a21oi_1 _14565_ (.A1(net54),
    .A2(_06659_),
    .Y(_06661_),
    .B1(_06660_));
 sg13g2_nor2_1 _14566_ (.A(net147),
    .B(_06661_),
    .Y(_06662_));
 sg13g2_a21oi_1 _14567_ (.A1(_06130_),
    .A2(net105),
    .Y(_00562_),
    .B1(_06662_));
 sg13g2_inv_1 _14568_ (.Y(_06663_),
    .A(_06131_));
 sg13g2_o21ai_1 _14569_ (.B1(_06130_),
    .Y(_06664_),
    .A1(_06158_),
    .A2(_06161_));
 sg13g2_nor3_1 _14570_ (.A(_06130_),
    .B(_06158_),
    .C(_06161_),
    .Y(_06665_));
 sg13g2_a21oi_1 _14571_ (.A1(_05631_),
    .A2(_06664_),
    .Y(_06666_),
    .B1(_06665_));
 sg13g2_xnor2_1 _14572_ (.Y(_06667_),
    .A(_05643_),
    .B(_06131_));
 sg13g2_xnor2_1 _14573_ (.Y(_06668_),
    .A(_06666_),
    .B(_06667_));
 sg13g2_nor2_1 _14574_ (.A(\clock_inst.sec_c[7] ),
    .B(net235),
    .Y(_06669_));
 sg13g2_a21oi_1 _14575_ (.A1(net94),
    .A2(_06668_),
    .Y(_06670_),
    .B1(_06669_));
 sg13g2_nand2_1 _14576_ (.Y(_06671_),
    .A(net142),
    .B(_06670_));
 sg13g2_o21ai_1 _14577_ (.B1(_06671_),
    .Y(_00563_),
    .A1(_06663_),
    .A2(net139));
 sg13g2_nor2_1 _14578_ (.A(_06173_),
    .B(_06169_),
    .Y(_06672_));
 sg13g2_xnor2_1 _14579_ (.Y(_06673_),
    .A(net26),
    .B(_06672_));
 sg13g2_nor2_1 _14580_ (.A(\clock_inst.sec_c[8] ),
    .B(net238),
    .Y(_06674_));
 sg13g2_a21oi_1 _14581_ (.A1(_06304_),
    .A2(_06673_),
    .Y(_06675_),
    .B1(_06674_));
 sg13g2_nor2_1 _14582_ (.A(_01347_),
    .B(_06675_),
    .Y(_06676_));
 sg13g2_a21oi_1 _14583_ (.A1(_06172_),
    .A2(net105),
    .Y(_00564_),
    .B1(_06676_));
 sg13g2_mux2_1 _14584_ (.A0(_06173_),
    .A1(_06169_),
    .S(net26),
    .X(_06677_));
 sg13g2_xor2_1 _14585_ (.B(_06677_),
    .A(_06176_),
    .X(_06678_));
 sg13g2_and2_1 _14586_ (.A(\clock_inst.sec_c[9] ),
    .B(net107),
    .X(_06679_));
 sg13g2_a21oi_1 _14587_ (.A1(net93),
    .A2(_06678_),
    .Y(_06680_),
    .B1(_06679_));
 sg13g2_nor2_1 _14588_ (.A(_06176_),
    .B(net144),
    .Y(_06681_));
 sg13g2_a21oi_1 _14589_ (.A1(net88),
    .A2(_06680_),
    .Y(_00565_),
    .B1(_06681_));
 sg13g2_nand2_1 _14590_ (.Y(_06682_),
    .A(\clock_inst.sec_a[0] ),
    .B(net355));
 sg13g2_xor2_1 _14591_ (.B(_06682_),
    .A(\clock_inst.sec_tile.e[0] ),
    .X(_06683_));
 sg13g2_o21ai_1 _14592_ (.B1(_06127_),
    .Y(_00566_),
    .A1(net135),
    .A2(_06683_));
 sg13g2_buf_1 _14593_ (.A(\clock_inst.sec_tile.e[10] ),
    .X(_06684_));
 sg13g2_buf_2 _14594_ (.A(\clock_inst.sec_tile.e[9] ),
    .X(_06685_));
 sg13g2_inv_1 _14595_ (.Y(_06686_),
    .A(\clock_inst.sec_a[3] ));
 sg13g2_inv_1 _14596_ (.Y(_06687_),
    .A(\clock_inst.sec_tile.e[3] ));
 sg13g2_buf_1 _14597_ (.A(\clock_inst.sec_tile.e[5] ),
    .X(_06688_));
 sg13g2_buf_1 _14598_ (.A(\clock_inst.sec_tile.e[4] ),
    .X(_06689_));
 sg13g2_o21ai_1 _14599_ (.B1(_06689_),
    .Y(_06690_),
    .A1(_05362_),
    .A2(_06688_));
 sg13g2_o21ai_1 _14600_ (.B1(\clock_inst.sec_a[4] ),
    .Y(_06691_),
    .A1(_05362_),
    .A2(_06688_));
 sg13g2_nand2_1 _14601_ (.Y(_06692_),
    .A(\clock_inst.sec_a[0] ),
    .B(\clock_inst.sec_tile.e[0] ));
 sg13g2_nor2_1 _14602_ (.A(\clock_inst.sec_a[1] ),
    .B(\clock_inst.sec_tile.e[1] ),
    .Y(_06693_));
 sg13g2_nand2_1 _14603_ (.Y(_06694_),
    .A(\clock_inst.sec_a[1] ),
    .B(\clock_inst.sec_tile.e[1] ));
 sg13g2_o21ai_1 _14604_ (.B1(_06694_),
    .Y(_06695_),
    .A1(_06692_),
    .A2(_06693_));
 sg13g2_or2_1 _14605_ (.X(_06696_),
    .B(\clock_inst.sec_tile.e[2] ),
    .A(_05113_));
 sg13g2_and2_1 _14606_ (.A(_05113_),
    .B(\clock_inst.sec_tile.e[2] ),
    .X(_06697_));
 sg13g2_a221oi_1 _14607_ (.B2(_06696_),
    .C1(_06697_),
    .B1(_06695_),
    .A1(\clock_inst.sec_a[3] ),
    .Y(_06698_),
    .A2(\clock_inst.sec_tile.e[3] ));
 sg13g2_a221oi_1 _14608_ (.B2(_06691_),
    .C1(_06698_),
    .B1(_06690_),
    .A1(_06686_),
    .Y(_06699_),
    .A2(_06687_));
 sg13g2_buf_2 _14609_ (.A(_06699_),
    .X(_06700_));
 sg13g2_nor2_1 _14610_ (.A(_05362_),
    .B(_06688_),
    .Y(_06701_));
 sg13g2_nand2_1 _14611_ (.Y(_06702_),
    .A(\clock_inst.sec_a[4] ),
    .B(_06689_));
 sg13g2_nand2_1 _14612_ (.Y(_06703_),
    .A(_05362_),
    .B(_06688_));
 sg13g2_o21ai_1 _14613_ (.B1(_06703_),
    .Y(_06704_),
    .A1(_06701_),
    .A2(_06702_));
 sg13g2_buf_1 _14614_ (.A(_06704_),
    .X(_06705_));
 sg13g2_buf_1 _14615_ (.A(\clock_inst.sec_tile.e[6] ),
    .X(_06706_));
 sg13g2_inv_1 _14616_ (.Y(_06707_),
    .A(_06706_));
 sg13g2_nor2_1 _14617_ (.A(_05392_),
    .B(\clock_inst.sec_tile.e[7] ),
    .Y(_06708_));
 sg13g2_nor2_1 _14618_ (.A(_06707_),
    .B(_06708_),
    .Y(_06709_));
 sg13g2_o21ai_1 _14619_ (.B1(_06709_),
    .Y(_06710_),
    .A1(_06700_),
    .A2(_06705_));
 sg13g2_inv_1 _14620_ (.Y(_06711_),
    .A(\clock_inst.sec_a[6] ));
 sg13g2_nor2_1 _14621_ (.A(_06711_),
    .B(_06708_),
    .Y(_06712_));
 sg13g2_o21ai_1 _14622_ (.B1(_06712_),
    .Y(_06713_),
    .A1(_06700_),
    .A2(_06705_));
 sg13g2_nor3_1 _14623_ (.A(_06711_),
    .B(_06707_),
    .C(_06708_),
    .Y(_06714_));
 sg13g2_a21oi_1 _14624_ (.A1(_05392_),
    .A2(\clock_inst.sec_tile.e[7] ),
    .Y(_06715_),
    .B1(_06714_));
 sg13g2_nand3_1 _14625_ (.B(_06713_),
    .C(_06715_),
    .A(_06710_),
    .Y(_06716_));
 sg13g2_buf_2 _14626_ (.A(_06716_),
    .X(_06717_));
 sg13g2_nor2b_1 _14627_ (.A(_04935_),
    .B_N(\clock_inst.sec_tile.e[8] ),
    .Y(_06718_));
 sg13g2_and4_1 _14628_ (.A(_06685_),
    .B(_01815_),
    .C(_06717_),
    .D(_06718_),
    .X(_06719_));
 sg13g2_nand2b_1 _14629_ (.Y(_06720_),
    .B(_04935_),
    .A_N(\clock_inst.sec_tile.e[8] ));
 sg13g2_nor4_1 _14630_ (.A(_06685_),
    .B(net542),
    .C(_06717_),
    .D(_06720_),
    .Y(_06721_));
 sg13g2_nor3_1 _14631_ (.A(_06684_),
    .B(_06719_),
    .C(_06721_),
    .Y(_06722_));
 sg13g2_o21ai_1 _14632_ (.B1(_06684_),
    .Y(_06723_),
    .A1(_06719_),
    .A2(_06721_));
 sg13g2_nand2b_1 _14633_ (.Y(_06724_),
    .B(_06723_),
    .A_N(_06722_));
 sg13g2_nand2_1 _14634_ (.Y(_06725_),
    .A(_06128_),
    .B(net94));
 sg13g2_nand2_1 _14635_ (.Y(_06726_),
    .A(_06129_),
    .B(net94));
 sg13g2_mux2_1 _14636_ (.A0(_06725_),
    .A1(_06726_),
    .S(_06177_),
    .X(_06727_));
 sg13g2_a21oi_1 _14637_ (.A1(\clock_inst.sec_c[10] ),
    .A2(net43),
    .Y(_06728_),
    .B1(net138));
 sg13g2_a22oi_1 _14638_ (.Y(_00567_),
    .B1(_06727_),
    .B2(_06728_),
    .A2(_06724_),
    .A1(_01062_));
 sg13g2_buf_1 _14639_ (.A(_06717_),
    .X(_06729_));
 sg13g2_and3_1 _14640_ (.X(_06730_),
    .A(_06685_),
    .B(_06684_),
    .C(_06718_));
 sg13g2_nand2_1 _14641_ (.Y(_06731_),
    .A(net25),
    .B(_06730_));
 sg13g2_or4_1 _14642_ (.A(_06685_),
    .B(_06684_),
    .C(_06717_),
    .D(_06720_),
    .X(_06732_));
 sg13g2_a21oi_1 _14643_ (.A1(_06731_),
    .A2(_06732_),
    .Y(_06733_),
    .B1(net447));
 sg13g2_xnor2_1 _14644_ (.Y(_06734_),
    .A(\clock_inst.sec_tile.e[11] ),
    .B(_06733_));
 sg13g2_nand2_1 _14645_ (.Y(_06735_),
    .A(_06188_),
    .B(net157));
 sg13g2_a221oi_1 _14646_ (.B2(_06175_),
    .C1(_06735_),
    .B1(_06183_),
    .A1(_06171_),
    .Y(_06736_),
    .A2(_06185_));
 sg13g2_a21oi_1 _14647_ (.A1(_06187_),
    .A2(_06189_),
    .Y(_06737_),
    .B1(_06736_));
 sg13g2_a21oi_1 _14648_ (.A1(\clock_inst.sec_c[11] ),
    .A2(net43),
    .Y(_06738_),
    .B1(net138));
 sg13g2_a22oi_1 _14649_ (.Y(_00568_),
    .B1(_06737_),
    .B2(_06738_),
    .A2(_06734_),
    .A1(net111));
 sg13g2_buf_1 _14650_ (.A(\clock_inst.sec_tile.e[12] ),
    .X(_06739_));
 sg13g2_nor4_2 _14651_ (.A(_06685_),
    .B(_06684_),
    .C(\clock_inst.sec_tile.e[11] ),
    .Y(_06740_),
    .D(_06720_));
 sg13g2_nand2_1 _14652_ (.Y(_06741_),
    .A(_01796_),
    .B(_06740_));
 sg13g2_and2_1 _14653_ (.A(\clock_inst.sec_tile.e[11] ),
    .B(_06730_),
    .X(_06742_));
 sg13g2_buf_1 _14654_ (.A(_06742_),
    .X(_06743_));
 sg13g2_nand3_1 _14655_ (.B(net25),
    .C(_06743_),
    .A(net442),
    .Y(_06744_));
 sg13g2_o21ai_1 _14656_ (.B1(_06744_),
    .Y(_06745_),
    .A1(net25),
    .A2(_06741_));
 sg13g2_xnor2_1 _14657_ (.Y(_06746_),
    .A(_06739_),
    .B(_06745_));
 sg13g2_a21oi_1 _14658_ (.A1(net63),
    .A2(_06746_),
    .Y(_00569_),
    .B1(_06201_));
 sg13g2_buf_1 _14659_ (.A(\clock_inst.sec_tile.e[13] ),
    .X(_06747_));
 sg13g2_nor2_1 _14660_ (.A(_06739_),
    .B(_01675_),
    .Y(_06748_));
 sg13g2_nand2_1 _14661_ (.Y(_06749_),
    .A(_06740_),
    .B(_06748_));
 sg13g2_nor2_1 _14662_ (.A(_06729_),
    .B(_06749_),
    .Y(_06750_));
 sg13g2_and4_1 _14663_ (.A(_06739_),
    .B(_01728_),
    .C(_06717_),
    .D(_06743_),
    .X(_06751_));
 sg13g2_buf_1 _14664_ (.A(_06751_),
    .X(_06752_));
 sg13g2_nor2_1 _14665_ (.A(_06750_),
    .B(_06752_),
    .Y(_06753_));
 sg13g2_xor2_1 _14666_ (.B(_06753_),
    .A(_06747_),
    .X(_06754_));
 sg13g2_a22oi_1 _14667_ (.Y(_00570_),
    .B1(_06754_),
    .B2(net78),
    .A2(_06210_),
    .A1(_06209_));
 sg13g2_buf_1 _14668_ (.A(\clock_inst.sec_tile.e[14] ),
    .X(_06755_));
 sg13g2_nor3_1 _14669_ (.A(_06747_),
    .B(_06729_),
    .C(_06749_),
    .Y(_06756_));
 sg13g2_a21oi_1 _14670_ (.A1(_06747_),
    .A2(_06752_),
    .Y(_06757_),
    .B1(_06756_));
 sg13g2_xnor2_1 _14671_ (.Y(_06758_),
    .A(_06755_),
    .B(_06757_));
 sg13g2_mux2_1 _14672_ (.A0(_06217_),
    .A1(_06758_),
    .S(net83),
    .X(_00571_));
 sg13g2_and2_1 _14673_ (.A(_06747_),
    .B(_06755_),
    .X(_06759_));
 sg13g2_nor4_1 _14674_ (.A(_06747_),
    .B(_06755_),
    .C(_06717_),
    .D(_06749_),
    .Y(_06760_));
 sg13g2_a21oi_1 _14675_ (.A1(_06752_),
    .A2(_06759_),
    .Y(_06761_),
    .B1(_06760_));
 sg13g2_xnor2_1 _14676_ (.Y(_06762_),
    .A(\clock_inst.sec_tile.e[15] ),
    .B(_06761_));
 sg13g2_mux2_1 _14677_ (.A0(_06224_),
    .A1(_06762_),
    .S(net83),
    .X(_00572_));
 sg13g2_nor3_1 _14678_ (.A(_06747_),
    .B(_06755_),
    .C(\clock_inst.sec_tile.e[15] ),
    .Y(_06763_));
 sg13g2_nand3_1 _14679_ (.B(_06748_),
    .C(_06763_),
    .A(_06740_),
    .Y(_06764_));
 sg13g2_nor2b_1 _14680_ (.A(_04935_),
    .B_N(\clock_inst.sec_tile.e[15] ),
    .Y(_06765_));
 sg13g2_and4_1 _14681_ (.A(_06739_),
    .B(_01728_),
    .C(_06759_),
    .D(_06765_),
    .X(_06766_));
 sg13g2_o21ai_1 _14682_ (.B1(_06766_),
    .Y(_06767_),
    .A1(_06743_),
    .A2(_06740_));
 sg13g2_mux2_1 _14683_ (.A0(_06764_),
    .A1(_06767_),
    .S(net25),
    .X(_06768_));
 sg13g2_xor2_1 _14684_ (.B(_06768_),
    .A(\clock_inst.sec_tile.e[16] ),
    .X(_06769_));
 sg13g2_a22oi_1 _14685_ (.Y(_00573_),
    .B1(_06769_),
    .B2(net78),
    .A2(_06231_),
    .A1(_06230_));
 sg13g2_nand3_1 _14686_ (.B(_06748_),
    .C(_06763_),
    .A(_06740_),
    .Y(_06770_));
 sg13g2_nor3_1 _14687_ (.A(\clock_inst.sec_tile.e[16] ),
    .B(net25),
    .C(_06770_),
    .Y(_06771_));
 sg13g2_nand4_1 _14688_ (.B(net25),
    .C(_06743_),
    .A(\clock_inst.sec_tile.e[16] ),
    .Y(_06772_),
    .D(_06766_));
 sg13g2_nand2b_1 _14689_ (.Y(_06773_),
    .B(_06772_),
    .A_N(_06771_));
 sg13g2_xnor2_1 _14690_ (.Y(_06774_),
    .A(\clock_inst.sec_tile.e[17] ),
    .B(_06773_));
 sg13g2_a22oi_1 _14691_ (.Y(_00574_),
    .B1(_06774_),
    .B2(net79),
    .A2(_06240_),
    .A1(_06239_));
 sg13g2_buf_2 _14692_ (.A(\clock_inst.sec_tile.e[18] ),
    .X(_06775_));
 sg13g2_nor2_1 _14693_ (.A(_06775_),
    .B(net80),
    .Y(_06776_));
 sg13g2_a22oi_1 _14694_ (.Y(_06777_),
    .B1(_01802_),
    .B2(_06775_),
    .A2(net49),
    .A1(_06241_));
 sg13g2_nor2b_1 _14695_ (.A(_06777_),
    .B_N(_05001_),
    .Y(_06778_));
 sg13g2_a221oi_1 _14696_ (.B2(_06241_),
    .C1(_05001_),
    .B1(_01805_),
    .A1(_06775_),
    .Y(_06779_),
    .A2(net154));
 sg13g2_nor3_1 _14697_ (.A(_06776_),
    .B(_06778_),
    .C(_06779_),
    .Y(_00575_));
 sg13g2_nand2_1 _14698_ (.Y(_06780_),
    .A(net559),
    .B(_06775_));
 sg13g2_xor2_1 _14699_ (.B(_06780_),
    .A(_05046_),
    .X(_06781_));
 sg13g2_nor2_1 _14700_ (.A(net405),
    .B(_06781_),
    .Y(_06782_));
 sg13g2_xnor2_1 _14701_ (.Y(_06783_),
    .A(\clock_inst.sec_tile.e[19] ),
    .B(_06782_));
 sg13g2_a21oi_1 _14702_ (.A1(net63),
    .A2(_06783_),
    .Y(_00576_),
    .B1(_06252_));
 sg13g2_xnor2_1 _14703_ (.Y(_06784_),
    .A(_05048_),
    .B(_06692_));
 sg13g2_nor2_1 _14704_ (.A(net405),
    .B(_06784_),
    .Y(_06785_));
 sg13g2_xnor2_1 _14705_ (.Y(_06786_),
    .A(\clock_inst.sec_tile.e[1] ),
    .B(_06785_));
 sg13g2_a21oi_1 _14706_ (.A1(net63),
    .A2(_06786_),
    .Y(_00577_),
    .B1(_06258_));
 sg13g2_buf_1 _14707_ (.A(\clock_inst.sec_tile.e[20] ),
    .X(_06787_));
 sg13g2_a22oi_1 _14708_ (.Y(_06788_),
    .B1(_05046_),
    .B2(\clock_inst.sec_tile.e[19] ),
    .A2(_06775_),
    .A1(net559));
 sg13g2_nor2_1 _14709_ (.A(_05046_),
    .B(\clock_inst.sec_tile.e[19] ),
    .Y(_06789_));
 sg13g2_nor2_1 _14710_ (.A(_06788_),
    .B(_06789_),
    .Y(_06790_));
 sg13g2_xnor2_1 _14711_ (.Y(_06791_),
    .A(_05090_),
    .B(_06790_));
 sg13g2_nor2_1 _14712_ (.A(net405),
    .B(_06791_),
    .Y(_06792_));
 sg13g2_xnor2_1 _14713_ (.Y(_06793_),
    .A(_06787_),
    .B(_06792_));
 sg13g2_a21oi_1 _14714_ (.A1(net63),
    .A2(_06793_),
    .Y(_00578_),
    .B1(_06268_));
 sg13g2_buf_1 _14715_ (.A(\clock_inst.sec_tile.e[21] ),
    .X(_06794_));
 sg13g2_or2_1 _14716_ (.X(_06795_),
    .B(_06787_),
    .A(_05090_));
 sg13g2_nand2_1 _14717_ (.Y(_06796_),
    .A(_05090_),
    .B(_06787_));
 sg13g2_o21ai_1 _14718_ (.B1(_06796_),
    .Y(_06797_),
    .A1(_06788_),
    .A2(_06789_));
 sg13g2_and2_1 _14719_ (.A(_06795_),
    .B(_06797_),
    .X(_06798_));
 sg13g2_buf_2 _14720_ (.A(_06798_),
    .X(_06799_));
 sg13g2_xnor2_1 _14721_ (.Y(_06800_),
    .A(net372),
    .B(_06799_));
 sg13g2_nor2_1 _14722_ (.A(net405),
    .B(_06800_),
    .Y(_06801_));
 sg13g2_xnor2_1 _14723_ (.Y(_06802_),
    .A(net555),
    .B(_06801_));
 sg13g2_a21oi_1 _14724_ (.A1(_04792_),
    .A2(_06802_),
    .Y(_00579_),
    .B1(_06282_));
 sg13g2_buf_1 _14725_ (.A(\clock_inst.sec_tile.e[22] ),
    .X(_06803_));
 sg13g2_nor2_1 _14726_ (.A(net555),
    .B(_06799_),
    .Y(_06804_));
 sg13g2_nor2b_1 _14727_ (.A(net457),
    .B_N(net555),
    .Y(_06805_));
 sg13g2_a22oi_1 _14728_ (.Y(_06806_),
    .B1(_06805_),
    .B2(_06799_),
    .A2(_06804_),
    .A1(net372));
 sg13g2_nor2_1 _14729_ (.A(net405),
    .B(_06806_),
    .Y(_06807_));
 sg13g2_xnor2_1 _14730_ (.Y(_06808_),
    .A(_06803_),
    .B(_06807_));
 sg13g2_a21oi_1 _14731_ (.A1(net63),
    .A2(_06808_),
    .Y(_00580_),
    .B1(_06292_));
 sg13g2_nand3_1 _14732_ (.B(_06799_),
    .C(_06805_),
    .A(_06803_),
    .Y(_06809_));
 sg13g2_nand3b_1 _14733_ (.B(_06804_),
    .C(net372),
    .Y(_06810_),
    .A_N(_06803_));
 sg13g2_a21oi_1 _14734_ (.A1(_06809_),
    .A2(_06810_),
    .Y(_06811_),
    .B1(net447));
 sg13g2_xnor2_1 _14735_ (.Y(_06812_),
    .A(\clock_inst.sec_tile.e[23] ),
    .B(_06811_));
 sg13g2_a21oi_1 _14736_ (.A1(net63),
    .A2(_06812_),
    .Y(_00581_),
    .B1(_06301_));
 sg13g2_buf_1 _14737_ (.A(\clock_inst.sec_tile.e[24] ),
    .X(_06813_));
 sg13g2_and4_1 _14738_ (.A(_06803_),
    .B(\clock_inst.sec_tile.e[23] ),
    .C(_06795_),
    .D(_06797_),
    .X(_06814_));
 sg13g2_buf_1 _14739_ (.A(_06814_),
    .X(_06815_));
 sg13g2_or2_1 _14740_ (.X(_06816_),
    .B(_06815_),
    .A(net523));
 sg13g2_nor2_1 _14741_ (.A(_06803_),
    .B(\clock_inst.sec_tile.e[23] ),
    .Y(_06817_));
 sg13g2_nand2b_1 _14742_ (.Y(_06818_),
    .B(_06817_),
    .A_N(_06799_));
 sg13g2_a22oi_1 _14743_ (.Y(_06819_),
    .B1(_06818_),
    .B2(net523),
    .A2(_06816_),
    .A1(_06794_));
 sg13g2_xnor2_1 _14744_ (.Y(_06820_),
    .A(net455),
    .B(_06819_));
 sg13g2_nor2_1 _14745_ (.A(net405),
    .B(_06820_),
    .Y(_06821_));
 sg13g2_xnor2_1 _14746_ (.Y(_06822_),
    .A(_06813_),
    .B(_06821_));
 sg13g2_a21oi_1 _14747_ (.A1(_04792_),
    .A2(_06822_),
    .Y(_00582_),
    .B1(_06313_));
 sg13g2_nor4_1 _14748_ (.A(net455),
    .B(net555),
    .C(_06813_),
    .D(_06818_),
    .Y(_06823_));
 sg13g2_inv_1 _14749_ (.Y(_06824_),
    .A(_06813_));
 sg13g2_nor3_1 _14750_ (.A(net372),
    .B(_06824_),
    .C(_06819_),
    .Y(_06825_));
 sg13g2_o21ai_1 _14751_ (.B1(net443),
    .Y(_06826_),
    .A1(_06823_),
    .A2(_06825_));
 sg13g2_xor2_1 _14752_ (.B(_06826_),
    .A(\clock_inst.sec_tile.e[25] ),
    .X(_06827_));
 sg13g2_xnor2_1 _14753_ (.Y(_06828_),
    .A(_06314_),
    .B(_06320_));
 sg13g2_o21ai_1 _14754_ (.B1(net233),
    .Y(_06829_),
    .A1(\clock_inst.sec_c[25] ),
    .A2(net54));
 sg13g2_a21o_1 _14755_ (.A2(_06828_),
    .A1(net50),
    .B1(_06829_),
    .X(_06830_));
 sg13g2_o21ai_1 _14756_ (.B1(_06830_),
    .Y(_00583_),
    .A1(net135),
    .A2(_06827_));
 sg13g2_buf_1 _14757_ (.A(\clock_inst.sec_tile.e[26] ),
    .X(_06831_));
 sg13g2_and2_1 _14758_ (.A(_06813_),
    .B(\clock_inst.sec_tile.e[25] ),
    .X(_06832_));
 sg13g2_buf_1 _14759_ (.A(_06832_),
    .X(_06833_));
 sg13g2_a21o_1 _14760_ (.A2(_06833_),
    .A1(_06815_),
    .B1(net523),
    .X(_06834_));
 sg13g2_nor2_1 _14761_ (.A(_06813_),
    .B(\clock_inst.sec_tile.e[25] ),
    .Y(_06835_));
 sg13g2_nand3b_1 _14762_ (.B(_06817_),
    .C(_06835_),
    .Y(_06836_),
    .A_N(_06799_));
 sg13g2_a22oi_1 _14763_ (.Y(_06837_),
    .B1(_06836_),
    .B2(net523),
    .A2(_06834_),
    .A1(net555));
 sg13g2_buf_2 _14764_ (.A(_06837_),
    .X(_06838_));
 sg13g2_xnor2_1 _14765_ (.Y(_06839_),
    .A(_06545_),
    .B(_06838_));
 sg13g2_nor2_1 _14766_ (.A(net446),
    .B(_06839_),
    .Y(_06840_));
 sg13g2_xnor2_1 _14767_ (.Y(_06841_),
    .A(net554),
    .B(_06840_));
 sg13g2_o21ai_1 _14768_ (.B1(_06337_),
    .Y(_00584_),
    .A1(_02131_),
    .A2(_06841_));
 sg13g2_buf_2 _14769_ (.A(\clock_inst.sec_tile.e[27] ),
    .X(_06842_));
 sg13g2_and2_1 _14770_ (.A(_05090_),
    .B(_06787_),
    .X(_06843_));
 sg13g2_nor2_1 _14771_ (.A(_05090_),
    .B(_06787_),
    .Y(_06844_));
 sg13g2_nor3_1 _14772_ (.A(_06788_),
    .B(_06789_),
    .C(_06844_),
    .Y(_06845_));
 sg13g2_nand2_1 _14773_ (.Y(_06846_),
    .A(_06817_),
    .B(_06835_));
 sg13g2_or4_1 _14774_ (.A(net555),
    .B(_06843_),
    .C(_06845_),
    .D(_06846_),
    .X(_06847_));
 sg13g2_buf_1 _14775_ (.A(_06847_),
    .X(_06848_));
 sg13g2_nor3_1 _14776_ (.A(_06545_),
    .B(net554),
    .C(_06848_),
    .Y(_06849_));
 sg13g2_nand4_1 _14777_ (.B(net554),
    .C(_06815_),
    .A(net555),
    .Y(_06850_),
    .D(_06833_));
 sg13g2_nor2_1 _14778_ (.A(net372),
    .B(_06850_),
    .Y(_06851_));
 sg13g2_o21ai_1 _14779_ (.B1(net355),
    .Y(_06852_),
    .A1(_06849_),
    .A2(_06851_));
 sg13g2_xor2_1 _14780_ (.B(_06852_),
    .A(_06842_),
    .X(_06853_));
 sg13g2_xnor2_1 _14781_ (.Y(_06854_),
    .A(_06347_),
    .B(_06343_));
 sg13g2_nand2_1 _14782_ (.Y(_06855_),
    .A(net45),
    .B(_06854_));
 sg13g2_a21oi_1 _14783_ (.A1(\clock_inst.sec_c[27] ),
    .A2(net43),
    .Y(_06856_),
    .B1(net138));
 sg13g2_a22oi_1 _14784_ (.Y(_00585_),
    .B1(_06855_),
    .B2(_06856_),
    .A2(_06853_),
    .A1(net111));
 sg13g2_buf_1 _14785_ (.A(_01686_),
    .X(_06857_));
 sg13g2_buf_1 _14786_ (.A(\clock_inst.sec_tile.e[28] ),
    .X(_06858_));
 sg13g2_nand2b_1 _14787_ (.Y(_06859_),
    .B(_05139_),
    .A_N(net554));
 sg13g2_nor2_1 _14788_ (.A(_06842_),
    .B(_06859_),
    .Y(_06860_));
 sg13g2_nand3_1 _14789_ (.B(net554),
    .C(_06842_),
    .A(_06544_),
    .Y(_06861_));
 sg13g2_nor2_1 _14790_ (.A(_06838_),
    .B(_06861_),
    .Y(_06862_));
 sg13g2_a21oi_1 _14791_ (.A1(_06838_),
    .A2(_06860_),
    .Y(_06863_),
    .B1(_06862_));
 sg13g2_nor2_1 _14792_ (.A(_04793_),
    .B(_06863_),
    .Y(_06864_));
 sg13g2_xnor2_1 _14793_ (.Y(_06865_),
    .A(_06858_),
    .B(_06864_));
 sg13g2_a21oi_1 _14794_ (.A1(net53),
    .A2(_06865_),
    .Y(_00586_),
    .B1(_06357_));
 sg13g2_buf_1 _14795_ (.A(\clock_inst.sec_tile.e[29] ),
    .X(_06866_));
 sg13g2_o21ai_1 _14796_ (.B1(net457),
    .Y(_06867_),
    .A1(net554),
    .A2(_06848_));
 sg13g2_o21ai_1 _14797_ (.B1(net523),
    .Y(_06868_),
    .A1(_06842_),
    .A2(_06858_));
 sg13g2_and4_1 _14798_ (.A(net555),
    .B(net554),
    .C(_06815_),
    .D(_06833_),
    .X(_06869_));
 sg13g2_nand3_1 _14799_ (.B(_06858_),
    .C(_06869_),
    .A(_06842_),
    .Y(_06870_));
 sg13g2_nand3_1 _14800_ (.B(_06868_),
    .C(_06870_),
    .A(_06867_),
    .Y(_06871_));
 sg13g2_xnor2_1 _14801_ (.Y(_06872_),
    .A(net372),
    .B(_06871_));
 sg13g2_nor2_1 _14802_ (.A(net405),
    .B(_06872_),
    .Y(_06873_));
 sg13g2_xnor2_1 _14803_ (.Y(_06874_),
    .A(_06866_),
    .B(_06873_));
 sg13g2_a21oi_1 _14804_ (.A1(net53),
    .A2(_06874_),
    .Y(_00587_),
    .B1(_06369_));
 sg13g2_buf_1 _14805_ (.A(net502),
    .X(_06875_));
 sg13g2_xnor2_1 _14806_ (.Y(_06876_),
    .A(_05113_),
    .B(_06695_));
 sg13g2_nor2_1 _14807_ (.A(net366),
    .B(_06876_),
    .Y(_06877_));
 sg13g2_xnor2_1 _14808_ (.Y(_06878_),
    .A(\clock_inst.sec_tile.e[2] ),
    .B(_06877_));
 sg13g2_a21oi_1 _14809_ (.A1(net53),
    .A2(_06878_),
    .Y(_00588_),
    .B1(_06376_));
 sg13g2_nand2_1 _14810_ (.Y(_06879_),
    .A(_05864_),
    .B(_01610_));
 sg13g2_buf_1 _14811_ (.A(_06879_),
    .X(_06880_));
 sg13g2_or3_1 _14812_ (.A(_06842_),
    .B(_06858_),
    .C(_06866_),
    .X(_06881_));
 sg13g2_buf_1 _14813_ (.A(_06881_),
    .X(_06882_));
 sg13g2_nor2_1 _14814_ (.A(_06859_),
    .B(_06882_),
    .Y(_06883_));
 sg13g2_nand2_1 _14815_ (.Y(_06884_),
    .A(_06858_),
    .B(_06866_));
 sg13g2_nor2_1 _14816_ (.A(_06861_),
    .B(_06884_),
    .Y(_06885_));
 sg13g2_nor2_1 _14817_ (.A(_06883_),
    .B(_06885_),
    .Y(_06886_));
 sg13g2_o21ai_1 _14818_ (.B1(net457),
    .Y(_06887_),
    .A1(net554),
    .A2(_06882_));
 sg13g2_o21ai_1 _14819_ (.B1(_06887_),
    .Y(_06888_),
    .A1(_06838_),
    .A2(_06886_));
 sg13g2_xnor2_1 _14820_ (.Y(_06889_),
    .A(_05142_),
    .B(_06888_));
 sg13g2_nand2_1 _14821_ (.Y(_06890_),
    .A(_06880_),
    .B(_06889_));
 sg13g2_buf_1 _14822_ (.A(\clock_inst.sec_tile.e[30] ),
    .X(_06891_));
 sg13g2_a21oi_1 _14823_ (.A1(net80),
    .A2(_06890_),
    .Y(_06892_),
    .B1(_06891_));
 sg13g2_nand2_1 _14824_ (.Y(_06893_),
    .A(_06891_),
    .B(net445));
 sg13g2_o21ai_1 _14825_ (.B1(net242),
    .Y(_06894_),
    .A1(_06889_),
    .A2(_06893_));
 sg13g2_and2_1 _14826_ (.A(_06880_),
    .B(_06894_),
    .X(_06895_));
 sg13g2_o21ai_1 _14827_ (.B1(_06386_),
    .Y(_00589_),
    .A1(_06892_),
    .A2(_06895_));
 sg13g2_buf_1 _14828_ (.A(\clock_inst.sec_tile.e[31] ),
    .X(_06896_));
 sg13g2_inv_1 _14829_ (.Y(_06897_),
    .A(_06896_));
 sg13g2_nor2_1 _14830_ (.A(net242),
    .B(net235),
    .Y(_06898_));
 sg13g2_nor4_1 _14831_ (.A(_06831_),
    .B(_06891_),
    .C(_06848_),
    .D(_06882_),
    .Y(_06899_));
 sg13g2_nand2b_1 _14832_ (.Y(_06900_),
    .B(_05140_),
    .A_N(_06891_));
 sg13g2_nor2b_1 _14833_ (.A(_05139_),
    .B_N(_06891_),
    .Y(_06901_));
 sg13g2_nand4_1 _14834_ (.B(_06858_),
    .C(_06866_),
    .A(_06842_),
    .Y(_06902_),
    .D(_06901_));
 sg13g2_o21ai_1 _14835_ (.B1(_06902_),
    .Y(_06903_),
    .A1(_06882_),
    .A2(_06900_));
 sg13g2_o21ai_1 _14836_ (.B1(_06903_),
    .Y(_06904_),
    .A1(_06831_),
    .A2(_06848_));
 sg13g2_nor3_1 _14837_ (.A(net457),
    .B(_06850_),
    .C(_06904_),
    .Y(_06905_));
 sg13g2_a21oi_1 _14838_ (.A1(_05142_),
    .A2(_06899_),
    .Y(_06906_),
    .B1(_06905_));
 sg13g2_nor3_1 _14839_ (.A(_06897_),
    .B(net501),
    .C(_06906_),
    .Y(_06907_));
 sg13g2_a21oi_1 _14840_ (.A1(_06897_),
    .A2(_06906_),
    .Y(_06908_),
    .B1(_06907_));
 sg13g2_a22oi_1 _14841_ (.Y(_06909_),
    .B1(_06908_),
    .B2(net136),
    .A2(_06898_),
    .A1(_05864_));
 sg13g2_nand2b_1 _14842_ (.Y(_06910_),
    .B(net23),
    .A_N(_06405_));
 sg13g2_a22oi_1 _14843_ (.Y(_00590_),
    .B1(_06909_),
    .B2(_06910_),
    .A2(net137),
    .A1(_06897_));
 sg13g2_nor2_1 _14844_ (.A(_06891_),
    .B(_06896_),
    .Y(_06911_));
 sg13g2_nand3_1 _14845_ (.B(_06883_),
    .C(_06911_),
    .A(_06835_),
    .Y(_06912_));
 sg13g2_nand2_1 _14846_ (.Y(_06913_),
    .A(_06896_),
    .B(_06901_));
 sg13g2_and2_1 _14847_ (.A(_06544_),
    .B(_06833_),
    .X(_06914_));
 sg13g2_a21oi_1 _14848_ (.A1(_05141_),
    .A2(_06835_),
    .Y(_06915_),
    .B1(_06914_));
 sg13g2_nor3_1 _14849_ (.A(_06819_),
    .B(_06886_),
    .C(_06915_),
    .Y(_06916_));
 sg13g2_mux2_1 _14850_ (.A0(_06912_),
    .A1(_06913_),
    .S(_06916_),
    .X(_06917_));
 sg13g2_nand2_1 _14851_ (.Y(_06918_),
    .A(_06880_),
    .B(_06917_));
 sg13g2_buf_1 _14852_ (.A(\clock_inst.sec_tile.e[32] ),
    .X(_06919_));
 sg13g2_a21oi_1 _14853_ (.A1(_01678_),
    .A2(_06918_),
    .Y(_06920_),
    .B1(_06919_));
 sg13g2_nand3b_1 _14854_ (.B(net357),
    .C(_06919_),
    .Y(_06921_),
    .A_N(_06917_));
 sg13g2_a21oi_1 _14855_ (.A1(net161),
    .A2(_06921_),
    .Y(_06922_),
    .B1(_06379_));
 sg13g2_o21ai_1 _14856_ (.B1(_06415_),
    .Y(_00591_),
    .A1(_06920_),
    .A2(_06922_));
 sg13g2_buf_1 _14857_ (.A(\clock_inst.sec_tile.e[33] ),
    .X(_06923_));
 sg13g2_inv_1 _14858_ (.Y(_06924_),
    .A(_06923_));
 sg13g2_nand3b_1 _14859_ (.B(_06911_),
    .C(_05140_),
    .Y(_06925_),
    .A_N(_06919_));
 sg13g2_or2_1 _14860_ (.X(_06926_),
    .B(_06925_),
    .A(_06866_));
 sg13g2_nand4_1 _14861_ (.B(_06896_),
    .C(_06919_),
    .A(_06866_),
    .Y(_06927_),
    .D(_06901_));
 sg13g2_mux2_1 _14862_ (.A0(_06926_),
    .A1(_06927_),
    .S(_06871_),
    .X(_06928_));
 sg13g2_a21o_1 _14863_ (.A2(_06928_),
    .A1(_06422_),
    .B1(net137),
    .X(_06929_));
 sg13g2_nand2_1 _14864_ (.Y(_06930_),
    .A(_06923_),
    .B(net442));
 sg13g2_o21ai_1 _14865_ (.B1(_01063_),
    .Y(_06931_),
    .A1(_06928_),
    .A2(_06930_));
 sg13g2_and2_1 _14866_ (.A(_06422_),
    .B(_06931_),
    .X(_06932_));
 sg13g2_a21oi_1 _14867_ (.A1(_06924_),
    .A2(_06929_),
    .Y(_00592_),
    .B1(_06932_));
 sg13g2_nand2_1 _14868_ (.Y(_06933_),
    .A(net236),
    .B(_06880_));
 sg13g2_buf_1 _14869_ (.A(\clock_inst.sec_tile.e[34] ),
    .X(_06934_));
 sg13g2_nand3_1 _14870_ (.B(net442),
    .C(_06880_),
    .A(_06934_),
    .Y(_06935_));
 sg13g2_nand2b_1 _14871_ (.Y(_06936_),
    .B(_06880_),
    .A_N(_06934_));
 sg13g2_or2_1 _14872_ (.X(_06937_),
    .B(_06925_),
    .A(_06923_));
 sg13g2_nand4_1 _14873_ (.B(_06919_),
    .C(_06923_),
    .A(_06896_),
    .Y(_06938_),
    .D(_06901_));
 sg13g2_mux2_1 _14874_ (.A0(_06937_),
    .A1(_06938_),
    .S(_06888_),
    .X(_06939_));
 sg13g2_mux2_1 _14875_ (.A0(_06935_),
    .A1(_06936_),
    .S(_06939_),
    .X(_06940_));
 sg13g2_nand2b_1 _14876_ (.Y(_06941_),
    .B(_02072_),
    .A_N(_06934_));
 sg13g2_nand3_1 _14877_ (.B(_06940_),
    .C(_06941_),
    .A(_06933_),
    .Y(_06942_));
 sg13g2_o21ai_1 _14878_ (.B1(_06942_),
    .Y(_00593_),
    .A1(net44),
    .A2(_06433_));
 sg13g2_nor3_1 _14879_ (.A(_06934_),
    .B(_06882_),
    .C(_06937_),
    .Y(_06943_));
 sg13g2_nand4_1 _14880_ (.B(_06919_),
    .C(_06923_),
    .A(_06896_),
    .Y(_06944_),
    .D(_06934_));
 sg13g2_nor4_1 _14881_ (.A(net457),
    .B(_06850_),
    .C(_06904_),
    .D(_06944_),
    .Y(_06945_));
 sg13g2_a21oi_1 _14882_ (.A1(_06904_),
    .A2(_06943_),
    .Y(_06946_),
    .B1(_06945_));
 sg13g2_a21oi_1 _14883_ (.A1(_06880_),
    .A2(_06946_),
    .Y(_06947_),
    .B1(_02072_));
 sg13g2_nor2_1 _14884_ (.A(\clock_inst.sec_tile.e[35] ),
    .B(_06947_),
    .Y(_06948_));
 sg13g2_nand3b_1 _14885_ (.B(net357),
    .C(\clock_inst.sec_tile.e[35] ),
    .Y(_06949_),
    .A_N(_06946_));
 sg13g2_a21oi_1 _14886_ (.A1(net161),
    .A2(_06949_),
    .Y(_06950_),
    .B1(_06379_));
 sg13g2_o21ai_1 _14887_ (.B1(_06442_),
    .Y(_00594_),
    .A1(_06948_),
    .A2(_06950_));
 sg13g2_nand2_1 _14888_ (.Y(_06951_),
    .A(\clock_inst.sec_a[36] ),
    .B(net355));
 sg13g2_xor2_1 _14889_ (.B(_06951_),
    .A(\clock_inst.sec_tile.e[36] ),
    .X(_06952_));
 sg13g2_o21ai_1 _14890_ (.B1(_06448_),
    .Y(_00595_),
    .A1(net135),
    .A2(_06952_));
 sg13g2_nand2_1 _14891_ (.Y(_06953_),
    .A(\clock_inst.sec_a[36] ),
    .B(\clock_inst.sec_tile.e[36] ));
 sg13g2_xnor2_1 _14892_ (.Y(_06954_),
    .A(_05178_),
    .B(_06953_));
 sg13g2_nor2_1 _14893_ (.A(net366),
    .B(_06954_),
    .Y(_06955_));
 sg13g2_xnor2_1 _14894_ (.Y(_06956_),
    .A(\clock_inst.sec_tile.e[37] ),
    .B(_06955_));
 sg13g2_a21oi_1 _14895_ (.A1(net53),
    .A2(_06956_),
    .Y(_00596_),
    .B1(_06456_));
 sg13g2_nor2_1 _14896_ (.A(\clock_inst.sec_a[37] ),
    .B(\clock_inst.sec_tile.e[37] ),
    .Y(_06957_));
 sg13g2_a22oi_1 _14897_ (.Y(_06958_),
    .B1(\clock_inst.sec_a[37] ),
    .B2(\clock_inst.sec_tile.e[37] ),
    .A2(\clock_inst.sec_tile.e[36] ),
    .A1(\clock_inst.sec_a[36] ));
 sg13g2_nor2_1 _14898_ (.A(_06957_),
    .B(_06958_),
    .Y(_06959_));
 sg13g2_xnor2_1 _14899_ (.Y(_06960_),
    .A(_05197_),
    .B(_06959_));
 sg13g2_nor2_1 _14900_ (.A(net366),
    .B(_06960_),
    .Y(_06961_));
 sg13g2_xnor2_1 _14901_ (.Y(_06962_),
    .A(\clock_inst.sec_tile.e[38] ),
    .B(_06961_));
 sg13g2_a21oi_1 _14902_ (.A1(net53),
    .A2(_06962_),
    .Y(_00597_),
    .B1(_06466_));
 sg13g2_buf_2 _14903_ (.A(\clock_inst.sec_tile.e[39] ),
    .X(_06963_));
 sg13g2_nor2_1 _14904_ (.A(_05197_),
    .B(\clock_inst.sec_tile.e[38] ),
    .Y(_06964_));
 sg13g2_or3_1 _14905_ (.A(_06957_),
    .B(_06958_),
    .C(_06964_),
    .X(_06965_));
 sg13g2_buf_1 _14906_ (.A(_06965_),
    .X(_06966_));
 sg13g2_nand2_1 _14907_ (.Y(_06967_),
    .A(_05197_),
    .B(\clock_inst.sec_tile.e[38] ));
 sg13g2_nand2_1 _14908_ (.Y(_06968_),
    .A(_06966_),
    .B(_06967_));
 sg13g2_xnor2_1 _14909_ (.Y(_06969_),
    .A(_05221_),
    .B(_06968_));
 sg13g2_nor2_1 _14910_ (.A(net366),
    .B(_06969_),
    .Y(_06970_));
 sg13g2_xnor2_1 _14911_ (.Y(_06971_),
    .A(_06963_),
    .B(_06970_));
 sg13g2_a21oi_1 _14912_ (.A1(net53),
    .A2(_06971_),
    .Y(_00598_),
    .B1(_06478_));
 sg13g2_a21oi_1 _14913_ (.A1(_06695_),
    .A2(_06696_),
    .Y(_06972_),
    .B1(_06697_));
 sg13g2_xnor2_1 _14914_ (.Y(_06973_),
    .A(_06686_),
    .B(_06972_));
 sg13g2_nor2_1 _14915_ (.A(net366),
    .B(_06973_),
    .Y(_06974_));
 sg13g2_xnor2_1 _14916_ (.Y(_06975_),
    .A(\clock_inst.sec_tile.e[3] ),
    .B(_06974_));
 sg13g2_a21oi_1 _14917_ (.A1(net53),
    .A2(_06975_),
    .Y(_00599_),
    .B1(_06485_));
 sg13g2_buf_2 _14918_ (.A(\clock_inst.sec_tile.e[40] ),
    .X(_06976_));
 sg13g2_a21o_1 _14919_ (.A2(_06968_),
    .A1(_06963_),
    .B1(_05221_),
    .X(_06977_));
 sg13g2_o21ai_1 _14920_ (.B1(_06977_),
    .Y(_06978_),
    .A1(_06963_),
    .A2(_06968_));
 sg13g2_xor2_1 _14921_ (.B(_06978_),
    .A(_05267_),
    .X(_06979_));
 sg13g2_nor2_1 _14922_ (.A(net366),
    .B(_06979_),
    .Y(_06980_));
 sg13g2_xnor2_1 _14923_ (.Y(_06981_),
    .A(_06976_),
    .B(_06980_));
 sg13g2_a21oi_1 _14924_ (.A1(net53),
    .A2(_06981_),
    .Y(_00600_),
    .B1(_06495_));
 sg13g2_buf_1 _14925_ (.A(\clock_inst.sec_tile.e[41] ),
    .X(_06982_));
 sg13g2_inv_1 _14926_ (.Y(_06983_),
    .A(_06982_));
 sg13g2_a22oi_1 _14927_ (.Y(_06984_),
    .B1(_05267_),
    .B2(_06976_),
    .A2(_06963_),
    .A1(_05221_));
 sg13g2_and2_1 _14928_ (.A(_06967_),
    .B(_06984_),
    .X(_06985_));
 sg13g2_nand2_1 _14929_ (.Y(_06986_),
    .A(_05267_),
    .B(_06976_));
 sg13g2_nor2_1 _14930_ (.A(_05221_),
    .B(_06963_),
    .Y(_06987_));
 sg13g2_nor2_1 _14931_ (.A(_05267_),
    .B(_06976_),
    .Y(_06988_));
 sg13g2_a21o_1 _14932_ (.A2(_06987_),
    .A1(_06986_),
    .B1(_06988_),
    .X(_06989_));
 sg13g2_a21o_1 _14933_ (.A2(_06985_),
    .A1(_06966_),
    .B1(_06989_),
    .X(_06990_));
 sg13g2_buf_1 _14934_ (.A(_06990_),
    .X(_06991_));
 sg13g2_xnor2_1 _14935_ (.Y(_06992_),
    .A(_05286_),
    .B(_06991_));
 sg13g2_nor2_1 _14936_ (.A(net501),
    .B(_06992_),
    .Y(_06993_));
 sg13g2_xnor2_1 _14937_ (.Y(_06994_),
    .A(_06983_),
    .B(_06993_));
 sg13g2_nor2_1 _14938_ (.A(net144),
    .B(_06994_),
    .Y(_06995_));
 sg13g2_a21oi_1 _14939_ (.A1(net88),
    .A2(_06502_),
    .Y(_00601_),
    .B1(_06995_));
 sg13g2_buf_1 _14940_ (.A(\clock_inst.sec_tile.e[42] ),
    .X(_06996_));
 sg13g2_inv_1 _14941_ (.Y(_06997_),
    .A(_06996_));
 sg13g2_inv_1 _14942_ (.Y(_06998_),
    .A(_05316_));
 sg13g2_a21oi_1 _14943_ (.A1(_06966_),
    .A2(_06985_),
    .Y(_06999_),
    .B1(_06989_));
 sg13g2_o21ai_1 _14944_ (.B1(\clock_inst.sec_a[41] ),
    .Y(_07000_),
    .A1(_06982_),
    .A2(_06999_));
 sg13g2_o21ai_1 _14945_ (.B1(_07000_),
    .Y(_07001_),
    .A1(_06983_),
    .A2(_06991_));
 sg13g2_xnor2_1 _14946_ (.Y(_07002_),
    .A(_06998_),
    .B(_07001_));
 sg13g2_nand2_1 _14947_ (.Y(_07003_),
    .A(net357),
    .B(_07002_));
 sg13g2_xnor2_1 _14948_ (.Y(_07004_),
    .A(_06997_),
    .B(_07003_));
 sg13g2_o21ai_1 _14949_ (.B1(_06516_),
    .Y(_00602_),
    .A1(net146),
    .A2(_07004_));
 sg13g2_buf_1 _14950_ (.A(\clock_inst.sec_tile.e[43] ),
    .X(_07005_));
 sg13g2_a221oi_1 _14951_ (.B2(_06997_),
    .C1(_06991_),
    .B1(_06998_),
    .A1(_05286_),
    .Y(_07006_),
    .A2(_06983_));
 sg13g2_nor2_1 _14952_ (.A(_05286_),
    .B(_06983_),
    .Y(_07007_));
 sg13g2_o21ai_1 _14953_ (.B1(_07007_),
    .Y(_07008_),
    .A1(_05316_),
    .A2(_06996_));
 sg13g2_o21ai_1 _14954_ (.B1(_07008_),
    .Y(_07009_),
    .A1(_06998_),
    .A2(_06997_));
 sg13g2_or2_1 _14955_ (.X(_07010_),
    .B(_07009_),
    .A(_07006_));
 sg13g2_buf_1 _14956_ (.A(_07010_),
    .X(_07011_));
 sg13g2_xnor2_1 _14957_ (.Y(_07012_),
    .A(_05318_),
    .B(_07011_));
 sg13g2_nand2_1 _14958_ (.Y(_07013_),
    .A(net443),
    .B(_07012_));
 sg13g2_xnor2_1 _14959_ (.Y(_07014_),
    .A(net553),
    .B(_07013_));
 sg13g2_nor2_1 _14960_ (.A(net144),
    .B(_07014_),
    .Y(_07015_));
 sg13g2_a21oi_1 _14961_ (.A1(net88),
    .A2(_06534_),
    .Y(_00603_),
    .B1(_07015_));
 sg13g2_buf_1 _14962_ (.A(\clock_inst.sec_tile.e[44] ),
    .X(_07016_));
 sg13g2_buf_1 _14963_ (.A(_07016_),
    .X(_07017_));
 sg13g2_nor3_1 _14964_ (.A(net553),
    .B(_07006_),
    .C(_07009_),
    .Y(_07018_));
 sg13g2_o21ai_1 _14965_ (.B1(net553),
    .Y(_07019_),
    .A1(_07006_),
    .A2(_07009_));
 sg13g2_o21ai_1 _14966_ (.B1(_07019_),
    .Y(_07020_),
    .A1(_05318_),
    .A2(_07018_));
 sg13g2_buf_2 _14967_ (.A(_07020_),
    .X(_07021_));
 sg13g2_buf_8 _14968_ (.A(_07021_),
    .X(_07022_));
 sg13g2_xnor2_1 _14969_ (.Y(_07023_),
    .A(net558),
    .B(net21));
 sg13g2_nor2_1 _14970_ (.A(_06875_),
    .B(_07023_),
    .Y(_07024_));
 sg13g2_xnor2_1 _14971_ (.Y(_07025_),
    .A(net519),
    .B(_07024_));
 sg13g2_a21oi_1 _14972_ (.A1(_06857_),
    .A2(_07025_),
    .Y(_00604_),
    .B1(_06552_));
 sg13g2_buf_2 _14973_ (.A(\clock_inst.sec_tile.e[45] ),
    .X(_07026_));
 sg13g2_nor2_1 _14974_ (.A(_05356_),
    .B(_07016_),
    .Y(_07027_));
 sg13g2_nor2b_1 _14975_ (.A(net558),
    .B_N(_07016_),
    .Y(_07028_));
 sg13g2_mux2_1 _14976_ (.A0(_07027_),
    .A1(_07028_),
    .S(net21),
    .X(_07029_));
 sg13g2_nand2_1 _14977_ (.Y(_07030_),
    .A(net355),
    .B(_07029_));
 sg13g2_xor2_1 _14978_ (.B(_07030_),
    .A(_07026_),
    .X(_07031_));
 sg13g2_xnor2_1 _14979_ (.Y(_07032_),
    .A(_06558_),
    .B(_06554_));
 sg13g2_nand2_1 _14980_ (.Y(_07033_),
    .A(net45),
    .B(_07032_));
 sg13g2_a21oi_1 _14981_ (.A1(\clock_inst.sec_c[45] ),
    .A2(net43),
    .Y(_07034_),
    .B1(net138));
 sg13g2_a22oi_1 _14982_ (.Y(_00605_),
    .B1(_07033_),
    .B2(_07034_),
    .A2(_07031_),
    .A1(net111));
 sg13g2_buf_1 _14983_ (.A(\clock_inst.sec_tile.e[46] ),
    .X(_07035_));
 sg13g2_nand3_1 _14984_ (.B(net21),
    .C(_07028_),
    .A(_07026_),
    .Y(_07036_));
 sg13g2_or4_1 _14985_ (.A(_05356_),
    .B(net519),
    .C(_07026_),
    .D(net21),
    .X(_07037_));
 sg13g2_a21oi_1 _14986_ (.A1(_07036_),
    .A2(_07037_),
    .Y(_07038_),
    .B1(net448));
 sg13g2_xnor2_1 _14987_ (.Y(_07039_),
    .A(_07035_),
    .B(_07038_));
 sg13g2_a22oi_1 _14988_ (.Y(_00606_),
    .B1(_07039_),
    .B2(net79),
    .A2(_06566_),
    .A1(_06565_));
 sg13g2_nor2_1 _14989_ (.A(_07026_),
    .B(_07035_),
    .Y(_07040_));
 sg13g2_and2_1 _14990_ (.A(_07026_),
    .B(_07035_),
    .X(_07041_));
 sg13g2_a22oi_1 _14991_ (.Y(_07042_),
    .B1(_07041_),
    .B2(_07028_),
    .A2(_07040_),
    .A1(_07027_));
 sg13g2_xnor2_1 _14992_ (.Y(_07043_),
    .A(\clock_inst.sec_a[43] ),
    .B(net553));
 sg13g2_nor2_1 _14993_ (.A(_07042_),
    .B(_07043_),
    .Y(_07044_));
 sg13g2_nand2_1 _14994_ (.Y(_07045_),
    .A(net519),
    .B(_07041_));
 sg13g2_nand2b_1 _14995_ (.Y(_07046_),
    .B(_07040_),
    .A_N(net519));
 sg13g2_a22oi_1 _14996_ (.Y(_07047_),
    .B1(net558),
    .B2(_07046_),
    .A2(net553),
    .A1(\clock_inst.sec_a[43] ));
 sg13g2_a21oi_1 _14997_ (.A1(_05356_),
    .A2(_07045_),
    .Y(_07048_),
    .B1(_07047_));
 sg13g2_a21o_1 _14998_ (.A2(_07044_),
    .A1(_07011_),
    .B1(_07048_),
    .X(_07049_));
 sg13g2_xnor2_1 _14999_ (.Y(_07050_),
    .A(net558),
    .B(_07049_));
 sg13g2_nor2_1 _15000_ (.A(net446),
    .B(_07050_),
    .Y(_07051_));
 sg13g2_xnor2_1 _15001_ (.Y(_07052_),
    .A(\clock_inst.sec_tile.e[47] ),
    .B(_07051_));
 sg13g2_xnor2_1 _15002_ (.Y(_07053_),
    .A(_06567_),
    .B(_06572_));
 sg13g2_o21ai_1 _15003_ (.B1(net233),
    .Y(_07054_),
    .A1(\clock_inst.sec_c[47] ),
    .A2(net101));
 sg13g2_a21o_1 _15004_ (.A2(_07053_),
    .A1(net50),
    .B1(_07054_),
    .X(_07055_));
 sg13g2_o21ai_1 _15005_ (.B1(_07055_),
    .Y(_00607_),
    .A1(net146),
    .A2(_07052_));
 sg13g2_buf_1 _15006_ (.A(\clock_inst.sec_tile.e[48] ),
    .X(_07056_));
 sg13g2_nor2_1 _15007_ (.A(_05356_),
    .B(\clock_inst.sec_tile.e[47] ),
    .Y(_07057_));
 sg13g2_nand2_1 _15008_ (.Y(_07058_),
    .A(_07040_),
    .B(_07057_));
 sg13g2_nor2_1 _15009_ (.A(net519),
    .B(_07058_),
    .Y(_07059_));
 sg13g2_nor2b_1 _15010_ (.A(net558),
    .B_N(\clock_inst.sec_tile.e[47] ),
    .Y(_07060_));
 sg13g2_nor2b_1 _15011_ (.A(_07045_),
    .B_N(_07060_),
    .Y(_07061_));
 sg13g2_mux2_1 _15012_ (.A0(_07059_),
    .A1(_07061_),
    .S(net21),
    .X(_07062_));
 sg13g2_nand2_1 _15013_ (.Y(_07063_),
    .A(net357),
    .B(_07062_));
 sg13g2_xor2_1 _15014_ (.B(_07063_),
    .A(_07056_),
    .X(_07064_));
 sg13g2_a22oi_1 _15015_ (.Y(_00608_),
    .B1(_07064_),
    .B2(net79),
    .A2(_06586_),
    .A1(_06585_));
 sg13g2_buf_2 _15016_ (.A(\clock_inst.sec_tile.e[49] ),
    .X(_07065_));
 sg13g2_or2_1 _15017_ (.X(_07066_),
    .B(_07058_),
    .A(_07056_));
 sg13g2_buf_1 _15018_ (.A(_07066_),
    .X(_07067_));
 sg13g2_nor2_1 _15019_ (.A(net519),
    .B(_07067_),
    .Y(_07068_));
 sg13g2_and2_1 _15020_ (.A(_07056_),
    .B(_07061_),
    .X(_07069_));
 sg13g2_mux2_1 _15021_ (.A0(_07068_),
    .A1(_07069_),
    .S(_07021_),
    .X(_07070_));
 sg13g2_nand3_1 _15022_ (.B(net357),
    .C(_07070_),
    .A(_07065_),
    .Y(_07071_));
 sg13g2_a221oi_1 _15023_ (.B2(net153),
    .C1(_06597_),
    .B1(_07071_),
    .A1(\clock_inst.sec_c[49] ),
    .Y(_07072_),
    .A2(net82));
 sg13g2_a21oi_1 _15024_ (.A1(\clock_inst.sec_c[49] ),
    .A2(_01610_),
    .Y(_07073_),
    .B1(_07065_));
 sg13g2_nand2b_1 _15025_ (.Y(_07074_),
    .B(_07073_),
    .A_N(_07070_));
 sg13g2_inv_1 _15026_ (.Y(_07075_),
    .A(_07065_));
 sg13g2_nand2_1 _15027_ (.Y(_07076_),
    .A(_07075_),
    .B(net137));
 sg13g2_o21ai_1 _15028_ (.B1(_07076_),
    .Y(_07077_),
    .A1(_06597_),
    .A2(_07074_));
 sg13g2_nor2_1 _15029_ (.A(_07072_),
    .B(_07077_),
    .Y(_00609_));
 sg13g2_xnor2_1 _15030_ (.Y(_07078_),
    .A(_06144_),
    .B(_06601_));
 sg13g2_nand2_1 _15031_ (.Y(_07079_),
    .A(net87),
    .B(_07078_));
 sg13g2_o21ai_1 _15032_ (.B1(_07079_),
    .Y(_07080_),
    .A1(\clock_inst.sec_c[4] ),
    .A2(net50));
 sg13g2_a21oi_1 _15033_ (.A1(_06686_),
    .A2(_06687_),
    .Y(_07081_),
    .B1(_06698_));
 sg13g2_xnor2_1 _15034_ (.Y(_07082_),
    .A(_05337_),
    .B(_07081_));
 sg13g2_nand2_1 _15035_ (.Y(_07083_),
    .A(net443),
    .B(_07082_));
 sg13g2_xnor2_1 _15036_ (.Y(_07084_),
    .A(_06689_),
    .B(_07083_));
 sg13g2_nor2_1 _15037_ (.A(net144),
    .B(_07084_),
    .Y(_07085_));
 sg13g2_a21oi_1 _15038_ (.A1(net88),
    .A2(_07080_),
    .Y(_00610_),
    .B1(_07085_));
 sg13g2_inv_1 _15039_ (.Y(_07086_),
    .A(\clock_inst.sec_tile.e[50] ));
 sg13g2_and3_1 _15040_ (.X(_07087_),
    .A(_07035_),
    .B(_07056_),
    .C(_07065_));
 sg13g2_nor3_1 _15041_ (.A(_07035_),
    .B(_07056_),
    .C(_07065_),
    .Y(_07088_));
 sg13g2_a22oi_1 _15042_ (.Y(_07089_),
    .B1(_07088_),
    .B2(_07057_),
    .A2(_07087_),
    .A1(_07060_));
 sg13g2_nor2b_1 _15043_ (.A(_07089_),
    .B_N(net519),
    .Y(_07090_));
 sg13g2_nand3_1 _15044_ (.B(_07086_),
    .C(_07090_),
    .A(_07026_),
    .Y(_07091_));
 sg13g2_mux2_1 _15045_ (.A0(_07086_),
    .A1(_07091_),
    .S(_07021_),
    .X(_07092_));
 sg13g2_or4_1 _15046_ (.A(_07017_),
    .B(_07065_),
    .C(\clock_inst.sec_tile.e[50] ),
    .D(_07067_),
    .X(_07093_));
 sg13g2_or2_1 _15047_ (.X(_07094_),
    .B(_07093_),
    .A(net21));
 sg13g2_o21ai_1 _15048_ (.B1(_07094_),
    .Y(_07095_),
    .A1(_05355_),
    .A2(_07092_));
 sg13g2_and3_1 _15049_ (.X(_07096_),
    .A(_05356_),
    .B(_07026_),
    .C(_07090_));
 sg13g2_nor4_1 _15050_ (.A(_07065_),
    .B(net21),
    .C(_07067_),
    .D(_07090_),
    .Y(_07097_));
 sg13g2_o21ai_1 _15051_ (.B1(net356),
    .Y(_07098_),
    .A1(_07096_),
    .A2(_07097_));
 sg13g2_a221oi_1 _15052_ (.B2(\clock_inst.sec_tile.e[50] ),
    .C1(net155),
    .B1(_07098_),
    .A1(net356),
    .Y(_07099_),
    .A2(_07095_));
 sg13g2_a21oi_1 _15053_ (.A1(_06610_),
    .A2(_06611_),
    .Y(_00611_),
    .B1(_07099_));
 sg13g2_buf_1 _15054_ (.A(\clock_inst.sec_tile.e[51] ),
    .X(_07100_));
 sg13g2_nor2_1 _15055_ (.A(_07075_),
    .B(_07086_),
    .Y(_07101_));
 sg13g2_and2_1 _15056_ (.A(_07056_),
    .B(_07101_),
    .X(_07102_));
 sg13g2_nand3_1 _15057_ (.B(_07060_),
    .C(_07102_),
    .A(_07049_),
    .Y(_07103_));
 sg13g2_a21oi_1 _15058_ (.A1(_07094_),
    .A2(_07103_),
    .Y(_07104_),
    .B1(net447));
 sg13g2_xnor2_1 _15059_ (.Y(_07105_),
    .A(_07100_),
    .B(_07104_));
 sg13g2_xnor2_1 _15060_ (.Y(_07106_),
    .A(_06623_),
    .B(_06619_));
 sg13g2_nand2_1 _15061_ (.Y(_07107_),
    .A(net45),
    .B(_07106_));
 sg13g2_a21oi_1 _15062_ (.A1(\clock_inst.sec_c[51] ),
    .A2(net47),
    .Y(_07108_),
    .B1(net136));
 sg13g2_a22oi_1 _15063_ (.Y(_00612_),
    .B1(_07107_),
    .B2(_07108_),
    .A2(_07105_),
    .A1(net111));
 sg13g2_or2_1 _15064_ (.X(_07109_),
    .B(_07059_),
    .A(_07061_));
 sg13g2_nand4_1 _15065_ (.B(net21),
    .C(_07102_),
    .A(_07100_),
    .Y(_07110_),
    .D(_07109_));
 sg13g2_or2_1 _15066_ (.X(_07111_),
    .B(_07093_),
    .A(_07100_));
 sg13g2_a221oi_1 _15067_ (.B2(_07111_),
    .C1(net446),
    .B1(_07110_),
    .A1(_05355_),
    .Y(_07112_),
    .A2(_07022_));
 sg13g2_xnor2_1 _15068_ (.Y(_07113_),
    .A(\clock_inst.sec_tile.e[52] ),
    .B(_07112_));
 sg13g2_a21oi_1 _15069_ (.A1(_06857_),
    .A2(_07113_),
    .Y(_00613_),
    .B1(_06635_));
 sg13g2_inv_1 _15070_ (.Y(_07114_),
    .A(\clock_inst.sec_tile.e[53] ));
 sg13g2_nor2_1 _15071_ (.A(net558),
    .B(_07017_),
    .Y(_07115_));
 sg13g2_or2_1 _15072_ (.X(_07116_),
    .B(net553),
    .A(_06996_));
 sg13g2_a21oi_1 _15073_ (.A1(_06982_),
    .A2(_06999_),
    .Y(_07117_),
    .B1(_07116_));
 sg13g2_or2_1 _15074_ (.X(_07118_),
    .B(net553),
    .A(_05316_));
 sg13g2_a21oi_1 _15075_ (.A1(_06982_),
    .A2(_06999_),
    .Y(_07119_),
    .B1(_07118_));
 sg13g2_o21ai_1 _15076_ (.B1(_07000_),
    .Y(_07120_),
    .A1(_07117_),
    .A2(_07119_));
 sg13g2_nor3_1 _15077_ (.A(_05316_),
    .B(_06996_),
    .C(net553),
    .Y(_07121_));
 sg13g2_nor2_1 _15078_ (.A(_05318_),
    .B(_07121_),
    .Y(_07122_));
 sg13g2_and2_1 _15079_ (.A(net558),
    .B(net519),
    .X(_07123_));
 sg13g2_a221oi_1 _15080_ (.B2(_07122_),
    .C1(_07123_),
    .B1(_07120_),
    .A1(_07005_),
    .Y(_07124_),
    .A2(_07011_));
 sg13g2_or2_1 _15081_ (.X(_07125_),
    .B(\clock_inst.sec_tile.e[52] ),
    .A(_07100_));
 sg13g2_nor4_1 _15082_ (.A(_07065_),
    .B(\clock_inst.sec_tile.e[50] ),
    .C(_07067_),
    .D(_07125_),
    .Y(_07126_));
 sg13g2_o21ai_1 _15083_ (.B1(_07126_),
    .Y(_07127_),
    .A1(_07115_),
    .A2(_07124_));
 sg13g2_and2_1 _15084_ (.A(_07100_),
    .B(\clock_inst.sec_tile.e[52] ),
    .X(_07128_));
 sg13g2_nand4_1 _15085_ (.B(_07069_),
    .C(_07101_),
    .A(_07022_),
    .Y(_07129_),
    .D(_07128_));
 sg13g2_nand2_1 _15086_ (.Y(_07130_),
    .A(_07127_),
    .B(_07129_));
 sg13g2_o21ai_1 _15087_ (.B1(net80),
    .Y(_07131_),
    .A1(_06648_),
    .A2(_07130_));
 sg13g2_nand2_1 _15088_ (.Y(_07132_),
    .A(\clock_inst.sec_tile.e[53] ),
    .B(net442));
 sg13g2_a21o_1 _15089_ (.A2(_07129_),
    .A1(_07127_),
    .B1(_07132_),
    .X(_07133_));
 sg13g2_a21oi_1 _15090_ (.A1(net145),
    .A2(_07133_),
    .Y(_07134_),
    .B1(_06648_));
 sg13g2_a21oi_1 _15091_ (.A1(_07114_),
    .A2(_07131_),
    .Y(_00614_),
    .B1(_07134_));
 sg13g2_a21o_1 _15092_ (.A2(_07081_),
    .A1(_06689_),
    .B1(\clock_inst.sec_a[4] ),
    .X(_07135_));
 sg13g2_o21ai_1 _15093_ (.B1(_07135_),
    .Y(_07136_),
    .A1(_06689_),
    .A2(_07081_));
 sg13g2_xor2_1 _15094_ (.B(_07136_),
    .A(_05362_),
    .X(_07137_));
 sg13g2_nor2_1 _15095_ (.A(net366),
    .B(_07137_),
    .Y(_07138_));
 sg13g2_xnor2_1 _15096_ (.Y(_07139_),
    .A(_06688_),
    .B(_07138_));
 sg13g2_a21oi_1 _15097_ (.A1(net75),
    .A2(_07139_),
    .Y(_00615_),
    .B1(_06656_));
 sg13g2_nor2_1 _15098_ (.A(_06700_),
    .B(_06705_),
    .Y(_07140_));
 sg13g2_xnor2_1 _15099_ (.Y(_07141_),
    .A(_06711_),
    .B(_07140_));
 sg13g2_nor2_1 _15100_ (.A(net366),
    .B(_07141_),
    .Y(_07142_));
 sg13g2_xnor2_1 _15101_ (.Y(_07143_),
    .A(_06706_),
    .B(_07142_));
 sg13g2_a21oi_1 _15102_ (.A1(net75),
    .A2(_07143_),
    .Y(_00616_),
    .B1(_06662_));
 sg13g2_nor3_1 _15103_ (.A(_06706_),
    .B(_06700_),
    .C(_06705_),
    .Y(_07144_));
 sg13g2_o21ai_1 _15104_ (.B1(_06706_),
    .Y(_07145_),
    .A1(_06700_),
    .A2(_06705_));
 sg13g2_o21ai_1 _15105_ (.B1(_07145_),
    .Y(_07146_),
    .A1(_06711_),
    .A2(_07144_));
 sg13g2_xnor2_1 _15106_ (.Y(_07147_),
    .A(_05392_),
    .B(_07146_));
 sg13g2_nor2_1 _15107_ (.A(net446),
    .B(_07147_),
    .Y(_07148_));
 sg13g2_xnor2_1 _15108_ (.Y(_07149_),
    .A(\clock_inst.sec_tile.e[7] ),
    .B(_07148_));
 sg13g2_o21ai_1 _15109_ (.B1(_06671_),
    .Y(_00617_),
    .A1(net146),
    .A2(_07149_));
 sg13g2_xnor2_1 _15110_ (.Y(_07150_),
    .A(_04935_),
    .B(net25));
 sg13g2_nor2_1 _15111_ (.A(_06875_),
    .B(_07150_),
    .Y(_07151_));
 sg13g2_xnor2_1 _15112_ (.Y(_07152_),
    .A(\clock_inst.sec_tile.e[8] ),
    .B(_07151_));
 sg13g2_a21oi_1 _15113_ (.A1(net75),
    .A2(_07152_),
    .Y(_00618_),
    .B1(_06676_));
 sg13g2_or2_1 _15114_ (.X(_07153_),
    .B(_06720_),
    .A(net542));
 sg13g2_nand2_1 _15115_ (.Y(_07154_),
    .A(_01815_),
    .B(_06718_));
 sg13g2_mux2_1 _15116_ (.A0(_07153_),
    .A1(_07154_),
    .S(net25),
    .X(_07155_));
 sg13g2_xnor2_1 _15117_ (.Y(_07156_),
    .A(_06685_),
    .B(_07155_));
 sg13g2_nor2_1 _15118_ (.A(net144),
    .B(_07156_),
    .Y(_07157_));
 sg13g2_a21oi_1 _15119_ (.A1(net88),
    .A2(_06680_),
    .Y(_00619_),
    .B1(_07157_));
 sg13g2_buf_1 _15120_ (.A(\clock_inst.frameno[4] ),
    .X(_07158_));
 sg13g2_nand2b_1 _15121_ (.Y(_07159_),
    .B(\clock_inst.frameno[6] ),
    .A_N(_07158_));
 sg13g2_buf_1 _15122_ (.A(\clock_inst.frameno[5] ),
    .X(_07160_));
 sg13g2_buf_1 _15123_ (.A(\clock_inst.frameno[3] ),
    .X(_07161_));
 sg13g2_nand2b_1 _15124_ (.Y(_07162_),
    .B(_07161_),
    .A_N(_07160_));
 sg13g2_buf_1 _15125_ (.A(\clock_inst.frameno[1] ),
    .X(_07163_));
 sg13g2_buf_1 _15126_ (.A(\clock_inst.frameno[0] ),
    .X(_07164_));
 sg13g2_nand2_1 _15127_ (.Y(_07165_),
    .A(_07163_),
    .B(_07164_));
 sg13g2_nor4_1 _15128_ (.A(\clock_inst.frameno[2] ),
    .B(_07159_),
    .C(_07162_),
    .D(_07165_),
    .Y(_07166_));
 sg13g2_buf_2 _15129_ (.A(_07166_),
    .X(_07167_));
 sg13g2_buf_1 _15130_ (.A(rst_n),
    .X(_07168_));
 sg13g2_buf_1 _15131_ (.A(_07168_),
    .X(_07169_));
 sg13g2_nand2b_1 _15132_ (.Y(_07170_),
    .B(net552),
    .A_N(_07167_));
 sg13g2_buf_1 _15133_ (.A(_07170_),
    .X(_07171_));
 sg13g2_and2_1 _15134_ (.A(net549),
    .B(_00000_),
    .X(_07172_));
 sg13g2_a21oi_1 _15135_ (.A1(net450),
    .A2(_07164_),
    .Y(_07173_),
    .B1(_07172_));
 sg13g2_nor2_1 _15136_ (.A(_07171_),
    .B(_07173_),
    .Y(_00004_));
 sg13g2_nand2_1 _15137_ (.Y(_07174_),
    .A(net549),
    .B(_07164_));
 sg13g2_xor2_1 _15138_ (.B(_07174_),
    .A(_07163_),
    .X(_07175_));
 sg13g2_nor2_1 _15139_ (.A(_07171_),
    .B(_07175_),
    .Y(_00005_));
 sg13g2_inv_1 _15140_ (.Y(_07176_),
    .A(\clock_inst.frameno[2] ));
 sg13g2_nand3_1 _15141_ (.B(_07163_),
    .C(_07164_),
    .A(net583),
    .Y(_07177_));
 sg13g2_xnor2_1 _15142_ (.Y(_07178_),
    .A(_07176_),
    .B(_07177_));
 sg13g2_nor2_1 _15143_ (.A(_07171_),
    .B(_07178_),
    .Y(_00006_));
 sg13g2_nor2_2 _15144_ (.A(_07176_),
    .B(_07177_),
    .Y(_07179_));
 sg13g2_xnor2_1 _15145_ (.Y(_07180_),
    .A(_07161_),
    .B(_07179_));
 sg13g2_nor2_1 _15146_ (.A(_07171_),
    .B(_07180_),
    .Y(_00007_));
 sg13g2_nand2_1 _15147_ (.Y(_07181_),
    .A(_07161_),
    .B(_07179_));
 sg13g2_xor2_1 _15148_ (.B(_07181_),
    .A(_07158_),
    .X(_07182_));
 sg13g2_nor2_1 _15149_ (.A(_07171_),
    .B(_07182_),
    .Y(_00008_));
 sg13g2_inv_2 _15150_ (.Y(_07183_),
    .A(_07168_));
 sg13g2_buf_1 _15151_ (.A(_07183_),
    .X(_07184_));
 sg13g2_nand3_1 _15152_ (.B(_07158_),
    .C(_07179_),
    .A(_07161_),
    .Y(_07185_));
 sg13g2_xor2_1 _15153_ (.B(_07185_),
    .A(_07160_),
    .X(_07186_));
 sg13g2_nor2_1 _15154_ (.A(net518),
    .B(_07186_),
    .Y(_00009_));
 sg13g2_nand4_1 _15155_ (.B(_07160_),
    .C(_07158_),
    .A(_07161_),
    .Y(_07187_),
    .D(_07179_));
 sg13g2_xor2_1 _15156_ (.B(_07187_),
    .A(\clock_inst.frameno[6] ),
    .X(_07188_));
 sg13g2_nor2_1 _15157_ (.A(_07171_),
    .B(_07188_),
    .Y(_00010_));
 sg13g2_nor3_2 _15158_ (.A(_02285_),
    .B(_02756_),
    .C(_02297_),
    .Y(_07189_));
 sg13g2_a21o_1 _15159_ (.A2(_07167_),
    .A1(net4),
    .B1(_07189_),
    .X(_07190_));
 sg13g2_buf_1 _15160_ (.A(_07190_),
    .X(_07191_));
 sg13g2_nand2_1 _15161_ (.Y(_07192_),
    .A(net547),
    .B(_07191_));
 sg13g2_xnor2_1 _15162_ (.Y(_07193_),
    .A(net504),
    .B(_07192_));
 sg13g2_nor2_1 _15163_ (.A(_07184_),
    .B(_07193_),
    .Y(_00012_));
 sg13g2_nand2_1 _15164_ (.Y(_07194_),
    .A(net545),
    .B(_07191_));
 sg13g2_a21oi_1 _15165_ (.A1(net545),
    .A2(_00743_),
    .Y(_07195_),
    .B1(net509));
 sg13g2_nor2_1 _15166_ (.A(_07183_),
    .B(_07195_),
    .Y(_07196_));
 sg13g2_o21ai_1 _15167_ (.B1(_07196_),
    .Y(_07197_),
    .A1(_00775_),
    .A2(_07194_));
 sg13g2_a21oi_1 _15168_ (.A1(net453),
    .A2(_07192_),
    .Y(_00013_),
    .B1(_07197_));
 sg13g2_nor3_1 _15169_ (.A(net461),
    .B(net460),
    .C(_04902_),
    .Y(_07198_));
 sg13g2_a21o_1 _15170_ (.A2(_07167_),
    .A1(net3),
    .B1(_07198_),
    .X(_07199_));
 sg13g2_buf_1 _15171_ (.A(_07199_),
    .X(_07200_));
 sg13g2_inv_1 _15172_ (.Y(_07201_),
    .A(_07200_));
 sg13g2_nand2_1 _15173_ (.Y(_07202_),
    .A(net205),
    .B(_07201_));
 sg13g2_nand2_1 _15174_ (.Y(_07203_),
    .A(_00002_),
    .B(_07200_));
 sg13g2_nand2b_1 _15175_ (.Y(_07204_),
    .B(net552),
    .A_N(_07189_));
 sg13g2_a21oi_1 _15176_ (.A1(_07202_),
    .A2(_07203_),
    .Y(_00416_),
    .B1(_07204_));
 sg13g2_nand2_1 _15177_ (.Y(_07205_),
    .A(net230),
    .B(_07200_));
 sg13g2_xnor2_1 _15178_ (.Y(_07206_),
    .A(net215),
    .B(_07205_));
 sg13g2_nor2_1 _15179_ (.A(_07204_),
    .B(_07206_),
    .Y(_00418_));
 sg13g2_nand2b_1 _15180_ (.Y(_07207_),
    .B(_07200_),
    .A_N(_02261_));
 sg13g2_or2_1 _15181_ (.X(_07208_),
    .B(_07207_),
    .A(net134));
 sg13g2_xnor2_1 _15182_ (.Y(_07209_),
    .A(net200),
    .B(_07208_));
 sg13g2_nor2_1 _15183_ (.A(_07204_),
    .B(_07209_),
    .Y(_00421_));
 sg13g2_nand2_1 _15184_ (.Y(_07210_),
    .A(_00001_),
    .B(_07167_));
 sg13g2_nand2b_1 _15185_ (.Y(_07211_),
    .B(net116),
    .A_N(_07167_));
 sg13g2_nand2b_1 _15186_ (.Y(_07212_),
    .B(net552),
    .A_N(_07198_));
 sg13g2_a21oi_1 _15187_ (.A1(_07210_),
    .A2(_07211_),
    .Y(_00620_),
    .B1(_07212_));
 sg13g2_and2_1 _15188_ (.A(_05329_),
    .B(_07167_),
    .X(_07213_));
 sg13g2_buf_1 _15189_ (.A(_07213_),
    .X(_07214_));
 sg13g2_xnor2_1 _15190_ (.Y(_07215_),
    .A(net118),
    .B(_07214_));
 sg13g2_nor2_1 _15191_ (.A(_07212_),
    .B(_07215_),
    .Y(_00622_));
 sg13g2_nand2_1 _15192_ (.Y(_07216_),
    .A(net184),
    .B(_07214_));
 sg13g2_xnor2_1 _15193_ (.Y(_07217_),
    .A(net58),
    .B(_07216_));
 sg13g2_nor2_1 _15194_ (.A(_07212_),
    .B(_07217_),
    .Y(_00623_));
 sg13g2_nor2b_1 _15195_ (.A(_04985_),
    .B_N(_07214_),
    .Y(_07218_));
 sg13g2_xnor2_1 _15196_ (.Y(_07219_),
    .A(net179),
    .B(_07218_));
 sg13g2_nor2_1 _15197_ (.A(_07212_),
    .B(_07219_),
    .Y(_00625_));
 sg13g2_nand4_1 _15198_ (.B(_01018_),
    .C(_01019_),
    .A(_01017_),
    .Y(_07220_),
    .D(_01014_));
 sg13g2_buf_1 _15199_ (.A(_07220_),
    .X(_07221_));
 sg13g2_nand2_1 _15200_ (.Y(_07222_),
    .A(\clock_inst.vga_inst.vga_x[4] ),
    .B(_01028_));
 sg13g2_nor2_1 _15201_ (.A(_07221_),
    .B(_07222_),
    .Y(_07223_));
 sg13g2_and2_1 _15202_ (.A(net574),
    .B(_07223_),
    .X(_07224_));
 sg13g2_buf_1 _15203_ (.A(_07224_),
    .X(_07225_));
 sg13g2_nor2b_1 _15204_ (.A(_01023_),
    .B_N(_01024_),
    .Y(_07226_));
 sg13g2_nand3b_1 _15205_ (.B(_07225_),
    .C(_07226_),
    .Y(_07227_),
    .A_N(_01015_));
 sg13g2_inv_1 _15206_ (.Y(_07228_),
    .A(_01028_));
 sg13g2_nand3_1 _15207_ (.B(net574),
    .C(_01016_),
    .A(_07228_),
    .Y(_07229_));
 sg13g2_nand3_1 _15208_ (.B(_01018_),
    .C(_01019_),
    .A(_01017_),
    .Y(_07230_));
 sg13g2_buf_1 _15209_ (.A(_07230_),
    .X(_07231_));
 sg13g2_or3_1 _15210_ (.A(_01026_),
    .B(_07229_),
    .C(_07231_),
    .X(_07232_));
 sg13g2_buf_2 _15211_ (.A(_07232_),
    .X(_07233_));
 sg13g2_nand2_1 _15212_ (.Y(_07234_),
    .A(_07168_),
    .B(_07233_));
 sg13g2_buf_2 _15213_ (.A(_07234_),
    .X(_07235_));
 sg13g2_a21o_1 _15214_ (.A2(_07227_),
    .A1(\clock_inst.vga_inst.vga_horizontal_visible ),
    .B1(_07235_),
    .X(_00627_));
 sg13g2_nand2_1 _15215_ (.Y(_07236_),
    .A(_01015_),
    .B(_07226_));
 sg13g2_nor4_1 _15216_ (.A(\clock_inst.vga_inst.vga_x[4] ),
    .B(_01028_),
    .C(_07221_),
    .D(_07236_),
    .Y(_07237_));
 sg13g2_mux2_1 _15217_ (.A0(\clock_inst.vga_hs ),
    .A1(net574),
    .S(_07237_),
    .X(_07238_));
 sg13g2_or2_1 _15218_ (.X(_00628_),
    .B(_07238_),
    .A(net518));
 sg13g2_and3_1 _15219_ (.X(_00632_),
    .A(net552),
    .B(_00003_),
    .C(_07233_));
 sg13g2_xnor2_1 _15220_ (.Y(_07239_),
    .A(_01017_),
    .B(_01018_));
 sg13g2_nor2_1 _15221_ (.A(net518),
    .B(_07239_),
    .Y(_00633_));
 sg13g2_nand2_1 _15222_ (.Y(_07240_),
    .A(_01017_),
    .B(_01018_));
 sg13g2_xor2_1 _15223_ (.B(_07240_),
    .A(_01019_),
    .X(_07241_));
 sg13g2_nor2_1 _15224_ (.A(net518),
    .B(_07241_),
    .Y(_00634_));
 sg13g2_xor2_1 _15225_ (.B(_07231_),
    .A(_01014_),
    .X(_07242_));
 sg13g2_nor2_1 _15226_ (.A(_07235_),
    .B(_07242_),
    .Y(_00635_));
 sg13g2_xnor2_1 _15227_ (.Y(_07243_),
    .A(_01022_),
    .B(_07221_));
 sg13g2_nor2_1 _15228_ (.A(_07235_),
    .B(_07243_),
    .Y(_00636_));
 sg13g2_nor2_1 _15229_ (.A(_01022_),
    .B(_07221_),
    .Y(_07244_));
 sg13g2_xnor2_1 _15230_ (.Y(_07245_),
    .A(_01028_),
    .B(_07244_));
 sg13g2_nor2_1 _15231_ (.A(_07235_),
    .B(_07245_),
    .Y(_00637_));
 sg13g2_xnor2_1 _15232_ (.Y(_07246_),
    .A(net574),
    .B(_07223_));
 sg13g2_nor2_1 _15233_ (.A(_07235_),
    .B(_07246_),
    .Y(_00638_));
 sg13g2_xnor2_1 _15234_ (.Y(_07247_),
    .A(_01015_),
    .B(_07225_));
 sg13g2_nor2_1 _15235_ (.A(_07235_),
    .B(_07247_),
    .Y(_00639_));
 sg13g2_nand2_1 _15236_ (.Y(_07248_),
    .A(_01015_),
    .B(_07225_));
 sg13g2_xor2_1 _15237_ (.B(_07248_),
    .A(_01023_),
    .X(_07249_));
 sg13g2_nor2_1 _15238_ (.A(_07235_),
    .B(_07249_),
    .Y(_00640_));
 sg13g2_nand3_1 _15239_ (.B(_01023_),
    .C(_07225_),
    .A(_01015_),
    .Y(_07250_));
 sg13g2_xor2_1 _15240_ (.B(_07250_),
    .A(_01024_),
    .X(_07251_));
 sg13g2_nor2_1 _15241_ (.A(_07235_),
    .B(_07251_),
    .Y(_00641_));
 sg13g2_a21oi_1 _15242_ (.A1(_00742_),
    .A2(_00679_),
    .Y(_07252_),
    .B1(_00881_));
 sg13g2_o21ai_1 _15243_ (.B1(_07169_),
    .Y(_07253_),
    .A1(net454),
    .A2(_07191_));
 sg13g2_a21o_1 _15244_ (.A2(_07252_),
    .A1(_07191_),
    .B1(_07253_),
    .X(_00011_));
 sg13g2_o21ai_1 _15245_ (.B1(_00678_),
    .Y(_07254_),
    .A1(net364),
    .A2(_07194_));
 sg13g2_a21oi_1 _15246_ (.A1(net510),
    .A2(_07192_),
    .Y(_07255_),
    .B1(net453));
 sg13g2_o21ai_1 _15247_ (.B1(_07169_),
    .Y(_07256_),
    .A1(net515),
    .A2(_07255_));
 sg13g2_a21o_1 _15248_ (.A2(_07254_),
    .A1(_00881_),
    .B1(_07256_),
    .X(_00014_));
 sg13g2_o21ai_1 _15249_ (.B1(_02816_),
    .Y(_07257_),
    .A1(net193),
    .A2(_07201_));
 sg13g2_a21o_1 _15250_ (.A2(_07257_),
    .A1(_07205_),
    .B1(net518),
    .X(_00417_));
 sg13g2_nor3_1 _15251_ (.A(_00002_),
    .B(_02413_),
    .C(_07201_),
    .Y(_07258_));
 sg13g2_xnor2_1 _15252_ (.Y(_07259_),
    .A(net214),
    .B(_07258_));
 sg13g2_o21ai_1 _15253_ (.B1(net552),
    .Y(_00419_),
    .A1(_07189_),
    .A2(_07259_));
 sg13g2_xnor2_1 _15254_ (.Y(_07260_),
    .A(net134),
    .B(_07207_));
 sg13g2_o21ai_1 _15255_ (.B1(net552),
    .Y(_00420_),
    .A1(_07189_),
    .A2(_07260_));
 sg13g2_nand2_1 _15256_ (.Y(_07261_),
    .A(net180),
    .B(_07167_));
 sg13g2_xnor2_1 _15257_ (.Y(_07262_),
    .A(net176),
    .B(_07261_));
 sg13g2_nand2_1 _15258_ (.Y(_00621_),
    .A(net552),
    .B(_07262_));
 sg13g2_a21oi_1 _15259_ (.A1(net176),
    .A2(_05568_),
    .Y(_07263_),
    .B1(_07214_));
 sg13g2_o21ai_1 _15260_ (.B1(net165),
    .Y(_07264_),
    .A1(net460),
    .A2(_07263_));
 sg13g2_a21oi_1 _15261_ (.A1(_05437_),
    .A2(_07214_),
    .Y(_07265_),
    .B1(_07183_));
 sg13g2_nand2_1 _15262_ (.Y(_00624_),
    .A(_07264_),
    .B(_07265_));
 sg13g2_nor2_1 _15263_ (.A(net518),
    .B(_07227_),
    .Y(_00626_));
 sg13g2_nor2_1 _15264_ (.A(_01046_),
    .B(_07233_),
    .Y(_07266_));
 sg13g2_nand4_1 _15265_ (.B(_01048_),
    .C(net573),
    .A(_01047_),
    .Y(_07267_),
    .D(_07266_));
 sg13g2_nor4_1 _15266_ (.A(_07184_),
    .B(net543),
    .C(_01067_),
    .D(_07267_),
    .Y(_00629_));
 sg13g2_inv_1 _15267_ (.Y(_07268_),
    .A(net573));
 sg13g2_nor4_2 _15268_ (.A(_01026_),
    .B(_01046_),
    .C(_07229_),
    .Y(_07269_),
    .D(_07231_));
 sg13g2_nand3_1 _15269_ (.B(_01048_),
    .C(_07269_),
    .A(_01047_),
    .Y(_07270_));
 sg13g2_nor2_2 _15270_ (.A(_07268_),
    .B(_07270_),
    .Y(_07271_));
 sg13g2_nand3b_1 _15271_ (.B(_01044_),
    .C(_07271_),
    .Y(_07272_),
    .A_N(_01038_));
 sg13g2_o21ai_1 _15272_ (.B1(_07168_),
    .Y(_07273_),
    .A1(net150),
    .A2(_07233_));
 sg13g2_buf_1 _15273_ (.A(_07273_),
    .X(_07274_));
 sg13g2_a21o_1 _15274_ (.A2(_07272_),
    .A1(\clock_inst.vga_inst.vga_vertical_visible ),
    .B1(_07274_),
    .X(_00630_));
 sg13g2_nand2_1 _15275_ (.Y(_07275_),
    .A(_07268_),
    .B(_01037_));
 sg13g2_nor2_1 _15276_ (.A(_01067_),
    .B(_07275_),
    .Y(_07276_));
 sg13g2_nand3_1 _15277_ (.B(_07269_),
    .C(_07276_),
    .A(_01049_),
    .Y(_07277_));
 sg13g2_inv_1 _15278_ (.Y(_07278_),
    .A(\clock_inst.vga_inst.vga_y[0] ));
 sg13g2_nand3b_1 _15279_ (.B(_07278_),
    .C(_01049_),
    .Y(_07279_),
    .A_N(_01045_));
 sg13g2_buf_1 _15280_ (.A(_07279_),
    .X(_07280_));
 sg13g2_nand2b_1 _15281_ (.Y(_07281_),
    .B(_07276_),
    .A_N(_07233_));
 sg13g2_o21ai_1 _15282_ (.B1(\clock_inst.vga_inst.vga_vs ),
    .Y(_07282_),
    .A1(_07280_),
    .A2(_07281_));
 sg13g2_nand3_1 _15283_ (.B(_07277_),
    .C(_07282_),
    .A(net552),
    .Y(_00631_));
 sg13g2_xnor2_1 _15284_ (.Y(_07283_),
    .A(_07278_),
    .B(_07233_));
 sg13g2_nor2_1 _15285_ (.A(net518),
    .B(_07283_),
    .Y(_00642_));
 sg13g2_nor2_1 _15286_ (.A(_07278_),
    .B(_07233_),
    .Y(_07284_));
 sg13g2_xnor2_1 _15287_ (.Y(_07285_),
    .A(_01045_),
    .B(_07284_));
 sg13g2_nor2_1 _15288_ (.A(net518),
    .B(_07285_),
    .Y(_00643_));
 sg13g2_xnor2_1 _15289_ (.Y(_07286_),
    .A(_01048_),
    .B(_07269_));
 sg13g2_nor2_1 _15290_ (.A(net24),
    .B(_07286_),
    .Y(_00644_));
 sg13g2_nand2_1 _15291_ (.Y(_07287_),
    .A(_01048_),
    .B(_07269_));
 sg13g2_xor2_1 _15292_ (.B(_07287_),
    .A(_01047_),
    .X(_07288_));
 sg13g2_nor2_1 _15293_ (.A(net24),
    .B(_07288_),
    .Y(_00645_));
 sg13g2_xnor2_1 _15294_ (.Y(_07289_),
    .A(_07268_),
    .B(_07270_));
 sg13g2_nor2_1 _15295_ (.A(net24),
    .B(_07289_),
    .Y(_00646_));
 sg13g2_xnor2_1 _15296_ (.Y(_07290_),
    .A(_01038_),
    .B(_07271_));
 sg13g2_nor2_1 _15297_ (.A(net24),
    .B(_07290_),
    .Y(_00647_));
 sg13g2_nand2_1 _15298_ (.Y(_07291_),
    .A(net543),
    .B(_07271_));
 sg13g2_xor2_1 _15299_ (.B(_07291_),
    .A(_01040_),
    .X(_07292_));
 sg13g2_nor2_1 _15300_ (.A(net24),
    .B(_07292_),
    .Y(_00648_));
 sg13g2_nand3_1 _15301_ (.B(_01040_),
    .C(_07271_),
    .A(net543),
    .Y(_07293_));
 sg13g2_xor2_1 _15302_ (.B(_07293_),
    .A(_01041_),
    .X(_07294_));
 sg13g2_nor2_1 _15303_ (.A(net24),
    .B(_07294_),
    .Y(_00649_));
 sg13g2_nand2_1 _15304_ (.Y(_07295_),
    .A(_01040_),
    .B(_01041_));
 sg13g2_nor2_1 _15305_ (.A(_07295_),
    .B(_07291_),
    .Y(_07296_));
 sg13g2_xnor2_1 _15306_ (.Y(_07297_),
    .A(_01042_),
    .B(_07296_));
 sg13g2_nor2_1 _15307_ (.A(net24),
    .B(_07297_),
    .Y(_00650_));
 sg13g2_nand2_1 _15308_ (.Y(_07298_),
    .A(_01042_),
    .B(_07296_));
 sg13g2_xor2_1 _15309_ (.B(_07298_),
    .A(_01039_),
    .X(_07299_));
 sg13g2_nor2_1 _15310_ (.A(net24),
    .B(_07299_),
    .Y(_00651_));
 sg13g2_nor4_1 _15311_ (.A(_01022_),
    .B(_01023_),
    .C(_01039_),
    .D(_01021_),
    .Y(_07300_));
 sg13g2_nor4_1 _15312_ (.A(_01042_),
    .B(_01065_),
    .C(_07295_),
    .D(_07280_),
    .Y(_07301_));
 sg13g2_nor2b_1 _15313_ (.A(net574),
    .B_N(_01024_),
    .Y(_07302_));
 sg13g2_nor2b_1 _15314_ (.A(_01048_),
    .B_N(_01047_),
    .Y(_07303_));
 sg13g2_nor3_1 _15315_ (.A(_01045_),
    .B(\clock_inst.vga_inst.vga_y[0] ),
    .C(_01041_),
    .Y(_07304_));
 sg13g2_nand4_1 _15316_ (.B(_01040_),
    .C(_07303_),
    .A(net543),
    .Y(_07305_),
    .D(_07304_));
 sg13g2_xnor2_1 _15317_ (.Y(_07306_),
    .A(net573),
    .B(_01042_));
 sg13g2_nor2_1 _15318_ (.A(_07305_),
    .B(_07306_),
    .Y(_07307_));
 sg13g2_nor2b_1 _15319_ (.A(_01024_),
    .B_N(net574),
    .Y(_07308_));
 sg13g2_a22oi_1 _15320_ (.Y(_07309_),
    .B1(_07307_),
    .B2(_07308_),
    .A2(_07302_),
    .A1(_07301_));
 sg13g2_a221oi_1 _15321_ (.B2(_07301_),
    .C1(_01028_),
    .B1(_07308_),
    .A1(_07302_),
    .Y(_07310_),
    .A2(_07307_));
 sg13g2_a21oi_1 _15322_ (.A1(_01028_),
    .A2(_07309_),
    .Y(_07311_),
    .B1(_07310_));
 sg13g2_or3_1 _15323_ (.A(\clock_inst.sec_tile.e[17] ),
    .B(\clock_inst.sec_tile.e[35] ),
    .C(\clock_inst.sec_tile.e[53] ),
    .X(_07312_));
 sg13g2_nand3_1 _15324_ (.B(_01015_),
    .C(_01020_),
    .A(_01014_),
    .Y(_07313_));
 sg13g2_nand2b_1 _15325_ (.Y(_07314_),
    .B(_01023_),
    .A_N(_01024_));
 sg13g2_nor4_1 _15326_ (.A(net574),
    .B(_07222_),
    .C(_07313_),
    .D(_07314_),
    .Y(_07315_));
 sg13g2_nand3_1 _15327_ (.B(_07228_),
    .C(_01027_),
    .A(_01022_),
    .Y(_07316_));
 sg13g2_nor4_1 _15328_ (.A(_01023_),
    .B(_01024_),
    .C(_07313_),
    .D(_07316_),
    .Y(_07317_));
 sg13g2_nor4_1 _15329_ (.A(net573),
    .B(net543),
    .C(_01067_),
    .D(_07280_),
    .Y(_07318_));
 sg13g2_nor2_1 _15330_ (.A(_01039_),
    .B(_07275_),
    .Y(_07319_));
 sg13g2_nor4_1 _15331_ (.A(_01040_),
    .B(_01041_),
    .C(_01042_),
    .D(_07280_),
    .Y(_07320_));
 sg13g2_nand3_1 _15332_ (.B(_07319_),
    .C(_07320_),
    .A(_07317_),
    .Y(_07321_));
 sg13g2_nand2b_1 _15333_ (.Y(_07322_),
    .B(_07321_),
    .A_N(_07318_));
 sg13g2_o21ai_1 _15334_ (.B1(_07322_),
    .Y(_07323_),
    .A1(_07315_),
    .A2(_07317_));
 sg13g2_nor4_1 _15335_ (.A(_01037_),
    .B(_01021_),
    .C(_07314_),
    .D(_07316_),
    .Y(_07324_));
 sg13g2_a21oi_1 _15336_ (.A1(net543),
    .A2(_07315_),
    .Y(_07325_),
    .B1(_07324_));
 sg13g2_nor3_1 _15337_ (.A(net573),
    .B(_01039_),
    .C(_07325_),
    .Y(_07326_));
 sg13g2_nand3_1 _15338_ (.B(net543),
    .C(_01039_),
    .A(net573),
    .Y(_07327_));
 sg13g2_nor4_1 _15339_ (.A(_01021_),
    .B(_07314_),
    .C(_07316_),
    .D(_07327_),
    .Y(_07328_));
 sg13g2_o21ai_1 _15340_ (.B1(_07320_),
    .Y(_07329_),
    .A1(_07326_),
    .A2(_07328_));
 sg13g2_nand3_1 _15341_ (.B(_07323_),
    .C(_07329_),
    .A(_07312_),
    .Y(_07330_));
 sg13g2_a21oi_1 _15342_ (.A1(_07300_),
    .A2(_07311_),
    .Y(_07331_),
    .B1(_07330_));
 sg13g2_nor2_1 _15343_ (.A(net448),
    .B(_07331_),
    .Y(_00652_));
 sg13g2_nor3_1 _15344_ (.A(\clock_inst.hour_tile.e[17] ),
    .B(\clock_inst.hour_tile.e[35] ),
    .C(\clock_inst.hour_tile.e[53] ),
    .Y(_07332_));
 sg13g2_nor3_2 _15345_ (.A(\clock_inst.min_tile.e[17] ),
    .B(\clock_inst.min_tile.e[35] ),
    .C(\clock_inst.min_tile.e[53] ),
    .Y(_07333_));
 sg13g2_nand2b_1 _15346_ (.Y(_07334_),
    .B(_07333_),
    .A_N(_07332_));
 sg13g2_a21oi_1 _15347_ (.A1(_07331_),
    .A2(_07334_),
    .Y(_00653_),
    .B1(net448));
 sg13g2_nor2_1 _15348_ (.A(_07333_),
    .B(_07332_),
    .Y(_07335_));
 sg13g2_a21oi_1 _15349_ (.A1(_07331_),
    .A2(_07335_),
    .Y(_00654_),
    .B1(net448));
 sg13g2_buf_2 _15350_ (.A(ui_in[0]),
    .X(_07336_));
 sg13g2_nand2_1 _15351_ (.Y(_07337_),
    .A(_07336_),
    .B(\clock_inst.vga_horizontal_blank_strobe ));
 sg13g2_inv_1 _15352_ (.Y(_07338_),
    .A(_07336_));
 sg13g2_nand2_1 _15353_ (.Y(_07339_),
    .A(_07164_),
    .B(_07338_));
 sg13g2_buf_1 _15354_ (.A(ui_in[1]),
    .X(_07340_));
 sg13g2_inv_1 _15355_ (.Y(_07341_),
    .A(_07340_));
 sg13g2_nor2_1 _15356_ (.A(net2),
    .B(net1),
    .Y(_07342_));
 sg13g2_buf_2 _15357_ (.A(_07342_),
    .X(_07343_));
 sg13g2_nand2_1 _15358_ (.Y(_07344_),
    .A(_07341_),
    .B(_07343_));
 sg13g2_a21oi_1 _15359_ (.A1(_07337_),
    .A2(_07339_),
    .Y(net5),
    .B1(_07344_));
 sg13g2_nand2_1 _15360_ (.Y(_07345_),
    .A(_07163_),
    .B(_07338_));
 sg13g2_a21oi_1 _15361_ (.A1(_07337_),
    .A2(_07345_),
    .Y(net6),
    .B1(_07344_));
 sg13g2_buf_1 _15362_ (.A(_07340_),
    .X(_07346_));
 sg13g2_nor2_1 _15363_ (.A(\clock_inst.frameno[2] ),
    .B(_07346_),
    .Y(_07347_));
 sg13g2_a21oi_1 _15364_ (.A1(_02711_),
    .A2(net551),
    .Y(_07348_),
    .B1(_07347_));
 sg13g2_nor2_2 _15365_ (.A(_07338_),
    .B(_07340_),
    .Y(_07349_));
 sg13g2_nand2_1 _15366_ (.Y(_07350_),
    .A(net163),
    .B(_07349_));
 sg13g2_o21ai_1 _15367_ (.B1(_07350_),
    .Y(_07351_),
    .A1(_07336_),
    .A2(_07348_));
 sg13g2_o21ai_1 _15368_ (.B1(_07343_),
    .Y(_07352_),
    .A1(_07338_),
    .A2(_07341_));
 sg13g2_buf_1 _15369_ (.A(_07352_),
    .X(_07353_));
 sg13g2_a22oi_1 _15370_ (.Y(net7),
    .B1(_07353_),
    .B2(_00675_),
    .A2(_07351_),
    .A1(_07343_));
 sg13g2_nor2_1 _15371_ (.A(_07161_),
    .B(net551),
    .Y(_07354_));
 sg13g2_a21oi_1 _15372_ (.A1(_02550_),
    .A2(net551),
    .Y(_07355_),
    .B1(_07354_));
 sg13g2_nand2_1 _15373_ (.Y(_07356_),
    .A(_05203_),
    .B(_07349_));
 sg13g2_o21ai_1 _15374_ (.B1(_07356_),
    .Y(_07357_),
    .A1(_07336_),
    .A2(_07355_));
 sg13g2_a22oi_1 _15375_ (.Y(net8),
    .B1(_07357_),
    .B2(_07343_),
    .A2(_07353_),
    .A1(_00790_));
 sg13g2_nor2_1 _15376_ (.A(_07158_),
    .B(net551),
    .Y(_07358_));
 sg13g2_a21oi_1 _15377_ (.A1(_02442_),
    .A2(net551),
    .Y(_07359_),
    .B1(_07358_));
 sg13g2_nand2_1 _15378_ (.Y(_07360_),
    .A(net170),
    .B(_07349_));
 sg13g2_o21ai_1 _15379_ (.B1(_07360_),
    .Y(_07361_),
    .A1(_07336_),
    .A2(_07359_));
 sg13g2_a22oi_1 _15380_ (.Y(net9),
    .B1(_07361_),
    .B2(_07343_),
    .A2(_07353_),
    .A1(_00680_));
 sg13g2_nor2_1 _15381_ (.A(_07160_),
    .B(net551),
    .Y(_07362_));
 sg13g2_a21oi_1 _15382_ (.A1(_02586_),
    .A2(net551),
    .Y(_07363_),
    .B1(_07362_));
 sg13g2_nand2_1 _15383_ (.Y(_07364_),
    .A(net58),
    .B(_07349_));
 sg13g2_o21ai_1 _15384_ (.B1(_07364_),
    .Y(_07365_),
    .A1(_07336_),
    .A2(_07363_));
 sg13g2_a22oi_1 _15385_ (.Y(net10),
    .B1(_07365_),
    .B2(_07343_),
    .A2(_07353_),
    .A1(_00672_));
 sg13g2_mux2_1 _15386_ (.A0(\clock_inst.frameno[6] ),
    .A1(_02415_),
    .S(_07346_),
    .X(_07366_));
 sg13g2_a22oi_1 _15387_ (.Y(_07367_),
    .B1(_07366_),
    .B2(_07338_),
    .A2(_07349_),
    .A1(_05393_));
 sg13g2_nor2b_1 _15388_ (.A(_07367_),
    .B_N(_07343_),
    .Y(net11));
 sg13g2_nor2_1 _15389_ (.A(_02664_),
    .B(_07336_),
    .Y(_07368_));
 sg13g2_a22oi_1 _15390_ (.Y(_07369_),
    .B1(_07368_),
    .B2(net551),
    .A2(_07349_),
    .A1(net179));
 sg13g2_nor2b_1 _15391_ (.A(_07369_),
    .B_N(_07343_),
    .Y(net12));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _15393_ (.A(net584),
    .X(uio_oe[0]));
 sg13g2_buf_1 _15394_ (.A(net585),
    .X(uio_oe[1]));
 sg13g2_buf_1 _15395_ (.A(net586),
    .X(uio_oe[2]));
 sg13g2_buf_1 _15396_ (.A(net587),
    .X(uio_oe[3]));
 sg13g2_buf_1 _15397_ (.A(net588),
    .X(uio_oe[4]));
 sg13g2_buf_1 _15398_ (.A(net589),
    .X(uio_oe[5]));
 sg13g2_buf_1 _15399_ (.A(net590),
    .X(uio_oe[6]));
 sg13g2_buf_1 _15400_ (.A(net591),
    .X(uio_oe[7]));
 sg13g2_buf_1 _15401_ (.A(net17),
    .X(net13));
 sg13g2_buf_1 _15402_ (.A(net18),
    .X(net14));
 sg13g2_buf_1 _15403_ (.A(net19),
    .X(net15));
 sg13g2_buf_1 _15404_ (.A(\clock_inst.vga_inst.vga_vs ),
    .X(net16));
 sg13g2_buf_1 _15405_ (.A(\clock_inst.vga_hs ),
    .X(net20));
 sg13g2_dfrbp_1 \clock_inst.frameno[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net592),
    .D(_00004_),
    .Q_N(_00000_),
    .Q(\clock_inst.frameno[0] ));
 sg13g2_dfrbp_1 \clock_inst.frameno[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net593),
    .D(_00005_),
    .Q_N(_08016_),
    .Q(\clock_inst.frameno[1] ));
 sg13g2_dfrbp_1 \clock_inst.frameno[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net594),
    .D(_00006_),
    .Q_N(_08015_),
    .Q(\clock_inst.frameno[2] ));
 sg13g2_dfrbp_1 \clock_inst.frameno[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net595),
    .D(_00007_),
    .Q_N(_08014_),
    .Q(\clock_inst.frameno[3] ));
 sg13g2_dfrbp_1 \clock_inst.frameno[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net596),
    .D(_00008_),
    .Q_N(_08013_),
    .Q(\clock_inst.frameno[4] ));
 sg13g2_dfrbp_1 \clock_inst.frameno[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net597),
    .D(_00009_),
    .Q_N(_08012_),
    .Q(\clock_inst.frameno[5] ));
 sg13g2_dfrbp_1 \clock_inst.frameno[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net598),
    .D(_00010_),
    .Q_N(_08011_),
    .Q(\clock_inst.frameno[6] ));
 sg13g2_dfrbp_1 \clock_inst.hour[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net599),
    .D(_00011_),
    .Q_N(_08010_),
    .Q(\clock_inst.hour[0] ));
 sg13g2_dfrbp_1 \clock_inst.hour[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net600),
    .D(_00012_),
    .Q_N(_08009_),
    .Q(\clock_inst.hour[1] ));
 sg13g2_dfrbp_1 \clock_inst.hour[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net601),
    .D(_00013_),
    .Q_N(_08008_),
    .Q(\clock_inst.hour[2] ));
 sg13g2_dfrbp_1 \clock_inst.hour[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net602),
    .D(_00014_),
    .Q_N(_08007_),
    .Q(\clock_inst.hour[3] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net603),
    .D(_00015_),
    .Q_N(_08006_),
    .Q(\clock_inst.hour_a[0] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[17]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net604),
    .D(_00016_),
    .Q_N(_08005_),
    .Q(\clock_inst.hour_a[10] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[19]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net605),
    .D(_00017_),
    .Q_N(_08004_),
    .Q(\clock_inst.hour_a[19] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net606),
    .D(_00018_),
    .Q_N(_08003_),
    .Q(\clock_inst.hour_a[1] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[20]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net607),
    .D(_00019_),
    .Q_N(_08002_),
    .Q(\clock_inst.hour_a[20] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[21]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net608),
    .D(_00020_),
    .Q_N(_08001_),
    .Q(\clock_inst.hour_a[21] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[22]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net609),
    .D(_00021_),
    .Q_N(_08000_),
    .Q(\clock_inst.hour_a[22] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[23]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net610),
    .D(_00022_),
    .Q_N(_07999_),
    .Q(\clock_inst.hour_a[23] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net611),
    .D(_00023_),
    .Q_N(_07998_),
    .Q(\clock_inst.hour_a[2] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[35]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net612),
    .D(_00024_),
    .Q_N(_07997_),
    .Q(\clock_inst.hour_a[24] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[36]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net613),
    .D(_00025_),
    .Q_N(_07996_),
    .Q(\clock_inst.hour_a[36] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[37]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net614),
    .D(_00026_),
    .Q_N(_07995_),
    .Q(\clock_inst.hour_a[37] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[38]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net615),
    .D(_00027_),
    .Q_N(_07994_),
    .Q(\clock_inst.hour_a[38] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[39]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net616),
    .D(_00028_),
    .Q_N(_07993_),
    .Q(\clock_inst.hour_a[39] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[3]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net617),
    .D(_00029_),
    .Q_N(_07992_),
    .Q(\clock_inst.hour_a[3] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[40]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net618),
    .D(_00030_),
    .Q_N(_07991_),
    .Q(\clock_inst.hour_a[40] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[41]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net619),
    .D(_00031_),
    .Q_N(_07990_),
    .Q(\clock_inst.hour_a[41] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[42]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net620),
    .D(_00032_),
    .Q_N(_07989_),
    .Q(\clock_inst.hour_a[42] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[43]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net621),
    .D(_00033_),
    .Q_N(_07988_),
    .Q(\clock_inst.hour_a[43] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[52]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net622),
    .D(_00034_),
    .Q_N(_07987_),
    .Q(\clock_inst.hour_a[44] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[5]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net623),
    .D(_00035_),
    .Q_N(_07986_),
    .Q(\clock_inst.hour_a[5] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[6]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net624),
    .D(_00036_),
    .Q_N(_07985_),
    .Q(\clock_inst.hour_a[6] ));
 sg13g2_dfrbp_1 \clock_inst.hour_a[7]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net625),
    .D(_00037_),
    .Q_N(_07984_),
    .Q(\clock_inst.hour_a[7] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net626),
    .D(_00038_),
    .Q_N(_07983_),
    .Q(\clock_inst.hour_b[0] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[17]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net627),
    .D(_00039_),
    .Q_N(_07982_),
    .Q(\clock_inst.hour_b[10] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[19]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net628),
    .D(_00040_),
    .Q_N(_07981_),
    .Q(\clock_inst.hour_b[19] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net629),
    .D(_00041_),
    .Q_N(_07980_),
    .Q(\clock_inst.hour_b[1] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[20]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net630),
    .D(_00042_),
    .Q_N(_07979_),
    .Q(\clock_inst.hour_b[20] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[22]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net631),
    .D(_00043_),
    .Q_N(_07978_),
    .Q(\clock_inst.hour_b[22] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[23]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net632),
    .D(_00044_),
    .Q_N(_07977_),
    .Q(\clock_inst.hour_b[23] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net633),
    .D(_00045_),
    .Q_N(_07976_),
    .Q(\clock_inst.hour_b[2] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[35]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net634),
    .D(_00046_),
    .Q_N(_07975_),
    .Q(\clock_inst.hour_b[21] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[36]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net635),
    .D(_00047_),
    .Q_N(_07974_),
    .Q(\clock_inst.hour_b[36] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[37]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net636),
    .D(_00048_),
    .Q_N(_07973_),
    .Q(\clock_inst.hour_b[37] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[38]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net637),
    .D(_00049_),
    .Q_N(_07972_),
    .Q(\clock_inst.hour_b[38] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[39]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net638),
    .D(_00050_),
    .Q_N(_07971_),
    .Q(\clock_inst.hour_b[39] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[40]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net639),
    .D(_00051_),
    .Q_N(_07970_),
    .Q(\clock_inst.hour_b[40] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[41]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net640),
    .D(_00052_),
    .Q_N(_07969_),
    .Q(\clock_inst.hour_b[41] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[42]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net641),
    .D(_00053_),
    .Q_N(_07968_),
    .Q(\clock_inst.hour_b[42] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[4]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net642),
    .D(_00054_),
    .Q_N(_07967_),
    .Q(\clock_inst.hour_b[4] ));
 sg13g2_dfrbp_1 \clock_inst.hour_b[5]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net643),
    .D(_00055_),
    .Q_N(_07966_),
    .Q(\clock_inst.hour_b[5] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net644),
    .D(_00056_),
    .Q_N(_07965_),
    .Q(\clock_inst.hour_c[10] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[11]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net645),
    .D(_00057_),
    .Q_N(_07964_),
    .Q(\clock_inst.hour_c[11] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[12]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net646),
    .D(_00058_),
    .Q_N(_07963_),
    .Q(\clock_inst.hour_c[12] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[13]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net647),
    .D(_00059_),
    .Q_N(_07962_),
    .Q(\clock_inst.hour_c[13] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[14]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net648),
    .D(_00060_),
    .Q_N(_07961_),
    .Q(\clock_inst.hour_c[14] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[15]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net649),
    .D(_00061_),
    .Q_N(_07960_),
    .Q(\clock_inst.hour_c[15] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[16]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net650),
    .D(_00062_),
    .Q_N(_07959_),
    .Q(\clock_inst.hour_c[16] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[17]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net651),
    .D(_00063_),
    .Q_N(_07958_),
    .Q(\clock_inst.hour_c[17] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[18]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net652),
    .D(_00064_),
    .Q_N(_07957_),
    .Q(\clock_inst.hour_a[18] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[19]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net653),
    .D(_00065_),
    .Q_N(_07956_),
    .Q(\clock_inst.hour_c[19] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[1]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net654),
    .D(_00066_),
    .Q_N(_07955_),
    .Q(\clock_inst.hour_c[1] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[21]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net655),
    .D(_00067_),
    .Q_N(_07954_),
    .Q(\clock_inst.hour_c[21] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[23]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net656),
    .D(_00068_),
    .Q_N(_07953_),
    .Q(\clock_inst.hour_c[23] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[24]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net657),
    .D(_00069_),
    .Q_N(_07952_),
    .Q(\clock_inst.hour_c[24] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[25]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net658),
    .D(_00070_),
    .Q_N(_07951_),
    .Q(\clock_inst.hour_c[25] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[26]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net659),
    .D(_00071_),
    .Q_N(_07950_),
    .Q(\clock_inst.hour_c[26] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[27]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net660),
    .D(_00072_),
    .Q_N(_07949_),
    .Q(\clock_inst.hour_c[27] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[28]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net661),
    .D(_00073_),
    .Q_N(_07948_),
    .Q(\clock_inst.hour_c[28] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[29]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net662),
    .D(_00074_),
    .Q_N(_07947_),
    .Q(\clock_inst.hour_c[29] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[30]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net663),
    .D(_00075_),
    .Q_N(_07946_),
    .Q(\clock_inst.hour_c[30] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[31]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net664),
    .D(_00076_),
    .Q_N(_07945_),
    .Q(\clock_inst.hour_a[4] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[32]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net665),
    .D(_00077_),
    .Q_N(_07944_),
    .Q(\clock_inst.hour_c[32] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[35]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net666),
    .D(_00078_),
    .Q_N(_07943_),
    .Q(\clock_inst.hour_c[33] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[36]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net667),
    .D(_00079_),
    .Q_N(_07942_),
    .Q(\clock_inst.hour_c[0] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[37]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net668),
    .D(_00080_),
    .Q_N(_07941_),
    .Q(\clock_inst.hour_c[37] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[39]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net669),
    .D(_00081_),
    .Q_N(_07940_),
    .Q(\clock_inst.hour_c[2] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[40]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net670),
    .D(_00082_),
    .Q_N(_07939_),
    .Q(\clock_inst.hour_c[40] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[41]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net671),
    .D(_00083_),
    .Q_N(_07938_),
    .Q(\clock_inst.hour_c[41] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[42]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net672),
    .D(_00084_),
    .Q_N(_07937_),
    .Q(\clock_inst.hour_c[42] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[43]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net673),
    .D(_00085_),
    .Q_N(_07936_),
    .Q(\clock_inst.hour_c[43] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[44]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net674),
    .D(_00086_),
    .Q_N(_07935_),
    .Q(\clock_inst.hour_c[44] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[45]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net675),
    .D(_00087_),
    .Q_N(_07934_),
    .Q(\clock_inst.hour_c[45] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[46]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net676),
    .D(_00088_),
    .Q_N(_07933_),
    .Q(\clock_inst.hour_c[46] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[49]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net677),
    .D(_00089_),
    .Q_N(_07932_),
    .Q(\clock_inst.hour_c[49] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[50]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net678),
    .D(_00090_),
    .Q_N(_07931_),
    .Q(\clock_inst.hour_c[50] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[51]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net679),
    .D(_00091_),
    .Q_N(_07930_),
    .Q(\clock_inst.hour_c[51] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[52]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net680),
    .D(_00092_),
    .Q_N(_07929_),
    .Q(\clock_inst.hour_c[52] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net681),
    .D(_00093_),
    .Q_N(_07928_),
    .Q(\clock_inst.hour_c[5] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[6]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net682),
    .D(_00094_),
    .Q_N(_07927_),
    .Q(\clock_inst.hour_c[6] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[7]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net683),
    .D(_00095_),
    .Q_N(_07926_),
    .Q(\clock_inst.hour_c[7] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[8]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net684),
    .D(_00096_),
    .Q_N(_07925_),
    .Q(\clock_inst.hour_c[8] ));
 sg13g2_dfrbp_1 \clock_inst.hour_c[9]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net685),
    .D(_00097_),
    .Q_N(_07924_),
    .Q(\clock_inst.hour_c[9] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net686),
    .D(_00098_),
    .Q_N(_07923_),
    .Q(\clock_inst.hour_tile.e0[0] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net687),
    .D(_00099_),
    .Q_N(_07922_),
    .Q(\clock_inst.hour_tile.e0[10] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[11]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net688),
    .D(_00100_),
    .Q_N(_07921_),
    .Q(\clock_inst.hour_tile.e0[11] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[12]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net689),
    .D(_00101_),
    .Q_N(_07920_),
    .Q(\clock_inst.hour_tile.e0[12] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[13]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net690),
    .D(_00102_),
    .Q_N(_07919_),
    .Q(\clock_inst.hour_tile.e0[13] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[14]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net691),
    .D(_00103_),
    .Q_N(_07918_),
    .Q(\clock_inst.hour_tile.e0[14] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[15]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net692),
    .D(_00104_),
    .Q_N(_07917_),
    .Q(\clock_inst.hour_tile.e0[15] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[16]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net693),
    .D(_00105_),
    .Q_N(_07916_),
    .Q(\clock_inst.hour_tile.e0[16] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[17]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net694),
    .D(_00106_),
    .Q_N(_07915_),
    .Q(\clock_inst.hour_tile.e0[17] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[18]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net695),
    .D(_00107_),
    .Q_N(_07914_),
    .Q(\clock_inst.hour_tile.e0[18] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[19]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net696),
    .D(_00108_),
    .Q_N(_07913_),
    .Q(\clock_inst.hour_tile.e0[19] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net697),
    .D(_00109_),
    .Q_N(_07912_),
    .Q(\clock_inst.hour_tile.e0[1] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[20]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net698),
    .D(_00110_),
    .Q_N(_07911_),
    .Q(\clock_inst.hour_tile.e0[20] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[21]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net699),
    .D(_00111_),
    .Q_N(_07910_),
    .Q(\clock_inst.hour_tile.e0[21] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[22]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net700),
    .D(_00112_),
    .Q_N(_07909_),
    .Q(\clock_inst.hour_tile.e0[22] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[23]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net701),
    .D(_00113_),
    .Q_N(_07908_),
    .Q(\clock_inst.hour_tile.e0[23] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[24]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net702),
    .D(_00114_),
    .Q_N(_07907_),
    .Q(\clock_inst.hour_tile.e0[24] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[25]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net703),
    .D(_00115_),
    .Q_N(_07906_),
    .Q(\clock_inst.hour_tile.e0[25] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[26]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net704),
    .D(_00116_),
    .Q_N(_07905_),
    .Q(\clock_inst.hour_tile.e0[26] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[27]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net705),
    .D(_00117_),
    .Q_N(_07904_),
    .Q(\clock_inst.hour_tile.e0[27] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[28]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net706),
    .D(_00118_),
    .Q_N(_07903_),
    .Q(\clock_inst.hour_tile.e0[28] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[29]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net707),
    .D(_00119_),
    .Q_N(_07902_),
    .Q(\clock_inst.hour_tile.e0[29] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net708),
    .D(_00120_),
    .Q_N(_07901_),
    .Q(\clock_inst.hour_tile.e0[2] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[30]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net709),
    .D(_00121_),
    .Q_N(_07900_),
    .Q(\clock_inst.hour_tile.e0[30] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[31]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net710),
    .D(_00122_),
    .Q_N(_07899_),
    .Q(\clock_inst.hour_tile.e0[31] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[32]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net711),
    .D(_00123_),
    .Q_N(_07898_),
    .Q(\clock_inst.hour_tile.e0[32] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[33]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net712),
    .D(_00124_),
    .Q_N(_07897_),
    .Q(\clock_inst.hour_tile.e0[33] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[34]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net713),
    .D(_00125_),
    .Q_N(_07896_),
    .Q(\clock_inst.hour_tile.e0[34] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[35]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net714),
    .D(_00126_),
    .Q_N(_07895_),
    .Q(\clock_inst.hour_tile.e0[35] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[36]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net715),
    .D(_00127_),
    .Q_N(_07894_),
    .Q(\clock_inst.hour_tile.e0[36] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[37]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net716),
    .D(_00128_),
    .Q_N(_07893_),
    .Q(\clock_inst.hour_tile.e0[37] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[38]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net717),
    .D(_00129_),
    .Q_N(_07892_),
    .Q(\clock_inst.hour_tile.e0[38] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[39]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net718),
    .D(_00130_),
    .Q_N(_07891_),
    .Q(\clock_inst.hour_tile.e0[39] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[3]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net719),
    .D(_00131_),
    .Q_N(_07890_),
    .Q(\clock_inst.hour_tile.e0[3] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[40]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net720),
    .D(_00132_),
    .Q_N(_07889_),
    .Q(\clock_inst.hour_tile.e0[40] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[41]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net721),
    .D(_00133_),
    .Q_N(_07888_),
    .Q(\clock_inst.hour_tile.e0[41] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[42]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net722),
    .D(_00134_),
    .Q_N(_07887_),
    .Q(\clock_inst.hour_tile.e0[42] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[43]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net723),
    .D(_00135_),
    .Q_N(_07886_),
    .Q(\clock_inst.hour_tile.e0[43] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[44]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net724),
    .D(_00136_),
    .Q_N(_07885_),
    .Q(\clock_inst.hour_tile.e0[44] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[45]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net725),
    .D(_00137_),
    .Q_N(_07884_),
    .Q(\clock_inst.hour_tile.e0[45] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[46]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net726),
    .D(_00138_),
    .Q_N(_07883_),
    .Q(\clock_inst.hour_tile.e0[46] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[47]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net727),
    .D(_00139_),
    .Q_N(_07882_),
    .Q(\clock_inst.hour_tile.e0[47] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[48]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net728),
    .D(_00140_),
    .Q_N(_07881_),
    .Q(\clock_inst.hour_tile.e0[48] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[49]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net729),
    .D(_00141_),
    .Q_N(_07880_),
    .Q(\clock_inst.hour_tile.e0[49] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[4]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net730),
    .D(_00142_),
    .Q_N(_07879_),
    .Q(\clock_inst.hour_tile.e0[4] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[50]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net731),
    .D(_00143_),
    .Q_N(_07878_),
    .Q(\clock_inst.hour_tile.e0[50] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[51]$_DFFE_PP_  (.CLK(clknet_4_10__leaf_clk),
    .RESET_B(net732),
    .D(_00144_),
    .Q_N(_07877_),
    .Q(\clock_inst.hour_tile.e0[51] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[52]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net733),
    .D(_00145_),
    .Q_N(_07876_),
    .Q(\clock_inst.hour_tile.e0[52] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[53]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net734),
    .D(_00146_),
    .Q_N(_07875_),
    .Q(\clock_inst.hour_tile.e0[53] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[5]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net735),
    .D(_00147_),
    .Q_N(_07874_),
    .Q(\clock_inst.hour_tile.e0[5] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[6]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net736),
    .D(_00148_),
    .Q_N(_07873_),
    .Q(\clock_inst.hour_tile.e0[6] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[7]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net737),
    .D(_00149_),
    .Q_N(_07872_),
    .Q(\clock_inst.hour_tile.e0[7] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[8]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net738),
    .D(_00150_),
    .Q_N(_07871_),
    .Q(\clock_inst.hour_tile.e0[8] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e0[9]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net739),
    .D(_00151_),
    .Q_N(_07870_),
    .Q(\clock_inst.hour_tile.e0[9] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net740),
    .D(_00152_),
    .Q_N(_07869_),
    .Q(\clock_inst.hour_tile.e[0] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[10]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net741),
    .D(_00153_),
    .Q_N(_07868_),
    .Q(\clock_inst.hour_tile.e[10] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[11]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net742),
    .D(_00154_),
    .Q_N(_07867_),
    .Q(\clock_inst.hour_tile.e[11] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[12]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net743),
    .D(_00155_),
    .Q_N(_07866_),
    .Q(\clock_inst.hour_tile.e[12] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[13]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net744),
    .D(_00156_),
    .Q_N(_07865_),
    .Q(\clock_inst.hour_tile.e[13] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[14]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net745),
    .D(_00157_),
    .Q_N(_07864_),
    .Q(\clock_inst.hour_tile.e[14] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[15]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net746),
    .D(_00158_),
    .Q_N(_07863_),
    .Q(\clock_inst.hour_tile.e[15] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[16]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net747),
    .D(_00159_),
    .Q_N(_07862_),
    .Q(\clock_inst.hour_tile.e[16] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[17]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net748),
    .D(_00160_),
    .Q_N(_07861_),
    .Q(\clock_inst.hour_tile.e[17] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[18]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net749),
    .D(_00161_),
    .Q_N(_07860_),
    .Q(\clock_inst.hour_tile.e[18] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[19]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net750),
    .D(_00162_),
    .Q_N(_07859_),
    .Q(\clock_inst.hour_tile.e[19] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net751),
    .D(_00163_),
    .Q_N(_07858_),
    .Q(\clock_inst.hour_tile.e[1] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[20]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net752),
    .D(_00164_),
    .Q_N(_07857_),
    .Q(\clock_inst.hour_tile.e[20] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[21]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net753),
    .D(_00165_),
    .Q_N(_07856_),
    .Q(\clock_inst.hour_tile.e[21] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[22]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net754),
    .D(_00166_),
    .Q_N(_07855_),
    .Q(\clock_inst.hour_tile.e[22] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[23]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net755),
    .D(_00167_),
    .Q_N(_07854_),
    .Q(\clock_inst.hour_tile.e[23] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[24]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net756),
    .D(_00168_),
    .Q_N(_07853_),
    .Q(\clock_inst.hour_tile.e[24] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[25]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net757),
    .D(_00169_),
    .Q_N(_07852_),
    .Q(\clock_inst.hour_tile.e[25] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[26]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net758),
    .D(_00170_),
    .Q_N(_07851_),
    .Q(\clock_inst.hour_tile.e[26] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[27]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net759),
    .D(_00171_),
    .Q_N(_07850_),
    .Q(\clock_inst.hour_tile.e[27] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[28]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net760),
    .D(_00172_),
    .Q_N(_07849_),
    .Q(\clock_inst.hour_tile.e[28] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[29]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net761),
    .D(_00173_),
    .Q_N(_07848_),
    .Q(\clock_inst.hour_tile.e[29] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net762),
    .D(_00174_),
    .Q_N(_07847_),
    .Q(\clock_inst.hour_tile.e[2] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[30]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net763),
    .D(_00175_),
    .Q_N(_07846_),
    .Q(\clock_inst.hour_tile.e[30] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[31]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net764),
    .D(_00176_),
    .Q_N(_07845_),
    .Q(\clock_inst.hour_tile.e[31] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[32]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net765),
    .D(_00177_),
    .Q_N(_07844_),
    .Q(\clock_inst.hour_tile.e[32] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[33]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net766),
    .D(_00178_),
    .Q_N(_07843_),
    .Q(\clock_inst.hour_tile.e[33] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[34]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net767),
    .D(_00179_),
    .Q_N(_07842_),
    .Q(\clock_inst.hour_tile.e[34] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[35]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net768),
    .D(_00180_),
    .Q_N(_07841_),
    .Q(\clock_inst.hour_tile.e[35] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[36]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net769),
    .D(_00181_),
    .Q_N(_07840_),
    .Q(\clock_inst.hour_tile.e[36] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[37]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net770),
    .D(_00182_),
    .Q_N(_07839_),
    .Q(\clock_inst.hour_tile.e[37] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[38]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net771),
    .D(_00183_),
    .Q_N(_07838_),
    .Q(\clock_inst.hour_tile.e[38] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[39]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net772),
    .D(_00184_),
    .Q_N(_07837_),
    .Q(\clock_inst.hour_tile.e[39] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[3]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net773),
    .D(_00185_),
    .Q_N(_07836_),
    .Q(\clock_inst.hour_tile.e[3] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[40]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net774),
    .D(_00186_),
    .Q_N(_07835_),
    .Q(\clock_inst.hour_tile.e[40] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[41]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net775),
    .D(_00187_),
    .Q_N(_07834_),
    .Q(\clock_inst.hour_tile.e[41] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[42]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net776),
    .D(_00188_),
    .Q_N(_07833_),
    .Q(\clock_inst.hour_tile.e[42] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[43]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net777),
    .D(_00189_),
    .Q_N(_07832_),
    .Q(\clock_inst.hour_tile.e[43] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[44]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net778),
    .D(_00190_),
    .Q_N(_07831_),
    .Q(\clock_inst.hour_tile.e[44] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[45]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net779),
    .D(_00191_),
    .Q_N(_07830_),
    .Q(\clock_inst.hour_tile.e[45] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[46]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net780),
    .D(_00192_),
    .Q_N(_07829_),
    .Q(\clock_inst.hour_tile.e[46] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[47]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net781),
    .D(_00193_),
    .Q_N(_07828_),
    .Q(\clock_inst.hour_tile.e[47] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[48]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net782),
    .D(_00194_),
    .Q_N(_07827_),
    .Q(\clock_inst.hour_tile.e[48] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[49]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net783),
    .D(_00195_),
    .Q_N(_07826_),
    .Q(\clock_inst.hour_tile.e[49] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[4]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net784),
    .D(_00196_),
    .Q_N(_07825_),
    .Q(\clock_inst.hour_tile.e[4] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[50]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net785),
    .D(_00197_),
    .Q_N(_07824_),
    .Q(\clock_inst.hour_tile.e[50] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[51]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net786),
    .D(_00198_),
    .Q_N(_07823_),
    .Q(\clock_inst.hour_tile.e[51] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[52]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net787),
    .D(_00199_),
    .Q_N(_07822_),
    .Q(\clock_inst.hour_tile.e[52] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[53]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net788),
    .D(_00200_),
    .Q_N(_07821_),
    .Q(\clock_inst.hour_tile.e[53] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net789),
    .D(_00201_),
    .Q_N(_07820_),
    .Q(\clock_inst.hour_tile.e[5] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[6]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net790),
    .D(_00202_),
    .Q_N(_07819_),
    .Q(\clock_inst.hour_tile.e[6] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net791),
    .D(_00203_),
    .Q_N(_07818_),
    .Q(\clock_inst.hour_tile.e[7] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[8]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net792),
    .D(_00204_),
    .Q_N(_07817_),
    .Q(\clock_inst.hour_tile.e[8] ));
 sg13g2_dfrbp_1 \clock_inst.hour_tile.e[9]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net793),
    .D(_00205_),
    .Q_N(_07816_),
    .Q(\clock_inst.hour_tile.e[9] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[0]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net794),
    .D(_00206_),
    .Q_N(_07815_),
    .Q(\clock_inst.min_a[0] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[17]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net795),
    .D(_00207_),
    .Q_N(_07814_),
    .Q(\clock_inst.min_a[10] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[18]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net796),
    .D(_00208_),
    .Q_N(_07813_),
    .Q(\clock_inst.min_a[18] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[19]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net797),
    .D(_00209_),
    .Q_N(_07812_),
    .Q(\clock_inst.min_a[19] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[1]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net798),
    .D(_00210_),
    .Q_N(_07811_),
    .Q(\clock_inst.min_a[1] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[20]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net799),
    .D(_00211_),
    .Q_N(_07810_),
    .Q(\clock_inst.min_a[20] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[21]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net800),
    .D(_00212_),
    .Q_N(_07809_),
    .Q(\clock_inst.min_a[21] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[22]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net801),
    .D(_00213_),
    .Q_N(_07808_),
    .Q(\clock_inst.min_a[22] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[23]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net802),
    .D(_00214_),
    .Q_N(_07807_),
    .Q(\clock_inst.min_a[23] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[2]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net803),
    .D(_00215_),
    .Q_N(_07806_),
    .Q(\clock_inst.min_a[2] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[35]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net804),
    .D(_00216_),
    .Q_N(_07805_),
    .Q(\clock_inst.min_a[24] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[36]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net805),
    .D(_00217_),
    .Q_N(_07804_),
    .Q(\clock_inst.min_a[36] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[37]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net806),
    .D(_00218_),
    .Q_N(_07803_),
    .Q(\clock_inst.min_a[37] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[38]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net807),
    .D(_00219_),
    .Q_N(_07802_),
    .Q(\clock_inst.min_a[38] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[39]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net808),
    .D(_00220_),
    .Q_N(_07801_),
    .Q(\clock_inst.min_a[39] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[3]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net809),
    .D(_00221_),
    .Q_N(_07800_),
    .Q(\clock_inst.min_a[3] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[40]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net810),
    .D(_00222_),
    .Q_N(_07799_),
    .Q(\clock_inst.min_a[40] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[41]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net811),
    .D(_00223_),
    .Q_N(_07798_),
    .Q(\clock_inst.min_a[41] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[42]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net812),
    .D(_00224_),
    .Q_N(_07797_),
    .Q(\clock_inst.min_a[42] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[43]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net813),
    .D(_00225_),
    .Q_N(_07796_),
    .Q(\clock_inst.min_a[43] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[44]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net814),
    .D(_00226_),
    .Q_N(_07795_),
    .Q(\clock_inst.min_a[44] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[4]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net815),
    .D(_00227_),
    .Q_N(_07794_),
    .Q(\clock_inst.min_a[4] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[52]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net816),
    .D(_00228_),
    .Q_N(_07793_),
    .Q(\clock_inst.min_a[45] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[5]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net817),
    .D(_00229_),
    .Q_N(_07792_),
    .Q(\clock_inst.min_a[5] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[6]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net818),
    .D(_00230_),
    .Q_N(_07791_),
    .Q(\clock_inst.min_a[6] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net819),
    .D(_00231_),
    .Q_N(_07790_),
    .Q(\clock_inst.min_a[7] ));
 sg13g2_dfrbp_1 \clock_inst.min_a[8]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net820),
    .D(_00232_),
    .Q_N(_07789_),
    .Q(\clock_inst.min_a[8] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[0]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net821),
    .D(_00233_),
    .Q_N(_07788_),
    .Q(\clock_inst.min_b[0] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[17]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net822),
    .D(_00234_),
    .Q_N(_07787_),
    .Q(\clock_inst.min_b[10] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[19]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net823),
    .D(_00235_),
    .Q_N(_07786_),
    .Q(\clock_inst.min_b[19] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[1]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net824),
    .D(_00236_),
    .Q_N(_07785_),
    .Q(\clock_inst.min_b[1] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[20]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net825),
    .D(_00237_),
    .Q_N(_07784_),
    .Q(\clock_inst.min_b[20] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[21]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net826),
    .D(_00238_),
    .Q_N(_07783_),
    .Q(\clock_inst.min_b[21] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[22]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net827),
    .D(_00239_),
    .Q_N(_07782_),
    .Q(\clock_inst.min_b[22] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[23]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net828),
    .D(_00240_),
    .Q_N(_07781_),
    .Q(\clock_inst.min_b[23] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[2]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net829),
    .D(_00241_),
    .Q_N(_07780_),
    .Q(\clock_inst.min_b[2] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[35]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net830),
    .D(_00242_),
    .Q_N(_07779_),
    .Q(\clock_inst.min_b[24] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[36]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net831),
    .D(_00243_),
    .Q_N(_07778_),
    .Q(\clock_inst.min_b[36] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[37]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net832),
    .D(_00244_),
    .Q_N(_07777_),
    .Q(\clock_inst.min_b[37] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[38]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net833),
    .D(_00245_),
    .Q_N(_07776_),
    .Q(\clock_inst.min_b[38] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[39]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net834),
    .D(_00246_),
    .Q_N(_07775_),
    .Q(\clock_inst.min_b[39] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[3]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net835),
    .D(_00247_),
    .Q_N(_07774_),
    .Q(\clock_inst.min_b[3] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[40]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net836),
    .D(_00248_),
    .Q_N(_07773_),
    .Q(\clock_inst.min_b[40] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[41]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net837),
    .D(_00249_),
    .Q_N(_07772_),
    .Q(\clock_inst.min_b[41] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[42]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net838),
    .D(_00250_),
    .Q_N(_07771_),
    .Q(\clock_inst.min_b[42] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[43]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net839),
    .D(_00251_),
    .Q_N(_07770_),
    .Q(\clock_inst.min_b[43] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[44]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net840),
    .D(_00252_),
    .Q_N(_07769_),
    .Q(\clock_inst.min_b[44] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[4]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net841),
    .D(_00253_),
    .Q_N(_07768_),
    .Q(\clock_inst.min_b[4] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[5]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net842),
    .D(_00254_),
    .Q_N(_07767_),
    .Q(\clock_inst.min_b[5] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[6]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net843),
    .D(_00255_),
    .Q_N(_07766_),
    .Q(\clock_inst.min_b[6] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net844),
    .D(_00256_),
    .Q_N(_07765_),
    .Q(\clock_inst.min_b[7] ));
 sg13g2_dfrbp_1 \clock_inst.min_b[8]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net845),
    .D(_00257_),
    .Q_N(_07764_),
    .Q(\clock_inst.min_b[8] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[0]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net846),
    .D(_00258_),
    .Q_N(_07763_),
    .Q(\clock_inst.min_c[0] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[10]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net847),
    .D(_00259_),
    .Q_N(_07762_),
    .Q(\clock_inst.min_c[10] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net848),
    .D(_00260_),
    .Q_N(_07761_),
    .Q(\clock_inst.min_c[11] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[12]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net849),
    .D(_00261_),
    .Q_N(_07760_),
    .Q(\clock_inst.min_c[12] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[13]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net850),
    .D(_00262_),
    .Q_N(_07759_),
    .Q(\clock_inst.min_c[13] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[14]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net851),
    .D(_00263_),
    .Q_N(_07758_),
    .Q(\clock_inst.min_c[14] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[15]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net852),
    .D(_00264_),
    .Q_N(_07757_),
    .Q(\clock_inst.min_c[15] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[16]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net853),
    .D(_00265_),
    .Q_N(_07756_),
    .Q(\clock_inst.min_c[16] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[17]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net854),
    .D(_00266_),
    .Q_N(_07755_),
    .Q(\clock_inst.min_c[17] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[19]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net855),
    .D(_00267_),
    .Q_N(_07754_),
    .Q(\clock_inst.min_c[19] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[1]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net856),
    .D(_00268_),
    .Q_N(_07753_),
    .Q(\clock_inst.min_c[1] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[21]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net857),
    .D(_00269_),
    .Q_N(_07752_),
    .Q(\clock_inst.min_c[21] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[22]$_DFFE_PP_  (.CLK(clknet_4_0__leaf_clk),
    .RESET_B(net858),
    .D(_00270_),
    .Q_N(_07751_),
    .Q(\clock_inst.min_c[22] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[23]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net859),
    .D(_00271_),
    .Q_N(_07750_),
    .Q(\clock_inst.min_c[23] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[24]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net860),
    .D(_00272_),
    .Q_N(_07749_),
    .Q(\clock_inst.min_c[24] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[25]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net861),
    .D(_00273_),
    .Q_N(_07748_),
    .Q(\clock_inst.min_c[25] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[26]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net862),
    .D(_00274_),
    .Q_N(_07747_),
    .Q(\clock_inst.min_c[26] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[27]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net863),
    .D(_00275_),
    .Q_N(_07746_),
    .Q(\clock_inst.min_c[27] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[28]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net864),
    .D(_00276_),
    .Q_N(_07745_),
    .Q(\clock_inst.min_c[28] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[29]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net865),
    .D(_00277_),
    .Q_N(_07744_),
    .Q(\clock_inst.min_c[29] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net866),
    .D(_00278_),
    .Q_N(_07743_),
    .Q(\clock_inst.min_c[2] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[30]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net867),
    .D(_00279_),
    .Q_N(_07742_),
    .Q(\clock_inst.min_c[30] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[31]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net868),
    .D(_00280_),
    .Q_N(_07741_),
    .Q(\clock_inst.min_c[31] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[32]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net869),
    .D(_00281_),
    .Q_N(_07740_),
    .Q(\clock_inst.min_c[32] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[35]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net870),
    .D(_00282_),
    .Q_N(_07739_),
    .Q(\clock_inst.min_c[33] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[36]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net871),
    .D(_00283_),
    .Q_N(_07738_),
    .Q(\clock_inst.min_c[36] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[37]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net872),
    .D(_00284_),
    .Q_N(_07737_),
    .Q(\clock_inst.min_c[37] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[38]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net873),
    .D(_00285_),
    .Q_N(_07736_),
    .Q(\clock_inst.min_c[38] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[39]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net874),
    .D(_00286_),
    .Q_N(_07735_),
    .Q(\clock_inst.min_c[39] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[3]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net875),
    .D(_00287_),
    .Q_N(_07734_),
    .Q(\clock_inst.min_c[3] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[40]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net876),
    .D(_00288_),
    .Q_N(_07733_),
    .Q(\clock_inst.min_c[40] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[41]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net877),
    .D(_00289_),
    .Q_N(_07732_),
    .Q(\clock_inst.min_c[41] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[42]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net878),
    .D(_00290_),
    .Q_N(_07731_),
    .Q(\clock_inst.min_c[42] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[43]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net879),
    .D(_00291_),
    .Q_N(_07730_),
    .Q(\clock_inst.min_c[43] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[44]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net880),
    .D(_00292_),
    .Q_N(_07729_),
    .Q(\clock_inst.min_c[44] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[45]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net881),
    .D(_00293_),
    .Q_N(_07728_),
    .Q(\clock_inst.min_c[45] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[46]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net882),
    .D(_00294_),
    .Q_N(_07727_),
    .Q(\clock_inst.min_c[46] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[47]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net883),
    .D(_00295_),
    .Q_N(_07726_),
    .Q(\clock_inst.min_c[47] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[48]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net884),
    .D(_00296_),
    .Q_N(_07725_),
    .Q(\clock_inst.min_c[48] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[49]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net885),
    .D(_00297_),
    .Q_N(_07724_),
    .Q(\clock_inst.min_c[49] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[4]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net886),
    .D(_00298_),
    .Q_N(_07723_),
    .Q(\clock_inst.min_c[4] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[50]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net887),
    .D(_00299_),
    .Q_N(_07722_),
    .Q(\clock_inst.min_c[50] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[51]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net888),
    .D(_00300_),
    .Q_N(_07721_),
    .Q(\clock_inst.min_c[51] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[52]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net889),
    .D(_00301_),
    .Q_N(_07720_),
    .Q(\clock_inst.min_c[52] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[53]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net890),
    .D(_00302_),
    .Q_N(_07719_),
    .Q(\clock_inst.min_c[53] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net891),
    .D(_00303_),
    .Q_N(_07718_),
    .Q(\clock_inst.min_c[5] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[6]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net892),
    .D(_00304_),
    .Q_N(_07717_),
    .Q(\clock_inst.min_c[6] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[7]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net893),
    .D(_00305_),
    .Q_N(_07716_),
    .Q(\clock_inst.min_c[7] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[8]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net894),
    .D(_00306_),
    .Q_N(_07715_),
    .Q(\clock_inst.min_c[8] ));
 sg13g2_dfrbp_1 \clock_inst.min_c[9]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net895),
    .D(_00307_),
    .Q_N(_07714_),
    .Q(\clock_inst.min_c[9] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[0]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net896),
    .D(_00308_),
    .Q_N(_07713_),
    .Q(\clock_inst.min_tile.e0[0] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[10]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net897),
    .D(_00309_),
    .Q_N(_07712_),
    .Q(\clock_inst.min_tile.e0[10] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[11]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net898),
    .D(_00310_),
    .Q_N(_07711_),
    .Q(\clock_inst.min_tile.e0[11] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[12]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net899),
    .D(_00311_),
    .Q_N(_07710_),
    .Q(\clock_inst.min_tile.e0[12] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[13]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net900),
    .D(_00312_),
    .Q_N(_07709_),
    .Q(\clock_inst.min_tile.e0[13] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[14]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net901),
    .D(_00313_),
    .Q_N(_07708_),
    .Q(\clock_inst.min_tile.e0[14] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[15]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net902),
    .D(_00314_),
    .Q_N(_07707_),
    .Q(\clock_inst.min_tile.e0[15] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[16]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net903),
    .D(_00315_),
    .Q_N(_07706_),
    .Q(\clock_inst.min_tile.e0[16] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[17]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net904),
    .D(_00316_),
    .Q_N(_07705_),
    .Q(\clock_inst.min_tile.e0[17] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[18]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net905),
    .D(_00317_),
    .Q_N(_07704_),
    .Q(\clock_inst.min_tile.e0[18] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[19]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net906),
    .D(_00318_),
    .Q_N(_07703_),
    .Q(\clock_inst.min_tile.e0[19] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[1]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net907),
    .D(_00319_),
    .Q_N(_07702_),
    .Q(\clock_inst.min_tile.e0[1] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[20]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net908),
    .D(_00320_),
    .Q_N(_07701_),
    .Q(\clock_inst.min_tile.e0[20] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[21]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net909),
    .D(_00321_),
    .Q_N(_07700_),
    .Q(\clock_inst.min_tile.e0[21] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[22]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net910),
    .D(_00322_),
    .Q_N(_07699_),
    .Q(\clock_inst.min_tile.e0[22] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[23]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net911),
    .D(_00323_),
    .Q_N(_07698_),
    .Q(\clock_inst.min_tile.e0[23] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[24]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net912),
    .D(_00324_),
    .Q_N(_07697_),
    .Q(\clock_inst.min_tile.e0[24] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[25]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net913),
    .D(_00325_),
    .Q_N(_07696_),
    .Q(\clock_inst.min_tile.e0[25] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[26]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net914),
    .D(_00326_),
    .Q_N(_07695_),
    .Q(\clock_inst.min_tile.e0[26] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[27]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net915),
    .D(_00327_),
    .Q_N(_07694_),
    .Q(\clock_inst.min_tile.e0[27] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[28]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net916),
    .D(_00328_),
    .Q_N(_07693_),
    .Q(\clock_inst.min_tile.e0[28] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[29]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net917),
    .D(_00329_),
    .Q_N(_07692_),
    .Q(\clock_inst.min_tile.e0[29] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[2]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net918),
    .D(_00330_),
    .Q_N(_07691_),
    .Q(\clock_inst.min_tile.e0[2] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[30]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net919),
    .D(_00331_),
    .Q_N(_07690_),
    .Q(\clock_inst.min_tile.e0[30] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[31]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net920),
    .D(_00332_),
    .Q_N(_07689_),
    .Q(\clock_inst.min_tile.e0[31] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[32]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net921),
    .D(_00333_),
    .Q_N(_07688_),
    .Q(\clock_inst.min_tile.e0[32] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[33]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net922),
    .D(_00334_),
    .Q_N(_07687_),
    .Q(\clock_inst.min_tile.e0[33] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[34]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net923),
    .D(_00335_),
    .Q_N(_07686_),
    .Q(\clock_inst.min_tile.e0[34] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[35]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net924),
    .D(_00336_),
    .Q_N(_07685_),
    .Q(\clock_inst.min_tile.e0[35] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[36]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net925),
    .D(_00337_),
    .Q_N(_07684_),
    .Q(\clock_inst.min_tile.e0[36] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[37]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net926),
    .D(_00338_),
    .Q_N(_07683_),
    .Q(\clock_inst.min_tile.e0[37] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[38]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net927),
    .D(_00339_),
    .Q_N(_07682_),
    .Q(\clock_inst.min_tile.e0[38] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[39]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net928),
    .D(_00340_),
    .Q_N(_07681_),
    .Q(\clock_inst.min_tile.e0[39] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[3]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net929),
    .D(_00341_),
    .Q_N(_07680_),
    .Q(\clock_inst.min_tile.e0[3] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[40]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net930),
    .D(_00342_),
    .Q_N(_07679_),
    .Q(\clock_inst.min_tile.e0[40] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[41]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net931),
    .D(_00343_),
    .Q_N(_07678_),
    .Q(\clock_inst.min_tile.e0[41] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[42]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net932),
    .D(_00344_),
    .Q_N(_07677_),
    .Q(\clock_inst.min_tile.e0[42] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[43]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net933),
    .D(_00345_),
    .Q_N(_07676_),
    .Q(\clock_inst.min_tile.e0[43] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[44]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net934),
    .D(_00346_),
    .Q_N(_07675_),
    .Q(\clock_inst.min_tile.e0[44] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[45]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net935),
    .D(_00347_),
    .Q_N(_07674_),
    .Q(\clock_inst.min_tile.e0[45] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[46]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net936),
    .D(_00348_),
    .Q_N(_07673_),
    .Q(\clock_inst.min_tile.e0[46] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[47]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net937),
    .D(_00349_),
    .Q_N(_07672_),
    .Q(\clock_inst.min_tile.e0[47] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[48]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net938),
    .D(_00350_),
    .Q_N(_07671_),
    .Q(\clock_inst.min_tile.e0[48] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[49]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net939),
    .D(_00351_),
    .Q_N(_07670_),
    .Q(\clock_inst.min_tile.e0[49] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[4]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net940),
    .D(_00352_),
    .Q_N(_07669_),
    .Q(\clock_inst.min_tile.e0[4] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[50]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net941),
    .D(_00353_),
    .Q_N(_07668_),
    .Q(\clock_inst.min_tile.e0[50] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[51]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net942),
    .D(_00354_),
    .Q_N(_07667_),
    .Q(\clock_inst.min_tile.e0[51] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[52]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net943),
    .D(_00355_),
    .Q_N(_07666_),
    .Q(\clock_inst.min_tile.e0[52] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[53]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net944),
    .D(_00356_),
    .Q_N(_07665_),
    .Q(\clock_inst.min_tile.e0[53] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[5]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net945),
    .D(_00357_),
    .Q_N(_07664_),
    .Q(\clock_inst.min_tile.e0[5] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[6]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net946),
    .D(_00358_),
    .Q_N(_07663_),
    .Q(\clock_inst.min_tile.e0[6] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[7]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net947),
    .D(_00359_),
    .Q_N(_07662_),
    .Q(\clock_inst.min_tile.e0[7] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[8]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net948),
    .D(_00360_),
    .Q_N(_07661_),
    .Q(\clock_inst.min_tile.e0[8] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e0[9]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net949),
    .D(_00361_),
    .Q_N(_07660_),
    .Q(\clock_inst.min_tile.e0[9] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[0]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net950),
    .D(_00362_),
    .Q_N(_07659_),
    .Q(\clock_inst.min_tile.e[0] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[10]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net951),
    .D(_00363_),
    .Q_N(_07658_),
    .Q(\clock_inst.min_tile.e[10] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[11]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net952),
    .D(_00364_),
    .Q_N(_07657_),
    .Q(\clock_inst.min_tile.e[11] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[12]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net953),
    .D(_00365_),
    .Q_N(_07656_),
    .Q(\clock_inst.min_tile.e[12] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[13]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net954),
    .D(_00366_),
    .Q_N(_07655_),
    .Q(\clock_inst.min_tile.e[13] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[14]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net955),
    .D(_00367_),
    .Q_N(_07654_),
    .Q(\clock_inst.min_tile.e[14] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[15]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net956),
    .D(_00368_),
    .Q_N(_07653_),
    .Q(\clock_inst.min_tile.e[15] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[16]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net957),
    .D(_00369_),
    .Q_N(_07652_),
    .Q(\clock_inst.min_tile.e[16] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[17]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net958),
    .D(_00370_),
    .Q_N(_07651_),
    .Q(\clock_inst.min_tile.e[17] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[18]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net959),
    .D(_00371_),
    .Q_N(_07650_),
    .Q(\clock_inst.min_tile.e[18] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[19]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net960),
    .D(_00372_),
    .Q_N(_07649_),
    .Q(\clock_inst.min_tile.e[19] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[1]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net961),
    .D(_00373_),
    .Q_N(_07648_),
    .Q(\clock_inst.min_tile.e[1] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[20]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net962),
    .D(_00374_),
    .Q_N(_07647_),
    .Q(\clock_inst.min_tile.e[20] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[21]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net963),
    .D(_00375_),
    .Q_N(_07646_),
    .Q(\clock_inst.min_tile.e[21] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[22]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net964),
    .D(_00376_),
    .Q_N(_07645_),
    .Q(\clock_inst.min_tile.e[22] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[23]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net965),
    .D(_00377_),
    .Q_N(_07644_),
    .Q(\clock_inst.min_tile.e[23] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[24]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net966),
    .D(_00378_),
    .Q_N(_07643_),
    .Q(\clock_inst.min_tile.e[24] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[25]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net967),
    .D(_00379_),
    .Q_N(_07642_),
    .Q(\clock_inst.min_tile.e[25] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[26]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net968),
    .D(_00380_),
    .Q_N(_07641_),
    .Q(\clock_inst.min_tile.e[26] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[27]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net969),
    .D(_00381_),
    .Q_N(_07640_),
    .Q(\clock_inst.min_tile.e[27] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[28]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net970),
    .D(_00382_),
    .Q_N(_07639_),
    .Q(\clock_inst.min_tile.e[28] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[29]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net971),
    .D(_00383_),
    .Q_N(_07638_),
    .Q(\clock_inst.min_tile.e[29] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[2]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net972),
    .D(_00384_),
    .Q_N(_07637_),
    .Q(\clock_inst.min_tile.e[2] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[30]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net973),
    .D(_00385_),
    .Q_N(_07636_),
    .Q(\clock_inst.min_tile.e[30] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[31]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net974),
    .D(_00386_),
    .Q_N(_07635_),
    .Q(\clock_inst.min_tile.e[31] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[32]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net975),
    .D(_00387_),
    .Q_N(_07634_),
    .Q(\clock_inst.min_tile.e[32] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[33]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net976),
    .D(_00388_),
    .Q_N(_07633_),
    .Q(\clock_inst.min_tile.e[33] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[34]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net977),
    .D(_00389_),
    .Q_N(_07632_),
    .Q(\clock_inst.min_tile.e[34] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[35]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net978),
    .D(_00390_),
    .Q_N(_07631_),
    .Q(\clock_inst.min_tile.e[35] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[36]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net979),
    .D(_00391_),
    .Q_N(_07630_),
    .Q(\clock_inst.min_tile.e[36] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[37]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net980),
    .D(_00392_),
    .Q_N(_07629_),
    .Q(\clock_inst.min_tile.e[37] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[38]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net981),
    .D(_00393_),
    .Q_N(_07628_),
    .Q(\clock_inst.min_tile.e[38] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[39]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net982),
    .D(_00394_),
    .Q_N(_07627_),
    .Q(\clock_inst.min_tile.e[39] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[3]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net983),
    .D(_00395_),
    .Q_N(_07626_),
    .Q(\clock_inst.min_tile.e[3] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[40]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net984),
    .D(_00396_),
    .Q_N(_07625_),
    .Q(\clock_inst.min_tile.e[40] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[41]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net985),
    .D(_00397_),
    .Q_N(_07624_),
    .Q(\clock_inst.min_tile.e[41] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[42]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net986),
    .D(_00398_),
    .Q_N(_07623_),
    .Q(\clock_inst.min_tile.e[42] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[43]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net987),
    .D(_00399_),
    .Q_N(_07622_),
    .Q(\clock_inst.min_tile.e[43] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[44]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net988),
    .D(_00400_),
    .Q_N(_07621_),
    .Q(\clock_inst.min_tile.e[44] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[45]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net989),
    .D(_00401_),
    .Q_N(_07620_),
    .Q(\clock_inst.min_tile.e[45] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[46]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net990),
    .D(_00402_),
    .Q_N(_07619_),
    .Q(\clock_inst.min_tile.e[46] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[47]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net991),
    .D(_00403_),
    .Q_N(_07618_),
    .Q(\clock_inst.min_tile.e[47] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[48]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net992),
    .D(_00404_),
    .Q_N(_07617_),
    .Q(\clock_inst.min_tile.e[48] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[49]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net993),
    .D(_00405_),
    .Q_N(_07616_),
    .Q(\clock_inst.min_tile.e[49] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[4]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net994),
    .D(_00406_),
    .Q_N(_07615_),
    .Q(\clock_inst.min_tile.e[4] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[50]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net995),
    .D(_00407_),
    .Q_N(_07614_),
    .Q(\clock_inst.min_tile.e[50] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[51]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net996),
    .D(_00408_),
    .Q_N(_07613_),
    .Q(\clock_inst.min_tile.e[51] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[52]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net997),
    .D(_00409_),
    .Q_N(_07612_),
    .Q(\clock_inst.min_tile.e[52] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[53]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net998),
    .D(_00410_),
    .Q_N(_07611_),
    .Q(\clock_inst.min_tile.e[53] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[5]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net999),
    .D(_00411_),
    .Q_N(_07610_),
    .Q(\clock_inst.min_tile.e[5] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[6]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1000),
    .D(_00412_),
    .Q_N(_07609_),
    .Q(\clock_inst.min_tile.e[6] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[7]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1001),
    .D(_00413_),
    .Q_N(_07608_),
    .Q(\clock_inst.min_tile.e[7] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[8]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1002),
    .D(_00414_),
    .Q_N(_07607_),
    .Q(\clock_inst.min_tile.e[8] ));
 sg13g2_dfrbp_1 \clock_inst.min_tile.e[9]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1003),
    .D(_00415_),
    .Q_N(_07606_),
    .Q(\clock_inst.min_tile.e[9] ));
 sg13g2_dfrbp_1 \clock_inst.minute[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1004),
    .D(_00416_),
    .Q_N(_00002_),
    .Q(\clock_inst.minute[0] ));
 sg13g2_dfrbp_1 \clock_inst.minute[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1005),
    .D(_00417_),
    .Q_N(_07605_),
    .Q(\clock_inst.minute[1] ));
 sg13g2_dfrbp_1 \clock_inst.minute[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1006),
    .D(_00418_),
    .Q_N(_07604_),
    .Q(\clock_inst.minute[2] ));
 sg13g2_dfrbp_1 \clock_inst.minute[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1007),
    .D(_00419_),
    .Q_N(_07603_),
    .Q(\clock_inst.minute[3] ));
 sg13g2_dfrbp_1 \clock_inst.minute[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1008),
    .D(_00420_),
    .Q_N(_07602_),
    .Q(\clock_inst.minute[4] ));
 sg13g2_dfrbp_1 \clock_inst.minute[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1009),
    .D(_00421_),
    .Q_N(_07601_),
    .Q(\clock_inst.minute[5] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1010),
    .D(_00422_),
    .Q_N(_07600_),
    .Q(\clock_inst.sec_a[0] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[17]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1011),
    .D(_00423_),
    .Q_N(_07599_),
    .Q(\clock_inst.sec_a[10] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[18]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1012),
    .D(_00424_),
    .Q_N(_07598_),
    .Q(\clock_inst.sec_a[18] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[19]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1013),
    .D(_00425_),
    .Q_N(_07597_),
    .Q(\clock_inst.sec_a[19] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1014),
    .D(_00426_),
    .Q_N(_07596_),
    .Q(\clock_inst.sec_a[1] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[20]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1015),
    .D(_00427_),
    .Q_N(_07595_),
    .Q(\clock_inst.sec_a[20] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1016),
    .D(_00428_),
    .Q_N(_07594_),
    .Q(\clock_inst.sec_a[2] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[35]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1017),
    .D(_00429_),
    .Q_N(_07593_),
    .Q(\clock_inst.sec_a[21] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[36]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1018),
    .D(_00430_),
    .Q_N(_07592_),
    .Q(\clock_inst.sec_a[36] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[37]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1019),
    .D(_00431_),
    .Q_N(_07591_),
    .Q(\clock_inst.sec_a[37] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[38]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1020),
    .D(_00432_),
    .Q_N(_07590_),
    .Q(\clock_inst.sec_a[38] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[39]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1021),
    .D(_00433_),
    .Q_N(_07589_),
    .Q(\clock_inst.sec_a[39] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1022),
    .D(_00434_),
    .Q_N(_07588_),
    .Q(\clock_inst.sec_a[3] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[40]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1023),
    .D(_00435_),
    .Q_N(_07587_),
    .Q(\clock_inst.sec_a[40] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[41]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1024),
    .D(_00436_),
    .Q_N(_07586_),
    .Q(\clock_inst.sec_a[41] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[42]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1025),
    .D(_00437_),
    .Q_N(_07585_),
    .Q(\clock_inst.sec_a[42] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[43]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1026),
    .D(_00438_),
    .Q_N(_07584_),
    .Q(\clock_inst.sec_a[43] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1027),
    .D(_00439_),
    .Q_N(_07583_),
    .Q(\clock_inst.sec_a[4] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[52]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1028),
    .D(_00440_),
    .Q_N(_07582_),
    .Q(\clock_inst.sec_a[44] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[5]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1029),
    .D(_00441_),
    .Q_N(_07581_),
    .Q(\clock_inst.sec_a[5] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[6]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1030),
    .D(_00442_),
    .Q_N(_07580_),
    .Q(\clock_inst.sec_a[6] ));
 sg13g2_dfrbp_1 \clock_inst.sec_a[7]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1031),
    .D(_00443_),
    .Q_N(_07579_),
    .Q(\clock_inst.sec_a[7] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1032),
    .D(_00444_),
    .Q_N(_07578_),
    .Q(\clock_inst.sec_b[0] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[17]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1033),
    .D(_00445_),
    .Q_N(_07577_),
    .Q(\clock_inst.sec_b[10] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[19]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1034),
    .D(_00446_),
    .Q_N(_07576_),
    .Q(\clock_inst.sec_b[19] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1035),
    .D(_00447_),
    .Q_N(_07575_),
    .Q(\clock_inst.sec_b[1] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[20]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1036),
    .D(_00448_),
    .Q_N(_07574_),
    .Q(\clock_inst.sec_b[20] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[2]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1037),
    .D(_00449_),
    .Q_N(_07573_),
    .Q(\clock_inst.sec_b[2] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[35]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1038),
    .D(_00450_),
    .Q_N(_07572_),
    .Q(\clock_inst.sec_b[21] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[36]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1039),
    .D(_00451_),
    .Q_N(_07571_),
    .Q(\clock_inst.sec_b[36] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[37]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1040),
    .D(_00452_),
    .Q_N(_07570_),
    .Q(\clock_inst.sec_b[37] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[38]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1041),
    .D(_00453_),
    .Q_N(_07569_),
    .Q(\clock_inst.sec_b[38] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[39]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1042),
    .D(_00454_),
    .Q_N(_07568_),
    .Q(\clock_inst.sec_b[39] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[3]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1043),
    .D(_00455_),
    .Q_N(_07567_),
    .Q(\clock_inst.sec_b[3] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[40]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1044),
    .D(_00456_),
    .Q_N(_07566_),
    .Q(\clock_inst.sec_b[40] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[41]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1045),
    .D(_00457_),
    .Q_N(_07565_),
    .Q(\clock_inst.sec_b[41] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[42]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1046),
    .D(_00458_),
    .Q_N(_07564_),
    .Q(\clock_inst.sec_b[42] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[43]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1047),
    .D(_00459_),
    .Q_N(_07563_),
    .Q(\clock_inst.sec_b[43] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[4]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1048),
    .D(_00460_),
    .Q_N(_07562_),
    .Q(\clock_inst.sec_b[4] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[5]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1049),
    .D(_00461_),
    .Q_N(_07561_),
    .Q(\clock_inst.sec_b[5] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1050),
    .D(_00462_),
    .Q_N(_07560_),
    .Q(\clock_inst.sec_b[6] ));
 sg13g2_dfrbp_1 \clock_inst.sec_b[7]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1051),
    .D(_00463_),
    .Q_N(_07559_),
    .Q(\clock_inst.sec_b[7] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1052),
    .D(_00464_),
    .Q_N(_07558_),
    .Q(\clock_inst.sec_c[0] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[10]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1053),
    .D(_00465_),
    .Q_N(_07557_),
    .Q(\clock_inst.sec_c[10] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[11]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1054),
    .D(_00466_),
    .Q_N(_07556_),
    .Q(\clock_inst.sec_c[11] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[12]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1055),
    .D(_00467_),
    .Q_N(_07555_),
    .Q(\clock_inst.sec_c[12] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[13]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1056),
    .D(_00468_),
    .Q_N(_07554_),
    .Q(\clock_inst.sec_c[13] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[14]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1057),
    .D(_00469_),
    .Q_N(_07553_),
    .Q(\clock_inst.sec_c[14] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[15]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1058),
    .D(_00470_),
    .Q_N(_07552_),
    .Q(\clock_inst.sec_c[15] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[16]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1059),
    .D(_00471_),
    .Q_N(_07551_),
    .Q(\clock_inst.sec_c[16] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[17]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1060),
    .D(_00472_),
    .Q_N(_07550_),
    .Q(\clock_inst.sec_c[17] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[19]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1061),
    .D(_00473_),
    .Q_N(_07549_),
    .Q(\clock_inst.sec_c[19] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1062),
    .D(_00474_),
    .Q_N(_07548_),
    .Q(\clock_inst.sec_c[1] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[20]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1063),
    .D(_00475_),
    .Q_N(_07547_),
    .Q(\clock_inst.sec_c[20] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[21]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1064),
    .D(_00476_),
    .Q_N(_07546_),
    .Q(\clock_inst.sec_c[21] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[22]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1065),
    .D(_00477_),
    .Q_N(_07545_),
    .Q(\clock_inst.sec_c[22] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[23]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1066),
    .D(_00478_),
    .Q_N(_07544_),
    .Q(\clock_inst.sec_c[23] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[24]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1067),
    .D(_00479_),
    .Q_N(_07543_),
    .Q(\clock_inst.sec_c[24] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[25]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1068),
    .D(_00480_),
    .Q_N(_07542_),
    .Q(\clock_inst.sec_c[25] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[26]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1069),
    .D(_00481_),
    .Q_N(_07541_),
    .Q(\clock_inst.sec_c[26] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[27]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1070),
    .D(_00482_),
    .Q_N(_07540_),
    .Q(\clock_inst.sec_c[27] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[28]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1071),
    .D(_00483_),
    .Q_N(_07539_),
    .Q(\clock_inst.sec_c[28] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[29]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1072),
    .D(_00484_),
    .Q_N(_07538_),
    .Q(\clock_inst.sec_c[29] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[2]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1073),
    .D(_00485_),
    .Q_N(_07537_),
    .Q(\clock_inst.sec_c[2] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[35]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1074),
    .D(_00486_),
    .Q_N(_07536_),
    .Q(\clock_inst.sec_c[30] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[36]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1075),
    .D(_00487_),
    .Q_N(_07535_),
    .Q(\clock_inst.sec_c[36] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[37]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1076),
    .D(_00488_),
    .Q_N(_07534_),
    .Q(\clock_inst.sec_c[37] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[38]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1077),
    .D(_00489_),
    .Q_N(_07533_),
    .Q(\clock_inst.sec_c[38] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[39]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1078),
    .D(_00490_),
    .Q_N(_07532_),
    .Q(\clock_inst.sec_c[39] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[3]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1079),
    .D(_00491_),
    .Q_N(_07531_),
    .Q(\clock_inst.sec_c[3] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[40]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1080),
    .D(_00492_),
    .Q_N(_07530_),
    .Q(\clock_inst.sec_c[40] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[41]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1081),
    .D(_00493_),
    .Q_N(_07529_),
    .Q(\clock_inst.sec_c[41] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[42]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1082),
    .D(_00494_),
    .Q_N(_07528_),
    .Q(\clock_inst.sec_c[42] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[43]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1083),
    .D(_00495_),
    .Q_N(_07527_),
    .Q(\clock_inst.sec_c[43] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[44]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1084),
    .D(_00496_),
    .Q_N(_07526_),
    .Q(\clock_inst.sec_c[44] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[45]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1085),
    .D(_00497_),
    .Q_N(_07525_),
    .Q(\clock_inst.sec_c[45] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[46]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1086),
    .D(_00498_),
    .Q_N(_07524_),
    .Q(\clock_inst.sec_c[46] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[47]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1087),
    .D(_00499_),
    .Q_N(_07523_),
    .Q(\clock_inst.sec_c[47] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[48]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1088),
    .D(_00500_),
    .Q_N(_07522_),
    .Q(\clock_inst.sec_c[48] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[49]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1089),
    .D(_00501_),
    .Q_N(_07521_),
    .Q(\clock_inst.sec_c[49] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[4]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1090),
    .D(_00502_),
    .Q_N(_07520_),
    .Q(\clock_inst.sec_c[4] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[50]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1091),
    .D(_00503_),
    .Q_N(_07519_),
    .Q(\clock_inst.sec_c[50] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[51]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1092),
    .D(_00504_),
    .Q_N(_07518_),
    .Q(\clock_inst.sec_c[51] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[52]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1093),
    .D(_00505_),
    .Q_N(_07517_),
    .Q(\clock_inst.sec_c[52] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[53]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1094),
    .D(_00506_),
    .Q_N(_07516_),
    .Q(\clock_inst.sec_c[53] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[5]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1095),
    .D(_00507_),
    .Q_N(_07515_),
    .Q(\clock_inst.sec_c[5] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1096),
    .D(_00508_),
    .Q_N(_07514_),
    .Q(\clock_inst.sec_c[6] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[7]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1097),
    .D(_00509_),
    .Q_N(_07513_),
    .Q(\clock_inst.sec_c[7] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[8]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1098),
    .D(_00510_),
    .Q_N(_07512_),
    .Q(\clock_inst.sec_c[8] ));
 sg13g2_dfrbp_1 \clock_inst.sec_c[9]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1099),
    .D(_00511_),
    .Q_N(_07511_),
    .Q(\clock_inst.sec_c[9] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1100),
    .D(_00512_),
    .Q_N(_07510_),
    .Q(\clock_inst.sec_tile.e0[0] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[10]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1101),
    .D(_00513_),
    .Q_N(_07509_),
    .Q(\clock_inst.sec_tile.e0[10] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[11]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1102),
    .D(_00514_),
    .Q_N(_07508_),
    .Q(\clock_inst.sec_tile.e0[11] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[12]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1103),
    .D(_00515_),
    .Q_N(_07507_),
    .Q(\clock_inst.sec_tile.e0[12] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[13]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1104),
    .D(_00516_),
    .Q_N(_07506_),
    .Q(\clock_inst.sec_tile.e0[13] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[14]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1105),
    .D(_00517_),
    .Q_N(_07505_),
    .Q(\clock_inst.sec_tile.e0[14] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[15]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1106),
    .D(_00518_),
    .Q_N(_07504_),
    .Q(\clock_inst.sec_tile.e0[15] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[16]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1107),
    .D(_00519_),
    .Q_N(_07503_),
    .Q(\clock_inst.sec_tile.e0[16] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[17]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1108),
    .D(_00520_),
    .Q_N(_07502_),
    .Q(\clock_inst.sec_tile.e0[17] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[18]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1109),
    .D(_00521_),
    .Q_N(_07501_),
    .Q(\clock_inst.sec_tile.e0[18] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[19]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1110),
    .D(_00522_),
    .Q_N(_07500_),
    .Q(\clock_inst.sec_tile.e0[19] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[1]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1111),
    .D(_00523_),
    .Q_N(_07499_),
    .Q(\clock_inst.sec_tile.e0[1] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[20]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1112),
    .D(_00524_),
    .Q_N(_07498_),
    .Q(\clock_inst.sec_tile.e0[20] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[21]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1113),
    .D(_00525_),
    .Q_N(_07497_),
    .Q(\clock_inst.sec_tile.e0[21] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[22]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1114),
    .D(_00526_),
    .Q_N(_07496_),
    .Q(\clock_inst.sec_tile.e0[22] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1115),
    .D(_00527_),
    .Q_N(_07495_),
    .Q(\clock_inst.sec_tile.e0[23] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[24]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1116),
    .D(_00528_),
    .Q_N(_07494_),
    .Q(\clock_inst.sec_tile.e0[24] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[25]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1117),
    .D(_00529_),
    .Q_N(_07493_),
    .Q(\clock_inst.sec_tile.e0[25] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[26]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1118),
    .D(_00530_),
    .Q_N(_07492_),
    .Q(\clock_inst.sec_tile.e0[26] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1119),
    .D(_00531_),
    .Q_N(_07491_),
    .Q(\clock_inst.sec_tile.e0[27] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[28]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1120),
    .D(_00532_),
    .Q_N(_07490_),
    .Q(\clock_inst.sec_tile.e0[28] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[29]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1121),
    .D(_00533_),
    .Q_N(_07489_),
    .Q(\clock_inst.sec_tile.e0[29] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[2]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1122),
    .D(_00534_),
    .Q_N(_07488_),
    .Q(\clock_inst.sec_tile.e0[2] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[30]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1123),
    .D(_00535_),
    .Q_N(_07487_),
    .Q(\clock_inst.sec_tile.e0[30] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[31]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1124),
    .D(_00536_),
    .Q_N(_07486_),
    .Q(\clock_inst.sec_tile.e0[31] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[32]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1125),
    .D(_00537_),
    .Q_N(_07485_),
    .Q(\clock_inst.sec_tile.e0[32] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[33]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1126),
    .D(_00538_),
    .Q_N(_07484_),
    .Q(\clock_inst.sec_tile.e0[33] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[34]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1127),
    .D(_00539_),
    .Q_N(_07483_),
    .Q(\clock_inst.sec_tile.e0[34] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[35]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1128),
    .D(_00540_),
    .Q_N(_07482_),
    .Q(\clock_inst.sec_tile.e0[35] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[36]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1129),
    .D(_00541_),
    .Q_N(_07481_),
    .Q(\clock_inst.sec_tile.e0[36] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[37]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1130),
    .D(_00542_),
    .Q_N(_07480_),
    .Q(\clock_inst.sec_tile.e0[37] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[38]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1131),
    .D(_00543_),
    .Q_N(_07479_),
    .Q(\clock_inst.sec_tile.e0[38] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[39]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1132),
    .D(_00544_),
    .Q_N(_07478_),
    .Q(\clock_inst.sec_tile.e0[39] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1133),
    .D(_00545_),
    .Q_N(_07477_),
    .Q(\clock_inst.sec_tile.e0[3] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[40]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1134),
    .D(_00546_),
    .Q_N(_07476_),
    .Q(\clock_inst.sec_tile.e0[40] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[41]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1135),
    .D(_00547_),
    .Q_N(_07475_),
    .Q(\clock_inst.sec_tile.e0[41] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[42]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1136),
    .D(_00548_),
    .Q_N(_07474_),
    .Q(\clock_inst.sec_tile.e0[42] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[43]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1137),
    .D(_00549_),
    .Q_N(_07473_),
    .Q(\clock_inst.sec_tile.e0[43] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[44]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1138),
    .D(_00550_),
    .Q_N(_07472_),
    .Q(\clock_inst.sec_tile.e0[44] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[45]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1139),
    .D(_00551_),
    .Q_N(_07471_),
    .Q(\clock_inst.sec_tile.e0[45] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[46]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1140),
    .D(_00552_),
    .Q_N(_07470_),
    .Q(\clock_inst.sec_tile.e0[46] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[47]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1141),
    .D(_00553_),
    .Q_N(_07469_),
    .Q(\clock_inst.sec_tile.e0[47] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[48]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1142),
    .D(_00554_),
    .Q_N(_07468_),
    .Q(\clock_inst.sec_tile.e0[48] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[49]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1143),
    .D(_00555_),
    .Q_N(_07467_),
    .Q(\clock_inst.sec_tile.e0[49] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[4]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1144),
    .D(_00556_),
    .Q_N(_07466_),
    .Q(\clock_inst.sec_tile.e0[4] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[50]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1145),
    .D(_00557_),
    .Q_N(_07465_),
    .Q(\clock_inst.sec_tile.e0[50] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[51]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1146),
    .D(_00558_),
    .Q_N(_07464_),
    .Q(\clock_inst.sec_tile.e0[51] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[52]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1147),
    .D(_00559_),
    .Q_N(_07463_),
    .Q(\clock_inst.sec_tile.e0[52] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[53]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1148),
    .D(_00560_),
    .Q_N(_07462_),
    .Q(\clock_inst.sec_tile.e0[53] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1149),
    .D(_00561_),
    .Q_N(_07461_),
    .Q(\clock_inst.sec_tile.e0[5] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[6]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1150),
    .D(_00562_),
    .Q_N(_07460_),
    .Q(\clock_inst.sec_tile.e0[6] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1151),
    .D(_00563_),
    .Q_N(_07459_),
    .Q(\clock_inst.sec_tile.e0[7] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[8]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1152),
    .D(_00564_),
    .Q_N(_07458_),
    .Q(\clock_inst.sec_tile.e0[8] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e0[9]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1153),
    .D(_00565_),
    .Q_N(_07457_),
    .Q(\clock_inst.sec_tile.e0[9] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1154),
    .D(_00566_),
    .Q_N(_07456_),
    .Q(\clock_inst.sec_tile.e[0] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[10]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1155),
    .D(_00567_),
    .Q_N(_07455_),
    .Q(\clock_inst.sec_tile.e[10] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[11]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1156),
    .D(_00568_),
    .Q_N(_07454_),
    .Q(\clock_inst.sec_tile.e[11] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[12]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1157),
    .D(_00569_),
    .Q_N(_07453_),
    .Q(\clock_inst.sec_tile.e[12] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[13]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1158),
    .D(_00570_),
    .Q_N(_07452_),
    .Q(\clock_inst.sec_tile.e[13] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[14]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1159),
    .D(_00571_),
    .Q_N(_07451_),
    .Q(\clock_inst.sec_tile.e[14] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[15]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1160),
    .D(_00572_),
    .Q_N(_07450_),
    .Q(\clock_inst.sec_tile.e[15] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[16]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1161),
    .D(_00573_),
    .Q_N(_07449_),
    .Q(\clock_inst.sec_tile.e[16] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[17]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1162),
    .D(_00574_),
    .Q_N(_07448_),
    .Q(\clock_inst.sec_tile.e[17] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[18]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1163),
    .D(_00575_),
    .Q_N(_07447_),
    .Q(\clock_inst.sec_tile.e[18] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[19]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1164),
    .D(_00576_),
    .Q_N(_07446_),
    .Q(\clock_inst.sec_tile.e[19] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1165),
    .D(_00577_),
    .Q_N(_07445_),
    .Q(\clock_inst.sec_tile.e[1] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[20]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1166),
    .D(_00578_),
    .Q_N(_07444_),
    .Q(\clock_inst.sec_tile.e[20] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[21]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1167),
    .D(_00579_),
    .Q_N(_07443_),
    .Q(\clock_inst.sec_tile.e[21] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[22]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1168),
    .D(_00580_),
    .Q_N(_07442_),
    .Q(\clock_inst.sec_tile.e[22] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[23]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1169),
    .D(_00581_),
    .Q_N(_07441_),
    .Q(\clock_inst.sec_tile.e[23] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[24]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1170),
    .D(_00582_),
    .Q_N(_07440_),
    .Q(\clock_inst.sec_tile.e[24] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[25]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1171),
    .D(_00583_),
    .Q_N(_07439_),
    .Q(\clock_inst.sec_tile.e[25] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[26]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1172),
    .D(_00584_),
    .Q_N(_07438_),
    .Q(\clock_inst.sec_tile.e[26] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[27]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1173),
    .D(_00585_),
    .Q_N(_07437_),
    .Q(\clock_inst.sec_tile.e[27] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[28]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1174),
    .D(_00586_),
    .Q_N(_07436_),
    .Q(\clock_inst.sec_tile.e[28] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[29]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1175),
    .D(_00587_),
    .Q_N(_07435_),
    .Q(\clock_inst.sec_tile.e[29] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[2]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1176),
    .D(_00588_),
    .Q_N(_07434_),
    .Q(\clock_inst.sec_tile.e[2] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[30]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1177),
    .D(_00589_),
    .Q_N(_07433_),
    .Q(\clock_inst.sec_tile.e[30] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[31]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1178),
    .D(_00590_),
    .Q_N(_07432_),
    .Q(\clock_inst.sec_tile.e[31] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[32]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1179),
    .D(_00591_),
    .Q_N(_07431_),
    .Q(\clock_inst.sec_tile.e[32] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[33]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1180),
    .D(_00592_),
    .Q_N(_07430_),
    .Q(\clock_inst.sec_tile.e[33] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[34]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1181),
    .D(_00593_),
    .Q_N(_07429_),
    .Q(\clock_inst.sec_tile.e[34] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[35]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1182),
    .D(_00594_),
    .Q_N(_07428_),
    .Q(\clock_inst.sec_tile.e[35] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[36]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1183),
    .D(_00595_),
    .Q_N(_07427_),
    .Q(\clock_inst.sec_tile.e[36] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[37]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1184),
    .D(_00596_),
    .Q_N(_07426_),
    .Q(\clock_inst.sec_tile.e[37] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[38]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1185),
    .D(_00597_),
    .Q_N(_07425_),
    .Q(\clock_inst.sec_tile.e[38] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[39]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1186),
    .D(_00598_),
    .Q_N(_07424_),
    .Q(\clock_inst.sec_tile.e[39] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1187),
    .D(_00599_),
    .Q_N(_07423_),
    .Q(\clock_inst.sec_tile.e[3] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[40]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1188),
    .D(_00600_),
    .Q_N(_07422_),
    .Q(\clock_inst.sec_tile.e[40] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[41]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1189),
    .D(_00601_),
    .Q_N(_07421_),
    .Q(\clock_inst.sec_tile.e[41] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[42]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1190),
    .D(_00602_),
    .Q_N(_07420_),
    .Q(\clock_inst.sec_tile.e[42] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[43]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1191),
    .D(_00603_),
    .Q_N(_07419_),
    .Q(\clock_inst.sec_tile.e[43] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[44]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1192),
    .D(_00604_),
    .Q_N(_07418_),
    .Q(\clock_inst.sec_tile.e[44] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[45]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1193),
    .D(_00605_),
    .Q_N(_07417_),
    .Q(\clock_inst.sec_tile.e[45] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[46]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1194),
    .D(_00606_),
    .Q_N(_07416_),
    .Q(\clock_inst.sec_tile.e[46] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[47]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1195),
    .D(_00607_),
    .Q_N(_07415_),
    .Q(\clock_inst.sec_tile.e[47] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[48]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1196),
    .D(_00608_),
    .Q_N(_07414_),
    .Q(\clock_inst.sec_tile.e[48] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[49]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1197),
    .D(_00609_),
    .Q_N(_07413_),
    .Q(\clock_inst.sec_tile.e[49] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[4]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1198),
    .D(_00610_),
    .Q_N(_07412_),
    .Q(\clock_inst.sec_tile.e[4] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[50]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1199),
    .D(_00611_),
    .Q_N(_07411_),
    .Q(\clock_inst.sec_tile.e[50] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[51]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1200),
    .D(_00612_),
    .Q_N(_07410_),
    .Q(\clock_inst.sec_tile.e[51] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[52]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1201),
    .D(_00613_),
    .Q_N(_07409_),
    .Q(\clock_inst.sec_tile.e[52] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[53]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1202),
    .D(_00614_),
    .Q_N(_07408_),
    .Q(\clock_inst.sec_tile.e[53] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[5]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1203),
    .D(_00615_),
    .Q_N(_07407_),
    .Q(\clock_inst.sec_tile.e[5] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[6]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1204),
    .D(_00616_),
    .Q_N(_07406_),
    .Q(\clock_inst.sec_tile.e[6] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[7]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1205),
    .D(_00617_),
    .Q_N(_07405_),
    .Q(\clock_inst.sec_tile.e[7] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[8]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1206),
    .D(_00618_),
    .Q_N(_07404_),
    .Q(\clock_inst.sec_tile.e[8] ));
 sg13g2_dfrbp_1 \clock_inst.sec_tile.e[9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1207),
    .D(_00619_),
    .Q_N(_07403_),
    .Q(\clock_inst.sec_tile.e[9] ));
 sg13g2_dfrbp_1 \clock_inst.second[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1208),
    .D(_00620_),
    .Q_N(_00001_),
    .Q(\clock_inst.second[0] ));
 sg13g2_dfrbp_1 \clock_inst.second[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1209),
    .D(_00621_),
    .Q_N(_07402_),
    .Q(\clock_inst.second[1] ));
 sg13g2_dfrbp_1 \clock_inst.second[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1210),
    .D(_00622_),
    .Q_N(_07401_),
    .Q(\clock_inst.second[2] ));
 sg13g2_dfrbp_1 \clock_inst.second[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1211),
    .D(_00623_),
    .Q_N(_07400_),
    .Q(\clock_inst.second[3] ));
 sg13g2_dfrbp_1 \clock_inst.second[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1212),
    .D(_00624_),
    .Q_N(_07399_),
    .Q(\clock_inst.second[4] ));
 sg13g2_dfrbp_1 \clock_inst.second[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1213),
    .D(_00625_),
    .Q_N(_07398_),
    .Q(\clock_inst.second[5] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_horizontal_blank_strobe$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1214),
    .D(_00626_),
    .Q_N(_07397_),
    .Q(\clock_inst.vga_horizontal_blank_strobe ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_horizontal_visible$_SDFFE_PP1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1215),
    .D(_00627_),
    .Q_N(_07396_),
    .Q(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_hs$_SDFFE_PP1N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1216),
    .D(_00628_),
    .Q_N(_07395_),
    .Q(\clock_inst.vga_hs ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_vertical_blank_strobe$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1217),
    .D(_00629_),
    .Q_N(_07394_),
    .Q(\clock_inst.vga_inst.vga_vertical_blank_strobe ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_vertical_visible$_SDFFE_PN1P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1218),
    .D(_00630_),
    .Q_N(_07393_),
    .Q(\clock_inst.vga_inst.vga_vertical_visible ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_vs$_SDFFE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1219),
    .D(_00631_),
    .Q_N(_07392_),
    .Q(\clock_inst.vga_inst.vga_vs ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[0]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1220),
    .D(_00632_),
    .Q_N(_00003_),
    .Q(\clock_inst.vga_inst.vga_x[0] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[1]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1221),
    .D(_00633_),
    .Q_N(_07391_),
    .Q(\clock_inst.vga_inst.vga_x[1] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[2]$_SDFF_PP0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1222),
    .D(_00634_),
    .Q_N(_07390_),
    .Q(\clock_inst.vga_inst.vga_x[2] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[3]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1223),
    .D(_00635_),
    .Q_N(_07389_),
    .Q(\clock_inst.vga_inst.vga_x[3] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[4]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1224),
    .D(_00636_),
    .Q_N(_07388_),
    .Q(\clock_inst.vga_inst.vga_x[4] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[5]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1225),
    .D(_00637_),
    .Q_N(_07387_),
    .Q(\clock_inst.vga_inst.vga_x[5] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[6]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1226),
    .D(_00638_),
    .Q_N(_07386_),
    .Q(\clock_inst.vga_inst.vga_x[6] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[7]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1227),
    .D(_00639_),
    .Q_N(_07385_),
    .Q(\clock_inst.vga_inst.vga_x[7] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[8]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1228),
    .D(_00640_),
    .Q_N(_07384_),
    .Q(\clock_inst.vga_inst.vga_x[8] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_x[9]$_SDFF_PP0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1229),
    .D(_00641_),
    .Q_N(_07383_),
    .Q(\clock_inst.vga_inst.vga_x[9] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1230),
    .D(_00642_),
    .Q_N(_07382_),
    .Q(\clock_inst.vga_inst.vga_y[0] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1231),
    .D(_00643_),
    .Q_N(_07381_),
    .Q(\clock_inst.vga_inst.vga_y[1] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1232),
    .D(_00644_),
    .Q_N(_07380_),
    .Q(\clock_inst.vga_inst.vga_y[2] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1233),
    .D(_00645_),
    .Q_N(_07379_),
    .Q(\clock_inst.vga_inst.vga_y[3] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1234),
    .D(_00646_),
    .Q_N(_07378_),
    .Q(\clock_inst.vga_inst.vga_y[4] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1235),
    .D(_00647_),
    .Q_N(_07377_),
    .Q(\clock_inst.vga_inst.vga_y[5] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1236),
    .D(_00648_),
    .Q_N(_07376_),
    .Q(\clock_inst.vga_inst.vga_y[6] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1237),
    .D(_00649_),
    .Q_N(_07375_),
    .Q(\clock_inst.vga_inst.vga_y[7] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1238),
    .D(_00650_),
    .Q_N(_07374_),
    .Q(\clock_inst.vga_inst.vga_y[8] ));
 sg13g2_dfrbp_1 \clock_inst.vga_inst.vga_y[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1239),
    .D(_00651_),
    .Q_N(_07373_),
    .Q(\clock_inst.vga_inst.vga_y[9] ));
 sg13g2_dfrbp_1 \clock_inst.vga_rgb[1]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1240),
    .D(_00652_),
    .Q_N(_07372_),
    .Q(net19));
 sg13g2_dfrbp_1 \clock_inst.vga_rgb[3]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1241),
    .D(_00653_),
    .Q_N(_07371_),
    .Q(net18));
 sg13g2_dfrbp_1 \clock_inst.vga_rgb[4]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1242),
    .D(_00654_),
    .Q_N(_07370_),
    .Q(net17));
 sg13g2_buf_1 input1 (.A(ui_in[2]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[7]),
    .X(net4));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[0]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[1]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[2]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[3]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[4]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[5]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[6]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[7]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[0]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[1]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[2]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[3]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[4]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[5]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[6]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout21 (.A(_07022_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_05006_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_01241_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_07274_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_06729_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_06184_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_05092_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_03225_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_03163_),
    .X(net29));
 sg13g2_buf_4 fanout30 (.X(net30),
    .A(_03023_));
 sg13g2_buf_2 fanout31 (.A(_02971_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_02871_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_02783_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_02736_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_02538_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_02520_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02429_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02351_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02251_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_02247_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_02172_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_02042_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_01925_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_01583_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_01573_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_01545_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_01471_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_01393_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_01240_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_01213_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_01203_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_01186_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_06857_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_06304_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_06272_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_05768_),
    .X(net56));
 sg13g2_buf_4 fanout57 (.X(net57),
    .A(_05360_));
 sg13g2_buf_2 fanout58 (.A(_05327_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_05319_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_05049_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_04933_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_04825_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_04792_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_04602_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_04420_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_04146_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_04134_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_03953_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_03671_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_02535_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_02350_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_02246_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_02171_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_01990_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_01914_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_01913_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_01844_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_01787_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_01687_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_01679_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_01654_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_01611_),
    .X(net82));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_01590_));
 sg13g2_buf_2 fanout84 (.A(_01519_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_01504_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_01492_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_01460_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_01458_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_01443_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_01377_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_01360_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_01356_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_01350_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_01279_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_01275_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_01263_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_01252_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_01247_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_01239_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_01230_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_01222_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_01216_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_01212_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_01202_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_01177_),
    .X(net105));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_01166_));
 sg13g2_buf_2 fanout107 (.A(_01162_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_01137_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_01120_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_01072_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_01062_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_01034_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_06260_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_05559_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_05321_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_05250_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_05231_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_05134_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_05091_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_05002_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_04950_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_04938_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_04937_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_04066_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_03918_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_03894_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_03845_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_02816_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_02747_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_02586_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_02550_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_02548_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_02430_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_02272_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_02131_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_02101_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_02073_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_01926_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_01746_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_01686_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_01655_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_01641_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_01559_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_01472_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_01409_),
    .X(net145));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(_01381_));
 sg13g2_buf_2 fanout147 (.A(_01347_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_01310_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_01293_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_01215_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_01201_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_01179_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_01176_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_01152_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_01138_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_01136_),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(_01130_));
 sg13g2_buf_2 fanout158 (.A(_01119_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_01071_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_01064_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_01061_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_01033_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_05616_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_05475_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_05393_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_05346_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_05330_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_05320_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_05303_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_05301_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_05256_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_05253_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_05245_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_05236_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_05225_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_05203_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_05173_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_05146_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_05136_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_05118_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_05093_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_05087_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_05080_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_05043_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_05021_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_05011_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_04970_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_04967_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_04953_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_04943_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_04936_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_04831_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_03090_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_02896_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_02874_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_02773_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_02767_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_02746_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_02711_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_02664_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_02649_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_02589_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_02585_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_02557_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_02544_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_02539_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_02527_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_02517_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_02509_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_02503_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_02483_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_02478_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_02475_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_02463_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_02442_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_02434_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_02407_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_02403_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_02382_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_02379_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_02376_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_02374_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_02373_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_02371_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_02365_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_02340_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_02295_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_02278_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_02270_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_02268_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_02236_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_01527_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_01380_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_01297_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_01284_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_01248_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_01210_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_01178_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_01151_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_01135_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_01070_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_01063_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_01055_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_01032_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_00663_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_06276_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_05704_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_05323_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_05298_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_05269_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_05262_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_05247_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_05241_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_05234_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_05202_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_05199_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_05169_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_05165_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_05154_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_05145_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_05131_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_05123_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_05102_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_05094_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_05067_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_05062_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_05057_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_05042_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_05032_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_05030_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_05022_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_05020_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_05016_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_05014_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_04987_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_04982_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_04979_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_04974_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_04966_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_04961_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_04957_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_04955_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_04952_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_04947_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_04945_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_04942_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_04941_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_04915_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_04904_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_04888_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_04866_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_04849_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_04844_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_04830_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_03033_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_02833_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_02772_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_02751_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_02716_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_02677_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_02639_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_02610_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_02608_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_02601_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_02584_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_02570_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_02561_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_02558_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_02545_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_02516_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_02501_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_02492_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_02488_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_02486_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_02473_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_02469_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_02465_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_02462_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_02456_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_02452_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_02448_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_02437_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_02432_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_02418_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_02416_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_02415_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_02410_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_02406_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_02402_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_02398_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_02391_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_02375_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_02364_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_02359_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_02339_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_02322_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_02315_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_02304_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_02281_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_02277_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_02274_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_02269_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_02267_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_02266_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_02264_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_02242_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_02239_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_02235_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_02234_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_02232_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_02225_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_02191_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_02188_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_02185_),
    .X(net354));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(_02061_));
 sg13g2_buf_2 fanout356 (.A(_01965_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_01797_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_00943_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_00837_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_00825_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_00763_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_00691_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_00687_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_00674_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_00662_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_06875_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_05251_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_05205_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_05186_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_05156_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_05144_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_05142_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_05127_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_05098_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_05073_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_05068_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_05036_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_05029_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_05019_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_05008_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_04996_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_04973_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_04960_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_04956_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_04954_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_04951_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_04944_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_04940_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_04914_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_04909_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_04906_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_04898_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_04894_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_04887_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_04878_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_04873_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_04871_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_04868_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_04862_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_04858_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_04857_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_04848_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_04839_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_04829_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_04793_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_04445_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_02606_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_02580_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_02576_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_02523_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_02491_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_02481_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_02454_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_02436_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_02431_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_02411_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_02409_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_02405_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_02401_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_02384_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_02356_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_02334_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_02323_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_02321_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_02303_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_02273_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_02265_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_02241_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_02238_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_02224_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_02223_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_02219_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_02211_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_02209_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_02206_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_02201_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_02198_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_02195_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_02187_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_02184_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_02003_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_01964_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_01816_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_01811_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_01796_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_01778_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_01743_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_01682_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_00845_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_00748_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_00703_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_00685_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_00680_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_00675_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_06545_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_05214_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_05141_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_04972_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_04929_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_04921_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_04919_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_04913_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_04907_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_04886_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_04875_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_04874_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_04872_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_04867_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_04861_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_04853_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_04847_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_04842_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_04841_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_04834_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_04828_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_04818_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_03892_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_02740_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_02569_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_02355_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_02329_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_02320_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_02302_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_02292_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_02286_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_02240_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_02226_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_02222_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_02218_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_02215_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_02203_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_02197_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_02194_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_02192_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_02189_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_02186_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_02183_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_02177_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_01815_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_01728_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_01681_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_01677_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_00881_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_00790_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_00777_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_00767_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_00746_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_00742_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_00737_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_00718_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_00709_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_00695_),
    .X(net512));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(_00689_));
 sg13g2_buf_2 fanout514 (.A(_00684_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_00672_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_00668_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_00666_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_07184_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_07017_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_06277_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_06270_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_05487_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_05140_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_04912_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_04855_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_04854_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_04850_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_04846_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_04833_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_04827_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_04165_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_02866_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_02782_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_02282_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_02250_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_02217_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_02214_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_02212_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_02182_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_02176_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_02173_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_01676_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_01038_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_00858_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_00735_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_00732_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_00698_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_00694_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_00683_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_00677_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_07346_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_07169_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_07005_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_06831_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_06794_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_06387_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_05486_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_05355_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_05001_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_04816_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_04810_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_04475_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_04464_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_04444_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_04266_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_02958_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_02853_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_02567_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_02249_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_02161_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_02153_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_01725_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_01036_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_01027_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_00925_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_00857_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_00827_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_00800_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_00752_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_00670_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_00664_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_00657_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_00656_),
    .X(net583));
 sg13g2_tiehi _15393__584 (.L_HI(net584));
 sg13g2_tiehi _15394__585 (.L_HI(net585));
 sg13g2_tiehi _15395__586 (.L_HI(net586));
 sg13g2_tiehi _15396__587 (.L_HI(net587));
 sg13g2_tiehi _15397__588 (.L_HI(net588));
 sg13g2_tiehi _15398__589 (.L_HI(net589));
 sg13g2_tiehi _15399__590 (.L_HI(net590));
 sg13g2_tiehi _15400__591 (.L_HI(net591));
 sg13g2_tiehi \clock_inst.frameno[0]$_SDFFE_PP0P__592  (.L_HI(net592));
 sg13g2_tiehi \clock_inst.frameno[1]$_SDFFE_PP0P__593  (.L_HI(net593));
 sg13g2_tiehi \clock_inst.frameno[2]$_SDFFE_PP0P__594  (.L_HI(net594));
 sg13g2_tiehi \clock_inst.frameno[3]$_SDFFE_PP0P__595  (.L_HI(net595));
 sg13g2_tiehi \clock_inst.frameno[4]$_SDFFE_PP0P__596  (.L_HI(net596));
 sg13g2_tiehi \clock_inst.frameno[5]$_SDFFE_PP0P__597  (.L_HI(net597));
 sg13g2_tiehi \clock_inst.frameno[6]$_SDFFE_PP0P__598  (.L_HI(net598));
 sg13g2_tiehi \clock_inst.hour[0]$_SDFFE_PN1P__599  (.L_HI(net599));
 sg13g2_tiehi \clock_inst.hour[1]$_SDFFE_PP0N__600  (.L_HI(net600));
 sg13g2_tiehi \clock_inst.hour[2]$_SDFFE_PP0N__601  (.L_HI(net601));
 sg13g2_tiehi \clock_inst.hour[3]$_SDFFE_PN1P__602  (.L_HI(net602));
 sg13g2_tiehi \clock_inst.hour_a[0]$_DFFE_PP__603  (.L_HI(net603));
 sg13g2_tiehi \clock_inst.hour_a[17]$_DFFE_PP__604  (.L_HI(net604));
 sg13g2_tiehi \clock_inst.hour_a[19]$_DFFE_PP__605  (.L_HI(net605));
 sg13g2_tiehi \clock_inst.hour_a[1]$_DFFE_PP__606  (.L_HI(net606));
 sg13g2_tiehi \clock_inst.hour_a[20]$_DFFE_PP__607  (.L_HI(net607));
 sg13g2_tiehi \clock_inst.hour_a[21]$_DFFE_PP__608  (.L_HI(net608));
 sg13g2_tiehi \clock_inst.hour_a[22]$_DFFE_PP__609  (.L_HI(net609));
 sg13g2_tiehi \clock_inst.hour_a[23]$_DFFE_PP__610  (.L_HI(net610));
 sg13g2_tiehi \clock_inst.hour_a[2]$_DFFE_PP__611  (.L_HI(net611));
 sg13g2_tiehi \clock_inst.hour_a[35]$_DFFE_PP__612  (.L_HI(net612));
 sg13g2_tiehi \clock_inst.hour_a[36]$_DFFE_PP__613  (.L_HI(net613));
 sg13g2_tiehi \clock_inst.hour_a[37]$_DFFE_PP__614  (.L_HI(net614));
 sg13g2_tiehi \clock_inst.hour_a[38]$_DFFE_PP__615  (.L_HI(net615));
 sg13g2_tiehi \clock_inst.hour_a[39]$_DFFE_PP__616  (.L_HI(net616));
 sg13g2_tiehi \clock_inst.hour_a[3]$_DFFE_PP__617  (.L_HI(net617));
 sg13g2_tiehi \clock_inst.hour_a[40]$_DFFE_PP__618  (.L_HI(net618));
 sg13g2_tiehi \clock_inst.hour_a[41]$_DFFE_PP__619  (.L_HI(net619));
 sg13g2_tiehi \clock_inst.hour_a[42]$_DFFE_PP__620  (.L_HI(net620));
 sg13g2_tiehi \clock_inst.hour_a[43]$_DFFE_PP__621  (.L_HI(net621));
 sg13g2_tiehi \clock_inst.hour_a[52]$_DFFE_PP__622  (.L_HI(net622));
 sg13g2_tiehi \clock_inst.hour_a[5]$_DFFE_PP__623  (.L_HI(net623));
 sg13g2_tiehi \clock_inst.hour_a[6]$_DFFE_PP__624  (.L_HI(net624));
 sg13g2_tiehi \clock_inst.hour_a[7]$_DFFE_PP__625  (.L_HI(net625));
 sg13g2_tiehi \clock_inst.hour_b[0]$_DFFE_PP__626  (.L_HI(net626));
 sg13g2_tiehi \clock_inst.hour_b[17]$_DFFE_PP__627  (.L_HI(net627));
 sg13g2_tiehi \clock_inst.hour_b[19]$_DFFE_PP__628  (.L_HI(net628));
 sg13g2_tiehi \clock_inst.hour_b[1]$_DFFE_PP__629  (.L_HI(net629));
 sg13g2_tiehi \clock_inst.hour_b[20]$_DFFE_PP__630  (.L_HI(net630));
 sg13g2_tiehi \clock_inst.hour_b[22]$_DFFE_PP__631  (.L_HI(net631));
 sg13g2_tiehi \clock_inst.hour_b[23]$_DFFE_PP__632  (.L_HI(net632));
 sg13g2_tiehi \clock_inst.hour_b[2]$_DFFE_PP__633  (.L_HI(net633));
 sg13g2_tiehi \clock_inst.hour_b[35]$_DFFE_PP__634  (.L_HI(net634));
 sg13g2_tiehi \clock_inst.hour_b[36]$_DFFE_PP__635  (.L_HI(net635));
 sg13g2_tiehi \clock_inst.hour_b[37]$_DFFE_PP__636  (.L_HI(net636));
 sg13g2_tiehi \clock_inst.hour_b[38]$_DFFE_PP__637  (.L_HI(net637));
 sg13g2_tiehi \clock_inst.hour_b[39]$_DFFE_PP__638  (.L_HI(net638));
 sg13g2_tiehi \clock_inst.hour_b[40]$_DFFE_PP__639  (.L_HI(net639));
 sg13g2_tiehi \clock_inst.hour_b[41]$_DFFE_PP__640  (.L_HI(net640));
 sg13g2_tiehi \clock_inst.hour_b[42]$_DFFE_PP__641  (.L_HI(net641));
 sg13g2_tiehi \clock_inst.hour_b[4]$_DFFE_PP__642  (.L_HI(net642));
 sg13g2_tiehi \clock_inst.hour_b[5]$_DFFE_PP__643  (.L_HI(net643));
 sg13g2_tiehi \clock_inst.hour_c[10]$_DFFE_PP__644  (.L_HI(net644));
 sg13g2_tiehi \clock_inst.hour_c[11]$_DFFE_PP__645  (.L_HI(net645));
 sg13g2_tiehi \clock_inst.hour_c[12]$_DFFE_PP__646  (.L_HI(net646));
 sg13g2_tiehi \clock_inst.hour_c[13]$_DFFE_PP__647  (.L_HI(net647));
 sg13g2_tiehi \clock_inst.hour_c[14]$_DFFE_PP__648  (.L_HI(net648));
 sg13g2_tiehi \clock_inst.hour_c[15]$_DFFE_PP__649  (.L_HI(net649));
 sg13g2_tiehi \clock_inst.hour_c[16]$_DFFE_PP__650  (.L_HI(net650));
 sg13g2_tiehi \clock_inst.hour_c[17]$_DFFE_PP__651  (.L_HI(net651));
 sg13g2_tiehi \clock_inst.hour_c[18]$_DFFE_PP__652  (.L_HI(net652));
 sg13g2_tiehi \clock_inst.hour_c[19]$_DFFE_PP__653  (.L_HI(net653));
 sg13g2_tiehi \clock_inst.hour_c[1]$_DFFE_PP__654  (.L_HI(net654));
 sg13g2_tiehi \clock_inst.hour_c[21]$_DFFE_PP__655  (.L_HI(net655));
 sg13g2_tiehi \clock_inst.hour_c[23]$_DFFE_PP__656  (.L_HI(net656));
 sg13g2_tiehi \clock_inst.hour_c[24]$_DFFE_PP__657  (.L_HI(net657));
 sg13g2_tiehi \clock_inst.hour_c[25]$_DFFE_PP__658  (.L_HI(net658));
 sg13g2_tiehi \clock_inst.hour_c[26]$_DFFE_PP__659  (.L_HI(net659));
 sg13g2_tiehi \clock_inst.hour_c[27]$_DFFE_PP__660  (.L_HI(net660));
 sg13g2_tiehi \clock_inst.hour_c[28]$_DFFE_PP__661  (.L_HI(net661));
 sg13g2_tiehi \clock_inst.hour_c[29]$_DFFE_PP__662  (.L_HI(net662));
 sg13g2_tiehi \clock_inst.hour_c[30]$_DFFE_PP__663  (.L_HI(net663));
 sg13g2_tiehi \clock_inst.hour_c[31]$_DFFE_PP__664  (.L_HI(net664));
 sg13g2_tiehi \clock_inst.hour_c[32]$_DFFE_PP__665  (.L_HI(net665));
 sg13g2_tiehi \clock_inst.hour_c[35]$_DFFE_PP__666  (.L_HI(net666));
 sg13g2_tiehi \clock_inst.hour_c[36]$_DFFE_PP__667  (.L_HI(net667));
 sg13g2_tiehi \clock_inst.hour_c[37]$_DFFE_PP__668  (.L_HI(net668));
 sg13g2_tiehi \clock_inst.hour_c[39]$_DFFE_PP__669  (.L_HI(net669));
 sg13g2_tiehi \clock_inst.hour_c[40]$_DFFE_PP__670  (.L_HI(net670));
 sg13g2_tiehi \clock_inst.hour_c[41]$_DFFE_PP__671  (.L_HI(net671));
 sg13g2_tiehi \clock_inst.hour_c[42]$_DFFE_PP__672  (.L_HI(net672));
 sg13g2_tiehi \clock_inst.hour_c[43]$_DFFE_PP__673  (.L_HI(net673));
 sg13g2_tiehi \clock_inst.hour_c[44]$_DFFE_PP__674  (.L_HI(net674));
 sg13g2_tiehi \clock_inst.hour_c[45]$_DFFE_PP__675  (.L_HI(net675));
 sg13g2_tiehi \clock_inst.hour_c[46]$_DFFE_PP__676  (.L_HI(net676));
 sg13g2_tiehi \clock_inst.hour_c[49]$_DFFE_PP__677  (.L_HI(net677));
 sg13g2_tiehi \clock_inst.hour_c[50]$_DFFE_PP__678  (.L_HI(net678));
 sg13g2_tiehi \clock_inst.hour_c[51]$_DFFE_PP__679  (.L_HI(net679));
 sg13g2_tiehi \clock_inst.hour_c[52]$_DFFE_PP__680  (.L_HI(net680));
 sg13g2_tiehi \clock_inst.hour_c[5]$_DFFE_PP__681  (.L_HI(net681));
 sg13g2_tiehi \clock_inst.hour_c[6]$_DFFE_PP__682  (.L_HI(net682));
 sg13g2_tiehi \clock_inst.hour_c[7]$_DFFE_PP__683  (.L_HI(net683));
 sg13g2_tiehi \clock_inst.hour_c[8]$_DFFE_PP__684  (.L_HI(net684));
 sg13g2_tiehi \clock_inst.hour_c[9]$_DFFE_PP__685  (.L_HI(net685));
 sg13g2_tiehi \clock_inst.hour_tile.e0[0]$_DFFE_PP__686  (.L_HI(net686));
 sg13g2_tiehi \clock_inst.hour_tile.e0[10]$_DFFE_PP__687  (.L_HI(net687));
 sg13g2_tiehi \clock_inst.hour_tile.e0[11]$_DFFE_PP__688  (.L_HI(net688));
 sg13g2_tiehi \clock_inst.hour_tile.e0[12]$_DFFE_PP__689  (.L_HI(net689));
 sg13g2_tiehi \clock_inst.hour_tile.e0[13]$_DFFE_PP__690  (.L_HI(net690));
 sg13g2_tiehi \clock_inst.hour_tile.e0[14]$_DFFE_PP__691  (.L_HI(net691));
 sg13g2_tiehi \clock_inst.hour_tile.e0[15]$_DFFE_PP__692  (.L_HI(net692));
 sg13g2_tiehi \clock_inst.hour_tile.e0[16]$_DFFE_PP__693  (.L_HI(net693));
 sg13g2_tiehi \clock_inst.hour_tile.e0[17]$_DFFE_PP__694  (.L_HI(net694));
 sg13g2_tiehi \clock_inst.hour_tile.e0[18]$_DFFE_PP__695  (.L_HI(net695));
 sg13g2_tiehi \clock_inst.hour_tile.e0[19]$_DFFE_PP__696  (.L_HI(net696));
 sg13g2_tiehi \clock_inst.hour_tile.e0[1]$_DFFE_PP__697  (.L_HI(net697));
 sg13g2_tiehi \clock_inst.hour_tile.e0[20]$_SDFFCE_PP0P__698  (.L_HI(net698));
 sg13g2_tiehi \clock_inst.hour_tile.e0[21]$_DFFE_PP__699  (.L_HI(net699));
 sg13g2_tiehi \clock_inst.hour_tile.e0[22]$_SDFFCE_PP0P__700  (.L_HI(net700));
 sg13g2_tiehi \clock_inst.hour_tile.e0[23]$_DFFE_PP__701  (.L_HI(net701));
 sg13g2_tiehi \clock_inst.hour_tile.e0[24]$_DFFE_PP__702  (.L_HI(net702));
 sg13g2_tiehi \clock_inst.hour_tile.e0[25]$_DFFE_PP__703  (.L_HI(net703));
 sg13g2_tiehi \clock_inst.hour_tile.e0[26]$_DFFE_PP__704  (.L_HI(net704));
 sg13g2_tiehi \clock_inst.hour_tile.e0[27]$_DFFE_PP__705  (.L_HI(net705));
 sg13g2_tiehi \clock_inst.hour_tile.e0[28]$_DFFE_PP__706  (.L_HI(net706));
 sg13g2_tiehi \clock_inst.hour_tile.e0[29]$_DFFE_PP__707  (.L_HI(net707));
 sg13g2_tiehi \clock_inst.hour_tile.e0[2]$_DFFE_PP__708  (.L_HI(net708));
 sg13g2_tiehi \clock_inst.hour_tile.e0[30]$_DFFE_PP__709  (.L_HI(net709));
 sg13g2_tiehi \clock_inst.hour_tile.e0[31]$_DFFE_PP__710  (.L_HI(net710));
 sg13g2_tiehi \clock_inst.hour_tile.e0[32]$_DFFE_PP__711  (.L_HI(net711));
 sg13g2_tiehi \clock_inst.hour_tile.e0[33]$_DFFE_PP__712  (.L_HI(net712));
 sg13g2_tiehi \clock_inst.hour_tile.e0[34]$_DFFE_PP__713  (.L_HI(net713));
 sg13g2_tiehi \clock_inst.hour_tile.e0[35]$_DFFE_PP__714  (.L_HI(net714));
 sg13g2_tiehi \clock_inst.hour_tile.e0[36]$_DFFE_PP__715  (.L_HI(net715));
 sg13g2_tiehi \clock_inst.hour_tile.e0[37]$_DFFE_PP__716  (.L_HI(net716));
 sg13g2_tiehi \clock_inst.hour_tile.e0[38]$_DFFE_PP__717  (.L_HI(net717));
 sg13g2_tiehi \clock_inst.hour_tile.e0[39]$_DFFE_PP__718  (.L_HI(net718));
 sg13g2_tiehi \clock_inst.hour_tile.e0[3]$_DFFE_PP__719  (.L_HI(net719));
 sg13g2_tiehi \clock_inst.hour_tile.e0[40]$_DFFE_PP__720  (.L_HI(net720));
 sg13g2_tiehi \clock_inst.hour_tile.e0[41]$_DFFE_PP__721  (.L_HI(net721));
 sg13g2_tiehi \clock_inst.hour_tile.e0[42]$_DFFE_PP__722  (.L_HI(net722));
 sg13g2_tiehi \clock_inst.hour_tile.e0[43]$_DFFE_PP__723  (.L_HI(net723));
 sg13g2_tiehi \clock_inst.hour_tile.e0[44]$_DFFE_PP__724  (.L_HI(net724));
 sg13g2_tiehi \clock_inst.hour_tile.e0[45]$_DFFE_PP__725  (.L_HI(net725));
 sg13g2_tiehi \clock_inst.hour_tile.e0[46]$_DFFE_PP__726  (.L_HI(net726));
 sg13g2_tiehi \clock_inst.hour_tile.e0[47]$_SDFFCE_PP1P__727  (.L_HI(net727));
 sg13g2_tiehi \clock_inst.hour_tile.e0[48]$_SDFFCE_PP0P__728  (.L_HI(net728));
 sg13g2_tiehi \clock_inst.hour_tile.e0[49]$_DFFE_PP__729  (.L_HI(net729));
 sg13g2_tiehi \clock_inst.hour_tile.e0[4]$_DFFE_PP__730  (.L_HI(net730));
 sg13g2_tiehi \clock_inst.hour_tile.e0[50]$_DFFE_PP__731  (.L_HI(net731));
 sg13g2_tiehi \clock_inst.hour_tile.e0[51]$_DFFE_PP__732  (.L_HI(net732));
 sg13g2_tiehi \clock_inst.hour_tile.e0[52]$_DFFE_PP__733  (.L_HI(net733));
 sg13g2_tiehi \clock_inst.hour_tile.e0[53]$_DFFE_PP__734  (.L_HI(net734));
 sg13g2_tiehi \clock_inst.hour_tile.e0[5]$_DFFE_PP__735  (.L_HI(net735));
 sg13g2_tiehi \clock_inst.hour_tile.e0[6]$_DFFE_PP__736  (.L_HI(net736));
 sg13g2_tiehi \clock_inst.hour_tile.e0[7]$_DFFE_PP__737  (.L_HI(net737));
 sg13g2_tiehi \clock_inst.hour_tile.e0[8]$_DFFE_PP__738  (.L_HI(net738));
 sg13g2_tiehi \clock_inst.hour_tile.e0[9]$_DFFE_PP__739  (.L_HI(net739));
 sg13g2_tiehi \clock_inst.hour_tile.e[0]$_DFFE_PP__740  (.L_HI(net740));
 sg13g2_tiehi \clock_inst.hour_tile.e[10]$_DFFE_PP__741  (.L_HI(net741));
 sg13g2_tiehi \clock_inst.hour_tile.e[11]$_DFFE_PP__742  (.L_HI(net742));
 sg13g2_tiehi \clock_inst.hour_tile.e[12]$_DFFE_PP__743  (.L_HI(net743));
 sg13g2_tiehi \clock_inst.hour_tile.e[13]$_DFFE_PP__744  (.L_HI(net744));
 sg13g2_tiehi \clock_inst.hour_tile.e[14]$_DFFE_PP__745  (.L_HI(net745));
 sg13g2_tiehi \clock_inst.hour_tile.e[15]$_DFFE_PP__746  (.L_HI(net746));
 sg13g2_tiehi \clock_inst.hour_tile.e[16]$_DFFE_PP__747  (.L_HI(net747));
 sg13g2_tiehi \clock_inst.hour_tile.e[17]$_DFFE_PP__748  (.L_HI(net748));
 sg13g2_tiehi \clock_inst.hour_tile.e[18]$_DFFE_PP__749  (.L_HI(net749));
 sg13g2_tiehi \clock_inst.hour_tile.e[19]$_DFFE_PP__750  (.L_HI(net750));
 sg13g2_tiehi \clock_inst.hour_tile.e[1]$_DFFE_PP__751  (.L_HI(net751));
 sg13g2_tiehi \clock_inst.hour_tile.e[20]$_SDFFCE_PP0P__752  (.L_HI(net752));
 sg13g2_tiehi \clock_inst.hour_tile.e[21]$_DFFE_PP__753  (.L_HI(net753));
 sg13g2_tiehi \clock_inst.hour_tile.e[22]$_SDFFCE_PP0P__754  (.L_HI(net754));
 sg13g2_tiehi \clock_inst.hour_tile.e[23]$_DFFE_PP__755  (.L_HI(net755));
 sg13g2_tiehi \clock_inst.hour_tile.e[24]$_DFFE_PP__756  (.L_HI(net756));
 sg13g2_tiehi \clock_inst.hour_tile.e[25]$_DFFE_PP__757  (.L_HI(net757));
 sg13g2_tiehi \clock_inst.hour_tile.e[26]$_DFFE_PP__758  (.L_HI(net758));
 sg13g2_tiehi \clock_inst.hour_tile.e[27]$_DFFE_PP__759  (.L_HI(net759));
 sg13g2_tiehi \clock_inst.hour_tile.e[28]$_DFFE_PP__760  (.L_HI(net760));
 sg13g2_tiehi \clock_inst.hour_tile.e[29]$_DFFE_PP__761  (.L_HI(net761));
 sg13g2_tiehi \clock_inst.hour_tile.e[2]$_DFFE_PP__762  (.L_HI(net762));
 sg13g2_tiehi \clock_inst.hour_tile.e[30]$_DFFE_PP__763  (.L_HI(net763));
 sg13g2_tiehi \clock_inst.hour_tile.e[31]$_DFFE_PP__764  (.L_HI(net764));
 sg13g2_tiehi \clock_inst.hour_tile.e[32]$_DFFE_PP__765  (.L_HI(net765));
 sg13g2_tiehi \clock_inst.hour_tile.e[33]$_DFFE_PP__766  (.L_HI(net766));
 sg13g2_tiehi \clock_inst.hour_tile.e[34]$_DFFE_PP__767  (.L_HI(net767));
 sg13g2_tiehi \clock_inst.hour_tile.e[35]$_DFFE_PP__768  (.L_HI(net768));
 sg13g2_tiehi \clock_inst.hour_tile.e[36]$_DFFE_PP__769  (.L_HI(net769));
 sg13g2_tiehi \clock_inst.hour_tile.e[37]$_DFFE_PP__770  (.L_HI(net770));
 sg13g2_tiehi \clock_inst.hour_tile.e[38]$_DFFE_PP__771  (.L_HI(net771));
 sg13g2_tiehi \clock_inst.hour_tile.e[39]$_DFFE_PP__772  (.L_HI(net772));
 sg13g2_tiehi \clock_inst.hour_tile.e[3]$_DFFE_PP__773  (.L_HI(net773));
 sg13g2_tiehi \clock_inst.hour_tile.e[40]$_DFFE_PP__774  (.L_HI(net774));
 sg13g2_tiehi \clock_inst.hour_tile.e[41]$_DFFE_PP__775  (.L_HI(net775));
 sg13g2_tiehi \clock_inst.hour_tile.e[42]$_DFFE_PP__776  (.L_HI(net776));
 sg13g2_tiehi \clock_inst.hour_tile.e[43]$_DFFE_PP__777  (.L_HI(net777));
 sg13g2_tiehi \clock_inst.hour_tile.e[44]$_DFFE_PP__778  (.L_HI(net778));
 sg13g2_tiehi \clock_inst.hour_tile.e[45]$_DFFE_PP__779  (.L_HI(net779));
 sg13g2_tiehi \clock_inst.hour_tile.e[46]$_DFFE_PP__780  (.L_HI(net780));
 sg13g2_tiehi \clock_inst.hour_tile.e[47]$_SDFFCE_PP1P__781  (.L_HI(net781));
 sg13g2_tiehi \clock_inst.hour_tile.e[48]$_SDFFCE_PP0P__782  (.L_HI(net782));
 sg13g2_tiehi \clock_inst.hour_tile.e[49]$_DFFE_PP__783  (.L_HI(net783));
 sg13g2_tiehi \clock_inst.hour_tile.e[4]$_DFFE_PP__784  (.L_HI(net784));
 sg13g2_tiehi \clock_inst.hour_tile.e[50]$_DFFE_PP__785  (.L_HI(net785));
 sg13g2_tiehi \clock_inst.hour_tile.e[51]$_DFFE_PP__786  (.L_HI(net786));
 sg13g2_tiehi \clock_inst.hour_tile.e[52]$_DFFE_PP__787  (.L_HI(net787));
 sg13g2_tiehi \clock_inst.hour_tile.e[53]$_DFFE_PP__788  (.L_HI(net788));
 sg13g2_tiehi \clock_inst.hour_tile.e[5]$_DFFE_PP__789  (.L_HI(net789));
 sg13g2_tiehi \clock_inst.hour_tile.e[6]$_DFFE_PP__790  (.L_HI(net790));
 sg13g2_tiehi \clock_inst.hour_tile.e[7]$_DFFE_PP__791  (.L_HI(net791));
 sg13g2_tiehi \clock_inst.hour_tile.e[8]$_DFFE_PP__792  (.L_HI(net792));
 sg13g2_tiehi \clock_inst.hour_tile.e[9]$_DFFE_PP__793  (.L_HI(net793));
 sg13g2_tiehi \clock_inst.min_a[0]$_DFFE_PP__794  (.L_HI(net794));
 sg13g2_tiehi \clock_inst.min_a[17]$_DFFE_PP__795  (.L_HI(net795));
 sg13g2_tiehi \clock_inst.min_a[18]$_DFFE_PP__796  (.L_HI(net796));
 sg13g2_tiehi \clock_inst.min_a[19]$_DFFE_PP__797  (.L_HI(net797));
 sg13g2_tiehi \clock_inst.min_a[1]$_DFFE_PP__798  (.L_HI(net798));
 sg13g2_tiehi \clock_inst.min_a[20]$_DFFE_PP__799  (.L_HI(net799));
 sg13g2_tiehi \clock_inst.min_a[21]$_DFFE_PP__800  (.L_HI(net800));
 sg13g2_tiehi \clock_inst.min_a[22]$_DFFE_PP__801  (.L_HI(net801));
 sg13g2_tiehi \clock_inst.min_a[23]$_DFFE_PP__802  (.L_HI(net802));
 sg13g2_tiehi \clock_inst.min_a[2]$_DFFE_PP__803  (.L_HI(net803));
 sg13g2_tiehi \clock_inst.min_a[35]$_DFFE_PP__804  (.L_HI(net804));
 sg13g2_tiehi \clock_inst.min_a[36]$_DFFE_PP__805  (.L_HI(net805));
 sg13g2_tiehi \clock_inst.min_a[37]$_DFFE_PP__806  (.L_HI(net806));
 sg13g2_tiehi \clock_inst.min_a[38]$_DFFE_PP__807  (.L_HI(net807));
 sg13g2_tiehi \clock_inst.min_a[39]$_DFFE_PP__808  (.L_HI(net808));
 sg13g2_tiehi \clock_inst.min_a[3]$_DFFE_PP__809  (.L_HI(net809));
 sg13g2_tiehi \clock_inst.min_a[40]$_DFFE_PP__810  (.L_HI(net810));
 sg13g2_tiehi \clock_inst.min_a[41]$_DFFE_PP__811  (.L_HI(net811));
 sg13g2_tiehi \clock_inst.min_a[42]$_DFFE_PP__812  (.L_HI(net812));
 sg13g2_tiehi \clock_inst.min_a[43]$_DFFE_PP__813  (.L_HI(net813));
 sg13g2_tiehi \clock_inst.min_a[44]$_DFFE_PP__814  (.L_HI(net814));
 sg13g2_tiehi \clock_inst.min_a[4]$_DFFE_PP__815  (.L_HI(net815));
 sg13g2_tiehi \clock_inst.min_a[52]$_DFFE_PP__816  (.L_HI(net816));
 sg13g2_tiehi \clock_inst.min_a[5]$_DFFE_PP__817  (.L_HI(net817));
 sg13g2_tiehi \clock_inst.min_a[6]$_DFFE_PP__818  (.L_HI(net818));
 sg13g2_tiehi \clock_inst.min_a[7]$_DFFE_PP__819  (.L_HI(net819));
 sg13g2_tiehi \clock_inst.min_a[8]$_DFFE_PP__820  (.L_HI(net820));
 sg13g2_tiehi \clock_inst.min_b[0]$_DFFE_PP__821  (.L_HI(net821));
 sg13g2_tiehi \clock_inst.min_b[17]$_DFFE_PP__822  (.L_HI(net822));
 sg13g2_tiehi \clock_inst.min_b[19]$_DFFE_PP__823  (.L_HI(net823));
 sg13g2_tiehi \clock_inst.min_b[1]$_DFFE_PP__824  (.L_HI(net824));
 sg13g2_tiehi \clock_inst.min_b[20]$_DFFE_PP__825  (.L_HI(net825));
 sg13g2_tiehi \clock_inst.min_b[21]$_DFFE_PP__826  (.L_HI(net826));
 sg13g2_tiehi \clock_inst.min_b[22]$_DFFE_PP__827  (.L_HI(net827));
 sg13g2_tiehi \clock_inst.min_b[23]$_DFFE_PP__828  (.L_HI(net828));
 sg13g2_tiehi \clock_inst.min_b[2]$_DFFE_PP__829  (.L_HI(net829));
 sg13g2_tiehi \clock_inst.min_b[35]$_DFFE_PP__830  (.L_HI(net830));
 sg13g2_tiehi \clock_inst.min_b[36]$_DFFE_PP__831  (.L_HI(net831));
 sg13g2_tiehi \clock_inst.min_b[37]$_DFFE_PP__832  (.L_HI(net832));
 sg13g2_tiehi \clock_inst.min_b[38]$_DFFE_PP__833  (.L_HI(net833));
 sg13g2_tiehi \clock_inst.min_b[39]$_DFFE_PP__834  (.L_HI(net834));
 sg13g2_tiehi \clock_inst.min_b[3]$_DFFE_PP__835  (.L_HI(net835));
 sg13g2_tiehi \clock_inst.min_b[40]$_DFFE_PP__836  (.L_HI(net836));
 sg13g2_tiehi \clock_inst.min_b[41]$_DFFE_PP__837  (.L_HI(net837));
 sg13g2_tiehi \clock_inst.min_b[42]$_DFFE_PP__838  (.L_HI(net838));
 sg13g2_tiehi \clock_inst.min_b[43]$_DFFE_PP__839  (.L_HI(net839));
 sg13g2_tiehi \clock_inst.min_b[44]$_DFFE_PP__840  (.L_HI(net840));
 sg13g2_tiehi \clock_inst.min_b[4]$_DFFE_PP__841  (.L_HI(net841));
 sg13g2_tiehi \clock_inst.min_b[5]$_DFFE_PP__842  (.L_HI(net842));
 sg13g2_tiehi \clock_inst.min_b[6]$_DFFE_PP__843  (.L_HI(net843));
 sg13g2_tiehi \clock_inst.min_b[7]$_DFFE_PP__844  (.L_HI(net844));
 sg13g2_tiehi \clock_inst.min_b[8]$_DFFE_PP__845  (.L_HI(net845));
 sg13g2_tiehi \clock_inst.min_c[0]$_DFFE_PP__846  (.L_HI(net846));
 sg13g2_tiehi \clock_inst.min_c[10]$_DFFE_PP__847  (.L_HI(net847));
 sg13g2_tiehi \clock_inst.min_c[11]$_DFFE_PP__848  (.L_HI(net848));
 sg13g2_tiehi \clock_inst.min_c[12]$_DFFE_PP__849  (.L_HI(net849));
 sg13g2_tiehi \clock_inst.min_c[13]$_DFFE_PP__850  (.L_HI(net850));
 sg13g2_tiehi \clock_inst.min_c[14]$_DFFE_PP__851  (.L_HI(net851));
 sg13g2_tiehi \clock_inst.min_c[15]$_DFFE_PP__852  (.L_HI(net852));
 sg13g2_tiehi \clock_inst.min_c[16]$_DFFE_PP__853  (.L_HI(net853));
 sg13g2_tiehi \clock_inst.min_c[17]$_DFFE_PP__854  (.L_HI(net854));
 sg13g2_tiehi \clock_inst.min_c[19]$_DFFE_PP__855  (.L_HI(net855));
 sg13g2_tiehi \clock_inst.min_c[1]$_DFFE_PP__856  (.L_HI(net856));
 sg13g2_tiehi \clock_inst.min_c[21]$_DFFE_PP__857  (.L_HI(net857));
 sg13g2_tiehi \clock_inst.min_c[22]$_DFFE_PP__858  (.L_HI(net858));
 sg13g2_tiehi \clock_inst.min_c[23]$_DFFE_PP__859  (.L_HI(net859));
 sg13g2_tiehi \clock_inst.min_c[24]$_DFFE_PP__860  (.L_HI(net860));
 sg13g2_tiehi \clock_inst.min_c[25]$_DFFE_PP__861  (.L_HI(net861));
 sg13g2_tiehi \clock_inst.min_c[26]$_DFFE_PP__862  (.L_HI(net862));
 sg13g2_tiehi \clock_inst.min_c[27]$_DFFE_PP__863  (.L_HI(net863));
 sg13g2_tiehi \clock_inst.min_c[28]$_DFFE_PP__864  (.L_HI(net864));
 sg13g2_tiehi \clock_inst.min_c[29]$_DFFE_PP__865  (.L_HI(net865));
 sg13g2_tiehi \clock_inst.min_c[2]$_DFFE_PP__866  (.L_HI(net866));
 sg13g2_tiehi \clock_inst.min_c[30]$_DFFE_PP__867  (.L_HI(net867));
 sg13g2_tiehi \clock_inst.min_c[31]$_DFFE_PP__868  (.L_HI(net868));
 sg13g2_tiehi \clock_inst.min_c[32]$_DFFE_PP__869  (.L_HI(net869));
 sg13g2_tiehi \clock_inst.min_c[35]$_DFFE_PP__870  (.L_HI(net870));
 sg13g2_tiehi \clock_inst.min_c[36]$_DFFE_PP__871  (.L_HI(net871));
 sg13g2_tiehi \clock_inst.min_c[37]$_DFFE_PP__872  (.L_HI(net872));
 sg13g2_tiehi \clock_inst.min_c[38]$_DFFE_PP__873  (.L_HI(net873));
 sg13g2_tiehi \clock_inst.min_c[39]$_DFFE_PP__874  (.L_HI(net874));
 sg13g2_tiehi \clock_inst.min_c[3]$_DFFE_PP__875  (.L_HI(net875));
 sg13g2_tiehi \clock_inst.min_c[40]$_DFFE_PP__876  (.L_HI(net876));
 sg13g2_tiehi \clock_inst.min_c[41]$_DFFE_PP__877  (.L_HI(net877));
 sg13g2_tiehi \clock_inst.min_c[42]$_DFFE_PP__878  (.L_HI(net878));
 sg13g2_tiehi \clock_inst.min_c[43]$_DFFE_PP__879  (.L_HI(net879));
 sg13g2_tiehi \clock_inst.min_c[44]$_DFFE_PP__880  (.L_HI(net880));
 sg13g2_tiehi \clock_inst.min_c[45]$_DFFE_PP__881  (.L_HI(net881));
 sg13g2_tiehi \clock_inst.min_c[46]$_DFFE_PP__882  (.L_HI(net882));
 sg13g2_tiehi \clock_inst.min_c[47]$_DFFE_PP__883  (.L_HI(net883));
 sg13g2_tiehi \clock_inst.min_c[48]$_DFFE_PP__884  (.L_HI(net884));
 sg13g2_tiehi \clock_inst.min_c[49]$_DFFE_PP__885  (.L_HI(net885));
 sg13g2_tiehi \clock_inst.min_c[4]$_DFFE_PP__886  (.L_HI(net886));
 sg13g2_tiehi \clock_inst.min_c[50]$_DFFE_PP__887  (.L_HI(net887));
 sg13g2_tiehi \clock_inst.min_c[51]$_DFFE_PP__888  (.L_HI(net888));
 sg13g2_tiehi \clock_inst.min_c[52]$_DFFE_PP__889  (.L_HI(net889));
 sg13g2_tiehi \clock_inst.min_c[53]$_DFFE_PP__890  (.L_HI(net890));
 sg13g2_tiehi \clock_inst.min_c[5]$_DFFE_PP__891  (.L_HI(net891));
 sg13g2_tiehi \clock_inst.min_c[6]$_DFFE_PP__892  (.L_HI(net892));
 sg13g2_tiehi \clock_inst.min_c[7]$_DFFE_PP__893  (.L_HI(net893));
 sg13g2_tiehi \clock_inst.min_c[8]$_DFFE_PP__894  (.L_HI(net894));
 sg13g2_tiehi \clock_inst.min_c[9]$_DFFE_PP__895  (.L_HI(net895));
 sg13g2_tiehi \clock_inst.min_tile.e0[0]$_DFFE_PP__896  (.L_HI(net896));
 sg13g2_tiehi \clock_inst.min_tile.e0[10]$_DFFE_PP__897  (.L_HI(net897));
 sg13g2_tiehi \clock_inst.min_tile.e0[11]$_DFFE_PP__898  (.L_HI(net898));
 sg13g2_tiehi \clock_inst.min_tile.e0[12]$_DFFE_PP__899  (.L_HI(net899));
 sg13g2_tiehi \clock_inst.min_tile.e0[13]$_DFFE_PP__900  (.L_HI(net900));
 sg13g2_tiehi \clock_inst.min_tile.e0[14]$_DFFE_PP__901  (.L_HI(net901));
 sg13g2_tiehi \clock_inst.min_tile.e0[15]$_DFFE_PP__902  (.L_HI(net902));
 sg13g2_tiehi \clock_inst.min_tile.e0[16]$_DFFE_PP__903  (.L_HI(net903));
 sg13g2_tiehi \clock_inst.min_tile.e0[17]$_DFFE_PP__904  (.L_HI(net904));
 sg13g2_tiehi \clock_inst.min_tile.e0[18]$_DFFE_PP__905  (.L_HI(net905));
 sg13g2_tiehi \clock_inst.min_tile.e0[19]$_DFFE_PP__906  (.L_HI(net906));
 sg13g2_tiehi \clock_inst.min_tile.e0[1]$_DFFE_PP__907  (.L_HI(net907));
 sg13g2_tiehi \clock_inst.min_tile.e0[20]$_SDFFCE_PP0P__908  (.L_HI(net908));
 sg13g2_tiehi \clock_inst.min_tile.e0[21]$_DFFE_PP__909  (.L_HI(net909));
 sg13g2_tiehi \clock_inst.min_tile.e0[22]$_DFFE_PP__910  (.L_HI(net910));
 sg13g2_tiehi \clock_inst.min_tile.e0[23]$_DFFE_PP__911  (.L_HI(net911));
 sg13g2_tiehi \clock_inst.min_tile.e0[24]$_DFFE_PP__912  (.L_HI(net912));
 sg13g2_tiehi \clock_inst.min_tile.e0[25]$_DFFE_PP__913  (.L_HI(net913));
 sg13g2_tiehi \clock_inst.min_tile.e0[26]$_DFFE_PP__914  (.L_HI(net914));
 sg13g2_tiehi \clock_inst.min_tile.e0[27]$_DFFE_PP__915  (.L_HI(net915));
 sg13g2_tiehi \clock_inst.min_tile.e0[28]$_DFFE_PP__916  (.L_HI(net916));
 sg13g2_tiehi \clock_inst.min_tile.e0[29]$_DFFE_PP__917  (.L_HI(net917));
 sg13g2_tiehi \clock_inst.min_tile.e0[2]$_DFFE_PP__918  (.L_HI(net918));
 sg13g2_tiehi \clock_inst.min_tile.e0[30]$_DFFE_PP__919  (.L_HI(net919));
 sg13g2_tiehi \clock_inst.min_tile.e0[31]$_DFFE_PP__920  (.L_HI(net920));
 sg13g2_tiehi \clock_inst.min_tile.e0[32]$_DFFE_PP__921  (.L_HI(net921));
 sg13g2_tiehi \clock_inst.min_tile.e0[33]$_DFFE_PP__922  (.L_HI(net922));
 sg13g2_tiehi \clock_inst.min_tile.e0[34]$_DFFE_PP__923  (.L_HI(net923));
 sg13g2_tiehi \clock_inst.min_tile.e0[35]$_DFFE_PP__924  (.L_HI(net924));
 sg13g2_tiehi \clock_inst.min_tile.e0[36]$_DFFE_PP__925  (.L_HI(net925));
 sg13g2_tiehi \clock_inst.min_tile.e0[37]$_DFFE_PP__926  (.L_HI(net926));
 sg13g2_tiehi \clock_inst.min_tile.e0[38]$_DFFE_PP__927  (.L_HI(net927));
 sg13g2_tiehi \clock_inst.min_tile.e0[39]$_DFFE_PP__928  (.L_HI(net928));
 sg13g2_tiehi \clock_inst.min_tile.e0[3]$_DFFE_PP__929  (.L_HI(net929));
 sg13g2_tiehi \clock_inst.min_tile.e0[40]$_DFFE_PP__930  (.L_HI(net930));
 sg13g2_tiehi \clock_inst.min_tile.e0[41]$_DFFE_PP__931  (.L_HI(net931));
 sg13g2_tiehi \clock_inst.min_tile.e0[42]$_DFFE_PP__932  (.L_HI(net932));
 sg13g2_tiehi \clock_inst.min_tile.e0[43]$_DFFE_PP__933  (.L_HI(net933));
 sg13g2_tiehi \clock_inst.min_tile.e0[44]$_DFFE_PP__934  (.L_HI(net934));
 sg13g2_tiehi \clock_inst.min_tile.e0[45]$_DFFE_PP__935  (.L_HI(net935));
 sg13g2_tiehi \clock_inst.min_tile.e0[46]$_DFFE_PP__936  (.L_HI(net936));
 sg13g2_tiehi \clock_inst.min_tile.e0[47]$_DFFE_PP__937  (.L_HI(net937));
 sg13g2_tiehi \clock_inst.min_tile.e0[48]$_DFFE_PP__938  (.L_HI(net938));
 sg13g2_tiehi \clock_inst.min_tile.e0[49]$_DFFE_PP__939  (.L_HI(net939));
 sg13g2_tiehi \clock_inst.min_tile.e0[4]$_DFFE_PP__940  (.L_HI(net940));
 sg13g2_tiehi \clock_inst.min_tile.e0[50]$_DFFE_PP__941  (.L_HI(net941));
 sg13g2_tiehi \clock_inst.min_tile.e0[51]$_DFFE_PP__942  (.L_HI(net942));
 sg13g2_tiehi \clock_inst.min_tile.e0[52]$_DFFE_PP__943  (.L_HI(net943));
 sg13g2_tiehi \clock_inst.min_tile.e0[53]$_DFFE_PP__944  (.L_HI(net944));
 sg13g2_tiehi \clock_inst.min_tile.e0[5]$_DFFE_PP__945  (.L_HI(net945));
 sg13g2_tiehi \clock_inst.min_tile.e0[6]$_DFFE_PP__946  (.L_HI(net946));
 sg13g2_tiehi \clock_inst.min_tile.e0[7]$_DFFE_PP__947  (.L_HI(net947));
 sg13g2_tiehi \clock_inst.min_tile.e0[8]$_DFFE_PP__948  (.L_HI(net948));
 sg13g2_tiehi \clock_inst.min_tile.e0[9]$_DFFE_PP__949  (.L_HI(net949));
 sg13g2_tiehi \clock_inst.min_tile.e[0]$_DFFE_PP__950  (.L_HI(net950));
 sg13g2_tiehi \clock_inst.min_tile.e[10]$_DFFE_PP__951  (.L_HI(net951));
 sg13g2_tiehi \clock_inst.min_tile.e[11]$_DFFE_PP__952  (.L_HI(net952));
 sg13g2_tiehi \clock_inst.min_tile.e[12]$_DFFE_PP__953  (.L_HI(net953));
 sg13g2_tiehi \clock_inst.min_tile.e[13]$_DFFE_PP__954  (.L_HI(net954));
 sg13g2_tiehi \clock_inst.min_tile.e[14]$_DFFE_PP__955  (.L_HI(net955));
 sg13g2_tiehi \clock_inst.min_tile.e[15]$_DFFE_PP__956  (.L_HI(net956));
 sg13g2_tiehi \clock_inst.min_tile.e[16]$_DFFE_PP__957  (.L_HI(net957));
 sg13g2_tiehi \clock_inst.min_tile.e[17]$_DFFE_PP__958  (.L_HI(net958));
 sg13g2_tiehi \clock_inst.min_tile.e[18]$_DFFE_PP__959  (.L_HI(net959));
 sg13g2_tiehi \clock_inst.min_tile.e[19]$_DFFE_PP__960  (.L_HI(net960));
 sg13g2_tiehi \clock_inst.min_tile.e[1]$_DFFE_PP__961  (.L_HI(net961));
 sg13g2_tiehi \clock_inst.min_tile.e[20]$_SDFFCE_PP0P__962  (.L_HI(net962));
 sg13g2_tiehi \clock_inst.min_tile.e[21]$_DFFE_PP__963  (.L_HI(net963));
 sg13g2_tiehi \clock_inst.min_tile.e[22]$_DFFE_PP__964  (.L_HI(net964));
 sg13g2_tiehi \clock_inst.min_tile.e[23]$_DFFE_PP__965  (.L_HI(net965));
 sg13g2_tiehi \clock_inst.min_tile.e[24]$_DFFE_PP__966  (.L_HI(net966));
 sg13g2_tiehi \clock_inst.min_tile.e[25]$_DFFE_PP__967  (.L_HI(net967));
 sg13g2_tiehi \clock_inst.min_tile.e[26]$_DFFE_PP__968  (.L_HI(net968));
 sg13g2_tiehi \clock_inst.min_tile.e[27]$_DFFE_PP__969  (.L_HI(net969));
 sg13g2_tiehi \clock_inst.min_tile.e[28]$_DFFE_PP__970  (.L_HI(net970));
 sg13g2_tiehi \clock_inst.min_tile.e[29]$_DFFE_PP__971  (.L_HI(net971));
 sg13g2_tiehi \clock_inst.min_tile.e[2]$_DFFE_PP__972  (.L_HI(net972));
 sg13g2_tiehi \clock_inst.min_tile.e[30]$_DFFE_PP__973  (.L_HI(net973));
 sg13g2_tiehi \clock_inst.min_tile.e[31]$_DFFE_PP__974  (.L_HI(net974));
 sg13g2_tiehi \clock_inst.min_tile.e[32]$_DFFE_PP__975  (.L_HI(net975));
 sg13g2_tiehi \clock_inst.min_tile.e[33]$_DFFE_PP__976  (.L_HI(net976));
 sg13g2_tiehi \clock_inst.min_tile.e[34]$_DFFE_PP__977  (.L_HI(net977));
 sg13g2_tiehi \clock_inst.min_tile.e[35]$_DFFE_PP__978  (.L_HI(net978));
 sg13g2_tiehi \clock_inst.min_tile.e[36]$_DFFE_PP__979  (.L_HI(net979));
 sg13g2_tiehi \clock_inst.min_tile.e[37]$_DFFE_PP__980  (.L_HI(net980));
 sg13g2_tiehi \clock_inst.min_tile.e[38]$_DFFE_PP__981  (.L_HI(net981));
 sg13g2_tiehi \clock_inst.min_tile.e[39]$_DFFE_PP__982  (.L_HI(net982));
 sg13g2_tiehi \clock_inst.min_tile.e[3]$_DFFE_PP__983  (.L_HI(net983));
 sg13g2_tiehi \clock_inst.min_tile.e[40]$_DFFE_PP__984  (.L_HI(net984));
 sg13g2_tiehi \clock_inst.min_tile.e[41]$_DFFE_PP__985  (.L_HI(net985));
 sg13g2_tiehi \clock_inst.min_tile.e[42]$_DFFE_PP__986  (.L_HI(net986));
 sg13g2_tiehi \clock_inst.min_tile.e[43]$_DFFE_PP__987  (.L_HI(net987));
 sg13g2_tiehi \clock_inst.min_tile.e[44]$_DFFE_PP__988  (.L_HI(net988));
 sg13g2_tiehi \clock_inst.min_tile.e[45]$_DFFE_PP__989  (.L_HI(net989));
 sg13g2_tiehi \clock_inst.min_tile.e[46]$_DFFE_PP__990  (.L_HI(net990));
 sg13g2_tiehi \clock_inst.min_tile.e[47]$_DFFE_PP__991  (.L_HI(net991));
 sg13g2_tiehi \clock_inst.min_tile.e[48]$_DFFE_PP__992  (.L_HI(net992));
 sg13g2_tiehi \clock_inst.min_tile.e[49]$_DFFE_PP__993  (.L_HI(net993));
 sg13g2_tiehi \clock_inst.min_tile.e[4]$_DFFE_PP__994  (.L_HI(net994));
 sg13g2_tiehi \clock_inst.min_tile.e[50]$_DFFE_PP__995  (.L_HI(net995));
 sg13g2_tiehi \clock_inst.min_tile.e[51]$_DFFE_PP__996  (.L_HI(net996));
 sg13g2_tiehi \clock_inst.min_tile.e[52]$_DFFE_PP__997  (.L_HI(net997));
 sg13g2_tiehi \clock_inst.min_tile.e[53]$_DFFE_PP__998  (.L_HI(net998));
 sg13g2_tiehi \clock_inst.min_tile.e[5]$_DFFE_PP__999  (.L_HI(net999));
 sg13g2_tiehi \clock_inst.min_tile.e[6]$_DFFE_PP__1000  (.L_HI(net1000));
 sg13g2_tiehi \clock_inst.min_tile.e[7]$_DFFE_PP__1001  (.L_HI(net1001));
 sg13g2_tiehi \clock_inst.min_tile.e[8]$_DFFE_PP__1002  (.L_HI(net1002));
 sg13g2_tiehi \clock_inst.min_tile.e[9]$_DFFE_PP__1003  (.L_HI(net1003));
 sg13g2_tiehi \clock_inst.minute[0]$_SDFFE_PP0N__1004  (.L_HI(net1004));
 sg13g2_tiehi \clock_inst.minute[1]$_SDFFE_PN1P__1005  (.L_HI(net1005));
 sg13g2_tiehi \clock_inst.minute[2]$_SDFFE_PP0N__1006  (.L_HI(net1006));
 sg13g2_tiehi \clock_inst.minute[3]$_SDFFE_PN1P__1007  (.L_HI(net1007));
 sg13g2_tiehi \clock_inst.minute[4]$_SDFFE_PN1P__1008  (.L_HI(net1008));
 sg13g2_tiehi \clock_inst.minute[5]$_SDFFE_PP0N__1009  (.L_HI(net1009));
 sg13g2_tiehi \clock_inst.sec_a[0]$_DFFE_PP__1010  (.L_HI(net1010));
 sg13g2_tiehi \clock_inst.sec_a[17]$_DFFE_PP__1011  (.L_HI(net1011));
 sg13g2_tiehi \clock_inst.sec_a[18]$_DFFE_PP__1012  (.L_HI(net1012));
 sg13g2_tiehi \clock_inst.sec_a[19]$_DFFE_PP__1013  (.L_HI(net1013));
 sg13g2_tiehi \clock_inst.sec_a[1]$_DFFE_PP__1014  (.L_HI(net1014));
 sg13g2_tiehi \clock_inst.sec_a[20]$_DFFE_PP__1015  (.L_HI(net1015));
 sg13g2_tiehi \clock_inst.sec_a[2]$_DFFE_PP__1016  (.L_HI(net1016));
 sg13g2_tiehi \clock_inst.sec_a[35]$_DFFE_PP__1017  (.L_HI(net1017));
 sg13g2_tiehi \clock_inst.sec_a[36]$_DFFE_PP__1018  (.L_HI(net1018));
 sg13g2_tiehi \clock_inst.sec_a[37]$_DFFE_PP__1019  (.L_HI(net1019));
 sg13g2_tiehi \clock_inst.sec_a[38]$_DFFE_PP__1020  (.L_HI(net1020));
 sg13g2_tiehi \clock_inst.sec_a[39]$_DFFE_PP__1021  (.L_HI(net1021));
 sg13g2_tiehi \clock_inst.sec_a[3]$_DFFE_PP__1022  (.L_HI(net1022));
 sg13g2_tiehi \clock_inst.sec_a[40]$_DFFE_PP__1023  (.L_HI(net1023));
 sg13g2_tiehi \clock_inst.sec_a[41]$_DFFE_PP__1024  (.L_HI(net1024));
 sg13g2_tiehi \clock_inst.sec_a[42]$_DFFE_PP__1025  (.L_HI(net1025));
 sg13g2_tiehi \clock_inst.sec_a[43]$_DFFE_PP__1026  (.L_HI(net1026));
 sg13g2_tiehi \clock_inst.sec_a[4]$_DFFE_PP__1027  (.L_HI(net1027));
 sg13g2_tiehi \clock_inst.sec_a[52]$_DFFE_PP__1028  (.L_HI(net1028));
 sg13g2_tiehi \clock_inst.sec_a[5]$_DFFE_PP__1029  (.L_HI(net1029));
 sg13g2_tiehi \clock_inst.sec_a[6]$_DFFE_PP__1030  (.L_HI(net1030));
 sg13g2_tiehi \clock_inst.sec_a[7]$_DFFE_PP__1031  (.L_HI(net1031));
 sg13g2_tiehi \clock_inst.sec_b[0]$_DFFE_PP__1032  (.L_HI(net1032));
 sg13g2_tiehi \clock_inst.sec_b[17]$_DFFE_PP__1033  (.L_HI(net1033));
 sg13g2_tiehi \clock_inst.sec_b[19]$_DFFE_PP__1034  (.L_HI(net1034));
 sg13g2_tiehi \clock_inst.sec_b[1]$_DFFE_PP__1035  (.L_HI(net1035));
 sg13g2_tiehi \clock_inst.sec_b[20]$_DFFE_PP__1036  (.L_HI(net1036));
 sg13g2_tiehi \clock_inst.sec_b[2]$_DFFE_PP__1037  (.L_HI(net1037));
 sg13g2_tiehi \clock_inst.sec_b[35]$_DFFE_PP__1038  (.L_HI(net1038));
 sg13g2_tiehi \clock_inst.sec_b[36]$_DFFE_PP__1039  (.L_HI(net1039));
 sg13g2_tiehi \clock_inst.sec_b[37]$_DFFE_PP__1040  (.L_HI(net1040));
 sg13g2_tiehi \clock_inst.sec_b[38]$_DFFE_PP__1041  (.L_HI(net1041));
 sg13g2_tiehi \clock_inst.sec_b[39]$_DFFE_PP__1042  (.L_HI(net1042));
 sg13g2_tiehi \clock_inst.sec_b[3]$_DFFE_PP__1043  (.L_HI(net1043));
 sg13g2_tiehi \clock_inst.sec_b[40]$_DFFE_PP__1044  (.L_HI(net1044));
 sg13g2_tiehi \clock_inst.sec_b[41]$_DFFE_PP__1045  (.L_HI(net1045));
 sg13g2_tiehi \clock_inst.sec_b[42]$_DFFE_PP__1046  (.L_HI(net1046));
 sg13g2_tiehi \clock_inst.sec_b[43]$_DFFE_PP__1047  (.L_HI(net1047));
 sg13g2_tiehi \clock_inst.sec_b[4]$_DFFE_PP__1048  (.L_HI(net1048));
 sg13g2_tiehi \clock_inst.sec_b[5]$_DFFE_PP__1049  (.L_HI(net1049));
 sg13g2_tiehi \clock_inst.sec_b[6]$_DFFE_PP__1050  (.L_HI(net1050));
 sg13g2_tiehi \clock_inst.sec_b[7]$_DFFE_PP__1051  (.L_HI(net1051));
 sg13g2_tiehi \clock_inst.sec_c[0]$_DFFE_PP__1052  (.L_HI(net1052));
 sg13g2_tiehi \clock_inst.sec_c[10]$_DFFE_PP__1053  (.L_HI(net1053));
 sg13g2_tiehi \clock_inst.sec_c[11]$_DFFE_PP__1054  (.L_HI(net1054));
 sg13g2_tiehi \clock_inst.sec_c[12]$_DFFE_PP__1055  (.L_HI(net1055));
 sg13g2_tiehi \clock_inst.sec_c[13]$_DFFE_PP__1056  (.L_HI(net1056));
 sg13g2_tiehi \clock_inst.sec_c[14]$_DFFE_PP__1057  (.L_HI(net1057));
 sg13g2_tiehi \clock_inst.sec_c[15]$_DFFE_PP__1058  (.L_HI(net1058));
 sg13g2_tiehi \clock_inst.sec_c[16]$_DFFE_PP__1059  (.L_HI(net1059));
 sg13g2_tiehi \clock_inst.sec_c[17]$_DFFE_PP__1060  (.L_HI(net1060));
 sg13g2_tiehi \clock_inst.sec_c[19]$_DFFE_PP__1061  (.L_HI(net1061));
 sg13g2_tiehi \clock_inst.sec_c[1]$_DFFE_PP__1062  (.L_HI(net1062));
 sg13g2_tiehi \clock_inst.sec_c[20]$_DFFE_PP__1063  (.L_HI(net1063));
 sg13g2_tiehi \clock_inst.sec_c[21]$_DFFE_PP__1064  (.L_HI(net1064));
 sg13g2_tiehi \clock_inst.sec_c[22]$_DFFE_PP__1065  (.L_HI(net1065));
 sg13g2_tiehi \clock_inst.sec_c[23]$_DFFE_PP__1066  (.L_HI(net1066));
 sg13g2_tiehi \clock_inst.sec_c[24]$_DFFE_PP__1067  (.L_HI(net1067));
 sg13g2_tiehi \clock_inst.sec_c[25]$_DFFE_PP__1068  (.L_HI(net1068));
 sg13g2_tiehi \clock_inst.sec_c[26]$_DFFE_PP__1069  (.L_HI(net1069));
 sg13g2_tiehi \clock_inst.sec_c[27]$_DFFE_PP__1070  (.L_HI(net1070));
 sg13g2_tiehi \clock_inst.sec_c[28]$_DFFE_PP__1071  (.L_HI(net1071));
 sg13g2_tiehi \clock_inst.sec_c[29]$_DFFE_PP__1072  (.L_HI(net1072));
 sg13g2_tiehi \clock_inst.sec_c[2]$_DFFE_PP__1073  (.L_HI(net1073));
 sg13g2_tiehi \clock_inst.sec_c[35]$_DFFE_PP__1074  (.L_HI(net1074));
 sg13g2_tiehi \clock_inst.sec_c[36]$_DFFE_PP__1075  (.L_HI(net1075));
 sg13g2_tiehi \clock_inst.sec_c[37]$_DFFE_PP__1076  (.L_HI(net1076));
 sg13g2_tiehi \clock_inst.sec_c[38]$_DFFE_PP__1077  (.L_HI(net1077));
 sg13g2_tiehi \clock_inst.sec_c[39]$_DFFE_PP__1078  (.L_HI(net1078));
 sg13g2_tiehi \clock_inst.sec_c[3]$_DFFE_PP__1079  (.L_HI(net1079));
 sg13g2_tiehi \clock_inst.sec_c[40]$_DFFE_PP__1080  (.L_HI(net1080));
 sg13g2_tiehi \clock_inst.sec_c[41]$_DFFE_PP__1081  (.L_HI(net1081));
 sg13g2_tiehi \clock_inst.sec_c[42]$_DFFE_PP__1082  (.L_HI(net1082));
 sg13g2_tiehi \clock_inst.sec_c[43]$_DFFE_PP__1083  (.L_HI(net1083));
 sg13g2_tiehi \clock_inst.sec_c[44]$_DFFE_PP__1084  (.L_HI(net1084));
 sg13g2_tiehi \clock_inst.sec_c[45]$_DFFE_PP__1085  (.L_HI(net1085));
 sg13g2_tiehi \clock_inst.sec_c[46]$_DFFE_PP__1086  (.L_HI(net1086));
 sg13g2_tiehi \clock_inst.sec_c[47]$_DFFE_PP__1087  (.L_HI(net1087));
 sg13g2_tiehi \clock_inst.sec_c[48]$_DFFE_PP__1088  (.L_HI(net1088));
 sg13g2_tiehi \clock_inst.sec_c[49]$_DFFE_PP__1089  (.L_HI(net1089));
 sg13g2_tiehi \clock_inst.sec_c[4]$_DFFE_PP__1090  (.L_HI(net1090));
 sg13g2_tiehi \clock_inst.sec_c[50]$_DFFE_PP__1091  (.L_HI(net1091));
 sg13g2_tiehi \clock_inst.sec_c[51]$_DFFE_PP__1092  (.L_HI(net1092));
 sg13g2_tiehi \clock_inst.sec_c[52]$_DFFE_PP__1093  (.L_HI(net1093));
 sg13g2_tiehi \clock_inst.sec_c[53]$_DFFE_PP__1094  (.L_HI(net1094));
 sg13g2_tiehi \clock_inst.sec_c[5]$_DFFE_PP__1095  (.L_HI(net1095));
 sg13g2_tiehi \clock_inst.sec_c[6]$_DFFE_PP__1096  (.L_HI(net1096));
 sg13g2_tiehi \clock_inst.sec_c[7]$_DFFE_PP__1097  (.L_HI(net1097));
 sg13g2_tiehi \clock_inst.sec_c[8]$_DFFE_PP__1098  (.L_HI(net1098));
 sg13g2_tiehi \clock_inst.sec_c[9]$_DFFE_PP__1099  (.L_HI(net1099));
 sg13g2_tiehi \clock_inst.sec_tile.e0[0]$_DFFE_PP__1100  (.L_HI(net1100));
 sg13g2_tiehi \clock_inst.sec_tile.e0[10]$_DFFE_PP__1101  (.L_HI(net1101));
 sg13g2_tiehi \clock_inst.sec_tile.e0[11]$_DFFE_PP__1102  (.L_HI(net1102));
 sg13g2_tiehi \clock_inst.sec_tile.e0[12]$_DFFE_PP__1103  (.L_HI(net1103));
 sg13g2_tiehi \clock_inst.sec_tile.e0[13]$_DFFE_PP__1104  (.L_HI(net1104));
 sg13g2_tiehi \clock_inst.sec_tile.e0[14]$_DFFE_PP__1105  (.L_HI(net1105));
 sg13g2_tiehi \clock_inst.sec_tile.e0[15]$_DFFE_PP__1106  (.L_HI(net1106));
 sg13g2_tiehi \clock_inst.sec_tile.e0[16]$_DFFE_PP__1107  (.L_HI(net1107));
 sg13g2_tiehi \clock_inst.sec_tile.e0[17]$_DFFE_PP__1108  (.L_HI(net1108));
 sg13g2_tiehi \clock_inst.sec_tile.e0[18]$_DFFE_PP__1109  (.L_HI(net1109));
 sg13g2_tiehi \clock_inst.sec_tile.e0[19]$_DFFE_PP__1110  (.L_HI(net1110));
 sg13g2_tiehi \clock_inst.sec_tile.e0[1]$_DFFE_PP__1111  (.L_HI(net1111));
 sg13g2_tiehi \clock_inst.sec_tile.e0[20]$_DFFE_PP__1112  (.L_HI(net1112));
 sg13g2_tiehi \clock_inst.sec_tile.e0[21]$_DFFE_PP__1113  (.L_HI(net1113));
 sg13g2_tiehi \clock_inst.sec_tile.e0[22]$_DFFE_PP__1114  (.L_HI(net1114));
 sg13g2_tiehi \clock_inst.sec_tile.e0[23]$_DFFE_PP__1115  (.L_HI(net1115));
 sg13g2_tiehi \clock_inst.sec_tile.e0[24]$_DFFE_PP__1116  (.L_HI(net1116));
 sg13g2_tiehi \clock_inst.sec_tile.e0[25]$_DFFE_PP__1117  (.L_HI(net1117));
 sg13g2_tiehi \clock_inst.sec_tile.e0[26]$_DFFE_PP__1118  (.L_HI(net1118));
 sg13g2_tiehi \clock_inst.sec_tile.e0[27]$_DFFE_PP__1119  (.L_HI(net1119));
 sg13g2_tiehi \clock_inst.sec_tile.e0[28]$_DFFE_PP__1120  (.L_HI(net1120));
 sg13g2_tiehi \clock_inst.sec_tile.e0[29]$_DFFE_PP__1121  (.L_HI(net1121));
 sg13g2_tiehi \clock_inst.sec_tile.e0[2]$_DFFE_PP__1122  (.L_HI(net1122));
 sg13g2_tiehi \clock_inst.sec_tile.e0[30]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \clock_inst.sec_tile.e0[31]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \clock_inst.sec_tile.e0[32]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \clock_inst.sec_tile.e0[33]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \clock_inst.sec_tile.e0[34]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \clock_inst.sec_tile.e0[35]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \clock_inst.sec_tile.e0[36]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \clock_inst.sec_tile.e0[37]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \clock_inst.sec_tile.e0[38]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \clock_inst.sec_tile.e0[39]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \clock_inst.sec_tile.e0[3]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \clock_inst.sec_tile.e0[40]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \clock_inst.sec_tile.e0[41]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \clock_inst.sec_tile.e0[42]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \clock_inst.sec_tile.e0[43]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \clock_inst.sec_tile.e0[44]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \clock_inst.sec_tile.e0[45]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \clock_inst.sec_tile.e0[46]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \clock_inst.sec_tile.e0[47]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \clock_inst.sec_tile.e0[48]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \clock_inst.sec_tile.e0[49]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \clock_inst.sec_tile.e0[4]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \clock_inst.sec_tile.e0[50]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \clock_inst.sec_tile.e0[51]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \clock_inst.sec_tile.e0[52]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \clock_inst.sec_tile.e0[53]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \clock_inst.sec_tile.e0[5]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \clock_inst.sec_tile.e0[6]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \clock_inst.sec_tile.e0[7]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \clock_inst.sec_tile.e0[8]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \clock_inst.sec_tile.e0[9]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \clock_inst.sec_tile.e[0]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \clock_inst.sec_tile.e[10]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \clock_inst.sec_tile.e[11]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \clock_inst.sec_tile.e[12]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \clock_inst.sec_tile.e[13]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \clock_inst.sec_tile.e[14]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \clock_inst.sec_tile.e[15]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \clock_inst.sec_tile.e[16]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \clock_inst.sec_tile.e[17]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \clock_inst.sec_tile.e[18]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \clock_inst.sec_tile.e[19]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \clock_inst.sec_tile.e[1]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \clock_inst.sec_tile.e[20]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \clock_inst.sec_tile.e[21]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \clock_inst.sec_tile.e[22]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \clock_inst.sec_tile.e[23]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \clock_inst.sec_tile.e[24]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \clock_inst.sec_tile.e[25]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \clock_inst.sec_tile.e[26]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \clock_inst.sec_tile.e[27]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \clock_inst.sec_tile.e[28]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \clock_inst.sec_tile.e[29]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \clock_inst.sec_tile.e[2]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \clock_inst.sec_tile.e[30]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \clock_inst.sec_tile.e[31]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \clock_inst.sec_tile.e[32]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \clock_inst.sec_tile.e[33]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \clock_inst.sec_tile.e[34]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \clock_inst.sec_tile.e[35]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \clock_inst.sec_tile.e[36]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \clock_inst.sec_tile.e[37]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \clock_inst.sec_tile.e[38]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \clock_inst.sec_tile.e[39]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \clock_inst.sec_tile.e[3]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \clock_inst.sec_tile.e[40]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \clock_inst.sec_tile.e[41]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \clock_inst.sec_tile.e[42]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \clock_inst.sec_tile.e[43]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \clock_inst.sec_tile.e[44]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \clock_inst.sec_tile.e[45]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \clock_inst.sec_tile.e[46]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \clock_inst.sec_tile.e[47]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \clock_inst.sec_tile.e[48]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \clock_inst.sec_tile.e[49]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \clock_inst.sec_tile.e[4]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \clock_inst.sec_tile.e[50]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \clock_inst.sec_tile.e[51]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \clock_inst.sec_tile.e[52]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \clock_inst.sec_tile.e[53]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \clock_inst.sec_tile.e[5]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \clock_inst.sec_tile.e[6]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \clock_inst.sec_tile.e[7]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \clock_inst.sec_tile.e[8]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \clock_inst.sec_tile.e[9]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \clock_inst.second[0]$_SDFFE_PP0N__1208  (.L_HI(net1208));
 sg13g2_tiehi \clock_inst.second[1]$_SDFFE_PN1P__1209  (.L_HI(net1209));
 sg13g2_tiehi \clock_inst.second[2]$_SDFFE_PP0N__1210  (.L_HI(net1210));
 sg13g2_tiehi \clock_inst.second[3]$_SDFFE_PP0N__1211  (.L_HI(net1211));
 sg13g2_tiehi \clock_inst.second[4]$_SDFFE_PN1P__1212  (.L_HI(net1212));
 sg13g2_tiehi \clock_inst.second[5]$_SDFFE_PP0N__1213  (.L_HI(net1213));
 sg13g2_tiehi \clock_inst.vga_inst.vga_horizontal_blank_strobe$_SDFF_PN0__1214  (.L_HI(net1214));
 sg13g2_tiehi \clock_inst.vga_inst.vga_horizontal_visible$_SDFFE_PP1P__1215  (.L_HI(net1215));
 sg13g2_tiehi \clock_inst.vga_inst.vga_hs$_SDFFE_PP1N__1216  (.L_HI(net1216));
 sg13g2_tiehi \clock_inst.vga_inst.vga_vertical_blank_strobe$_SDFF_PN0__1217  (.L_HI(net1217));
 sg13g2_tiehi \clock_inst.vga_inst.vga_vertical_visible$_SDFFE_PN1P__1218  (.L_HI(net1218));
 sg13g2_tiehi \clock_inst.vga_inst.vga_vs$_SDFFE_PN1P__1219  (.L_HI(net1219));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[0]$_SDFF_PP0__1220  (.L_HI(net1220));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[1]$_SDFF_PP0__1221  (.L_HI(net1221));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[2]$_SDFF_PP0__1222  (.L_HI(net1222));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[3]$_SDFF_PP0__1223  (.L_HI(net1223));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[4]$_SDFF_PP0__1224  (.L_HI(net1224));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[5]$_SDFF_PP0__1225  (.L_HI(net1225));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[6]$_SDFF_PP0__1226  (.L_HI(net1226));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[7]$_SDFF_PP0__1227  (.L_HI(net1227));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[8]$_SDFF_PP0__1228  (.L_HI(net1228));
 sg13g2_tiehi \clock_inst.vga_inst.vga_x[9]$_SDFF_PP0__1229  (.L_HI(net1229));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[0]$_SDFFE_PN0P__1230  (.L_HI(net1230));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[1]$_SDFFE_PN0P__1231  (.L_HI(net1231));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[2]$_SDFFE_PN0P__1232  (.L_HI(net1232));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[3]$_SDFFE_PN0P__1233  (.L_HI(net1233));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[4]$_SDFFE_PN0P__1234  (.L_HI(net1234));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[5]$_SDFFE_PN0P__1235  (.L_HI(net1235));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[6]$_SDFFE_PN0P__1236  (.L_HI(net1236));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[7]$_SDFFE_PN0P__1237  (.L_HI(net1237));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[8]$_SDFFE_PN0P__1238  (.L_HI(net1238));
 sg13g2_tiehi \clock_inst.vga_inst.vga_y[9]$_SDFFE_PN0P__1239  (.L_HI(net1239));
 sg13g2_tiehi \clock_inst.vga_rgb[1]$_SDFF_PN0__1240  (.L_HI(net1240));
 sg13g2_tiehi \clock_inst.vga_rgb[3]$_SDFF_PN0__1241  (.L_HI(net1241));
 sg13g2_tiehi \clock_inst.vga_rgb[4]$_SDFF_PN0__1242  (.L_HI(net1242));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_4_0__f_clk (.X(clknet_4_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_4_1__f_clk (.X(clknet_4_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_4_2__f_clk (.X(clknet_4_2__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_4_3__f_clk (.X(clknet_4_3__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_4_4__f_clk (.X(clknet_4_4__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_4_5__f_clk (.X(clknet_4_5__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_4_6__f_clk (.X(clknet_4_6__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_4_7__f_clk (.X(clknet_4_7__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_4_8__f_clk (.X(clknet_4_8__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_4_9__f_clk (.X(clknet_4_9__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_4_10__f_clk (.X(clknet_4_10__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_4_11__f_clk (.X(clknet_4_11__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_4_12__f_clk (.X(clknet_4_12__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_4_13__f_clk (.X(clknet_4_13__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_4_14__f_clk (.X(clknet_4_14__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_4_15__f_clk (.X(clknet_4_15__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_9__leaf_clk));
 sg13g2_inv_2 clkload2 (.A(clknet_4_10__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_leaf_94_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_95_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_0_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_leaf_97_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_6_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_57_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_83_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_84_clk));
 sg13g2_buf_16 clkload13 (.A(clknet_leaf_10_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_14_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_15_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_20_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_21_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_73_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_74_clk));
 sg13g2_inv_4 clkload22 (.A(clknet_leaf_76_clk));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_80_clk));
 sg13g2_buf_8 clkload24 (.A(clknet_leaf_58_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_59_clk));
 sg13g2_buf_8 clkload26 (.A(clknet_leaf_60_clk));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_61_clk));
 sg13g2_buf_8 clkload28 (.A(clknet_leaf_81_clk));
 sg13g2_inv_2 clkload29 (.A(clknet_leaf_67_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_69_clk));
 sg13g2_inv_4 clkload31 (.A(clknet_leaf_70_clk));
 sg13g2_buf_8 clkload32 (.A(clknet_leaf_72_clk));
 sg13g2_inv_2 clkload33 (.A(clknet_leaf_51_clk));
 sg13g2_buf_16 clkload34 (.A(clknet_leaf_62_clk));
 sg13g2_buf_8 clkload35 (.A(clknet_leaf_64_clk));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_65_clk));
 sg13g2_inv_1 clkload37 (.A(clknet_leaf_30_clk));
 sg13g2_inv_4 clkload38 (.A(clknet_leaf_45_clk));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_54_clk));
 sg13g2_buf_16 clkload40 (.A(clknet_leaf_56_clk));
 sg13g2_inv_1 clkload41 (.A(clknet_leaf_31_clk));
 sg13g2_buf_8 clkload42 (.A(clknet_leaf_32_clk));
 sg13g2_inv_4 clkload43 (.A(clknet_leaf_46_clk));
 sg13g2_inv_2 clkload44 (.A(clknet_leaf_48_clk));
 sg13g2_inv_1 clkload45 (.A(clknet_leaf_41_clk));
 sg13g2_inv_4 clkload46 (.A(clknet_leaf_44_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00216_));
 sg13g2_antennanp ANTENNA_2 (.A(_00216_));
 sg13g2_antennanp ANTENNA_3 (.A(_00242_));
 sg13g2_antennanp ANTENNA_4 (.A(_00419_));
 sg13g2_antennanp ANTENNA_5 (.A(_00419_));
 sg13g2_antennanp ANTENNA_6 (.A(_00438_));
 sg13g2_antennanp ANTENNA_7 (.A(_00438_));
 sg13g2_antennanp ANTENNA_8 (.A(_00656_));
 sg13g2_antennanp ANTENNA_9 (.A(_00656_));
 sg13g2_antennanp ANTENNA_10 (.A(_00656_));
 sg13g2_antennanp ANTENNA_11 (.A(_00672_));
 sg13g2_antennanp ANTENNA_12 (.A(_00672_));
 sg13g2_antennanp ANTENNA_13 (.A(_00672_));
 sg13g2_antennanp ANTENNA_14 (.A(_00672_));
 sg13g2_antennanp ANTENNA_15 (.A(_00675_));
 sg13g2_antennanp ANTENNA_16 (.A(_00675_));
 sg13g2_antennanp ANTENNA_17 (.A(_00675_));
 sg13g2_antennanp ANTENNA_18 (.A(_00675_));
 sg13g2_antennanp ANTENNA_19 (.A(_00680_));
 sg13g2_antennanp ANTENNA_20 (.A(_00680_));
 sg13g2_antennanp ANTENNA_21 (.A(_00680_));
 sg13g2_antennanp ANTENNA_22 (.A(_00680_));
 sg13g2_antennanp ANTENNA_23 (.A(_00680_));
 sg13g2_antennanp ANTENNA_24 (.A(_00680_));
 sg13g2_antennanp ANTENNA_25 (.A(_00683_));
 sg13g2_antennanp ANTENNA_26 (.A(_00683_));
 sg13g2_antennanp ANTENNA_27 (.A(_00683_));
 sg13g2_antennanp ANTENNA_28 (.A(_00683_));
 sg13g2_antennanp ANTENNA_29 (.A(_00683_));
 sg13g2_antennanp ANTENNA_30 (.A(_00689_));
 sg13g2_antennanp ANTENNA_31 (.A(_00689_));
 sg13g2_antennanp ANTENNA_32 (.A(_00689_));
 sg13g2_antennanp ANTENNA_33 (.A(_00689_));
 sg13g2_antennanp ANTENNA_34 (.A(_00689_));
 sg13g2_antennanp ANTENNA_35 (.A(_00790_));
 sg13g2_antennanp ANTENNA_36 (.A(_00790_));
 sg13g2_antennanp ANTENNA_37 (.A(_00790_));
 sg13g2_antennanp ANTENNA_38 (.A(_01030_));
 sg13g2_antennanp ANTENNA_39 (.A(_01030_));
 sg13g2_antennanp ANTENNA_40 (.A(_01051_));
 sg13g2_antennanp ANTENNA_41 (.A(_01053_));
 sg13g2_antennanp ANTENNA_42 (.A(_01053_));
 sg13g2_antennanp ANTENNA_43 (.A(_01056_));
 sg13g2_antennanp ANTENNA_44 (.A(_01056_));
 sg13g2_antennanp ANTENNA_45 (.A(_01061_));
 sg13g2_antennanp ANTENNA_46 (.A(_01061_));
 sg13g2_antennanp ANTENNA_47 (.A(_01061_));
 sg13g2_antennanp ANTENNA_48 (.A(_01070_));
 sg13g2_antennanp ANTENNA_49 (.A(_01070_));
 sg13g2_antennanp ANTENNA_50 (.A(_01070_));
 sg13g2_antennanp ANTENNA_51 (.A(_01071_));
 sg13g2_antennanp ANTENNA_52 (.A(_01071_));
 sg13g2_antennanp ANTENNA_53 (.A(_01071_));
 sg13g2_antennanp ANTENNA_54 (.A(_01071_));
 sg13g2_antennanp ANTENNA_55 (.A(_01071_));
 sg13g2_antennanp ANTENNA_56 (.A(_01071_));
 sg13g2_antennanp ANTENNA_57 (.A(_01151_));
 sg13g2_antennanp ANTENNA_58 (.A(_01151_));
 sg13g2_antennanp ANTENNA_59 (.A(_01151_));
 sg13g2_antennanp ANTENNA_60 (.A(_01178_));
 sg13g2_antennanp ANTENNA_61 (.A(_01178_));
 sg13g2_antennanp ANTENNA_62 (.A(_01178_));
 sg13g2_antennanp ANTENNA_63 (.A(_01178_));
 sg13g2_antennanp ANTENNA_64 (.A(_01212_));
 sg13g2_antennanp ANTENNA_65 (.A(_01212_));
 sg13g2_antennanp ANTENNA_66 (.A(_01212_));
 sg13g2_antennanp ANTENNA_67 (.A(_01252_));
 sg13g2_antennanp ANTENNA_68 (.A(_01252_));
 sg13g2_antennanp ANTENNA_69 (.A(_01252_));
 sg13g2_antennanp ANTENNA_70 (.A(_01252_));
 sg13g2_antennanp ANTENNA_71 (.A(_01360_));
 sg13g2_antennanp ANTENNA_72 (.A(_01360_));
 sg13g2_antennanp ANTENNA_73 (.A(_01360_));
 sg13g2_antennanp ANTENNA_74 (.A(_01458_));
 sg13g2_antennanp ANTENNA_75 (.A(_01458_));
 sg13g2_antennanp ANTENNA_76 (.A(_01458_));
 sg13g2_antennanp ANTENNA_77 (.A(_01458_));
 sg13g2_antennanp ANTENNA_78 (.A(_01519_));
 sg13g2_antennanp ANTENNA_79 (.A(_01519_));
 sg13g2_antennanp ANTENNA_80 (.A(_01519_));
 sg13g2_antennanp ANTENNA_81 (.A(_01527_));
 sg13g2_antennanp ANTENNA_82 (.A(_01527_));
 sg13g2_antennanp ANTENNA_83 (.A(_01527_));
 sg13g2_antennanp ANTENNA_84 (.A(_01655_));
 sg13g2_antennanp ANTENNA_85 (.A(_01655_));
 sg13g2_antennanp ANTENNA_86 (.A(_01655_));
 sg13g2_antennanp ANTENNA_87 (.A(_01655_));
 sg13g2_antennanp ANTENNA_88 (.A(_01655_));
 sg13g2_antennanp ANTENNA_89 (.A(_01655_));
 sg13g2_antennanp ANTENNA_90 (.A(_01655_));
 sg13g2_antennanp ANTENNA_91 (.A(_01655_));
 sg13g2_antennanp ANTENNA_92 (.A(_01655_));
 sg13g2_antennanp ANTENNA_93 (.A(_01675_));
 sg13g2_antennanp ANTENNA_94 (.A(_01675_));
 sg13g2_antennanp ANTENNA_95 (.A(_01675_));
 sg13g2_antennanp ANTENNA_96 (.A(_01675_));
 sg13g2_antennanp ANTENNA_97 (.A(_01675_));
 sg13g2_antennanp ANTENNA_98 (.A(_01676_));
 sg13g2_antennanp ANTENNA_99 (.A(_01676_));
 sg13g2_antennanp ANTENNA_100 (.A(_01676_));
 sg13g2_antennanp ANTENNA_101 (.A(_01726_));
 sg13g2_antennanp ANTENNA_102 (.A(_01726_));
 sg13g2_antennanp ANTENNA_103 (.A(_01844_));
 sg13g2_antennanp ANTENNA_104 (.A(_01844_));
 sg13g2_antennanp ANTENNA_105 (.A(_01844_));
 sg13g2_antennanp ANTENNA_106 (.A(_02251_));
 sg13g2_antennanp ANTENNA_107 (.A(_02251_));
 sg13g2_antennanp ANTENNA_108 (.A(_02251_));
 sg13g2_antennanp ANTENNA_109 (.A(_02395_));
 sg13g2_antennanp ANTENNA_110 (.A(_02519_));
 sg13g2_antennanp ANTENNA_111 (.A(_02567_));
 sg13g2_antennanp ANTENNA_112 (.A(_02567_));
 sg13g2_antennanp ANTENNA_113 (.A(_02567_));
 sg13g2_antennanp ANTENNA_114 (.A(_02569_));
 sg13g2_antennanp ANTENNA_115 (.A(_02569_));
 sg13g2_antennanp ANTENNA_116 (.A(_02569_));
 sg13g2_antennanp ANTENNA_117 (.A(_02569_));
 sg13g2_antennanp ANTENNA_118 (.A(_02934_));
 sg13g2_antennanp ANTENNA_119 (.A(_02934_));
 sg13g2_antennanp ANTENNA_120 (.A(_02934_));
 sg13g2_antennanp ANTENNA_121 (.A(_02942_));
 sg13g2_antennanp ANTENNA_122 (.A(_02942_));
 sg13g2_antennanp ANTENNA_123 (.A(_02959_));
 sg13g2_antennanp ANTENNA_124 (.A(_02959_));
 sg13g2_antennanp ANTENNA_125 (.A(_02959_));
 sg13g2_antennanp ANTENNA_126 (.A(_02959_));
 sg13g2_antennanp ANTENNA_127 (.A(_02959_));
 sg13g2_antennanp ANTENNA_128 (.A(_02959_));
 sg13g2_antennanp ANTENNA_129 (.A(_02959_));
 sg13g2_antennanp ANTENNA_130 (.A(_03065_));
 sg13g2_antennanp ANTENNA_131 (.A(_03065_));
 sg13g2_antennanp ANTENNA_132 (.A(_03278_));
 sg13g2_antennanp ANTENNA_133 (.A(_03304_));
 sg13g2_antennanp ANTENNA_134 (.A(_03304_));
 sg13g2_antennanp ANTENNA_135 (.A(_03354_));
 sg13g2_antennanp ANTENNA_136 (.A(_03354_));
 sg13g2_antennanp ANTENNA_137 (.A(_03354_));
 sg13g2_antennanp ANTENNA_138 (.A(_03397_));
 sg13g2_antennanp ANTENNA_139 (.A(_03397_));
 sg13g2_antennanp ANTENNA_140 (.A(_03397_));
 sg13g2_antennanp ANTENNA_141 (.A(_03535_));
 sg13g2_antennanp ANTENNA_142 (.A(_03644_));
 sg13g2_antennanp ANTENNA_143 (.A(_05221_));
 sg13g2_antennanp ANTENNA_144 (.A(_05221_));
 sg13g2_antennanp ANTENNA_145 (.A(_05221_));
 sg13g2_antennanp ANTENNA_146 (.A(_05221_));
 sg13g2_antennanp ANTENNA_147 (.A(_05221_));
 sg13g2_antennanp ANTENNA_148 (.A(_05221_));
 sg13g2_antennanp ANTENNA_149 (.A(_05300_));
 sg13g2_antennanp ANTENNA_150 (.A(_05300_));
 sg13g2_antennanp ANTENNA_151 (.A(_05424_));
 sg13g2_antennanp ANTENNA_152 (.A(_05424_));
 sg13g2_antennanp ANTENNA_153 (.A(_05424_));
 sg13g2_antennanp ANTENNA_154 (.A(_05424_));
 sg13g2_antennanp ANTENNA_155 (.A(_05424_));
 sg13g2_antennanp ANTENNA_156 (.A(_05864_));
 sg13g2_antennanp ANTENNA_157 (.A(_05864_));
 sg13g2_antennanp ANTENNA_158 (.A(_05864_));
 sg13g2_antennanp ANTENNA_159 (.A(_05864_));
 sg13g2_antennanp ANTENNA_160 (.A(_05864_));
 sg13g2_antennanp ANTENNA_161 (.A(_05864_));
 sg13g2_antennanp ANTENNA_162 (.A(_06065_));
 sg13g2_antennanp ANTENNA_163 (.A(_07183_));
 sg13g2_antennanp ANTENNA_164 (.A(_07183_));
 sg13g2_antennanp ANTENNA_165 (.A(_07183_));
 sg13g2_antennanp ANTENNA_166 (.A(_07183_));
 sg13g2_antennanp ANTENNA_167 (.A(_07183_));
 sg13g2_antennanp ANTENNA_168 (.A(_07183_));
 sg13g2_antennanp ANTENNA_169 (.A(_07183_));
 sg13g2_antennanp ANTENNA_170 (.A(_07183_));
 sg13g2_antennanp ANTENNA_171 (.A(_07184_));
 sg13g2_antennanp ANTENNA_172 (.A(_07184_));
 sg13g2_antennanp ANTENNA_173 (.A(_07184_));
 sg13g2_antennanp ANTENNA_174 (.A(_07184_));
 sg13g2_antennanp ANTENNA_175 (.A(_07190_));
 sg13g2_antennanp ANTENNA_176 (.A(_07312_));
 sg13g2_antennanp ANTENNA_177 (.A(_07334_));
 sg13g2_antennanp ANTENNA_178 (.A(_07334_));
 sg13g2_antennanp ANTENNA_179 (.A(_07335_));
 sg13g2_antennanp ANTENNA_180 (.A(_07335_));
 sg13g2_antennanp ANTENNA_181 (.A(clk));
 sg13g2_antennanp ANTENNA_182 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_183 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_184 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_185 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_186 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_187 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_188 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_189 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_190 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_191 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_192 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_193 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_194 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_195 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_196 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_197 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_198 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_199 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_200 (.A(\clock_inst.min_c[50] ));
 sg13g2_antennanp ANTENNA_201 (.A(\clock_inst.min_c[50] ));
 sg13g2_antennanp ANTENNA_202 (.A(\clock_inst.min_c[50] ));
 sg13g2_antennanp ANTENNA_203 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_204 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_205 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_206 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_207 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_208 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_209 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_210 (.A(\clock_inst.sec_c[25] ));
 sg13g2_antennanp ANTENNA_211 (.A(\clock_inst.sec_c[25] ));
 sg13g2_antennanp ANTENNA_212 (.A(\clock_inst.sec_c[25] ));
 sg13g2_antennanp ANTENNA_213 (.A(\clock_inst.sec_c[25] ));
 sg13g2_antennanp ANTENNA_214 (.A(\clock_inst.sec_c[45] ));
 sg13g2_antennanp ANTENNA_215 (.A(\clock_inst.sec_c[45] ));
 sg13g2_antennanp ANTENNA_216 (.A(\clock_inst.sec_c[45] ));
 sg13g2_antennanp ANTENNA_217 (.A(\clock_inst.sec_c[45] ));
 sg13g2_antennanp ANTENNA_218 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_219 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_220 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_221 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_222 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_223 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_224 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_225 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_226 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_227 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_228 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_229 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_230 (.A(net74));
 sg13g2_antennanp ANTENNA_231 (.A(net74));
 sg13g2_antennanp ANTENNA_232 (.A(net74));
 sg13g2_antennanp ANTENNA_233 (.A(net74));
 sg13g2_antennanp ANTENNA_234 (.A(net74));
 sg13g2_antennanp ANTENNA_235 (.A(net74));
 sg13g2_antennanp ANTENNA_236 (.A(net74));
 sg13g2_antennanp ANTENNA_237 (.A(net74));
 sg13g2_antennanp ANTENNA_238 (.A(net74));
 sg13g2_antennanp ANTENNA_239 (.A(net83));
 sg13g2_antennanp ANTENNA_240 (.A(net83));
 sg13g2_antennanp ANTENNA_241 (.A(net83));
 sg13g2_antennanp ANTENNA_242 (.A(net83));
 sg13g2_antennanp ANTENNA_243 (.A(net83));
 sg13g2_antennanp ANTENNA_244 (.A(net83));
 sg13g2_antennanp ANTENNA_245 (.A(net83));
 sg13g2_antennanp ANTENNA_246 (.A(net83));
 sg13g2_antennanp ANTENNA_247 (.A(net91));
 sg13g2_antennanp ANTENNA_248 (.A(net91));
 sg13g2_antennanp ANTENNA_249 (.A(net91));
 sg13g2_antennanp ANTENNA_250 (.A(net91));
 sg13g2_antennanp ANTENNA_251 (.A(net91));
 sg13g2_antennanp ANTENNA_252 (.A(net91));
 sg13g2_antennanp ANTENNA_253 (.A(net91));
 sg13g2_antennanp ANTENNA_254 (.A(net91));
 sg13g2_antennanp ANTENNA_255 (.A(net91));
 sg13g2_antennanp ANTENNA_256 (.A(net94));
 sg13g2_antennanp ANTENNA_257 (.A(net94));
 sg13g2_antennanp ANTENNA_258 (.A(net94));
 sg13g2_antennanp ANTENNA_259 (.A(net94));
 sg13g2_antennanp ANTENNA_260 (.A(net94));
 sg13g2_antennanp ANTENNA_261 (.A(net94));
 sg13g2_antennanp ANTENNA_262 (.A(net94));
 sg13g2_antennanp ANTENNA_263 (.A(net94));
 sg13g2_antennanp ANTENNA_264 (.A(net94));
 sg13g2_antennanp ANTENNA_265 (.A(net157));
 sg13g2_antennanp ANTENNA_266 (.A(net157));
 sg13g2_antennanp ANTENNA_267 (.A(net157));
 sg13g2_antennanp ANTENNA_268 (.A(net157));
 sg13g2_antennanp ANTENNA_269 (.A(net157));
 sg13g2_antennanp ANTENNA_270 (.A(net157));
 sg13g2_antennanp ANTENNA_271 (.A(net157));
 sg13g2_antennanp ANTENNA_272 (.A(net157));
 sg13g2_antennanp ANTENNA_273 (.A(net159));
 sg13g2_antennanp ANTENNA_274 (.A(net159));
 sg13g2_antennanp ANTENNA_275 (.A(net159));
 sg13g2_antennanp ANTENNA_276 (.A(net159));
 sg13g2_antennanp ANTENNA_277 (.A(net159));
 sg13g2_antennanp ANTENNA_278 (.A(net159));
 sg13g2_antennanp ANTENNA_279 (.A(net159));
 sg13g2_antennanp ANTENNA_280 (.A(net159));
 sg13g2_antennanp ANTENNA_281 (.A(net159));
 sg13g2_antennanp ANTENNA_282 (.A(net239));
 sg13g2_antennanp ANTENNA_283 (.A(net239));
 sg13g2_antennanp ANTENNA_284 (.A(net239));
 sg13g2_antennanp ANTENNA_285 (.A(net239));
 sg13g2_antennanp ANTENNA_286 (.A(net239));
 sg13g2_antennanp ANTENNA_287 (.A(net239));
 sg13g2_antennanp ANTENNA_288 (.A(net239));
 sg13g2_antennanp ANTENNA_289 (.A(net239));
 sg13g2_antennanp ANTENNA_290 (.A(net239));
 sg13g2_antennanp ANTENNA_291 (.A(net513));
 sg13g2_antennanp ANTENNA_292 (.A(net513));
 sg13g2_antennanp ANTENNA_293 (.A(net513));
 sg13g2_antennanp ANTENNA_294 (.A(net513));
 sg13g2_antennanp ANTENNA_295 (.A(net513));
 sg13g2_antennanp ANTENNA_296 (.A(net513));
 sg13g2_antennanp ANTENNA_297 (.A(net513));
 sg13g2_antennanp ANTENNA_298 (.A(net513));
 sg13g2_antennanp ANTENNA_299 (.A(net513));
 sg13g2_antennanp ANTENNA_300 (.A(net513));
 sg13g2_antennanp ANTENNA_301 (.A(net513));
 sg13g2_antennanp ANTENNA_302 (.A(net513));
 sg13g2_antennanp ANTENNA_303 (.A(net513));
 sg13g2_antennanp ANTENNA_304 (.A(net513));
 sg13g2_antennanp ANTENNA_305 (.A(net513));
 sg13g2_antennanp ANTENNA_306 (.A(net513));
 sg13g2_antennanp ANTENNA_307 (.A(net513));
 sg13g2_antennanp ANTENNA_308 (.A(net513));
 sg13g2_antennanp ANTENNA_309 (.A(net513));
 sg13g2_antennanp ANTENNA_310 (.A(net513));
 sg13g2_antennanp ANTENNA_311 (.A(net513));
 sg13g2_antennanp ANTENNA_312 (.A(net513));
 sg13g2_antennanp ANTENNA_313 (.A(net513));
 sg13g2_antennanp ANTENNA_314 (.A(net549));
 sg13g2_antennanp ANTENNA_315 (.A(net549));
 sg13g2_antennanp ANTENNA_316 (.A(net549));
 sg13g2_antennanp ANTENNA_317 (.A(net549));
 sg13g2_antennanp ANTENNA_318 (.A(net549));
 sg13g2_antennanp ANTENNA_319 (.A(net549));
 sg13g2_antennanp ANTENNA_320 (.A(net549));
 sg13g2_antennanp ANTENNA_321 (.A(net549));
 sg13g2_antennanp ANTENNA_322 (.A(net549));
 sg13g2_antennanp ANTENNA_323 (.A(net583));
 sg13g2_antennanp ANTENNA_324 (.A(net583));
 sg13g2_antennanp ANTENNA_325 (.A(net583));
 sg13g2_antennanp ANTENNA_326 (.A(net583));
 sg13g2_antennanp ANTENNA_327 (.A(net583));
 sg13g2_antennanp ANTENNA_328 (.A(net583));
 sg13g2_antennanp ANTENNA_329 (.A(net583));
 sg13g2_antennanp ANTENNA_330 (.A(net583));
 sg13g2_antennanp ANTENNA_331 (.A(net583));
 sg13g2_antennanp ANTENNA_332 (.A(net583));
 sg13g2_antennanp ANTENNA_333 (.A(net583));
 sg13g2_antennanp ANTENNA_334 (.A(net583));
 sg13g2_antennanp ANTENNA_335 (.A(net583));
 sg13g2_antennanp ANTENNA_336 (.A(net583));
 sg13g2_antennanp ANTENNA_337 (.A(net583));
 sg13g2_antennanp ANTENNA_338 (.A(net583));
 sg13g2_antennanp ANTENNA_339 (.A(net583));
 sg13g2_antennanp ANTENNA_340 (.A(net583));
 sg13g2_antennanp ANTENNA_341 (.A(net583));
 sg13g2_antennanp ANTENNA_342 (.A(net583));
 sg13g2_antennanp ANTENNA_343 (.A(net583));
 sg13g2_antennanp ANTENNA_344 (.A(_00216_));
 sg13g2_antennanp ANTENNA_345 (.A(_00216_));
 sg13g2_antennanp ANTENNA_346 (.A(_00242_));
 sg13g2_antennanp ANTENNA_347 (.A(_00242_));
 sg13g2_antennanp ANTENNA_348 (.A(_00419_));
 sg13g2_antennanp ANTENNA_349 (.A(_00419_));
 sg13g2_antennanp ANTENNA_350 (.A(_00656_));
 sg13g2_antennanp ANTENNA_351 (.A(_00656_));
 sg13g2_antennanp ANTENNA_352 (.A(_00656_));
 sg13g2_antennanp ANTENNA_353 (.A(_00656_));
 sg13g2_antennanp ANTENNA_354 (.A(_00656_));
 sg13g2_antennanp ANTENNA_355 (.A(_00680_));
 sg13g2_antennanp ANTENNA_356 (.A(_00680_));
 sg13g2_antennanp ANTENNA_357 (.A(_00680_));
 sg13g2_antennanp ANTENNA_358 (.A(_00680_));
 sg13g2_antennanp ANTENNA_359 (.A(_00680_));
 sg13g2_antennanp ANTENNA_360 (.A(_00680_));
 sg13g2_antennanp ANTENNA_361 (.A(_00683_));
 sg13g2_antennanp ANTENNA_362 (.A(_00683_));
 sg13g2_antennanp ANTENNA_363 (.A(_00683_));
 sg13g2_antennanp ANTENNA_364 (.A(_00683_));
 sg13g2_antennanp ANTENNA_365 (.A(_00683_));
 sg13g2_antennanp ANTENNA_366 (.A(_00790_));
 sg13g2_antennanp ANTENNA_367 (.A(_00790_));
 sg13g2_antennanp ANTENNA_368 (.A(_00790_));
 sg13g2_antennanp ANTENNA_369 (.A(_00790_));
 sg13g2_antennanp ANTENNA_370 (.A(_00790_));
 sg13g2_antennanp ANTENNA_371 (.A(_00790_));
 sg13g2_antennanp ANTENNA_372 (.A(_00790_));
 sg13g2_antennanp ANTENNA_373 (.A(_01030_));
 sg13g2_antennanp ANTENNA_374 (.A(_01030_));
 sg13g2_antennanp ANTENNA_375 (.A(_01051_));
 sg13g2_antennanp ANTENNA_376 (.A(_01056_));
 sg13g2_antennanp ANTENNA_377 (.A(_01056_));
 sg13g2_antennanp ANTENNA_378 (.A(_01070_));
 sg13g2_antennanp ANTENNA_379 (.A(_01070_));
 sg13g2_antennanp ANTENNA_380 (.A(_01070_));
 sg13g2_antennanp ANTENNA_381 (.A(_01071_));
 sg13g2_antennanp ANTENNA_382 (.A(_01071_));
 sg13g2_antennanp ANTENNA_383 (.A(_01071_));
 sg13g2_antennanp ANTENNA_384 (.A(_01071_));
 sg13g2_antennanp ANTENNA_385 (.A(_01178_));
 sg13g2_antennanp ANTENNA_386 (.A(_01178_));
 sg13g2_antennanp ANTENNA_387 (.A(_01178_));
 sg13g2_antennanp ANTENNA_388 (.A(_01178_));
 sg13g2_antennanp ANTENNA_389 (.A(_01212_));
 sg13g2_antennanp ANTENNA_390 (.A(_01212_));
 sg13g2_antennanp ANTENNA_391 (.A(_01212_));
 sg13g2_antennanp ANTENNA_392 (.A(_01252_));
 sg13g2_antennanp ANTENNA_393 (.A(_01252_));
 sg13g2_antennanp ANTENNA_394 (.A(_01252_));
 sg13g2_antennanp ANTENNA_395 (.A(_01252_));
 sg13g2_antennanp ANTENNA_396 (.A(_01360_));
 sg13g2_antennanp ANTENNA_397 (.A(_01360_));
 sg13g2_antennanp ANTENNA_398 (.A(_01360_));
 sg13g2_antennanp ANTENNA_399 (.A(_01675_));
 sg13g2_antennanp ANTENNA_400 (.A(_01675_));
 sg13g2_antennanp ANTENNA_401 (.A(_01675_));
 sg13g2_antennanp ANTENNA_402 (.A(_01675_));
 sg13g2_antennanp ANTENNA_403 (.A(_01675_));
 sg13g2_antennanp ANTENNA_404 (.A(_01676_));
 sg13g2_antennanp ANTENNA_405 (.A(_01676_));
 sg13g2_antennanp ANTENNA_406 (.A(_01676_));
 sg13g2_antennanp ANTENNA_407 (.A(_01676_));
 sg13g2_antennanp ANTENNA_408 (.A(_01726_));
 sg13g2_antennanp ANTENNA_409 (.A(_01844_));
 sg13g2_antennanp ANTENNA_410 (.A(_01844_));
 sg13g2_antennanp ANTENNA_411 (.A(_01844_));
 sg13g2_antennanp ANTENNA_412 (.A(_02395_));
 sg13g2_antennanp ANTENNA_413 (.A(_02519_));
 sg13g2_antennanp ANTENNA_414 (.A(_02567_));
 sg13g2_antennanp ANTENNA_415 (.A(_02567_));
 sg13g2_antennanp ANTENNA_416 (.A(_02567_));
 sg13g2_antennanp ANTENNA_417 (.A(_02934_));
 sg13g2_antennanp ANTENNA_418 (.A(_02942_));
 sg13g2_antennanp ANTENNA_419 (.A(_02942_));
 sg13g2_antennanp ANTENNA_420 (.A(_03065_));
 sg13g2_antennanp ANTENNA_421 (.A(_03065_));
 sg13g2_antennanp ANTENNA_422 (.A(_03278_));
 sg13g2_antennanp ANTENNA_423 (.A(_03304_));
 sg13g2_antennanp ANTENNA_424 (.A(_03304_));
 sg13g2_antennanp ANTENNA_425 (.A(_03354_));
 sg13g2_antennanp ANTENNA_426 (.A(_03354_));
 sg13g2_antennanp ANTENNA_427 (.A(_03354_));
 sg13g2_antennanp ANTENNA_428 (.A(_03397_));
 sg13g2_antennanp ANTENNA_429 (.A(_03397_));
 sg13g2_antennanp ANTENNA_430 (.A(_03397_));
 sg13g2_antennanp ANTENNA_431 (.A(_03535_));
 sg13g2_antennanp ANTENNA_432 (.A(_03644_));
 sg13g2_antennanp ANTENNA_433 (.A(_05221_));
 sg13g2_antennanp ANTENNA_434 (.A(_05221_));
 sg13g2_antennanp ANTENNA_435 (.A(_05221_));
 sg13g2_antennanp ANTENNA_436 (.A(_05221_));
 sg13g2_antennanp ANTENNA_437 (.A(_05221_));
 sg13g2_antennanp ANTENNA_438 (.A(_05221_));
 sg13g2_antennanp ANTENNA_439 (.A(_05300_));
 sg13g2_antennanp ANTENNA_440 (.A(_05300_));
 sg13g2_antennanp ANTENNA_441 (.A(_05424_));
 sg13g2_antennanp ANTENNA_442 (.A(_05424_));
 sg13g2_antennanp ANTENNA_443 (.A(_05424_));
 sg13g2_antennanp ANTENNA_444 (.A(_05424_));
 sg13g2_antennanp ANTENNA_445 (.A(_05424_));
 sg13g2_antennanp ANTENNA_446 (.A(_05864_));
 sg13g2_antennanp ANTENNA_447 (.A(_05864_));
 sg13g2_antennanp ANTENNA_448 (.A(_05864_));
 sg13g2_antennanp ANTENNA_449 (.A(_05864_));
 sg13g2_antennanp ANTENNA_450 (.A(_05864_));
 sg13g2_antennanp ANTENNA_451 (.A(_05864_));
 sg13g2_antennanp ANTENNA_452 (.A(_06065_));
 sg13g2_antennanp ANTENNA_453 (.A(_07183_));
 sg13g2_antennanp ANTENNA_454 (.A(_07183_));
 sg13g2_antennanp ANTENNA_455 (.A(_07183_));
 sg13g2_antennanp ANTENNA_456 (.A(_07183_));
 sg13g2_antennanp ANTENNA_457 (.A(_07183_));
 sg13g2_antennanp ANTENNA_458 (.A(_07183_));
 sg13g2_antennanp ANTENNA_459 (.A(_07183_));
 sg13g2_antennanp ANTENNA_460 (.A(_07183_));
 sg13g2_antennanp ANTENNA_461 (.A(_07183_));
 sg13g2_antennanp ANTENNA_462 (.A(_07183_));
 sg13g2_antennanp ANTENNA_463 (.A(_07184_));
 sg13g2_antennanp ANTENNA_464 (.A(_07184_));
 sg13g2_antennanp ANTENNA_465 (.A(_07184_));
 sg13g2_antennanp ANTENNA_466 (.A(_07184_));
 sg13g2_antennanp ANTENNA_467 (.A(_07190_));
 sg13g2_antennanp ANTENNA_468 (.A(_07190_));
 sg13g2_antennanp ANTENNA_469 (.A(_07312_));
 sg13g2_antennanp ANTENNA_470 (.A(_07334_));
 sg13g2_antennanp ANTENNA_471 (.A(_07334_));
 sg13g2_antennanp ANTENNA_472 (.A(_07335_));
 sg13g2_antennanp ANTENNA_473 (.A(_07335_));
 sg13g2_antennanp ANTENNA_474 (.A(clk));
 sg13g2_antennanp ANTENNA_475 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_476 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_477 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_478 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_479 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_480 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_481 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_482 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_483 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_484 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_485 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_486 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_487 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_488 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_489 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_490 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_491 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_492 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_493 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_494 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_495 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_496 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_497 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_498 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_499 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_500 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_501 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_502 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_503 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_504 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_505 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_506 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_507 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_508 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_509 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_510 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_511 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_512 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_513 (.A(net74));
 sg13g2_antennanp ANTENNA_514 (.A(net74));
 sg13g2_antennanp ANTENNA_515 (.A(net74));
 sg13g2_antennanp ANTENNA_516 (.A(net74));
 sg13g2_antennanp ANTENNA_517 (.A(net74));
 sg13g2_antennanp ANTENNA_518 (.A(net74));
 sg13g2_antennanp ANTENNA_519 (.A(net74));
 sg13g2_antennanp ANTENNA_520 (.A(net74));
 sg13g2_antennanp ANTENNA_521 (.A(net74));
 sg13g2_antennanp ANTENNA_522 (.A(net83));
 sg13g2_antennanp ANTENNA_523 (.A(net83));
 sg13g2_antennanp ANTENNA_524 (.A(net83));
 sg13g2_antennanp ANTENNA_525 (.A(net83));
 sg13g2_antennanp ANTENNA_526 (.A(net83));
 sg13g2_antennanp ANTENNA_527 (.A(net83));
 sg13g2_antennanp ANTENNA_528 (.A(net83));
 sg13g2_antennanp ANTENNA_529 (.A(net83));
 sg13g2_antennanp ANTENNA_530 (.A(net83));
 sg13g2_antennanp ANTENNA_531 (.A(net83));
 sg13g2_antennanp ANTENNA_532 (.A(net83));
 sg13g2_antennanp ANTENNA_533 (.A(net83));
 sg13g2_antennanp ANTENNA_534 (.A(net83));
 sg13g2_antennanp ANTENNA_535 (.A(net83));
 sg13g2_antennanp ANTENNA_536 (.A(net83));
 sg13g2_antennanp ANTENNA_537 (.A(net83));
 sg13g2_antennanp ANTENNA_538 (.A(net83));
 sg13g2_antennanp ANTENNA_539 (.A(net83));
 sg13g2_antennanp ANTENNA_540 (.A(net157));
 sg13g2_antennanp ANTENNA_541 (.A(net157));
 sg13g2_antennanp ANTENNA_542 (.A(net157));
 sg13g2_antennanp ANTENNA_543 (.A(net157));
 sg13g2_antennanp ANTENNA_544 (.A(net157));
 sg13g2_antennanp ANTENNA_545 (.A(net157));
 sg13g2_antennanp ANTENNA_546 (.A(net157));
 sg13g2_antennanp ANTENNA_547 (.A(net157));
 sg13g2_antennanp ANTENNA_548 (.A(net159));
 sg13g2_antennanp ANTENNA_549 (.A(net159));
 sg13g2_antennanp ANTENNA_550 (.A(net159));
 sg13g2_antennanp ANTENNA_551 (.A(net159));
 sg13g2_antennanp ANTENNA_552 (.A(net159));
 sg13g2_antennanp ANTENNA_553 (.A(net159));
 sg13g2_antennanp ANTENNA_554 (.A(net159));
 sg13g2_antennanp ANTENNA_555 (.A(net159));
 sg13g2_antennanp ANTENNA_556 (.A(net159));
 sg13g2_antennanp ANTENNA_557 (.A(net239));
 sg13g2_antennanp ANTENNA_558 (.A(net239));
 sg13g2_antennanp ANTENNA_559 (.A(net239));
 sg13g2_antennanp ANTENNA_560 (.A(net239));
 sg13g2_antennanp ANTENNA_561 (.A(net239));
 sg13g2_antennanp ANTENNA_562 (.A(net239));
 sg13g2_antennanp ANTENNA_563 (.A(net239));
 sg13g2_antennanp ANTENNA_564 (.A(net239));
 sg13g2_antennanp ANTENNA_565 (.A(net239));
 sg13g2_antennanp ANTENNA_566 (.A(net513));
 sg13g2_antennanp ANTENNA_567 (.A(net513));
 sg13g2_antennanp ANTENNA_568 (.A(net513));
 sg13g2_antennanp ANTENNA_569 (.A(net513));
 sg13g2_antennanp ANTENNA_570 (.A(net513));
 sg13g2_antennanp ANTENNA_571 (.A(net513));
 sg13g2_antennanp ANTENNA_572 (.A(net513));
 sg13g2_antennanp ANTENNA_573 (.A(net513));
 sg13g2_antennanp ANTENNA_574 (.A(net513));
 sg13g2_antennanp ANTENNA_575 (.A(net549));
 sg13g2_antennanp ANTENNA_576 (.A(net549));
 sg13g2_antennanp ANTENNA_577 (.A(net549));
 sg13g2_antennanp ANTENNA_578 (.A(net549));
 sg13g2_antennanp ANTENNA_579 (.A(net549));
 sg13g2_antennanp ANTENNA_580 (.A(net549));
 sg13g2_antennanp ANTENNA_581 (.A(net549));
 sg13g2_antennanp ANTENNA_582 (.A(net549));
 sg13g2_antennanp ANTENNA_583 (.A(net549));
 sg13g2_antennanp ANTENNA_584 (.A(net583));
 sg13g2_antennanp ANTENNA_585 (.A(net583));
 sg13g2_antennanp ANTENNA_586 (.A(net583));
 sg13g2_antennanp ANTENNA_587 (.A(net583));
 sg13g2_antennanp ANTENNA_588 (.A(net583));
 sg13g2_antennanp ANTENNA_589 (.A(net583));
 sg13g2_antennanp ANTENNA_590 (.A(net583));
 sg13g2_antennanp ANTENNA_591 (.A(net583));
 sg13g2_antennanp ANTENNA_592 (.A(net583));
 sg13g2_antennanp ANTENNA_593 (.A(net583));
 sg13g2_antennanp ANTENNA_594 (.A(net583));
 sg13g2_antennanp ANTENNA_595 (.A(net583));
 sg13g2_antennanp ANTENNA_596 (.A(net583));
 sg13g2_antennanp ANTENNA_597 (.A(net583));
 sg13g2_antennanp ANTENNA_598 (.A(net583));
 sg13g2_antennanp ANTENNA_599 (.A(net583));
 sg13g2_antennanp ANTENNA_600 (.A(net583));
 sg13g2_antennanp ANTENNA_601 (.A(net583));
 sg13g2_antennanp ANTENNA_602 (.A(net583));
 sg13g2_antennanp ANTENNA_603 (.A(net583));
 sg13g2_antennanp ANTENNA_604 (.A(net583));
 sg13g2_antennanp ANTENNA_605 (.A(_00216_));
 sg13g2_antennanp ANTENNA_606 (.A(_00216_));
 sg13g2_antennanp ANTENNA_607 (.A(_00242_));
 sg13g2_antennanp ANTENNA_608 (.A(_00242_));
 sg13g2_antennanp ANTENNA_609 (.A(_00419_));
 sg13g2_antennanp ANTENNA_610 (.A(_00419_));
 sg13g2_antennanp ANTENNA_611 (.A(_00656_));
 sg13g2_antennanp ANTENNA_612 (.A(_00656_));
 sg13g2_antennanp ANTENNA_613 (.A(_00656_));
 sg13g2_antennanp ANTENNA_614 (.A(_00680_));
 sg13g2_antennanp ANTENNA_615 (.A(_00680_));
 sg13g2_antennanp ANTENNA_616 (.A(_00680_));
 sg13g2_antennanp ANTENNA_617 (.A(_00680_));
 sg13g2_antennanp ANTENNA_618 (.A(_00683_));
 sg13g2_antennanp ANTENNA_619 (.A(_00683_));
 sg13g2_antennanp ANTENNA_620 (.A(_00683_));
 sg13g2_antennanp ANTENNA_621 (.A(_01051_));
 sg13g2_antennanp ANTENNA_622 (.A(_01056_));
 sg13g2_antennanp ANTENNA_623 (.A(_01056_));
 sg13g2_antennanp ANTENNA_624 (.A(_01070_));
 sg13g2_antennanp ANTENNA_625 (.A(_01070_));
 sg13g2_antennanp ANTENNA_626 (.A(_01071_));
 sg13g2_antennanp ANTENNA_627 (.A(_01071_));
 sg13g2_antennanp ANTENNA_628 (.A(_01071_));
 sg13g2_antennanp ANTENNA_629 (.A(_01071_));
 sg13g2_antennanp ANTENNA_630 (.A(_01178_));
 sg13g2_antennanp ANTENNA_631 (.A(_01178_));
 sg13g2_antennanp ANTENNA_632 (.A(_01178_));
 sg13g2_antennanp ANTENNA_633 (.A(_01178_));
 sg13g2_antennanp ANTENNA_634 (.A(_01212_));
 sg13g2_antennanp ANTENNA_635 (.A(_01212_));
 sg13g2_antennanp ANTENNA_636 (.A(_01212_));
 sg13g2_antennanp ANTENNA_637 (.A(_01252_));
 sg13g2_antennanp ANTENNA_638 (.A(_01252_));
 sg13g2_antennanp ANTENNA_639 (.A(_01252_));
 sg13g2_antennanp ANTENNA_640 (.A(_01252_));
 sg13g2_antennanp ANTENNA_641 (.A(_01360_));
 sg13g2_antennanp ANTENNA_642 (.A(_01360_));
 sg13g2_antennanp ANTENNA_643 (.A(_01360_));
 sg13g2_antennanp ANTENNA_644 (.A(_01675_));
 sg13g2_antennanp ANTENNA_645 (.A(_01675_));
 sg13g2_antennanp ANTENNA_646 (.A(_01675_));
 sg13g2_antennanp ANTENNA_647 (.A(_01675_));
 sg13g2_antennanp ANTENNA_648 (.A(_01675_));
 sg13g2_antennanp ANTENNA_649 (.A(_01676_));
 sg13g2_antennanp ANTENNA_650 (.A(_01676_));
 sg13g2_antennanp ANTENNA_651 (.A(_01676_));
 sg13g2_antennanp ANTENNA_652 (.A(_01676_));
 sg13g2_antennanp ANTENNA_653 (.A(_01726_));
 sg13g2_antennanp ANTENNA_654 (.A(_01844_));
 sg13g2_antennanp ANTENNA_655 (.A(_01844_));
 sg13g2_antennanp ANTENNA_656 (.A(_01844_));
 sg13g2_antennanp ANTENNA_657 (.A(_02395_));
 sg13g2_antennanp ANTENNA_658 (.A(_02519_));
 sg13g2_antennanp ANTENNA_659 (.A(_02567_));
 sg13g2_antennanp ANTENNA_660 (.A(_02567_));
 sg13g2_antennanp ANTENNA_661 (.A(_02567_));
 sg13g2_antennanp ANTENNA_662 (.A(_02934_));
 sg13g2_antennanp ANTENNA_663 (.A(_02942_));
 sg13g2_antennanp ANTENNA_664 (.A(_02942_));
 sg13g2_antennanp ANTENNA_665 (.A(_03065_));
 sg13g2_antennanp ANTENNA_666 (.A(_03065_));
 sg13g2_antennanp ANTENNA_667 (.A(_03278_));
 sg13g2_antennanp ANTENNA_668 (.A(_03304_));
 sg13g2_antennanp ANTENNA_669 (.A(_03304_));
 sg13g2_antennanp ANTENNA_670 (.A(_03354_));
 sg13g2_antennanp ANTENNA_671 (.A(_03354_));
 sg13g2_antennanp ANTENNA_672 (.A(_03354_));
 sg13g2_antennanp ANTENNA_673 (.A(_03397_));
 sg13g2_antennanp ANTENNA_674 (.A(_03397_));
 sg13g2_antennanp ANTENNA_675 (.A(_03397_));
 sg13g2_antennanp ANTENNA_676 (.A(_03535_));
 sg13g2_antennanp ANTENNA_677 (.A(_03644_));
 sg13g2_antennanp ANTENNA_678 (.A(_05221_));
 sg13g2_antennanp ANTENNA_679 (.A(_05221_));
 sg13g2_antennanp ANTENNA_680 (.A(_05221_));
 sg13g2_antennanp ANTENNA_681 (.A(_05221_));
 sg13g2_antennanp ANTENNA_682 (.A(_05221_));
 sg13g2_antennanp ANTENNA_683 (.A(_05221_));
 sg13g2_antennanp ANTENNA_684 (.A(_05300_));
 sg13g2_antennanp ANTENNA_685 (.A(_05300_));
 sg13g2_antennanp ANTENNA_686 (.A(_05424_));
 sg13g2_antennanp ANTENNA_687 (.A(_05424_));
 sg13g2_antennanp ANTENNA_688 (.A(_05424_));
 sg13g2_antennanp ANTENNA_689 (.A(_05424_));
 sg13g2_antennanp ANTENNA_690 (.A(_05424_));
 sg13g2_antennanp ANTENNA_691 (.A(_05864_));
 sg13g2_antennanp ANTENNA_692 (.A(_05864_));
 sg13g2_antennanp ANTENNA_693 (.A(_05864_));
 sg13g2_antennanp ANTENNA_694 (.A(_05864_));
 sg13g2_antennanp ANTENNA_695 (.A(_05864_));
 sg13g2_antennanp ANTENNA_696 (.A(_05864_));
 sg13g2_antennanp ANTENNA_697 (.A(_06065_));
 sg13g2_antennanp ANTENNA_698 (.A(_07183_));
 sg13g2_antennanp ANTENNA_699 (.A(_07183_));
 sg13g2_antennanp ANTENNA_700 (.A(_07183_));
 sg13g2_antennanp ANTENNA_701 (.A(_07183_));
 sg13g2_antennanp ANTENNA_702 (.A(_07183_));
 sg13g2_antennanp ANTENNA_703 (.A(_07183_));
 sg13g2_antennanp ANTENNA_704 (.A(_07183_));
 sg13g2_antennanp ANTENNA_705 (.A(_07183_));
 sg13g2_antennanp ANTENNA_706 (.A(_07183_));
 sg13g2_antennanp ANTENNA_707 (.A(_07183_));
 sg13g2_antennanp ANTENNA_708 (.A(_07190_));
 sg13g2_antennanp ANTENNA_709 (.A(_07312_));
 sg13g2_antennanp ANTENNA_710 (.A(_07334_));
 sg13g2_antennanp ANTENNA_711 (.A(_07334_));
 sg13g2_antennanp ANTENNA_712 (.A(_07335_));
 sg13g2_antennanp ANTENNA_713 (.A(_07335_));
 sg13g2_antennanp ANTENNA_714 (.A(clk));
 sg13g2_antennanp ANTENNA_715 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_716 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_717 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_718 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_719 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_720 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_721 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_722 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_723 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_724 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_725 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_726 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_727 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_728 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_729 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_730 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_731 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_732 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_733 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_734 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_735 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_736 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_737 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_738 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_739 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_740 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_741 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_742 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_743 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_744 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_745 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_746 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_747 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_748 (.A(\clock_inst.sec_c[49] ));
 sg13g2_antennanp ANTENNA_749 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_750 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_751 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_752 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_753 (.A(net74));
 sg13g2_antennanp ANTENNA_754 (.A(net74));
 sg13g2_antennanp ANTENNA_755 (.A(net74));
 sg13g2_antennanp ANTENNA_756 (.A(net74));
 sg13g2_antennanp ANTENNA_757 (.A(net74));
 sg13g2_antennanp ANTENNA_758 (.A(net74));
 sg13g2_antennanp ANTENNA_759 (.A(net74));
 sg13g2_antennanp ANTENNA_760 (.A(net74));
 sg13g2_antennanp ANTENNA_761 (.A(net74));
 sg13g2_antennanp ANTENNA_762 (.A(net83));
 sg13g2_antennanp ANTENNA_763 (.A(net83));
 sg13g2_antennanp ANTENNA_764 (.A(net83));
 sg13g2_antennanp ANTENNA_765 (.A(net83));
 sg13g2_antennanp ANTENNA_766 (.A(net83));
 sg13g2_antennanp ANTENNA_767 (.A(net83));
 sg13g2_antennanp ANTENNA_768 (.A(net83));
 sg13g2_antennanp ANTENNA_769 (.A(net83));
 sg13g2_antennanp ANTENNA_770 (.A(net83));
 sg13g2_antennanp ANTENNA_771 (.A(net83));
 sg13g2_antennanp ANTENNA_772 (.A(net83));
 sg13g2_antennanp ANTENNA_773 (.A(net83));
 sg13g2_antennanp ANTENNA_774 (.A(net83));
 sg13g2_antennanp ANTENNA_775 (.A(net83));
 sg13g2_antennanp ANTENNA_776 (.A(net83));
 sg13g2_antennanp ANTENNA_777 (.A(net83));
 sg13g2_antennanp ANTENNA_778 (.A(net83));
 sg13g2_antennanp ANTENNA_779 (.A(net83));
 sg13g2_antennanp ANTENNA_780 (.A(net157));
 sg13g2_antennanp ANTENNA_781 (.A(net157));
 sg13g2_antennanp ANTENNA_782 (.A(net157));
 sg13g2_antennanp ANTENNA_783 (.A(net157));
 sg13g2_antennanp ANTENNA_784 (.A(net157));
 sg13g2_antennanp ANTENNA_785 (.A(net157));
 sg13g2_antennanp ANTENNA_786 (.A(net157));
 sg13g2_antennanp ANTENNA_787 (.A(net157));
 sg13g2_antennanp ANTENNA_788 (.A(net159));
 sg13g2_antennanp ANTENNA_789 (.A(net159));
 sg13g2_antennanp ANTENNA_790 (.A(net159));
 sg13g2_antennanp ANTENNA_791 (.A(net159));
 sg13g2_antennanp ANTENNA_792 (.A(net159));
 sg13g2_antennanp ANTENNA_793 (.A(net159));
 sg13g2_antennanp ANTENNA_794 (.A(net159));
 sg13g2_antennanp ANTENNA_795 (.A(net159));
 sg13g2_antennanp ANTENNA_796 (.A(net159));
 sg13g2_antennanp ANTENNA_797 (.A(net239));
 sg13g2_antennanp ANTENNA_798 (.A(net239));
 sg13g2_antennanp ANTENNA_799 (.A(net239));
 sg13g2_antennanp ANTENNA_800 (.A(net239));
 sg13g2_antennanp ANTENNA_801 (.A(net239));
 sg13g2_antennanp ANTENNA_802 (.A(net239));
 sg13g2_antennanp ANTENNA_803 (.A(net239));
 sg13g2_antennanp ANTENNA_804 (.A(net239));
 sg13g2_antennanp ANTENNA_805 (.A(net239));
 sg13g2_antennanp ANTENNA_806 (.A(net513));
 sg13g2_antennanp ANTENNA_807 (.A(net513));
 sg13g2_antennanp ANTENNA_808 (.A(net513));
 sg13g2_antennanp ANTENNA_809 (.A(net513));
 sg13g2_antennanp ANTENNA_810 (.A(net513));
 sg13g2_antennanp ANTENNA_811 (.A(net513));
 sg13g2_antennanp ANTENNA_812 (.A(net513));
 sg13g2_antennanp ANTENNA_813 (.A(net513));
 sg13g2_antennanp ANTENNA_814 (.A(net513));
 sg13g2_antennanp ANTENNA_815 (.A(net549));
 sg13g2_antennanp ANTENNA_816 (.A(net549));
 sg13g2_antennanp ANTENNA_817 (.A(net549));
 sg13g2_antennanp ANTENNA_818 (.A(net549));
 sg13g2_antennanp ANTENNA_819 (.A(net549));
 sg13g2_antennanp ANTENNA_820 (.A(net549));
 sg13g2_antennanp ANTENNA_821 (.A(net549));
 sg13g2_antennanp ANTENNA_822 (.A(net549));
 sg13g2_antennanp ANTENNA_823 (.A(net549));
 sg13g2_antennanp ANTENNA_824 (.A(net583));
 sg13g2_antennanp ANTENNA_825 (.A(net583));
 sg13g2_antennanp ANTENNA_826 (.A(net583));
 sg13g2_antennanp ANTENNA_827 (.A(net583));
 sg13g2_antennanp ANTENNA_828 (.A(net583));
 sg13g2_antennanp ANTENNA_829 (.A(net583));
 sg13g2_antennanp ANTENNA_830 (.A(net583));
 sg13g2_antennanp ANTENNA_831 (.A(net583));
 sg13g2_antennanp ANTENNA_832 (.A(net583));
 sg13g2_antennanp ANTENNA_833 (.A(net583));
 sg13g2_antennanp ANTENNA_834 (.A(net583));
 sg13g2_antennanp ANTENNA_835 (.A(net583));
 sg13g2_antennanp ANTENNA_836 (.A(net583));
 sg13g2_antennanp ANTENNA_837 (.A(net583));
 sg13g2_antennanp ANTENNA_838 (.A(net583));
 sg13g2_antennanp ANTENNA_839 (.A(net583));
 sg13g2_antennanp ANTENNA_840 (.A(net583));
 sg13g2_antennanp ANTENNA_841 (.A(net583));
 sg13g2_antennanp ANTENNA_842 (.A(net583));
 sg13g2_antennanp ANTENNA_843 (.A(net583));
 sg13g2_antennanp ANTENNA_844 (.A(net583));
 sg13g2_antennanp ANTENNA_845 (.A(_00216_));
 sg13g2_antennanp ANTENNA_846 (.A(_00216_));
 sg13g2_antennanp ANTENNA_847 (.A(_00242_));
 sg13g2_antennanp ANTENNA_848 (.A(_00242_));
 sg13g2_antennanp ANTENNA_849 (.A(_00419_));
 sg13g2_antennanp ANTENNA_850 (.A(_00419_));
 sg13g2_antennanp ANTENNA_851 (.A(_00656_));
 sg13g2_antennanp ANTENNA_852 (.A(_00656_));
 sg13g2_antennanp ANTENNA_853 (.A(_00656_));
 sg13g2_antennanp ANTENNA_854 (.A(_00680_));
 sg13g2_antennanp ANTENNA_855 (.A(_00680_));
 sg13g2_antennanp ANTENNA_856 (.A(_00680_));
 sg13g2_antennanp ANTENNA_857 (.A(_00680_));
 sg13g2_antennanp ANTENNA_858 (.A(_00680_));
 sg13g2_antennanp ANTENNA_859 (.A(_00680_));
 sg13g2_antennanp ANTENNA_860 (.A(_00680_));
 sg13g2_antennanp ANTENNA_861 (.A(_00680_));
 sg13g2_antennanp ANTENNA_862 (.A(_00680_));
 sg13g2_antennanp ANTENNA_863 (.A(_00683_));
 sg13g2_antennanp ANTENNA_864 (.A(_00683_));
 sg13g2_antennanp ANTENNA_865 (.A(_00683_));
 sg13g2_antennanp ANTENNA_866 (.A(_01051_));
 sg13g2_antennanp ANTENNA_867 (.A(_01056_));
 sg13g2_antennanp ANTENNA_868 (.A(_01056_));
 sg13g2_antennanp ANTENNA_869 (.A(_01070_));
 sg13g2_antennanp ANTENNA_870 (.A(_01070_));
 sg13g2_antennanp ANTENNA_871 (.A(_01071_));
 sg13g2_antennanp ANTENNA_872 (.A(_01071_));
 sg13g2_antennanp ANTENNA_873 (.A(_01071_));
 sg13g2_antennanp ANTENNA_874 (.A(_01071_));
 sg13g2_antennanp ANTENNA_875 (.A(_01178_));
 sg13g2_antennanp ANTENNA_876 (.A(_01178_));
 sg13g2_antennanp ANTENNA_877 (.A(_01178_));
 sg13g2_antennanp ANTENNA_878 (.A(_01178_));
 sg13g2_antennanp ANTENNA_879 (.A(_01212_));
 sg13g2_antennanp ANTENNA_880 (.A(_01212_));
 sg13g2_antennanp ANTENNA_881 (.A(_01212_));
 sg13g2_antennanp ANTENNA_882 (.A(_01252_));
 sg13g2_antennanp ANTENNA_883 (.A(_01252_));
 sg13g2_antennanp ANTENNA_884 (.A(_01252_));
 sg13g2_antennanp ANTENNA_885 (.A(_01252_));
 sg13g2_antennanp ANTENNA_886 (.A(_01360_));
 sg13g2_antennanp ANTENNA_887 (.A(_01360_));
 sg13g2_antennanp ANTENNA_888 (.A(_01360_));
 sg13g2_antennanp ANTENNA_889 (.A(_01675_));
 sg13g2_antennanp ANTENNA_890 (.A(_01675_));
 sg13g2_antennanp ANTENNA_891 (.A(_01675_));
 sg13g2_antennanp ANTENNA_892 (.A(_01675_));
 sg13g2_antennanp ANTENNA_893 (.A(_01675_));
 sg13g2_antennanp ANTENNA_894 (.A(_01676_));
 sg13g2_antennanp ANTENNA_895 (.A(_01676_));
 sg13g2_antennanp ANTENNA_896 (.A(_01676_));
 sg13g2_antennanp ANTENNA_897 (.A(_01676_));
 sg13g2_antennanp ANTENNA_898 (.A(_01726_));
 sg13g2_antennanp ANTENNA_899 (.A(_01726_));
 sg13g2_antennanp ANTENNA_900 (.A(_01844_));
 sg13g2_antennanp ANTENNA_901 (.A(_01844_));
 sg13g2_antennanp ANTENNA_902 (.A(_01844_));
 sg13g2_antennanp ANTENNA_903 (.A(_02395_));
 sg13g2_antennanp ANTENNA_904 (.A(_02519_));
 sg13g2_antennanp ANTENNA_905 (.A(_02567_));
 sg13g2_antennanp ANTENNA_906 (.A(_02567_));
 sg13g2_antennanp ANTENNA_907 (.A(_02567_));
 sg13g2_antennanp ANTENNA_908 (.A(_02934_));
 sg13g2_antennanp ANTENNA_909 (.A(_02942_));
 sg13g2_antennanp ANTENNA_910 (.A(_02942_));
 sg13g2_antennanp ANTENNA_911 (.A(_03065_));
 sg13g2_antennanp ANTENNA_912 (.A(_03065_));
 sg13g2_antennanp ANTENNA_913 (.A(_03278_));
 sg13g2_antennanp ANTENNA_914 (.A(_03304_));
 sg13g2_antennanp ANTENNA_915 (.A(_03304_));
 sg13g2_antennanp ANTENNA_916 (.A(_03354_));
 sg13g2_antennanp ANTENNA_917 (.A(_03354_));
 sg13g2_antennanp ANTENNA_918 (.A(_03354_));
 sg13g2_antennanp ANTENNA_919 (.A(_03397_));
 sg13g2_antennanp ANTENNA_920 (.A(_03397_));
 sg13g2_antennanp ANTENNA_921 (.A(_03397_));
 sg13g2_antennanp ANTENNA_922 (.A(_03535_));
 sg13g2_antennanp ANTENNA_923 (.A(_03644_));
 sg13g2_antennanp ANTENNA_924 (.A(_05221_));
 sg13g2_antennanp ANTENNA_925 (.A(_05221_));
 sg13g2_antennanp ANTENNA_926 (.A(_05221_));
 sg13g2_antennanp ANTENNA_927 (.A(_05221_));
 sg13g2_antennanp ANTENNA_928 (.A(_05221_));
 sg13g2_antennanp ANTENNA_929 (.A(_05221_));
 sg13g2_antennanp ANTENNA_930 (.A(_05300_));
 sg13g2_antennanp ANTENNA_931 (.A(_05424_));
 sg13g2_antennanp ANTENNA_932 (.A(_05424_));
 sg13g2_antennanp ANTENNA_933 (.A(_05424_));
 sg13g2_antennanp ANTENNA_934 (.A(_05424_));
 sg13g2_antennanp ANTENNA_935 (.A(_05424_));
 sg13g2_antennanp ANTENNA_936 (.A(_06065_));
 sg13g2_antennanp ANTENNA_937 (.A(_07183_));
 sg13g2_antennanp ANTENNA_938 (.A(_07183_));
 sg13g2_antennanp ANTENNA_939 (.A(_07183_));
 sg13g2_antennanp ANTENNA_940 (.A(_07183_));
 sg13g2_antennanp ANTENNA_941 (.A(_07183_));
 sg13g2_antennanp ANTENNA_942 (.A(_07183_));
 sg13g2_antennanp ANTENNA_943 (.A(_07183_));
 sg13g2_antennanp ANTENNA_944 (.A(_07183_));
 sg13g2_antennanp ANTENNA_945 (.A(_07183_));
 sg13g2_antennanp ANTENNA_946 (.A(_07183_));
 sg13g2_antennanp ANTENNA_947 (.A(_07190_));
 sg13g2_antennanp ANTENNA_948 (.A(_07312_));
 sg13g2_antennanp ANTENNA_949 (.A(_07334_));
 sg13g2_antennanp ANTENNA_950 (.A(_07334_));
 sg13g2_antennanp ANTENNA_951 (.A(_07335_));
 sg13g2_antennanp ANTENNA_952 (.A(_07335_));
 sg13g2_antennanp ANTENNA_953 (.A(clk));
 sg13g2_antennanp ANTENNA_954 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_955 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_956 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_957 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_958 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_959 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_960 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_961 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_962 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_963 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_964 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_965 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_966 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_967 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_968 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_969 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_970 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_971 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_972 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_973 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_974 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_975 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_976 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_977 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_978 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_979 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_980 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_981 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_982 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_983 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_984 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_985 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_986 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_987 (.A(net74));
 sg13g2_antennanp ANTENNA_988 (.A(net74));
 sg13g2_antennanp ANTENNA_989 (.A(net74));
 sg13g2_antennanp ANTENNA_990 (.A(net74));
 sg13g2_antennanp ANTENNA_991 (.A(net74));
 sg13g2_antennanp ANTENNA_992 (.A(net74));
 sg13g2_antennanp ANTENNA_993 (.A(net74));
 sg13g2_antennanp ANTENNA_994 (.A(net74));
 sg13g2_antennanp ANTENNA_995 (.A(net74));
 sg13g2_antennanp ANTENNA_996 (.A(net157));
 sg13g2_antennanp ANTENNA_997 (.A(net157));
 sg13g2_antennanp ANTENNA_998 (.A(net157));
 sg13g2_antennanp ANTENNA_999 (.A(net157));
 sg13g2_antennanp ANTENNA_1000 (.A(net157));
 sg13g2_antennanp ANTENNA_1001 (.A(net157));
 sg13g2_antennanp ANTENNA_1002 (.A(net157));
 sg13g2_antennanp ANTENNA_1003 (.A(net157));
 sg13g2_antennanp ANTENNA_1004 (.A(net159));
 sg13g2_antennanp ANTENNA_1005 (.A(net159));
 sg13g2_antennanp ANTENNA_1006 (.A(net159));
 sg13g2_antennanp ANTENNA_1007 (.A(net159));
 sg13g2_antennanp ANTENNA_1008 (.A(net159));
 sg13g2_antennanp ANTENNA_1009 (.A(net159));
 sg13g2_antennanp ANTENNA_1010 (.A(net159));
 sg13g2_antennanp ANTENNA_1011 (.A(net159));
 sg13g2_antennanp ANTENNA_1012 (.A(net159));
 sg13g2_antennanp ANTENNA_1013 (.A(net513));
 sg13g2_antennanp ANTENNA_1014 (.A(net513));
 sg13g2_antennanp ANTENNA_1015 (.A(net513));
 sg13g2_antennanp ANTENNA_1016 (.A(net513));
 sg13g2_antennanp ANTENNA_1017 (.A(net513));
 sg13g2_antennanp ANTENNA_1018 (.A(net513));
 sg13g2_antennanp ANTENNA_1019 (.A(net513));
 sg13g2_antennanp ANTENNA_1020 (.A(net513));
 sg13g2_antennanp ANTENNA_1021 (.A(net513));
 sg13g2_antennanp ANTENNA_1022 (.A(net549));
 sg13g2_antennanp ANTENNA_1023 (.A(net549));
 sg13g2_antennanp ANTENNA_1024 (.A(net549));
 sg13g2_antennanp ANTENNA_1025 (.A(net549));
 sg13g2_antennanp ANTENNA_1026 (.A(net549));
 sg13g2_antennanp ANTENNA_1027 (.A(net549));
 sg13g2_antennanp ANTENNA_1028 (.A(net549));
 sg13g2_antennanp ANTENNA_1029 (.A(net549));
 sg13g2_antennanp ANTENNA_1030 (.A(net549));
 sg13g2_antennanp ANTENNA_1031 (.A(net583));
 sg13g2_antennanp ANTENNA_1032 (.A(net583));
 sg13g2_antennanp ANTENNA_1033 (.A(net583));
 sg13g2_antennanp ANTENNA_1034 (.A(net583));
 sg13g2_antennanp ANTENNA_1035 (.A(net583));
 sg13g2_antennanp ANTENNA_1036 (.A(net583));
 sg13g2_antennanp ANTENNA_1037 (.A(net583));
 sg13g2_antennanp ANTENNA_1038 (.A(net583));
 sg13g2_antennanp ANTENNA_1039 (.A(net583));
 sg13g2_antennanp ANTENNA_1040 (.A(net583));
 sg13g2_antennanp ANTENNA_1041 (.A(net583));
 sg13g2_antennanp ANTENNA_1042 (.A(net583));
 sg13g2_antennanp ANTENNA_1043 (.A(net583));
 sg13g2_antennanp ANTENNA_1044 (.A(net583));
 sg13g2_antennanp ANTENNA_1045 (.A(net583));
 sg13g2_antennanp ANTENNA_1046 (.A(net583));
 sg13g2_antennanp ANTENNA_1047 (.A(net583));
 sg13g2_antennanp ANTENNA_1048 (.A(net583));
 sg13g2_antennanp ANTENNA_1049 (.A(net583));
 sg13g2_antennanp ANTENNA_1050 (.A(_00216_));
 sg13g2_antennanp ANTENNA_1051 (.A(_00216_));
 sg13g2_antennanp ANTENNA_1052 (.A(_00242_));
 sg13g2_antennanp ANTENNA_1053 (.A(_00242_));
 sg13g2_antennanp ANTENNA_1054 (.A(_00419_));
 sg13g2_antennanp ANTENNA_1055 (.A(_00419_));
 sg13g2_antennanp ANTENNA_1056 (.A(_00656_));
 sg13g2_antennanp ANTENNA_1057 (.A(_00656_));
 sg13g2_antennanp ANTENNA_1058 (.A(_00656_));
 sg13g2_antennanp ANTENNA_1059 (.A(_00680_));
 sg13g2_antennanp ANTENNA_1060 (.A(_00680_));
 sg13g2_antennanp ANTENNA_1061 (.A(_00680_));
 sg13g2_antennanp ANTENNA_1062 (.A(_00680_));
 sg13g2_antennanp ANTENNA_1063 (.A(_00680_));
 sg13g2_antennanp ANTENNA_1064 (.A(_00680_));
 sg13g2_antennanp ANTENNA_1065 (.A(_00680_));
 sg13g2_antennanp ANTENNA_1066 (.A(_00680_));
 sg13g2_antennanp ANTENNA_1067 (.A(_00680_));
 sg13g2_antennanp ANTENNA_1068 (.A(_00683_));
 sg13g2_antennanp ANTENNA_1069 (.A(_00683_));
 sg13g2_antennanp ANTENNA_1070 (.A(_00683_));
 sg13g2_antennanp ANTENNA_1071 (.A(_00683_));
 sg13g2_antennanp ANTENNA_1072 (.A(_01051_));
 sg13g2_antennanp ANTENNA_1073 (.A(_01070_));
 sg13g2_antennanp ANTENNA_1074 (.A(_01070_));
 sg13g2_antennanp ANTENNA_1075 (.A(_01071_));
 sg13g2_antennanp ANTENNA_1076 (.A(_01071_));
 sg13g2_antennanp ANTENNA_1077 (.A(_01071_));
 sg13g2_antennanp ANTENNA_1078 (.A(_01071_));
 sg13g2_antennanp ANTENNA_1079 (.A(_01178_));
 sg13g2_antennanp ANTENNA_1080 (.A(_01178_));
 sg13g2_antennanp ANTENNA_1081 (.A(_01178_));
 sg13g2_antennanp ANTENNA_1082 (.A(_01178_));
 sg13g2_antennanp ANTENNA_1083 (.A(_01212_));
 sg13g2_antennanp ANTENNA_1084 (.A(_01212_));
 sg13g2_antennanp ANTENNA_1085 (.A(_01212_));
 sg13g2_antennanp ANTENNA_1086 (.A(_01252_));
 sg13g2_antennanp ANTENNA_1087 (.A(_01252_));
 sg13g2_antennanp ANTENNA_1088 (.A(_01252_));
 sg13g2_antennanp ANTENNA_1089 (.A(_01252_));
 sg13g2_antennanp ANTENNA_1090 (.A(_01360_));
 sg13g2_antennanp ANTENNA_1091 (.A(_01360_));
 sg13g2_antennanp ANTENNA_1092 (.A(_01360_));
 sg13g2_antennanp ANTENNA_1093 (.A(_01675_));
 sg13g2_antennanp ANTENNA_1094 (.A(_01675_));
 sg13g2_antennanp ANTENNA_1095 (.A(_01675_));
 sg13g2_antennanp ANTENNA_1096 (.A(_01675_));
 sg13g2_antennanp ANTENNA_1097 (.A(_01675_));
 sg13g2_antennanp ANTENNA_1098 (.A(_01676_));
 sg13g2_antennanp ANTENNA_1099 (.A(_01676_));
 sg13g2_antennanp ANTENNA_1100 (.A(_01676_));
 sg13g2_antennanp ANTENNA_1101 (.A(_01676_));
 sg13g2_antennanp ANTENNA_1102 (.A(_01726_));
 sg13g2_antennanp ANTENNA_1103 (.A(_01726_));
 sg13g2_antennanp ANTENNA_1104 (.A(_01844_));
 sg13g2_antennanp ANTENNA_1105 (.A(_01844_));
 sg13g2_antennanp ANTENNA_1106 (.A(_01844_));
 sg13g2_antennanp ANTENNA_1107 (.A(_02395_));
 sg13g2_antennanp ANTENNA_1108 (.A(_02519_));
 sg13g2_antennanp ANTENNA_1109 (.A(_02567_));
 sg13g2_antennanp ANTENNA_1110 (.A(_02567_));
 sg13g2_antennanp ANTENNA_1111 (.A(_02567_));
 sg13g2_antennanp ANTENNA_1112 (.A(_02934_));
 sg13g2_antennanp ANTENNA_1113 (.A(_02942_));
 sg13g2_antennanp ANTENNA_1114 (.A(_02942_));
 sg13g2_antennanp ANTENNA_1115 (.A(_03065_));
 sg13g2_antennanp ANTENNA_1116 (.A(_03065_));
 sg13g2_antennanp ANTENNA_1117 (.A(_03278_));
 sg13g2_antennanp ANTENNA_1118 (.A(_03304_));
 sg13g2_antennanp ANTENNA_1119 (.A(_03304_));
 sg13g2_antennanp ANTENNA_1120 (.A(_03354_));
 sg13g2_antennanp ANTENNA_1121 (.A(_03354_));
 sg13g2_antennanp ANTENNA_1122 (.A(_03354_));
 sg13g2_antennanp ANTENNA_1123 (.A(_03397_));
 sg13g2_antennanp ANTENNA_1124 (.A(_03397_));
 sg13g2_antennanp ANTENNA_1125 (.A(_03397_));
 sg13g2_antennanp ANTENNA_1126 (.A(_03535_));
 sg13g2_antennanp ANTENNA_1127 (.A(_03644_));
 sg13g2_antennanp ANTENNA_1128 (.A(_05221_));
 sg13g2_antennanp ANTENNA_1129 (.A(_05221_));
 sg13g2_antennanp ANTENNA_1130 (.A(_05221_));
 sg13g2_antennanp ANTENNA_1131 (.A(_05221_));
 sg13g2_antennanp ANTENNA_1132 (.A(_05221_));
 sg13g2_antennanp ANTENNA_1133 (.A(_05221_));
 sg13g2_antennanp ANTENNA_1134 (.A(_05300_));
 sg13g2_antennanp ANTENNA_1135 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1136 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1137 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1138 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1139 (.A(_05424_));
 sg13g2_antennanp ANTENNA_1140 (.A(_06065_));
 sg13g2_antennanp ANTENNA_1141 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1142 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1143 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1144 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1145 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1146 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1147 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1148 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1149 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1150 (.A(_07183_));
 sg13g2_antennanp ANTENNA_1151 (.A(_07190_));
 sg13g2_antennanp ANTENNA_1152 (.A(_07312_));
 sg13g2_antennanp ANTENNA_1153 (.A(_07334_));
 sg13g2_antennanp ANTENNA_1154 (.A(_07334_));
 sg13g2_antennanp ANTENNA_1155 (.A(_07335_));
 sg13g2_antennanp ANTENNA_1156 (.A(_07335_));
 sg13g2_antennanp ANTENNA_1157 (.A(clk));
 sg13g2_antennanp ANTENNA_1158 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_1159 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_1160 (.A(\clock_inst.min_c[12] ));
 sg13g2_antennanp ANTENNA_1161 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_1162 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_1163 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_1164 (.A(\clock_inst.min_c[14] ));
 sg13g2_antennanp ANTENNA_1165 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_1166 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_1167 (.A(\clock_inst.min_c[16] ));
 sg13g2_antennanp ANTENNA_1168 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_1169 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_1170 (.A(\clock_inst.min_c[22] ));
 sg13g2_antennanp ANTENNA_1171 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_1172 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_1173 (.A(\clock_inst.min_c[25] ));
 sg13g2_antennanp ANTENNA_1174 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_1175 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_1176 (.A(\clock_inst.min_c[27] ));
 sg13g2_antennanp ANTENNA_1177 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_1178 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_1179 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_1180 (.A(\clock_inst.sec_c[11] ));
 sg13g2_antennanp ANTENNA_1181 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_1182 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_1183 (.A(\clock_inst.sec_c[16] ));
 sg13g2_antennanp ANTENNA_1184 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_1185 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_1186 (.A(\clock_inst.sec_c[48] ));
 sg13g2_antennanp ANTENNA_1187 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_1188 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_1189 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_1190 (.A(\clock_inst.vga_inst.vga_horizontal_visible ));
 sg13g2_antennanp ANTENNA_1191 (.A(net74));
 sg13g2_antennanp ANTENNA_1192 (.A(net74));
 sg13g2_antennanp ANTENNA_1193 (.A(net74));
 sg13g2_antennanp ANTENNA_1194 (.A(net74));
 sg13g2_antennanp ANTENNA_1195 (.A(net74));
 sg13g2_antennanp ANTENNA_1196 (.A(net74));
 sg13g2_antennanp ANTENNA_1197 (.A(net74));
 sg13g2_antennanp ANTENNA_1198 (.A(net74));
 sg13g2_antennanp ANTENNA_1199 (.A(net74));
 sg13g2_antennanp ANTENNA_1200 (.A(net157));
 sg13g2_antennanp ANTENNA_1201 (.A(net157));
 sg13g2_antennanp ANTENNA_1202 (.A(net157));
 sg13g2_antennanp ANTENNA_1203 (.A(net157));
 sg13g2_antennanp ANTENNA_1204 (.A(net157));
 sg13g2_antennanp ANTENNA_1205 (.A(net157));
 sg13g2_antennanp ANTENNA_1206 (.A(net157));
 sg13g2_antennanp ANTENNA_1207 (.A(net157));
 sg13g2_antennanp ANTENNA_1208 (.A(net513));
 sg13g2_antennanp ANTENNA_1209 (.A(net513));
 sg13g2_antennanp ANTENNA_1210 (.A(net513));
 sg13g2_antennanp ANTENNA_1211 (.A(net513));
 sg13g2_antennanp ANTENNA_1212 (.A(net513));
 sg13g2_antennanp ANTENNA_1213 (.A(net513));
 sg13g2_antennanp ANTENNA_1214 (.A(net513));
 sg13g2_antennanp ANTENNA_1215 (.A(net513));
 sg13g2_antennanp ANTENNA_1216 (.A(net513));
 sg13g2_antennanp ANTENNA_1217 (.A(net549));
 sg13g2_antennanp ANTENNA_1218 (.A(net549));
 sg13g2_antennanp ANTENNA_1219 (.A(net549));
 sg13g2_antennanp ANTENNA_1220 (.A(net549));
 sg13g2_antennanp ANTENNA_1221 (.A(net549));
 sg13g2_antennanp ANTENNA_1222 (.A(net549));
 sg13g2_antennanp ANTENNA_1223 (.A(net549));
 sg13g2_antennanp ANTENNA_1224 (.A(net549));
 sg13g2_antennanp ANTENNA_1225 (.A(net549));
 sg13g2_antennanp ANTENNA_1226 (.A(net583));
 sg13g2_antennanp ANTENNA_1227 (.A(net583));
 sg13g2_antennanp ANTENNA_1228 (.A(net583));
 sg13g2_antennanp ANTENNA_1229 (.A(net583));
 sg13g2_antennanp ANTENNA_1230 (.A(net583));
 sg13g2_antennanp ANTENNA_1231 (.A(net583));
 sg13g2_antennanp ANTENNA_1232 (.A(net583));
 sg13g2_antennanp ANTENNA_1233 (.A(net583));
 sg13g2_antennanp ANTENNA_1234 (.A(net583));
 sg13g2_antennanp ANTENNA_1235 (.A(net583));
 sg13g2_antennanp ANTENNA_1236 (.A(net583));
 sg13g2_antennanp ANTENNA_1237 (.A(net583));
 sg13g2_antennanp ANTENNA_1238 (.A(net583));
 sg13g2_antennanp ANTENNA_1239 (.A(net583));
 sg13g2_antennanp ANTENNA_1240 (.A(net583));
 sg13g2_antennanp ANTENNA_1241 (.A(net583));
 sg13g2_antennanp ANTENNA_1242 (.A(net583));
 sg13g2_antennanp ANTENNA_1243 (.A(net583));
 sg13g2_antennanp ANTENNA_1244 (.A(net583));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_4 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_216 ();
 sg13g2_decap_8 FILLER_0_223 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_decap_4 FILLER_0_237 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_fill_2 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_8 FILLER_0_425 ();
 sg13g2_decap_8 FILLER_0_432 ();
 sg13g2_decap_8 FILLER_0_439 ();
 sg13g2_decap_8 FILLER_0_446 ();
 sg13g2_decap_8 FILLER_0_453 ();
 sg13g2_decap_4 FILLER_0_460 ();
 sg13g2_fill_2 FILLER_0_464 ();
 sg13g2_decap_8 FILLER_0_470 ();
 sg13g2_decap_8 FILLER_0_477 ();
 sg13g2_fill_2 FILLER_0_484 ();
 sg13g2_decap_4 FILLER_0_490 ();
 sg13g2_fill_1 FILLER_0_494 ();
 sg13g2_decap_4 FILLER_0_499 ();
 sg13g2_fill_2 FILLER_0_503 ();
 sg13g2_decap_8 FILLER_0_509 ();
 sg13g2_decap_8 FILLER_0_516 ();
 sg13g2_decap_8 FILLER_0_523 ();
 sg13g2_decap_8 FILLER_0_530 ();
 sg13g2_decap_8 FILLER_0_537 ();
 sg13g2_decap_8 FILLER_0_548 ();
 sg13g2_decap_8 FILLER_0_555 ();
 sg13g2_decap_8 FILLER_0_562 ();
 sg13g2_decap_8 FILLER_0_569 ();
 sg13g2_decap_8 FILLER_0_580 ();
 sg13g2_fill_2 FILLER_0_587 ();
 sg13g2_fill_1 FILLER_0_589 ();
 sg13g2_decap_8 FILLER_0_594 ();
 sg13g2_decap_8 FILLER_0_601 ();
 sg13g2_decap_8 FILLER_0_608 ();
 sg13g2_decap_8 FILLER_0_615 ();
 sg13g2_decap_8 FILLER_0_622 ();
 sg13g2_decap_8 FILLER_0_629 ();
 sg13g2_decap_8 FILLER_0_636 ();
 sg13g2_decap_8 FILLER_0_643 ();
 sg13g2_decap_8 FILLER_0_650 ();
 sg13g2_decap_4 FILLER_0_657 ();
 sg13g2_fill_1 FILLER_0_661 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_8 FILLER_0_673 ();
 sg13g2_decap_8 FILLER_0_680 ();
 sg13g2_decap_8 FILLER_0_687 ();
 sg13g2_decap_4 FILLER_0_694 ();
 sg13g2_fill_1 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_703 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_773 ();
 sg13g2_fill_2 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_786 ();
 sg13g2_decap_8 FILLER_0_793 ();
 sg13g2_decap_8 FILLER_0_800 ();
 sg13g2_decap_8 FILLER_0_807 ();
 sg13g2_decap_8 FILLER_0_814 ();
 sg13g2_decap_8 FILLER_0_821 ();
 sg13g2_decap_8 FILLER_0_828 ();
 sg13g2_decap_8 FILLER_0_835 ();
 sg13g2_fill_1 FILLER_0_842 ();
 sg13g2_fill_2 FILLER_0_853 ();
 sg13g2_fill_1 FILLER_0_855 ();
 sg13g2_fill_2 FILLER_0_865 ();
 sg13g2_decap_8 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_0_884 ();
 sg13g2_decap_8 FILLER_0_891 ();
 sg13g2_decap_8 FILLER_0_898 ();
 sg13g2_decap_8 FILLER_0_905 ();
 sg13g2_decap_8 FILLER_0_920 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_4 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_999 ();
 sg13g2_decap_8 FILLER_0_1006 ();
 sg13g2_decap_8 FILLER_0_1013 ();
 sg13g2_decap_8 FILLER_0_1024 ();
 sg13g2_decap_8 FILLER_0_1031 ();
 sg13g2_decap_8 FILLER_0_1038 ();
 sg13g2_decap_8 FILLER_0_1045 ();
 sg13g2_decap_8 FILLER_0_1052 ();
 sg13g2_decap_8 FILLER_0_1059 ();
 sg13g2_decap_8 FILLER_0_1066 ();
 sg13g2_decap_8 FILLER_0_1073 ();
 sg13g2_decap_8 FILLER_0_1080 ();
 sg13g2_decap_8 FILLER_0_1087 ();
 sg13g2_decap_8 FILLER_0_1094 ();
 sg13g2_decap_8 FILLER_0_1101 ();
 sg13g2_decap_8 FILLER_0_1108 ();
 sg13g2_fill_2 FILLER_0_1115 ();
 sg13g2_fill_1 FILLER_0_1117 ();
 sg13g2_decap_8 FILLER_0_1124 ();
 sg13g2_decap_8 FILLER_0_1131 ();
 sg13g2_decap_8 FILLER_0_1142 ();
 sg13g2_decap_8 FILLER_0_1149 ();
 sg13g2_decap_8 FILLER_0_1156 ();
 sg13g2_decap_8 FILLER_0_1163 ();
 sg13g2_decap_8 FILLER_0_1170 ();
 sg13g2_decap_8 FILLER_0_1181 ();
 sg13g2_decap_8 FILLER_0_1188 ();
 sg13g2_decap_8 FILLER_0_1195 ();
 sg13g2_decap_8 FILLER_0_1202 ();
 sg13g2_decap_8 FILLER_0_1213 ();
 sg13g2_decap_8 FILLER_0_1220 ();
 sg13g2_fill_2 FILLER_0_1227 ();
 sg13g2_decap_8 FILLER_0_1233 ();
 sg13g2_decap_8 FILLER_0_1240 ();
 sg13g2_decap_4 FILLER_0_1247 ();
 sg13g2_decap_8 FILLER_0_1263 ();
 sg13g2_decap_8 FILLER_0_1270 ();
 sg13g2_decap_8 FILLER_0_1277 ();
 sg13g2_decap_8 FILLER_0_1284 ();
 sg13g2_decap_8 FILLER_0_1291 ();
 sg13g2_decap_8 FILLER_0_1298 ();
 sg13g2_decap_4 FILLER_0_1305 ();
 sg13g2_decap_8 FILLER_0_1313 ();
 sg13g2_decap_8 FILLER_0_1320 ();
 sg13g2_decap_8 FILLER_0_1327 ();
 sg13g2_decap_8 FILLER_0_1334 ();
 sg13g2_decap_8 FILLER_0_1341 ();
 sg13g2_decap_8 FILLER_0_1348 ();
 sg13g2_decap_8 FILLER_0_1355 ();
 sg13g2_decap_8 FILLER_0_1362 ();
 sg13g2_decap_8 FILLER_0_1369 ();
 sg13g2_decap_8 FILLER_0_1376 ();
 sg13g2_decap_8 FILLER_0_1383 ();
 sg13g2_decap_8 FILLER_0_1390 ();
 sg13g2_decap_8 FILLER_0_1397 ();
 sg13g2_decap_8 FILLER_0_1404 ();
 sg13g2_decap_8 FILLER_0_1411 ();
 sg13g2_decap_8 FILLER_0_1418 ();
 sg13g2_decap_8 FILLER_0_1425 ();
 sg13g2_decap_8 FILLER_0_1432 ();
 sg13g2_decap_8 FILLER_0_1439 ();
 sg13g2_decap_8 FILLER_0_1446 ();
 sg13g2_decap_8 FILLER_0_1453 ();
 sg13g2_decap_8 FILLER_0_1460 ();
 sg13g2_decap_8 FILLER_0_1467 ();
 sg13g2_decap_8 FILLER_0_1474 ();
 sg13g2_decap_8 FILLER_0_1481 ();
 sg13g2_decap_8 FILLER_0_1488 ();
 sg13g2_decap_8 FILLER_0_1495 ();
 sg13g2_decap_8 FILLER_0_1502 ();
 sg13g2_decap_8 FILLER_0_1509 ();
 sg13g2_decap_8 FILLER_0_1516 ();
 sg13g2_decap_8 FILLER_0_1523 ();
 sg13g2_decap_8 FILLER_0_1530 ();
 sg13g2_decap_8 FILLER_0_1537 ();
 sg13g2_decap_8 FILLER_0_1544 ();
 sg13g2_decap_8 FILLER_0_1551 ();
 sg13g2_decap_8 FILLER_0_1558 ();
 sg13g2_decap_8 FILLER_0_1565 ();
 sg13g2_decap_8 FILLER_0_1572 ();
 sg13g2_decap_8 FILLER_0_1579 ();
 sg13g2_decap_8 FILLER_0_1586 ();
 sg13g2_decap_8 FILLER_0_1593 ();
 sg13g2_decap_8 FILLER_0_1600 ();
 sg13g2_decap_8 FILLER_0_1607 ();
 sg13g2_decap_8 FILLER_0_1614 ();
 sg13g2_decap_8 FILLER_0_1621 ();
 sg13g2_decap_8 FILLER_0_1628 ();
 sg13g2_decap_8 FILLER_0_1635 ();
 sg13g2_decap_8 FILLER_0_1642 ();
 sg13g2_decap_8 FILLER_0_1649 ();
 sg13g2_decap_8 FILLER_0_1656 ();
 sg13g2_decap_8 FILLER_0_1663 ();
 sg13g2_decap_8 FILLER_0_1670 ();
 sg13g2_decap_8 FILLER_0_1677 ();
 sg13g2_decap_8 FILLER_0_1684 ();
 sg13g2_decap_8 FILLER_0_1691 ();
 sg13g2_decap_8 FILLER_0_1698 ();
 sg13g2_decap_8 FILLER_0_1705 ();
 sg13g2_decap_8 FILLER_0_1712 ();
 sg13g2_decap_8 FILLER_0_1719 ();
 sg13g2_decap_8 FILLER_0_1726 ();
 sg13g2_decap_8 FILLER_0_1733 ();
 sg13g2_decap_8 FILLER_0_1740 ();
 sg13g2_decap_8 FILLER_0_1747 ();
 sg13g2_decap_8 FILLER_0_1754 ();
 sg13g2_decap_8 FILLER_0_1761 ();
 sg13g2_decap_4 FILLER_0_1768 ();
 sg13g2_fill_2 FILLER_0_1772 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_fill_2 FILLER_1_105 ();
 sg13g2_fill_1 FILLER_1_107 ();
 sg13g2_decap_4 FILLER_1_116 ();
 sg13g2_fill_1 FILLER_1_120 ();
 sg13g2_decap_8 FILLER_1_125 ();
 sg13g2_decap_8 FILLER_1_132 ();
 sg13g2_decap_8 FILLER_1_139 ();
 sg13g2_decap_8 FILLER_1_146 ();
 sg13g2_decap_8 FILLER_1_153 ();
 sg13g2_fill_1 FILLER_1_160 ();
 sg13g2_fill_2 FILLER_1_165 ();
 sg13g2_fill_1 FILLER_1_167 ();
 sg13g2_decap_8 FILLER_1_173 ();
 sg13g2_decap_8 FILLER_1_180 ();
 sg13g2_decap_8 FILLER_1_187 ();
 sg13g2_fill_2 FILLER_1_194 ();
 sg13g2_fill_1 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_205 ();
 sg13g2_decap_4 FILLER_1_212 ();
 sg13g2_fill_2 FILLER_1_216 ();
 sg13g2_fill_1 FILLER_1_223 ();
 sg13g2_fill_2 FILLER_1_228 ();
 sg13g2_fill_1 FILLER_1_230 ();
 sg13g2_fill_2 FILLER_1_237 ();
 sg13g2_fill_1 FILLER_1_239 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_4 FILLER_1_266 ();
 sg13g2_fill_2 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_fill_2 FILLER_1_301 ();
 sg13g2_decap_4 FILLER_1_321 ();
 sg13g2_fill_1 FILLER_1_325 ();
 sg13g2_decap_4 FILLER_1_330 ();
 sg13g2_fill_2 FILLER_1_334 ();
 sg13g2_decap_8 FILLER_1_340 ();
 sg13g2_decap_8 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_354 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_4 FILLER_1_375 ();
 sg13g2_fill_2 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_decap_8 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_1_435 ();
 sg13g2_decap_8 FILLER_1_442 ();
 sg13g2_decap_4 FILLER_1_449 ();
 sg13g2_fill_1 FILLER_1_458 ();
 sg13g2_fill_2 FILLER_1_490 ();
 sg13g2_fill_1 FILLER_1_492 ();
 sg13g2_decap_8 FILLER_1_528 ();
 sg13g2_fill_2 FILLER_1_535 ();
 sg13g2_fill_1 FILLER_1_537 ();
 sg13g2_decap_4 FILLER_1_572 ();
 sg13g2_fill_2 FILLER_1_581 ();
 sg13g2_fill_1 FILLER_1_583 ();
 sg13g2_decap_8 FILLER_1_610 ();
 sg13g2_fill_2 FILLER_1_617 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_4 FILLER_1_682 ();
 sg13g2_fill_2 FILLER_1_686 ();
 sg13g2_fill_2 FILLER_1_691 ();
 sg13g2_fill_2 FILLER_1_719 ();
 sg13g2_decap_4 FILLER_1_734 ();
 sg13g2_fill_1 FILLER_1_738 ();
 sg13g2_decap_8 FILLER_1_754 ();
 sg13g2_fill_1 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_806 ();
 sg13g2_decap_8 FILLER_1_813 ();
 sg13g2_fill_1 FILLER_1_820 ();
 sg13g2_fill_1 FILLER_1_831 ();
 sg13g2_decap_8 FILLER_1_856 ();
 sg13g2_fill_1 FILLER_1_863 ();
 sg13g2_fill_1 FILLER_1_872 ();
 sg13g2_fill_1 FILLER_1_877 ();
 sg13g2_fill_2 FILLER_1_883 ();
 sg13g2_decap_4 FILLER_1_893 ();
 sg13g2_fill_1 FILLER_1_897 ();
 sg13g2_decap_4 FILLER_1_903 ();
 sg13g2_fill_2 FILLER_1_907 ();
 sg13g2_decap_8 FILLER_1_939 ();
 sg13g2_decap_8 FILLER_1_946 ();
 sg13g2_decap_8 FILLER_1_953 ();
 sg13g2_fill_1 FILLER_1_960 ();
 sg13g2_decap_8 FILLER_1_970 ();
 sg13g2_fill_2 FILLER_1_977 ();
 sg13g2_fill_1 FILLER_1_979 ();
 sg13g2_decap_8 FILLER_1_984 ();
 sg13g2_fill_2 FILLER_1_991 ();
 sg13g2_decap_8 FILLER_1_998 ();
 sg13g2_decap_4 FILLER_1_1005 ();
 sg13g2_fill_2 FILLER_1_1009 ();
 sg13g2_decap_8 FILLER_1_1042 ();
 sg13g2_decap_4 FILLER_1_1049 ();
 sg13g2_fill_1 FILLER_1_1053 ();
 sg13g2_decap_4 FILLER_1_1060 ();
 sg13g2_decap_4 FILLER_1_1067 ();
 sg13g2_fill_2 FILLER_1_1071 ();
 sg13g2_decap_8 FILLER_1_1097 ();
 sg13g2_decap_8 FILLER_1_1104 ();
 sg13g2_fill_1 FILLER_1_1111 ();
 sg13g2_decap_8 FILLER_1_1161 ();
 sg13g2_fill_2 FILLER_1_1168 ();
 sg13g2_fill_1 FILLER_1_1170 ();
 sg13g2_decap_4 FILLER_1_1197 ();
 sg13g2_fill_1 FILLER_1_1201 ();
 sg13g2_fill_1 FILLER_1_1228 ();
 sg13g2_fill_1 FILLER_1_1241 ();
 sg13g2_decap_4 FILLER_1_1250 ();
 sg13g2_fill_1 FILLER_1_1254 ();
 sg13g2_fill_2 FILLER_1_1259 ();
 sg13g2_fill_1 FILLER_1_1261 ();
 sg13g2_decap_4 FILLER_1_1284 ();
 sg13g2_fill_2 FILLER_1_1292 ();
 sg13g2_decap_8 FILLER_1_1328 ();
 sg13g2_decap_8 FILLER_1_1335 ();
 sg13g2_decap_8 FILLER_1_1342 ();
 sg13g2_decap_8 FILLER_1_1349 ();
 sg13g2_decap_8 FILLER_1_1356 ();
 sg13g2_decap_8 FILLER_1_1363 ();
 sg13g2_decap_8 FILLER_1_1370 ();
 sg13g2_decap_8 FILLER_1_1377 ();
 sg13g2_decap_8 FILLER_1_1384 ();
 sg13g2_decap_8 FILLER_1_1391 ();
 sg13g2_decap_8 FILLER_1_1398 ();
 sg13g2_decap_8 FILLER_1_1405 ();
 sg13g2_decap_8 FILLER_1_1412 ();
 sg13g2_decap_8 FILLER_1_1419 ();
 sg13g2_decap_8 FILLER_1_1426 ();
 sg13g2_decap_8 FILLER_1_1433 ();
 sg13g2_decap_8 FILLER_1_1440 ();
 sg13g2_decap_8 FILLER_1_1447 ();
 sg13g2_decap_8 FILLER_1_1454 ();
 sg13g2_decap_8 FILLER_1_1461 ();
 sg13g2_decap_8 FILLER_1_1468 ();
 sg13g2_decap_8 FILLER_1_1475 ();
 sg13g2_decap_8 FILLER_1_1482 ();
 sg13g2_decap_8 FILLER_1_1489 ();
 sg13g2_decap_8 FILLER_1_1496 ();
 sg13g2_decap_8 FILLER_1_1503 ();
 sg13g2_decap_8 FILLER_1_1510 ();
 sg13g2_decap_8 FILLER_1_1517 ();
 sg13g2_decap_8 FILLER_1_1524 ();
 sg13g2_decap_8 FILLER_1_1531 ();
 sg13g2_decap_8 FILLER_1_1538 ();
 sg13g2_decap_8 FILLER_1_1545 ();
 sg13g2_decap_8 FILLER_1_1552 ();
 sg13g2_decap_8 FILLER_1_1559 ();
 sg13g2_decap_8 FILLER_1_1566 ();
 sg13g2_decap_8 FILLER_1_1573 ();
 sg13g2_decap_8 FILLER_1_1580 ();
 sg13g2_decap_8 FILLER_1_1587 ();
 sg13g2_decap_8 FILLER_1_1594 ();
 sg13g2_decap_8 FILLER_1_1601 ();
 sg13g2_decap_8 FILLER_1_1608 ();
 sg13g2_decap_8 FILLER_1_1615 ();
 sg13g2_decap_8 FILLER_1_1622 ();
 sg13g2_decap_8 FILLER_1_1629 ();
 sg13g2_decap_8 FILLER_1_1636 ();
 sg13g2_decap_8 FILLER_1_1643 ();
 sg13g2_decap_8 FILLER_1_1650 ();
 sg13g2_decap_8 FILLER_1_1657 ();
 sg13g2_decap_8 FILLER_1_1664 ();
 sg13g2_decap_8 FILLER_1_1671 ();
 sg13g2_decap_8 FILLER_1_1678 ();
 sg13g2_decap_8 FILLER_1_1685 ();
 sg13g2_decap_8 FILLER_1_1692 ();
 sg13g2_decap_8 FILLER_1_1699 ();
 sg13g2_decap_8 FILLER_1_1706 ();
 sg13g2_decap_8 FILLER_1_1713 ();
 sg13g2_decap_8 FILLER_1_1720 ();
 sg13g2_decap_8 FILLER_1_1727 ();
 sg13g2_decap_8 FILLER_1_1734 ();
 sg13g2_decap_8 FILLER_1_1741 ();
 sg13g2_decap_8 FILLER_1_1748 ();
 sg13g2_decap_8 FILLER_1_1755 ();
 sg13g2_decap_8 FILLER_1_1762 ();
 sg13g2_decap_4 FILLER_1_1769 ();
 sg13g2_fill_1 FILLER_1_1773 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_fill_1 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_96 ();
 sg13g2_decap_4 FILLER_2_103 ();
 sg13g2_decap_8 FILLER_2_111 ();
 sg13g2_fill_2 FILLER_2_118 ();
 sg13g2_decap_8 FILLER_2_125 ();
 sg13g2_fill_2 FILLER_2_132 ();
 sg13g2_fill_1 FILLER_2_134 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_fill_2 FILLER_2_151 ();
 sg13g2_fill_1 FILLER_2_153 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_fill_1 FILLER_2_181 ();
 sg13g2_decap_4 FILLER_2_187 ();
 sg13g2_fill_1 FILLER_2_191 ();
 sg13g2_fill_1 FILLER_2_225 ();
 sg13g2_decap_8 FILLER_2_250 ();
 sg13g2_decap_4 FILLER_2_257 ();
 sg13g2_fill_2 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_267 ();
 sg13g2_decap_8 FILLER_2_279 ();
 sg13g2_decap_4 FILLER_2_286 ();
 sg13g2_fill_1 FILLER_2_300 ();
 sg13g2_fill_2 FILLER_2_309 ();
 sg13g2_fill_1 FILLER_2_311 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_fill_1 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_341 ();
 sg13g2_decap_8 FILLER_2_348 ();
 sg13g2_fill_2 FILLER_2_355 ();
 sg13g2_fill_2 FILLER_2_366 ();
 sg13g2_fill_1 FILLER_2_368 ();
 sg13g2_fill_2 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_4 FILLER_2_395 ();
 sg13g2_fill_1 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_decap_4 FILLER_2_416 ();
 sg13g2_fill_1 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_2_433 ();
 sg13g2_decap_8 FILLER_2_440 ();
 sg13g2_decap_8 FILLER_2_447 ();
 sg13g2_decap_8 FILLER_2_454 ();
 sg13g2_decap_8 FILLER_2_461 ();
 sg13g2_decap_8 FILLER_2_468 ();
 sg13g2_decap_8 FILLER_2_475 ();
 sg13g2_decap_8 FILLER_2_482 ();
 sg13g2_decap_8 FILLER_2_489 ();
 sg13g2_decap_8 FILLER_2_496 ();
 sg13g2_decap_8 FILLER_2_503 ();
 sg13g2_decap_8 FILLER_2_514 ();
 sg13g2_decap_8 FILLER_2_521 ();
 sg13g2_decap_8 FILLER_2_528 ();
 sg13g2_decap_8 FILLER_2_535 ();
 sg13g2_decap_8 FILLER_2_542 ();
 sg13g2_fill_1 FILLER_2_549 ();
 sg13g2_decap_8 FILLER_2_594 ();
 sg13g2_decap_4 FILLER_2_601 ();
 sg13g2_decap_4 FILLER_2_610 ();
 sg13g2_decap_8 FILLER_2_645 ();
 sg13g2_decap_8 FILLER_2_652 ();
 sg13g2_decap_8 FILLER_2_659 ();
 sg13g2_decap_8 FILLER_2_666 ();
 sg13g2_fill_2 FILLER_2_673 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_fill_2 FILLER_2_707 ();
 sg13g2_fill_1 FILLER_2_709 ();
 sg13g2_fill_2 FILLER_2_718 ();
 sg13g2_fill_1 FILLER_2_720 ();
 sg13g2_fill_2 FILLER_2_725 ();
 sg13g2_fill_1 FILLER_2_727 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_fill_1 FILLER_2_760 ();
 sg13g2_decap_4 FILLER_2_774 ();
 sg13g2_fill_2 FILLER_2_790 ();
 sg13g2_fill_1 FILLER_2_792 ();
 sg13g2_fill_2 FILLER_2_803 ();
 sg13g2_fill_1 FILLER_2_810 ();
 sg13g2_fill_2 FILLER_2_816 ();
 sg13g2_fill_1 FILLER_2_818 ();
 sg13g2_decap_8 FILLER_2_824 ();
 sg13g2_decap_8 FILLER_2_831 ();
 sg13g2_decap_8 FILLER_2_838 ();
 sg13g2_decap_8 FILLER_2_845 ();
 sg13g2_decap_4 FILLER_2_852 ();
 sg13g2_fill_2 FILLER_2_856 ();
 sg13g2_decap_8 FILLER_2_870 ();
 sg13g2_decap_8 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_2_884 ();
 sg13g2_fill_1 FILLER_2_891 ();
 sg13g2_decap_4 FILLER_2_896 ();
 sg13g2_decap_8 FILLER_2_908 ();
 sg13g2_fill_1 FILLER_2_915 ();
 sg13g2_decap_8 FILLER_2_922 ();
 sg13g2_decap_8 FILLER_2_929 ();
 sg13g2_decap_8 FILLER_2_936 ();
 sg13g2_decap_8 FILLER_2_943 ();
 sg13g2_decap_8 FILLER_2_950 ();
 sg13g2_decap_8 FILLER_2_957 ();
 sg13g2_fill_2 FILLER_2_964 ();
 sg13g2_decap_8 FILLER_2_990 ();
 sg13g2_decap_8 FILLER_2_997 ();
 sg13g2_decap_8 FILLER_2_1004 ();
 sg13g2_decap_8 FILLER_2_1011 ();
 sg13g2_fill_2 FILLER_2_1018 ();
 sg13g2_fill_2 FILLER_2_1028 ();
 sg13g2_decap_4 FILLER_2_1035 ();
 sg13g2_fill_1 FILLER_2_1050 ();
 sg13g2_decap_8 FILLER_2_1059 ();
 sg13g2_fill_1 FILLER_2_1066 ();
 sg13g2_fill_2 FILLER_2_1074 ();
 sg13g2_decap_8 FILLER_2_1085 ();
 sg13g2_decap_8 FILLER_2_1092 ();
 sg13g2_decap_8 FILLER_2_1099 ();
 sg13g2_fill_2 FILLER_2_1106 ();
 sg13g2_fill_1 FILLER_2_1108 ();
 sg13g2_fill_1 FILLER_2_1135 ();
 sg13g2_decap_8 FILLER_2_1139 ();
 sg13g2_decap_8 FILLER_2_1146 ();
 sg13g2_decap_8 FILLER_2_1153 ();
 sg13g2_decap_4 FILLER_2_1160 ();
 sg13g2_decap_4 FILLER_2_1176 ();
 sg13g2_decap_8 FILLER_2_1188 ();
 sg13g2_fill_1 FILLER_2_1195 ();
 sg13g2_decap_8 FILLER_2_1205 ();
 sg13g2_decap_8 FILLER_2_1212 ();
 sg13g2_decap_8 FILLER_2_1219 ();
 sg13g2_decap_8 FILLER_2_1226 ();
 sg13g2_decap_8 FILLER_2_1233 ();
 sg13g2_decap_8 FILLER_2_1240 ();
 sg13g2_decap_8 FILLER_2_1247 ();
 sg13g2_decap_4 FILLER_2_1269 ();
 sg13g2_fill_2 FILLER_2_1273 ();
 sg13g2_decap_8 FILLER_2_1280 ();
 sg13g2_decap_8 FILLER_2_1287 ();
 sg13g2_fill_2 FILLER_2_1294 ();
 sg13g2_fill_1 FILLER_2_1296 ();
 sg13g2_decap_8 FILLER_2_1302 ();
 sg13g2_fill_1 FILLER_2_1309 ();
 sg13g2_decap_8 FILLER_2_1314 ();
 sg13g2_decap_8 FILLER_2_1321 ();
 sg13g2_decap_8 FILLER_2_1328 ();
 sg13g2_fill_2 FILLER_2_1335 ();
 sg13g2_decap_8 FILLER_2_1341 ();
 sg13g2_decap_8 FILLER_2_1348 ();
 sg13g2_decap_8 FILLER_2_1355 ();
 sg13g2_decap_8 FILLER_2_1362 ();
 sg13g2_decap_8 FILLER_2_1369 ();
 sg13g2_decap_8 FILLER_2_1376 ();
 sg13g2_decap_8 FILLER_2_1383 ();
 sg13g2_decap_8 FILLER_2_1390 ();
 sg13g2_decap_8 FILLER_2_1397 ();
 sg13g2_decap_4 FILLER_2_1404 ();
 sg13g2_decap_8 FILLER_2_1412 ();
 sg13g2_decap_8 FILLER_2_1419 ();
 sg13g2_decap_8 FILLER_2_1426 ();
 sg13g2_decap_8 FILLER_2_1433 ();
 sg13g2_decap_8 FILLER_2_1440 ();
 sg13g2_decap_8 FILLER_2_1447 ();
 sg13g2_decap_8 FILLER_2_1454 ();
 sg13g2_decap_8 FILLER_2_1461 ();
 sg13g2_decap_8 FILLER_2_1468 ();
 sg13g2_decap_8 FILLER_2_1475 ();
 sg13g2_decap_8 FILLER_2_1482 ();
 sg13g2_decap_8 FILLER_2_1489 ();
 sg13g2_decap_8 FILLER_2_1496 ();
 sg13g2_decap_8 FILLER_2_1503 ();
 sg13g2_decap_8 FILLER_2_1510 ();
 sg13g2_decap_8 FILLER_2_1517 ();
 sg13g2_decap_8 FILLER_2_1524 ();
 sg13g2_decap_8 FILLER_2_1531 ();
 sg13g2_decap_8 FILLER_2_1538 ();
 sg13g2_decap_8 FILLER_2_1545 ();
 sg13g2_decap_8 FILLER_2_1552 ();
 sg13g2_decap_8 FILLER_2_1559 ();
 sg13g2_decap_8 FILLER_2_1566 ();
 sg13g2_decap_8 FILLER_2_1573 ();
 sg13g2_decap_8 FILLER_2_1580 ();
 sg13g2_decap_8 FILLER_2_1587 ();
 sg13g2_decap_8 FILLER_2_1594 ();
 sg13g2_decap_8 FILLER_2_1601 ();
 sg13g2_decap_8 FILLER_2_1608 ();
 sg13g2_decap_8 FILLER_2_1615 ();
 sg13g2_decap_8 FILLER_2_1622 ();
 sg13g2_decap_8 FILLER_2_1629 ();
 sg13g2_decap_8 FILLER_2_1636 ();
 sg13g2_decap_8 FILLER_2_1643 ();
 sg13g2_decap_8 FILLER_2_1650 ();
 sg13g2_decap_8 FILLER_2_1657 ();
 sg13g2_decap_8 FILLER_2_1664 ();
 sg13g2_decap_8 FILLER_2_1671 ();
 sg13g2_decap_8 FILLER_2_1678 ();
 sg13g2_decap_8 FILLER_2_1685 ();
 sg13g2_decap_8 FILLER_2_1692 ();
 sg13g2_decap_8 FILLER_2_1699 ();
 sg13g2_decap_8 FILLER_2_1706 ();
 sg13g2_decap_8 FILLER_2_1713 ();
 sg13g2_decap_8 FILLER_2_1720 ();
 sg13g2_decap_8 FILLER_2_1727 ();
 sg13g2_decap_8 FILLER_2_1734 ();
 sg13g2_decap_8 FILLER_2_1741 ();
 sg13g2_decap_8 FILLER_2_1748 ();
 sg13g2_decap_8 FILLER_2_1755 ();
 sg13g2_decap_8 FILLER_2_1762 ();
 sg13g2_decap_4 FILLER_2_1769 ();
 sg13g2_fill_1 FILLER_2_1773 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_4 FILLER_3_84 ();
 sg13g2_fill_1 FILLER_3_88 ();
 sg13g2_decap_4 FILLER_3_101 ();
 sg13g2_decap_8 FILLER_3_115 ();
 sg13g2_decap_8 FILLER_3_122 ();
 sg13g2_decap_4 FILLER_3_129 ();
 sg13g2_fill_2 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_156 ();
 sg13g2_decap_8 FILLER_3_170 ();
 sg13g2_fill_2 FILLER_3_177 ();
 sg13g2_fill_1 FILLER_3_184 ();
 sg13g2_decap_4 FILLER_3_194 ();
 sg13g2_fill_2 FILLER_3_198 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_4 FILLER_3_221 ();
 sg13g2_fill_2 FILLER_3_225 ();
 sg13g2_decap_4 FILLER_3_232 ();
 sg13g2_fill_1 FILLER_3_236 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_fill_1 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_269 ();
 sg13g2_decap_8 FILLER_3_276 ();
 sg13g2_decap_4 FILLER_3_283 ();
 sg13g2_fill_1 FILLER_3_287 ();
 sg13g2_decap_4 FILLER_3_298 ();
 sg13g2_fill_1 FILLER_3_302 ();
 sg13g2_decap_8 FILLER_3_316 ();
 sg13g2_decap_8 FILLER_3_323 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_fill_2 FILLER_3_368 ();
 sg13g2_decap_4 FILLER_3_375 ();
 sg13g2_fill_2 FILLER_3_379 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_1 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_8 FILLER_3_424 ();
 sg13g2_decap_8 FILLER_3_431 ();
 sg13g2_fill_1 FILLER_3_438 ();
 sg13g2_decap_8 FILLER_3_451 ();
 sg13g2_decap_8 FILLER_3_458 ();
 sg13g2_fill_1 FILLER_3_465 ();
 sg13g2_decap_8 FILLER_3_470 ();
 sg13g2_decap_8 FILLER_3_477 ();
 sg13g2_fill_2 FILLER_3_484 ();
 sg13g2_fill_1 FILLER_3_486 ();
 sg13g2_fill_2 FILLER_3_491 ();
 sg13g2_fill_1 FILLER_3_498 ();
 sg13g2_fill_1 FILLER_3_525 ();
 sg13g2_fill_1 FILLER_3_530 ();
 sg13g2_fill_2 FILLER_3_557 ();
 sg13g2_fill_1 FILLER_3_564 ();
 sg13g2_decap_4 FILLER_3_570 ();
 sg13g2_fill_1 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_579 ();
 sg13g2_decap_4 FILLER_3_586 ();
 sg13g2_fill_1 FILLER_3_590 ();
 sg13g2_decap_8 FILLER_3_596 ();
 sg13g2_decap_4 FILLER_3_608 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_4 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_657 ();
 sg13g2_decap_4 FILLER_3_664 ();
 sg13g2_fill_2 FILLER_3_694 ();
 sg13g2_fill_1 FILLER_3_696 ();
 sg13g2_decap_8 FILLER_3_701 ();
 sg13g2_decap_8 FILLER_3_708 ();
 sg13g2_decap_8 FILLER_3_715 ();
 sg13g2_decap_8 FILLER_3_722 ();
 sg13g2_decap_8 FILLER_3_729 ();
 sg13g2_decap_8 FILLER_3_736 ();
 sg13g2_decap_8 FILLER_3_748 ();
 sg13g2_decap_8 FILLER_3_755 ();
 sg13g2_decap_8 FILLER_3_762 ();
 sg13g2_decap_8 FILLER_3_769 ();
 sg13g2_decap_4 FILLER_3_776 ();
 sg13g2_fill_1 FILLER_3_780 ();
 sg13g2_decap_8 FILLER_3_786 ();
 sg13g2_decap_8 FILLER_3_793 ();
 sg13g2_decap_4 FILLER_3_800 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_4 FILLER_3_833 ();
 sg13g2_fill_2 FILLER_3_842 ();
 sg13g2_fill_1 FILLER_3_844 ();
 sg13g2_decap_8 FILLER_3_849 ();
 sg13g2_decap_8 FILLER_3_856 ();
 sg13g2_decap_8 FILLER_3_863 ();
 sg13g2_decap_8 FILLER_3_870 ();
 sg13g2_decap_8 FILLER_3_877 ();
 sg13g2_fill_1 FILLER_3_884 ();
 sg13g2_decap_8 FILLER_3_889 ();
 sg13g2_decap_8 FILLER_3_896 ();
 sg13g2_decap_8 FILLER_3_903 ();
 sg13g2_decap_8 FILLER_3_945 ();
 sg13g2_decap_8 FILLER_3_952 ();
 sg13g2_decap_8 FILLER_3_959 ();
 sg13g2_decap_4 FILLER_3_966 ();
 sg13g2_fill_1 FILLER_3_970 ();
 sg13g2_decap_4 FILLER_3_976 ();
 sg13g2_fill_2 FILLER_3_988 ();
 sg13g2_fill_1 FILLER_3_999 ();
 sg13g2_decap_8 FILLER_3_1007 ();
 sg13g2_decap_4 FILLER_3_1014 ();
 sg13g2_decap_8 FILLER_3_1023 ();
 sg13g2_decap_4 FILLER_3_1030 ();
 sg13g2_fill_2 FILLER_3_1034 ();
 sg13g2_fill_1 FILLER_3_1050 ();
 sg13g2_fill_2 FILLER_3_1056 ();
 sg13g2_fill_1 FILLER_3_1077 ();
 sg13g2_decap_8 FILLER_3_1088 ();
 sg13g2_decap_4 FILLER_3_1095 ();
 sg13g2_fill_2 FILLER_3_1099 ();
 sg13g2_fill_2 FILLER_3_1115 ();
 sg13g2_decap_8 FILLER_3_1146 ();
 sg13g2_decap_8 FILLER_3_1153 ();
 sg13g2_fill_1 FILLER_3_1160 ();
 sg13g2_fill_2 FILLER_3_1172 ();
 sg13g2_decap_8 FILLER_3_1177 ();
 sg13g2_decap_8 FILLER_3_1184 ();
 sg13g2_decap_4 FILLER_3_1191 ();
 sg13g2_fill_2 FILLER_3_1195 ();
 sg13g2_decap_8 FILLER_3_1215 ();
 sg13g2_decap_4 FILLER_3_1222 ();
 sg13g2_fill_2 FILLER_3_1226 ();
 sg13g2_decap_8 FILLER_3_1232 ();
 sg13g2_decap_4 FILLER_3_1239 ();
 sg13g2_fill_2 FILLER_3_1243 ();
 sg13g2_decap_8 FILLER_3_1255 ();
 sg13g2_decap_8 FILLER_3_1262 ();
 sg13g2_decap_8 FILLER_3_1269 ();
 sg13g2_decap_8 FILLER_3_1276 ();
 sg13g2_decap_8 FILLER_3_1283 ();
 sg13g2_decap_8 FILLER_3_1295 ();
 sg13g2_fill_2 FILLER_3_1302 ();
 sg13g2_fill_2 FILLER_3_1312 ();
 sg13g2_fill_1 FILLER_3_1314 ();
 sg13g2_decap_8 FILLER_3_1358 ();
 sg13g2_decap_8 FILLER_3_1365 ();
 sg13g2_decap_8 FILLER_3_1372 ();
 sg13g2_decap_8 FILLER_3_1379 ();
 sg13g2_fill_2 FILLER_3_1386 ();
 sg13g2_fill_1 FILLER_3_1388 ();
 sg13g2_decap_8 FILLER_3_1393 ();
 sg13g2_fill_2 FILLER_3_1400 ();
 sg13g2_fill_1 FILLER_3_1402 ();
 sg13g2_decap_8 FILLER_3_1429 ();
 sg13g2_decap_8 FILLER_3_1436 ();
 sg13g2_decap_8 FILLER_3_1443 ();
 sg13g2_decap_8 FILLER_3_1450 ();
 sg13g2_decap_8 FILLER_3_1457 ();
 sg13g2_decap_8 FILLER_3_1464 ();
 sg13g2_decap_8 FILLER_3_1471 ();
 sg13g2_decap_8 FILLER_3_1478 ();
 sg13g2_decap_8 FILLER_3_1485 ();
 sg13g2_decap_8 FILLER_3_1492 ();
 sg13g2_decap_8 FILLER_3_1499 ();
 sg13g2_decap_8 FILLER_3_1506 ();
 sg13g2_decap_8 FILLER_3_1513 ();
 sg13g2_decap_8 FILLER_3_1520 ();
 sg13g2_decap_8 FILLER_3_1527 ();
 sg13g2_decap_8 FILLER_3_1534 ();
 sg13g2_decap_8 FILLER_3_1541 ();
 sg13g2_decap_8 FILLER_3_1548 ();
 sg13g2_decap_8 FILLER_3_1555 ();
 sg13g2_decap_8 FILLER_3_1562 ();
 sg13g2_decap_8 FILLER_3_1569 ();
 sg13g2_decap_8 FILLER_3_1576 ();
 sg13g2_decap_8 FILLER_3_1583 ();
 sg13g2_decap_8 FILLER_3_1590 ();
 sg13g2_decap_8 FILLER_3_1597 ();
 sg13g2_decap_8 FILLER_3_1604 ();
 sg13g2_decap_8 FILLER_3_1611 ();
 sg13g2_decap_8 FILLER_3_1618 ();
 sg13g2_decap_8 FILLER_3_1625 ();
 sg13g2_decap_8 FILLER_3_1632 ();
 sg13g2_decap_8 FILLER_3_1639 ();
 sg13g2_decap_8 FILLER_3_1646 ();
 sg13g2_decap_8 FILLER_3_1653 ();
 sg13g2_decap_8 FILLER_3_1660 ();
 sg13g2_decap_8 FILLER_3_1667 ();
 sg13g2_decap_8 FILLER_3_1674 ();
 sg13g2_decap_8 FILLER_3_1681 ();
 sg13g2_decap_8 FILLER_3_1688 ();
 sg13g2_decap_8 FILLER_3_1695 ();
 sg13g2_decap_8 FILLER_3_1702 ();
 sg13g2_decap_8 FILLER_3_1709 ();
 sg13g2_decap_8 FILLER_3_1716 ();
 sg13g2_decap_8 FILLER_3_1723 ();
 sg13g2_decap_8 FILLER_3_1730 ();
 sg13g2_decap_8 FILLER_3_1737 ();
 sg13g2_decap_8 FILLER_3_1744 ();
 sg13g2_decap_8 FILLER_3_1751 ();
 sg13g2_decap_8 FILLER_3_1758 ();
 sg13g2_decap_8 FILLER_3_1765 ();
 sg13g2_fill_2 FILLER_3_1772 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_4 FILLER_4_70 ();
 sg13g2_fill_2 FILLER_4_74 ();
 sg13g2_decap_4 FILLER_4_80 ();
 sg13g2_fill_2 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_104 ();
 sg13g2_fill_2 FILLER_4_111 ();
 sg13g2_decap_8 FILLER_4_117 ();
 sg13g2_decap_8 FILLER_4_124 ();
 sg13g2_decap_8 FILLER_4_131 ();
 sg13g2_decap_8 FILLER_4_138 ();
 sg13g2_decap_4 FILLER_4_150 ();
 sg13g2_fill_1 FILLER_4_154 ();
 sg13g2_decap_4 FILLER_4_160 ();
 sg13g2_decap_4 FILLER_4_168 ();
 sg13g2_fill_2 FILLER_4_183 ();
 sg13g2_fill_1 FILLER_4_185 ();
 sg13g2_fill_1 FILLER_4_198 ();
 sg13g2_decap_8 FILLER_4_215 ();
 sg13g2_fill_2 FILLER_4_222 ();
 sg13g2_fill_1 FILLER_4_224 ();
 sg13g2_fill_2 FILLER_4_237 ();
 sg13g2_fill_1 FILLER_4_244 ();
 sg13g2_fill_2 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_fill_2 FILLER_4_285 ();
 sg13g2_fill_2 FILLER_4_296 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_decap_4 FILLER_4_309 ();
 sg13g2_fill_2 FILLER_4_313 ();
 sg13g2_fill_1 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_353 ();
 sg13g2_fill_2 FILLER_4_360 ();
 sg13g2_fill_1 FILLER_4_362 ();
 sg13g2_fill_2 FILLER_4_374 ();
 sg13g2_decap_4 FILLER_4_380 ();
 sg13g2_fill_1 FILLER_4_389 ();
 sg13g2_fill_1 FILLER_4_394 ();
 sg13g2_fill_2 FILLER_4_400 ();
 sg13g2_fill_1 FILLER_4_407 ();
 sg13g2_decap_4 FILLER_4_426 ();
 sg13g2_fill_1 FILLER_4_430 ();
 sg13g2_decap_4 FILLER_4_436 ();
 sg13g2_decap_8 FILLER_4_463 ();
 sg13g2_decap_8 FILLER_4_470 ();
 sg13g2_decap_8 FILLER_4_477 ();
 sg13g2_decap_8 FILLER_4_484 ();
 sg13g2_decap_8 FILLER_4_491 ();
 sg13g2_decap_8 FILLER_4_498 ();
 sg13g2_fill_2 FILLER_4_505 ();
 sg13g2_fill_1 FILLER_4_507 ();
 sg13g2_decap_8 FILLER_4_512 ();
 sg13g2_decap_8 FILLER_4_519 ();
 sg13g2_decap_8 FILLER_4_526 ();
 sg13g2_decap_4 FILLER_4_533 ();
 sg13g2_fill_2 FILLER_4_537 ();
 sg13g2_decap_8 FILLER_4_543 ();
 sg13g2_decap_8 FILLER_4_550 ();
 sg13g2_decap_8 FILLER_4_561 ();
 sg13g2_decap_8 FILLER_4_568 ();
 sg13g2_decap_8 FILLER_4_575 ();
 sg13g2_decap_8 FILLER_4_582 ();
 sg13g2_decap_4 FILLER_4_589 ();
 sg13g2_decap_8 FILLER_4_597 ();
 sg13g2_decap_8 FILLER_4_604 ();
 sg13g2_decap_8 FILLER_4_611 ();
 sg13g2_decap_8 FILLER_4_618 ();
 sg13g2_decap_4 FILLER_4_625 ();
 sg13g2_fill_1 FILLER_4_629 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_4 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_676 ();
 sg13g2_fill_2 FILLER_4_683 ();
 sg13g2_fill_1 FILLER_4_685 ();
 sg13g2_decap_8 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_697 ();
 sg13g2_decap_8 FILLER_4_704 ();
 sg13g2_decap_4 FILLER_4_737 ();
 sg13g2_fill_2 FILLER_4_741 ();
 sg13g2_decap_4 FILLER_4_786 ();
 sg13g2_fill_2 FILLER_4_790 ();
 sg13g2_decap_8 FILLER_4_796 ();
 sg13g2_decap_4 FILLER_4_803 ();
 sg13g2_fill_1 FILLER_4_807 ();
 sg13g2_decap_8 FILLER_4_820 ();
 sg13g2_decap_8 FILLER_4_827 ();
 sg13g2_decap_4 FILLER_4_834 ();
 sg13g2_decap_8 FILLER_4_864 ();
 sg13g2_decap_8 FILLER_4_871 ();
 sg13g2_fill_1 FILLER_4_904 ();
 sg13g2_fill_2 FILLER_4_937 ();
 sg13g2_fill_1 FILLER_4_939 ();
 sg13g2_decap_8 FILLER_4_944 ();
 sg13g2_fill_1 FILLER_4_951 ();
 sg13g2_decap_8 FILLER_4_978 ();
 sg13g2_decap_8 FILLER_4_985 ();
 sg13g2_decap_4 FILLER_4_992 ();
 sg13g2_fill_2 FILLER_4_996 ();
 sg13g2_decap_8 FILLER_4_1013 ();
 sg13g2_decap_4 FILLER_4_1020 ();
 sg13g2_fill_2 FILLER_4_1036 ();
 sg13g2_fill_1 FILLER_4_1038 ();
 sg13g2_fill_2 FILLER_4_1047 ();
 sg13g2_decap_8 FILLER_4_1053 ();
 sg13g2_decap_4 FILLER_4_1060 ();
 sg13g2_fill_1 FILLER_4_1064 ();
 sg13g2_decap_8 FILLER_4_1071 ();
 sg13g2_fill_2 FILLER_4_1078 ();
 sg13g2_fill_1 FILLER_4_1080 ();
 sg13g2_fill_1 FILLER_4_1092 ();
 sg13g2_decap_8 FILLER_4_1097 ();
 sg13g2_decap_8 FILLER_4_1104 ();
 sg13g2_decap_8 FILLER_4_1111 ();
 sg13g2_fill_1 FILLER_4_1118 ();
 sg13g2_decap_4 FILLER_4_1159 ();
 sg13g2_fill_2 FILLER_4_1163 ();
 sg13g2_decap_4 FILLER_4_1169 ();
 sg13g2_fill_1 FILLER_4_1173 ();
 sg13g2_fill_2 FILLER_4_1179 ();
 sg13g2_fill_1 FILLER_4_1181 ();
 sg13g2_fill_2 FILLER_4_1214 ();
 sg13g2_decap_8 FILLER_4_1247 ();
 sg13g2_decap_8 FILLER_4_1254 ();
 sg13g2_decap_8 FILLER_4_1261 ();
 sg13g2_decap_8 FILLER_4_1298 ();
 sg13g2_decap_8 FILLER_4_1305 ();
 sg13g2_decap_8 FILLER_4_1312 ();
 sg13g2_fill_2 FILLER_4_1319 ();
 sg13g2_decap_8 FILLER_4_1326 ();
 sg13g2_decap_8 FILLER_4_1333 ();
 sg13g2_decap_8 FILLER_4_1340 ();
 sg13g2_fill_1 FILLER_4_1347 ();
 sg13g2_decap_8 FILLER_4_1362 ();
 sg13g2_decap_8 FILLER_4_1369 ();
 sg13g2_decap_4 FILLER_4_1402 ();
 sg13g2_fill_2 FILLER_4_1429 ();
 sg13g2_fill_1 FILLER_4_1431 ();
 sg13g2_decap_8 FILLER_4_1436 ();
 sg13g2_decap_8 FILLER_4_1443 ();
 sg13g2_decap_8 FILLER_4_1450 ();
 sg13g2_decap_8 FILLER_4_1457 ();
 sg13g2_decap_8 FILLER_4_1464 ();
 sg13g2_decap_8 FILLER_4_1471 ();
 sg13g2_decap_8 FILLER_4_1478 ();
 sg13g2_decap_8 FILLER_4_1485 ();
 sg13g2_decap_8 FILLER_4_1492 ();
 sg13g2_decap_8 FILLER_4_1499 ();
 sg13g2_decap_8 FILLER_4_1506 ();
 sg13g2_decap_8 FILLER_4_1513 ();
 sg13g2_decap_8 FILLER_4_1520 ();
 sg13g2_decap_8 FILLER_4_1527 ();
 sg13g2_decap_8 FILLER_4_1534 ();
 sg13g2_decap_8 FILLER_4_1541 ();
 sg13g2_decap_8 FILLER_4_1548 ();
 sg13g2_decap_8 FILLER_4_1555 ();
 sg13g2_decap_8 FILLER_4_1562 ();
 sg13g2_decap_8 FILLER_4_1569 ();
 sg13g2_decap_8 FILLER_4_1576 ();
 sg13g2_decap_8 FILLER_4_1583 ();
 sg13g2_decap_8 FILLER_4_1590 ();
 sg13g2_decap_8 FILLER_4_1597 ();
 sg13g2_decap_8 FILLER_4_1604 ();
 sg13g2_decap_8 FILLER_4_1611 ();
 sg13g2_decap_8 FILLER_4_1618 ();
 sg13g2_decap_8 FILLER_4_1625 ();
 sg13g2_decap_8 FILLER_4_1632 ();
 sg13g2_decap_8 FILLER_4_1639 ();
 sg13g2_decap_8 FILLER_4_1646 ();
 sg13g2_decap_8 FILLER_4_1653 ();
 sg13g2_decap_8 FILLER_4_1660 ();
 sg13g2_decap_8 FILLER_4_1667 ();
 sg13g2_decap_8 FILLER_4_1674 ();
 sg13g2_decap_8 FILLER_4_1681 ();
 sg13g2_decap_8 FILLER_4_1688 ();
 sg13g2_decap_8 FILLER_4_1695 ();
 sg13g2_decap_8 FILLER_4_1702 ();
 sg13g2_decap_8 FILLER_4_1709 ();
 sg13g2_decap_8 FILLER_4_1716 ();
 sg13g2_decap_8 FILLER_4_1723 ();
 sg13g2_decap_8 FILLER_4_1730 ();
 sg13g2_decap_8 FILLER_4_1737 ();
 sg13g2_decap_8 FILLER_4_1744 ();
 sg13g2_decap_8 FILLER_4_1751 ();
 sg13g2_decap_8 FILLER_4_1758 ();
 sg13g2_decap_8 FILLER_4_1765 ();
 sg13g2_fill_2 FILLER_4_1772 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_fill_1 FILLER_5_49 ();
 sg13g2_decap_4 FILLER_5_59 ();
 sg13g2_fill_1 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_73 ();
 sg13g2_fill_1 FILLER_5_80 ();
 sg13g2_fill_2 FILLER_5_89 ();
 sg13g2_fill_1 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_4 FILLER_5_109 ();
 sg13g2_fill_1 FILLER_5_113 ();
 sg13g2_fill_1 FILLER_5_119 ();
 sg13g2_decap_4 FILLER_5_124 ();
 sg13g2_decap_4 FILLER_5_133 ();
 sg13g2_decap_4 FILLER_5_143 ();
 sg13g2_fill_2 FILLER_5_151 ();
 sg13g2_fill_1 FILLER_5_153 ();
 sg13g2_fill_2 FILLER_5_163 ();
 sg13g2_decap_8 FILLER_5_170 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_192 ();
 sg13g2_decap_8 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_5_206 ();
 sg13g2_decap_4 FILLER_5_213 ();
 sg13g2_fill_2 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_4 FILLER_5_245 ();
 sg13g2_fill_2 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_8 FILLER_5_293 ();
 sg13g2_decap_4 FILLER_5_300 ();
 sg13g2_fill_1 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_fill_1 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_4 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_fill_2 FILLER_5_384 ();
 sg13g2_fill_1 FILLER_5_391 ();
 sg13g2_decap_4 FILLER_5_397 ();
 sg13g2_fill_1 FILLER_5_401 ();
 sg13g2_fill_2 FILLER_5_412 ();
 sg13g2_decap_8 FILLER_5_419 ();
 sg13g2_decap_8 FILLER_5_426 ();
 sg13g2_decap_8 FILLER_5_433 ();
 sg13g2_fill_1 FILLER_5_440 ();
 sg13g2_decap_8 FILLER_5_447 ();
 sg13g2_decap_8 FILLER_5_454 ();
 sg13g2_fill_2 FILLER_5_461 ();
 sg13g2_fill_1 FILLER_5_463 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_fill_2 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_533 ();
 sg13g2_decap_8 FILLER_5_540 ();
 sg13g2_fill_2 FILLER_5_551 ();
 sg13g2_fill_1 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_558 ();
 sg13g2_decap_8 FILLER_5_565 ();
 sg13g2_decap_8 FILLER_5_572 ();
 sg13g2_fill_2 FILLER_5_579 ();
 sg13g2_decap_4 FILLER_5_620 ();
 sg13g2_fill_1 FILLER_5_624 ();
 sg13g2_decap_8 FILLER_5_633 ();
 sg13g2_fill_2 FILLER_5_640 ();
 sg13g2_fill_1 FILLER_5_642 ();
 sg13g2_fill_1 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_653 ();
 sg13g2_decap_4 FILLER_5_660 ();
 sg13g2_fill_2 FILLER_5_664 ();
 sg13g2_decap_4 FILLER_5_675 ();
 sg13g2_fill_1 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_706 ();
 sg13g2_fill_2 FILLER_5_713 ();
 sg13g2_fill_1 FILLER_5_715 ();
 sg13g2_decap_4 FILLER_5_720 ();
 sg13g2_fill_1 FILLER_5_724 ();
 sg13g2_decap_8 FILLER_5_729 ();
 sg13g2_decap_8 FILLER_5_736 ();
 sg13g2_decap_8 FILLER_5_751 ();
 sg13g2_decap_8 FILLER_5_758 ();
 sg13g2_decap_4 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_773 ();
 sg13g2_decap_4 FILLER_5_780 ();
 sg13g2_fill_1 FILLER_5_784 ();
 sg13g2_fill_2 FILLER_5_811 ();
 sg13g2_decap_8 FILLER_5_818 ();
 sg13g2_decap_8 FILLER_5_825 ();
 sg13g2_decap_8 FILLER_5_832 ();
 sg13g2_decap_8 FILLER_5_839 ();
 sg13g2_fill_2 FILLER_5_846 ();
 sg13g2_decap_8 FILLER_5_852 ();
 sg13g2_decap_8 FILLER_5_859 ();
 sg13g2_decap_8 FILLER_5_866 ();
 sg13g2_decap_8 FILLER_5_873 ();
 sg13g2_fill_1 FILLER_5_880 ();
 sg13g2_decap_8 FILLER_5_889 ();
 sg13g2_decap_4 FILLER_5_896 ();
 sg13g2_decap_8 FILLER_5_904 ();
 sg13g2_fill_2 FILLER_5_911 ();
 sg13g2_decap_8 FILLER_5_917 ();
 sg13g2_decap_8 FILLER_5_924 ();
 sg13g2_decap_8 FILLER_5_931 ();
 sg13g2_decap_8 FILLER_5_938 ();
 sg13g2_fill_2 FILLER_5_945 ();
 sg13g2_decap_4 FILLER_5_955 ();
 sg13g2_fill_1 FILLER_5_959 ();
 sg13g2_decap_8 FILLER_5_964 ();
 sg13g2_fill_1 FILLER_5_971 ();
 sg13g2_decap_8 FILLER_5_976 ();
 sg13g2_decap_8 FILLER_5_983 ();
 sg13g2_decap_8 FILLER_5_990 ();
 sg13g2_decap_4 FILLER_5_997 ();
 sg13g2_decap_8 FILLER_5_1006 ();
 sg13g2_decap_8 FILLER_5_1013 ();
 sg13g2_decap_8 FILLER_5_1020 ();
 sg13g2_decap_8 FILLER_5_1027 ();
 sg13g2_decap_4 FILLER_5_1034 ();
 sg13g2_fill_1 FILLER_5_1038 ();
 sg13g2_decap_4 FILLER_5_1054 ();
 sg13g2_fill_1 FILLER_5_1058 ();
 sg13g2_decap_8 FILLER_5_1064 ();
 sg13g2_decap_8 FILLER_5_1071 ();
 sg13g2_decap_8 FILLER_5_1078 ();
 sg13g2_fill_2 FILLER_5_1090 ();
 sg13g2_fill_1 FILLER_5_1092 ();
 sg13g2_decap_4 FILLER_5_1101 ();
 sg13g2_fill_2 FILLER_5_1105 ();
 sg13g2_decap_8 FILLER_5_1110 ();
 sg13g2_decap_8 FILLER_5_1148 ();
 sg13g2_decap_8 FILLER_5_1155 ();
 sg13g2_decap_8 FILLER_5_1162 ();
 sg13g2_decap_4 FILLER_5_1169 ();
 sg13g2_decap_4 FILLER_5_1181 ();
 sg13g2_fill_2 FILLER_5_1185 ();
 sg13g2_decap_4 FILLER_5_1192 ();
 sg13g2_fill_1 FILLER_5_1196 ();
 sg13g2_decap_8 FILLER_5_1201 ();
 sg13g2_decap_4 FILLER_5_1208 ();
 sg13g2_fill_1 FILLER_5_1212 ();
 sg13g2_decap_4 FILLER_5_1218 ();
 sg13g2_fill_1 FILLER_5_1222 ();
 sg13g2_decap_8 FILLER_5_1228 ();
 sg13g2_decap_8 FILLER_5_1235 ();
 sg13g2_decap_8 FILLER_5_1242 ();
 sg13g2_decap_8 FILLER_5_1249 ();
 sg13g2_decap_8 FILLER_5_1256 ();
 sg13g2_decap_4 FILLER_5_1263 ();
 sg13g2_fill_1 FILLER_5_1267 ();
 sg13g2_decap_8 FILLER_5_1276 ();
 sg13g2_decap_8 FILLER_5_1283 ();
 sg13g2_fill_1 FILLER_5_1290 ();
 sg13g2_decap_8 FILLER_5_1295 ();
 sg13g2_decap_8 FILLER_5_1302 ();
 sg13g2_decap_8 FILLER_5_1313 ();
 sg13g2_fill_2 FILLER_5_1320 ();
 sg13g2_fill_1 FILLER_5_1322 ();
 sg13g2_decap_8 FILLER_5_1328 ();
 sg13g2_decap_8 FILLER_5_1335 ();
 sg13g2_fill_2 FILLER_5_1342 ();
 sg13g2_decap_8 FILLER_5_1359 ();
 sg13g2_decap_4 FILLER_5_1366 ();
 sg13g2_fill_1 FILLER_5_1370 ();
 sg13g2_decap_4 FILLER_5_1376 ();
 sg13g2_fill_1 FILLER_5_1380 ();
 sg13g2_decap_4 FILLER_5_1402 ();
 sg13g2_fill_1 FILLER_5_1424 ();
 sg13g2_decap_8 FILLER_5_1456 ();
 sg13g2_decap_8 FILLER_5_1463 ();
 sg13g2_decap_8 FILLER_5_1470 ();
 sg13g2_decap_8 FILLER_5_1477 ();
 sg13g2_decap_8 FILLER_5_1484 ();
 sg13g2_decap_8 FILLER_5_1491 ();
 sg13g2_decap_8 FILLER_5_1498 ();
 sg13g2_decap_8 FILLER_5_1505 ();
 sg13g2_decap_8 FILLER_5_1512 ();
 sg13g2_decap_8 FILLER_5_1519 ();
 sg13g2_decap_8 FILLER_5_1526 ();
 sg13g2_decap_8 FILLER_5_1533 ();
 sg13g2_decap_8 FILLER_5_1540 ();
 sg13g2_decap_8 FILLER_5_1547 ();
 sg13g2_decap_8 FILLER_5_1554 ();
 sg13g2_decap_8 FILLER_5_1561 ();
 sg13g2_decap_8 FILLER_5_1568 ();
 sg13g2_decap_8 FILLER_5_1575 ();
 sg13g2_decap_8 FILLER_5_1582 ();
 sg13g2_decap_8 FILLER_5_1589 ();
 sg13g2_decap_8 FILLER_5_1596 ();
 sg13g2_decap_8 FILLER_5_1603 ();
 sg13g2_decap_8 FILLER_5_1610 ();
 sg13g2_decap_8 FILLER_5_1617 ();
 sg13g2_decap_8 FILLER_5_1624 ();
 sg13g2_decap_8 FILLER_5_1631 ();
 sg13g2_decap_8 FILLER_5_1638 ();
 sg13g2_decap_8 FILLER_5_1645 ();
 sg13g2_decap_8 FILLER_5_1652 ();
 sg13g2_decap_8 FILLER_5_1659 ();
 sg13g2_decap_8 FILLER_5_1666 ();
 sg13g2_decap_8 FILLER_5_1673 ();
 sg13g2_decap_8 FILLER_5_1680 ();
 sg13g2_decap_8 FILLER_5_1687 ();
 sg13g2_decap_8 FILLER_5_1694 ();
 sg13g2_decap_8 FILLER_5_1701 ();
 sg13g2_decap_8 FILLER_5_1708 ();
 sg13g2_decap_8 FILLER_5_1715 ();
 sg13g2_decap_8 FILLER_5_1722 ();
 sg13g2_decap_8 FILLER_5_1729 ();
 sg13g2_decap_8 FILLER_5_1736 ();
 sg13g2_decap_8 FILLER_5_1743 ();
 sg13g2_decap_8 FILLER_5_1750 ();
 sg13g2_decap_8 FILLER_5_1757 ();
 sg13g2_decap_8 FILLER_5_1764 ();
 sg13g2_fill_2 FILLER_5_1771 ();
 sg13g2_fill_1 FILLER_5_1773 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_fill_2 FILLER_6_53 ();
 sg13g2_fill_1 FILLER_6_55 ();
 sg13g2_decap_4 FILLER_6_61 ();
 sg13g2_fill_1 FILLER_6_65 ();
 sg13g2_fill_2 FILLER_6_75 ();
 sg13g2_decap_8 FILLER_6_86 ();
 sg13g2_fill_2 FILLER_6_93 ();
 sg13g2_decap_8 FILLER_6_99 ();
 sg13g2_fill_1 FILLER_6_106 ();
 sg13g2_fill_2 FILLER_6_117 ();
 sg13g2_fill_1 FILLER_6_128 ();
 sg13g2_fill_2 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_decap_4 FILLER_6_153 ();
 sg13g2_decap_8 FILLER_6_162 ();
 sg13g2_decap_8 FILLER_6_169 ();
 sg13g2_fill_1 FILLER_6_176 ();
 sg13g2_fill_1 FILLER_6_195 ();
 sg13g2_decap_4 FILLER_6_209 ();
 sg13g2_fill_2 FILLER_6_213 ();
 sg13g2_fill_1 FILLER_6_233 ();
 sg13g2_decap_4 FILLER_6_239 ();
 sg13g2_fill_2 FILLER_6_243 ();
 sg13g2_fill_1 FILLER_6_254 ();
 sg13g2_decap_8 FILLER_6_265 ();
 sg13g2_decap_8 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_279 ();
 sg13g2_decap_8 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_293 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_fill_2 FILLER_6_319 ();
 sg13g2_decap_4 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_fill_2 FILLER_6_379 ();
 sg13g2_decap_4 FILLER_6_389 ();
 sg13g2_fill_2 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_fill_2 FILLER_6_424 ();
 sg13g2_fill_1 FILLER_6_426 ();
 sg13g2_decap_4 FILLER_6_435 ();
 sg13g2_fill_2 FILLER_6_439 ();
 sg13g2_decap_8 FILLER_6_449 ();
 sg13g2_fill_1 FILLER_6_456 ();
 sg13g2_decap_8 FILLER_6_465 ();
 sg13g2_decap_8 FILLER_6_472 ();
 sg13g2_fill_1 FILLER_6_479 ();
 sg13g2_decap_8 FILLER_6_484 ();
 sg13g2_decap_8 FILLER_6_491 ();
 sg13g2_decap_8 FILLER_6_498 ();
 sg13g2_decap_8 FILLER_6_505 ();
 sg13g2_decap_8 FILLER_6_512 ();
 sg13g2_decap_8 FILLER_6_519 ();
 sg13g2_decap_8 FILLER_6_526 ();
 sg13g2_fill_2 FILLER_6_543 ();
 sg13g2_decap_8 FILLER_6_575 ();
 sg13g2_decap_8 FILLER_6_582 ();
 sg13g2_decap_8 FILLER_6_589 ();
 sg13g2_decap_8 FILLER_6_596 ();
 sg13g2_decap_8 FILLER_6_603 ();
 sg13g2_decap_8 FILLER_6_610 ();
 sg13g2_decap_8 FILLER_6_617 ();
 sg13g2_fill_2 FILLER_6_624 ();
 sg13g2_fill_1 FILLER_6_626 ();
 sg13g2_fill_2 FILLER_6_632 ();
 sg13g2_fill_2 FILLER_6_639 ();
 sg13g2_decap_8 FILLER_6_667 ();
 sg13g2_decap_8 FILLER_6_674 ();
 sg13g2_decap_8 FILLER_6_681 ();
 sg13g2_fill_1 FILLER_6_688 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_fill_1 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_730 ();
 sg13g2_decap_8 FILLER_6_737 ();
 sg13g2_decap_8 FILLER_6_744 ();
 sg13g2_decap_8 FILLER_6_751 ();
 sg13g2_decap_8 FILLER_6_758 ();
 sg13g2_decap_8 FILLER_6_769 ();
 sg13g2_decap_8 FILLER_6_776 ();
 sg13g2_decap_8 FILLER_6_783 ();
 sg13g2_decap_8 FILLER_6_790 ();
 sg13g2_decap_8 FILLER_6_797 ();
 sg13g2_decap_8 FILLER_6_804 ();
 sg13g2_decap_8 FILLER_6_811 ();
 sg13g2_decap_8 FILLER_6_818 ();
 sg13g2_decap_8 FILLER_6_825 ();
 sg13g2_decap_8 FILLER_6_832 ();
 sg13g2_fill_2 FILLER_6_839 ();
 sg13g2_decap_4 FILLER_6_867 ();
 sg13g2_decap_8 FILLER_6_875 ();
 sg13g2_decap_8 FILLER_6_891 ();
 sg13g2_decap_4 FILLER_6_898 ();
 sg13g2_decap_8 FILLER_6_906 ();
 sg13g2_fill_1 FILLER_6_918 ();
 sg13g2_fill_2 FILLER_6_927 ();
 sg13g2_decap_4 FILLER_6_937 ();
 sg13g2_fill_2 FILLER_6_941 ();
 sg13g2_decap_4 FILLER_6_952 ();
 sg13g2_fill_1 FILLER_6_956 ();
 sg13g2_fill_1 FILLER_6_966 ();
 sg13g2_decap_8 FILLER_6_980 ();
 sg13g2_decap_8 FILLER_6_987 ();
 sg13g2_decap_4 FILLER_6_994 ();
 sg13g2_fill_2 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_4 FILLER_6_1019 ();
 sg13g2_fill_1 FILLER_6_1023 ();
 sg13g2_decap_8 FILLER_6_1028 ();
 sg13g2_decap_8 FILLER_6_1035 ();
 sg13g2_decap_8 FILLER_6_1042 ();
 sg13g2_fill_1 FILLER_6_1049 ();
 sg13g2_decap_8 FILLER_6_1055 ();
 sg13g2_decap_4 FILLER_6_1062 ();
 sg13g2_decap_8 FILLER_6_1071 ();
 sg13g2_fill_2 FILLER_6_1078 ();
 sg13g2_fill_1 FILLER_6_1080 ();
 sg13g2_decap_8 FILLER_6_1086 ();
 sg13g2_fill_1 FILLER_6_1093 ();
 sg13g2_decap_4 FILLER_6_1130 ();
 sg13g2_decap_8 FILLER_6_1164 ();
 sg13g2_fill_2 FILLER_6_1179 ();
 sg13g2_fill_1 FILLER_6_1181 ();
 sg13g2_fill_2 FILLER_6_1199 ();
 sg13g2_decap_8 FILLER_6_1205 ();
 sg13g2_fill_1 FILLER_6_1212 ();
 sg13g2_fill_2 FILLER_6_1242 ();
 sg13g2_decap_4 FILLER_6_1256 ();
 sg13g2_fill_2 FILLER_6_1260 ();
 sg13g2_decap_8 FILLER_6_1266 ();
 sg13g2_decap_8 FILLER_6_1273 ();
 sg13g2_decap_8 FILLER_6_1280 ();
 sg13g2_decap_8 FILLER_6_1287 ();
 sg13g2_decap_8 FILLER_6_1294 ();
 sg13g2_fill_1 FILLER_6_1301 ();
 sg13g2_decap_8 FILLER_6_1328 ();
 sg13g2_decap_8 FILLER_6_1335 ();
 sg13g2_decap_8 FILLER_6_1342 ();
 sg13g2_decap_8 FILLER_6_1349 ();
 sg13g2_fill_2 FILLER_6_1368 ();
 sg13g2_fill_1 FILLER_6_1374 ();
 sg13g2_decap_4 FILLER_6_1380 ();
 sg13g2_fill_1 FILLER_6_1384 ();
 sg13g2_fill_1 FILLER_6_1398 ();
 sg13g2_decap_8 FILLER_6_1422 ();
 sg13g2_decap_8 FILLER_6_1429 ();
 sg13g2_decap_8 FILLER_6_1436 ();
 sg13g2_decap_8 FILLER_6_1443 ();
 sg13g2_decap_8 FILLER_6_1450 ();
 sg13g2_decap_8 FILLER_6_1457 ();
 sg13g2_decap_8 FILLER_6_1464 ();
 sg13g2_decap_8 FILLER_6_1471 ();
 sg13g2_decap_8 FILLER_6_1478 ();
 sg13g2_decap_8 FILLER_6_1485 ();
 sg13g2_decap_8 FILLER_6_1492 ();
 sg13g2_decap_8 FILLER_6_1499 ();
 sg13g2_decap_8 FILLER_6_1506 ();
 sg13g2_decap_8 FILLER_6_1513 ();
 sg13g2_decap_8 FILLER_6_1520 ();
 sg13g2_decap_8 FILLER_6_1527 ();
 sg13g2_decap_8 FILLER_6_1534 ();
 sg13g2_decap_8 FILLER_6_1541 ();
 sg13g2_decap_8 FILLER_6_1548 ();
 sg13g2_decap_8 FILLER_6_1555 ();
 sg13g2_decap_8 FILLER_6_1562 ();
 sg13g2_decap_8 FILLER_6_1569 ();
 sg13g2_decap_8 FILLER_6_1576 ();
 sg13g2_decap_8 FILLER_6_1583 ();
 sg13g2_decap_8 FILLER_6_1590 ();
 sg13g2_decap_8 FILLER_6_1597 ();
 sg13g2_decap_8 FILLER_6_1604 ();
 sg13g2_decap_8 FILLER_6_1611 ();
 sg13g2_decap_8 FILLER_6_1618 ();
 sg13g2_decap_8 FILLER_6_1625 ();
 sg13g2_decap_8 FILLER_6_1632 ();
 sg13g2_decap_8 FILLER_6_1639 ();
 sg13g2_decap_8 FILLER_6_1646 ();
 sg13g2_decap_8 FILLER_6_1653 ();
 sg13g2_decap_8 FILLER_6_1660 ();
 sg13g2_decap_8 FILLER_6_1667 ();
 sg13g2_decap_8 FILLER_6_1674 ();
 sg13g2_decap_8 FILLER_6_1681 ();
 sg13g2_decap_8 FILLER_6_1688 ();
 sg13g2_decap_8 FILLER_6_1695 ();
 sg13g2_decap_8 FILLER_6_1702 ();
 sg13g2_decap_8 FILLER_6_1709 ();
 sg13g2_decap_8 FILLER_6_1716 ();
 sg13g2_decap_8 FILLER_6_1723 ();
 sg13g2_decap_8 FILLER_6_1730 ();
 sg13g2_decap_8 FILLER_6_1737 ();
 sg13g2_decap_8 FILLER_6_1744 ();
 sg13g2_decap_8 FILLER_6_1751 ();
 sg13g2_decap_8 FILLER_6_1758 ();
 sg13g2_decap_8 FILLER_6_1765 ();
 sg13g2_fill_2 FILLER_6_1772 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_4 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_44 ();
 sg13g2_fill_1 FILLER_7_70 ();
 sg13g2_decap_4 FILLER_7_85 ();
 sg13g2_fill_1 FILLER_7_89 ();
 sg13g2_fill_1 FILLER_7_95 ();
 sg13g2_decap_4 FILLER_7_106 ();
 sg13g2_fill_2 FILLER_7_110 ();
 sg13g2_decap_4 FILLER_7_117 ();
 sg13g2_fill_2 FILLER_7_121 ();
 sg13g2_decap_8 FILLER_7_128 ();
 sg13g2_decap_8 FILLER_7_135 ();
 sg13g2_fill_2 FILLER_7_142 ();
 sg13g2_fill_1 FILLER_7_144 ();
 sg13g2_decap_8 FILLER_7_158 ();
 sg13g2_decap_4 FILLER_7_165 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_decap_4 FILLER_7_176 ();
 sg13g2_fill_1 FILLER_7_180 ();
 sg13g2_fill_2 FILLER_7_191 ();
 sg13g2_fill_1 FILLER_7_193 ();
 sg13g2_decap_4 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_207 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_fill_1 FILLER_7_232 ();
 sg13g2_decap_4 FILLER_7_239 ();
 sg13g2_decap_8 FILLER_7_263 ();
 sg13g2_decap_8 FILLER_7_270 ();
 sg13g2_decap_8 FILLER_7_277 ();
 sg13g2_decap_8 FILLER_7_284 ();
 sg13g2_decap_8 FILLER_7_291 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_fill_1 FILLER_7_312 ();
 sg13g2_fill_2 FILLER_7_318 ();
 sg13g2_fill_2 FILLER_7_328 ();
 sg13g2_decap_4 FILLER_7_334 ();
 sg13g2_fill_2 FILLER_7_342 ();
 sg13g2_fill_1 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_fill_1 FILLER_7_357 ();
 sg13g2_fill_1 FILLER_7_363 ();
 sg13g2_fill_2 FILLER_7_368 ();
 sg13g2_fill_2 FILLER_7_375 ();
 sg13g2_fill_1 FILLER_7_377 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_fill_1 FILLER_7_390 ();
 sg13g2_decap_4 FILLER_7_401 ();
 sg13g2_fill_2 FILLER_7_405 ();
 sg13g2_decap_4 FILLER_7_412 ();
 sg13g2_fill_1 FILLER_7_416 ();
 sg13g2_fill_2 FILLER_7_423 ();
 sg13g2_fill_1 FILLER_7_425 ();
 sg13g2_decap_4 FILLER_7_429 ();
 sg13g2_fill_1 FILLER_7_433 ();
 sg13g2_fill_2 FILLER_7_458 ();
 sg13g2_fill_1 FILLER_7_470 ();
 sg13g2_decap_8 FILLER_7_475 ();
 sg13g2_decap_4 FILLER_7_482 ();
 sg13g2_decap_8 FILLER_7_491 ();
 sg13g2_decap_8 FILLER_7_498 ();
 sg13g2_decap_8 FILLER_7_505 ();
 sg13g2_decap_8 FILLER_7_512 ();
 sg13g2_decap_8 FILLER_7_519 ();
 sg13g2_decap_8 FILLER_7_526 ();
 sg13g2_decap_8 FILLER_7_533 ();
 sg13g2_fill_1 FILLER_7_540 ();
 sg13g2_decap_4 FILLER_7_590 ();
 sg13g2_fill_1 FILLER_7_594 ();
 sg13g2_fill_2 FILLER_7_599 ();
 sg13g2_decap_8 FILLER_7_636 ();
 sg13g2_fill_1 FILLER_7_643 ();
 sg13g2_decap_8 FILLER_7_661 ();
 sg13g2_decap_8 FILLER_7_668 ();
 sg13g2_decap_8 FILLER_7_675 ();
 sg13g2_decap_8 FILLER_7_711 ();
 sg13g2_fill_2 FILLER_7_718 ();
 sg13g2_fill_1 FILLER_7_720 ();
 sg13g2_fill_1 FILLER_7_726 ();
 sg13g2_decap_8 FILLER_7_731 ();
 sg13g2_fill_2 FILLER_7_738 ();
 sg13g2_fill_1 FILLER_7_740 ();
 sg13g2_decap_8 FILLER_7_745 ();
 sg13g2_decap_4 FILLER_7_752 ();
 sg13g2_fill_2 FILLER_7_756 ();
 sg13g2_fill_1 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_790 ();
 sg13g2_decap_8 FILLER_7_797 ();
 sg13g2_decap_8 FILLER_7_804 ();
 sg13g2_fill_1 FILLER_7_811 ();
 sg13g2_fill_1 FILLER_7_824 ();
 sg13g2_decap_8 FILLER_7_829 ();
 sg13g2_fill_2 FILLER_7_836 ();
 sg13g2_fill_1 FILLER_7_838 ();
 sg13g2_decap_8 FILLER_7_844 ();
 sg13g2_decap_8 FILLER_7_851 ();
 sg13g2_decap_8 FILLER_7_858 ();
 sg13g2_decap_8 FILLER_7_869 ();
 sg13g2_decap_4 FILLER_7_876 ();
 sg13g2_decap_8 FILLER_7_888 ();
 sg13g2_decap_4 FILLER_7_895 ();
 sg13g2_fill_1 FILLER_7_899 ();
 sg13g2_decap_8 FILLER_7_904 ();
 sg13g2_decap_8 FILLER_7_919 ();
 sg13g2_decap_8 FILLER_7_926 ();
 sg13g2_decap_8 FILLER_7_933 ();
 sg13g2_decap_8 FILLER_7_940 ();
 sg13g2_decap_8 FILLER_7_947 ();
 sg13g2_decap_8 FILLER_7_954 ();
 sg13g2_decap_8 FILLER_7_992 ();
 sg13g2_fill_2 FILLER_7_999 ();
 sg13g2_decap_8 FILLER_7_1027 ();
 sg13g2_fill_2 FILLER_7_1034 ();
 sg13g2_fill_2 FILLER_7_1050 ();
 sg13g2_decap_4 FILLER_7_1058 ();
 sg13g2_fill_1 FILLER_7_1062 ();
 sg13g2_decap_8 FILLER_7_1067 ();
 sg13g2_fill_1 FILLER_7_1079 ();
 sg13g2_decap_8 FILLER_7_1084 ();
 sg13g2_fill_2 FILLER_7_1091 ();
 sg13g2_fill_1 FILLER_7_1093 ();
 sg13g2_fill_2 FILLER_7_1099 ();
 sg13g2_decap_8 FILLER_7_1136 ();
 sg13g2_decap_8 FILLER_7_1143 ();
 sg13g2_decap_8 FILLER_7_1150 ();
 sg13g2_decap_8 FILLER_7_1157 ();
 sg13g2_decap_8 FILLER_7_1164 ();
 sg13g2_decap_8 FILLER_7_1171 ();
 sg13g2_fill_1 FILLER_7_1178 ();
 sg13g2_fill_2 FILLER_7_1193 ();
 sg13g2_fill_1 FILLER_7_1195 ();
 sg13g2_decap_8 FILLER_7_1201 ();
 sg13g2_decap_8 FILLER_7_1208 ();
 sg13g2_decap_8 FILLER_7_1215 ();
 sg13g2_decap_8 FILLER_7_1222 ();
 sg13g2_decap_8 FILLER_7_1229 ();
 sg13g2_decap_8 FILLER_7_1236 ();
 sg13g2_decap_8 FILLER_7_1243 ();
 sg13g2_decap_8 FILLER_7_1281 ();
 sg13g2_decap_8 FILLER_7_1288 ();
 sg13g2_decap_4 FILLER_7_1295 ();
 sg13g2_decap_8 FILLER_7_1315 ();
 sg13g2_decap_8 FILLER_7_1322 ();
 sg13g2_decap_4 FILLER_7_1329 ();
 sg13g2_fill_1 FILLER_7_1333 ();
 sg13g2_decap_8 FILLER_7_1342 ();
 sg13g2_fill_1 FILLER_7_1349 ();
 sg13g2_decap_8 FILLER_7_1361 ();
 sg13g2_fill_2 FILLER_7_1368 ();
 sg13g2_fill_1 FILLER_7_1370 ();
 sg13g2_fill_2 FILLER_7_1374 ();
 sg13g2_fill_1 FILLER_7_1376 ();
 sg13g2_fill_2 FILLER_7_1396 ();
 sg13g2_fill_1 FILLER_7_1403 ();
 sg13g2_decap_8 FILLER_7_1421 ();
 sg13g2_fill_2 FILLER_7_1428 ();
 sg13g2_decap_8 FILLER_7_1436 ();
 sg13g2_decap_8 FILLER_7_1443 ();
 sg13g2_decap_8 FILLER_7_1450 ();
 sg13g2_decap_8 FILLER_7_1457 ();
 sg13g2_decap_8 FILLER_7_1464 ();
 sg13g2_decap_8 FILLER_7_1471 ();
 sg13g2_decap_8 FILLER_7_1478 ();
 sg13g2_decap_4 FILLER_7_1485 ();
 sg13g2_fill_2 FILLER_7_1489 ();
 sg13g2_decap_8 FILLER_7_1495 ();
 sg13g2_decap_8 FILLER_7_1502 ();
 sg13g2_decap_8 FILLER_7_1509 ();
 sg13g2_decap_8 FILLER_7_1516 ();
 sg13g2_decap_8 FILLER_7_1523 ();
 sg13g2_decap_8 FILLER_7_1530 ();
 sg13g2_decap_8 FILLER_7_1537 ();
 sg13g2_decap_8 FILLER_7_1544 ();
 sg13g2_decap_8 FILLER_7_1551 ();
 sg13g2_decap_8 FILLER_7_1558 ();
 sg13g2_decap_8 FILLER_7_1565 ();
 sg13g2_decap_8 FILLER_7_1572 ();
 sg13g2_decap_8 FILLER_7_1579 ();
 sg13g2_decap_8 FILLER_7_1586 ();
 sg13g2_decap_8 FILLER_7_1593 ();
 sg13g2_decap_8 FILLER_7_1600 ();
 sg13g2_decap_8 FILLER_7_1607 ();
 sg13g2_decap_8 FILLER_7_1614 ();
 sg13g2_decap_8 FILLER_7_1621 ();
 sg13g2_decap_8 FILLER_7_1628 ();
 sg13g2_decap_8 FILLER_7_1635 ();
 sg13g2_decap_8 FILLER_7_1642 ();
 sg13g2_decap_8 FILLER_7_1649 ();
 sg13g2_decap_8 FILLER_7_1656 ();
 sg13g2_decap_8 FILLER_7_1663 ();
 sg13g2_decap_8 FILLER_7_1670 ();
 sg13g2_decap_8 FILLER_7_1677 ();
 sg13g2_decap_8 FILLER_7_1684 ();
 sg13g2_decap_8 FILLER_7_1691 ();
 sg13g2_decap_8 FILLER_7_1698 ();
 sg13g2_decap_8 FILLER_7_1705 ();
 sg13g2_decap_8 FILLER_7_1712 ();
 sg13g2_decap_8 FILLER_7_1719 ();
 sg13g2_decap_8 FILLER_7_1726 ();
 sg13g2_decap_8 FILLER_7_1733 ();
 sg13g2_decap_8 FILLER_7_1740 ();
 sg13g2_decap_8 FILLER_7_1747 ();
 sg13g2_decap_8 FILLER_7_1754 ();
 sg13g2_decap_8 FILLER_7_1761 ();
 sg13g2_decap_4 FILLER_7_1768 ();
 sg13g2_fill_2 FILLER_7_1772 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_4 FILLER_8_42 ();
 sg13g2_fill_2 FILLER_8_46 ();
 sg13g2_decap_4 FILLER_8_52 ();
 sg13g2_fill_1 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_62 ();
 sg13g2_fill_1 FILLER_8_77 ();
 sg13g2_fill_2 FILLER_8_82 ();
 sg13g2_fill_1 FILLER_8_88 ();
 sg13g2_decap_4 FILLER_8_94 ();
 sg13g2_fill_2 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_115 ();
 sg13g2_decap_4 FILLER_8_122 ();
 sg13g2_fill_1 FILLER_8_131 ();
 sg13g2_fill_2 FILLER_8_136 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_decap_4 FILLER_8_158 ();
 sg13g2_decap_4 FILLER_8_171 ();
 sg13g2_fill_1 FILLER_8_175 ();
 sg13g2_fill_2 FILLER_8_182 ();
 sg13g2_fill_1 FILLER_8_184 ();
 sg13g2_fill_2 FILLER_8_214 ();
 sg13g2_decap_4 FILLER_8_221 ();
 sg13g2_fill_2 FILLER_8_225 ();
 sg13g2_fill_2 FILLER_8_235 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_fill_1 FILLER_8_253 ();
 sg13g2_fill_2 FILLER_8_265 ();
 sg13g2_fill_1 FILLER_8_267 ();
 sg13g2_decap_8 FILLER_8_272 ();
 sg13g2_fill_2 FILLER_8_279 ();
 sg13g2_fill_1 FILLER_8_281 ();
 sg13g2_decap_8 FILLER_8_292 ();
 sg13g2_decap_4 FILLER_8_299 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_4 FILLER_8_314 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_decap_8 FILLER_8_325 ();
 sg13g2_decap_8 FILLER_8_332 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_fill_1 FILLER_8_365 ();
 sg13g2_fill_1 FILLER_8_370 ();
 sg13g2_fill_1 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_fill_1 FILLER_8_401 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_8_418 ();
 sg13g2_fill_1 FILLER_8_425 ();
 sg13g2_decap_8 FILLER_8_432 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_fill_2 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_fill_1 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_482 ();
 sg13g2_fill_2 FILLER_8_494 ();
 sg13g2_fill_1 FILLER_8_496 ();
 sg13g2_fill_2 FILLER_8_506 ();
 sg13g2_fill_1 FILLER_8_508 ();
 sg13g2_decap_4 FILLER_8_514 ();
 sg13g2_fill_1 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_524 ();
 sg13g2_decap_8 FILLER_8_531 ();
 sg13g2_decap_8 FILLER_8_538 ();
 sg13g2_decap_4 FILLER_8_545 ();
 sg13g2_fill_1 FILLER_8_549 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_4 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_590 ();
 sg13g2_decap_8 FILLER_8_597 ();
 sg13g2_decap_8 FILLER_8_604 ();
 sg13g2_decap_8 FILLER_8_615 ();
 sg13g2_decap_8 FILLER_8_622 ();
 sg13g2_fill_1 FILLER_8_629 ();
 sg13g2_fill_2 FILLER_8_635 ();
 sg13g2_decap_8 FILLER_8_667 ();
 sg13g2_fill_2 FILLER_8_674 ();
 sg13g2_fill_1 FILLER_8_676 ();
 sg13g2_decap_4 FILLER_8_682 ();
 sg13g2_decap_8 FILLER_8_690 ();
 sg13g2_decap_8 FILLER_8_697 ();
 sg13g2_decap_8 FILLER_8_704 ();
 sg13g2_decap_8 FILLER_8_711 ();
 sg13g2_fill_2 FILLER_8_718 ();
 sg13g2_decap_8 FILLER_8_746 ();
 sg13g2_decap_4 FILLER_8_753 ();
 sg13g2_fill_2 FILLER_8_757 ();
 sg13g2_decap_8 FILLER_8_766 ();
 sg13g2_decap_8 FILLER_8_773 ();
 sg13g2_decap_8 FILLER_8_780 ();
 sg13g2_decap_4 FILLER_8_787 ();
 sg13g2_fill_2 FILLER_8_791 ();
 sg13g2_fill_1 FILLER_8_797 ();
 sg13g2_decap_8 FILLER_8_829 ();
 sg13g2_fill_1 FILLER_8_836 ();
 sg13g2_fill_1 FILLER_8_841 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_2 FILLER_8_861 ();
 sg13g2_fill_1 FILLER_8_863 ();
 sg13g2_decap_8 FILLER_8_867 ();
 sg13g2_fill_2 FILLER_8_880 ();
 sg13g2_decap_8 FILLER_8_890 ();
 sg13g2_fill_2 FILLER_8_897 ();
 sg13g2_fill_1 FILLER_8_899 ();
 sg13g2_decap_8 FILLER_8_910 ();
 sg13g2_fill_2 FILLER_8_917 ();
 sg13g2_fill_1 FILLER_8_919 ();
 sg13g2_decap_4 FILLER_8_923 ();
 sg13g2_fill_1 FILLER_8_927 ();
 sg13g2_decap_8 FILLER_8_938 ();
 sg13g2_decap_8 FILLER_8_945 ();
 sg13g2_decap_8 FILLER_8_952 ();
 sg13g2_decap_8 FILLER_8_962 ();
 sg13g2_decap_4 FILLER_8_969 ();
 sg13g2_decap_8 FILLER_8_977 ();
 sg13g2_decap_8 FILLER_8_988 ();
 sg13g2_decap_8 FILLER_8_995 ();
 sg13g2_decap_8 FILLER_8_1007 ();
 sg13g2_decap_8 FILLER_8_1014 ();
 sg13g2_decap_8 FILLER_8_1021 ();
 sg13g2_decap_4 FILLER_8_1028 ();
 sg13g2_fill_2 FILLER_8_1032 ();
 sg13g2_decap_8 FILLER_8_1046 ();
 sg13g2_decap_8 FILLER_8_1053 ();
 sg13g2_decap_4 FILLER_8_1060 ();
 sg13g2_fill_2 FILLER_8_1064 ();
 sg13g2_decap_4 FILLER_8_1087 ();
 sg13g2_fill_1 FILLER_8_1091 ();
 sg13g2_fill_1 FILLER_8_1118 ();
 sg13g2_decap_8 FILLER_8_1129 ();
 sg13g2_decap_8 FILLER_8_1165 ();
 sg13g2_decap_8 FILLER_8_1172 ();
 sg13g2_fill_2 FILLER_8_1187 ();
 sg13g2_decap_8 FILLER_8_1192 ();
 sg13g2_decap_8 FILLER_8_1199 ();
 sg13g2_decap_4 FILLER_8_1206 ();
 sg13g2_decap_4 FILLER_8_1213 ();
 sg13g2_decap_8 FILLER_8_1243 ();
 sg13g2_decap_8 FILLER_8_1250 ();
 sg13g2_decap_8 FILLER_8_1257 ();
 sg13g2_decap_8 FILLER_8_1264 ();
 sg13g2_decap_8 FILLER_8_1271 ();
 sg13g2_decap_8 FILLER_8_1278 ();
 sg13g2_decap_8 FILLER_8_1285 ();
 sg13g2_decap_8 FILLER_8_1292 ();
 sg13g2_decap_8 FILLER_8_1299 ();
 sg13g2_fill_2 FILLER_8_1306 ();
 sg13g2_fill_1 FILLER_8_1317 ();
 sg13g2_decap_4 FILLER_8_1328 ();
 sg13g2_fill_1 FILLER_8_1332 ();
 sg13g2_fill_1 FILLER_8_1338 ();
 sg13g2_decap_4 FILLER_8_1350 ();
 sg13g2_fill_2 FILLER_8_1385 ();
 sg13g2_fill_2 FILLER_8_1397 ();
 sg13g2_fill_1 FILLER_8_1399 ();
 sg13g2_decap_4 FILLER_8_1410 ();
 sg13g2_fill_2 FILLER_8_1414 ();
 sg13g2_fill_1 FILLER_8_1427 ();
 sg13g2_decap_4 FILLER_8_1438 ();
 sg13g2_fill_1 FILLER_8_1442 ();
 sg13g2_decap_8 FILLER_8_1449 ();
 sg13g2_decap_8 FILLER_8_1456 ();
 sg13g2_decap_8 FILLER_8_1463 ();
 sg13g2_fill_2 FILLER_8_1470 ();
 sg13g2_decap_8 FILLER_8_1502 ();
 sg13g2_decap_8 FILLER_8_1509 ();
 sg13g2_decap_8 FILLER_8_1516 ();
 sg13g2_decap_8 FILLER_8_1523 ();
 sg13g2_decap_8 FILLER_8_1530 ();
 sg13g2_decap_8 FILLER_8_1537 ();
 sg13g2_decap_8 FILLER_8_1544 ();
 sg13g2_decap_8 FILLER_8_1551 ();
 sg13g2_decap_8 FILLER_8_1558 ();
 sg13g2_decap_8 FILLER_8_1565 ();
 sg13g2_decap_8 FILLER_8_1572 ();
 sg13g2_decap_8 FILLER_8_1579 ();
 sg13g2_decap_8 FILLER_8_1586 ();
 sg13g2_decap_8 FILLER_8_1593 ();
 sg13g2_decap_8 FILLER_8_1600 ();
 sg13g2_decap_8 FILLER_8_1607 ();
 sg13g2_decap_8 FILLER_8_1614 ();
 sg13g2_decap_8 FILLER_8_1621 ();
 sg13g2_decap_8 FILLER_8_1628 ();
 sg13g2_decap_8 FILLER_8_1635 ();
 sg13g2_decap_8 FILLER_8_1642 ();
 sg13g2_decap_8 FILLER_8_1649 ();
 sg13g2_decap_8 FILLER_8_1656 ();
 sg13g2_decap_8 FILLER_8_1663 ();
 sg13g2_decap_8 FILLER_8_1670 ();
 sg13g2_decap_8 FILLER_8_1677 ();
 sg13g2_decap_8 FILLER_8_1684 ();
 sg13g2_decap_8 FILLER_8_1691 ();
 sg13g2_decap_8 FILLER_8_1698 ();
 sg13g2_decap_8 FILLER_8_1705 ();
 sg13g2_decap_8 FILLER_8_1712 ();
 sg13g2_decap_8 FILLER_8_1719 ();
 sg13g2_decap_8 FILLER_8_1726 ();
 sg13g2_decap_8 FILLER_8_1733 ();
 sg13g2_decap_8 FILLER_8_1740 ();
 sg13g2_decap_8 FILLER_8_1747 ();
 sg13g2_decap_8 FILLER_8_1754 ();
 sg13g2_decap_8 FILLER_8_1761 ();
 sg13g2_decap_4 FILLER_8_1768 ();
 sg13g2_fill_2 FILLER_8_1772 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_37 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_67 ();
 sg13g2_fill_1 FILLER_9_75 ();
 sg13g2_fill_2 FILLER_9_91 ();
 sg13g2_fill_1 FILLER_9_93 ();
 sg13g2_decap_8 FILLER_9_136 ();
 sg13g2_fill_2 FILLER_9_143 ();
 sg13g2_decap_8 FILLER_9_150 ();
 sg13g2_decap_8 FILLER_9_157 ();
 sg13g2_fill_2 FILLER_9_164 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_172 ();
 sg13g2_decap_4 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_187 ();
 sg13g2_decap_4 FILLER_9_205 ();
 sg13g2_fill_2 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_decap_4 FILLER_9_236 ();
 sg13g2_decap_4 FILLER_9_249 ();
 sg13g2_fill_1 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_fill_1 FILLER_9_266 ();
 sg13g2_decap_4 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_296 ();
 sg13g2_fill_2 FILLER_9_314 ();
 sg13g2_fill_1 FILLER_9_320 ();
 sg13g2_fill_1 FILLER_9_326 ();
 sg13g2_decap_4 FILLER_9_340 ();
 sg13g2_fill_1 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_355 ();
 sg13g2_fill_1 FILLER_9_362 ();
 sg13g2_fill_2 FILLER_9_368 ();
 sg13g2_fill_1 FILLER_9_370 ();
 sg13g2_decap_4 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_decap_4 FILLER_9_408 ();
 sg13g2_fill_2 FILLER_9_417 ();
 sg13g2_fill_1 FILLER_9_424 ();
 sg13g2_fill_2 FILLER_9_435 ();
 sg13g2_fill_1 FILLER_9_437 ();
 sg13g2_decap_4 FILLER_9_448 ();
 sg13g2_fill_1 FILLER_9_452 ();
 sg13g2_fill_1 FILLER_9_461 ();
 sg13g2_decap_8 FILLER_9_471 ();
 sg13g2_fill_2 FILLER_9_478 ();
 sg13g2_decap_8 FILLER_9_484 ();
 sg13g2_decap_8 FILLER_9_491 ();
 sg13g2_decap_8 FILLER_9_498 ();
 sg13g2_decap_8 FILLER_9_505 ();
 sg13g2_decap_8 FILLER_9_512 ();
 sg13g2_decap_4 FILLER_9_519 ();
 sg13g2_fill_2 FILLER_9_523 ();
 sg13g2_decap_8 FILLER_9_530 ();
 sg13g2_decap_8 FILLER_9_537 ();
 sg13g2_decap_4 FILLER_9_544 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_fill_1 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_619 ();
 sg13g2_fill_2 FILLER_9_626 ();
 sg13g2_decap_4 FILLER_9_637 ();
 sg13g2_fill_2 FILLER_9_641 ();
 sg13g2_decap_8 FILLER_9_647 ();
 sg13g2_decap_8 FILLER_9_654 ();
 sg13g2_decap_8 FILLER_9_661 ();
 sg13g2_decap_4 FILLER_9_668 ();
 sg13g2_fill_2 FILLER_9_672 ();
 sg13g2_fill_1 FILLER_9_705 ();
 sg13g2_decap_8 FILLER_9_709 ();
 sg13g2_decap_8 FILLER_9_724 ();
 sg13g2_decap_8 FILLER_9_731 ();
 sg13g2_fill_2 FILLER_9_738 ();
 sg13g2_decap_8 FILLER_9_744 ();
 sg13g2_decap_8 FILLER_9_751 ();
 sg13g2_decap_8 FILLER_9_758 ();
 sg13g2_fill_2 FILLER_9_765 ();
 sg13g2_fill_1 FILLER_9_767 ();
 sg13g2_decap_8 FILLER_9_794 ();
 sg13g2_fill_2 FILLER_9_801 ();
 sg13g2_decap_4 FILLER_9_823 ();
 sg13g2_fill_2 FILLER_9_827 ();
 sg13g2_fill_2 FILLER_9_833 ();
 sg13g2_fill_1 FILLER_9_835 ();
 sg13g2_fill_2 FILLER_9_845 ();
 sg13g2_decap_8 FILLER_9_855 ();
 sg13g2_decap_8 FILLER_9_862 ();
 sg13g2_fill_2 FILLER_9_869 ();
 sg13g2_fill_1 FILLER_9_871 ();
 sg13g2_decap_4 FILLER_9_875 ();
 sg13g2_fill_1 FILLER_9_879 ();
 sg13g2_decap_8 FILLER_9_885 ();
 sg13g2_decap_8 FILLER_9_892 ();
 sg13g2_decap_8 FILLER_9_899 ();
 sg13g2_decap_8 FILLER_9_906 ();
 sg13g2_decap_8 FILLER_9_913 ();
 sg13g2_decap_8 FILLER_9_920 ();
 sg13g2_fill_2 FILLER_9_927 ();
 sg13g2_decap_4 FILLER_9_934 ();
 sg13g2_fill_1 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_955 ();
 sg13g2_decap_8 FILLER_9_962 ();
 sg13g2_decap_8 FILLER_9_969 ();
 sg13g2_fill_1 FILLER_9_976 ();
 sg13g2_decap_8 FILLER_9_981 ();
 sg13g2_decap_8 FILLER_9_988 ();
 sg13g2_decap_8 FILLER_9_995 ();
 sg13g2_decap_4 FILLER_9_1002 ();
 sg13g2_decap_4 FILLER_9_1032 ();
 sg13g2_decap_8 FILLER_9_1040 ();
 sg13g2_decap_8 FILLER_9_1047 ();
 sg13g2_decap_8 FILLER_9_1054 ();
 sg13g2_decap_4 FILLER_9_1061 ();
 sg13g2_fill_1 FILLER_9_1065 ();
 sg13g2_decap_8 FILLER_9_1078 ();
 sg13g2_decap_8 FILLER_9_1085 ();
 sg13g2_decap_4 FILLER_9_1092 ();
 sg13g2_fill_1 FILLER_9_1106 ();
 sg13g2_fill_1 FILLER_9_1117 ();
 sg13g2_decap_8 FILLER_9_1122 ();
 sg13g2_decap_8 FILLER_9_1129 ();
 sg13g2_decap_4 FILLER_9_1136 ();
 sg13g2_fill_2 FILLER_9_1140 ();
 sg13g2_decap_8 FILLER_9_1146 ();
 sg13g2_decap_8 FILLER_9_1153 ();
 sg13g2_decap_4 FILLER_9_1160 ();
 sg13g2_fill_1 FILLER_9_1164 ();
 sg13g2_decap_8 FILLER_9_1169 ();
 sg13g2_decap_8 FILLER_9_1176 ();
 sg13g2_decap_4 FILLER_9_1183 ();
 sg13g2_fill_2 FILLER_9_1187 ();
 sg13g2_decap_8 FILLER_9_1202 ();
 sg13g2_fill_1 FILLER_9_1209 ();
 sg13g2_fill_2 FILLER_9_1221 ();
 sg13g2_decap_8 FILLER_9_1233 ();
 sg13g2_fill_2 FILLER_9_1240 ();
 sg13g2_fill_1 FILLER_9_1242 ();
 sg13g2_fill_2 FILLER_9_1255 ();
 sg13g2_decap_8 FILLER_9_1261 ();
 sg13g2_fill_1 FILLER_9_1268 ();
 sg13g2_decap_8 FILLER_9_1273 ();
 sg13g2_decap_8 FILLER_9_1280 ();
 sg13g2_fill_2 FILLER_9_1287 ();
 sg13g2_fill_1 FILLER_9_1289 ();
 sg13g2_decap_8 FILLER_9_1294 ();
 sg13g2_fill_1 FILLER_9_1301 ();
 sg13g2_fill_2 FILLER_9_1312 ();
 sg13g2_fill_1 FILLER_9_1314 ();
 sg13g2_decap_8 FILLER_9_1328 ();
 sg13g2_decap_8 FILLER_9_1335 ();
 sg13g2_decap_8 FILLER_9_1342 ();
 sg13g2_decap_8 FILLER_9_1349 ();
 sg13g2_decap_8 FILLER_9_1356 ();
 sg13g2_decap_8 FILLER_9_1363 ();
 sg13g2_decap_8 FILLER_9_1370 ();
 sg13g2_decap_8 FILLER_9_1377 ();
 sg13g2_decap_4 FILLER_9_1384 ();
 sg13g2_fill_1 FILLER_9_1388 ();
 sg13g2_decap_8 FILLER_9_1396 ();
 sg13g2_decap_4 FILLER_9_1424 ();
 sg13g2_decap_8 FILLER_9_1433 ();
 sg13g2_decap_8 FILLER_9_1440 ();
 sg13g2_decap_8 FILLER_9_1447 ();
 sg13g2_decap_8 FILLER_9_1454 ();
 sg13g2_decap_8 FILLER_9_1461 ();
 sg13g2_decap_8 FILLER_9_1468 ();
 sg13g2_decap_8 FILLER_9_1475 ();
 sg13g2_decap_8 FILLER_9_1482 ();
 sg13g2_decap_8 FILLER_9_1489 ();
 sg13g2_decap_8 FILLER_9_1496 ();
 sg13g2_decap_8 FILLER_9_1503 ();
 sg13g2_decap_8 FILLER_9_1510 ();
 sg13g2_decap_8 FILLER_9_1517 ();
 sg13g2_decap_8 FILLER_9_1524 ();
 sg13g2_decap_8 FILLER_9_1531 ();
 sg13g2_decap_8 FILLER_9_1538 ();
 sg13g2_decap_8 FILLER_9_1545 ();
 sg13g2_decap_8 FILLER_9_1552 ();
 sg13g2_decap_8 FILLER_9_1559 ();
 sg13g2_decap_8 FILLER_9_1566 ();
 sg13g2_decap_8 FILLER_9_1573 ();
 sg13g2_decap_8 FILLER_9_1580 ();
 sg13g2_decap_8 FILLER_9_1587 ();
 sg13g2_decap_8 FILLER_9_1594 ();
 sg13g2_decap_8 FILLER_9_1601 ();
 sg13g2_decap_8 FILLER_9_1608 ();
 sg13g2_decap_8 FILLER_9_1615 ();
 sg13g2_decap_8 FILLER_9_1622 ();
 sg13g2_decap_8 FILLER_9_1629 ();
 sg13g2_decap_8 FILLER_9_1636 ();
 sg13g2_decap_8 FILLER_9_1643 ();
 sg13g2_decap_8 FILLER_9_1650 ();
 sg13g2_decap_8 FILLER_9_1657 ();
 sg13g2_decap_8 FILLER_9_1664 ();
 sg13g2_decap_8 FILLER_9_1671 ();
 sg13g2_decap_8 FILLER_9_1678 ();
 sg13g2_decap_8 FILLER_9_1685 ();
 sg13g2_decap_8 FILLER_9_1692 ();
 sg13g2_decap_8 FILLER_9_1699 ();
 sg13g2_decap_8 FILLER_9_1706 ();
 sg13g2_decap_8 FILLER_9_1713 ();
 sg13g2_decap_8 FILLER_9_1720 ();
 sg13g2_decap_8 FILLER_9_1727 ();
 sg13g2_decap_8 FILLER_9_1734 ();
 sg13g2_decap_8 FILLER_9_1741 ();
 sg13g2_decap_8 FILLER_9_1748 ();
 sg13g2_decap_8 FILLER_9_1755 ();
 sg13g2_decap_8 FILLER_9_1762 ();
 sg13g2_decap_4 FILLER_9_1769 ();
 sg13g2_fill_1 FILLER_9_1773 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_fill_2 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_37 ();
 sg13g2_decap_8 FILLER_10_44 ();
 sg13g2_fill_1 FILLER_10_51 ();
 sg13g2_fill_2 FILLER_10_57 ();
 sg13g2_decap_4 FILLER_10_75 ();
 sg13g2_fill_1 FILLER_10_83 ();
 sg13g2_decap_4 FILLER_10_98 ();
 sg13g2_fill_1 FILLER_10_102 ();
 sg13g2_fill_1 FILLER_10_114 ();
 sg13g2_fill_1 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_132 ();
 sg13g2_decap_8 FILLER_10_139 ();
 sg13g2_decap_8 FILLER_10_160 ();
 sg13g2_decap_8 FILLER_10_167 ();
 sg13g2_decap_8 FILLER_10_174 ();
 sg13g2_fill_2 FILLER_10_181 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_fill_2 FILLER_10_188 ();
 sg13g2_fill_1 FILLER_10_190 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_fill_2 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_240 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_decap_8 FILLER_10_253 ();
 sg13g2_decap_8 FILLER_10_264 ();
 sg13g2_fill_1 FILLER_10_271 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_decap_4 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_313 ();
 sg13g2_fill_2 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_332 ();
 sg13g2_fill_1 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_fill_2 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_fill_1 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_decap_8 FILLER_10_408 ();
 sg13g2_decap_4 FILLER_10_415 ();
 sg13g2_decap_4 FILLER_10_424 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_4 FILLER_10_445 ();
 sg13g2_fill_2 FILLER_10_449 ();
 sg13g2_decap_4 FILLER_10_467 ();
 sg13g2_fill_1 FILLER_10_471 ();
 sg13g2_decap_8 FILLER_10_477 ();
 sg13g2_fill_2 FILLER_10_484 ();
 sg13g2_fill_1 FILLER_10_486 ();
 sg13g2_decap_8 FILLER_10_493 ();
 sg13g2_decap_8 FILLER_10_500 ();
 sg13g2_decap_8 FILLER_10_507 ();
 sg13g2_decap_8 FILLER_10_514 ();
 sg13g2_fill_2 FILLER_10_521 ();
 sg13g2_fill_1 FILLER_10_523 ();
 sg13g2_decap_4 FILLER_10_529 ();
 sg13g2_fill_2 FILLER_10_533 ();
 sg13g2_decap_8 FILLER_10_541 ();
 sg13g2_decap_8 FILLER_10_548 ();
 sg13g2_decap_8 FILLER_10_555 ();
 sg13g2_decap_8 FILLER_10_562 ();
 sg13g2_fill_2 FILLER_10_569 ();
 sg13g2_decap_8 FILLER_10_575 ();
 sg13g2_decap_8 FILLER_10_582 ();
 sg13g2_decap_8 FILLER_10_603 ();
 sg13g2_fill_2 FILLER_10_610 ();
 sg13g2_fill_1 FILLER_10_612 ();
 sg13g2_decap_8 FILLER_10_617 ();
 sg13g2_fill_2 FILLER_10_624 ();
 sg13g2_decap_8 FILLER_10_635 ();
 sg13g2_decap_8 FILLER_10_642 ();
 sg13g2_decap_8 FILLER_10_649 ();
 sg13g2_fill_2 FILLER_10_656 ();
 sg13g2_decap_8 FILLER_10_662 ();
 sg13g2_fill_2 FILLER_10_669 ();
 sg13g2_fill_1 FILLER_10_671 ();
 sg13g2_decap_4 FILLER_10_676 ();
 sg13g2_fill_1 FILLER_10_680 ();
 sg13g2_decap_8 FILLER_10_685 ();
 sg13g2_decap_8 FILLER_10_692 ();
 sg13g2_decap_8 FILLER_10_699 ();
 sg13g2_decap_8 FILLER_10_706 ();
 sg13g2_fill_2 FILLER_10_725 ();
 sg13g2_fill_1 FILLER_10_727 ();
 sg13g2_fill_2 FILLER_10_746 ();
 sg13g2_fill_2 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_762 ();
 sg13g2_fill_1 FILLER_10_769 ();
 sg13g2_decap_4 FILLER_10_781 ();
 sg13g2_fill_1 FILLER_10_785 ();
 sg13g2_decap_8 FILLER_10_808 ();
 sg13g2_decap_4 FILLER_10_815 ();
 sg13g2_fill_2 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_824 ();
 sg13g2_decap_8 FILLER_10_831 ();
 sg13g2_fill_1 FILLER_10_838 ();
 sg13g2_fill_2 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_4 FILLER_10_861 ();
 sg13g2_fill_1 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_874 ();
 sg13g2_decap_8 FILLER_10_881 ();
 sg13g2_decap_8 FILLER_10_888 ();
 sg13g2_decap_4 FILLER_10_895 ();
 sg13g2_fill_2 FILLER_10_899 ();
 sg13g2_decap_8 FILLER_10_905 ();
 sg13g2_fill_2 FILLER_10_912 ();
 sg13g2_fill_1 FILLER_10_914 ();
 sg13g2_decap_4 FILLER_10_923 ();
 sg13g2_fill_1 FILLER_10_927 ();
 sg13g2_decap_4 FILLER_10_959 ();
 sg13g2_fill_1 FILLER_10_963 ();
 sg13g2_fill_1 FILLER_10_969 ();
 sg13g2_decap_8 FILLER_10_996 ();
 sg13g2_decap_4 FILLER_10_1003 ();
 sg13g2_fill_1 FILLER_10_1007 ();
 sg13g2_decap_8 FILLER_10_1017 ();
 sg13g2_decap_4 FILLER_10_1024 ();
 sg13g2_fill_2 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_10_1040 ();
 sg13g2_decap_8 FILLER_10_1047 ();
 sg13g2_decap_4 FILLER_10_1054 ();
 sg13g2_fill_1 FILLER_10_1058 ();
 sg13g2_fill_2 FILLER_10_1063 ();
 sg13g2_fill_2 FILLER_10_1071 ();
 sg13g2_fill_2 FILLER_10_1076 ();
 sg13g2_decap_8 FILLER_10_1090 ();
 sg13g2_fill_1 FILLER_10_1097 ();
 sg13g2_fill_2 FILLER_10_1104 ();
 sg13g2_fill_2 FILLER_10_1111 ();
 sg13g2_fill_1 FILLER_10_1113 ();
 sg13g2_fill_2 FILLER_10_1119 ();
 sg13g2_fill_1 FILLER_10_1121 ();
 sg13g2_fill_2 FILLER_10_1127 ();
 sg13g2_fill_2 FILLER_10_1138 ();
 sg13g2_fill_1 FILLER_10_1140 ();
 sg13g2_decap_8 FILLER_10_1149 ();
 sg13g2_fill_2 FILLER_10_1156 ();
 sg13g2_fill_1 FILLER_10_1158 ();
 sg13g2_decap_8 FILLER_10_1171 ();
 sg13g2_decap_8 FILLER_10_1178 ();
 sg13g2_decap_4 FILLER_10_1185 ();
 sg13g2_fill_2 FILLER_10_1189 ();
 sg13g2_decap_8 FILLER_10_1195 ();
 sg13g2_decap_4 FILLER_10_1202 ();
 sg13g2_fill_1 FILLER_10_1211 ();
 sg13g2_fill_1 FILLER_10_1224 ();
 sg13g2_decap_8 FILLER_10_1255 ();
 sg13g2_decap_4 FILLER_10_1288 ();
 sg13g2_decap_8 FILLER_10_1297 ();
 sg13g2_fill_1 FILLER_10_1304 ();
 sg13g2_decap_4 FILLER_10_1313 ();
 sg13g2_fill_2 FILLER_10_1317 ();
 sg13g2_decap_4 FILLER_10_1330 ();
 sg13g2_fill_2 FILLER_10_1334 ();
 sg13g2_decap_4 FILLER_10_1344 ();
 sg13g2_fill_2 FILLER_10_1364 ();
 sg13g2_decap_4 FILLER_10_1373 ();
 sg13g2_fill_1 FILLER_10_1377 ();
 sg13g2_decap_8 FILLER_10_1408 ();
 sg13g2_fill_2 FILLER_10_1415 ();
 sg13g2_fill_1 FILLER_10_1417 ();
 sg13g2_fill_1 FILLER_10_1423 ();
 sg13g2_fill_1 FILLER_10_1440 ();
 sg13g2_fill_2 FILLER_10_1455 ();
 sg13g2_fill_1 FILLER_10_1457 ();
 sg13g2_decap_4 FILLER_10_1462 ();
 sg13g2_fill_1 FILLER_10_1466 ();
 sg13g2_decap_8 FILLER_10_1471 ();
 sg13g2_decap_8 FILLER_10_1478 ();
 sg13g2_decap_8 FILLER_10_1485 ();
 sg13g2_decap_8 FILLER_10_1492 ();
 sg13g2_decap_8 FILLER_10_1499 ();
 sg13g2_decap_8 FILLER_10_1506 ();
 sg13g2_decap_8 FILLER_10_1513 ();
 sg13g2_decap_8 FILLER_10_1520 ();
 sg13g2_decap_8 FILLER_10_1527 ();
 sg13g2_decap_8 FILLER_10_1534 ();
 sg13g2_decap_8 FILLER_10_1541 ();
 sg13g2_decap_8 FILLER_10_1548 ();
 sg13g2_decap_8 FILLER_10_1555 ();
 sg13g2_decap_8 FILLER_10_1562 ();
 sg13g2_decap_8 FILLER_10_1569 ();
 sg13g2_decap_8 FILLER_10_1580 ();
 sg13g2_decap_8 FILLER_10_1587 ();
 sg13g2_decap_8 FILLER_10_1594 ();
 sg13g2_fill_2 FILLER_10_1601 ();
 sg13g2_fill_1 FILLER_10_1603 ();
 sg13g2_decap_8 FILLER_10_1608 ();
 sg13g2_decap_8 FILLER_10_1615 ();
 sg13g2_decap_8 FILLER_10_1622 ();
 sg13g2_decap_8 FILLER_10_1629 ();
 sg13g2_decap_8 FILLER_10_1636 ();
 sg13g2_decap_8 FILLER_10_1643 ();
 sg13g2_decap_8 FILLER_10_1650 ();
 sg13g2_decap_8 FILLER_10_1657 ();
 sg13g2_decap_8 FILLER_10_1664 ();
 sg13g2_decap_8 FILLER_10_1671 ();
 sg13g2_decap_8 FILLER_10_1678 ();
 sg13g2_decap_8 FILLER_10_1685 ();
 sg13g2_decap_8 FILLER_10_1692 ();
 sg13g2_decap_8 FILLER_10_1699 ();
 sg13g2_decap_8 FILLER_10_1706 ();
 sg13g2_decap_8 FILLER_10_1713 ();
 sg13g2_decap_8 FILLER_10_1720 ();
 sg13g2_decap_8 FILLER_10_1727 ();
 sg13g2_decap_8 FILLER_10_1734 ();
 sg13g2_decap_8 FILLER_10_1741 ();
 sg13g2_decap_8 FILLER_10_1748 ();
 sg13g2_decap_8 FILLER_10_1755 ();
 sg13g2_decap_8 FILLER_10_1762 ();
 sg13g2_decap_4 FILLER_10_1769 ();
 sg13g2_fill_1 FILLER_10_1773 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_fill_2 FILLER_11_49 ();
 sg13g2_fill_1 FILLER_11_51 ();
 sg13g2_fill_1 FILLER_11_61 ();
 sg13g2_decap_8 FILLER_11_67 ();
 sg13g2_fill_2 FILLER_11_74 ();
 sg13g2_fill_1 FILLER_11_76 ();
 sg13g2_fill_2 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_decap_4 FILLER_11_95 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_decap_8 FILLER_11_125 ();
 sg13g2_fill_2 FILLER_11_132 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_decap_8 FILLER_11_157 ();
 sg13g2_fill_2 FILLER_11_164 ();
 sg13g2_fill_1 FILLER_11_166 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_8 FILLER_11_184 ();
 sg13g2_decap_4 FILLER_11_191 ();
 sg13g2_fill_2 FILLER_11_204 ();
 sg13g2_fill_2 FILLER_11_210 ();
 sg13g2_decap_4 FILLER_11_222 ();
 sg13g2_decap_4 FILLER_11_231 ();
 sg13g2_fill_2 FILLER_11_240 ();
 sg13g2_decap_8 FILLER_11_254 ();
 sg13g2_fill_2 FILLER_11_261 ();
 sg13g2_fill_2 FILLER_11_269 ();
 sg13g2_fill_2 FILLER_11_276 ();
 sg13g2_fill_1 FILLER_11_278 ();
 sg13g2_fill_2 FILLER_11_284 ();
 sg13g2_decap_4 FILLER_11_291 ();
 sg13g2_fill_2 FILLER_11_295 ();
 sg13g2_decap_8 FILLER_11_302 ();
 sg13g2_decap_8 FILLER_11_309 ();
 sg13g2_decap_8 FILLER_11_316 ();
 sg13g2_decap_8 FILLER_11_323 ();
 sg13g2_fill_1 FILLER_11_330 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_fill_2 FILLER_11_350 ();
 sg13g2_fill_2 FILLER_11_360 ();
 sg13g2_decap_8 FILLER_11_377 ();
 sg13g2_decap_4 FILLER_11_384 ();
 sg13g2_fill_1 FILLER_11_388 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_4 FILLER_11_413 ();
 sg13g2_fill_1 FILLER_11_425 ();
 sg13g2_fill_2 FILLER_11_440 ();
 sg13g2_decap_4 FILLER_11_447 ();
 sg13g2_fill_1 FILLER_11_451 ();
 sg13g2_fill_1 FILLER_11_456 ();
 sg13g2_decap_8 FILLER_11_461 ();
 sg13g2_decap_8 FILLER_11_468 ();
 sg13g2_decap_8 FILLER_11_485 ();
 sg13g2_decap_4 FILLER_11_492 ();
 sg13g2_decap_8 FILLER_11_501 ();
 sg13g2_decap_8 FILLER_11_508 ();
 sg13g2_decap_8 FILLER_11_515 ();
 sg13g2_decap_8 FILLER_11_522 ();
 sg13g2_decap_8 FILLER_11_529 ();
 sg13g2_decap_8 FILLER_11_536 ();
 sg13g2_fill_2 FILLER_11_543 ();
 sg13g2_fill_1 FILLER_11_554 ();
 sg13g2_decap_8 FILLER_11_603 ();
 sg13g2_decap_4 FILLER_11_610 ();
 sg13g2_fill_2 FILLER_11_614 ();
 sg13g2_decap_8 FILLER_11_624 ();
 sg13g2_decap_4 FILLER_11_631 ();
 sg13g2_fill_1 FILLER_11_661 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_4 FILLER_11_711 ();
 sg13g2_fill_2 FILLER_11_715 ();
 sg13g2_fill_2 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_fill_1 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_741 ();
 sg13g2_decap_8 FILLER_11_748 ();
 sg13g2_decap_8 FILLER_11_755 ();
 sg13g2_decap_8 FILLER_11_762 ();
 sg13g2_decap_8 FILLER_11_773 ();
 sg13g2_decap_8 FILLER_11_780 ();
 sg13g2_decap_8 FILLER_11_787 ();
 sg13g2_decap_8 FILLER_11_794 ();
 sg13g2_decap_8 FILLER_11_801 ();
 sg13g2_fill_1 FILLER_11_808 ();
 sg13g2_decap_8 FILLER_11_822 ();
 sg13g2_fill_2 FILLER_11_829 ();
 sg13g2_fill_1 FILLER_11_844 ();
 sg13g2_decap_4 FILLER_11_852 ();
 sg13g2_decap_4 FILLER_11_860 ();
 sg13g2_fill_2 FILLER_11_864 ();
 sg13g2_decap_8 FILLER_11_871 ();
 sg13g2_decap_8 FILLER_11_878 ();
 sg13g2_decap_4 FILLER_11_885 ();
 sg13g2_fill_1 FILLER_11_889 ();
 sg13g2_decap_8 FILLER_11_894 ();
 sg13g2_decap_4 FILLER_11_901 ();
 sg13g2_fill_1 FILLER_11_905 ();
 sg13g2_decap_8 FILLER_11_924 ();
 sg13g2_decap_8 FILLER_11_931 ();
 sg13g2_decap_4 FILLER_11_941 ();
 sg13g2_decap_8 FILLER_11_953 ();
 sg13g2_decap_8 FILLER_11_960 ();
 sg13g2_decap_8 FILLER_11_967 ();
 sg13g2_decap_8 FILLER_11_974 ();
 sg13g2_fill_2 FILLER_11_981 ();
 sg13g2_decap_8 FILLER_11_988 ();
 sg13g2_decap_8 FILLER_11_995 ();
 sg13g2_decap_8 FILLER_11_1002 ();
 sg13g2_decap_4 FILLER_11_1009 ();
 sg13g2_fill_2 FILLER_11_1013 ();
 sg13g2_decap_4 FILLER_11_1019 ();
 sg13g2_fill_1 FILLER_11_1032 ();
 sg13g2_decap_8 FILLER_11_1038 ();
 sg13g2_decap_8 FILLER_11_1045 ();
 sg13g2_decap_8 FILLER_11_1052 ();
 sg13g2_decap_8 FILLER_11_1059 ();
 sg13g2_decap_4 FILLER_11_1066 ();
 sg13g2_decap_8 FILLER_11_1080 ();
 sg13g2_decap_8 FILLER_11_1087 ();
 sg13g2_decap_8 FILLER_11_1094 ();
 sg13g2_decap_8 FILLER_11_1101 ();
 sg13g2_fill_2 FILLER_11_1108 ();
 sg13g2_decap_8 FILLER_11_1117 ();
 sg13g2_decap_4 FILLER_11_1124 ();
 sg13g2_fill_2 FILLER_11_1128 ();
 sg13g2_decap_8 FILLER_11_1136 ();
 sg13g2_decap_4 FILLER_11_1143 ();
 sg13g2_fill_1 FILLER_11_1147 ();
 sg13g2_decap_8 FILLER_11_1197 ();
 sg13g2_fill_2 FILLER_11_1204 ();
 sg13g2_fill_1 FILLER_11_1206 ();
 sg13g2_decap_4 FILLER_11_1211 ();
 sg13g2_fill_1 FILLER_11_1221 ();
 sg13g2_decap_8 FILLER_11_1225 ();
 sg13g2_decap_8 FILLER_11_1232 ();
 sg13g2_decap_4 FILLER_11_1239 ();
 sg13g2_fill_2 FILLER_11_1243 ();
 sg13g2_decap_8 FILLER_11_1253 ();
 sg13g2_decap_8 FILLER_11_1260 ();
 sg13g2_decap_8 FILLER_11_1267 ();
 sg13g2_decap_8 FILLER_11_1274 ();
 sg13g2_decap_8 FILLER_11_1281 ();
 sg13g2_decap_8 FILLER_11_1288 ();
 sg13g2_decap_8 FILLER_11_1295 ();
 sg13g2_decap_8 FILLER_11_1302 ();
 sg13g2_decap_8 FILLER_11_1309 ();
 sg13g2_fill_1 FILLER_11_1316 ();
 sg13g2_decap_8 FILLER_11_1324 ();
 sg13g2_decap_8 FILLER_11_1331 ();
 sg13g2_fill_2 FILLER_11_1338 ();
 sg13g2_fill_1 FILLER_11_1340 ();
 sg13g2_decap_4 FILLER_11_1344 ();
 sg13g2_fill_2 FILLER_11_1348 ();
 sg13g2_fill_1 FILLER_11_1355 ();
 sg13g2_decap_4 FILLER_11_1361 ();
 sg13g2_fill_2 FILLER_11_1365 ();
 sg13g2_fill_2 FILLER_11_1384 ();
 sg13g2_decap_4 FILLER_11_1400 ();
 sg13g2_fill_2 FILLER_11_1409 ();
 sg13g2_fill_1 FILLER_11_1417 ();
 sg13g2_fill_1 FILLER_11_1425 ();
 sg13g2_fill_2 FILLER_11_1431 ();
 sg13g2_fill_2 FILLER_11_1440 ();
 sg13g2_fill_1 FILLER_11_1448 ();
 sg13g2_decap_4 FILLER_11_1459 ();
 sg13g2_fill_1 FILLER_11_1463 ();
 sg13g2_decap_8 FILLER_11_1469 ();
 sg13g2_decap_8 FILLER_11_1476 ();
 sg13g2_decap_8 FILLER_11_1483 ();
 sg13g2_decap_8 FILLER_11_1490 ();
 sg13g2_decap_8 FILLER_11_1497 ();
 sg13g2_decap_4 FILLER_11_1504 ();
 sg13g2_fill_2 FILLER_11_1508 ();
 sg13g2_decap_8 FILLER_11_1514 ();
 sg13g2_decap_8 FILLER_11_1521 ();
 sg13g2_decap_8 FILLER_11_1528 ();
 sg13g2_decap_4 FILLER_11_1535 ();
 sg13g2_decap_8 FILLER_11_1543 ();
 sg13g2_decap_8 FILLER_11_1550 ();
 sg13g2_decap_8 FILLER_11_1557 ();
 sg13g2_decap_4 FILLER_11_1564 ();
 sg13g2_fill_1 FILLER_11_1568 ();
 sg13g2_decap_8 FILLER_11_1595 ();
 sg13g2_decap_8 FILLER_11_1602 ();
 sg13g2_decap_8 FILLER_11_1609 ();
 sg13g2_decap_4 FILLER_11_1616 ();
 sg13g2_decap_8 FILLER_11_1624 ();
 sg13g2_decap_8 FILLER_11_1631 ();
 sg13g2_decap_8 FILLER_11_1638 ();
 sg13g2_decap_8 FILLER_11_1645 ();
 sg13g2_decap_8 FILLER_11_1652 ();
 sg13g2_decap_8 FILLER_11_1659 ();
 sg13g2_decap_8 FILLER_11_1666 ();
 sg13g2_decap_8 FILLER_11_1673 ();
 sg13g2_decap_8 FILLER_11_1680 ();
 sg13g2_decap_8 FILLER_11_1687 ();
 sg13g2_decap_8 FILLER_11_1694 ();
 sg13g2_decap_8 FILLER_11_1701 ();
 sg13g2_decap_8 FILLER_11_1708 ();
 sg13g2_decap_8 FILLER_11_1715 ();
 sg13g2_decap_8 FILLER_11_1722 ();
 sg13g2_decap_8 FILLER_11_1729 ();
 sg13g2_decap_8 FILLER_11_1736 ();
 sg13g2_decap_8 FILLER_11_1743 ();
 sg13g2_decap_8 FILLER_11_1750 ();
 sg13g2_decap_8 FILLER_11_1757 ();
 sg13g2_decap_8 FILLER_11_1764 ();
 sg13g2_fill_2 FILLER_11_1771 ();
 sg13g2_fill_1 FILLER_11_1773 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_4 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_43 ();
 sg13g2_decap_4 FILLER_12_50 ();
 sg13g2_fill_1 FILLER_12_54 ();
 sg13g2_decap_4 FILLER_12_60 ();
 sg13g2_fill_1 FILLER_12_64 ();
 sg13g2_fill_1 FILLER_12_70 ();
 sg13g2_fill_2 FILLER_12_76 ();
 sg13g2_fill_1 FILLER_12_78 ();
 sg13g2_decap_4 FILLER_12_97 ();
 sg13g2_fill_1 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_107 ();
 sg13g2_fill_2 FILLER_12_117 ();
 sg13g2_fill_1 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_125 ();
 sg13g2_decap_8 FILLER_12_132 ();
 sg13g2_fill_2 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_141 ();
 sg13g2_fill_2 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_164 ();
 sg13g2_decap_4 FILLER_12_171 ();
 sg13g2_fill_1 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_216 ();
 sg13g2_decap_4 FILLER_12_223 ();
 sg13g2_fill_2 FILLER_12_227 ();
 sg13g2_decap_4 FILLER_12_243 ();
 sg13g2_fill_2 FILLER_12_275 ();
 sg13g2_fill_1 FILLER_12_277 ();
 sg13g2_decap_4 FILLER_12_289 ();
 sg13g2_fill_2 FILLER_12_293 ();
 sg13g2_decap_8 FILLER_12_300 ();
 sg13g2_decap_8 FILLER_12_307 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_decap_4 FILLER_12_328 ();
 sg13g2_fill_1 FILLER_12_332 ();
 sg13g2_decap_8 FILLER_12_352 ();
 sg13g2_fill_2 FILLER_12_359 ();
 sg13g2_fill_1 FILLER_12_365 ();
 sg13g2_fill_1 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_fill_2 FILLER_12_388 ();
 sg13g2_fill_1 FILLER_12_390 ();
 sg13g2_fill_1 FILLER_12_396 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_12_415 ();
 sg13g2_decap_4 FILLER_12_422 ();
 sg13g2_fill_2 FILLER_12_426 ();
 sg13g2_fill_2 FILLER_12_436 ();
 sg13g2_fill_1 FILLER_12_438 ();
 sg13g2_decap_4 FILLER_12_443 ();
 sg13g2_fill_1 FILLER_12_447 ();
 sg13g2_decap_8 FILLER_12_453 ();
 sg13g2_decap_4 FILLER_12_460 ();
 sg13g2_fill_2 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_fill_1 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_501 ();
 sg13g2_fill_2 FILLER_12_508 ();
 sg13g2_fill_1 FILLER_12_510 ();
 sg13g2_decap_8 FILLER_12_516 ();
 sg13g2_decap_8 FILLER_12_523 ();
 sg13g2_decap_8 FILLER_12_530 ();
 sg13g2_decap_8 FILLER_12_537 ();
 sg13g2_decap_8 FILLER_12_544 ();
 sg13g2_decap_8 FILLER_12_551 ();
 sg13g2_decap_4 FILLER_12_558 ();
 sg13g2_decap_8 FILLER_12_566 ();
 sg13g2_decap_8 FILLER_12_573 ();
 sg13g2_decap_4 FILLER_12_580 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_fill_2 FILLER_12_623 ();
 sg13g2_fill_1 FILLER_12_625 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_fill_2 FILLER_12_648 ();
 sg13g2_fill_1 FILLER_12_650 ();
 sg13g2_decap_8 FILLER_12_656 ();
 sg13g2_decap_8 FILLER_12_663 ();
 sg13g2_decap_4 FILLER_12_670 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_4 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_722 ();
 sg13g2_decap_8 FILLER_12_729 ();
 sg13g2_decap_8 FILLER_12_775 ();
 sg13g2_fill_2 FILLER_12_782 ();
 sg13g2_decap_8 FILLER_12_815 ();
 sg13g2_decap_8 FILLER_12_822 ();
 sg13g2_decap_4 FILLER_12_829 ();
 sg13g2_fill_2 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_879 ();
 sg13g2_fill_1 FILLER_12_886 ();
 sg13g2_decap_8 FILLER_12_892 ();
 sg13g2_decap_8 FILLER_12_899 ();
 sg13g2_decap_4 FILLER_12_906 ();
 sg13g2_decap_4 FILLER_12_925 ();
 sg13g2_fill_2 FILLER_12_929 ();
 sg13g2_fill_2 FILLER_12_939 ();
 sg13g2_fill_1 FILLER_12_941 ();
 sg13g2_decap_8 FILLER_12_948 ();
 sg13g2_fill_2 FILLER_12_963 ();
 sg13g2_fill_2 FILLER_12_991 ();
 sg13g2_fill_2 FILLER_12_997 ();
 sg13g2_fill_2 FILLER_12_1007 ();
 sg13g2_fill_1 FILLER_12_1009 ();
 sg13g2_decap_8 FILLER_12_1035 ();
 sg13g2_decap_4 FILLER_12_1042 ();
 sg13g2_decap_8 FILLER_12_1054 ();
 sg13g2_fill_2 FILLER_12_1061 ();
 sg13g2_fill_2 FILLER_12_1071 ();
 sg13g2_decap_8 FILLER_12_1083 ();
 sg13g2_decap_8 FILLER_12_1090 ();
 sg13g2_decap_8 FILLER_12_1097 ();
 sg13g2_decap_4 FILLER_12_1104 ();
 sg13g2_decap_8 FILLER_12_1116 ();
 sg13g2_decap_4 FILLER_12_1123 ();
 sg13g2_decap_8 FILLER_12_1131 ();
 sg13g2_decap_8 FILLER_12_1138 ();
 sg13g2_fill_2 FILLER_12_1176 ();
 sg13g2_decap_8 FILLER_12_1181 ();
 sg13g2_decap_8 FILLER_12_1188 ();
 sg13g2_fill_2 FILLER_12_1195 ();
 sg13g2_fill_1 FILLER_12_1197 ();
 sg13g2_decap_8 FILLER_12_1224 ();
 sg13g2_decap_8 FILLER_12_1231 ();
 sg13g2_decap_8 FILLER_12_1238 ();
 sg13g2_decap_8 FILLER_12_1245 ();
 sg13g2_decap_8 FILLER_12_1252 ();
 sg13g2_fill_2 FILLER_12_1259 ();
 sg13g2_fill_1 FILLER_12_1261 ();
 sg13g2_fill_1 FILLER_12_1268 ();
 sg13g2_fill_1 FILLER_12_1273 ();
 sg13g2_decap_8 FILLER_12_1278 ();
 sg13g2_fill_1 FILLER_12_1285 ();
 sg13g2_fill_2 FILLER_12_1291 ();
 sg13g2_decap_8 FILLER_12_1323 ();
 sg13g2_decap_8 FILLER_12_1330 ();
 sg13g2_fill_2 FILLER_12_1337 ();
 sg13g2_decap_4 FILLER_12_1343 ();
 sg13g2_fill_1 FILLER_12_1347 ();
 sg13g2_decap_8 FILLER_12_1356 ();
 sg13g2_decap_8 FILLER_12_1363 ();
 sg13g2_fill_2 FILLER_12_1370 ();
 sg13g2_fill_1 FILLER_12_1372 ();
 sg13g2_decap_8 FILLER_12_1390 ();
 sg13g2_decap_8 FILLER_12_1397 ();
 sg13g2_fill_2 FILLER_12_1404 ();
 sg13g2_fill_1 FILLER_12_1406 ();
 sg13g2_fill_2 FILLER_12_1411 ();
 sg13g2_fill_2 FILLER_12_1423 ();
 sg13g2_fill_1 FILLER_12_1425 ();
 sg13g2_fill_1 FILLER_12_1434 ();
 sg13g2_fill_2 FILLER_12_1443 ();
 sg13g2_fill_2 FILLER_12_1450 ();
 sg13g2_decap_8 FILLER_12_1457 ();
 sg13g2_decap_8 FILLER_12_1464 ();
 sg13g2_decap_4 FILLER_12_1471 ();
 sg13g2_fill_2 FILLER_12_1475 ();
 sg13g2_decap_8 FILLER_12_1481 ();
 sg13g2_decap_8 FILLER_12_1488 ();
 sg13g2_decap_8 FILLER_12_1495 ();
 sg13g2_fill_2 FILLER_12_1502 ();
 sg13g2_decap_4 FILLER_12_1530 ();
 sg13g2_fill_1 FILLER_12_1534 ();
 sg13g2_decap_8 FILLER_12_1561 ();
 sg13g2_decap_8 FILLER_12_1568 ();
 sg13g2_decap_8 FILLER_12_1575 ();
 sg13g2_decap_8 FILLER_12_1582 ();
 sg13g2_fill_2 FILLER_12_1589 ();
 sg13g2_decap_8 FILLER_12_1604 ();
 sg13g2_decap_8 FILLER_12_1637 ();
 sg13g2_decap_8 FILLER_12_1644 ();
 sg13g2_decap_8 FILLER_12_1651 ();
 sg13g2_decap_8 FILLER_12_1658 ();
 sg13g2_decap_8 FILLER_12_1665 ();
 sg13g2_decap_8 FILLER_12_1672 ();
 sg13g2_decap_8 FILLER_12_1679 ();
 sg13g2_decap_8 FILLER_12_1686 ();
 sg13g2_decap_8 FILLER_12_1693 ();
 sg13g2_decap_8 FILLER_12_1700 ();
 sg13g2_decap_8 FILLER_12_1707 ();
 sg13g2_decap_8 FILLER_12_1714 ();
 sg13g2_decap_8 FILLER_12_1721 ();
 sg13g2_decap_8 FILLER_12_1728 ();
 sg13g2_decap_8 FILLER_12_1735 ();
 sg13g2_decap_8 FILLER_12_1742 ();
 sg13g2_decap_8 FILLER_12_1749 ();
 sg13g2_decap_8 FILLER_12_1756 ();
 sg13g2_decap_8 FILLER_12_1763 ();
 sg13g2_decap_4 FILLER_12_1770 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_32 ();
 sg13g2_decap_4 FILLER_13_37 ();
 sg13g2_fill_1 FILLER_13_45 ();
 sg13g2_decap_4 FILLER_13_55 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_fill_2 FILLER_13_102 ();
 sg13g2_fill_1 FILLER_13_104 ();
 sg13g2_decap_4 FILLER_13_111 ();
 sg13g2_decap_4 FILLER_13_119 ();
 sg13g2_fill_2 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_fill_2 FILLER_13_139 ();
 sg13g2_fill_2 FILLER_13_146 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_fill_2 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_187 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_209 ();
 sg13g2_decap_4 FILLER_13_215 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_230 ();
 sg13g2_fill_2 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_239 ();
 sg13g2_fill_2 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_fill_2 FILLER_13_254 ();
 sg13g2_fill_1 FILLER_13_256 ();
 sg13g2_decap_4 FILLER_13_265 ();
 sg13g2_fill_1 FILLER_13_269 ();
 sg13g2_decap_4 FILLER_13_280 ();
 sg13g2_fill_2 FILLER_13_284 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_fill_2 FILLER_13_297 ();
 sg13g2_decap_4 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_4 FILLER_13_336 ();
 sg13g2_fill_2 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_decap_4 FILLER_13_365 ();
 sg13g2_fill_1 FILLER_13_369 ();
 sg13g2_fill_2 FILLER_13_374 ();
 sg13g2_decap_4 FILLER_13_381 ();
 sg13g2_decap_4 FILLER_13_389 ();
 sg13g2_fill_1 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_4 FILLER_13_412 ();
 sg13g2_fill_2 FILLER_13_416 ();
 sg13g2_decap_4 FILLER_13_423 ();
 sg13g2_fill_1 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_433 ();
 sg13g2_decap_4 FILLER_13_440 ();
 sg13g2_decap_8 FILLER_13_449 ();
 sg13g2_fill_1 FILLER_13_456 ();
 sg13g2_decap_4 FILLER_13_472 ();
 sg13g2_decap_8 FILLER_13_481 ();
 sg13g2_fill_1 FILLER_13_488 ();
 sg13g2_decap_8 FILLER_13_494 ();
 sg13g2_decap_8 FILLER_13_501 ();
 sg13g2_decap_8 FILLER_13_508 ();
 sg13g2_decap_8 FILLER_13_515 ();
 sg13g2_decap_8 FILLER_13_522 ();
 sg13g2_decap_8 FILLER_13_529 ();
 sg13g2_decap_8 FILLER_13_536 ();
 sg13g2_fill_2 FILLER_13_543 ();
 sg13g2_fill_1 FILLER_13_545 ();
 sg13g2_decap_8 FILLER_13_572 ();
 sg13g2_decap_8 FILLER_13_579 ();
 sg13g2_decap_8 FILLER_13_591 ();
 sg13g2_decap_8 FILLER_13_598 ();
 sg13g2_decap_8 FILLER_13_605 ();
 sg13g2_decap_8 FILLER_13_612 ();
 sg13g2_decap_8 FILLER_13_619 ();
 sg13g2_decap_8 FILLER_13_626 ();
 sg13g2_decap_8 FILLER_13_633 ();
 sg13g2_fill_2 FILLER_13_645 ();
 sg13g2_fill_1 FILLER_13_647 ();
 sg13g2_fill_2 FILLER_13_678 ();
 sg13g2_fill_1 FILLER_13_680 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_4 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_727 ();
 sg13g2_decap_8 FILLER_13_734 ();
 sg13g2_decap_4 FILLER_13_741 ();
 sg13g2_fill_2 FILLER_13_745 ();
 sg13g2_decap_8 FILLER_13_751 ();
 sg13g2_decap_8 FILLER_13_758 ();
 sg13g2_decap_4 FILLER_13_765 ();
 sg13g2_decap_8 FILLER_13_773 ();
 sg13g2_decap_4 FILLER_13_780 ();
 sg13g2_fill_1 FILLER_13_784 ();
 sg13g2_fill_2 FILLER_13_792 ();
 sg13g2_decap_8 FILLER_13_807 ();
 sg13g2_decap_8 FILLER_13_814 ();
 sg13g2_decap_8 FILLER_13_821 ();
 sg13g2_decap_8 FILLER_13_828 ();
 sg13g2_decap_8 FILLER_13_835 ();
 sg13g2_decap_8 FILLER_13_842 ();
 sg13g2_decap_8 FILLER_13_849 ();
 sg13g2_decap_8 FILLER_13_856 ();
 sg13g2_decap_8 FILLER_13_863 ();
 sg13g2_decap_4 FILLER_13_870 ();
 sg13g2_fill_1 FILLER_13_874 ();
 sg13g2_decap_8 FILLER_13_880 ();
 sg13g2_decap_4 FILLER_13_913 ();
 sg13g2_fill_1 FILLER_13_917 ();
 sg13g2_decap_8 FILLER_13_922 ();
 sg13g2_decap_4 FILLER_13_929 ();
 sg13g2_decap_8 FILLER_13_950 ();
 sg13g2_decap_8 FILLER_13_957 ();
 sg13g2_decap_4 FILLER_13_964 ();
 sg13g2_fill_1 FILLER_13_968 ();
 sg13g2_decap_8 FILLER_13_974 ();
 sg13g2_decap_4 FILLER_13_981 ();
 sg13g2_fill_2 FILLER_13_985 ();
 sg13g2_decap_8 FILLER_13_992 ();
 sg13g2_decap_8 FILLER_13_999 ();
 sg13g2_decap_8 FILLER_13_1006 ();
 sg13g2_decap_8 FILLER_13_1013 ();
 sg13g2_decap_8 FILLER_13_1020 ();
 sg13g2_decap_8 FILLER_13_1027 ();
 sg13g2_decap_8 FILLER_13_1034 ();
 sg13g2_decap_8 FILLER_13_1041 ();
 sg13g2_decap_8 FILLER_13_1048 ();
 sg13g2_decap_4 FILLER_13_1055 ();
 sg13g2_decap_8 FILLER_13_1094 ();
 sg13g2_decap_8 FILLER_13_1101 ();
 sg13g2_decap_8 FILLER_13_1112 ();
 sg13g2_decap_8 FILLER_13_1145 ();
 sg13g2_decap_4 FILLER_13_1152 ();
 sg13g2_fill_2 FILLER_13_1156 ();
 sg13g2_decap_8 FILLER_13_1162 ();
 sg13g2_decap_8 FILLER_13_1169 ();
 sg13g2_decap_8 FILLER_13_1176 ();
 sg13g2_decap_8 FILLER_13_1183 ();
 sg13g2_decap_8 FILLER_13_1190 ();
 sg13g2_decap_8 FILLER_13_1197 ();
 sg13g2_decap_8 FILLER_13_1204 ();
 sg13g2_decap_8 FILLER_13_1211 ();
 sg13g2_decap_8 FILLER_13_1218 ();
 sg13g2_decap_8 FILLER_13_1225 ();
 sg13g2_decap_8 FILLER_13_1232 ();
 sg13g2_fill_1 FILLER_13_1239 ();
 sg13g2_decap_8 FILLER_13_1245 ();
 sg13g2_fill_1 FILLER_13_1257 ();
 sg13g2_decap_8 FILLER_13_1294 ();
 sg13g2_decap_8 FILLER_13_1301 ();
 sg13g2_decap_8 FILLER_13_1308 ();
 sg13g2_decap_8 FILLER_13_1315 ();
 sg13g2_decap_8 FILLER_13_1322 ();
 sg13g2_decap_8 FILLER_13_1329 ();
 sg13g2_decap_4 FILLER_13_1336 ();
 sg13g2_decap_8 FILLER_13_1371 ();
 sg13g2_decap_8 FILLER_13_1378 ();
 sg13g2_decap_8 FILLER_13_1385 ();
 sg13g2_decap_8 FILLER_13_1392 ();
 sg13g2_decap_8 FILLER_13_1399 ();
 sg13g2_decap_4 FILLER_13_1406 ();
 sg13g2_fill_2 FILLER_13_1410 ();
 sg13g2_decap_8 FILLER_13_1417 ();
 sg13g2_decap_8 FILLER_13_1424 ();
 sg13g2_fill_1 FILLER_13_1436 ();
 sg13g2_decap_8 FILLER_13_1447 ();
 sg13g2_fill_1 FILLER_13_1454 ();
 sg13g2_decap_4 FILLER_13_1459 ();
 sg13g2_fill_2 FILLER_13_1463 ();
 sg13g2_fill_1 FILLER_13_1469 ();
 sg13g2_decap_4 FILLER_13_1496 ();
 sg13g2_fill_2 FILLER_13_1500 ();
 sg13g2_decap_8 FILLER_13_1506 ();
 sg13g2_decap_8 FILLER_13_1513 ();
 sg13g2_decap_8 FILLER_13_1520 ();
 sg13g2_fill_2 FILLER_13_1527 ();
 sg13g2_decap_8 FILLER_13_1533 ();
 sg13g2_decap_8 FILLER_13_1540 ();
 sg13g2_decap_8 FILLER_13_1547 ();
 sg13g2_decap_4 FILLER_13_1554 ();
 sg13g2_fill_2 FILLER_13_1558 ();
 sg13g2_fill_2 FILLER_13_1573 ();
 sg13g2_fill_1 FILLER_13_1575 ();
 sg13g2_fill_2 FILLER_13_1581 ();
 sg13g2_fill_1 FILLER_13_1583 ();
 sg13g2_decap_8 FILLER_13_1615 ();
 sg13g2_decap_8 FILLER_13_1622 ();
 sg13g2_decap_8 FILLER_13_1634 ();
 sg13g2_decap_8 FILLER_13_1641 ();
 sg13g2_fill_1 FILLER_13_1648 ();
 sg13g2_decap_8 FILLER_13_1675 ();
 sg13g2_decap_8 FILLER_13_1682 ();
 sg13g2_decap_8 FILLER_13_1689 ();
 sg13g2_decap_8 FILLER_13_1696 ();
 sg13g2_decap_8 FILLER_13_1703 ();
 sg13g2_decap_8 FILLER_13_1710 ();
 sg13g2_decap_8 FILLER_13_1717 ();
 sg13g2_decap_8 FILLER_13_1724 ();
 sg13g2_decap_8 FILLER_13_1731 ();
 sg13g2_decap_8 FILLER_13_1738 ();
 sg13g2_decap_8 FILLER_13_1745 ();
 sg13g2_decap_8 FILLER_13_1752 ();
 sg13g2_decap_8 FILLER_13_1759 ();
 sg13g2_decap_8 FILLER_13_1766 ();
 sg13g2_fill_1 FILLER_13_1773 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_4 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_54 ();
 sg13g2_decap_4 FILLER_14_61 ();
 sg13g2_fill_2 FILLER_14_65 ();
 sg13g2_fill_1 FILLER_14_71 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_93 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_104 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_decap_4 FILLER_14_126 ();
 sg13g2_fill_2 FILLER_14_130 ();
 sg13g2_decap_4 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_fill_2 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_165 ();
 sg13g2_fill_2 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_4 FILLER_14_196 ();
 sg13g2_fill_2 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_fill_2 FILLER_14_229 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_decap_8 FILLER_14_262 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_fill_1 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_fill_2 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_4 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_fill_2 FILLER_14_371 ();
 sg13g2_fill_2 FILLER_14_379 ();
 sg13g2_fill_2 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_410 ();
 sg13g2_decap_4 FILLER_14_417 ();
 sg13g2_decap_4 FILLER_14_432 ();
 sg13g2_decap_4 FILLER_14_446 ();
 sg13g2_fill_1 FILLER_14_450 ();
 sg13g2_decap_8 FILLER_14_463 ();
 sg13g2_decap_8 FILLER_14_470 ();
 sg13g2_fill_1 FILLER_14_477 ();
 sg13g2_decap_8 FILLER_14_488 ();
 sg13g2_decap_8 FILLER_14_495 ();
 sg13g2_decap_8 FILLER_14_502 ();
 sg13g2_decap_8 FILLER_14_509 ();
 sg13g2_decap_8 FILLER_14_516 ();
 sg13g2_decap_8 FILLER_14_523 ();
 sg13g2_decap_8 FILLER_14_530 ();
 sg13g2_decap_8 FILLER_14_537 ();
 sg13g2_decap_8 FILLER_14_544 ();
 sg13g2_fill_1 FILLER_14_551 ();
 sg13g2_decap_4 FILLER_14_566 ();
 sg13g2_fill_1 FILLER_14_570 ();
 sg13g2_decap_8 FILLER_14_575 ();
 sg13g2_decap_8 FILLER_14_582 ();
 sg13g2_decap_8 FILLER_14_593 ();
 sg13g2_decap_4 FILLER_14_600 ();
 sg13g2_fill_2 FILLER_14_604 ();
 sg13g2_fill_2 FILLER_14_611 ();
 sg13g2_decap_8 FILLER_14_643 ();
 sg13g2_fill_2 FILLER_14_650 ();
 sg13g2_fill_1 FILLER_14_652 ();
 sg13g2_decap_8 FILLER_14_657 ();
 sg13g2_decap_8 FILLER_14_664 ();
 sg13g2_decap_4 FILLER_14_671 ();
 sg13g2_decap_8 FILLER_14_678 ();
 sg13g2_fill_2 FILLER_14_685 ();
 sg13g2_decap_8 FILLER_14_691 ();
 sg13g2_decap_8 FILLER_14_698 ();
 sg13g2_fill_2 FILLER_14_705 ();
 sg13g2_fill_2 FILLER_14_719 ();
 sg13g2_fill_1 FILLER_14_721 ();
 sg13g2_decap_4 FILLER_14_730 ();
 sg13g2_fill_1 FILLER_14_734 ();
 sg13g2_decap_8 FILLER_14_739 ();
 sg13g2_decap_8 FILLER_14_746 ();
 sg13g2_decap_8 FILLER_14_753 ();
 sg13g2_fill_2 FILLER_14_760 ();
 sg13g2_fill_1 FILLER_14_762 ();
 sg13g2_decap_8 FILLER_14_767 ();
 sg13g2_fill_2 FILLER_14_774 ();
 sg13g2_fill_1 FILLER_14_776 ();
 sg13g2_decap_8 FILLER_14_781 ();
 sg13g2_decap_4 FILLER_14_788 ();
 sg13g2_fill_2 FILLER_14_792 ();
 sg13g2_decap_4 FILLER_14_820 ();
 sg13g2_decap_8 FILLER_14_857 ();
 sg13g2_fill_2 FILLER_14_864 ();
 sg13g2_decap_8 FILLER_14_871 ();
 sg13g2_decap_8 FILLER_14_878 ();
 sg13g2_decap_8 FILLER_14_885 ();
 sg13g2_fill_1 FILLER_14_892 ();
 sg13g2_decap_8 FILLER_14_897 ();
 sg13g2_decap_8 FILLER_14_904 ();
 sg13g2_decap_8 FILLER_14_911 ();
 sg13g2_decap_8 FILLER_14_918 ();
 sg13g2_decap_8 FILLER_14_925 ();
 sg13g2_decap_4 FILLER_14_932 ();
 sg13g2_fill_1 FILLER_14_936 ();
 sg13g2_decap_8 FILLER_14_953 ();
 sg13g2_decap_8 FILLER_14_960 ();
 sg13g2_decap_8 FILLER_14_967 ();
 sg13g2_decap_8 FILLER_14_974 ();
 sg13g2_decap_8 FILLER_14_981 ();
 sg13g2_fill_1 FILLER_14_1014 ();
 sg13g2_decap_8 FILLER_14_1019 ();
 sg13g2_decap_4 FILLER_14_1026 ();
 sg13g2_fill_1 FILLER_14_1030 ();
 sg13g2_decap_8 FILLER_14_1034 ();
 sg13g2_decap_4 FILLER_14_1041 ();
 sg13g2_fill_1 FILLER_14_1045 ();
 sg13g2_decap_8 FILLER_14_1066 ();
 sg13g2_decap_8 FILLER_14_1073 ();
 sg13g2_decap_8 FILLER_14_1080 ();
 sg13g2_decap_4 FILLER_14_1087 ();
 sg13g2_fill_2 FILLER_14_1091 ();
 sg13g2_fill_2 FILLER_14_1096 ();
 sg13g2_fill_1 FILLER_14_1098 ();
 sg13g2_decap_8 FILLER_14_1118 ();
 sg13g2_fill_1 FILLER_14_1125 ();
 sg13g2_decap_8 FILLER_14_1130 ();
 sg13g2_fill_1 FILLER_14_1137 ();
 sg13g2_decap_8 FILLER_14_1142 ();
 sg13g2_decap_8 FILLER_14_1149 ();
 sg13g2_decap_8 FILLER_14_1156 ();
 sg13g2_decap_8 FILLER_14_1163 ();
 sg13g2_decap_8 FILLER_14_1170 ();
 sg13g2_decap_8 FILLER_14_1177 ();
 sg13g2_fill_2 FILLER_14_1184 ();
 sg13g2_decap_4 FILLER_14_1191 ();
 sg13g2_fill_1 FILLER_14_1195 ();
 sg13g2_fill_2 FILLER_14_1200 ();
 sg13g2_decap_8 FILLER_14_1228 ();
 sg13g2_fill_1 FILLER_14_1235 ();
 sg13g2_fill_2 FILLER_14_1246 ();
 sg13g2_decap_8 FILLER_14_1264 ();
 sg13g2_decap_4 FILLER_14_1271 ();
 sg13g2_fill_2 FILLER_14_1275 ();
 sg13g2_decap_8 FILLER_14_1281 ();
 sg13g2_decap_8 FILLER_14_1288 ();
 sg13g2_decap_8 FILLER_14_1295 ();
 sg13g2_decap_8 FILLER_14_1302 ();
 sg13g2_fill_2 FILLER_14_1309 ();
 sg13g2_decap_8 FILLER_14_1315 ();
 sg13g2_fill_2 FILLER_14_1322 ();
 sg13g2_fill_1 FILLER_14_1324 ();
 sg13g2_decap_4 FILLER_14_1341 ();
 sg13g2_fill_2 FILLER_14_1345 ();
 sg13g2_decap_8 FILLER_14_1351 ();
 sg13g2_decap_8 FILLER_14_1358 ();
 sg13g2_decap_8 FILLER_14_1365 ();
 sg13g2_fill_1 FILLER_14_1372 ();
 sg13g2_decap_8 FILLER_14_1390 ();
 sg13g2_decap_8 FILLER_14_1397 ();
 sg13g2_decap_4 FILLER_14_1404 ();
 sg13g2_fill_2 FILLER_14_1408 ();
 sg13g2_decap_8 FILLER_14_1417 ();
 sg13g2_decap_8 FILLER_14_1424 ();
 sg13g2_fill_1 FILLER_14_1431 ();
 sg13g2_decap_8 FILLER_14_1437 ();
 sg13g2_decap_8 FILLER_14_1444 ();
 sg13g2_fill_1 FILLER_14_1451 ();
 sg13g2_decap_4 FILLER_14_1460 ();
 sg13g2_fill_2 FILLER_14_1464 ();
 sg13g2_decap_8 FILLER_14_1474 ();
 sg13g2_decap_8 FILLER_14_1481 ();
 sg13g2_decap_8 FILLER_14_1488 ();
 sg13g2_decap_8 FILLER_14_1543 ();
 sg13g2_fill_2 FILLER_14_1550 ();
 sg13g2_fill_1 FILLER_14_1556 ();
 sg13g2_decap_4 FILLER_14_1562 ();
 sg13g2_fill_2 FILLER_14_1566 ();
 sg13g2_fill_2 FILLER_14_1574 ();
 sg13g2_decap_8 FILLER_14_1582 ();
 sg13g2_fill_2 FILLER_14_1589 ();
 sg13g2_fill_1 FILLER_14_1591 ();
 sg13g2_fill_2 FILLER_14_1596 ();
 sg13g2_decap_8 FILLER_14_1609 ();
 sg13g2_fill_2 FILLER_14_1616 ();
 sg13g2_decap_8 FILLER_14_1640 ();
 sg13g2_decap_8 FILLER_14_1647 ();
 sg13g2_fill_1 FILLER_14_1654 ();
 sg13g2_fill_2 FILLER_14_1659 ();
 sg13g2_decap_8 FILLER_14_1674 ();
 sg13g2_decap_8 FILLER_14_1681 ();
 sg13g2_decap_8 FILLER_14_1688 ();
 sg13g2_decap_8 FILLER_14_1695 ();
 sg13g2_decap_8 FILLER_14_1702 ();
 sg13g2_decap_8 FILLER_14_1709 ();
 sg13g2_decap_8 FILLER_14_1716 ();
 sg13g2_decap_8 FILLER_14_1723 ();
 sg13g2_decap_8 FILLER_14_1730 ();
 sg13g2_decap_8 FILLER_14_1737 ();
 sg13g2_decap_8 FILLER_14_1744 ();
 sg13g2_decap_8 FILLER_14_1751 ();
 sg13g2_decap_8 FILLER_14_1758 ();
 sg13g2_decap_8 FILLER_14_1765 ();
 sg13g2_fill_2 FILLER_14_1772 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_4 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_4 FILLER_15_56 ();
 sg13g2_fill_2 FILLER_15_60 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_fill_2 FILLER_15_95 ();
 sg13g2_fill_1 FILLER_15_97 ();
 sg13g2_decap_4 FILLER_15_102 ();
 sg13g2_fill_2 FILLER_15_106 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_133 ();
 sg13g2_fill_1 FILLER_15_135 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_fill_2 FILLER_15_173 ();
 sg13g2_fill_1 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_188 ();
 sg13g2_decap_4 FILLER_15_195 ();
 sg13g2_fill_1 FILLER_15_199 ();
 sg13g2_decap_4 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_215 ();
 sg13g2_fill_2 FILLER_15_234 ();
 sg13g2_fill_2 FILLER_15_260 ();
 sg13g2_fill_1 FILLER_15_262 ();
 sg13g2_decap_4 FILLER_15_274 ();
 sg13g2_fill_2 FILLER_15_278 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_decap_4 FILLER_15_298 ();
 sg13g2_fill_2 FILLER_15_302 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_319 ();
 sg13g2_decap_4 FILLER_15_326 ();
 sg13g2_decap_4 FILLER_15_339 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_fill_2 FILLER_15_367 ();
 sg13g2_fill_1 FILLER_15_369 ();
 sg13g2_decap_4 FILLER_15_380 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_fill_2 FILLER_15_390 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_decap_8 FILLER_15_429 ();
 sg13g2_fill_1 FILLER_15_436 ();
 sg13g2_fill_1 FILLER_15_441 ();
 sg13g2_decap_4 FILLER_15_455 ();
 sg13g2_fill_2 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_467 ();
 sg13g2_decap_8 FILLER_15_474 ();
 sg13g2_decap_4 FILLER_15_481 ();
 sg13g2_fill_2 FILLER_15_490 ();
 sg13g2_fill_1 FILLER_15_492 ();
 sg13g2_decap_8 FILLER_15_501 ();
 sg13g2_decap_8 FILLER_15_508 ();
 sg13g2_decap_8 FILLER_15_515 ();
 sg13g2_decap_8 FILLER_15_522 ();
 sg13g2_decap_8 FILLER_15_529 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_decap_8 FILLER_15_564 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_fill_2 FILLER_15_578 ();
 sg13g2_fill_1 FILLER_15_580 ();
 sg13g2_decap_8 FILLER_15_607 ();
 sg13g2_fill_2 FILLER_15_614 ();
 sg13g2_fill_1 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_621 ();
 sg13g2_decap_8 FILLER_15_628 ();
 sg13g2_decap_8 FILLER_15_635 ();
 sg13g2_decap_8 FILLER_15_642 ();
 sg13g2_decap_8 FILLER_15_649 ();
 sg13g2_decap_8 FILLER_15_656 ();
 sg13g2_decap_4 FILLER_15_663 ();
 sg13g2_fill_1 FILLER_15_667 ();
 sg13g2_fill_2 FILLER_15_673 ();
 sg13g2_decap_4 FILLER_15_680 ();
 sg13g2_fill_2 FILLER_15_684 ();
 sg13g2_fill_1 FILLER_15_689 ();
 sg13g2_fill_1 FILLER_15_703 ();
 sg13g2_decap_8 FILLER_15_708 ();
 sg13g2_decap_8 FILLER_15_715 ();
 sg13g2_fill_2 FILLER_15_722 ();
 sg13g2_fill_2 FILLER_15_754 ();
 sg13g2_decap_8 FILLER_15_782 ();
 sg13g2_decap_8 FILLER_15_789 ();
 sg13g2_decap_8 FILLER_15_796 ();
 sg13g2_decap_8 FILLER_15_803 ();
 sg13g2_decap_8 FILLER_15_810 ();
 sg13g2_decap_8 FILLER_15_817 ();
 sg13g2_decap_8 FILLER_15_824 ();
 sg13g2_decap_8 FILLER_15_831 ();
 sg13g2_fill_2 FILLER_15_838 ();
 sg13g2_decap_8 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_851 ();
 sg13g2_decap_8 FILLER_15_858 ();
 sg13g2_fill_1 FILLER_15_865 ();
 sg13g2_decap_8 FILLER_15_895 ();
 sg13g2_decap_8 FILLER_15_902 ();
 sg13g2_fill_2 FILLER_15_909 ();
 sg13g2_fill_1 FILLER_15_911 ();
 sg13g2_decap_8 FILLER_15_916 ();
 sg13g2_decap_8 FILLER_15_923 ();
 sg13g2_decap_8 FILLER_15_930 ();
 sg13g2_fill_2 FILLER_15_937 ();
 sg13g2_decap_8 FILLER_15_954 ();
 sg13g2_decap_8 FILLER_15_961 ();
 sg13g2_fill_2 FILLER_15_968 ();
 sg13g2_decap_8 FILLER_15_989 ();
 sg13g2_decap_8 FILLER_15_1000 ();
 sg13g2_fill_1 FILLER_15_1007 ();
 sg13g2_decap_4 FILLER_15_1018 ();
 sg13g2_fill_1 FILLER_15_1022 ();
 sg13g2_fill_1 FILLER_15_1027 ();
 sg13g2_decap_8 FILLER_15_1044 ();
 sg13g2_fill_1 FILLER_15_1051 ();
 sg13g2_fill_2 FILLER_15_1061 ();
 sg13g2_fill_1 FILLER_15_1063 ();
 sg13g2_decap_8 FILLER_15_1098 ();
 sg13g2_decap_8 FILLER_15_1105 ();
 sg13g2_decap_8 FILLER_15_1112 ();
 sg13g2_fill_1 FILLER_15_1145 ();
 sg13g2_fill_1 FILLER_15_1160 ();
 sg13g2_decap_8 FILLER_15_1174 ();
 sg13g2_decap_8 FILLER_15_1181 ();
 sg13g2_decap_4 FILLER_15_1188 ();
 sg13g2_fill_2 FILLER_15_1192 ();
 sg13g2_fill_2 FILLER_15_1200 ();
 sg13g2_decap_4 FILLER_15_1220 ();
 sg13g2_fill_2 FILLER_15_1224 ();
 sg13g2_fill_2 FILLER_15_1231 ();
 sg13g2_fill_1 FILLER_15_1233 ();
 sg13g2_decap_8 FILLER_15_1237 ();
 sg13g2_decap_4 FILLER_15_1244 ();
 sg13g2_fill_2 FILLER_15_1248 ();
 sg13g2_decap_8 FILLER_15_1262 ();
 sg13g2_decap_8 FILLER_15_1269 ();
 sg13g2_decap_8 FILLER_15_1276 ();
 sg13g2_decap_8 FILLER_15_1283 ();
 sg13g2_decap_8 FILLER_15_1290 ();
 sg13g2_fill_2 FILLER_15_1297 ();
 sg13g2_fill_1 FILLER_15_1304 ();
 sg13g2_fill_2 FILLER_15_1308 ();
 sg13g2_fill_1 FILLER_15_1310 ();
 sg13g2_decap_8 FILLER_15_1345 ();
 sg13g2_decap_4 FILLER_15_1352 ();
 sg13g2_fill_2 FILLER_15_1356 ();
 sg13g2_decap_8 FILLER_15_1362 ();
 sg13g2_decap_4 FILLER_15_1369 ();
 sg13g2_fill_1 FILLER_15_1373 ();
 sg13g2_decap_8 FILLER_15_1393 ();
 sg13g2_decap_8 FILLER_15_1400 ();
 sg13g2_fill_1 FILLER_15_1407 ();
 sg13g2_decap_8 FILLER_15_1413 ();
 sg13g2_decap_8 FILLER_15_1420 ();
 sg13g2_decap_8 FILLER_15_1427 ();
 sg13g2_decap_8 FILLER_15_1439 ();
 sg13g2_decap_8 FILLER_15_1446 ();
 sg13g2_decap_8 FILLER_15_1453 ();
 sg13g2_fill_2 FILLER_15_1460 ();
 sg13g2_fill_1 FILLER_15_1462 ();
 sg13g2_decap_8 FILLER_15_1489 ();
 sg13g2_decap_4 FILLER_15_1496 ();
 sg13g2_fill_2 FILLER_15_1500 ();
 sg13g2_decap_4 FILLER_15_1549 ();
 sg13g2_fill_1 FILLER_15_1553 ();
 sg13g2_decap_8 FILLER_15_1560 ();
 sg13g2_decap_8 FILLER_15_1567 ();
 sg13g2_fill_1 FILLER_15_1574 ();
 sg13g2_decap_8 FILLER_15_1583 ();
 sg13g2_decap_8 FILLER_15_1590 ();
 sg13g2_fill_2 FILLER_15_1597 ();
 sg13g2_fill_1 FILLER_15_1599 ();
 sg13g2_decap_8 FILLER_15_1605 ();
 sg13g2_fill_2 FILLER_15_1612 ();
 sg13g2_decap_8 FILLER_15_1622 ();
 sg13g2_decap_4 FILLER_15_1629 ();
 sg13g2_fill_1 FILLER_15_1633 ();
 sg13g2_fill_2 FILLER_15_1639 ();
 sg13g2_decap_8 FILLER_15_1647 ();
 sg13g2_decap_8 FILLER_15_1654 ();
 sg13g2_fill_2 FILLER_15_1661 ();
 sg13g2_fill_1 FILLER_15_1663 ();
 sg13g2_fill_2 FILLER_15_1683 ();
 sg13g2_fill_1 FILLER_15_1685 ();
 sg13g2_decap_8 FILLER_15_1689 ();
 sg13g2_fill_2 FILLER_15_1696 ();
 sg13g2_decap_8 FILLER_15_1702 ();
 sg13g2_decap_8 FILLER_15_1709 ();
 sg13g2_decap_8 FILLER_15_1716 ();
 sg13g2_decap_8 FILLER_15_1723 ();
 sg13g2_decap_8 FILLER_15_1730 ();
 sg13g2_decap_8 FILLER_15_1737 ();
 sg13g2_decap_8 FILLER_15_1744 ();
 sg13g2_decap_8 FILLER_15_1751 ();
 sg13g2_decap_8 FILLER_15_1758 ();
 sg13g2_decap_8 FILLER_15_1765 ();
 sg13g2_fill_2 FILLER_15_1772 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_21 ();
 sg13g2_fill_1 FILLER_16_25 ();
 sg13g2_decap_4 FILLER_16_30 ();
 sg13g2_fill_1 FILLER_16_34 ();
 sg13g2_decap_4 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_53 ();
 sg13g2_fill_2 FILLER_16_58 ();
 sg13g2_fill_1 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_71 ();
 sg13g2_decap_8 FILLER_16_78 ();
 sg13g2_fill_2 FILLER_16_89 ();
 sg13g2_fill_1 FILLER_16_91 ();
 sg13g2_fill_2 FILLER_16_97 ();
 sg13g2_fill_1 FILLER_16_109 ();
 sg13g2_fill_2 FILLER_16_119 ();
 sg13g2_decap_4 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_131 ();
 sg13g2_fill_1 FILLER_16_141 ();
 sg13g2_fill_2 FILLER_16_157 ();
 sg13g2_decap_8 FILLER_16_173 ();
 sg13g2_fill_1 FILLER_16_180 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_4 FILLER_16_200 ();
 sg13g2_fill_2 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_fill_1 FILLER_16_218 ();
 sg13g2_decap_4 FILLER_16_224 ();
 sg13g2_fill_1 FILLER_16_228 ();
 sg13g2_decap_4 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_237 ();
 sg13g2_decap_8 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_250 ();
 sg13g2_decap_8 FILLER_16_257 ();
 sg13g2_decap_8 FILLER_16_264 ();
 sg13g2_decap_8 FILLER_16_271 ();
 sg13g2_decap_8 FILLER_16_285 ();
 sg13g2_decap_4 FILLER_16_292 ();
 sg13g2_fill_2 FILLER_16_296 ();
 sg13g2_decap_4 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_8 FILLER_16_360 ();
 sg13g2_decap_4 FILLER_16_367 ();
 sg13g2_fill_2 FILLER_16_371 ();
 sg13g2_fill_2 FILLER_16_396 ();
 sg13g2_fill_1 FILLER_16_398 ();
 sg13g2_decap_8 FILLER_16_404 ();
 sg13g2_decap_4 FILLER_16_411 ();
 sg13g2_decap_8 FILLER_16_425 ();
 sg13g2_decap_4 FILLER_16_432 ();
 sg13g2_fill_2 FILLER_16_436 ();
 sg13g2_decap_4 FILLER_16_456 ();
 sg13g2_fill_2 FILLER_16_460 ();
 sg13g2_decap_8 FILLER_16_502 ();
 sg13g2_decap_8 FILLER_16_509 ();
 sg13g2_decap_8 FILLER_16_516 ();
 sg13g2_fill_1 FILLER_16_523 ();
 sg13g2_fill_1 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_566 ();
 sg13g2_decap_4 FILLER_16_583 ();
 sg13g2_fill_2 FILLER_16_587 ();
 sg13g2_decap_8 FILLER_16_593 ();
 sg13g2_decap_8 FILLER_16_600 ();
 sg13g2_decap_8 FILLER_16_607 ();
 sg13g2_fill_2 FILLER_16_614 ();
 sg13g2_fill_2 FILLER_16_621 ();
 sg13g2_fill_2 FILLER_16_627 ();
 sg13g2_fill_1 FILLER_16_629 ();
 sg13g2_decap_8 FILLER_16_634 ();
 sg13g2_decap_8 FILLER_16_641 ();
 sg13g2_decap_8 FILLER_16_652 ();
 sg13g2_decap_4 FILLER_16_659 ();
 sg13g2_fill_1 FILLER_16_663 ();
 sg13g2_fill_2 FILLER_16_694 ();
 sg13g2_fill_1 FILLER_16_696 ();
 sg13g2_decap_8 FILLER_16_703 ();
 sg13g2_decap_4 FILLER_16_710 ();
 sg13g2_fill_1 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_725 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_decap_8 FILLER_16_753 ();
 sg13g2_decap_8 FILLER_16_760 ();
 sg13g2_decap_8 FILLER_16_767 ();
 sg13g2_decap_8 FILLER_16_774 ();
 sg13g2_decap_4 FILLER_16_781 ();
 sg13g2_fill_2 FILLER_16_785 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_4 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_838 ();
 sg13g2_fill_1 FILLER_16_845 ();
 sg13g2_decap_8 FILLER_16_856 ();
 sg13g2_fill_2 FILLER_16_863 ();
 sg13g2_fill_1 FILLER_16_865 ();
 sg13g2_decap_8 FILLER_16_869 ();
 sg13g2_fill_1 FILLER_16_876 ();
 sg13g2_decap_8 FILLER_16_881 ();
 sg13g2_decap_8 FILLER_16_888 ();
 sg13g2_decap_4 FILLER_16_895 ();
 sg13g2_fill_1 FILLER_16_899 ();
 sg13g2_decap_4 FILLER_16_934 ();
 sg13g2_fill_1 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_944 ();
 sg13g2_decap_8 FILLER_16_951 ();
 sg13g2_fill_2 FILLER_16_958 ();
 sg13g2_decap_8 FILLER_16_977 ();
 sg13g2_fill_1 FILLER_16_984 ();
 sg13g2_decap_8 FILLER_16_989 ();
 sg13g2_decap_8 FILLER_16_996 ();
 sg13g2_decap_4 FILLER_16_1022 ();
 sg13g2_fill_1 FILLER_16_1026 ();
 sg13g2_decap_8 FILLER_16_1049 ();
 sg13g2_decap_8 FILLER_16_1056 ();
 sg13g2_decap_8 FILLER_16_1063 ();
 sg13g2_fill_2 FILLER_16_1070 ();
 sg13g2_fill_1 FILLER_16_1072 ();
 sg13g2_decap_8 FILLER_16_1077 ();
 sg13g2_decap_8 FILLER_16_1084 ();
 sg13g2_decap_8 FILLER_16_1091 ();
 sg13g2_fill_2 FILLER_16_1098 ();
 sg13g2_decap_8 FILLER_16_1105 ();
 sg13g2_decap_4 FILLER_16_1112 ();
 sg13g2_fill_2 FILLER_16_1125 ();
 sg13g2_decap_8 FILLER_16_1140 ();
 sg13g2_decap_8 FILLER_16_1147 ();
 sg13g2_fill_1 FILLER_16_1154 ();
 sg13g2_fill_2 FILLER_16_1181 ();
 sg13g2_fill_1 FILLER_16_1183 ();
 sg13g2_decap_4 FILLER_16_1188 ();
 sg13g2_fill_2 FILLER_16_1192 ();
 sg13g2_decap_4 FILLER_16_1204 ();
 sg13g2_fill_1 FILLER_16_1208 ();
 sg13g2_decap_8 FILLER_16_1217 ();
 sg13g2_decap_8 FILLER_16_1224 ();
 sg13g2_fill_1 FILLER_16_1231 ();
 sg13g2_fill_2 FILLER_16_1264 ();
 sg13g2_fill_1 FILLER_16_1266 ();
 sg13g2_decap_8 FILLER_16_1271 ();
 sg13g2_fill_2 FILLER_16_1278 ();
 sg13g2_fill_1 FILLER_16_1280 ();
 sg13g2_decap_4 FILLER_16_1286 ();
 sg13g2_fill_2 FILLER_16_1290 ();
 sg13g2_decap_8 FILLER_16_1295 ();
 sg13g2_fill_1 FILLER_16_1317 ();
 sg13g2_decap_8 FILLER_16_1323 ();
 sg13g2_decap_8 FILLER_16_1330 ();
 sg13g2_fill_1 FILLER_16_1356 ();
 sg13g2_decap_8 FILLER_16_1362 ();
 sg13g2_decap_8 FILLER_16_1369 ();
 sg13g2_fill_1 FILLER_16_1376 ();
 sg13g2_fill_1 FILLER_16_1407 ();
 sg13g2_fill_2 FILLER_16_1416 ();
 sg13g2_fill_2 FILLER_16_1421 ();
 sg13g2_decap_8 FILLER_16_1431 ();
 sg13g2_decap_4 FILLER_16_1438 ();
 sg13g2_decap_8 FILLER_16_1446 ();
 sg13g2_decap_8 FILLER_16_1453 ();
 sg13g2_decap_8 FILLER_16_1460 ();
 sg13g2_decap_8 FILLER_16_1467 ();
 sg13g2_decap_8 FILLER_16_1474 ();
 sg13g2_decap_8 FILLER_16_1481 ();
 sg13g2_decap_8 FILLER_16_1488 ();
 sg13g2_decap_8 FILLER_16_1495 ();
 sg13g2_decap_4 FILLER_16_1502 ();
 sg13g2_fill_1 FILLER_16_1523 ();
 sg13g2_decap_4 FILLER_16_1534 ();
 sg13g2_decap_8 FILLER_16_1549 ();
 sg13g2_decap_8 FILLER_16_1556 ();
 sg13g2_decap_8 FILLER_16_1563 ();
 sg13g2_decap_4 FILLER_16_1570 ();
 sg13g2_fill_2 FILLER_16_1574 ();
 sg13g2_decap_4 FILLER_16_1581 ();
 sg13g2_fill_2 FILLER_16_1585 ();
 sg13g2_decap_8 FILLER_16_1593 ();
 sg13g2_fill_1 FILLER_16_1600 ();
 sg13g2_fill_1 FILLER_16_1607 ();
 sg13g2_fill_1 FILLER_16_1613 ();
 sg13g2_fill_1 FILLER_16_1619 ();
 sg13g2_fill_1 FILLER_16_1631 ();
 sg13g2_decap_8 FILLER_16_1636 ();
 sg13g2_decap_8 FILLER_16_1643 ();
 sg13g2_decap_8 FILLER_16_1650 ();
 sg13g2_decap_8 FILLER_16_1657 ();
 sg13g2_decap_8 FILLER_16_1664 ();
 sg13g2_decap_4 FILLER_16_1671 ();
 sg13g2_fill_2 FILLER_16_1675 ();
 sg13g2_fill_1 FILLER_16_1680 ();
 sg13g2_fill_2 FILLER_16_1689 ();
 sg13g2_decap_8 FILLER_16_1717 ();
 sg13g2_decap_8 FILLER_16_1724 ();
 sg13g2_decap_8 FILLER_16_1731 ();
 sg13g2_decap_8 FILLER_16_1738 ();
 sg13g2_decap_8 FILLER_16_1745 ();
 sg13g2_decap_8 FILLER_16_1752 ();
 sg13g2_decap_8 FILLER_16_1759 ();
 sg13g2_decap_8 FILLER_16_1766 ();
 sg13g2_fill_1 FILLER_16_1773 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_4 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_39 ();
 sg13g2_fill_2 FILLER_17_49 ();
 sg13g2_fill_1 FILLER_17_51 ();
 sg13g2_fill_2 FILLER_17_57 ();
 sg13g2_fill_2 FILLER_17_76 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_fill_1 FILLER_17_89 ();
 sg13g2_fill_1 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_fill_2 FILLER_17_113 ();
 sg13g2_fill_1 FILLER_17_115 ();
 sg13g2_decap_8 FILLER_17_121 ();
 sg13g2_decap_8 FILLER_17_128 ();
 sg13g2_fill_2 FILLER_17_135 ();
 sg13g2_decap_4 FILLER_17_142 ();
 sg13g2_fill_1 FILLER_17_146 ();
 sg13g2_decap_4 FILLER_17_153 ();
 sg13g2_fill_2 FILLER_17_162 ();
 sg13g2_decap_4 FILLER_17_169 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_fill_2 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_4 FILLER_17_245 ();
 sg13g2_fill_1 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_274 ();
 sg13g2_decap_8 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_317 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_4 FILLER_17_331 ();
 sg13g2_fill_2 FILLER_17_335 ();
 sg13g2_fill_2 FILLER_17_341 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_fill_1 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_4 FILLER_17_377 ();
 sg13g2_fill_1 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_fill_1 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_426 ();
 sg13g2_fill_1 FILLER_17_433 ();
 sg13g2_decap_4 FILLER_17_438 ();
 sg13g2_fill_1 FILLER_17_442 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_fill_2 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_496 ();
 sg13g2_decap_8 FILLER_17_503 ();
 sg13g2_decap_4 FILLER_17_510 ();
 sg13g2_fill_2 FILLER_17_514 ();
 sg13g2_fill_1 FILLER_17_520 ();
 sg13g2_fill_2 FILLER_17_542 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_fill_2 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_568 ();
 sg13g2_decap_8 FILLER_17_575 ();
 sg13g2_decap_4 FILLER_17_582 ();
 sg13g2_decap_8 FILLER_17_615 ();
 sg13g2_decap_8 FILLER_17_653 ();
 sg13g2_decap_8 FILLER_17_660 ();
 sg13g2_decap_4 FILLER_17_667 ();
 sg13g2_decap_8 FILLER_17_675 ();
 sg13g2_decap_8 FILLER_17_682 ();
 sg13g2_decap_8 FILLER_17_689 ();
 sg13g2_decap_4 FILLER_17_696 ();
 sg13g2_fill_2 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_705 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_739 ();
 sg13g2_decap_8 FILLER_17_746 ();
 sg13g2_decap_8 FILLER_17_753 ();
 sg13g2_decap_8 FILLER_17_760 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_decap_8 FILLER_17_818 ();
 sg13g2_decap_8 FILLER_17_825 ();
 sg13g2_fill_1 FILLER_17_832 ();
 sg13g2_fill_1 FILLER_17_846 ();
 sg13g2_fill_2 FILLER_17_864 ();
 sg13g2_fill_1 FILLER_17_878 ();
 sg13g2_decap_8 FILLER_17_883 ();
 sg13g2_decap_8 FILLER_17_890 ();
 sg13g2_decap_8 FILLER_17_897 ();
 sg13g2_fill_1 FILLER_17_904 ();
 sg13g2_decap_8 FILLER_17_908 ();
 sg13g2_decap_8 FILLER_17_915 ();
 sg13g2_fill_2 FILLER_17_922 ();
 sg13g2_fill_1 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_17_933 ();
 sg13g2_decap_8 FILLER_17_940 ();
 sg13g2_decap_8 FILLER_17_947 ();
 sg13g2_fill_2 FILLER_17_954 ();
 sg13g2_fill_1 FILLER_17_956 ();
 sg13g2_fill_2 FILLER_17_1014 ();
 sg13g2_fill_1 FILLER_17_1041 ();
 sg13g2_decap_8 FILLER_17_1073 ();
 sg13g2_fill_2 FILLER_17_1088 ();
 sg13g2_fill_1 FILLER_17_1090 ();
 sg13g2_decap_4 FILLER_17_1110 ();
 sg13g2_fill_1 FILLER_17_1125 ();
 sg13g2_decap_8 FILLER_17_1152 ();
 sg13g2_decap_4 FILLER_17_1159 ();
 sg13g2_fill_1 FILLER_17_1175 ();
 sg13g2_decap_8 FILLER_17_1186 ();
 sg13g2_decap_8 FILLER_17_1193 ();
 sg13g2_decap_8 FILLER_17_1200 ();
 sg13g2_decap_8 FILLER_17_1207 ();
 sg13g2_decap_4 FILLER_17_1218 ();
 sg13g2_fill_1 FILLER_17_1222 ();
 sg13g2_decap_4 FILLER_17_1226 ();
 sg13g2_fill_2 FILLER_17_1230 ();
 sg13g2_fill_1 FILLER_17_1236 ();
 sg13g2_fill_1 FILLER_17_1259 ();
 sg13g2_decap_4 FILLER_17_1264 ();
 sg13g2_fill_1 FILLER_17_1268 ();
 sg13g2_fill_1 FILLER_17_1283 ();
 sg13g2_fill_1 FILLER_17_1296 ();
 sg13g2_decap_4 FILLER_17_1313 ();
 sg13g2_decap_8 FILLER_17_1327 ();
 sg13g2_decap_8 FILLER_17_1334 ();
 sg13g2_fill_2 FILLER_17_1341 ();
 sg13g2_decap_8 FILLER_17_1353 ();
 sg13g2_decap_8 FILLER_17_1360 ();
 sg13g2_decap_8 FILLER_17_1372 ();
 sg13g2_decap_8 FILLER_17_1379 ();
 sg13g2_decap_8 FILLER_17_1386 ();
 sg13g2_decap_8 FILLER_17_1393 ();
 sg13g2_decap_8 FILLER_17_1400 ();
 sg13g2_decap_8 FILLER_17_1407 ();
 sg13g2_fill_1 FILLER_17_1414 ();
 sg13g2_decap_8 FILLER_17_1460 ();
 sg13g2_decap_8 FILLER_17_1472 ();
 sg13g2_decap_8 FILLER_17_1479 ();
 sg13g2_decap_8 FILLER_17_1486 ();
 sg13g2_decap_4 FILLER_17_1493 ();
 sg13g2_fill_2 FILLER_17_1497 ();
 sg13g2_decap_8 FILLER_17_1511 ();
 sg13g2_fill_2 FILLER_17_1518 ();
 sg13g2_fill_1 FILLER_17_1520 ();
 sg13g2_fill_2 FILLER_17_1527 ();
 sg13g2_fill_1 FILLER_17_1529 ();
 sg13g2_fill_1 FILLER_17_1537 ();
 sg13g2_fill_1 FILLER_17_1542 ();
 sg13g2_decap_8 FILLER_17_1547 ();
 sg13g2_decap_8 FILLER_17_1554 ();
 sg13g2_decap_8 FILLER_17_1561 ();
 sg13g2_decap_8 FILLER_17_1568 ();
 sg13g2_fill_1 FILLER_17_1575 ();
 sg13g2_decap_8 FILLER_17_1581 ();
 sg13g2_decap_8 FILLER_17_1588 ();
 sg13g2_decap_8 FILLER_17_1595 ();
 sg13g2_decap_4 FILLER_17_1602 ();
 sg13g2_fill_2 FILLER_17_1606 ();
 sg13g2_fill_2 FILLER_17_1611 ();
 sg13g2_fill_2 FILLER_17_1636 ();
 sg13g2_decap_4 FILLER_17_1646 ();
 sg13g2_decap_4 FILLER_17_1655 ();
 sg13g2_decap_8 FILLER_17_1667 ();
 sg13g2_fill_1 FILLER_17_1684 ();
 sg13g2_fill_1 FILLER_17_1688 ();
 sg13g2_decap_8 FILLER_17_1700 ();
 sg13g2_decap_8 FILLER_17_1707 ();
 sg13g2_fill_2 FILLER_17_1714 ();
 sg13g2_decap_8 FILLER_17_1720 ();
 sg13g2_decap_8 FILLER_17_1727 ();
 sg13g2_decap_8 FILLER_17_1734 ();
 sg13g2_decap_8 FILLER_17_1741 ();
 sg13g2_decap_8 FILLER_17_1748 ();
 sg13g2_decap_8 FILLER_17_1755 ();
 sg13g2_decap_8 FILLER_17_1762 ();
 sg13g2_decap_4 FILLER_17_1769 ();
 sg13g2_fill_1 FILLER_17_1773 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_fill_2 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_41 ();
 sg13g2_fill_1 FILLER_18_46 ();
 sg13g2_decap_4 FILLER_18_51 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_66 ();
 sg13g2_fill_1 FILLER_18_68 ();
 sg13g2_decap_4 FILLER_18_74 ();
 sg13g2_fill_2 FILLER_18_78 ();
 sg13g2_fill_1 FILLER_18_90 ();
 sg13g2_decap_4 FILLER_18_97 ();
 sg13g2_fill_2 FILLER_18_101 ();
 sg13g2_decap_8 FILLER_18_114 ();
 sg13g2_fill_2 FILLER_18_126 ();
 sg13g2_fill_2 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_135 ();
 sg13g2_decap_4 FILLER_18_146 ();
 sg13g2_fill_1 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_160 ();
 sg13g2_decap_4 FILLER_18_172 ();
 sg13g2_fill_2 FILLER_18_176 ();
 sg13g2_decap_4 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_202 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_223 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_fill_2 FILLER_18_241 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_254 ();
 sg13g2_decap_8 FILLER_18_274 ();
 sg13g2_decap_8 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_288 ();
 sg13g2_fill_2 FILLER_18_295 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_2 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_4 FILLER_18_341 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_decap_4 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_4 FILLER_18_387 ();
 sg13g2_fill_2 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_fill_2 FILLER_18_404 ();
 sg13g2_decap_4 FILLER_18_421 ();
 sg13g2_fill_2 FILLER_18_425 ();
 sg13g2_decap_8 FILLER_18_432 ();
 sg13g2_decap_4 FILLER_18_439 ();
 sg13g2_decap_4 FILLER_18_447 ();
 sg13g2_fill_2 FILLER_18_451 ();
 sg13g2_decap_8 FILLER_18_458 ();
 sg13g2_decap_8 FILLER_18_465 ();
 sg13g2_fill_1 FILLER_18_472 ();
 sg13g2_decap_8 FILLER_18_481 ();
 sg13g2_decap_8 FILLER_18_498 ();
 sg13g2_decap_8 FILLER_18_505 ();
 sg13g2_decap_4 FILLER_18_512 ();
 sg13g2_fill_1 FILLER_18_516 ();
 sg13g2_decap_4 FILLER_18_521 ();
 sg13g2_fill_1 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_530 ();
 sg13g2_decap_8 FILLER_18_537 ();
 sg13g2_decap_8 FILLER_18_544 ();
 sg13g2_decap_8 FILLER_18_551 ();
 sg13g2_decap_8 FILLER_18_558 ();
 sg13g2_decap_8 FILLER_18_565 ();
 sg13g2_decap_8 FILLER_18_572 ();
 sg13g2_decap_8 FILLER_18_605 ();
 sg13g2_decap_8 FILLER_18_612 ();
 sg13g2_fill_2 FILLER_18_619 ();
 sg13g2_fill_1 FILLER_18_621 ();
 sg13g2_decap_8 FILLER_18_626 ();
 sg13g2_decap_8 FILLER_18_633 ();
 sg13g2_decap_4 FILLER_18_640 ();
 sg13g2_decap_8 FILLER_18_648 ();
 sg13g2_decap_4 FILLER_18_655 ();
 sg13g2_fill_1 FILLER_18_659 ();
 sg13g2_fill_2 FILLER_18_664 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_4 FILLER_18_693 ();
 sg13g2_fill_2 FILLER_18_697 ();
 sg13g2_decap_8 FILLER_18_708 ();
 sg13g2_fill_1 FILLER_18_715 ();
 sg13g2_decap_4 FILLER_18_720 ();
 sg13g2_fill_1 FILLER_18_724 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_fill_2 FILLER_18_777 ();
 sg13g2_fill_1 FILLER_18_779 ();
 sg13g2_decap_4 FILLER_18_784 ();
 sg13g2_fill_1 FILLER_18_788 ();
 sg13g2_decap_4 FILLER_18_792 ();
 sg13g2_fill_2 FILLER_18_796 ();
 sg13g2_decap_8 FILLER_18_802 ();
 sg13g2_decap_8 FILLER_18_809 ();
 sg13g2_decap_4 FILLER_18_816 ();
 sg13g2_fill_2 FILLER_18_820 ();
 sg13g2_fill_2 FILLER_18_835 ();
 sg13g2_decap_4 FILLER_18_841 ();
 sg13g2_fill_1 FILLER_18_845 ();
 sg13g2_fill_2 FILLER_18_858 ();
 sg13g2_decap_8 FILLER_18_898 ();
 sg13g2_decap_8 FILLER_18_910 ();
 sg13g2_decap_4 FILLER_18_921 ();
 sg13g2_decap_8 FILLER_18_928 ();
 sg13g2_decap_8 FILLER_18_935 ();
 sg13g2_decap_8 FILLER_18_942 ();
 sg13g2_decap_4 FILLER_18_949 ();
 sg13g2_fill_2 FILLER_18_962 ();
 sg13g2_fill_1 FILLER_18_964 ();
 sg13g2_decap_8 FILLER_18_970 ();
 sg13g2_fill_2 FILLER_18_977 ();
 sg13g2_fill_1 FILLER_18_979 ();
 sg13g2_decap_8 FILLER_18_988 ();
 sg13g2_decap_8 FILLER_18_995 ();
 sg13g2_decap_4 FILLER_18_1002 ();
 sg13g2_fill_2 FILLER_18_1006 ();
 sg13g2_fill_2 FILLER_18_1048 ();
 sg13g2_decap_8 FILLER_18_1058 ();
 sg13g2_decap_8 FILLER_18_1065 ();
 sg13g2_decap_8 FILLER_18_1072 ();
 sg13g2_decap_8 FILLER_18_1079 ();
 sg13g2_decap_8 FILLER_18_1086 ();
 sg13g2_fill_2 FILLER_18_1093 ();
 sg13g2_fill_1 FILLER_18_1095 ();
 sg13g2_fill_2 FILLER_18_1100 ();
 sg13g2_decap_8 FILLER_18_1106 ();
 sg13g2_fill_2 FILLER_18_1113 ();
 sg13g2_fill_1 FILLER_18_1115 ();
 sg13g2_decap_8 FILLER_18_1123 ();
 sg13g2_fill_1 FILLER_18_1130 ();
 sg13g2_decap_8 FILLER_18_1139 ();
 sg13g2_decap_8 FILLER_18_1146 ();
 sg13g2_decap_8 FILLER_18_1153 ();
 sg13g2_decap_8 FILLER_18_1195 ();
 sg13g2_decap_8 FILLER_18_1202 ();
 sg13g2_decap_8 FILLER_18_1209 ();
 sg13g2_decap_8 FILLER_18_1216 ();
 sg13g2_decap_8 FILLER_18_1223 ();
 sg13g2_fill_2 FILLER_18_1230 ();
 sg13g2_fill_1 FILLER_18_1248 ();
 sg13g2_decap_8 FILLER_18_1257 ();
 sg13g2_decap_4 FILLER_18_1264 ();
 sg13g2_fill_1 FILLER_18_1268 ();
 sg13g2_decap_8 FILLER_18_1274 ();
 sg13g2_decap_8 FILLER_18_1281 ();
 sg13g2_decap_8 FILLER_18_1288 ();
 sg13g2_decap_8 FILLER_18_1295 ();
 sg13g2_fill_1 FILLER_18_1302 ();
 sg13g2_decap_8 FILLER_18_1314 ();
 sg13g2_decap_8 FILLER_18_1326 ();
 sg13g2_decap_4 FILLER_18_1333 ();
 sg13g2_fill_2 FILLER_18_1337 ();
 sg13g2_fill_2 FILLER_18_1349 ();
 sg13g2_fill_1 FILLER_18_1351 ();
 sg13g2_decap_8 FILLER_18_1361 ();
 sg13g2_fill_1 FILLER_18_1368 ();
 sg13g2_decap_4 FILLER_18_1373 ();
 sg13g2_fill_2 FILLER_18_1377 ();
 sg13g2_fill_1 FILLER_18_1401 ();
 sg13g2_decap_8 FILLER_18_1412 ();
 sg13g2_decap_8 FILLER_18_1419 ();
 sg13g2_decap_8 FILLER_18_1426 ();
 sg13g2_decap_4 FILLER_18_1433 ();
 sg13g2_fill_2 FILLER_18_1437 ();
 sg13g2_decap_4 FILLER_18_1443 ();
 sg13g2_fill_1 FILLER_18_1447 ();
 sg13g2_decap_8 FILLER_18_1453 ();
 sg13g2_decap_8 FILLER_18_1460 ();
 sg13g2_decap_8 FILLER_18_1467 ();
 sg13g2_decap_8 FILLER_18_1474 ();
 sg13g2_decap_8 FILLER_18_1481 ();
 sg13g2_decap_8 FILLER_18_1488 ();
 sg13g2_decap_8 FILLER_18_1495 ();
 sg13g2_decap_4 FILLER_18_1502 ();
 sg13g2_decap_4 FILLER_18_1515 ();
 sg13g2_fill_2 FILLER_18_1519 ();
 sg13g2_decap_4 FILLER_18_1524 ();
 sg13g2_fill_2 FILLER_18_1528 ();
 sg13g2_fill_2 FILLER_18_1535 ();
 sg13g2_fill_1 FILLER_18_1537 ();
 sg13g2_decap_8 FILLER_18_1554 ();
 sg13g2_fill_1 FILLER_18_1561 ();
 sg13g2_decap_8 FILLER_18_1567 ();
 sg13g2_fill_1 FILLER_18_1574 ();
 sg13g2_fill_1 FILLER_18_1588 ();
 sg13g2_fill_2 FILLER_18_1619 ();
 sg13g2_fill_2 FILLER_18_1626 ();
 sg13g2_fill_1 FILLER_18_1632 ();
 sg13g2_decap_8 FILLER_18_1636 ();
 sg13g2_decap_8 FILLER_18_1643 ();
 sg13g2_decap_8 FILLER_18_1650 ();
 sg13g2_decap_8 FILLER_18_1657 ();
 sg13g2_decap_8 FILLER_18_1664 ();
 sg13g2_fill_2 FILLER_18_1680 ();
 sg13g2_fill_1 FILLER_18_1689 ();
 sg13g2_decap_4 FILLER_18_1703 ();
 sg13g2_fill_2 FILLER_18_1707 ();
 sg13g2_decap_8 FILLER_18_1735 ();
 sg13g2_decap_8 FILLER_18_1742 ();
 sg13g2_decap_8 FILLER_18_1749 ();
 sg13g2_decap_8 FILLER_18_1756 ();
 sg13g2_decap_8 FILLER_18_1763 ();
 sg13g2_decap_4 FILLER_18_1770 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_4 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_48 ();
 sg13g2_fill_1 FILLER_19_52 ();
 sg13g2_decap_4 FILLER_19_58 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_fill_2 FILLER_19_75 ();
 sg13g2_decap_4 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_85 ();
 sg13g2_fill_2 FILLER_19_91 ();
 sg13g2_fill_2 FILLER_19_112 ();
 sg13g2_fill_1 FILLER_19_114 ();
 sg13g2_decap_8 FILLER_19_134 ();
 sg13g2_fill_2 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_148 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_fill_2 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_171 ();
 sg13g2_decap_4 FILLER_19_183 ();
 sg13g2_fill_1 FILLER_19_187 ();
 sg13g2_decap_4 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_230 ();
 sg13g2_fill_2 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_251 ();
 sg13g2_decap_4 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_262 ();
 sg13g2_decap_4 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_273 ();
 sg13g2_decap_4 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_decap_4 FILLER_19_289 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_decap_4 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_329 ();
 sg13g2_fill_2 FILLER_19_336 ();
 sg13g2_decap_4 FILLER_19_342 ();
 sg13g2_decap_4 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_355 ();
 sg13g2_fill_1 FILLER_19_361 ();
 sg13g2_decap_4 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_4 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_4 FILLER_19_455 ();
 sg13g2_fill_1 FILLER_19_459 ();
 sg13g2_decap_8 FILLER_19_465 ();
 sg13g2_fill_2 FILLER_19_482 ();
 sg13g2_fill_2 FILLER_19_488 ();
 sg13g2_fill_1 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_499 ();
 sg13g2_decap_8 FILLER_19_506 ();
 sg13g2_decap_8 FILLER_19_513 ();
 sg13g2_decap_8 FILLER_19_520 ();
 sg13g2_decap_8 FILLER_19_527 ();
 sg13g2_decap_8 FILLER_19_534 ();
 sg13g2_fill_2 FILLER_19_541 ();
 sg13g2_decap_4 FILLER_19_549 ();
 sg13g2_fill_2 FILLER_19_553 ();
 sg13g2_decap_4 FILLER_19_561 ();
 sg13g2_fill_2 FILLER_19_565 ();
 sg13g2_decap_4 FILLER_19_570 ();
 sg13g2_fill_2 FILLER_19_574 ();
 sg13g2_decap_4 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_641 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_4 FILLER_19_700 ();
 sg13g2_fill_2 FILLER_19_704 ();
 sg13g2_decap_8 FILLER_19_712 ();
 sg13g2_decap_4 FILLER_19_723 ();
 sg13g2_fill_1 FILLER_19_727 ();
 sg13g2_decap_8 FILLER_19_732 ();
 sg13g2_decap_4 FILLER_19_739 ();
 sg13g2_fill_2 FILLER_19_743 ();
 sg13g2_decap_8 FILLER_19_748 ();
 sg13g2_decap_4 FILLER_19_755 ();
 sg13g2_fill_1 FILLER_19_759 ();
 sg13g2_decap_8 FILLER_19_764 ();
 sg13g2_decap_4 FILLER_19_771 ();
 sg13g2_fill_1 FILLER_19_775 ();
 sg13g2_decap_4 FILLER_19_788 ();
 sg13g2_fill_1 FILLER_19_805 ();
 sg13g2_fill_1 FILLER_19_810 ();
 sg13g2_decap_8 FILLER_19_816 ();
 sg13g2_decap_4 FILLER_19_823 ();
 sg13g2_fill_2 FILLER_19_827 ();
 sg13g2_decap_8 FILLER_19_834 ();
 sg13g2_fill_1 FILLER_19_841 ();
 sg13g2_decap_8 FILLER_19_876 ();
 sg13g2_fill_1 FILLER_19_883 ();
 sg13g2_decap_8 FILLER_19_889 ();
 sg13g2_decap_8 FILLER_19_896 ();
 sg13g2_decap_4 FILLER_19_903 ();
 sg13g2_fill_2 FILLER_19_907 ();
 sg13g2_decap_8 FILLER_19_935 ();
 sg13g2_decap_8 FILLER_19_942 ();
 sg13g2_decap_8 FILLER_19_949 ();
 sg13g2_fill_2 FILLER_19_956 ();
 sg13g2_fill_1 FILLER_19_958 ();
 sg13g2_decap_8 FILLER_19_989 ();
 sg13g2_decap_8 FILLER_19_996 ();
 sg13g2_fill_1 FILLER_19_1003 ();
 sg13g2_fill_2 FILLER_19_1013 ();
 sg13g2_decap_8 FILLER_19_1020 ();
 sg13g2_decap_8 FILLER_19_1027 ();
 sg13g2_decap_4 FILLER_19_1034 ();
 sg13g2_fill_2 FILLER_19_1038 ();
 sg13g2_decap_8 FILLER_19_1044 ();
 sg13g2_decap_8 FILLER_19_1051 ();
 sg13g2_decap_8 FILLER_19_1058 ();
 sg13g2_fill_2 FILLER_19_1070 ();
 sg13g2_decap_8 FILLER_19_1081 ();
 sg13g2_decap_8 FILLER_19_1088 ();
 sg13g2_decap_4 FILLER_19_1095 ();
 sg13g2_decap_4 FILLER_19_1104 ();
 sg13g2_fill_1 FILLER_19_1108 ();
 sg13g2_decap_8 FILLER_19_1116 ();
 sg13g2_decap_4 FILLER_19_1123 ();
 sg13g2_fill_1 FILLER_19_1127 ();
 sg13g2_decap_8 FILLER_19_1133 ();
 sg13g2_fill_2 FILLER_19_1140 ();
 sg13g2_fill_1 FILLER_19_1142 ();
 sg13g2_fill_2 FILLER_19_1147 ();
 sg13g2_decap_8 FILLER_19_1154 ();
 sg13g2_decap_8 FILLER_19_1161 ();
 sg13g2_decap_8 FILLER_19_1168 ();
 sg13g2_fill_2 FILLER_19_1175 ();
 sg13g2_decap_8 FILLER_19_1227 ();
 sg13g2_decap_4 FILLER_19_1234 ();
 sg13g2_fill_2 FILLER_19_1238 ();
 sg13g2_decap_4 FILLER_19_1254 ();
 sg13g2_fill_1 FILLER_19_1258 ();
 sg13g2_decap_4 FILLER_19_1263 ();
 sg13g2_fill_2 FILLER_19_1267 ();
 sg13g2_decap_8 FILLER_19_1279 ();
 sg13g2_decap_8 FILLER_19_1315 ();
 sg13g2_decap_8 FILLER_19_1322 ();
 sg13g2_decap_8 FILLER_19_1329 ();
 sg13g2_decap_4 FILLER_19_1336 ();
 sg13g2_fill_2 FILLER_19_1340 ();
 sg13g2_decap_8 FILLER_19_1358 ();
 sg13g2_decap_4 FILLER_19_1365 ();
 sg13g2_fill_2 FILLER_19_1395 ();
 sg13g2_decap_8 FILLER_19_1401 ();
 sg13g2_decap_8 FILLER_19_1408 ();
 sg13g2_decap_8 FILLER_19_1415 ();
 sg13g2_decap_8 FILLER_19_1422 ();
 sg13g2_decap_4 FILLER_19_1429 ();
 sg13g2_fill_2 FILLER_19_1433 ();
 sg13g2_fill_1 FILLER_19_1445 ();
 sg13g2_decap_8 FILLER_19_1454 ();
 sg13g2_fill_2 FILLER_19_1461 ();
 sg13g2_fill_1 FILLER_19_1463 ();
 sg13g2_decap_8 FILLER_19_1468 ();
 sg13g2_decap_8 FILLER_19_1475 ();
 sg13g2_decap_8 FILLER_19_1482 ();
 sg13g2_fill_2 FILLER_19_1501 ();
 sg13g2_fill_2 FILLER_19_1540 ();
 sg13g2_decap_4 FILLER_19_1547 ();
 sg13g2_fill_2 FILLER_19_1551 ();
 sg13g2_decap_8 FILLER_19_1557 ();
 sg13g2_decap_8 FILLER_19_1564 ();
 sg13g2_decap_8 FILLER_19_1571 ();
 sg13g2_decap_8 FILLER_19_1578 ();
 sg13g2_decap_4 FILLER_19_1585 ();
 sg13g2_fill_2 FILLER_19_1589 ();
 sg13g2_fill_2 FILLER_19_1595 ();
 sg13g2_fill_1 FILLER_19_1597 ();
 sg13g2_decap_4 FILLER_19_1601 ();
 sg13g2_fill_1 FILLER_19_1605 ();
 sg13g2_fill_2 FILLER_19_1626 ();
 sg13g2_fill_1 FILLER_19_1628 ();
 sg13g2_decap_8 FILLER_19_1634 ();
 sg13g2_decap_8 FILLER_19_1641 ();
 sg13g2_fill_1 FILLER_19_1648 ();
 sg13g2_fill_2 FILLER_19_1656 ();
 sg13g2_fill_1 FILLER_19_1658 ();
 sg13g2_fill_2 FILLER_19_1664 ();
 sg13g2_fill_1 FILLER_19_1681 ();
 sg13g2_decap_4 FILLER_19_1700 ();
 sg13g2_fill_2 FILLER_19_1704 ();
 sg13g2_decap_8 FILLER_19_1719 ();
 sg13g2_decap_8 FILLER_19_1726 ();
 sg13g2_decap_8 FILLER_19_1733 ();
 sg13g2_decap_8 FILLER_19_1740 ();
 sg13g2_decap_8 FILLER_19_1747 ();
 sg13g2_decap_8 FILLER_19_1754 ();
 sg13g2_decap_8 FILLER_19_1761 ();
 sg13g2_decap_4 FILLER_19_1768 ();
 sg13g2_fill_2 FILLER_19_1772 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_decap_4 FILLER_20_44 ();
 sg13g2_fill_1 FILLER_20_48 ();
 sg13g2_fill_2 FILLER_20_54 ();
 sg13g2_fill_1 FILLER_20_56 ();
 sg13g2_decap_4 FILLER_20_61 ();
 sg13g2_decap_4 FILLER_20_69 ();
 sg13g2_fill_2 FILLER_20_73 ();
 sg13g2_decap_4 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_85 ();
 sg13g2_decap_4 FILLER_20_91 ();
 sg13g2_fill_2 FILLER_20_95 ();
 sg13g2_fill_1 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_116 ();
 sg13g2_fill_2 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_143 ();
 sg13g2_decap_4 FILLER_20_150 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_decap_4 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_194 ();
 sg13g2_decap_8 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_211 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_fill_2 FILLER_20_230 ();
 sg13g2_decap_8 FILLER_20_236 ();
 sg13g2_decap_8 FILLER_20_243 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_fill_2 FILLER_20_271 ();
 sg13g2_fill_1 FILLER_20_279 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_4 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_330 ();
 sg13g2_fill_2 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_338 ();
 sg13g2_decap_4 FILLER_20_344 ();
 sg13g2_fill_2 FILLER_20_353 ();
 sg13g2_fill_1 FILLER_20_355 ();
 sg13g2_decap_4 FILLER_20_361 ();
 sg13g2_fill_1 FILLER_20_365 ();
 sg13g2_fill_2 FILLER_20_376 ();
 sg13g2_fill_1 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_386 ();
 sg13g2_fill_1 FILLER_20_392 ();
 sg13g2_fill_1 FILLER_20_398 ();
 sg13g2_fill_2 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_416 ();
 sg13g2_fill_2 FILLER_20_422 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_fill_1 FILLER_20_443 ();
 sg13g2_decap_4 FILLER_20_449 ();
 sg13g2_fill_2 FILLER_20_453 ();
 sg13g2_fill_2 FILLER_20_460 ();
 sg13g2_fill_2 FILLER_20_473 ();
 sg13g2_decap_4 FILLER_20_484 ();
 sg13g2_decap_4 FILLER_20_493 ();
 sg13g2_fill_1 FILLER_20_497 ();
 sg13g2_decap_4 FILLER_20_503 ();
 sg13g2_fill_2 FILLER_20_512 ();
 sg13g2_decap_8 FILLER_20_533 ();
 sg13g2_fill_2 FILLER_20_540 ();
 sg13g2_decap_8 FILLER_20_545 ();
 sg13g2_decap_8 FILLER_20_552 ();
 sg13g2_decap_8 FILLER_20_559 ();
 sg13g2_decap_8 FILLER_20_566 ();
 sg13g2_decap_8 FILLER_20_573 ();
 sg13g2_decap_4 FILLER_20_580 ();
 sg13g2_fill_2 FILLER_20_584 ();
 sg13g2_decap_8 FILLER_20_591 ();
 sg13g2_decap_8 FILLER_20_598 ();
 sg13g2_decap_8 FILLER_20_605 ();
 sg13g2_decap_8 FILLER_20_612 ();
 sg13g2_decap_8 FILLER_20_619 ();
 sg13g2_decap_8 FILLER_20_626 ();
 sg13g2_decap_8 FILLER_20_633 ();
 sg13g2_decap_8 FILLER_20_640 ();
 sg13g2_fill_1 FILLER_20_647 ();
 sg13g2_decap_8 FILLER_20_654 ();
 sg13g2_decap_8 FILLER_20_661 ();
 sg13g2_decap_8 FILLER_20_668 ();
 sg13g2_decap_8 FILLER_20_675 ();
 sg13g2_decap_4 FILLER_20_682 ();
 sg13g2_fill_1 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_691 ();
 sg13g2_decap_8 FILLER_20_698 ();
 sg13g2_decap_8 FILLER_20_705 ();
 sg13g2_decap_8 FILLER_20_712 ();
 sg13g2_fill_2 FILLER_20_719 ();
 sg13g2_fill_1 FILLER_20_747 ();
 sg13g2_fill_2 FILLER_20_779 ();
 sg13g2_fill_1 FILLER_20_781 ();
 sg13g2_fill_1 FILLER_20_790 ();
 sg13g2_decap_4 FILLER_20_799 ();
 sg13g2_fill_1 FILLER_20_803 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_4 FILLER_20_819 ();
 sg13g2_fill_1 FILLER_20_823 ();
 sg13g2_decap_8 FILLER_20_839 ();
 sg13g2_decap_8 FILLER_20_846 ();
 sg13g2_decap_8 FILLER_20_853 ();
 sg13g2_decap_4 FILLER_20_860 ();
 sg13g2_fill_2 FILLER_20_864 ();
 sg13g2_fill_2 FILLER_20_896 ();
 sg13g2_decap_8 FILLER_20_902 ();
 sg13g2_decap_8 FILLER_20_909 ();
 sg13g2_decap_8 FILLER_20_916 ();
 sg13g2_decap_4 FILLER_20_923 ();
 sg13g2_fill_2 FILLER_20_931 ();
 sg13g2_decap_8 FILLER_20_938 ();
 sg13g2_decap_8 FILLER_20_945 ();
 sg13g2_decap_8 FILLER_20_952 ();
 sg13g2_decap_8 FILLER_20_959 ();
 sg13g2_decap_8 FILLER_20_966 ();
 sg13g2_decap_8 FILLER_20_973 ();
 sg13g2_decap_8 FILLER_20_980 ();
 sg13g2_decap_8 FILLER_20_987 ();
 sg13g2_decap_8 FILLER_20_994 ();
 sg13g2_decap_4 FILLER_20_1001 ();
 sg13g2_fill_2 FILLER_20_1005 ();
 sg13g2_decap_8 FILLER_20_1022 ();
 sg13g2_fill_2 FILLER_20_1033 ();
 sg13g2_fill_1 FILLER_20_1035 ();
 sg13g2_fill_2 FILLER_20_1044 ();
 sg13g2_fill_1 FILLER_20_1046 ();
 sg13g2_decap_8 FILLER_20_1050 ();
 sg13g2_decap_4 FILLER_20_1057 ();
 sg13g2_fill_1 FILLER_20_1061 ();
 sg13g2_fill_2 FILLER_20_1080 ();
 sg13g2_fill_1 FILLER_20_1082 ();
 sg13g2_decap_8 FILLER_20_1087 ();
 sg13g2_decap_8 FILLER_20_1094 ();
 sg13g2_decap_4 FILLER_20_1124 ();
 sg13g2_decap_8 FILLER_20_1134 ();
 sg13g2_fill_2 FILLER_20_1141 ();
 sg13g2_fill_1 FILLER_20_1143 ();
 sg13g2_decap_8 FILLER_20_1152 ();
 sg13g2_decap_8 FILLER_20_1159 ();
 sg13g2_decap_8 FILLER_20_1166 ();
 sg13g2_decap_8 FILLER_20_1173 ();
 sg13g2_decap_8 FILLER_20_1180 ();
 sg13g2_fill_2 FILLER_20_1187 ();
 sg13g2_fill_1 FILLER_20_1189 ();
 sg13g2_decap_8 FILLER_20_1194 ();
 sg13g2_decap_8 FILLER_20_1201 ();
 sg13g2_decap_8 FILLER_20_1208 ();
 sg13g2_fill_2 FILLER_20_1215 ();
 sg13g2_decap_8 FILLER_20_1225 ();
 sg13g2_decap_8 FILLER_20_1232 ();
 sg13g2_decap_8 FILLER_20_1247 ();
 sg13g2_decap_8 FILLER_20_1254 ();
 sg13g2_decap_8 FILLER_20_1261 ();
 sg13g2_decap_8 FILLER_20_1268 ();
 sg13g2_decap_8 FILLER_20_1275 ();
 sg13g2_decap_8 FILLER_20_1282 ();
 sg13g2_decap_4 FILLER_20_1289 ();
 sg13g2_fill_1 FILLER_20_1293 ();
 sg13g2_fill_2 FILLER_20_1314 ();
 sg13g2_decap_8 FILLER_20_1320 ();
 sg13g2_decap_8 FILLER_20_1327 ();
 sg13g2_decap_8 FILLER_20_1334 ();
 sg13g2_decap_8 FILLER_20_1341 ();
 sg13g2_decap_8 FILLER_20_1348 ();
 sg13g2_decap_8 FILLER_20_1355 ();
 sg13g2_decap_8 FILLER_20_1362 ();
 sg13g2_decap_8 FILLER_20_1369 ();
 sg13g2_decap_8 FILLER_20_1376 ();
 sg13g2_decap_4 FILLER_20_1383 ();
 sg13g2_decap_8 FILLER_20_1391 ();
 sg13g2_decap_8 FILLER_20_1398 ();
 sg13g2_decap_8 FILLER_20_1405 ();
 sg13g2_decap_8 FILLER_20_1412 ();
 sg13g2_decap_8 FILLER_20_1419 ();
 sg13g2_decap_8 FILLER_20_1426 ();
 sg13g2_decap_8 FILLER_20_1433 ();
 sg13g2_decap_8 FILLER_20_1470 ();
 sg13g2_decap_8 FILLER_20_1477 ();
 sg13g2_decap_8 FILLER_20_1484 ();
 sg13g2_decap_8 FILLER_20_1491 ();
 sg13g2_decap_8 FILLER_20_1498 ();
 sg13g2_fill_1 FILLER_20_1505 ();
 sg13g2_decap_8 FILLER_20_1514 ();
 sg13g2_decap_8 FILLER_20_1521 ();
 sg13g2_decap_8 FILLER_20_1528 ();
 sg13g2_decap_8 FILLER_20_1535 ();
 sg13g2_fill_2 FILLER_20_1542 ();
 sg13g2_decap_8 FILLER_20_1570 ();
 sg13g2_decap_8 FILLER_20_1584 ();
 sg13g2_fill_2 FILLER_20_1591 ();
 sg13g2_fill_1 FILLER_20_1598 ();
 sg13g2_fill_1 FILLER_20_1603 ();
 sg13g2_fill_1 FILLER_20_1614 ();
 sg13g2_decap_8 FILLER_20_1627 ();
 sg13g2_decap_8 FILLER_20_1634 ();
 sg13g2_decap_8 FILLER_20_1641 ();
 sg13g2_decap_8 FILLER_20_1648 ();
 sg13g2_decap_8 FILLER_20_1655 ();
 sg13g2_decap_8 FILLER_20_1662 ();
 sg13g2_decap_8 FILLER_20_1669 ();
 sg13g2_fill_1 FILLER_20_1676 ();
 sg13g2_decap_8 FILLER_20_1681 ();
 sg13g2_fill_2 FILLER_20_1688 ();
 sg13g2_fill_1 FILLER_20_1690 ();
 sg13g2_decap_4 FILLER_20_1701 ();
 sg13g2_fill_2 FILLER_20_1705 ();
 sg13g2_decap_8 FILLER_20_1715 ();
 sg13g2_decap_8 FILLER_20_1722 ();
 sg13g2_fill_2 FILLER_20_1729 ();
 sg13g2_decap_8 FILLER_20_1740 ();
 sg13g2_decap_8 FILLER_20_1747 ();
 sg13g2_decap_8 FILLER_20_1754 ();
 sg13g2_decap_8 FILLER_20_1761 ();
 sg13g2_decap_4 FILLER_20_1768 ();
 sg13g2_fill_2 FILLER_20_1772 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_decap_4 FILLER_21_46 ();
 sg13g2_fill_2 FILLER_21_50 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_4 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_78 ();
 sg13g2_fill_2 FILLER_21_85 ();
 sg13g2_fill_1 FILLER_21_92 ();
 sg13g2_fill_1 FILLER_21_112 ();
 sg13g2_decap_4 FILLER_21_119 ();
 sg13g2_fill_1 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_129 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_4 FILLER_21_147 ();
 sg13g2_fill_1 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_4 FILLER_21_168 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_decap_4 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_fill_2 FILLER_21_209 ();
 sg13g2_decap_4 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_221 ();
 sg13g2_decap_4 FILLER_21_246 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_fill_2 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_fill_2 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_322 ();
 sg13g2_fill_2 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_347 ();
 sg13g2_fill_2 FILLER_21_354 ();
 sg13g2_fill_1 FILLER_21_356 ();
 sg13g2_decap_4 FILLER_21_363 ();
 sg13g2_fill_1 FILLER_21_367 ();
 sg13g2_fill_2 FILLER_21_373 ();
 sg13g2_fill_2 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_382 ();
 sg13g2_decap_4 FILLER_21_393 ();
 sg13g2_fill_2 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_fill_2 FILLER_21_420 ();
 sg13g2_fill_1 FILLER_21_422 ();
 sg13g2_decap_4 FILLER_21_428 ();
 sg13g2_fill_1 FILLER_21_432 ();
 sg13g2_fill_2 FILLER_21_442 ();
 sg13g2_fill_2 FILLER_21_454 ();
 sg13g2_decap_8 FILLER_21_470 ();
 sg13g2_decap_4 FILLER_21_477 ();
 sg13g2_fill_2 FILLER_21_481 ();
 sg13g2_decap_8 FILLER_21_492 ();
 sg13g2_decap_8 FILLER_21_499 ();
 sg13g2_decap_8 FILLER_21_506 ();
 sg13g2_decap_8 FILLER_21_513 ();
 sg13g2_decap_8 FILLER_21_520 ();
 sg13g2_decap_4 FILLER_21_527 ();
 sg13g2_fill_1 FILLER_21_531 ();
 sg13g2_decap_8 FILLER_21_562 ();
 sg13g2_decap_8 FILLER_21_569 ();
 sg13g2_decap_8 FILLER_21_576 ();
 sg13g2_decap_8 FILLER_21_583 ();
 sg13g2_fill_2 FILLER_21_590 ();
 sg13g2_decap_4 FILLER_21_597 ();
 sg13g2_fill_1 FILLER_21_601 ();
 sg13g2_fill_2 FILLER_21_612 ();
 sg13g2_fill_2 FILLER_21_640 ();
 sg13g2_decap_4 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_715 ();
 sg13g2_fill_1 FILLER_21_722 ();
 sg13g2_decap_8 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_746 ();
 sg13g2_decap_8 FILLER_21_753 ();
 sg13g2_decap_8 FILLER_21_760 ();
 sg13g2_decap_8 FILLER_21_767 ();
 sg13g2_decap_8 FILLER_21_774 ();
 sg13g2_decap_8 FILLER_21_781 ();
 sg13g2_fill_2 FILLER_21_788 ();
 sg13g2_fill_1 FILLER_21_790 ();
 sg13g2_decap_8 FILLER_21_795 ();
 sg13g2_decap_8 FILLER_21_802 ();
 sg13g2_decap_4 FILLER_21_809 ();
 sg13g2_fill_2 FILLER_21_813 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_21_868 ();
 sg13g2_decap_8 FILLER_21_875 ();
 sg13g2_decap_8 FILLER_21_882 ();
 sg13g2_decap_8 FILLER_21_889 ();
 sg13g2_decap_8 FILLER_21_896 ();
 sg13g2_decap_8 FILLER_21_903 ();
 sg13g2_fill_1 FILLER_21_910 ();
 sg13g2_decap_4 FILLER_21_915 ();
 sg13g2_fill_1 FILLER_21_919 ();
 sg13g2_fill_2 FILLER_21_946 ();
 sg13g2_fill_1 FILLER_21_948 ();
 sg13g2_decap_4 FILLER_21_953 ();
 sg13g2_decap_8 FILLER_21_964 ();
 sg13g2_decap_8 FILLER_21_971 ();
 sg13g2_fill_1 FILLER_21_978 ();
 sg13g2_decap_8 FILLER_21_983 ();
 sg13g2_decap_4 FILLER_21_990 ();
 sg13g2_decap_8 FILLER_21_997 ();
 sg13g2_fill_2 FILLER_21_1004 ();
 sg13g2_fill_1 FILLER_21_1006 ();
 sg13g2_decap_8 FILLER_21_1012 ();
 sg13g2_decap_8 FILLER_21_1019 ();
 sg13g2_decap_8 FILLER_21_1026 ();
 sg13g2_decap_8 FILLER_21_1033 ();
 sg13g2_decap_8 FILLER_21_1040 ();
 sg13g2_decap_8 FILLER_21_1047 ();
 sg13g2_decap_8 FILLER_21_1054 ();
 sg13g2_fill_2 FILLER_21_1061 ();
 sg13g2_decap_4 FILLER_21_1072 ();
 sg13g2_decap_8 FILLER_21_1081 ();
 sg13g2_decap_8 FILLER_21_1088 ();
 sg13g2_decap_8 FILLER_21_1095 ();
 sg13g2_decap_8 FILLER_21_1102 ();
 sg13g2_fill_2 FILLER_21_1109 ();
 sg13g2_decap_4 FILLER_21_1123 ();
 sg13g2_fill_2 FILLER_21_1127 ();
 sg13g2_decap_8 FILLER_21_1137 ();
 sg13g2_fill_2 FILLER_21_1144 ();
 sg13g2_fill_1 FILLER_21_1146 ();
 sg13g2_decap_8 FILLER_21_1166 ();
 sg13g2_decap_8 FILLER_21_1173 ();
 sg13g2_fill_2 FILLER_21_1180 ();
 sg13g2_fill_1 FILLER_21_1182 ();
 sg13g2_decap_8 FILLER_21_1188 ();
 sg13g2_fill_1 FILLER_21_1205 ();
 sg13g2_decap_4 FILLER_21_1210 ();
 sg13g2_fill_1 FILLER_21_1214 ();
 sg13g2_decap_8 FILLER_21_1225 ();
 sg13g2_decap_8 FILLER_21_1232 ();
 sg13g2_decap_8 FILLER_21_1244 ();
 sg13g2_decap_8 FILLER_21_1251 ();
 sg13g2_decap_8 FILLER_21_1258 ();
 sg13g2_decap_8 FILLER_21_1265 ();
 sg13g2_decap_8 FILLER_21_1272 ();
 sg13g2_decap_8 FILLER_21_1279 ();
 sg13g2_decap_8 FILLER_21_1286 ();
 sg13g2_decap_4 FILLER_21_1293 ();
 sg13g2_decap_8 FILLER_21_1302 ();
 sg13g2_decap_8 FILLER_21_1309 ();
 sg13g2_decap_8 FILLER_21_1316 ();
 sg13g2_decap_8 FILLER_21_1323 ();
 sg13g2_decap_8 FILLER_21_1330 ();
 sg13g2_decap_4 FILLER_21_1343 ();
 sg13g2_fill_2 FILLER_21_1347 ();
 sg13g2_decap_8 FILLER_21_1362 ();
 sg13g2_fill_2 FILLER_21_1369 ();
 sg13g2_decap_8 FILLER_21_1408 ();
 sg13g2_fill_2 FILLER_21_1415 ();
 sg13g2_decap_8 FILLER_21_1421 ();
 sg13g2_decap_8 FILLER_21_1428 ();
 sg13g2_decap_8 FILLER_21_1435 ();
 sg13g2_decap_8 FILLER_21_1442 ();
 sg13g2_decap_8 FILLER_21_1453 ();
 sg13g2_decap_8 FILLER_21_1460 ();
 sg13g2_decap_8 FILLER_21_1467 ();
 sg13g2_decap_4 FILLER_21_1474 ();
 sg13g2_fill_1 FILLER_21_1478 ();
 sg13g2_decap_8 FILLER_21_1483 ();
 sg13g2_decap_8 FILLER_21_1490 ();
 sg13g2_decap_8 FILLER_21_1497 ();
 sg13g2_decap_8 FILLER_21_1504 ();
 sg13g2_decap_8 FILLER_21_1511 ();
 sg13g2_decap_8 FILLER_21_1518 ();
 sg13g2_decap_4 FILLER_21_1525 ();
 sg13g2_decap_8 FILLER_21_1533 ();
 sg13g2_decap_8 FILLER_21_1540 ();
 sg13g2_decap_8 FILLER_21_1547 ();
 sg13g2_decap_8 FILLER_21_1554 ();
 sg13g2_fill_1 FILLER_21_1561 ();
 sg13g2_decap_4 FILLER_21_1570 ();
 sg13g2_decap_8 FILLER_21_1583 ();
 sg13g2_decap_8 FILLER_21_1590 ();
 sg13g2_fill_2 FILLER_21_1602 ();
 sg13g2_decap_4 FILLER_21_1610 ();
 sg13g2_decap_8 FILLER_21_1619 ();
 sg13g2_decap_8 FILLER_21_1626 ();
 sg13g2_fill_2 FILLER_21_1633 ();
 sg13g2_decap_4 FILLER_21_1665 ();
 sg13g2_fill_1 FILLER_21_1669 ();
 sg13g2_decap_8 FILLER_21_1696 ();
 sg13g2_decap_4 FILLER_21_1703 ();
 sg13g2_fill_2 FILLER_21_1707 ();
 sg13g2_decap_8 FILLER_21_1714 ();
 sg13g2_fill_2 FILLER_21_1721 ();
 sg13g2_fill_1 FILLER_21_1723 ();
 sg13g2_decap_8 FILLER_21_1750 ();
 sg13g2_decap_8 FILLER_21_1757 ();
 sg13g2_decap_8 FILLER_21_1764 ();
 sg13g2_fill_2 FILLER_21_1771 ();
 sg13g2_fill_1 FILLER_21_1773 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_39 ();
 sg13g2_decap_4 FILLER_22_45 ();
 sg13g2_fill_1 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_59 ();
 sg13g2_decap_8 FILLER_22_66 ();
 sg13g2_decap_8 FILLER_22_73 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_fill_2 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_129 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_decap_4 FILLER_22_146 ();
 sg13g2_decap_4 FILLER_22_155 ();
 sg13g2_decap_8 FILLER_22_162 ();
 sg13g2_decap_8 FILLER_22_169 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_4 FILLER_22_231 ();
 sg13g2_fill_1 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_4 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_256 ();
 sg13g2_fill_2 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_281 ();
 sg13g2_fill_2 FILLER_22_287 ();
 sg13g2_fill_2 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_300 ();
 sg13g2_fill_1 FILLER_22_307 ();
 sg13g2_fill_2 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_325 ();
 sg13g2_decap_4 FILLER_22_332 ();
 sg13g2_fill_1 FILLER_22_336 ();
 sg13g2_decap_4 FILLER_22_348 ();
 sg13g2_fill_2 FILLER_22_352 ();
 sg13g2_decap_8 FILLER_22_358 ();
 sg13g2_decap_4 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_4 FILLER_22_402 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_decap_4 FILLER_22_414 ();
 sg13g2_fill_2 FILLER_22_423 ();
 sg13g2_fill_2 FILLER_22_430 ();
 sg13g2_fill_1 FILLER_22_432 ();
 sg13g2_decap_4 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_fill_2 FILLER_22_525 ();
 sg13g2_fill_1 FILLER_22_527 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_fill_2 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_561 ();
 sg13g2_decap_8 FILLER_22_568 ();
 sg13g2_decap_4 FILLER_22_575 ();
 sg13g2_fill_1 FILLER_22_579 ();
 sg13g2_decap_8 FILLER_22_583 ();
 sg13g2_decap_8 FILLER_22_590 ();
 sg13g2_decap_8 FILLER_22_597 ();
 sg13g2_decap_8 FILLER_22_604 ();
 sg13g2_decap_8 FILLER_22_611 ();
 sg13g2_fill_2 FILLER_22_618 ();
 sg13g2_fill_1 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_625 ();
 sg13g2_decap_8 FILLER_22_632 ();
 sg13g2_decap_8 FILLER_22_639 ();
 sg13g2_decap_8 FILLER_22_646 ();
 sg13g2_decap_4 FILLER_22_653 ();
 sg13g2_fill_2 FILLER_22_657 ();
 sg13g2_decap_8 FILLER_22_663 ();
 sg13g2_decap_8 FILLER_22_670 ();
 sg13g2_decap_8 FILLER_22_677 ();
 sg13g2_decap_8 FILLER_22_684 ();
 sg13g2_decap_8 FILLER_22_691 ();
 sg13g2_decap_8 FILLER_22_698 ();
 sg13g2_decap_8 FILLER_22_705 ();
 sg13g2_decap_4 FILLER_22_712 ();
 sg13g2_fill_2 FILLER_22_716 ();
 sg13g2_decap_4 FILLER_22_721 ();
 sg13g2_fill_2 FILLER_22_725 ();
 sg13g2_decap_4 FILLER_22_755 ();
 sg13g2_fill_2 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_795 ();
 sg13g2_decap_8 FILLER_22_802 ();
 sg13g2_fill_1 FILLER_22_809 ();
 sg13g2_fill_2 FILLER_22_826 ();
 sg13g2_fill_2 FILLER_22_847 ();
 sg13g2_fill_1 FILLER_22_849 ();
 sg13g2_decap_8 FILLER_22_855 ();
 sg13g2_decap_4 FILLER_22_862 ();
 sg13g2_fill_1 FILLER_22_866 ();
 sg13g2_decap_8 FILLER_22_875 ();
 sg13g2_decap_8 FILLER_22_882 ();
 sg13g2_decap_8 FILLER_22_889 ();
 sg13g2_decap_8 FILLER_22_896 ();
 sg13g2_fill_2 FILLER_22_903 ();
 sg13g2_fill_1 FILLER_22_905 ();
 sg13g2_decap_8 FILLER_22_910 ();
 sg13g2_fill_2 FILLER_22_917 ();
 sg13g2_decap_8 FILLER_22_924 ();
 sg13g2_decap_8 FILLER_22_931 ();
 sg13g2_decap_8 FILLER_22_938 ();
 sg13g2_fill_1 FILLER_22_945 ();
 sg13g2_fill_2 FILLER_22_950 ();
 sg13g2_fill_1 FILLER_22_952 ();
 sg13g2_decap_8 FILLER_22_965 ();
 sg13g2_fill_2 FILLER_22_998 ();
 sg13g2_fill_1 FILLER_22_1000 ();
 sg13g2_decap_8 FILLER_22_1031 ();
 sg13g2_fill_1 FILLER_22_1038 ();
 sg13g2_decap_4 FILLER_22_1044 ();
 sg13g2_decap_4 FILLER_22_1058 ();
 sg13g2_fill_2 FILLER_22_1062 ();
 sg13g2_fill_2 FILLER_22_1080 ();
 sg13g2_fill_1 FILLER_22_1082 ();
 sg13g2_fill_2 FILLER_22_1109 ();
 sg13g2_decap_8 FILLER_22_1127 ();
 sg13g2_fill_2 FILLER_22_1134 ();
 sg13g2_decap_8 FILLER_22_1140 ();
 sg13g2_fill_1 FILLER_22_1147 ();
 sg13g2_fill_2 FILLER_22_1154 ();
 sg13g2_fill_1 FILLER_22_1156 ();
 sg13g2_fill_2 FILLER_22_1160 ();
 sg13g2_fill_1 FILLER_22_1162 ();
 sg13g2_decap_8 FILLER_22_1168 ();
 sg13g2_decap_8 FILLER_22_1175 ();
 sg13g2_decap_8 FILLER_22_1182 ();
 sg13g2_fill_2 FILLER_22_1208 ();
 sg13g2_decap_8 FILLER_22_1223 ();
 sg13g2_decap_4 FILLER_22_1230 ();
 sg13g2_decap_4 FILLER_22_1275 ();
 sg13g2_fill_1 FILLER_22_1279 ();
 sg13g2_fill_2 FILLER_22_1288 ();
 sg13g2_decap_4 FILLER_22_1294 ();
 sg13g2_fill_1 FILLER_22_1304 ();
 sg13g2_fill_1 FILLER_22_1310 ();
 sg13g2_decap_8 FILLER_22_1328 ();
 sg13g2_fill_1 FILLER_22_1335 ();
 sg13g2_decap_4 FILLER_22_1341 ();
 sg13g2_decap_8 FILLER_22_1355 ();
 sg13g2_decap_8 FILLER_22_1362 ();
 sg13g2_fill_2 FILLER_22_1369 ();
 sg13g2_decap_8 FILLER_22_1376 ();
 sg13g2_fill_2 FILLER_22_1383 ();
 sg13g2_decap_8 FILLER_22_1389 ();
 sg13g2_decap_8 FILLER_22_1396 ();
 sg13g2_decap_8 FILLER_22_1403 ();
 sg13g2_decap_8 FILLER_22_1436 ();
 sg13g2_fill_2 FILLER_22_1443 ();
 sg13g2_decap_8 FILLER_22_1462 ();
 sg13g2_fill_2 FILLER_22_1469 ();
 sg13g2_fill_1 FILLER_22_1471 ();
 sg13g2_decap_8 FILLER_22_1498 ();
 sg13g2_decap_4 FILLER_22_1505 ();
 sg13g2_fill_2 FILLER_22_1509 ();
 sg13g2_decap_8 FILLER_22_1515 ();
 sg13g2_decap_8 FILLER_22_1522 ();
 sg13g2_decap_8 FILLER_22_1529 ();
 sg13g2_decap_8 FILLER_22_1536 ();
 sg13g2_fill_2 FILLER_22_1543 ();
 sg13g2_decap_8 FILLER_22_1551 ();
 sg13g2_decap_8 FILLER_22_1558 ();
 sg13g2_decap_8 FILLER_22_1565 ();
 sg13g2_decap_8 FILLER_22_1572 ();
 sg13g2_decap_8 FILLER_22_1579 ();
 sg13g2_decap_8 FILLER_22_1586 ();
 sg13g2_decap_8 FILLER_22_1593 ();
 sg13g2_decap_8 FILLER_22_1600 ();
 sg13g2_fill_2 FILLER_22_1607 ();
 sg13g2_decap_8 FILLER_22_1614 ();
 sg13g2_decap_8 FILLER_22_1621 ();
 sg13g2_decap_8 FILLER_22_1628 ();
 sg13g2_decap_8 FILLER_22_1635 ();
 sg13g2_decap_4 FILLER_22_1642 ();
 sg13g2_fill_2 FILLER_22_1646 ();
 sg13g2_fill_2 FILLER_22_1652 ();
 sg13g2_fill_1 FILLER_22_1654 ();
 sg13g2_decap_4 FILLER_22_1669 ();
 sg13g2_fill_1 FILLER_22_1673 ();
 sg13g2_decap_8 FILLER_22_1681 ();
 sg13g2_fill_1 FILLER_22_1693 ();
 sg13g2_decap_8 FILLER_22_1698 ();
 sg13g2_fill_2 FILLER_22_1705 ();
 sg13g2_fill_1 FILLER_22_1707 ();
 sg13g2_decap_8 FILLER_22_1712 ();
 sg13g2_decap_8 FILLER_22_1719 ();
 sg13g2_decap_8 FILLER_22_1726 ();
 sg13g2_decap_8 FILLER_22_1733 ();
 sg13g2_decap_8 FILLER_22_1740 ();
 sg13g2_decap_8 FILLER_22_1747 ();
 sg13g2_decap_8 FILLER_22_1754 ();
 sg13g2_decap_8 FILLER_22_1761 ();
 sg13g2_decap_4 FILLER_22_1768 ();
 sg13g2_fill_2 FILLER_22_1772 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_30 ();
 sg13g2_fill_1 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_47 ();
 sg13g2_decap_4 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_61 ();
 sg13g2_fill_2 FILLER_23_68 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_2 FILLER_23_89 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_fill_1 FILLER_23_102 ();
 sg13g2_fill_2 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_111 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_fill_2 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_148 ();
 sg13g2_decap_8 FILLER_23_155 ();
 sg13g2_decap_8 FILLER_23_162 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_fill_1 FILLER_23_179 ();
 sg13g2_fill_2 FILLER_23_185 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_4 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_246 ();
 sg13g2_decap_4 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_325 ();
 sg13g2_decap_4 FILLER_23_332 ();
 sg13g2_fill_1 FILLER_23_336 ();
 sg13g2_fill_1 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_decap_4 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_363 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_fill_2 FILLER_23_384 ();
 sg13g2_fill_1 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_fill_1 FILLER_23_409 ();
 sg13g2_decap_8 FILLER_23_415 ();
 sg13g2_decap_8 FILLER_23_422 ();
 sg13g2_decap_4 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_decap_8 FILLER_23_452 ();
 sg13g2_fill_1 FILLER_23_472 ();
 sg13g2_decap_8 FILLER_23_482 ();
 sg13g2_decap_8 FILLER_23_489 ();
 sg13g2_decap_8 FILLER_23_496 ();
 sg13g2_decap_8 FILLER_23_509 ();
 sg13g2_fill_2 FILLER_23_516 ();
 sg13g2_fill_1 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_548 ();
 sg13g2_decap_4 FILLER_23_555 ();
 sg13g2_decap_8 FILLER_23_585 ();
 sg13g2_decap_8 FILLER_23_618 ();
 sg13g2_decap_8 FILLER_23_625 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_4 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_701 ();
 sg13g2_decap_8 FILLER_23_708 ();
 sg13g2_fill_2 FILLER_23_715 ();
 sg13g2_decap_4 FILLER_23_721 ();
 sg13g2_decap_4 FILLER_23_730 ();
 sg13g2_fill_1 FILLER_23_734 ();
 sg13g2_decap_8 FILLER_23_739 ();
 sg13g2_decap_8 FILLER_23_746 ();
 sg13g2_decap_4 FILLER_23_753 ();
 sg13g2_fill_1 FILLER_23_757 ();
 sg13g2_decap_8 FILLER_23_766 ();
 sg13g2_decap_8 FILLER_23_773 ();
 sg13g2_decap_8 FILLER_23_780 ();
 sg13g2_decap_8 FILLER_23_787 ();
 sg13g2_decap_8 FILLER_23_794 ();
 sg13g2_decap_8 FILLER_23_801 ();
 sg13g2_decap_8 FILLER_23_808 ();
 sg13g2_decap_8 FILLER_23_815 ();
 sg13g2_decap_8 FILLER_23_822 ();
 sg13g2_fill_1 FILLER_23_829 ();
 sg13g2_decap_8 FILLER_23_834 ();
 sg13g2_decap_8 FILLER_23_841 ();
 sg13g2_decap_8 FILLER_23_848 ();
 sg13g2_decap_4 FILLER_23_855 ();
 sg13g2_fill_1 FILLER_23_859 ();
 sg13g2_fill_2 FILLER_23_871 ();
 sg13g2_decap_8 FILLER_23_878 ();
 sg13g2_decap_8 FILLER_23_885 ();
 sg13g2_decap_8 FILLER_23_892 ();
 sg13g2_decap_8 FILLER_23_899 ();
 sg13g2_decap_8 FILLER_23_906 ();
 sg13g2_decap_4 FILLER_23_913 ();
 sg13g2_fill_1 FILLER_23_917 ();
 sg13g2_decap_4 FILLER_23_940 ();
 sg13g2_fill_2 FILLER_23_954 ();
 sg13g2_fill_1 FILLER_23_956 ();
 sg13g2_decap_8 FILLER_23_967 ();
 sg13g2_fill_2 FILLER_23_974 ();
 sg13g2_decap_8 FILLER_23_981 ();
 sg13g2_decap_8 FILLER_23_988 ();
 sg13g2_decap_8 FILLER_23_995 ();
 sg13g2_fill_2 FILLER_23_1002 ();
 sg13g2_fill_1 FILLER_23_1004 ();
 sg13g2_decap_8 FILLER_23_1010 ();
 sg13g2_decap_8 FILLER_23_1017 ();
 sg13g2_fill_2 FILLER_23_1024 ();
 sg13g2_decap_8 FILLER_23_1044 ();
 sg13g2_decap_8 FILLER_23_1051 ();
 sg13g2_decap_8 FILLER_23_1058 ();
 sg13g2_fill_2 FILLER_23_1065 ();
 sg13g2_decap_8 FILLER_23_1077 ();
 sg13g2_decap_8 FILLER_23_1084 ();
 sg13g2_decap_4 FILLER_23_1095 ();
 sg13g2_decap_8 FILLER_23_1103 ();
 sg13g2_fill_1 FILLER_23_1110 ();
 sg13g2_fill_2 FILLER_23_1122 ();
 sg13g2_decap_8 FILLER_23_1150 ();
 sg13g2_decap_8 FILLER_23_1217 ();
 sg13g2_decap_8 FILLER_23_1224 ();
 sg13g2_decap_8 FILLER_23_1231 ();
 sg13g2_decap_8 FILLER_23_1238 ();
 sg13g2_decap_4 FILLER_23_1245 ();
 sg13g2_fill_2 FILLER_23_1249 ();
 sg13g2_decap_8 FILLER_23_1255 ();
 sg13g2_decap_8 FILLER_23_1262 ();
 sg13g2_decap_8 FILLER_23_1269 ();
 sg13g2_fill_2 FILLER_23_1292 ();
 sg13g2_fill_1 FILLER_23_1294 ();
 sg13g2_decap_4 FILLER_23_1300 ();
 sg13g2_fill_1 FILLER_23_1304 ();
 sg13g2_fill_1 FILLER_23_1314 ();
 sg13g2_decap_8 FILLER_23_1319 ();
 sg13g2_decap_4 FILLER_23_1326 ();
 sg13g2_fill_2 FILLER_23_1330 ();
 sg13g2_decap_8 FILLER_23_1336 ();
 sg13g2_decap_4 FILLER_23_1343 ();
 sg13g2_fill_2 FILLER_23_1347 ();
 sg13g2_decap_8 FILLER_23_1379 ();
 sg13g2_decap_8 FILLER_23_1386 ();
 sg13g2_decap_8 FILLER_23_1393 ();
 sg13g2_fill_1 FILLER_23_1400 ();
 sg13g2_decap_8 FILLER_23_1404 ();
 sg13g2_decap_8 FILLER_23_1411 ();
 sg13g2_decap_8 FILLER_23_1423 ();
 sg13g2_decap_8 FILLER_23_1430 ();
 sg13g2_decap_4 FILLER_23_1437 ();
 sg13g2_fill_2 FILLER_23_1441 ();
 sg13g2_decap_4 FILLER_23_1469 ();
 sg13g2_decap_8 FILLER_23_1477 ();
 sg13g2_decap_8 FILLER_23_1484 ();
 sg13g2_fill_1 FILLER_23_1491 ();
 sg13g2_decap_4 FILLER_23_1497 ();
 sg13g2_fill_2 FILLER_23_1501 ();
 sg13g2_decap_8 FILLER_23_1533 ();
 sg13g2_fill_2 FILLER_23_1540 ();
 sg13g2_fill_1 FILLER_23_1542 ();
 sg13g2_decap_8 FILLER_23_1547 ();
 sg13g2_decap_8 FILLER_23_1554 ();
 sg13g2_fill_2 FILLER_23_1561 ();
 sg13g2_fill_2 FILLER_23_1589 ();
 sg13g2_fill_1 FILLER_23_1608 ();
 sg13g2_decap_8 FILLER_23_1613 ();
 sg13g2_fill_2 FILLER_23_1620 ();
 sg13g2_fill_1 FILLER_23_1622 ();
 sg13g2_fill_1 FILLER_23_1628 ();
 sg13g2_fill_1 FILLER_23_1635 ();
 sg13g2_fill_1 FILLER_23_1641 ();
 sg13g2_fill_1 FILLER_23_1646 ();
 sg13g2_fill_2 FILLER_23_1655 ();
 sg13g2_fill_2 FILLER_23_1679 ();
 sg13g2_fill_2 FILLER_23_1696 ();
 sg13g2_decap_8 FILLER_23_1703 ();
 sg13g2_decap_8 FILLER_23_1710 ();
 sg13g2_decap_8 FILLER_23_1717 ();
 sg13g2_decap_8 FILLER_23_1724 ();
 sg13g2_decap_8 FILLER_23_1731 ();
 sg13g2_decap_8 FILLER_23_1738 ();
 sg13g2_decap_8 FILLER_23_1745 ();
 sg13g2_decap_8 FILLER_23_1752 ();
 sg13g2_decap_8 FILLER_23_1759 ();
 sg13g2_decap_8 FILLER_23_1766 ();
 sg13g2_fill_1 FILLER_23_1773 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_65 ();
 sg13g2_decap_8 FILLER_24_72 ();
 sg13g2_fill_2 FILLER_24_79 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_93 ();
 sg13g2_fill_2 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_fill_1 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_decap_4 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_204 ();
 sg13g2_decap_4 FILLER_24_210 ();
 sg13g2_fill_1 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_fill_2 FILLER_24_263 ();
 sg13g2_decap_4 FILLER_24_270 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_fill_2 FILLER_24_324 ();
 sg13g2_decap_4 FILLER_24_331 ();
 sg13g2_fill_2 FILLER_24_335 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_fill_2 FILLER_24_389 ();
 sg13g2_decap_4 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_2 FILLER_24_414 ();
 sg13g2_decap_4 FILLER_24_421 ();
 sg13g2_decap_8 FILLER_24_430 ();
 sg13g2_fill_2 FILLER_24_437 ();
 sg13g2_fill_1 FILLER_24_439 ();
 sg13g2_decap_8 FILLER_24_445 ();
 sg13g2_decap_4 FILLER_24_452 ();
 sg13g2_fill_2 FILLER_24_456 ();
 sg13g2_decap_8 FILLER_24_471 ();
 sg13g2_decap_8 FILLER_24_478 ();
 sg13g2_decap_8 FILLER_24_485 ();
 sg13g2_decap_8 FILLER_24_492 ();
 sg13g2_decap_8 FILLER_24_499 ();
 sg13g2_fill_2 FILLER_24_506 ();
 sg13g2_fill_1 FILLER_24_508 ();
 sg13g2_decap_8 FILLER_24_524 ();
 sg13g2_decap_8 FILLER_24_535 ();
 sg13g2_decap_8 FILLER_24_542 ();
 sg13g2_decap_8 FILLER_24_549 ();
 sg13g2_decap_8 FILLER_24_556 ();
 sg13g2_fill_2 FILLER_24_563 ();
 sg13g2_decap_8 FILLER_24_569 ();
 sg13g2_decap_4 FILLER_24_576 ();
 sg13g2_fill_1 FILLER_24_580 ();
 sg13g2_decap_8 FILLER_24_586 ();
 sg13g2_decap_4 FILLER_24_593 ();
 sg13g2_fill_1 FILLER_24_597 ();
 sg13g2_decap_8 FILLER_24_628 ();
 sg13g2_fill_1 FILLER_24_635 ();
 sg13g2_decap_8 FILLER_24_640 ();
 sg13g2_decap_8 FILLER_24_647 ();
 sg13g2_decap_8 FILLER_24_654 ();
 sg13g2_decap_4 FILLER_24_661 ();
 sg13g2_fill_2 FILLER_24_665 ();
 sg13g2_fill_1 FILLER_24_674 ();
 sg13g2_decap_4 FILLER_24_705 ();
 sg13g2_fill_1 FILLER_24_709 ();
 sg13g2_decap_8 FILLER_24_736 ();
 sg13g2_decap_8 FILLER_24_743 ();
 sg13g2_decap_4 FILLER_24_750 ();
 sg13g2_fill_2 FILLER_24_759 ();
 sg13g2_fill_1 FILLER_24_761 ();
 sg13g2_decap_8 FILLER_24_766 ();
 sg13g2_decap_8 FILLER_24_773 ();
 sg13g2_fill_1 FILLER_24_780 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_fill_2 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_4 FILLER_24_847 ();
 sg13g2_fill_1 FILLER_24_851 ();
 sg13g2_fill_2 FILLER_24_856 ();
 sg13g2_fill_1 FILLER_24_858 ();
 sg13g2_fill_2 FILLER_24_864 ();
 sg13g2_decap_8 FILLER_24_878 ();
 sg13g2_decap_8 FILLER_24_885 ();
 sg13g2_fill_1 FILLER_24_892 ();
 sg13g2_decap_8 FILLER_24_898 ();
 sg13g2_decap_4 FILLER_24_905 ();
 sg13g2_fill_1 FILLER_24_909 ();
 sg13g2_decap_8 FILLER_24_920 ();
 sg13g2_fill_2 FILLER_24_944 ();
 sg13g2_fill_1 FILLER_24_946 ();
 sg13g2_decap_8 FILLER_24_951 ();
 sg13g2_decap_8 FILLER_24_958 ();
 sg13g2_decap_8 FILLER_24_965 ();
 sg13g2_fill_2 FILLER_24_972 ();
 sg13g2_decap_4 FILLER_24_979 ();
 sg13g2_fill_1 FILLER_24_983 ();
 sg13g2_decap_4 FILLER_24_995 ();
 sg13g2_fill_1 FILLER_24_999 ();
 sg13g2_decap_8 FILLER_24_1010 ();
 sg13g2_decap_8 FILLER_24_1017 ();
 sg13g2_decap_8 FILLER_24_1024 ();
 sg13g2_fill_1 FILLER_24_1047 ();
 sg13g2_fill_2 FILLER_24_1056 ();
 sg13g2_fill_2 FILLER_24_1062 ();
 sg13g2_fill_1 FILLER_24_1070 ();
 sg13g2_fill_1 FILLER_24_1084 ();
 sg13g2_decap_8 FILLER_24_1116 ();
 sg13g2_decap_8 FILLER_24_1123 ();
 sg13g2_fill_2 FILLER_24_1130 ();
 sg13g2_decap_8 FILLER_24_1136 ();
 sg13g2_decap_8 FILLER_24_1143 ();
 sg13g2_decap_8 FILLER_24_1150 ();
 sg13g2_decap_8 FILLER_24_1157 ();
 sg13g2_decap_8 FILLER_24_1168 ();
 sg13g2_decap_8 FILLER_24_1175 ();
 sg13g2_decap_8 FILLER_24_1182 ();
 sg13g2_decap_8 FILLER_24_1189 ();
 sg13g2_fill_1 FILLER_24_1196 ();
 sg13g2_decap_8 FILLER_24_1228 ();
 sg13g2_fill_2 FILLER_24_1235 ();
 sg13g2_fill_1 FILLER_24_1242 ();
 sg13g2_decap_8 FILLER_24_1261 ();
 sg13g2_decap_8 FILLER_24_1268 ();
 sg13g2_fill_1 FILLER_24_1275 ();
 sg13g2_fill_2 FILLER_24_1287 ();
 sg13g2_fill_1 FILLER_24_1289 ();
 sg13g2_decap_4 FILLER_24_1305 ();
 sg13g2_decap_8 FILLER_24_1335 ();
 sg13g2_decap_8 FILLER_24_1342 ();
 sg13g2_decap_8 FILLER_24_1349 ();
 sg13g2_fill_2 FILLER_24_1356 ();
 sg13g2_fill_1 FILLER_24_1358 ();
 sg13g2_decap_8 FILLER_24_1363 ();
 sg13g2_decap_8 FILLER_24_1370 ();
 sg13g2_fill_1 FILLER_24_1382 ();
 sg13g2_fill_1 FILLER_24_1412 ();
 sg13g2_decap_8 FILLER_24_1418 ();
 sg13g2_decap_4 FILLER_24_1425 ();
 sg13g2_fill_2 FILLER_24_1429 ();
 sg13g2_decap_4 FILLER_24_1446 ();
 sg13g2_fill_1 FILLER_24_1450 ();
 sg13g2_decap_8 FILLER_24_1455 ();
 sg13g2_decap_8 FILLER_24_1462 ();
 sg13g2_fill_1 FILLER_24_1469 ();
 sg13g2_decap_8 FILLER_24_1494 ();
 sg13g2_decap_4 FILLER_24_1501 ();
 sg13g2_decap_8 FILLER_24_1513 ();
 sg13g2_decap_8 FILLER_24_1520 ();
 sg13g2_decap_4 FILLER_24_1527 ();
 sg13g2_decap_4 FILLER_24_1536 ();
 sg13g2_fill_1 FILLER_24_1540 ();
 sg13g2_decap_4 FILLER_24_1545 ();
 sg13g2_fill_1 FILLER_24_1549 ();
 sg13g2_decap_4 FILLER_24_1556 ();
 sg13g2_fill_1 FILLER_24_1560 ();
 sg13g2_fill_2 FILLER_24_1566 ();
 sg13g2_fill_1 FILLER_24_1568 ();
 sg13g2_decap_8 FILLER_24_1573 ();
 sg13g2_decap_4 FILLER_24_1580 ();
 sg13g2_decap_8 FILLER_24_1588 ();
 sg13g2_decap_8 FILLER_24_1595 ();
 sg13g2_decap_8 FILLER_24_1602 ();
 sg13g2_decap_4 FILLER_24_1609 ();
 sg13g2_fill_1 FILLER_24_1613 ();
 sg13g2_decap_4 FILLER_24_1625 ();
 sg13g2_fill_2 FILLER_24_1629 ();
 sg13g2_decap_8 FILLER_24_1634 ();
 sg13g2_decap_8 FILLER_24_1641 ();
 sg13g2_decap_8 FILLER_24_1648 ();
 sg13g2_fill_2 FILLER_24_1655 ();
 sg13g2_decap_8 FILLER_24_1661 ();
 sg13g2_decap_8 FILLER_24_1668 ();
 sg13g2_decap_8 FILLER_24_1675 ();
 sg13g2_decap_8 FILLER_24_1682 ();
 sg13g2_decap_8 FILLER_24_1689 ();
 sg13g2_decap_4 FILLER_24_1696 ();
 sg13g2_fill_2 FILLER_24_1700 ();
 sg13g2_decap_8 FILLER_24_1715 ();
 sg13g2_decap_8 FILLER_24_1722 ();
 sg13g2_decap_8 FILLER_24_1729 ();
 sg13g2_fill_1 FILLER_24_1736 ();
 sg13g2_decap_8 FILLER_24_1741 ();
 sg13g2_decap_8 FILLER_24_1748 ();
 sg13g2_decap_8 FILLER_24_1755 ();
 sg13g2_decap_8 FILLER_24_1762 ();
 sg13g2_decap_4 FILLER_24_1769 ();
 sg13g2_fill_1 FILLER_24_1773 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_18 ();
 sg13g2_decap_4 FILLER_25_24 ();
 sg13g2_fill_1 FILLER_25_33 ();
 sg13g2_decap_4 FILLER_25_38 ();
 sg13g2_fill_2 FILLER_25_46 ();
 sg13g2_fill_1 FILLER_25_48 ();
 sg13g2_decap_4 FILLER_25_59 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_2 FILLER_25_89 ();
 sg13g2_fill_2 FILLER_25_95 ();
 sg13g2_decap_4 FILLER_25_106 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_fill_2 FILLER_25_120 ();
 sg13g2_fill_2 FILLER_25_127 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_fill_2 FILLER_25_143 ();
 sg13g2_fill_1 FILLER_25_145 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_decap_4 FILLER_25_157 ();
 sg13g2_fill_1 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_fill_1 FILLER_25_186 ();
 sg13g2_decap_4 FILLER_25_197 ();
 sg13g2_decap_8 FILLER_25_206 ();
 sg13g2_decap_4 FILLER_25_213 ();
 sg13g2_decap_4 FILLER_25_222 ();
 sg13g2_decap_4 FILLER_25_231 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_240 ();
 sg13g2_fill_2 FILLER_25_247 ();
 sg13g2_decap_8 FILLER_25_253 ();
 sg13g2_decap_8 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_fill_2 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_292 ();
 sg13g2_decap_8 FILLER_25_299 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_fill_2 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_25_360 ();
 sg13g2_decap_8 FILLER_25_374 ();
 sg13g2_decap_4 FILLER_25_381 ();
 sg13g2_fill_1 FILLER_25_385 ();
 sg13g2_fill_1 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_fill_2 FILLER_25_413 ();
 sg13g2_fill_2 FILLER_25_420 ();
 sg13g2_fill_1 FILLER_25_422 ();
 sg13g2_decap_8 FILLER_25_426 ();
 sg13g2_decap_4 FILLER_25_433 ();
 sg13g2_fill_2 FILLER_25_437 ();
 sg13g2_decap_8 FILLER_25_444 ();
 sg13g2_fill_1 FILLER_25_459 ();
 sg13g2_decap_8 FILLER_25_465 ();
 sg13g2_fill_2 FILLER_25_472 ();
 sg13g2_fill_1 FILLER_25_474 ();
 sg13g2_decap_8 FILLER_25_480 ();
 sg13g2_decap_8 FILLER_25_487 ();
 sg13g2_fill_2 FILLER_25_494 ();
 sg13g2_fill_1 FILLER_25_496 ();
 sg13g2_decap_8 FILLER_25_548 ();
 sg13g2_decap_4 FILLER_25_555 ();
 sg13g2_fill_1 FILLER_25_590 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_4 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_645 ();
 sg13g2_decap_8 FILLER_25_652 ();
 sg13g2_decap_8 FILLER_25_659 ();
 sg13g2_decap_8 FILLER_25_666 ();
 sg13g2_decap_8 FILLER_25_673 ();
 sg13g2_fill_1 FILLER_25_680 ();
 sg13g2_decap_8 FILLER_25_698 ();
 sg13g2_decap_8 FILLER_25_705 ();
 sg13g2_decap_8 FILLER_25_712 ();
 sg13g2_fill_1 FILLER_25_719 ();
 sg13g2_decap_8 FILLER_25_725 ();
 sg13g2_decap_8 FILLER_25_732 ();
 sg13g2_fill_2 FILLER_25_739 ();
 sg13g2_fill_1 FILLER_25_741 ();
 sg13g2_decap_8 FILLER_25_745 ();
 sg13g2_fill_2 FILLER_25_752 ();
 sg13g2_fill_1 FILLER_25_754 ();
 sg13g2_decap_8 FILLER_25_781 ();
 sg13g2_decap_4 FILLER_25_788 ();
 sg13g2_fill_1 FILLER_25_792 ();
 sg13g2_decap_8 FILLER_25_797 ();
 sg13g2_decap_8 FILLER_25_804 ();
 sg13g2_decap_8 FILLER_25_811 ();
 sg13g2_decap_8 FILLER_25_818 ();
 sg13g2_fill_2 FILLER_25_825 ();
 sg13g2_fill_1 FILLER_25_831 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_4 FILLER_25_854 ();
 sg13g2_fill_1 FILLER_25_858 ();
 sg13g2_decap_4 FILLER_25_863 ();
 sg13g2_fill_2 FILLER_25_867 ();
 sg13g2_decap_8 FILLER_25_881 ();
 sg13g2_fill_1 FILLER_25_888 ();
 sg13g2_decap_8 FILLER_25_896 ();
 sg13g2_fill_2 FILLER_25_903 ();
 sg13g2_fill_1 FILLER_25_905 ();
 sg13g2_decap_4 FILLER_25_925 ();
 sg13g2_fill_2 FILLER_25_929 ();
 sg13g2_fill_2 FILLER_25_936 ();
 sg13g2_fill_1 FILLER_25_938 ();
 sg13g2_decap_8 FILLER_25_948 ();
 sg13g2_fill_2 FILLER_25_955 ();
 sg13g2_fill_2 FILLER_25_963 ();
 sg13g2_decap_8 FILLER_25_969 ();
 sg13g2_decap_8 FILLER_25_976 ();
 sg13g2_fill_2 FILLER_25_983 ();
 sg13g2_fill_2 FILLER_25_996 ();
 sg13g2_decap_8 FILLER_25_1009 ();
 sg13g2_decap_4 FILLER_25_1016 ();
 sg13g2_fill_2 FILLER_25_1020 ();
 sg13g2_fill_1 FILLER_25_1049 ();
 sg13g2_fill_2 FILLER_25_1067 ();
 sg13g2_decap_8 FILLER_25_1098 ();
 sg13g2_decap_8 FILLER_25_1105 ();
 sg13g2_decap_8 FILLER_25_1112 ();
 sg13g2_decap_8 FILLER_25_1119 ();
 sg13g2_decap_8 FILLER_25_1126 ();
 sg13g2_decap_4 FILLER_25_1133 ();
 sg13g2_fill_2 FILLER_25_1137 ();
 sg13g2_decap_8 FILLER_25_1143 ();
 sg13g2_decap_8 FILLER_25_1150 ();
 sg13g2_decap_8 FILLER_25_1157 ();
 sg13g2_decap_4 FILLER_25_1164 ();
 sg13g2_fill_2 FILLER_25_1197 ();
 sg13g2_decap_8 FILLER_25_1230 ();
 sg13g2_decap_8 FILLER_25_1237 ();
 sg13g2_decap_8 FILLER_25_1244 ();
 sg13g2_fill_1 FILLER_25_1256 ();
 sg13g2_decap_8 FILLER_25_1260 ();
 sg13g2_decap_8 FILLER_25_1267 ();
 sg13g2_decap_8 FILLER_25_1300 ();
 sg13g2_decap_8 FILLER_25_1307 ();
 sg13g2_decap_8 FILLER_25_1314 ();
 sg13g2_decap_8 FILLER_25_1321 ();
 sg13g2_decap_8 FILLER_25_1328 ();
 sg13g2_decap_8 FILLER_25_1335 ();
 sg13g2_decap_8 FILLER_25_1342 ();
 sg13g2_fill_1 FILLER_25_1349 ();
 sg13g2_decap_8 FILLER_25_1376 ();
 sg13g2_decap_8 FILLER_25_1383 ();
 sg13g2_decap_8 FILLER_25_1390 ();
 sg13g2_decap_8 FILLER_25_1397 ();
 sg13g2_decap_8 FILLER_25_1404 ();
 sg13g2_decap_8 FILLER_25_1411 ();
 sg13g2_decap_8 FILLER_25_1418 ();
 sg13g2_fill_1 FILLER_25_1425 ();
 sg13g2_fill_2 FILLER_25_1436 ();
 sg13g2_fill_1 FILLER_25_1438 ();
 sg13g2_decap_8 FILLER_25_1470 ();
 sg13g2_fill_2 FILLER_25_1481 ();
 sg13g2_fill_1 FILLER_25_1505 ();
 sg13g2_fill_2 FILLER_25_1525 ();
 sg13g2_fill_1 FILLER_25_1527 ();
 sg13g2_decap_8 FILLER_25_1540 ();
 sg13g2_fill_2 FILLER_25_1547 ();
 sg13g2_fill_2 FILLER_25_1553 ();
 sg13g2_fill_1 FILLER_25_1555 ();
 sg13g2_decap_8 FILLER_25_1564 ();
 sg13g2_decap_8 FILLER_25_1571 ();
 sg13g2_decap_8 FILLER_25_1578 ();
 sg13g2_decap_8 FILLER_25_1585 ();
 sg13g2_decap_8 FILLER_25_1596 ();
 sg13g2_decap_4 FILLER_25_1603 ();
 sg13g2_fill_2 FILLER_25_1612 ();
 sg13g2_decap_4 FILLER_25_1625 ();
 sg13g2_fill_2 FILLER_25_1629 ();
 sg13g2_decap_8 FILLER_25_1635 ();
 sg13g2_decap_8 FILLER_25_1642 ();
 sg13g2_decap_8 FILLER_25_1649 ();
 sg13g2_decap_8 FILLER_25_1656 ();
 sg13g2_fill_2 FILLER_25_1663 ();
 sg13g2_fill_1 FILLER_25_1665 ();
 sg13g2_fill_1 FILLER_25_1680 ();
 sg13g2_decap_8 FILLER_25_1685 ();
 sg13g2_decap_8 FILLER_25_1692 ();
 sg13g2_fill_2 FILLER_25_1699 ();
 sg13g2_decap_4 FILLER_25_1710 ();
 sg13g2_decap_4 FILLER_25_1726 ();
 sg13g2_decap_8 FILLER_25_1756 ();
 sg13g2_decap_8 FILLER_25_1763 ();
 sg13g2_decap_4 FILLER_25_1770 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_4 FILLER_26_21 ();
 sg13g2_fill_2 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_40 ();
 sg13g2_fill_2 FILLER_26_47 ();
 sg13g2_fill_1 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_55 ();
 sg13g2_decap_8 FILLER_26_62 ();
 sg13g2_decap_4 FILLER_26_73 ();
 sg13g2_fill_2 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_fill_2 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_119 ();
 sg13g2_decap_4 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_145 ();
 sg13g2_fill_1 FILLER_26_160 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_197 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_fill_2 FILLER_26_220 ();
 sg13g2_decap_4 FILLER_26_227 ();
 sg13g2_fill_2 FILLER_26_241 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_272 ();
 sg13g2_fill_2 FILLER_26_279 ();
 sg13g2_decap_4 FILLER_26_291 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_fill_2 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_fill_2 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_decap_4 FILLER_26_377 ();
 sg13g2_fill_1 FILLER_26_381 ();
 sg13g2_fill_2 FILLER_26_388 ();
 sg13g2_decap_4 FILLER_26_400 ();
 sg13g2_decap_8 FILLER_26_408 ();
 sg13g2_fill_2 FILLER_26_415 ();
 sg13g2_fill_1 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_442 ();
 sg13g2_decap_8 FILLER_26_451 ();
 sg13g2_decap_8 FILLER_26_458 ();
 sg13g2_fill_2 FILLER_26_465 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_fill_1 FILLER_26_518 ();
 sg13g2_decap_4 FILLER_26_560 ();
 sg13g2_decap_4 FILLER_26_570 ();
 sg13g2_fill_1 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_579 ();
 sg13g2_decap_8 FILLER_26_586 ();
 sg13g2_decap_8 FILLER_26_593 ();
 sg13g2_fill_1 FILLER_26_600 ();
 sg13g2_fill_2 FILLER_26_610 ();
 sg13g2_fill_1 FILLER_26_612 ();
 sg13g2_decap_4 FILLER_26_617 ();
 sg13g2_fill_2 FILLER_26_621 ();
 sg13g2_fill_2 FILLER_26_632 ();
 sg13g2_fill_1 FILLER_26_665 ();
 sg13g2_fill_1 FILLER_26_671 ();
 sg13g2_fill_1 FILLER_26_676 ();
 sg13g2_fill_1 FILLER_26_703 ();
 sg13g2_decap_4 FILLER_26_713 ();
 sg13g2_fill_1 FILLER_26_717 ();
 sg13g2_decap_4 FILLER_26_723 ();
 sg13g2_fill_1 FILLER_26_727 ();
 sg13g2_fill_2 FILLER_26_732 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_fill_2 FILLER_26_803 ();
 sg13g2_fill_1 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_fill_1 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_841 ();
 sg13g2_decap_8 FILLER_26_848 ();
 sg13g2_decap_8 FILLER_26_855 ();
 sg13g2_fill_1 FILLER_26_862 ();
 sg13g2_fill_2 FILLER_26_871 ();
 sg13g2_fill_1 FILLER_26_873 ();
 sg13g2_decap_8 FILLER_26_882 ();
 sg13g2_fill_2 FILLER_26_893 ();
 sg13g2_decap_8 FILLER_26_900 ();
 sg13g2_decap_8 FILLER_26_907 ();
 sg13g2_decap_8 FILLER_26_914 ();
 sg13g2_decap_8 FILLER_26_921 ();
 sg13g2_decap_8 FILLER_26_928 ();
 sg13g2_fill_2 FILLER_26_935 ();
 sg13g2_fill_1 FILLER_26_937 ();
 sg13g2_decap_4 FILLER_26_955 ();
 sg13g2_decap_8 FILLER_26_973 ();
 sg13g2_decap_4 FILLER_26_980 ();
 sg13g2_fill_2 FILLER_26_995 ();
 sg13g2_fill_1 FILLER_26_997 ();
 sg13g2_decap_4 FILLER_26_1003 ();
 sg13g2_fill_1 FILLER_26_1007 ();
 sg13g2_fill_1 FILLER_26_1012 ();
 sg13g2_fill_2 FILLER_26_1019 ();
 sg13g2_fill_1 FILLER_26_1021 ();
 sg13g2_fill_2 FILLER_26_1034 ();
 sg13g2_fill_2 FILLER_26_1052 ();
 sg13g2_fill_2 FILLER_26_1059 ();
 sg13g2_fill_1 FILLER_26_1079 ();
 sg13g2_decap_8 FILLER_26_1089 ();
 sg13g2_decap_8 FILLER_26_1096 ();
 sg13g2_decap_8 FILLER_26_1103 ();
 sg13g2_decap_8 FILLER_26_1114 ();
 sg13g2_decap_4 FILLER_26_1121 ();
 sg13g2_decap_8 FILLER_26_1158 ();
 sg13g2_decap_4 FILLER_26_1165 ();
 sg13g2_fill_2 FILLER_26_1169 ();
 sg13g2_fill_1 FILLER_26_1187 ();
 sg13g2_decap_8 FILLER_26_1204 ();
 sg13g2_fill_1 FILLER_26_1229 ();
 sg13g2_decap_8 FILLER_26_1237 ();
 sg13g2_decap_8 FILLER_26_1244 ();
 sg13g2_fill_2 FILLER_26_1251 ();
 sg13g2_fill_1 FILLER_26_1279 ();
 sg13g2_decap_8 FILLER_26_1284 ();
 sg13g2_decap_8 FILLER_26_1291 ();
 sg13g2_decap_8 FILLER_26_1298 ();
 sg13g2_decap_8 FILLER_26_1305 ();
 sg13g2_decap_4 FILLER_26_1312 ();
 sg13g2_decap_8 FILLER_26_1320 ();
 sg13g2_decap_8 FILLER_26_1327 ();
 sg13g2_decap_4 FILLER_26_1334 ();
 sg13g2_fill_2 FILLER_26_1342 ();
 sg13g2_fill_1 FILLER_26_1344 ();
 sg13g2_decap_4 FILLER_26_1354 ();
 sg13g2_decap_8 FILLER_26_1362 ();
 sg13g2_fill_1 FILLER_26_1369 ();
 sg13g2_decap_8 FILLER_26_1382 ();
 sg13g2_fill_2 FILLER_26_1389 ();
 sg13g2_fill_1 FILLER_26_1391 ();
 sg13g2_decap_8 FILLER_26_1396 ();
 sg13g2_decap_8 FILLER_26_1403 ();
 sg13g2_decap_8 FILLER_26_1410 ();
 sg13g2_decap_8 FILLER_26_1417 ();
 sg13g2_decap_8 FILLER_26_1424 ();
 sg13g2_fill_1 FILLER_26_1431 ();
 sg13g2_decap_8 FILLER_26_1436 ();
 sg13g2_decap_8 FILLER_26_1443 ();
 sg13g2_decap_8 FILLER_26_1450 ();
 sg13g2_decap_8 FILLER_26_1457 ();
 sg13g2_decap_8 FILLER_26_1464 ();
 sg13g2_decap_8 FILLER_26_1471 ();
 sg13g2_decap_8 FILLER_26_1478 ();
 sg13g2_decap_8 FILLER_26_1485 ();
 sg13g2_decap_8 FILLER_26_1492 ();
 sg13g2_decap_8 FILLER_26_1499 ();
 sg13g2_decap_8 FILLER_26_1506 ();
 sg13g2_decap_8 FILLER_26_1517 ();
 sg13g2_decap_8 FILLER_26_1524 ();
 sg13g2_decap_8 FILLER_26_1536 ();
 sg13g2_fill_1 FILLER_26_1543 ();
 sg13g2_decap_8 FILLER_26_1551 ();
 sg13g2_decap_8 FILLER_26_1558 ();
 sg13g2_decap_8 FILLER_26_1627 ();
 sg13g2_decap_4 FILLER_26_1634 ();
 sg13g2_fill_2 FILLER_26_1638 ();
 sg13g2_fill_1 FILLER_26_1666 ();
 sg13g2_fill_2 FILLER_26_1672 ();
 sg13g2_decap_4 FILLER_26_1682 ();
 sg13g2_fill_1 FILLER_26_1686 ();
 sg13g2_fill_2 FILLER_26_1704 ();
 sg13g2_decap_8 FILLER_26_1715 ();
 sg13g2_decap_8 FILLER_26_1722 ();
 sg13g2_decap_8 FILLER_26_1729 ();
 sg13g2_decap_8 FILLER_26_1736 ();
 sg13g2_decap_8 FILLER_26_1743 ();
 sg13g2_decap_8 FILLER_26_1750 ();
 sg13g2_decap_8 FILLER_26_1757 ();
 sg13g2_decap_8 FILLER_26_1764 ();
 sg13g2_fill_2 FILLER_26_1771 ();
 sg13g2_fill_1 FILLER_26_1773 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_35 ();
 sg13g2_fill_1 FILLER_27_37 ();
 sg13g2_decap_8 FILLER_27_46 ();
 sg13g2_decap_8 FILLER_27_53 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_decap_4 FILLER_27_66 ();
 sg13g2_fill_2 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_81 ();
 sg13g2_decap_8 FILLER_27_88 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_decap_4 FILLER_27_149 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_decap_4 FILLER_27_173 ();
 sg13g2_fill_2 FILLER_27_177 ();
 sg13g2_decap_4 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_decap_4 FILLER_27_228 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_decap_4 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_252 ();
 sg13g2_fill_1 FILLER_27_258 ();
 sg13g2_decap_8 FILLER_27_265 ();
 sg13g2_decap_8 FILLER_27_272 ();
 sg13g2_decap_4 FILLER_27_279 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_312 ();
 sg13g2_decap_8 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_4 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_decap_4 FILLER_27_363 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_397 ();
 sg13g2_fill_1 FILLER_27_404 ();
 sg13g2_decap_8 FILLER_27_418 ();
 sg13g2_fill_2 FILLER_27_425 ();
 sg13g2_fill_2 FILLER_27_444 ();
 sg13g2_decap_8 FILLER_27_464 ();
 sg13g2_decap_8 FILLER_27_471 ();
 sg13g2_decap_8 FILLER_27_478 ();
 sg13g2_decap_8 FILLER_27_485 ();
 sg13g2_decap_4 FILLER_27_492 ();
 sg13g2_fill_2 FILLER_27_496 ();
 sg13g2_fill_2 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_510 ();
 sg13g2_decap_8 FILLER_27_517 ();
 sg13g2_fill_1 FILLER_27_527 ();
 sg13g2_decap_8 FILLER_27_534 ();
 sg13g2_fill_2 FILLER_27_541 ();
 sg13g2_fill_2 FILLER_27_582 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_4 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_632 ();
 sg13g2_decap_8 FILLER_27_639 ();
 sg13g2_decap_8 FILLER_27_646 ();
 sg13g2_decap_8 FILLER_27_653 ();
 sg13g2_fill_2 FILLER_27_660 ();
 sg13g2_decap_8 FILLER_27_666 ();
 sg13g2_decap_8 FILLER_27_673 ();
 sg13g2_decap_8 FILLER_27_680 ();
 sg13g2_decap_8 FILLER_27_687 ();
 sg13g2_decap_8 FILLER_27_694 ();
 sg13g2_decap_4 FILLER_27_701 ();
 sg13g2_fill_2 FILLER_27_705 ();
 sg13g2_decap_4 FILLER_27_711 ();
 sg13g2_fill_2 FILLER_27_724 ();
 sg13g2_fill_2 FILLER_27_734 ();
 sg13g2_fill_1 FILLER_27_736 ();
 sg13g2_decap_4 FILLER_27_750 ();
 sg13g2_fill_1 FILLER_27_754 ();
 sg13g2_fill_1 FILLER_27_763 ();
 sg13g2_decap_4 FILLER_27_794 ();
 sg13g2_fill_1 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_825 ();
 sg13g2_decap_4 FILLER_27_832 ();
 sg13g2_fill_2 FILLER_27_836 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_8 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_decap_8 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_912 ();
 sg13g2_decap_8 FILLER_27_919 ();
 sg13g2_decap_8 FILLER_27_926 ();
 sg13g2_decap_8 FILLER_27_933 ();
 sg13g2_decap_8 FILLER_27_940 ();
 sg13g2_decap_8 FILLER_27_947 ();
 sg13g2_fill_2 FILLER_27_954 ();
 sg13g2_decap_8 FILLER_27_972 ();
 sg13g2_decap_8 FILLER_27_979 ();
 sg13g2_fill_2 FILLER_27_986 ();
 sg13g2_decap_8 FILLER_27_993 ();
 sg13g2_decap_8 FILLER_27_1000 ();
 sg13g2_decap_4 FILLER_27_1007 ();
 sg13g2_fill_1 FILLER_27_1021 ();
 sg13g2_decap_4 FILLER_27_1028 ();
 sg13g2_fill_1 FILLER_27_1032 ();
 sg13g2_decap_4 FILLER_27_1042 ();
 sg13g2_fill_1 FILLER_27_1046 ();
 sg13g2_fill_1 FILLER_27_1057 ();
 sg13g2_fill_1 FILLER_27_1063 ();
 sg13g2_decap_8 FILLER_27_1090 ();
 sg13g2_decap_8 FILLER_27_1097 ();
 sg13g2_fill_1 FILLER_27_1104 ();
 sg13g2_decap_8 FILLER_27_1120 ();
 sg13g2_fill_2 FILLER_27_1127 ();
 sg13g2_fill_1 FILLER_27_1129 ();
 sg13g2_fill_1 FILLER_27_1145 ();
 sg13g2_fill_2 FILLER_27_1172 ();
 sg13g2_fill_2 FILLER_27_1182 ();
 sg13g2_fill_2 FILLER_27_1201 ();
 sg13g2_fill_2 FILLER_27_1212 ();
 sg13g2_decap_8 FILLER_27_1228 ();
 sg13g2_fill_2 FILLER_27_1235 ();
 sg13g2_fill_1 FILLER_27_1260 ();
 sg13g2_decap_8 FILLER_27_1265 ();
 sg13g2_decap_8 FILLER_27_1272 ();
 sg13g2_decap_8 FILLER_27_1279 ();
 sg13g2_decap_8 FILLER_27_1286 ();
 sg13g2_decap_8 FILLER_27_1293 ();
 sg13g2_decap_8 FILLER_27_1313 ();
 sg13g2_decap_8 FILLER_27_1320 ();
 sg13g2_decap_8 FILLER_27_1327 ();
 sg13g2_decap_4 FILLER_27_1334 ();
 sg13g2_fill_1 FILLER_27_1338 ();
 sg13g2_fill_1 FILLER_27_1344 ();
 sg13g2_decap_8 FILLER_27_1357 ();
 sg13g2_decap_8 FILLER_27_1415 ();
 sg13g2_decap_4 FILLER_27_1422 ();
 sg13g2_decap_4 FILLER_27_1452 ();
 sg13g2_fill_1 FILLER_27_1456 ();
 sg13g2_fill_1 FILLER_27_1465 ();
 sg13g2_decap_4 FILLER_27_1477 ();
 sg13g2_fill_2 FILLER_27_1481 ();
 sg13g2_fill_1 FILLER_27_1488 ();
 sg13g2_fill_1 FILLER_27_1494 ();
 sg13g2_decap_8 FILLER_27_1508 ();
 sg13g2_fill_1 FILLER_27_1515 ();
 sg13g2_fill_1 FILLER_27_1521 ();
 sg13g2_fill_1 FILLER_27_1533 ();
 sg13g2_fill_1 FILLER_27_1540 ();
 sg13g2_fill_1 FILLER_27_1547 ();
 sg13g2_decap_8 FILLER_27_1553 ();
 sg13g2_decap_8 FILLER_27_1560 ();
 sg13g2_decap_8 FILLER_27_1567 ();
 sg13g2_decap_8 FILLER_27_1574 ();
 sg13g2_decap_8 FILLER_27_1581 ();
 sg13g2_decap_8 FILLER_27_1588 ();
 sg13g2_decap_8 FILLER_27_1595 ();
 sg13g2_decap_8 FILLER_27_1602 ();
 sg13g2_decap_8 FILLER_27_1609 ();
 sg13g2_decap_8 FILLER_27_1616 ();
 sg13g2_decap_4 FILLER_27_1623 ();
 sg13g2_fill_1 FILLER_27_1627 ();
 sg13g2_decap_8 FILLER_27_1632 ();
 sg13g2_decap_4 FILLER_27_1639 ();
 sg13g2_fill_1 FILLER_27_1643 ();
 sg13g2_decap_8 FILLER_27_1648 ();
 sg13g2_decap_8 FILLER_27_1655 ();
 sg13g2_decap_4 FILLER_27_1662 ();
 sg13g2_fill_1 FILLER_27_1666 ();
 sg13g2_decap_8 FILLER_27_1671 ();
 sg13g2_decap_8 FILLER_27_1678 ();
 sg13g2_decap_8 FILLER_27_1685 ();
 sg13g2_fill_2 FILLER_27_1692 ();
 sg13g2_decap_8 FILLER_27_1698 ();
 sg13g2_fill_2 FILLER_27_1713 ();
 sg13g2_decap_8 FILLER_27_1725 ();
 sg13g2_decap_8 FILLER_27_1732 ();
 sg13g2_decap_8 FILLER_27_1739 ();
 sg13g2_decap_8 FILLER_27_1746 ();
 sg13g2_decap_8 FILLER_27_1753 ();
 sg13g2_decap_8 FILLER_27_1760 ();
 sg13g2_decap_8 FILLER_27_1767 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_34 ();
 sg13g2_decap_4 FILLER_28_47 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_decap_4 FILLER_28_68 ();
 sg13g2_fill_2 FILLER_28_72 ();
 sg13g2_decap_4 FILLER_28_87 ();
 sg13g2_decap_4 FILLER_28_95 ();
 sg13g2_fill_1 FILLER_28_99 ();
 sg13g2_decap_8 FILLER_28_104 ();
 sg13g2_decap_8 FILLER_28_111 ();
 sg13g2_decap_8 FILLER_28_118 ();
 sg13g2_decap_8 FILLER_28_125 ();
 sg13g2_decap_4 FILLER_28_132 ();
 sg13g2_fill_2 FILLER_28_136 ();
 sg13g2_decap_8 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_165 ();
 sg13g2_decap_8 FILLER_28_180 ();
 sg13g2_decap_8 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_decap_4 FILLER_28_205 ();
 sg13g2_fill_2 FILLER_28_209 ();
 sg13g2_fill_2 FILLER_28_220 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_228 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_4 FILLER_28_248 ();
 sg13g2_decap_4 FILLER_28_257 ();
 sg13g2_fill_1 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_271 ();
 sg13g2_decap_4 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_285 ();
 sg13g2_decap_4 FILLER_28_291 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_decap_4 FILLER_28_307 ();
 sg13g2_fill_1 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_decap_4 FILLER_28_341 ();
 sg13g2_decap_4 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_387 ();
 sg13g2_fill_2 FILLER_28_393 ();
 sg13g2_fill_1 FILLER_28_395 ();
 sg13g2_fill_1 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_28_411 ();
 sg13g2_fill_2 FILLER_28_418 ();
 sg13g2_fill_2 FILLER_28_430 ();
 sg13g2_decap_4 FILLER_28_437 ();
 sg13g2_decap_8 FILLER_28_453 ();
 sg13g2_decap_8 FILLER_28_460 ();
 sg13g2_decap_8 FILLER_28_472 ();
 sg13g2_decap_8 FILLER_28_479 ();
 sg13g2_decap_8 FILLER_28_486 ();
 sg13g2_decap_4 FILLER_28_493 ();
 sg13g2_fill_2 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_fill_2 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_545 ();
 sg13g2_decap_4 FILLER_28_552 ();
 sg13g2_fill_2 FILLER_28_556 ();
 sg13g2_fill_2 FILLER_28_562 ();
 sg13g2_fill_1 FILLER_28_564 ();
 sg13g2_decap_4 FILLER_28_603 ();
 sg13g2_fill_1 FILLER_28_607 ();
 sg13g2_decap_8 FILLER_28_612 ();
 sg13g2_decap_8 FILLER_28_619 ();
 sg13g2_fill_1 FILLER_28_626 ();
 sg13g2_fill_1 FILLER_28_634 ();
 sg13g2_fill_1 FILLER_28_661 ();
 sg13g2_decap_4 FILLER_28_667 ();
 sg13g2_fill_2 FILLER_28_671 ();
 sg13g2_decap_8 FILLER_28_699 ();
 sg13g2_decap_4 FILLER_28_706 ();
 sg13g2_fill_1 FILLER_28_710 ();
 sg13g2_fill_2 FILLER_28_716 ();
 sg13g2_fill_1 FILLER_28_718 ();
 sg13g2_decap_8 FILLER_28_723 ();
 sg13g2_decap_8 FILLER_28_730 ();
 sg13g2_decap_4 FILLER_28_737 ();
 sg13g2_fill_1 FILLER_28_741 ();
 sg13g2_decap_8 FILLER_28_746 ();
 sg13g2_decap_8 FILLER_28_753 ();
 sg13g2_fill_1 FILLER_28_760 ();
 sg13g2_decap_4 FILLER_28_765 ();
 sg13g2_fill_2 FILLER_28_769 ();
 sg13g2_decap_8 FILLER_28_775 ();
 sg13g2_decap_8 FILLER_28_782 ();
 sg13g2_fill_2 FILLER_28_789 ();
 sg13g2_fill_1 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_808 ();
 sg13g2_decap_8 FILLER_28_815 ();
 sg13g2_fill_2 FILLER_28_822 ();
 sg13g2_decap_8 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_fill_1 FILLER_28_858 ();
 sg13g2_decap_4 FILLER_28_863 ();
 sg13g2_fill_2 FILLER_28_879 ();
 sg13g2_decap_4 FILLER_28_885 ();
 sg13g2_decap_8 FILLER_28_893 ();
 sg13g2_fill_2 FILLER_28_900 ();
 sg13g2_decap_8 FILLER_28_907 ();
 sg13g2_decap_8 FILLER_28_914 ();
 sg13g2_fill_1 FILLER_28_921 ();
 sg13g2_decap_8 FILLER_28_926 ();
 sg13g2_decap_8 FILLER_28_933 ();
 sg13g2_fill_2 FILLER_28_953 ();
 sg13g2_decap_8 FILLER_28_971 ();
 sg13g2_decap_8 FILLER_28_978 ();
 sg13g2_decap_4 FILLER_28_985 ();
 sg13g2_fill_2 FILLER_28_1005 ();
 sg13g2_decap_8 FILLER_28_1011 ();
 sg13g2_fill_2 FILLER_28_1018 ();
 sg13g2_fill_1 FILLER_28_1020 ();
 sg13g2_decap_8 FILLER_28_1029 ();
 sg13g2_decap_4 FILLER_28_1036 ();
 sg13g2_fill_2 FILLER_28_1040 ();
 sg13g2_decap_8 FILLER_28_1046 ();
 sg13g2_decap_8 FILLER_28_1053 ();
 sg13g2_decap_8 FILLER_28_1060 ();
 sg13g2_decap_4 FILLER_28_1067 ();
 sg13g2_fill_1 FILLER_28_1071 ();
 sg13g2_decap_8 FILLER_28_1091 ();
 sg13g2_decap_8 FILLER_28_1098 ();
 sg13g2_fill_2 FILLER_28_1105 ();
 sg13g2_decap_8 FILLER_28_1114 ();
 sg13g2_decap_8 FILLER_28_1121 ();
 sg13g2_decap_4 FILLER_28_1128 ();
 sg13g2_fill_2 FILLER_28_1147 ();
 sg13g2_fill_1 FILLER_28_1153 ();
 sg13g2_decap_8 FILLER_28_1158 ();
 sg13g2_decap_8 FILLER_28_1165 ();
 sg13g2_decap_8 FILLER_28_1172 ();
 sg13g2_decap_8 FILLER_28_1179 ();
 sg13g2_decap_8 FILLER_28_1186 ();
 sg13g2_decap_4 FILLER_28_1193 ();
 sg13g2_fill_2 FILLER_28_1212 ();
 sg13g2_decap_8 FILLER_28_1219 ();
 sg13g2_decap_8 FILLER_28_1226 ();
 sg13g2_fill_2 FILLER_28_1262 ();
 sg13g2_fill_1 FILLER_28_1264 ();
 sg13g2_decap_8 FILLER_28_1283 ();
 sg13g2_decap_8 FILLER_28_1290 ();
 sg13g2_decap_8 FILLER_28_1302 ();
 sg13g2_fill_1 FILLER_28_1309 ();
 sg13g2_decap_8 FILLER_28_1315 ();
 sg13g2_decap_8 FILLER_28_1322 ();
 sg13g2_decap_8 FILLER_28_1329 ();
 sg13g2_decap_8 FILLER_28_1336 ();
 sg13g2_decap_8 FILLER_28_1343 ();
 sg13g2_decap_8 FILLER_28_1350 ();
 sg13g2_decap_8 FILLER_28_1357 ();
 sg13g2_decap_8 FILLER_28_1364 ();
 sg13g2_fill_2 FILLER_28_1371 ();
 sg13g2_fill_1 FILLER_28_1373 ();
 sg13g2_decap_8 FILLER_28_1388 ();
 sg13g2_decap_4 FILLER_28_1395 ();
 sg13g2_fill_1 FILLER_28_1399 ();
 sg13g2_decap_8 FILLER_28_1407 ();
 sg13g2_decap_8 FILLER_28_1414 ();
 sg13g2_decap_8 FILLER_28_1421 ();
 sg13g2_fill_1 FILLER_28_1428 ();
 sg13g2_decap_8 FILLER_28_1434 ();
 sg13g2_decap_8 FILLER_28_1441 ();
 sg13g2_decap_8 FILLER_28_1448 ();
 sg13g2_decap_4 FILLER_28_1455 ();
 sg13g2_decap_4 FILLER_28_1474 ();
 sg13g2_decap_4 FILLER_28_1495 ();
 sg13g2_fill_1 FILLER_28_1499 ();
 sg13g2_decap_8 FILLER_28_1505 ();
 sg13g2_fill_2 FILLER_28_1512 ();
 sg13g2_fill_1 FILLER_28_1514 ();
 sg13g2_decap_8 FILLER_28_1520 ();
 sg13g2_decap_8 FILLER_28_1527 ();
 sg13g2_fill_1 FILLER_28_1534 ();
 sg13g2_fill_2 FILLER_28_1542 ();
 sg13g2_fill_1 FILLER_28_1544 ();
 sg13g2_fill_2 FILLER_28_1553 ();
 sg13g2_fill_1 FILLER_28_1555 ();
 sg13g2_decap_8 FILLER_28_1560 ();
 sg13g2_decap_8 FILLER_28_1567 ();
 sg13g2_decap_8 FILLER_28_1574 ();
 sg13g2_decap_8 FILLER_28_1581 ();
 sg13g2_fill_1 FILLER_28_1588 ();
 sg13g2_decap_4 FILLER_28_1593 ();
 sg13g2_fill_1 FILLER_28_1597 ();
 sg13g2_decap_8 FILLER_28_1624 ();
 sg13g2_decap_8 FILLER_28_1631 ();
 sg13g2_decap_8 FILLER_28_1638 ();
 sg13g2_decap_4 FILLER_28_1645 ();
 sg13g2_decap_8 FILLER_28_1653 ();
 sg13g2_decap_4 FILLER_28_1660 ();
 sg13g2_fill_1 FILLER_28_1664 ();
 sg13g2_decap_8 FILLER_28_1670 ();
 sg13g2_fill_2 FILLER_28_1677 ();
 sg13g2_fill_1 FILLER_28_1679 ();
 sg13g2_decap_8 FILLER_28_1684 ();
 sg13g2_fill_1 FILLER_28_1691 ();
 sg13g2_decap_8 FILLER_28_1695 ();
 sg13g2_decap_8 FILLER_28_1702 ();
 sg13g2_decap_8 FILLER_28_1709 ();
 sg13g2_decap_8 FILLER_28_1716 ();
 sg13g2_decap_8 FILLER_28_1723 ();
 sg13g2_decap_8 FILLER_28_1730 ();
 sg13g2_decap_8 FILLER_28_1737 ();
 sg13g2_decap_8 FILLER_28_1744 ();
 sg13g2_decap_8 FILLER_28_1751 ();
 sg13g2_decap_8 FILLER_28_1758 ();
 sg13g2_decap_8 FILLER_28_1765 ();
 sg13g2_fill_2 FILLER_28_1772 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_fill_2 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_44 ();
 sg13g2_decap_4 FILLER_29_54 ();
 sg13g2_fill_2 FILLER_29_58 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_75 ();
 sg13g2_fill_1 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_87 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_fill_1 FILLER_29_101 ();
 sg13g2_decap_4 FILLER_29_115 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_125 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_decap_8 FILLER_29_139 ();
 sg13g2_decap_4 FILLER_29_146 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_157 ();
 sg13g2_fill_2 FILLER_29_164 ();
 sg13g2_fill_1 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_decap_4 FILLER_29_195 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_decap_4 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_208 ();
 sg13g2_decap_4 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_218 ();
 sg13g2_decap_8 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_240 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_decap_4 FILLER_29_248 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_265 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_decap_4 FILLER_29_283 ();
 sg13g2_decap_4 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_300 ();
 sg13g2_decap_8 FILLER_29_307 ();
 sg13g2_decap_4 FILLER_29_314 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_decap_4 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_343 ();
 sg13g2_decap_4 FILLER_29_349 ();
 sg13g2_fill_2 FILLER_29_353 ();
 sg13g2_decap_8 FILLER_29_366 ();
 sg13g2_decap_8 FILLER_29_373 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_2 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_decap_4 FILLER_29_395 ();
 sg13g2_fill_2 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_29_414 ();
 sg13g2_fill_2 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_431 ();
 sg13g2_fill_1 FILLER_29_433 ();
 sg13g2_decap_8 FILLER_29_439 ();
 sg13g2_decap_8 FILLER_29_446 ();
 sg13g2_fill_1 FILLER_29_458 ();
 sg13g2_decap_8 FILLER_29_468 ();
 sg13g2_decap_8 FILLER_29_475 ();
 sg13g2_decap_8 FILLER_29_482 ();
 sg13g2_decap_8 FILLER_29_489 ();
 sg13g2_decap_8 FILLER_29_496 ();
 sg13g2_decap_8 FILLER_29_503 ();
 sg13g2_decap_8 FILLER_29_510 ();
 sg13g2_decap_8 FILLER_29_517 ();
 sg13g2_decap_4 FILLER_29_524 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_4 FILLER_29_546 ();
 sg13g2_fill_2 FILLER_29_550 ();
 sg13g2_fill_2 FILLER_29_557 ();
 sg13g2_decap_8 FILLER_29_576 ();
 sg13g2_decap_8 FILLER_29_583 ();
 sg13g2_decap_4 FILLER_29_590 ();
 sg13g2_fill_2 FILLER_29_594 ();
 sg13g2_decap_8 FILLER_29_627 ();
 sg13g2_decap_8 FILLER_29_634 ();
 sg13g2_decap_8 FILLER_29_645 ();
 sg13g2_decap_8 FILLER_29_652 ();
 sg13g2_decap_8 FILLER_29_659 ();
 sg13g2_decap_8 FILLER_29_666 ();
 sg13g2_decap_4 FILLER_29_673 ();
 sg13g2_fill_2 FILLER_29_677 ();
 sg13g2_decap_8 FILLER_29_683 ();
 sg13g2_decap_8 FILLER_29_690 ();
 sg13g2_decap_8 FILLER_29_697 ();
 sg13g2_fill_2 FILLER_29_704 ();
 sg13g2_decap_8 FILLER_29_718 ();
 sg13g2_decap_8 FILLER_29_725 ();
 sg13g2_decap_8 FILLER_29_732 ();
 sg13g2_decap_8 FILLER_29_739 ();
 sg13g2_fill_1 FILLER_29_751 ();
 sg13g2_decap_8 FILLER_29_778 ();
 sg13g2_decap_4 FILLER_29_785 ();
 sg13g2_decap_4 FILLER_29_820 ();
 sg13g2_decap_8 FILLER_29_829 ();
 sg13g2_fill_2 FILLER_29_836 ();
 sg13g2_decap_8 FILLER_29_869 ();
 sg13g2_fill_1 FILLER_29_881 ();
 sg13g2_fill_1 FILLER_29_941 ();
 sg13g2_decap_8 FILLER_29_972 ();
 sg13g2_decap_4 FILLER_29_979 ();
 sg13g2_fill_1 FILLER_29_983 ();
 sg13g2_fill_2 FILLER_29_1001 ();
 sg13g2_fill_1 FILLER_29_1003 ();
 sg13g2_decap_8 FILLER_29_1009 ();
 sg13g2_decap_8 FILLER_29_1016 ();
 sg13g2_decap_4 FILLER_29_1023 ();
 sg13g2_decap_8 FILLER_29_1059 ();
 sg13g2_decap_4 FILLER_29_1066 ();
 sg13g2_fill_2 FILLER_29_1070 ();
 sg13g2_decap_8 FILLER_29_1076 ();
 sg13g2_decap_8 FILLER_29_1083 ();
 sg13g2_decap_4 FILLER_29_1090 ();
 sg13g2_fill_2 FILLER_29_1094 ();
 sg13g2_decap_8 FILLER_29_1100 ();
 sg13g2_decap_8 FILLER_29_1116 ();
 sg13g2_decap_8 FILLER_29_1123 ();
 sg13g2_decap_8 FILLER_29_1130 ();
 sg13g2_decap_4 FILLER_29_1137 ();
 sg13g2_fill_2 FILLER_29_1153 ();
 sg13g2_decap_8 FILLER_29_1164 ();
 sg13g2_decap_8 FILLER_29_1171 ();
 sg13g2_decap_8 FILLER_29_1178 ();
 sg13g2_decap_4 FILLER_29_1185 ();
 sg13g2_fill_2 FILLER_29_1189 ();
 sg13g2_decap_8 FILLER_29_1208 ();
 sg13g2_decap_8 FILLER_29_1215 ();
 sg13g2_decap_8 FILLER_29_1222 ();
 sg13g2_decap_4 FILLER_29_1229 ();
 sg13g2_decap_8 FILLER_29_1247 ();
 sg13g2_fill_2 FILLER_29_1254 ();
 sg13g2_decap_8 FILLER_29_1261 ();
 sg13g2_decap_8 FILLER_29_1268 ();
 sg13g2_decap_8 FILLER_29_1275 ();
 sg13g2_decap_8 FILLER_29_1282 ();
 sg13g2_decap_8 FILLER_29_1289 ();
 sg13g2_fill_1 FILLER_29_1296 ();
 sg13g2_decap_8 FILLER_29_1315 ();
 sg13g2_decap_8 FILLER_29_1322 ();
 sg13g2_decap_4 FILLER_29_1329 ();
 sg13g2_fill_2 FILLER_29_1333 ();
 sg13g2_decap_8 FILLER_29_1365 ();
 sg13g2_decap_8 FILLER_29_1372 ();
 sg13g2_decap_8 FILLER_29_1379 ();
 sg13g2_decap_8 FILLER_29_1386 ();
 sg13g2_decap_8 FILLER_29_1393 ();
 sg13g2_fill_2 FILLER_29_1400 ();
 sg13g2_fill_1 FILLER_29_1402 ();
 sg13g2_decap_8 FILLER_29_1411 ();
 sg13g2_decap_4 FILLER_29_1418 ();
 sg13g2_decap_8 FILLER_29_1426 ();
 sg13g2_decap_8 FILLER_29_1433 ();
 sg13g2_decap_8 FILLER_29_1440 ();
 sg13g2_decap_8 FILLER_29_1447 ();
 sg13g2_decap_4 FILLER_29_1454 ();
 sg13g2_fill_1 FILLER_29_1458 ();
 sg13g2_decap_8 FILLER_29_1464 ();
 sg13g2_decap_4 FILLER_29_1471 ();
 sg13g2_fill_2 FILLER_29_1475 ();
 sg13g2_decap_4 FILLER_29_1493 ();
 sg13g2_decap_8 FILLER_29_1502 ();
 sg13g2_decap_8 FILLER_29_1513 ();
 sg13g2_decap_8 FILLER_29_1520 ();
 sg13g2_decap_8 FILLER_29_1527 ();
 sg13g2_decap_8 FILLER_29_1534 ();
 sg13g2_fill_2 FILLER_29_1541 ();
 sg13g2_fill_1 FILLER_29_1543 ();
 sg13g2_fill_2 FILLER_29_1550 ();
 sg13g2_fill_1 FILLER_29_1552 ();
 sg13g2_decap_8 FILLER_29_1560 ();
 sg13g2_decap_8 FILLER_29_1567 ();
 sg13g2_decap_8 FILLER_29_1574 ();
 sg13g2_decap_8 FILLER_29_1594 ();
 sg13g2_decap_4 FILLER_29_1601 ();
 sg13g2_fill_1 FILLER_29_1605 ();
 sg13g2_decap_8 FILLER_29_1610 ();
 sg13g2_decap_4 FILLER_29_1617 ();
 sg13g2_fill_1 FILLER_29_1621 ();
 sg13g2_decap_8 FILLER_29_1652 ();
 sg13g2_decap_4 FILLER_29_1659 ();
 sg13g2_fill_2 FILLER_29_1663 ();
 sg13g2_fill_2 FILLER_29_1671 ();
 sg13g2_decap_8 FILLER_29_1703 ();
 sg13g2_decap_4 FILLER_29_1710 ();
 sg13g2_fill_2 FILLER_29_1714 ();
 sg13g2_decap_8 FILLER_29_1746 ();
 sg13g2_decap_8 FILLER_29_1753 ();
 sg13g2_decap_8 FILLER_29_1760 ();
 sg13g2_decap_8 FILLER_29_1767 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_67 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_80 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_decap_4 FILLER_30_92 ();
 sg13g2_decap_4 FILLER_30_100 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_decap_4 FILLER_30_114 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_decap_4 FILLER_30_124 ();
 sg13g2_decap_4 FILLER_30_132 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_1 FILLER_30_141 ();
 sg13g2_decap_8 FILLER_30_151 ();
 sg13g2_decap_4 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_fill_2 FILLER_30_213 ();
 sg13g2_decap_4 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_4 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_289 ();
 sg13g2_fill_1 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_317 ();
 sg13g2_fill_1 FILLER_30_324 ();
 sg13g2_decap_4 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_379 ();
 sg13g2_fill_2 FILLER_30_385 ();
 sg13g2_fill_1 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_4 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_418 ();
 sg13g2_fill_2 FILLER_30_424 ();
 sg13g2_decap_4 FILLER_30_436 ();
 sg13g2_fill_2 FILLER_30_440 ();
 sg13g2_fill_1 FILLER_30_457 ();
 sg13g2_fill_2 FILLER_30_462 ();
 sg13g2_fill_1 FILLER_30_464 ();
 sg13g2_decap_8 FILLER_30_470 ();
 sg13g2_decap_8 FILLER_30_477 ();
 sg13g2_decap_8 FILLER_30_484 ();
 sg13g2_decap_8 FILLER_30_491 ();
 sg13g2_decap_4 FILLER_30_498 ();
 sg13g2_decap_4 FILLER_30_511 ();
 sg13g2_fill_1 FILLER_30_515 ();
 sg13g2_decap_4 FILLER_30_555 ();
 sg13g2_decap_8 FILLER_30_585 ();
 sg13g2_decap_8 FILLER_30_592 ();
 sg13g2_decap_8 FILLER_30_599 ();
 sg13g2_decap_8 FILLER_30_606 ();
 sg13g2_fill_2 FILLER_30_613 ();
 sg13g2_decap_8 FILLER_30_629 ();
 sg13g2_decap_8 FILLER_30_636 ();
 sg13g2_decap_4 FILLER_30_643 ();
 sg13g2_fill_2 FILLER_30_647 ();
 sg13g2_decap_8 FILLER_30_682 ();
 sg13g2_decap_8 FILLER_30_689 ();
 sg13g2_decap_4 FILLER_30_696 ();
 sg13g2_fill_1 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_709 ();
 sg13g2_decap_8 FILLER_30_716 ();
 sg13g2_decap_4 FILLER_30_723 ();
 sg13g2_decap_8 FILLER_30_731 ();
 sg13g2_fill_2 FILLER_30_738 ();
 sg13g2_fill_1 FILLER_30_740 ();
 sg13g2_fill_2 FILLER_30_744 ();
 sg13g2_decap_8 FILLER_30_750 ();
 sg13g2_decap_8 FILLER_30_757 ();
 sg13g2_decap_8 FILLER_30_764 ();
 sg13g2_decap_8 FILLER_30_771 ();
 sg13g2_decap_8 FILLER_30_778 ();
 sg13g2_fill_2 FILLER_30_785 ();
 sg13g2_decap_4 FILLER_30_791 ();
 sg13g2_fill_1 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_fill_2 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_853 ();
 sg13g2_decap_8 FILLER_30_860 ();
 sg13g2_decap_8 FILLER_30_867 ();
 sg13g2_decap_8 FILLER_30_883 ();
 sg13g2_decap_8 FILLER_30_890 ();
 sg13g2_decap_8 FILLER_30_897 ();
 sg13g2_decap_8 FILLER_30_904 ();
 sg13g2_decap_8 FILLER_30_911 ();
 sg13g2_decap_8 FILLER_30_918 ();
 sg13g2_decap_8 FILLER_30_925 ();
 sg13g2_decap_4 FILLER_30_932 ();
 sg13g2_fill_2 FILLER_30_936 ();
 sg13g2_fill_1 FILLER_30_943 ();
 sg13g2_decap_8 FILLER_30_950 ();
 sg13g2_decap_8 FILLER_30_957 ();
 sg13g2_decap_8 FILLER_30_964 ();
 sg13g2_decap_8 FILLER_30_971 ();
 sg13g2_decap_8 FILLER_30_978 ();
 sg13g2_fill_2 FILLER_30_985 ();
 sg13g2_decap_8 FILLER_30_1018 ();
 sg13g2_decap_8 FILLER_30_1025 ();
 sg13g2_decap_8 FILLER_30_1032 ();
 sg13g2_decap_8 FILLER_30_1039 ();
 sg13g2_decap_8 FILLER_30_1046 ();
 sg13g2_decap_8 FILLER_30_1053 ();
 sg13g2_decap_8 FILLER_30_1060 ();
 sg13g2_decap_8 FILLER_30_1067 ();
 sg13g2_decap_4 FILLER_30_1079 ();
 sg13g2_fill_1 FILLER_30_1083 ();
 sg13g2_decap_4 FILLER_30_1115 ();
 sg13g2_fill_1 FILLER_30_1119 ();
 sg13g2_decap_4 FILLER_30_1123 ();
 sg13g2_fill_2 FILLER_30_1127 ();
 sg13g2_decap_8 FILLER_30_1137 ();
 sg13g2_fill_2 FILLER_30_1144 ();
 sg13g2_fill_1 FILLER_30_1146 ();
 sg13g2_decap_4 FILLER_30_1154 ();
 sg13g2_fill_1 FILLER_30_1158 ();
 sg13g2_decap_8 FILLER_30_1164 ();
 sg13g2_decap_8 FILLER_30_1176 ();
 sg13g2_decap_8 FILLER_30_1183 ();
 sg13g2_decap_8 FILLER_30_1190 ();
 sg13g2_fill_2 FILLER_30_1197 ();
 sg13g2_decap_8 FILLER_30_1207 ();
 sg13g2_decap_4 FILLER_30_1214 ();
 sg13g2_fill_2 FILLER_30_1218 ();
 sg13g2_decap_8 FILLER_30_1224 ();
 sg13g2_decap_8 FILLER_30_1231 ();
 sg13g2_decap_8 FILLER_30_1267 ();
 sg13g2_decap_8 FILLER_30_1274 ();
 sg13g2_decap_8 FILLER_30_1281 ();
 sg13g2_decap_8 FILLER_30_1288 ();
 sg13g2_fill_2 FILLER_30_1295 ();
 sg13g2_decap_8 FILLER_30_1301 ();
 sg13g2_fill_2 FILLER_30_1308 ();
 sg13g2_fill_1 FILLER_30_1310 ();
 sg13g2_decap_8 FILLER_30_1337 ();
 sg13g2_decap_4 FILLER_30_1344 ();
 sg13g2_fill_1 FILLER_30_1348 ();
 sg13g2_fill_2 FILLER_30_1359 ();
 sg13g2_decap_8 FILLER_30_1366 ();
 sg13g2_fill_2 FILLER_30_1373 ();
 sg13g2_fill_1 FILLER_30_1396 ();
 sg13g2_decap_8 FILLER_30_1445 ();
 sg13g2_decap_4 FILLER_30_1452 ();
 sg13g2_fill_1 FILLER_30_1456 ();
 sg13g2_fill_1 FILLER_30_1463 ();
 sg13g2_fill_1 FILLER_30_1469 ();
 sg13g2_fill_1 FILLER_30_1480 ();
 sg13g2_fill_2 FILLER_30_1486 ();
 sg13g2_fill_1 FILLER_30_1488 ();
 sg13g2_decap_4 FILLER_30_1532 ();
 sg13g2_decap_8 FILLER_30_1548 ();
 sg13g2_fill_2 FILLER_30_1555 ();
 sg13g2_decap_8 FILLER_30_1568 ();
 sg13g2_decap_4 FILLER_30_1575 ();
 sg13g2_fill_1 FILLER_30_1579 ();
 sg13g2_decap_4 FILLER_30_1589 ();
 sg13g2_fill_2 FILLER_30_1593 ();
 sg13g2_decap_8 FILLER_30_1605 ();
 sg13g2_fill_1 FILLER_30_1612 ();
 sg13g2_decap_8 FILLER_30_1621 ();
 sg13g2_decap_8 FILLER_30_1628 ();
 sg13g2_decap_8 FILLER_30_1635 ();
 sg13g2_fill_1 FILLER_30_1642 ();
 sg13g2_fill_2 FILLER_30_1648 ();
 sg13g2_fill_1 FILLER_30_1650 ();
 sg13g2_fill_2 FILLER_30_1660 ();
 sg13g2_decap_8 FILLER_30_1688 ();
 sg13g2_decap_8 FILLER_30_1695 ();
 sg13g2_decap_8 FILLER_30_1702 ();
 sg13g2_decap_8 FILLER_30_1709 ();
 sg13g2_decap_4 FILLER_30_1716 ();
 sg13g2_fill_2 FILLER_30_1720 ();
 sg13g2_decap_8 FILLER_30_1736 ();
 sg13g2_decap_8 FILLER_30_1743 ();
 sg13g2_decap_8 FILLER_30_1750 ();
 sg13g2_decap_8 FILLER_30_1757 ();
 sg13g2_decap_8 FILLER_30_1764 ();
 sg13g2_fill_2 FILLER_30_1771 ();
 sg13g2_fill_1 FILLER_30_1773 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_16 ();
 sg13g2_fill_2 FILLER_31_43 ();
 sg13g2_fill_1 FILLER_31_45 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_decap_4 FILLER_31_62 ();
 sg13g2_fill_2 FILLER_31_66 ();
 sg13g2_decap_4 FILLER_31_73 ();
 sg13g2_fill_2 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_90 ();
 sg13g2_fill_2 FILLER_31_99 ();
 sg13g2_fill_1 FILLER_31_101 ();
 sg13g2_decap_4 FILLER_31_106 ();
 sg13g2_decap_4 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_134 ();
 sg13g2_decap_8 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_159 ();
 sg13g2_fill_2 FILLER_31_164 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_176 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_fill_1 FILLER_31_193 ();
 sg13g2_decap_4 FILLER_31_205 ();
 sg13g2_decap_8 FILLER_31_218 ();
 sg13g2_decap_4 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_decap_8 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_247 ();
 sg13g2_decap_4 FILLER_31_254 ();
 sg13g2_decap_4 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_8 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_310 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_4 FILLER_31_336 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_4 FILLER_31_402 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_decap_4 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_31_463 ();
 sg13g2_fill_1 FILLER_31_470 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_4 FILLER_31_504 ();
 sg13g2_fill_2 FILLER_31_508 ();
 sg13g2_decap_8 FILLER_31_516 ();
 sg13g2_decap_8 FILLER_31_523 ();
 sg13g2_decap_8 FILLER_31_530 ();
 sg13g2_decap_8 FILLER_31_537 ();
 sg13g2_decap_4 FILLER_31_544 ();
 sg13g2_fill_2 FILLER_31_553 ();
 sg13g2_decap_8 FILLER_31_564 ();
 sg13g2_decap_8 FILLER_31_571 ();
 sg13g2_decap_8 FILLER_31_583 ();
 sg13g2_decap_8 FILLER_31_590 ();
 sg13g2_decap_4 FILLER_31_597 ();
 sg13g2_fill_1 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_635 ();
 sg13g2_decap_8 FILLER_31_642 ();
 sg13g2_decap_8 FILLER_31_649 ();
 sg13g2_decap_4 FILLER_31_656 ();
 sg13g2_fill_2 FILLER_31_660 ();
 sg13g2_decap_8 FILLER_31_666 ();
 sg13g2_decap_4 FILLER_31_673 ();
 sg13g2_fill_2 FILLER_31_677 ();
 sg13g2_decap_4 FILLER_31_700 ();
 sg13g2_fill_2 FILLER_31_704 ();
 sg13g2_fill_1 FILLER_31_711 ();
 sg13g2_fill_2 FILLER_31_717 ();
 sg13g2_decap_8 FILLER_31_747 ();
 sg13g2_decap_8 FILLER_31_754 ();
 sg13g2_decap_8 FILLER_31_761 ();
 sg13g2_decap_4 FILLER_31_768 ();
 sg13g2_fill_1 FILLER_31_772 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_4 FILLER_31_784 ();
 sg13g2_fill_1 FILLER_31_788 ();
 sg13g2_fill_2 FILLER_31_793 ();
 sg13g2_fill_1 FILLER_31_795 ();
 sg13g2_decap_4 FILLER_31_801 ();
 sg13g2_fill_1 FILLER_31_805 ();
 sg13g2_fill_2 FILLER_31_809 ();
 sg13g2_fill_1 FILLER_31_811 ();
 sg13g2_decap_8 FILLER_31_846 ();
 sg13g2_decap_8 FILLER_31_853 ();
 sg13g2_decap_8 FILLER_31_860 ();
 sg13g2_decap_4 FILLER_31_867 ();
 sg13g2_decap_8 FILLER_31_881 ();
 sg13g2_decap_4 FILLER_31_888 ();
 sg13g2_fill_2 FILLER_31_902 ();
 sg13g2_fill_1 FILLER_31_904 ();
 sg13g2_decap_8 FILLER_31_910 ();
 sg13g2_decap_8 FILLER_31_917 ();
 sg13g2_decap_8 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_4 FILLER_31_938 ();
 sg13g2_fill_2 FILLER_31_942 ();
 sg13g2_decap_8 FILLER_31_950 ();
 sg13g2_decap_8 FILLER_31_957 ();
 sg13g2_decap_8 FILLER_31_964 ();
 sg13g2_decap_8 FILLER_31_971 ();
 sg13g2_fill_2 FILLER_31_978 ();
 sg13g2_decap_8 FILLER_31_991 ();
 sg13g2_decap_8 FILLER_31_998 ();
 sg13g2_decap_8 FILLER_31_1005 ();
 sg13g2_decap_8 FILLER_31_1012 ();
 sg13g2_fill_2 FILLER_31_1019 ();
 sg13g2_fill_1 FILLER_31_1021 ();
 sg13g2_decap_4 FILLER_31_1026 ();
 sg13g2_decap_8 FILLER_31_1036 ();
 sg13g2_fill_1 FILLER_31_1043 ();
 sg13g2_decap_8 FILLER_31_1048 ();
 sg13g2_decap_8 FILLER_31_1055 ();
 sg13g2_decap_8 FILLER_31_1062 ();
 sg13g2_decap_8 FILLER_31_1069 ();
 sg13g2_fill_1 FILLER_31_1076 ();
 sg13g2_decap_8 FILLER_31_1118 ();
 sg13g2_decap_8 FILLER_31_1125 ();
 sg13g2_decap_4 FILLER_31_1132 ();
 sg13g2_fill_1 FILLER_31_1144 ();
 sg13g2_decap_4 FILLER_31_1171 ();
 sg13g2_fill_1 FILLER_31_1175 ();
 sg13g2_fill_1 FILLER_31_1181 ();
 sg13g2_decap_8 FILLER_31_1190 ();
 sg13g2_decap_8 FILLER_31_1197 ();
 sg13g2_decap_8 FILLER_31_1204 ();
 sg13g2_fill_2 FILLER_31_1211 ();
 sg13g2_decap_8 FILLER_31_1217 ();
 sg13g2_decap_8 FILLER_31_1224 ();
 sg13g2_fill_2 FILLER_31_1231 ();
 sg13g2_fill_2 FILLER_31_1265 ();
 sg13g2_fill_1 FILLER_31_1267 ();
 sg13g2_fill_2 FILLER_31_1282 ();
 sg13g2_decap_4 FILLER_31_1289 ();
 sg13g2_decap_8 FILLER_31_1297 ();
 sg13g2_decap_8 FILLER_31_1304 ();
 sg13g2_decap_4 FILLER_31_1311 ();
 sg13g2_fill_2 FILLER_31_1324 ();
 sg13g2_fill_1 FILLER_31_1326 ();
 sg13g2_fill_2 FILLER_31_1330 ();
 sg13g2_fill_1 FILLER_31_1332 ();
 sg13g2_decap_8 FILLER_31_1344 ();
 sg13g2_decap_4 FILLER_31_1351 ();
 sg13g2_fill_1 FILLER_31_1355 ();
 sg13g2_decap_8 FILLER_31_1365 ();
 sg13g2_fill_1 FILLER_31_1372 ();
 sg13g2_decap_4 FILLER_31_1383 ();
 sg13g2_fill_2 FILLER_31_1387 ();
 sg13g2_decap_8 FILLER_31_1393 ();
 sg13g2_decap_4 FILLER_31_1400 ();
 sg13g2_decap_4 FILLER_31_1412 ();
 sg13g2_fill_2 FILLER_31_1416 ();
 sg13g2_decap_8 FILLER_31_1423 ();
 sg13g2_fill_1 FILLER_31_1430 ();
 sg13g2_decap_8 FILLER_31_1443 ();
 sg13g2_decap_8 FILLER_31_1450 ();
 sg13g2_decap_4 FILLER_31_1457 ();
 sg13g2_decap_8 FILLER_31_1471 ();
 sg13g2_fill_1 FILLER_31_1478 ();
 sg13g2_decap_8 FILLER_31_1483 ();
 sg13g2_fill_2 FILLER_31_1490 ();
 sg13g2_decap_8 FILLER_31_1517 ();
 sg13g2_decap_8 FILLER_31_1524 ();
 sg13g2_decap_8 FILLER_31_1531 ();
 sg13g2_decap_8 FILLER_31_1538 ();
 sg13g2_decap_8 FILLER_31_1545 ();
 sg13g2_decap_8 FILLER_31_1552 ();
 sg13g2_decap_8 FILLER_31_1559 ();
 sg13g2_decap_4 FILLER_31_1566 ();
 sg13g2_fill_2 FILLER_31_1570 ();
 sg13g2_decap_8 FILLER_31_1589 ();
 sg13g2_decap_8 FILLER_31_1596 ();
 sg13g2_fill_2 FILLER_31_1611 ();
 sg13g2_fill_2 FILLER_31_1618 ();
 sg13g2_decap_8 FILLER_31_1624 ();
 sg13g2_decap_8 FILLER_31_1631 ();
 sg13g2_decap_8 FILLER_31_1638 ();
 sg13g2_fill_2 FILLER_31_1645 ();
 sg13g2_fill_2 FILLER_31_1665 ();
 sg13g2_fill_1 FILLER_31_1667 ();
 sg13g2_decap_8 FILLER_31_1700 ();
 sg13g2_decap_8 FILLER_31_1707 ();
 sg13g2_fill_2 FILLER_31_1714 ();
 sg13g2_decap_4 FILLER_31_1721 ();
 sg13g2_decap_8 FILLER_31_1736 ();
 sg13g2_decap_8 FILLER_31_1743 ();
 sg13g2_decap_8 FILLER_31_1750 ();
 sg13g2_decap_8 FILLER_31_1757 ();
 sg13g2_decap_8 FILLER_31_1764 ();
 sg13g2_fill_2 FILLER_31_1771 ();
 sg13g2_fill_1 FILLER_31_1773 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_27 ();
 sg13g2_fill_1 FILLER_32_31 ();
 sg13g2_decap_8 FILLER_32_39 ();
 sg13g2_decap_8 FILLER_32_46 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_decap_8 FILLER_32_59 ();
 sg13g2_decap_8 FILLER_32_66 ();
 sg13g2_decap_8 FILLER_32_73 ();
 sg13g2_decap_8 FILLER_32_80 ();
 sg13g2_fill_2 FILLER_32_87 ();
 sg13g2_decap_8 FILLER_32_93 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_153 ();
 sg13g2_decap_8 FILLER_32_160 ();
 sg13g2_decap_8 FILLER_32_167 ();
 sg13g2_decap_8 FILLER_32_174 ();
 sg13g2_decap_8 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_188 ();
 sg13g2_decap_8 FILLER_32_195 ();
 sg13g2_decap_8 FILLER_32_202 ();
 sg13g2_decap_8 FILLER_32_209 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_248 ();
 sg13g2_decap_8 FILLER_32_255 ();
 sg13g2_fill_2 FILLER_32_262 ();
 sg13g2_decap_4 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_303 ();
 sg13g2_decap_4 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_decap_4 FILLER_32_320 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_fill_1 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_345 ();
 sg13g2_decap_8 FILLER_32_352 ();
 sg13g2_fill_2 FILLER_32_359 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_4 FILLER_32_396 ();
 sg13g2_fill_1 FILLER_32_400 ();
 sg13g2_fill_1 FILLER_32_405 ();
 sg13g2_fill_1 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_416 ();
 sg13g2_fill_1 FILLER_32_423 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_fill_2 FILLER_32_442 ();
 sg13g2_fill_2 FILLER_32_451 ();
 sg13g2_fill_1 FILLER_32_456 ();
 sg13g2_fill_1 FILLER_32_461 ();
 sg13g2_decap_8 FILLER_32_472 ();
 sg13g2_decap_8 FILLER_32_479 ();
 sg13g2_decap_4 FILLER_32_486 ();
 sg13g2_fill_1 FILLER_32_546 ();
 sg13g2_fill_1 FILLER_32_577 ();
 sg13g2_fill_2 FILLER_32_582 ();
 sg13g2_fill_1 FILLER_32_584 ();
 sg13g2_decap_8 FILLER_32_650 ();
 sg13g2_decap_8 FILLER_32_657 ();
 sg13g2_fill_2 FILLER_32_664 ();
 sg13g2_fill_1 FILLER_32_666 ();
 sg13g2_decap_8 FILLER_32_680 ();
 sg13g2_decap_8 FILLER_32_687 ();
 sg13g2_decap_8 FILLER_32_694 ();
 sg13g2_decap_8 FILLER_32_709 ();
 sg13g2_fill_2 FILLER_32_716 ();
 sg13g2_fill_2 FILLER_32_722 ();
 sg13g2_fill_1 FILLER_32_724 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_fill_1 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_741 ();
 sg13g2_decap_8 FILLER_32_748 ();
 sg13g2_fill_1 FILLER_32_755 ();
 sg13g2_fill_2 FILLER_32_763 ();
 sg13g2_fill_1 FILLER_32_765 ();
 sg13g2_decap_8 FILLER_32_792 ();
 sg13g2_decap_4 FILLER_32_807 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_decap_4 FILLER_32_822 ();
 sg13g2_fill_2 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_832 ();
 sg13g2_decap_8 FILLER_32_839 ();
 sg13g2_fill_2 FILLER_32_846 ();
 sg13g2_decap_8 FILLER_32_851 ();
 sg13g2_decap_8 FILLER_32_858 ();
 sg13g2_decap_8 FILLER_32_865 ();
 sg13g2_fill_2 FILLER_32_872 ();
 sg13g2_decap_4 FILLER_32_885 ();
 sg13g2_fill_2 FILLER_32_889 ();
 sg13g2_decap_4 FILLER_32_934 ();
 sg13g2_fill_1 FILLER_32_938 ();
 sg13g2_fill_1 FILLER_32_944 ();
 sg13g2_decap_8 FILLER_32_951 ();
 sg13g2_decap_8 FILLER_32_958 ();
 sg13g2_decap_8 FILLER_32_965 ();
 sg13g2_decap_8 FILLER_32_972 ();
 sg13g2_fill_1 FILLER_32_983 ();
 sg13g2_decap_8 FILLER_32_990 ();
 sg13g2_decap_4 FILLER_32_997 ();
 sg13g2_fill_1 FILLER_32_1001 ();
 sg13g2_decap_8 FILLER_32_1007 ();
 sg13g2_decap_4 FILLER_32_1014 ();
 sg13g2_fill_1 FILLER_32_1018 ();
 sg13g2_fill_1 FILLER_32_1033 ();
 sg13g2_decap_8 FILLER_32_1063 ();
 sg13g2_decap_8 FILLER_32_1070 ();
 sg13g2_decap_8 FILLER_32_1077 ();
 sg13g2_fill_1 FILLER_32_1096 ();
 sg13g2_fill_1 FILLER_32_1101 ();
 sg13g2_decap_8 FILLER_32_1106 ();
 sg13g2_decap_8 FILLER_32_1113 ();
 sg13g2_decap_8 FILLER_32_1120 ();
 sg13g2_decap_8 FILLER_32_1127 ();
 sg13g2_decap_8 FILLER_32_1134 ();
 sg13g2_decap_8 FILLER_32_1141 ();
 sg13g2_decap_4 FILLER_32_1148 ();
 sg13g2_decap_8 FILLER_32_1156 ();
 sg13g2_decap_8 FILLER_32_1163 ();
 sg13g2_fill_2 FILLER_32_1170 ();
 sg13g2_fill_1 FILLER_32_1172 ();
 sg13g2_decap_4 FILLER_32_1199 ();
 sg13g2_fill_2 FILLER_32_1203 ();
 sg13g2_decap_8 FILLER_32_1210 ();
 sg13g2_decap_8 FILLER_32_1217 ();
 sg13g2_decap_4 FILLER_32_1224 ();
 sg13g2_fill_2 FILLER_32_1228 ();
 sg13g2_fill_1 FILLER_32_1239 ();
 sg13g2_decap_4 FILLER_32_1248 ();
 sg13g2_decap_8 FILLER_32_1256 ();
 sg13g2_decap_8 FILLER_32_1263 ();
 sg13g2_decap_8 FILLER_32_1270 ();
 sg13g2_decap_8 FILLER_32_1277 ();
 sg13g2_decap_8 FILLER_32_1284 ();
 sg13g2_decap_8 FILLER_32_1291 ();
 sg13g2_decap_8 FILLER_32_1298 ();
 sg13g2_decap_8 FILLER_32_1305 ();
 sg13g2_decap_8 FILLER_32_1332 ();
 sg13g2_decap_4 FILLER_32_1339 ();
 sg13g2_fill_1 FILLER_32_1343 ();
 sg13g2_fill_1 FILLER_32_1349 ();
 sg13g2_decap_4 FILLER_32_1362 ();
 sg13g2_fill_2 FILLER_32_1366 ();
 sg13g2_decap_8 FILLER_32_1376 ();
 sg13g2_fill_2 FILLER_32_1383 ();
 sg13g2_fill_1 FILLER_32_1385 ();
 sg13g2_decap_8 FILLER_32_1391 ();
 sg13g2_decap_8 FILLER_32_1398 ();
 sg13g2_decap_4 FILLER_32_1411 ();
 sg13g2_fill_1 FILLER_32_1418 ();
 sg13g2_decap_4 FILLER_32_1424 ();
 sg13g2_fill_2 FILLER_32_1428 ();
 sg13g2_decap_8 FILLER_32_1442 ();
 sg13g2_decap_8 FILLER_32_1449 ();
 sg13g2_decap_8 FILLER_32_1456 ();
 sg13g2_fill_1 FILLER_32_1463 ();
 sg13g2_decap_4 FILLER_32_1468 ();
 sg13g2_decap_4 FILLER_32_1502 ();
 sg13g2_decap_8 FILLER_32_1536 ();
 sg13g2_decap_4 FILLER_32_1543 ();
 sg13g2_fill_2 FILLER_32_1547 ();
 sg13g2_decap_4 FILLER_32_1568 ();
 sg13g2_fill_2 FILLER_32_1572 ();
 sg13g2_fill_2 FILLER_32_1579 ();
 sg13g2_fill_2 FILLER_32_1588 ();
 sg13g2_fill_1 FILLER_32_1595 ();
 sg13g2_decap_8 FILLER_32_1605 ();
 sg13g2_decap_8 FILLER_32_1612 ();
 sg13g2_decap_8 FILLER_32_1619 ();
 sg13g2_fill_1 FILLER_32_1626 ();
 sg13g2_decap_8 FILLER_32_1641 ();
 sg13g2_fill_2 FILLER_32_1652 ();
 sg13g2_fill_1 FILLER_32_1654 ();
 sg13g2_decap_8 FILLER_32_1659 ();
 sg13g2_decap_8 FILLER_32_1666 ();
 sg13g2_decap_8 FILLER_32_1673 ();
 sg13g2_decap_8 FILLER_32_1680 ();
 sg13g2_decap_8 FILLER_32_1687 ();
 sg13g2_decap_8 FILLER_32_1694 ();
 sg13g2_decap_4 FILLER_32_1701 ();
 sg13g2_decap_8 FILLER_32_1713 ();
 sg13g2_decap_4 FILLER_32_1720 ();
 sg13g2_fill_2 FILLER_32_1739 ();
 sg13g2_fill_2 FILLER_32_1771 ();
 sg13g2_fill_1 FILLER_32_1773 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_fill_2 FILLER_33_32 ();
 sg13g2_decap_4 FILLER_33_46 ();
 sg13g2_fill_1 FILLER_33_50 ();
 sg13g2_decap_8 FILLER_33_64 ();
 sg13g2_fill_2 FILLER_33_71 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_95 ();
 sg13g2_decap_8 FILLER_33_102 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_decap_4 FILLER_33_115 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_130 ();
 sg13g2_decap_4 FILLER_33_137 ();
 sg13g2_decap_8 FILLER_33_162 ();
 sg13g2_decap_8 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_184 ();
 sg13g2_decap_4 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_decap_4 FILLER_33_255 ();
 sg13g2_decap_8 FILLER_33_267 ();
 sg13g2_decap_8 FILLER_33_274 ();
 sg13g2_decap_4 FILLER_33_281 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_decap_8 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_336 ();
 sg13g2_decap_4 FILLER_33_351 ();
 sg13g2_decap_4 FILLER_33_363 ();
 sg13g2_decap_8 FILLER_33_375 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_fill_1 FILLER_33_403 ();
 sg13g2_decap_8 FILLER_33_410 ();
 sg13g2_decap_8 FILLER_33_417 ();
 sg13g2_decap_8 FILLER_33_424 ();
 sg13g2_fill_2 FILLER_33_431 ();
 sg13g2_fill_1 FILLER_33_443 ();
 sg13g2_decap_8 FILLER_33_463 ();
 sg13g2_fill_1 FILLER_33_470 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_fill_1 FILLER_33_511 ();
 sg13g2_decap_4 FILLER_33_516 ();
 sg13g2_fill_2 FILLER_33_520 ();
 sg13g2_decap_8 FILLER_33_526 ();
 sg13g2_decap_8 FILLER_33_533 ();
 sg13g2_decap_8 FILLER_33_540 ();
 sg13g2_decap_8 FILLER_33_547 ();
 sg13g2_fill_2 FILLER_33_554 ();
 sg13g2_fill_1 FILLER_33_556 ();
 sg13g2_decap_8 FILLER_33_564 ();
 sg13g2_decap_8 FILLER_33_571 ();
 sg13g2_decap_8 FILLER_33_578 ();
 sg13g2_decap_8 FILLER_33_594 ();
 sg13g2_decap_8 FILLER_33_601 ();
 sg13g2_decap_4 FILLER_33_608 ();
 sg13g2_fill_1 FILLER_33_619 ();
 sg13g2_fill_2 FILLER_33_625 ();
 sg13g2_decap_8 FILLER_33_636 ();
 sg13g2_decap_8 FILLER_33_643 ();
 sg13g2_decap_4 FILLER_33_650 ();
 sg13g2_fill_2 FILLER_33_654 ();
 sg13g2_fill_2 FILLER_33_687 ();
 sg13g2_fill_1 FILLER_33_689 ();
 sg13g2_decap_4 FILLER_33_694 ();
 sg13g2_fill_2 FILLER_33_698 ();
 sg13g2_decap_8 FILLER_33_704 ();
 sg13g2_decap_8 FILLER_33_711 ();
 sg13g2_fill_2 FILLER_33_718 ();
 sg13g2_decap_4 FILLER_33_729 ();
 sg13g2_fill_1 FILLER_33_733 ();
 sg13g2_decap_8 FILLER_33_739 ();
 sg13g2_fill_1 FILLER_33_746 ();
 sg13g2_decap_8 FILLER_33_753 ();
 sg13g2_decap_8 FILLER_33_760 ();
 sg13g2_decap_8 FILLER_33_767 ();
 sg13g2_decap_8 FILLER_33_774 ();
 sg13g2_decap_8 FILLER_33_781 ();
 sg13g2_fill_2 FILLER_33_788 ();
 sg13g2_fill_1 FILLER_33_790 ();
 sg13g2_fill_2 FILLER_33_799 ();
 sg13g2_decap_8 FILLER_33_820 ();
 sg13g2_fill_1 FILLER_33_827 ();
 sg13g2_decap_8 FILLER_33_832 ();
 sg13g2_decap_8 FILLER_33_839 ();
 sg13g2_fill_2 FILLER_33_846 ();
 sg13g2_decap_8 FILLER_33_855 ();
 sg13g2_decap_4 FILLER_33_862 ();
 sg13g2_fill_1 FILLER_33_866 ();
 sg13g2_decap_8 FILLER_33_876 ();
 sg13g2_fill_1 FILLER_33_883 ();
 sg13g2_decap_4 FILLER_33_897 ();
 sg13g2_fill_1 FILLER_33_901 ();
 sg13g2_fill_2 FILLER_33_930 ();
 sg13g2_fill_1 FILLER_33_932 ();
 sg13g2_decap_8 FILLER_33_942 ();
 sg13g2_decap_8 FILLER_33_949 ();
 sg13g2_decap_8 FILLER_33_956 ();
 sg13g2_decap_8 FILLER_33_963 ();
 sg13g2_decap_4 FILLER_33_970 ();
 sg13g2_fill_2 FILLER_33_974 ();
 sg13g2_fill_1 FILLER_33_989 ();
 sg13g2_decap_8 FILLER_33_994 ();
 sg13g2_decap_8 FILLER_33_1001 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_decap_8 FILLER_33_1015 ();
 sg13g2_fill_1 FILLER_33_1022 ();
 sg13g2_decap_8 FILLER_33_1028 ();
 sg13g2_decap_4 FILLER_33_1050 ();
 sg13g2_fill_1 FILLER_33_1054 ();
 sg13g2_decap_8 FILLER_33_1067 ();
 sg13g2_decap_8 FILLER_33_1074 ();
 sg13g2_fill_1 FILLER_33_1081 ();
 sg13g2_fill_1 FILLER_33_1092 ();
 sg13g2_decap_4 FILLER_33_1096 ();
 sg13g2_fill_1 FILLER_33_1100 ();
 sg13g2_decap_8 FILLER_33_1116 ();
 sg13g2_decap_8 FILLER_33_1123 ();
 sg13g2_decap_4 FILLER_33_1130 ();
 sg13g2_fill_2 FILLER_33_1134 ();
 sg13g2_fill_2 FILLER_33_1174 ();
 sg13g2_decap_8 FILLER_33_1194 ();
 sg13g2_decap_4 FILLER_33_1201 ();
 sg13g2_fill_1 FILLER_33_1205 ();
 sg13g2_decap_8 FILLER_33_1215 ();
 sg13g2_decap_8 FILLER_33_1222 ();
 sg13g2_fill_1 FILLER_33_1229 ();
 sg13g2_decap_8 FILLER_33_1240 ();
 sg13g2_decap_8 FILLER_33_1247 ();
 sg13g2_fill_2 FILLER_33_1254 ();
 sg13g2_fill_1 FILLER_33_1256 ();
 sg13g2_fill_1 FILLER_33_1261 ();
 sg13g2_fill_2 FILLER_33_1266 ();
 sg13g2_fill_1 FILLER_33_1268 ();
 sg13g2_decap_8 FILLER_33_1273 ();
 sg13g2_fill_1 FILLER_33_1280 ();
 sg13g2_fill_2 FILLER_33_1290 ();
 sg13g2_fill_1 FILLER_33_1292 ();
 sg13g2_fill_2 FILLER_33_1298 ();
 sg13g2_decap_4 FILLER_33_1305 ();
 sg13g2_fill_2 FILLER_33_1317 ();
 sg13g2_decap_4 FILLER_33_1327 ();
 sg13g2_decap_4 FILLER_33_1337 ();
 sg13g2_decap_8 FILLER_33_1347 ();
 sg13g2_fill_1 FILLER_33_1354 ();
 sg13g2_decap_8 FILLER_33_1360 ();
 sg13g2_decap_4 FILLER_33_1367 ();
 sg13g2_fill_2 FILLER_33_1382 ();
 sg13g2_fill_1 FILLER_33_1384 ();
 sg13g2_decap_8 FILLER_33_1393 ();
 sg13g2_decap_4 FILLER_33_1400 ();
 sg13g2_fill_1 FILLER_33_1404 ();
 sg13g2_fill_2 FILLER_33_1411 ();
 sg13g2_fill_1 FILLER_33_1413 ();
 sg13g2_decap_4 FILLER_33_1420 ();
 sg13g2_fill_2 FILLER_33_1424 ();
 sg13g2_decap_8 FILLER_33_1434 ();
 sg13g2_decap_8 FILLER_33_1441 ();
 sg13g2_decap_8 FILLER_33_1448 ();
 sg13g2_decap_8 FILLER_33_1455 ();
 sg13g2_decap_8 FILLER_33_1462 ();
 sg13g2_decap_8 FILLER_33_1469 ();
 sg13g2_decap_8 FILLER_33_1476 ();
 sg13g2_decap_8 FILLER_33_1483 ();
 sg13g2_decap_8 FILLER_33_1490 ();
 sg13g2_decap_8 FILLER_33_1497 ();
 sg13g2_fill_2 FILLER_33_1504 ();
 sg13g2_fill_2 FILLER_33_1519 ();
 sg13g2_decap_8 FILLER_33_1525 ();
 sg13g2_decap_8 FILLER_33_1532 ();
 sg13g2_decap_8 FILLER_33_1539 ();
 sg13g2_decap_8 FILLER_33_1546 ();
 sg13g2_decap_4 FILLER_33_1553 ();
 sg13g2_fill_2 FILLER_33_1557 ();
 sg13g2_decap_4 FILLER_33_1567 ();
 sg13g2_fill_1 FILLER_33_1571 ();
 sg13g2_decap_8 FILLER_33_1577 ();
 sg13g2_decap_8 FILLER_33_1589 ();
 sg13g2_decap_8 FILLER_33_1596 ();
 sg13g2_fill_2 FILLER_33_1603 ();
 sg13g2_decap_8 FILLER_33_1609 ();
 sg13g2_decap_8 FILLER_33_1616 ();
 sg13g2_decap_4 FILLER_33_1623 ();
 sg13g2_fill_1 FILLER_33_1640 ();
 sg13g2_decap_8 FILLER_33_1667 ();
 sg13g2_decap_8 FILLER_33_1674 ();
 sg13g2_fill_1 FILLER_33_1681 ();
 sg13g2_fill_1 FILLER_33_1691 ();
 sg13g2_decap_8 FILLER_33_1696 ();
 sg13g2_decap_4 FILLER_33_1703 ();
 sg13g2_fill_2 FILLER_33_1716 ();
 sg13g2_fill_1 FILLER_33_1718 ();
 sg13g2_fill_1 FILLER_33_1724 ();
 sg13g2_fill_2 FILLER_33_1739 ();
 sg13g2_decap_8 FILLER_33_1754 ();
 sg13g2_decap_8 FILLER_33_1761 ();
 sg13g2_decap_4 FILLER_33_1768 ();
 sg13g2_fill_2 FILLER_33_1772 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_11 ();
 sg13g2_fill_2 FILLER_34_16 ();
 sg13g2_fill_1 FILLER_34_18 ();
 sg13g2_fill_2 FILLER_34_63 ();
 sg13g2_fill_1 FILLER_34_65 ();
 sg13g2_decap_4 FILLER_34_92 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_123 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_fill_2 FILLER_34_156 ();
 sg13g2_decap_8 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_decap_8 FILLER_34_179 ();
 sg13g2_decap_8 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_34_193 ();
 sg13g2_decap_8 FILLER_34_200 ();
 sg13g2_decap_4 FILLER_34_207 ();
 sg13g2_fill_1 FILLER_34_211 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_227 ();
 sg13g2_decap_8 FILLER_34_234 ();
 sg13g2_decap_8 FILLER_34_241 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_255 ();
 sg13g2_fill_2 FILLER_34_262 ();
 sg13g2_fill_1 FILLER_34_264 ();
 sg13g2_decap_8 FILLER_34_270 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_decap_4 FILLER_34_305 ();
 sg13g2_fill_2 FILLER_34_309 ();
 sg13g2_decap_8 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_345 ();
 sg13g2_decap_8 FILLER_34_352 ();
 sg13g2_decap_8 FILLER_34_359 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_decap_4 FILLER_34_380 ();
 sg13g2_fill_2 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_390 ();
 sg13g2_decap_4 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_401 ();
 sg13g2_decap_8 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_34_412 ();
 sg13g2_decap_8 FILLER_34_419 ();
 sg13g2_decap_4 FILLER_34_426 ();
 sg13g2_fill_2 FILLER_34_430 ();
 sg13g2_fill_2 FILLER_34_442 ();
 sg13g2_decap_4 FILLER_34_447 ();
 sg13g2_fill_2 FILLER_34_451 ();
 sg13g2_decap_8 FILLER_34_456 ();
 sg13g2_fill_2 FILLER_34_463 ();
 sg13g2_fill_1 FILLER_34_465 ();
 sg13g2_decap_4 FILLER_34_471 ();
 sg13g2_fill_2 FILLER_34_475 ();
 sg13g2_decap_8 FILLER_34_495 ();
 sg13g2_decap_4 FILLER_34_502 ();
 sg13g2_fill_2 FILLER_34_506 ();
 sg13g2_decap_8 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_532 ();
 sg13g2_decap_8 FILLER_34_539 ();
 sg13g2_decap_8 FILLER_34_546 ();
 sg13g2_decap_8 FILLER_34_553 ();
 sg13g2_decap_8 FILLER_34_560 ();
 sg13g2_decap_8 FILLER_34_567 ();
 sg13g2_decap_8 FILLER_34_574 ();
 sg13g2_decap_8 FILLER_34_581 ();
 sg13g2_decap_8 FILLER_34_588 ();
 sg13g2_fill_1 FILLER_34_595 ();
 sg13g2_decap_8 FILLER_34_600 ();
 sg13g2_fill_2 FILLER_34_607 ();
 sg13g2_decap_8 FILLER_34_614 ();
 sg13g2_decap_8 FILLER_34_621 ();
 sg13g2_decap_8 FILLER_34_628 ();
 sg13g2_decap_8 FILLER_34_635 ();
 sg13g2_decap_8 FILLER_34_642 ();
 sg13g2_decap_8 FILLER_34_649 ();
 sg13g2_decap_4 FILLER_34_656 ();
 sg13g2_fill_2 FILLER_34_660 ();
 sg13g2_decap_8 FILLER_34_666 ();
 sg13g2_decap_8 FILLER_34_673 ();
 sg13g2_decap_4 FILLER_34_680 ();
 sg13g2_fill_1 FILLER_34_684 ();
 sg13g2_fill_2 FILLER_34_697 ();
 sg13g2_fill_1 FILLER_34_699 ();
 sg13g2_decap_8 FILLER_34_712 ();
 sg13g2_decap_8 FILLER_34_719 ();
 sg13g2_decap_8 FILLER_34_726 ();
 sg13g2_fill_1 FILLER_34_733 ();
 sg13g2_fill_2 FILLER_34_744 ();
 sg13g2_fill_1 FILLER_34_746 ();
 sg13g2_decap_8 FILLER_34_765 ();
 sg13g2_decap_8 FILLER_34_772 ();
 sg13g2_decap_8 FILLER_34_779 ();
 sg13g2_decap_4 FILLER_34_786 ();
 sg13g2_fill_1 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_decap_8 FILLER_34_840 ();
 sg13g2_fill_2 FILLER_34_847 ();
 sg13g2_fill_1 FILLER_34_849 ();
 sg13g2_fill_1 FILLER_34_858 ();
 sg13g2_decap_8 FILLER_34_868 ();
 sg13g2_decap_8 FILLER_34_875 ();
 sg13g2_decap_8 FILLER_34_882 ();
 sg13g2_decap_8 FILLER_34_889 ();
 sg13g2_fill_2 FILLER_34_896 ();
 sg13g2_fill_1 FILLER_34_898 ();
 sg13g2_fill_1 FILLER_34_905 ();
 sg13g2_decap_8 FILLER_34_912 ();
 sg13g2_decap_8 FILLER_34_919 ();
 sg13g2_fill_2 FILLER_34_930 ();
 sg13g2_fill_1 FILLER_34_932 ();
 sg13g2_decap_8 FILLER_34_941 ();
 sg13g2_decap_4 FILLER_34_953 ();
 sg13g2_decap_8 FILLER_34_965 ();
 sg13g2_decap_8 FILLER_34_972 ();
 sg13g2_decap_4 FILLER_34_982 ();
 sg13g2_fill_2 FILLER_34_986 ();
 sg13g2_decap_4 FILLER_34_992 ();
 sg13g2_decap_8 FILLER_34_1000 ();
 sg13g2_decap_4 FILLER_34_1007 ();
 sg13g2_fill_1 FILLER_34_1011 ();
 sg13g2_fill_2 FILLER_34_1027 ();
 sg13g2_fill_1 FILLER_34_1037 ();
 sg13g2_decap_4 FILLER_34_1044 ();
 sg13g2_fill_2 FILLER_34_1053 ();
 sg13g2_decap_8 FILLER_34_1060 ();
 sg13g2_decap_8 FILLER_34_1067 ();
 sg13g2_decap_4 FILLER_34_1074 ();
 sg13g2_fill_1 FILLER_34_1078 ();
 sg13g2_fill_1 FILLER_34_1089 ();
 sg13g2_fill_2 FILLER_34_1099 ();
 sg13g2_decap_8 FILLER_34_1110 ();
 sg13g2_decap_8 FILLER_34_1117 ();
 sg13g2_fill_2 FILLER_34_1124 ();
 sg13g2_decap_8 FILLER_34_1147 ();
 sg13g2_decap_8 FILLER_34_1154 ();
 sg13g2_fill_2 FILLER_34_1161 ();
 sg13g2_fill_1 FILLER_34_1163 ();
 sg13g2_fill_2 FILLER_34_1172 ();
 sg13g2_fill_2 FILLER_34_1179 ();
 sg13g2_decap_8 FILLER_34_1195 ();
 sg13g2_decap_4 FILLER_34_1202 ();
 sg13g2_fill_2 FILLER_34_1206 ();
 sg13g2_decap_4 FILLER_34_1212 ();
 sg13g2_fill_1 FILLER_34_1216 ();
 sg13g2_fill_1 FILLER_34_1222 ();
 sg13g2_fill_2 FILLER_34_1228 ();
 sg13g2_fill_1 FILLER_34_1230 ();
 sg13g2_decap_4 FILLER_34_1236 ();
 sg13g2_fill_2 FILLER_34_1240 ();
 sg13g2_fill_2 FILLER_34_1246 ();
 sg13g2_fill_1 FILLER_34_1248 ();
 sg13g2_decap_8 FILLER_34_1254 ();
 sg13g2_fill_2 FILLER_34_1269 ();
 sg13g2_fill_2 FILLER_34_1282 ();
 sg13g2_fill_1 FILLER_34_1284 ();
 sg13g2_decap_8 FILLER_34_1303 ();
 sg13g2_decap_8 FILLER_34_1310 ();
 sg13g2_decap_4 FILLER_34_1317 ();
 sg13g2_fill_2 FILLER_34_1321 ();
 sg13g2_fill_2 FILLER_34_1341 ();
 sg13g2_fill_1 FILLER_34_1343 ();
 sg13g2_decap_8 FILLER_34_1349 ();
 sg13g2_decap_8 FILLER_34_1356 ();
 sg13g2_decap_4 FILLER_34_1363 ();
 sg13g2_fill_1 FILLER_34_1367 ();
 sg13g2_decap_4 FILLER_34_1379 ();
 sg13g2_fill_1 FILLER_34_1383 ();
 sg13g2_fill_2 FILLER_34_1388 ();
 sg13g2_decap_8 FILLER_34_1394 ();
 sg13g2_decap_4 FILLER_34_1401 ();
 sg13g2_fill_2 FILLER_34_1405 ();
 sg13g2_decap_8 FILLER_34_1413 ();
 sg13g2_decap_8 FILLER_34_1420 ();
 sg13g2_decap_8 FILLER_34_1427 ();
 sg13g2_decap_8 FILLER_34_1434 ();
 sg13g2_decap_4 FILLER_34_1441 ();
 sg13g2_decap_8 FILLER_34_1489 ();
 sg13g2_decap_8 FILLER_34_1496 ();
 sg13g2_fill_2 FILLER_34_1503 ();
 sg13g2_decap_4 FILLER_34_1520 ();
 sg13g2_decap_8 FILLER_34_1578 ();
 sg13g2_decap_8 FILLER_34_1589 ();
 sg13g2_decap_4 FILLER_34_1596 ();
 sg13g2_fill_2 FILLER_34_1600 ();
 sg13g2_decap_8 FILLER_34_1610 ();
 sg13g2_decap_8 FILLER_34_1617 ();
 sg13g2_decap_4 FILLER_34_1624 ();
 sg13g2_fill_2 FILLER_34_1628 ();
 sg13g2_fill_2 FILLER_34_1635 ();
 sg13g2_fill_1 FILLER_34_1637 ();
 sg13g2_decap_8 FILLER_34_1641 ();
 sg13g2_decap_8 FILLER_34_1648 ();
 sg13g2_fill_2 FILLER_34_1655 ();
 sg13g2_fill_1 FILLER_34_1657 ();
 sg13g2_decap_8 FILLER_34_1662 ();
 sg13g2_decap_4 FILLER_34_1669 ();
 sg13g2_fill_1 FILLER_34_1673 ();
 sg13g2_decap_4 FILLER_34_1679 ();
 sg13g2_fill_1 FILLER_34_1683 ();
 sg13g2_decap_8 FILLER_34_1692 ();
 sg13g2_decap_8 FILLER_34_1699 ();
 sg13g2_decap_4 FILLER_34_1714 ();
 sg13g2_fill_2 FILLER_34_1718 ();
 sg13g2_decap_8 FILLER_34_1742 ();
 sg13g2_decap_8 FILLER_34_1749 ();
 sg13g2_decap_8 FILLER_34_1756 ();
 sg13g2_decap_8 FILLER_34_1763 ();
 sg13g2_decap_4 FILLER_34_1770 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_109 ();
 sg13g2_decap_8 FILLER_35_116 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_decap_8 FILLER_35_130 ();
 sg13g2_decap_8 FILLER_35_137 ();
 sg13g2_fill_1 FILLER_35_144 ();
 sg13g2_decap_8 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_156 ();
 sg13g2_decap_8 FILLER_35_163 ();
 sg13g2_decap_8 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_decap_8 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_191 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_decap_8 FILLER_35_205 ();
 sg13g2_decap_8 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_219 ();
 sg13g2_decap_8 FILLER_35_226 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_244 ();
 sg13g2_decap_8 FILLER_35_251 ();
 sg13g2_decap_8 FILLER_35_258 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_272 ();
 sg13g2_decap_8 FILLER_35_279 ();
 sg13g2_fill_1 FILLER_35_286 ();
 sg13g2_decap_8 FILLER_35_362 ();
 sg13g2_decap_8 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_376 ();
 sg13g2_fill_1 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_410 ();
 sg13g2_decap_8 FILLER_35_417 ();
 sg13g2_fill_2 FILLER_35_424 ();
 sg13g2_fill_1 FILLER_35_426 ();
 sg13g2_decap_8 FILLER_35_453 ();
 sg13g2_decap_8 FILLER_35_460 ();
 sg13g2_fill_2 FILLER_35_467 ();
 sg13g2_fill_1 FILLER_35_495 ();
 sg13g2_fill_1 FILLER_35_500 ();
 sg13g2_fill_2 FILLER_35_505 ();
 sg13g2_decap_4 FILLER_35_546 ();
 sg13g2_fill_2 FILLER_35_550 ();
 sg13g2_decap_4 FILLER_35_583 ();
 sg13g2_fill_1 FILLER_35_587 ();
 sg13g2_decap_8 FILLER_35_614 ();
 sg13g2_decap_8 FILLER_35_621 ();
 sg13g2_decap_4 FILLER_35_628 ();
 sg13g2_decap_8 FILLER_35_658 ();
 sg13g2_decap_4 FILLER_35_665 ();
 sg13g2_fill_2 FILLER_35_669 ();
 sg13g2_decap_8 FILLER_35_684 ();
 sg13g2_decap_8 FILLER_35_691 ();
 sg13g2_fill_2 FILLER_35_698 ();
 sg13g2_fill_1 FILLER_35_700 ();
 sg13g2_fill_1 FILLER_35_714 ();
 sg13g2_fill_2 FILLER_35_718 ();
 sg13g2_fill_1 FILLER_35_720 ();
 sg13g2_fill_2 FILLER_35_729 ();
 sg13g2_fill_1 FILLER_35_731 ();
 sg13g2_decap_8 FILLER_35_740 ();
 sg13g2_decap_8 FILLER_35_747 ();
 sg13g2_decap_4 FILLER_35_754 ();
 sg13g2_fill_2 FILLER_35_758 ();
 sg13g2_decap_8 FILLER_35_765 ();
 sg13g2_decap_8 FILLER_35_772 ();
 sg13g2_fill_2 FILLER_35_779 ();
 sg13g2_fill_1 FILLER_35_781 ();
 sg13g2_fill_2 FILLER_35_795 ();
 sg13g2_fill_1 FILLER_35_797 ();
 sg13g2_decap_8 FILLER_35_825 ();
 sg13g2_decap_4 FILLER_35_832 ();
 sg13g2_fill_1 FILLER_35_836 ();
 sg13g2_fill_1 FILLER_35_863 ();
 sg13g2_fill_1 FILLER_35_875 ();
 sg13g2_fill_1 FILLER_35_881 ();
 sg13g2_fill_1 FILLER_35_887 ();
 sg13g2_fill_2 FILLER_35_897 ();
 sg13g2_fill_1 FILLER_35_899 ();
 sg13g2_decap_8 FILLER_35_914 ();
 sg13g2_decap_8 FILLER_35_921 ();
 sg13g2_fill_2 FILLER_35_928 ();
 sg13g2_fill_1 FILLER_35_930 ();
 sg13g2_fill_2 FILLER_35_942 ();
 sg13g2_fill_1 FILLER_35_944 ();
 sg13g2_decap_8 FILLER_35_961 ();
 sg13g2_fill_2 FILLER_35_968 ();
 sg13g2_decap_4 FILLER_35_988 ();
 sg13g2_fill_1 FILLER_35_992 ();
 sg13g2_decap_4 FILLER_35_998 ();
 sg13g2_fill_1 FILLER_35_1002 ();
 sg13g2_decap_4 FILLER_35_1007 ();
 sg13g2_decap_8 FILLER_35_1025 ();
 sg13g2_fill_2 FILLER_35_1032 ();
 sg13g2_fill_1 FILLER_35_1034 ();
 sg13g2_fill_1 FILLER_35_1042 ();
 sg13g2_decap_8 FILLER_35_1049 ();
 sg13g2_decap_8 FILLER_35_1056 ();
 sg13g2_decap_8 FILLER_35_1063 ();
 sg13g2_decap_8 FILLER_35_1070 ();
 sg13g2_decap_8 FILLER_35_1077 ();
 sg13g2_decap_4 FILLER_35_1084 ();
 sg13g2_fill_2 FILLER_35_1088 ();
 sg13g2_decap_8 FILLER_35_1105 ();
 sg13g2_decap_8 FILLER_35_1112 ();
 sg13g2_decap_4 FILLER_35_1119 ();
 sg13g2_fill_1 FILLER_35_1123 ();
 sg13g2_fill_1 FILLER_35_1129 ();
 sg13g2_decap_8 FILLER_35_1148 ();
 sg13g2_fill_2 FILLER_35_1155 ();
 sg13g2_fill_1 FILLER_35_1157 ();
 sg13g2_fill_1 FILLER_35_1179 ();
 sg13g2_fill_1 FILLER_35_1186 ();
 sg13g2_decap_4 FILLER_35_1191 ();
 sg13g2_fill_2 FILLER_35_1195 ();
 sg13g2_decap_4 FILLER_35_1202 ();
 sg13g2_fill_2 FILLER_35_1206 ();
 sg13g2_fill_2 FILLER_35_1213 ();
 sg13g2_fill_1 FILLER_35_1215 ();
 sg13g2_decap_8 FILLER_35_1220 ();
 sg13g2_decap_8 FILLER_35_1227 ();
 sg13g2_decap_4 FILLER_35_1234 ();
 sg13g2_fill_2 FILLER_35_1238 ();
 sg13g2_decap_8 FILLER_35_1245 ();
 sg13g2_fill_2 FILLER_35_1252 ();
 sg13g2_fill_1 FILLER_35_1254 ();
 sg13g2_decap_8 FILLER_35_1285 ();
 sg13g2_decap_8 FILLER_35_1292 ();
 sg13g2_decap_8 FILLER_35_1299 ();
 sg13g2_decap_8 FILLER_35_1306 ();
 sg13g2_decap_4 FILLER_35_1313 ();
 sg13g2_fill_2 FILLER_35_1317 ();
 sg13g2_fill_1 FILLER_35_1333 ();
 sg13g2_decap_8 FILLER_35_1345 ();
 sg13g2_fill_2 FILLER_35_1357 ();
 sg13g2_fill_1 FILLER_35_1359 ();
 sg13g2_fill_1 FILLER_35_1364 ();
 sg13g2_fill_2 FILLER_35_1379 ();
 sg13g2_fill_1 FILLER_35_1381 ();
 sg13g2_fill_2 FILLER_35_1391 ();
 sg13g2_decap_4 FILLER_35_1396 ();
 sg13g2_decap_4 FILLER_35_1403 ();
 sg13g2_decap_8 FILLER_35_1434 ();
 sg13g2_decap_4 FILLER_35_1441 ();
 sg13g2_fill_1 FILLER_35_1445 ();
 sg13g2_fill_2 FILLER_35_1450 ();
 sg13g2_fill_1 FILLER_35_1452 ();
 sg13g2_fill_2 FILLER_35_1461 ();
 sg13g2_fill_1 FILLER_35_1463 ();
 sg13g2_decap_8 FILLER_35_1473 ();
 sg13g2_decap_8 FILLER_35_1480 ();
 sg13g2_decap_8 FILLER_35_1487 ();
 sg13g2_decap_8 FILLER_35_1494 ();
 sg13g2_decap_4 FILLER_35_1501 ();
 sg13g2_decap_8 FILLER_35_1509 ();
 sg13g2_decap_4 FILLER_35_1516 ();
 sg13g2_fill_1 FILLER_35_1520 ();
 sg13g2_decap_8 FILLER_35_1526 ();
 sg13g2_decap_8 FILLER_35_1533 ();
 sg13g2_fill_1 FILLER_35_1540 ();
 sg13g2_decap_8 FILLER_35_1545 ();
 sg13g2_decap_8 FILLER_35_1552 ();
 sg13g2_decap_8 FILLER_35_1559 ();
 sg13g2_decap_4 FILLER_35_1566 ();
 sg13g2_fill_2 FILLER_35_1570 ();
 sg13g2_fill_2 FILLER_35_1576 ();
 sg13g2_decap_8 FILLER_35_1583 ();
 sg13g2_decap_8 FILLER_35_1590 ();
 sg13g2_decap_4 FILLER_35_1597 ();
 sg13g2_fill_1 FILLER_35_1637 ();
 sg13g2_fill_1 FILLER_35_1646 ();
 sg13g2_decap_4 FILLER_35_1651 ();
 sg13g2_fill_1 FILLER_35_1655 ();
 sg13g2_fill_2 FILLER_35_1669 ();
 sg13g2_fill_1 FILLER_35_1671 ();
 sg13g2_decap_8 FILLER_35_1676 ();
 sg13g2_fill_1 FILLER_35_1683 ();
 sg13g2_decap_8 FILLER_35_1692 ();
 sg13g2_decap_8 FILLER_35_1699 ();
 sg13g2_decap_8 FILLER_35_1710 ();
 sg13g2_decap_8 FILLER_35_1717 ();
 sg13g2_decap_8 FILLER_35_1737 ();
 sg13g2_decap_8 FILLER_35_1744 ();
 sg13g2_decap_8 FILLER_35_1751 ();
 sg13g2_decap_8 FILLER_35_1758 ();
 sg13g2_decap_8 FILLER_35_1765 ();
 sg13g2_fill_2 FILLER_35_1772 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_4 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_25 ();
 sg13g2_decap_4 FILLER_36_53 ();
 sg13g2_fill_2 FILLER_36_57 ();
 sg13g2_fill_2 FILLER_36_89 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_decap_8 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_decap_8 FILLER_36_164 ();
 sg13g2_decap_4 FILLER_36_171 ();
 sg13g2_fill_2 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_decap_8 FILLER_36_236 ();
 sg13g2_decap_8 FILLER_36_243 ();
 sg13g2_fill_2 FILLER_36_250 ();
 sg13g2_fill_1 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_257 ();
 sg13g2_decap_8 FILLER_36_264 ();
 sg13g2_decap_8 FILLER_36_271 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_decap_8 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_decap_4 FILLER_36_306 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_decap_4 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_decap_8 FILLER_36_346 ();
 sg13g2_decap_8 FILLER_36_353 ();
 sg13g2_decap_8 FILLER_36_360 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_fill_1 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_8 FILLER_36_424 ();
 sg13g2_decap_4 FILLER_36_431 ();
 sg13g2_decap_8 FILLER_36_439 ();
 sg13g2_decap_8 FILLER_36_446 ();
 sg13g2_decap_8 FILLER_36_453 ();
 sg13g2_decap_8 FILLER_36_460 ();
 sg13g2_decap_8 FILLER_36_467 ();
 sg13g2_decap_8 FILLER_36_474 ();
 sg13g2_decap_8 FILLER_36_481 ();
 sg13g2_decap_4 FILLER_36_488 ();
 sg13g2_decap_8 FILLER_36_507 ();
 sg13g2_decap_8 FILLER_36_514 ();
 sg13g2_decap_8 FILLER_36_521 ();
 sg13g2_decap_8 FILLER_36_528 ();
 sg13g2_decap_8 FILLER_36_535 ();
 sg13g2_decap_8 FILLER_36_542 ();
 sg13g2_decap_8 FILLER_36_549 ();
 sg13g2_fill_2 FILLER_36_556 ();
 sg13g2_decap_8 FILLER_36_562 ();
 sg13g2_decap_8 FILLER_36_569 ();
 sg13g2_decap_8 FILLER_36_576 ();
 sg13g2_decap_8 FILLER_36_583 ();
 sg13g2_decap_8 FILLER_36_590 ();
 sg13g2_decap_8 FILLER_36_597 ();
 sg13g2_decap_8 FILLER_36_604 ();
 sg13g2_decap_8 FILLER_36_611 ();
 sg13g2_decap_8 FILLER_36_618 ();
 sg13g2_decap_8 FILLER_36_625 ();
 sg13g2_decap_4 FILLER_36_632 ();
 sg13g2_fill_1 FILLER_36_636 ();
 sg13g2_decap_8 FILLER_36_641 ();
 sg13g2_decap_4 FILLER_36_648 ();
 sg13g2_fill_1 FILLER_36_652 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_fill_1 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_699 ();
 sg13g2_decap_4 FILLER_36_706 ();
 sg13g2_fill_1 FILLER_36_710 ();
 sg13g2_fill_2 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_738 ();
 sg13g2_decap_8 FILLER_36_745 ();
 sg13g2_decap_8 FILLER_36_752 ();
 sg13g2_decap_8 FILLER_36_759 ();
 sg13g2_decap_8 FILLER_36_766 ();
 sg13g2_decap_8 FILLER_36_773 ();
 sg13g2_fill_2 FILLER_36_780 ();
 sg13g2_decap_8 FILLER_36_795 ();
 sg13g2_decap_8 FILLER_36_802 ();
 sg13g2_decap_4 FILLER_36_809 ();
 sg13g2_fill_2 FILLER_36_813 ();
 sg13g2_decap_8 FILLER_36_827 ();
 sg13g2_fill_2 FILLER_36_834 ();
 sg13g2_fill_1 FILLER_36_836 ();
 sg13g2_fill_1 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_858 ();
 sg13g2_decap_8 FILLER_36_865 ();
 sg13g2_decap_8 FILLER_36_872 ();
 sg13g2_decap_8 FILLER_36_879 ();
 sg13g2_decap_8 FILLER_36_886 ();
 sg13g2_fill_2 FILLER_36_893 ();
 sg13g2_fill_2 FILLER_36_903 ();
 sg13g2_fill_1 FILLER_36_915 ();
 sg13g2_decap_8 FILLER_36_946 ();
 sg13g2_decap_8 FILLER_36_953 ();
 sg13g2_decap_4 FILLER_36_960 ();
 sg13g2_fill_1 FILLER_36_964 ();
 sg13g2_decap_4 FILLER_36_970 ();
 sg13g2_fill_1 FILLER_36_974 ();
 sg13g2_decap_8 FILLER_36_980 ();
 sg13g2_fill_2 FILLER_36_987 ();
 sg13g2_decap_8 FILLER_36_993 ();
 sg13g2_decap_4 FILLER_36_1000 ();
 sg13g2_fill_2 FILLER_36_1031 ();
 sg13g2_fill_1 FILLER_36_1033 ();
 sg13g2_decap_8 FILLER_36_1043 ();
 sg13g2_decap_4 FILLER_36_1050 ();
 sg13g2_decap_4 FILLER_36_1061 ();
 sg13g2_fill_1 FILLER_36_1065 ();
 sg13g2_decap_4 FILLER_36_1070 ();
 sg13g2_fill_1 FILLER_36_1074 ();
 sg13g2_decap_8 FILLER_36_1080 ();
 sg13g2_decap_8 FILLER_36_1087 ();
 sg13g2_decap_8 FILLER_36_1094 ();
 sg13g2_fill_2 FILLER_36_1101 ();
 sg13g2_fill_2 FILLER_36_1108 ();
 sg13g2_decap_8 FILLER_36_1149 ();
 sg13g2_decap_8 FILLER_36_1156 ();
 sg13g2_decap_8 FILLER_36_1178 ();
 sg13g2_fill_2 FILLER_36_1185 ();
 sg13g2_fill_1 FILLER_36_1187 ();
 sg13g2_decap_4 FILLER_36_1193 ();
 sg13g2_fill_2 FILLER_36_1197 ();
 sg13g2_decap_8 FILLER_36_1215 ();
 sg13g2_decap_8 FILLER_36_1222 ();
 sg13g2_decap_8 FILLER_36_1229 ();
 sg13g2_decap_8 FILLER_36_1236 ();
 sg13g2_decap_8 FILLER_36_1243 ();
 sg13g2_fill_1 FILLER_36_1283 ();
 sg13g2_decap_8 FILLER_36_1296 ();
 sg13g2_decap_8 FILLER_36_1303 ();
 sg13g2_decap_8 FILLER_36_1310 ();
 sg13g2_fill_2 FILLER_36_1317 ();
 sg13g2_decap_8 FILLER_36_1331 ();
 sg13g2_decap_8 FILLER_36_1338 ();
 sg13g2_decap_8 FILLER_36_1345 ();
 sg13g2_fill_2 FILLER_36_1352 ();
 sg13g2_fill_2 FILLER_36_1371 ();
 sg13g2_decap_8 FILLER_36_1396 ();
 sg13g2_decap_4 FILLER_36_1403 ();
 sg13g2_decap_4 FILLER_36_1415 ();
 sg13g2_fill_2 FILLER_36_1433 ();
 sg13g2_decap_4 FILLER_36_1475 ();
 sg13g2_decap_8 FILLER_36_1496 ();
 sg13g2_decap_8 FILLER_36_1503 ();
 sg13g2_fill_2 FILLER_36_1510 ();
 sg13g2_decap_8 FILLER_36_1517 ();
 sg13g2_decap_8 FILLER_36_1524 ();
 sg13g2_decap_8 FILLER_36_1531 ();
 sg13g2_decap_8 FILLER_36_1538 ();
 sg13g2_decap_8 FILLER_36_1545 ();
 sg13g2_decap_4 FILLER_36_1556 ();
 sg13g2_fill_1 FILLER_36_1560 ();
 sg13g2_decap_8 FILLER_36_1590 ();
 sg13g2_fill_2 FILLER_36_1597 ();
 sg13g2_fill_2 FILLER_36_1603 ();
 sg13g2_decap_8 FILLER_36_1608 ();
 sg13g2_fill_2 FILLER_36_1615 ();
 sg13g2_decap_8 FILLER_36_1621 ();
 sg13g2_decap_8 FILLER_36_1628 ();
 sg13g2_decap_8 FILLER_36_1635 ();
 sg13g2_decap_8 FILLER_36_1646 ();
 sg13g2_decap_8 FILLER_36_1653 ();
 sg13g2_fill_2 FILLER_36_1660 ();
 sg13g2_fill_1 FILLER_36_1662 ();
 sg13g2_fill_1 FILLER_36_1667 ();
 sg13g2_decap_4 FILLER_36_1673 ();
 sg13g2_fill_1 FILLER_36_1677 ();
 sg13g2_fill_2 FILLER_36_1704 ();
 sg13g2_decap_8 FILLER_36_1725 ();
 sg13g2_fill_2 FILLER_36_1732 ();
 sg13g2_fill_2 FILLER_36_1738 ();
 sg13g2_fill_1 FILLER_36_1740 ();
 sg13g2_fill_2 FILLER_36_1744 ();
 sg13g2_fill_2 FILLER_36_1772 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_4 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_32 ();
 sg13g2_decap_8 FILLER_37_38 ();
 sg13g2_fill_2 FILLER_37_45 ();
 sg13g2_decap_8 FILLER_37_52 ();
 sg13g2_decap_8 FILLER_37_59 ();
 sg13g2_decap_8 FILLER_37_66 ();
 sg13g2_decap_8 FILLER_37_73 ();
 sg13g2_decap_8 FILLER_37_80 ();
 sg13g2_decap_8 FILLER_37_87 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_decap_8 FILLER_37_99 ();
 sg13g2_decap_8 FILLER_37_106 ();
 sg13g2_decap_8 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_120 ();
 sg13g2_fill_1 FILLER_37_122 ();
 sg13g2_decap_8 FILLER_37_127 ();
 sg13g2_decap_4 FILLER_37_134 ();
 sg13g2_fill_2 FILLER_37_138 ();
 sg13g2_decap_8 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_160 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_fill_2 FILLER_37_190 ();
 sg13g2_fill_1 FILLER_37_192 ();
 sg13g2_decap_8 FILLER_37_198 ();
 sg13g2_decap_8 FILLER_37_205 ();
 sg13g2_decap_8 FILLER_37_212 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_fill_2 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_decap_8 FILLER_37_283 ();
 sg13g2_decap_8 FILLER_37_290 ();
 sg13g2_decap_8 FILLER_37_297 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_decap_8 FILLER_37_311 ();
 sg13g2_decap_8 FILLER_37_318 ();
 sg13g2_decap_8 FILLER_37_325 ();
 sg13g2_decap_8 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_decap_8 FILLER_37_353 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_fill_2 FILLER_37_400 ();
 sg13g2_decap_4 FILLER_37_431 ();
 sg13g2_fill_2 FILLER_37_435 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_fill_2 FILLER_37_490 ();
 sg13g2_fill_1 FILLER_37_499 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_511 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_fill_1 FILLER_37_525 ();
 sg13g2_fill_2 FILLER_37_556 ();
 sg13g2_fill_1 FILLER_37_558 ();
 sg13g2_decap_8 FILLER_37_563 ();
 sg13g2_decap_8 FILLER_37_570 ();
 sg13g2_fill_2 FILLER_37_577 ();
 sg13g2_fill_2 FILLER_37_592 ();
 sg13g2_decap_8 FILLER_37_598 ();
 sg13g2_decap_8 FILLER_37_605 ();
 sg13g2_decap_4 FILLER_37_612 ();
 sg13g2_fill_1 FILLER_37_616 ();
 sg13g2_fill_1 FILLER_37_625 ();
 sg13g2_decap_4 FILLER_37_635 ();
 sg13g2_fill_1 FILLER_37_639 ();
 sg13g2_decap_4 FILLER_37_670 ();
 sg13g2_fill_2 FILLER_37_674 ();
 sg13g2_decap_8 FILLER_37_680 ();
 sg13g2_decap_8 FILLER_37_687 ();
 sg13g2_decap_8 FILLER_37_694 ();
 sg13g2_decap_8 FILLER_37_701 ();
 sg13g2_decap_8 FILLER_37_708 ();
 sg13g2_decap_8 FILLER_37_715 ();
 sg13g2_decap_8 FILLER_37_722 ();
 sg13g2_decap_8 FILLER_37_729 ();
 sg13g2_decap_8 FILLER_37_736 ();
 sg13g2_decap_8 FILLER_37_743 ();
 sg13g2_decap_4 FILLER_37_750 ();
 sg13g2_decap_8 FILLER_37_780 ();
 sg13g2_decap_8 FILLER_37_787 ();
 sg13g2_fill_2 FILLER_37_794 ();
 sg13g2_decap_8 FILLER_37_822 ();
 sg13g2_decap_8 FILLER_37_829 ();
 sg13g2_fill_2 FILLER_37_836 ();
 sg13g2_decap_8 FILLER_37_842 ();
 sg13g2_fill_2 FILLER_37_849 ();
 sg13g2_fill_1 FILLER_37_851 ();
 sg13g2_decap_8 FILLER_37_856 ();
 sg13g2_decap_4 FILLER_37_863 ();
 sg13g2_fill_1 FILLER_37_867 ();
 sg13g2_decap_8 FILLER_37_872 ();
 sg13g2_decap_8 FILLER_37_879 ();
 sg13g2_decap_8 FILLER_37_886 ();
 sg13g2_decap_8 FILLER_37_893 ();
 sg13g2_fill_2 FILLER_37_900 ();
 sg13g2_decap_8 FILLER_37_906 ();
 sg13g2_fill_2 FILLER_37_913 ();
 sg13g2_decap_8 FILLER_37_919 ();
 sg13g2_decap_8 FILLER_37_926 ();
 sg13g2_decap_8 FILLER_37_933 ();
 sg13g2_decap_8 FILLER_37_940 ();
 sg13g2_decap_8 FILLER_37_947 ();
 sg13g2_decap_4 FILLER_37_954 ();
 sg13g2_decap_8 FILLER_37_962 ();
 sg13g2_decap_8 FILLER_37_969 ();
 sg13g2_decap_4 FILLER_37_976 ();
 sg13g2_fill_1 FILLER_37_980 ();
 sg13g2_decap_4 FILLER_37_1007 ();
 sg13g2_decap_8 FILLER_37_1015 ();
 sg13g2_fill_1 FILLER_37_1022 ();
 sg13g2_fill_1 FILLER_37_1033 ();
 sg13g2_decap_8 FILLER_37_1039 ();
 sg13g2_decap_8 FILLER_37_1046 ();
 sg13g2_decap_4 FILLER_37_1053 ();
 sg13g2_fill_2 FILLER_37_1057 ();
 sg13g2_decap_8 FILLER_37_1085 ();
 sg13g2_decap_8 FILLER_37_1092 ();
 sg13g2_decap_8 FILLER_37_1099 ();
 sg13g2_decap_8 FILLER_37_1106 ();
 sg13g2_fill_2 FILLER_37_1113 ();
 sg13g2_decap_8 FILLER_37_1119 ();
 sg13g2_decap_8 FILLER_37_1126 ();
 sg13g2_decap_8 FILLER_37_1133 ();
 sg13g2_decap_8 FILLER_37_1140 ();
 sg13g2_decap_8 FILLER_37_1147 ();
 sg13g2_decap_8 FILLER_37_1154 ();
 sg13g2_fill_1 FILLER_37_1161 ();
 sg13g2_decap_8 FILLER_37_1172 ();
 sg13g2_fill_1 FILLER_37_1179 ();
 sg13g2_decap_8 FILLER_37_1184 ();
 sg13g2_decap_8 FILLER_37_1191 ();
 sg13g2_decap_4 FILLER_37_1198 ();
 sg13g2_fill_1 FILLER_37_1202 ();
 sg13g2_decap_4 FILLER_37_1207 ();
 sg13g2_fill_1 FILLER_37_1211 ();
 sg13g2_decap_8 FILLER_37_1217 ();
 sg13g2_decap_8 FILLER_37_1224 ();
 sg13g2_decap_4 FILLER_37_1231 ();
 sg13g2_fill_2 FILLER_37_1235 ();
 sg13g2_fill_2 FILLER_37_1245 ();
 sg13g2_fill_1 FILLER_37_1251 ();
 sg13g2_fill_1 FILLER_37_1260 ();
 sg13g2_fill_1 FILLER_37_1266 ();
 sg13g2_decap_8 FILLER_37_1277 ();
 sg13g2_decap_8 FILLER_37_1284 ();
 sg13g2_decap_8 FILLER_37_1291 ();
 sg13g2_decap_8 FILLER_37_1298 ();
 sg13g2_decap_8 FILLER_37_1305 ();
 sg13g2_fill_2 FILLER_37_1312 ();
 sg13g2_decap_8 FILLER_37_1344 ();
 sg13g2_decap_4 FILLER_37_1351 ();
 sg13g2_fill_1 FILLER_37_1355 ();
 sg13g2_fill_1 FILLER_37_1365 ();
 sg13g2_fill_1 FILLER_37_1370 ();
 sg13g2_fill_2 FILLER_37_1384 ();
 sg13g2_fill_1 FILLER_37_1386 ();
 sg13g2_fill_1 FILLER_37_1391 ();
 sg13g2_decap_8 FILLER_37_1397 ();
 sg13g2_decap_8 FILLER_37_1404 ();
 sg13g2_decap_8 FILLER_37_1411 ();
 sg13g2_decap_4 FILLER_37_1418 ();
 sg13g2_decap_8 FILLER_37_1427 ();
 sg13g2_decap_8 FILLER_37_1434 ();
 sg13g2_decap_4 FILLER_37_1441 ();
 sg13g2_fill_1 FILLER_37_1445 ();
 sg13g2_decap_8 FILLER_37_1450 ();
 sg13g2_decap_8 FILLER_37_1457 ();
 sg13g2_decap_8 FILLER_37_1464 ();
 sg13g2_fill_2 FILLER_37_1471 ();
 sg13g2_decap_4 FILLER_37_1507 ();
 sg13g2_decap_8 FILLER_37_1515 ();
 sg13g2_fill_1 FILLER_37_1522 ();
 sg13g2_fill_1 FILLER_37_1527 ();
 sg13g2_decap_8 FILLER_37_1532 ();
 sg13g2_decap_8 FILLER_37_1539 ();
 sg13g2_decap_4 FILLER_37_1546 ();
 sg13g2_fill_1 FILLER_37_1550 ();
 sg13g2_decap_4 FILLER_37_1556 ();
 sg13g2_fill_2 FILLER_37_1571 ();
 sg13g2_decap_8 FILLER_37_1590 ();
 sg13g2_fill_2 FILLER_37_1597 ();
 sg13g2_fill_1 FILLER_37_1604 ();
 sg13g2_decap_8 FILLER_37_1613 ();
 sg13g2_decap_8 FILLER_37_1620 ();
 sg13g2_decap_8 FILLER_37_1627 ();
 sg13g2_decap_8 FILLER_37_1660 ();
 sg13g2_fill_2 FILLER_37_1667 ();
 sg13g2_fill_1 FILLER_37_1669 ();
 sg13g2_decap_8 FILLER_37_1674 ();
 sg13g2_decap_8 FILLER_37_1681 ();
 sg13g2_decap_8 FILLER_37_1688 ();
 sg13g2_decap_8 FILLER_37_1695 ();
 sg13g2_decap_4 FILLER_37_1702 ();
 sg13g2_decap_8 FILLER_37_1711 ();
 sg13g2_decap_8 FILLER_37_1722 ();
 sg13g2_decap_8 FILLER_37_1729 ();
 sg13g2_decap_4 FILLER_37_1736 ();
 sg13g2_decap_8 FILLER_37_1745 ();
 sg13g2_fill_1 FILLER_37_1752 ();
 sg13g2_decap_8 FILLER_37_1757 ();
 sg13g2_decap_8 FILLER_37_1764 ();
 sg13g2_fill_2 FILLER_37_1771 ();
 sg13g2_fill_1 FILLER_37_1773 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_fill_2 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_55 ();
 sg13g2_decap_8 FILLER_38_62 ();
 sg13g2_decap_8 FILLER_38_69 ();
 sg13g2_decap_8 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_83 ();
 sg13g2_fill_2 FILLER_38_87 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_8 FILLER_38_100 ();
 sg13g2_decap_8 FILLER_38_107 ();
 sg13g2_decap_8 FILLER_38_114 ();
 sg13g2_fill_2 FILLER_38_121 ();
 sg13g2_fill_1 FILLER_38_123 ();
 sg13g2_decap_8 FILLER_38_129 ();
 sg13g2_decap_8 FILLER_38_136 ();
 sg13g2_fill_2 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_153 ();
 sg13g2_decap_4 FILLER_38_163 ();
 sg13g2_fill_1 FILLER_38_167 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_decap_4 FILLER_38_249 ();
 sg13g2_fill_2 FILLER_38_261 ();
 sg13g2_decap_8 FILLER_38_283 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_decap_8 FILLER_38_297 ();
 sg13g2_decap_8 FILLER_38_304 ();
 sg13g2_decap_8 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_318 ();
 sg13g2_decap_8 FILLER_38_325 ();
 sg13g2_decap_8 FILLER_38_332 ();
 sg13g2_decap_8 FILLER_38_339 ();
 sg13g2_decap_8 FILLER_38_346 ();
 sg13g2_decap_8 FILLER_38_353 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_fill_1 FILLER_38_375 ();
 sg13g2_decap_4 FILLER_38_379 ();
 sg13g2_decap_4 FILLER_38_388 ();
 sg13g2_fill_2 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_38_456 ();
 sg13g2_fill_1 FILLER_38_463 ();
 sg13g2_fill_2 FILLER_38_493 ();
 sg13g2_decap_8 FILLER_38_524 ();
 sg13g2_decap_4 FILLER_38_531 ();
 sg13g2_decap_8 FILLER_38_539 ();
 sg13g2_decap_8 FILLER_38_546 ();
 sg13g2_decap_8 FILLER_38_579 ();
 sg13g2_fill_1 FILLER_38_586 ();
 sg13g2_decap_8 FILLER_38_638 ();
 sg13g2_decap_8 FILLER_38_649 ();
 sg13g2_decap_8 FILLER_38_656 ();
 sg13g2_decap_8 FILLER_38_663 ();
 sg13g2_decap_8 FILLER_38_670 ();
 sg13g2_fill_2 FILLER_38_677 ();
 sg13g2_decap_8 FILLER_38_694 ();
 sg13g2_decap_8 FILLER_38_701 ();
 sg13g2_decap_4 FILLER_38_708 ();
 sg13g2_decap_8 FILLER_38_716 ();
 sg13g2_decap_8 FILLER_38_723 ();
 sg13g2_decap_8 FILLER_38_730 ();
 sg13g2_decap_8 FILLER_38_737 ();
 sg13g2_fill_2 FILLER_38_744 ();
 sg13g2_fill_2 FILLER_38_758 ();
 sg13g2_decap_8 FILLER_38_767 ();
 sg13g2_decap_8 FILLER_38_774 ();
 sg13g2_decap_8 FILLER_38_781 ();
 sg13g2_decap_8 FILLER_38_788 ();
 sg13g2_decap_4 FILLER_38_795 ();
 sg13g2_fill_1 FILLER_38_799 ();
 sg13g2_decap_8 FILLER_38_804 ();
 sg13g2_decap_8 FILLER_38_811 ();
 sg13g2_decap_8 FILLER_38_818 ();
 sg13g2_decap_8 FILLER_38_825 ();
 sg13g2_decap_8 FILLER_38_832 ();
 sg13g2_fill_1 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_871 ();
 sg13g2_fill_2 FILLER_38_878 ();
 sg13g2_decap_8 FILLER_38_911 ();
 sg13g2_fill_1 FILLER_38_918 ();
 sg13g2_decap_8 FILLER_38_923 ();
 sg13g2_decap_8 FILLER_38_930 ();
 sg13g2_decap_8 FILLER_38_937 ();
 sg13g2_decap_8 FILLER_38_944 ();
 sg13g2_decap_8 FILLER_38_977 ();
 sg13g2_decap_8 FILLER_38_984 ();
 sg13g2_decap_8 FILLER_38_991 ();
 sg13g2_decap_8 FILLER_38_998 ();
 sg13g2_decap_8 FILLER_38_1009 ();
 sg13g2_decap_8 FILLER_38_1016 ();
 sg13g2_decap_8 FILLER_38_1023 ();
 sg13g2_decap_8 FILLER_38_1030 ();
 sg13g2_decap_8 FILLER_38_1037 ();
 sg13g2_decap_8 FILLER_38_1044 ();
 sg13g2_decap_8 FILLER_38_1051 ();
 sg13g2_decap_8 FILLER_38_1058 ();
 sg13g2_fill_2 FILLER_38_1065 ();
 sg13g2_fill_1 FILLER_38_1067 ();
 sg13g2_decap_8 FILLER_38_1076 ();
 sg13g2_decap_8 FILLER_38_1083 ();
 sg13g2_decap_4 FILLER_38_1090 ();
 sg13g2_fill_2 FILLER_38_1094 ();
 sg13g2_decap_8 FILLER_38_1100 ();
 sg13g2_fill_1 FILLER_38_1107 ();
 sg13g2_decap_8 FILLER_38_1116 ();
 sg13g2_decap_8 FILLER_38_1123 ();
 sg13g2_decap_8 FILLER_38_1130 ();
 sg13g2_decap_8 FILLER_38_1137 ();
 sg13g2_decap_8 FILLER_38_1144 ();
 sg13g2_decap_8 FILLER_38_1151 ();
 sg13g2_decap_4 FILLER_38_1158 ();
 sg13g2_fill_1 FILLER_38_1162 ();
 sg13g2_decap_8 FILLER_38_1189 ();
 sg13g2_decap_8 FILLER_38_1196 ();
 sg13g2_decap_8 FILLER_38_1207 ();
 sg13g2_fill_2 FILLER_38_1214 ();
 sg13g2_fill_1 FILLER_38_1216 ();
 sg13g2_decap_8 FILLER_38_1221 ();
 sg13g2_fill_2 FILLER_38_1228 ();
 sg13g2_fill_1 FILLER_38_1230 ();
 sg13g2_decap_8 FILLER_38_1241 ();
 sg13g2_decap_8 FILLER_38_1248 ();
 sg13g2_fill_2 FILLER_38_1255 ();
 sg13g2_decap_8 FILLER_38_1279 ();
 sg13g2_decap_8 FILLER_38_1286 ();
 sg13g2_decap_8 FILLER_38_1293 ();
 sg13g2_decap_8 FILLER_38_1300 ();
 sg13g2_decap_8 FILLER_38_1307 ();
 sg13g2_decap_8 FILLER_38_1314 ();
 sg13g2_decap_8 FILLER_38_1325 ();
 sg13g2_decap_8 FILLER_38_1332 ();
 sg13g2_decap_8 FILLER_38_1339 ();
 sg13g2_decap_8 FILLER_38_1346 ();
 sg13g2_fill_2 FILLER_38_1353 ();
 sg13g2_fill_1 FILLER_38_1355 ();
 sg13g2_decap_8 FILLER_38_1360 ();
 sg13g2_decap_8 FILLER_38_1367 ();
 sg13g2_decap_8 FILLER_38_1374 ();
 sg13g2_decap_4 FILLER_38_1381 ();
 sg13g2_decap_8 FILLER_38_1389 ();
 sg13g2_decap_8 FILLER_38_1396 ();
 sg13g2_decap_8 FILLER_38_1403 ();
 sg13g2_decap_8 FILLER_38_1410 ();
 sg13g2_decap_8 FILLER_38_1417 ();
 sg13g2_decap_4 FILLER_38_1424 ();
 sg13g2_decap_8 FILLER_38_1432 ();
 sg13g2_decap_4 FILLER_38_1439 ();
 sg13g2_fill_2 FILLER_38_1443 ();
 sg13g2_decap_8 FILLER_38_1449 ();
 sg13g2_decap_8 FILLER_38_1456 ();
 sg13g2_decap_8 FILLER_38_1463 ();
 sg13g2_decap_8 FILLER_38_1470 ();
 sg13g2_decap_8 FILLER_38_1477 ();
 sg13g2_decap_8 FILLER_38_1484 ();
 sg13g2_decap_8 FILLER_38_1491 ();
 sg13g2_decap_4 FILLER_38_1498 ();
 sg13g2_fill_2 FILLER_38_1502 ();
 sg13g2_decap_8 FILLER_38_1530 ();
 sg13g2_decap_8 FILLER_38_1537 ();
 sg13g2_fill_2 FILLER_38_1544 ();
 sg13g2_fill_1 FILLER_38_1566 ();
 sg13g2_fill_2 FILLER_38_1597 ();
 sg13g2_fill_1 FILLER_38_1599 ();
 sg13g2_decap_8 FILLER_38_1629 ();
 sg13g2_decap_8 FILLER_38_1636 ();
 sg13g2_decap_8 FILLER_38_1643 ();
 sg13g2_fill_2 FILLER_38_1650 ();
 sg13g2_fill_1 FILLER_38_1652 ();
 sg13g2_decap_8 FILLER_38_1656 ();
 sg13g2_decap_8 FILLER_38_1663 ();
 sg13g2_decap_8 FILLER_38_1670 ();
 sg13g2_decap_8 FILLER_38_1677 ();
 sg13g2_decap_8 FILLER_38_1684 ();
 sg13g2_decap_8 FILLER_38_1691 ();
 sg13g2_decap_4 FILLER_38_1698 ();
 sg13g2_fill_1 FILLER_38_1702 ();
 sg13g2_fill_2 FILLER_38_1737 ();
 sg13g2_decap_8 FILLER_38_1758 ();
 sg13g2_decap_8 FILLER_38_1765 ();
 sg13g2_fill_2 FILLER_38_1772 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_4 FILLER_39_28 ();
 sg13g2_fill_2 FILLER_39_32 ();
 sg13g2_fill_2 FILLER_39_38 ();
 sg13g2_decap_8 FILLER_39_48 ();
 sg13g2_decap_4 FILLER_39_55 ();
 sg13g2_fill_1 FILLER_39_59 ();
 sg13g2_decap_8 FILLER_39_68 ();
 sg13g2_decap_8 FILLER_39_75 ();
 sg13g2_decap_4 FILLER_39_82 ();
 sg13g2_decap_4 FILLER_39_95 ();
 sg13g2_fill_1 FILLER_39_114 ();
 sg13g2_fill_2 FILLER_39_119 ();
 sg13g2_fill_1 FILLER_39_121 ();
 sg13g2_fill_2 FILLER_39_129 ();
 sg13g2_fill_1 FILLER_39_131 ();
 sg13g2_fill_1 FILLER_39_148 ();
 sg13g2_decap_4 FILLER_39_153 ();
 sg13g2_fill_2 FILLER_39_157 ();
 sg13g2_decap_8 FILLER_39_172 ();
 sg13g2_decap_8 FILLER_39_179 ();
 sg13g2_decap_4 FILLER_39_186 ();
 sg13g2_fill_2 FILLER_39_199 ();
 sg13g2_fill_2 FILLER_39_205 ();
 sg13g2_decap_4 FILLER_39_211 ();
 sg13g2_decap_8 FILLER_39_233 ();
 sg13g2_decap_8 FILLER_39_240 ();
 sg13g2_decap_8 FILLER_39_247 ();
 sg13g2_fill_2 FILLER_39_254 ();
 sg13g2_fill_2 FILLER_39_261 ();
 sg13g2_fill_2 FILLER_39_268 ();
 sg13g2_decap_8 FILLER_39_275 ();
 sg13g2_decap_8 FILLER_39_282 ();
 sg13g2_decap_8 FILLER_39_289 ();
 sg13g2_decap_8 FILLER_39_296 ();
 sg13g2_fill_2 FILLER_39_303 ();
 sg13g2_fill_1 FILLER_39_305 ();
 sg13g2_decap_8 FILLER_39_311 ();
 sg13g2_decap_8 FILLER_39_318 ();
 sg13g2_decap_4 FILLER_39_325 ();
 sg13g2_decap_4 FILLER_39_342 ();
 sg13g2_fill_2 FILLER_39_346 ();
 sg13g2_decap_4 FILLER_39_361 ();
 sg13g2_fill_1 FILLER_39_365 ();
 sg13g2_fill_2 FILLER_39_370 ();
 sg13g2_decap_8 FILLER_39_377 ();
 sg13g2_fill_2 FILLER_39_384 ();
 sg13g2_fill_1 FILLER_39_386 ();
 sg13g2_decap_4 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_39_409 ();
 sg13g2_decap_8 FILLER_39_416 ();
 sg13g2_decap_8 FILLER_39_423 ();
 sg13g2_decap_8 FILLER_39_430 ();
 sg13g2_decap_8 FILLER_39_437 ();
 sg13g2_decap_8 FILLER_39_444 ();
 sg13g2_fill_2 FILLER_39_451 ();
 sg13g2_decap_8 FILLER_39_456 ();
 sg13g2_decap_8 FILLER_39_463 ();
 sg13g2_fill_1 FILLER_39_470 ();
 sg13g2_fill_2 FILLER_39_475 ();
 sg13g2_decap_4 FILLER_39_483 ();
 sg13g2_fill_2 FILLER_39_487 ();
 sg13g2_decap_8 FILLER_39_495 ();
 sg13g2_decap_4 FILLER_39_502 ();
 sg13g2_decap_8 FILLER_39_509 ();
 sg13g2_fill_1 FILLER_39_516 ();
 sg13g2_decap_8 FILLER_39_521 ();
 sg13g2_decap_4 FILLER_39_528 ();
 sg13g2_fill_2 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_538 ();
 sg13g2_decap_8 FILLER_39_545 ();
 sg13g2_decap_8 FILLER_39_552 ();
 sg13g2_decap_8 FILLER_39_559 ();
 sg13g2_decap_8 FILLER_39_566 ();
 sg13g2_decap_8 FILLER_39_573 ();
 sg13g2_decap_8 FILLER_39_580 ();
 sg13g2_decap_8 FILLER_39_587 ();
 sg13g2_decap_4 FILLER_39_594 ();
 sg13g2_fill_2 FILLER_39_598 ();
 sg13g2_decap_8 FILLER_39_604 ();
 sg13g2_decap_4 FILLER_39_611 ();
 sg13g2_decap_8 FILLER_39_619 ();
 sg13g2_decap_8 FILLER_39_626 ();
 sg13g2_decap_8 FILLER_39_633 ();
 sg13g2_decap_8 FILLER_39_640 ();
 sg13g2_decap_8 FILLER_39_647 ();
 sg13g2_decap_8 FILLER_39_654 ();
 sg13g2_decap_4 FILLER_39_661 ();
 sg13g2_fill_1 FILLER_39_665 ();
 sg13g2_fill_2 FILLER_39_691 ();
 sg13g2_decap_8 FILLER_39_731 ();
 sg13g2_decap_8 FILLER_39_738 ();
 sg13g2_fill_2 FILLER_39_745 ();
 sg13g2_fill_1 FILLER_39_759 ();
 sg13g2_fill_2 FILLER_39_765 ();
 sg13g2_decap_8 FILLER_39_801 ();
 sg13g2_decap_8 FILLER_39_808 ();
 sg13g2_decap_4 FILLER_39_815 ();
 sg13g2_decap_8 FILLER_39_823 ();
 sg13g2_decap_8 FILLER_39_830 ();
 sg13g2_decap_8 FILLER_39_837 ();
 sg13g2_decap_8 FILLER_39_844 ();
 sg13g2_decap_8 FILLER_39_851 ();
 sg13g2_decap_8 FILLER_39_858 ();
 sg13g2_decap_8 FILLER_39_865 ();
 sg13g2_fill_2 FILLER_39_872 ();
 sg13g2_fill_1 FILLER_39_874 ();
 sg13g2_decap_8 FILLER_39_894 ();
 sg13g2_decap_8 FILLER_39_901 ();
 sg13g2_fill_2 FILLER_39_908 ();
 sg13g2_fill_1 FILLER_39_910 ();
 sg13g2_decap_8 FILLER_39_915 ();
 sg13g2_decap_8 FILLER_39_922 ();
 sg13g2_decap_8 FILLER_39_929 ();
 sg13g2_decap_8 FILLER_39_936 ();
 sg13g2_decap_8 FILLER_39_943 ();
 sg13g2_decap_8 FILLER_39_950 ();
 sg13g2_decap_8 FILLER_39_957 ();
 sg13g2_decap_8 FILLER_39_964 ();
 sg13g2_decap_8 FILLER_39_971 ();
 sg13g2_decap_8 FILLER_39_978 ();
 sg13g2_decap_8 FILLER_39_985 ();
 sg13g2_fill_1 FILLER_39_992 ();
 sg13g2_decap_8 FILLER_39_1017 ();
 sg13g2_decap_8 FILLER_39_1024 ();
 sg13g2_decap_8 FILLER_39_1031 ();
 sg13g2_fill_2 FILLER_39_1038 ();
 sg13g2_fill_1 FILLER_39_1040 ();
 sg13g2_decap_8 FILLER_39_1050 ();
 sg13g2_decap_8 FILLER_39_1057 ();
 sg13g2_fill_1 FILLER_39_1064 ();
 sg13g2_decap_8 FILLER_39_1091 ();
 sg13g2_decap_8 FILLER_39_1128 ();
 sg13g2_decap_8 FILLER_39_1135 ();
 sg13g2_fill_2 FILLER_39_1142 ();
 sg13g2_fill_1 FILLER_39_1144 ();
 sg13g2_decap_4 FILLER_39_1150 ();
 sg13g2_fill_1 FILLER_39_1154 ();
 sg13g2_decap_8 FILLER_39_1159 ();
 sg13g2_fill_2 FILLER_39_1166 ();
 sg13g2_decap_4 FILLER_39_1176 ();
 sg13g2_decap_8 FILLER_39_1185 ();
 sg13g2_decap_4 FILLER_39_1192 ();
 sg13g2_fill_2 FILLER_39_1196 ();
 sg13g2_decap_8 FILLER_39_1207 ();
 sg13g2_fill_1 FILLER_39_1214 ();
 sg13g2_decap_4 FILLER_39_1226 ();
 sg13g2_fill_2 FILLER_39_1230 ();
 sg13g2_fill_2 FILLER_39_1258 ();
 sg13g2_fill_1 FILLER_39_1263 ();
 sg13g2_fill_1 FILLER_39_1270 ();
 sg13g2_fill_1 FILLER_39_1278 ();
 sg13g2_decap_4 FILLER_39_1283 ();
 sg13g2_fill_2 FILLER_39_1287 ();
 sg13g2_fill_1 FILLER_39_1318 ();
 sg13g2_decap_8 FILLER_39_1323 ();
 sg13g2_decap_8 FILLER_39_1330 ();
 sg13g2_decap_8 FILLER_39_1337 ();
 sg13g2_decap_8 FILLER_39_1344 ();
 sg13g2_decap_8 FILLER_39_1351 ();
 sg13g2_decap_8 FILLER_39_1358 ();
 sg13g2_decap_8 FILLER_39_1365 ();
 sg13g2_decap_8 FILLER_39_1372 ();
 sg13g2_fill_1 FILLER_39_1379 ();
 sg13g2_decap_8 FILLER_39_1383 ();
 sg13g2_fill_2 FILLER_39_1390 ();
 sg13g2_fill_1 FILLER_39_1392 ();
 sg13g2_decap_4 FILLER_39_1397 ();
 sg13g2_fill_2 FILLER_39_1401 ();
 sg13g2_fill_1 FILLER_39_1407 ();
 sg13g2_fill_1 FILLER_39_1434 ();
 sg13g2_fill_1 FILLER_39_1464 ();
 sg13g2_fill_1 FILLER_39_1468 ();
 sg13g2_decap_8 FILLER_39_1504 ();
 sg13g2_decap_8 FILLER_39_1511 ();
 sg13g2_decap_8 FILLER_39_1518 ();
 sg13g2_decap_8 FILLER_39_1525 ();
 sg13g2_decap_8 FILLER_39_1532 ();
 sg13g2_decap_8 FILLER_39_1539 ();
 sg13g2_decap_8 FILLER_39_1546 ();
 sg13g2_decap_8 FILLER_39_1553 ();
 sg13g2_decap_4 FILLER_39_1560 ();
 sg13g2_decap_8 FILLER_39_1569 ();
 sg13g2_decap_8 FILLER_39_1576 ();
 sg13g2_decap_8 FILLER_39_1583 ();
 sg13g2_decap_8 FILLER_39_1590 ();
 sg13g2_fill_1 FILLER_39_1597 ();
 sg13g2_decap_8 FILLER_39_1604 ();
 sg13g2_decap_8 FILLER_39_1611 ();
 sg13g2_decap_8 FILLER_39_1618 ();
 sg13g2_decap_4 FILLER_39_1625 ();
 sg13g2_fill_2 FILLER_39_1635 ();
 sg13g2_decap_8 FILLER_39_1640 ();
 sg13g2_decap_8 FILLER_39_1647 ();
 sg13g2_decap_8 FILLER_39_1654 ();
 sg13g2_decap_8 FILLER_39_1661 ();
 sg13g2_decap_8 FILLER_39_1668 ();
 sg13g2_decap_8 FILLER_39_1675 ();
 sg13g2_decap_8 FILLER_39_1682 ();
 sg13g2_fill_1 FILLER_39_1689 ();
 sg13g2_decap_8 FILLER_39_1711 ();
 sg13g2_decap_8 FILLER_39_1718 ();
 sg13g2_decap_8 FILLER_39_1725 ();
 sg13g2_decap_8 FILLER_39_1732 ();
 sg13g2_decap_4 FILLER_39_1770 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_fill_1 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_43 ();
 sg13g2_fill_2 FILLER_40_50 ();
 sg13g2_decap_4 FILLER_40_60 ();
 sg13g2_fill_2 FILLER_40_68 ();
 sg13g2_fill_1 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_75 ();
 sg13g2_decap_4 FILLER_40_82 ();
 sg13g2_fill_1 FILLER_40_86 ();
 sg13g2_decap_4 FILLER_40_100 ();
 sg13g2_fill_1 FILLER_40_108 ();
 sg13g2_decap_4 FILLER_40_118 ();
 sg13g2_fill_2 FILLER_40_122 ();
 sg13g2_decap_8 FILLER_40_137 ();
 sg13g2_decap_8 FILLER_40_144 ();
 sg13g2_decap_8 FILLER_40_151 ();
 sg13g2_decap_8 FILLER_40_158 ();
 sg13g2_decap_8 FILLER_40_165 ();
 sg13g2_decap_8 FILLER_40_172 ();
 sg13g2_fill_1 FILLER_40_188 ();
 sg13g2_fill_2 FILLER_40_199 ();
 sg13g2_fill_2 FILLER_40_206 ();
 sg13g2_fill_1 FILLER_40_208 ();
 sg13g2_fill_1 FILLER_40_213 ();
 sg13g2_decap_4 FILLER_40_219 ();
 sg13g2_fill_2 FILLER_40_223 ();
 sg13g2_decap_8 FILLER_40_229 ();
 sg13g2_decap_8 FILLER_40_236 ();
 sg13g2_decap_8 FILLER_40_243 ();
 sg13g2_decap_4 FILLER_40_250 ();
 sg13g2_fill_1 FILLER_40_254 ();
 sg13g2_decap_4 FILLER_40_260 ();
 sg13g2_decap_4 FILLER_40_284 ();
 sg13g2_fill_1 FILLER_40_288 ();
 sg13g2_decap_8 FILLER_40_293 ();
 sg13g2_decap_4 FILLER_40_300 ();
 sg13g2_fill_1 FILLER_40_304 ();
 sg13g2_decap_4 FILLER_40_325 ();
 sg13g2_fill_2 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_337 ();
 sg13g2_fill_2 FILLER_40_344 ();
 sg13g2_fill_1 FILLER_40_346 ();
 sg13g2_fill_2 FILLER_40_361 ();
 sg13g2_fill_1 FILLER_40_363 ();
 sg13g2_decap_8 FILLER_40_368 ();
 sg13g2_decap_4 FILLER_40_391 ();
 sg13g2_fill_2 FILLER_40_395 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_decap_8 FILLER_40_409 ();
 sg13g2_decap_8 FILLER_40_416 ();
 sg13g2_decap_4 FILLER_40_423 ();
 sg13g2_fill_1 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_fill_2 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_454 ();
 sg13g2_decap_8 FILLER_40_461 ();
 sg13g2_decap_8 FILLER_40_468 ();
 sg13g2_decap_8 FILLER_40_475 ();
 sg13g2_decap_8 FILLER_40_482 ();
 sg13g2_decap_8 FILLER_40_489 ();
 sg13g2_decap_8 FILLER_40_500 ();
 sg13g2_decap_8 FILLER_40_507 ();
 sg13g2_decap_8 FILLER_40_514 ();
 sg13g2_decap_4 FILLER_40_521 ();
 sg13g2_fill_2 FILLER_40_525 ();
 sg13g2_decap_8 FILLER_40_557 ();
 sg13g2_decap_8 FILLER_40_564 ();
 sg13g2_fill_2 FILLER_40_571 ();
 sg13g2_decap_8 FILLER_40_602 ();
 sg13g2_decap_8 FILLER_40_609 ();
 sg13g2_decap_4 FILLER_40_620 ();
 sg13g2_fill_2 FILLER_40_624 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_8 FILLER_40_644 ();
 sg13g2_decap_8 FILLER_40_651 ();
 sg13g2_fill_2 FILLER_40_658 ();
 sg13g2_fill_1 FILLER_40_660 ();
 sg13g2_decap_8 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_679 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_decap_8 FILLER_40_693 ();
 sg13g2_decap_8 FILLER_40_700 ();
 sg13g2_fill_2 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_714 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_728 ();
 sg13g2_decap_4 FILLER_40_735 ();
 sg13g2_fill_1 FILLER_40_739 ();
 sg13g2_fill_2 FILLER_40_748 ();
 sg13g2_fill_1 FILLER_40_750 ();
 sg13g2_decap_8 FILLER_40_755 ();
 sg13g2_decap_8 FILLER_40_762 ();
 sg13g2_fill_2 FILLER_40_777 ();
 sg13g2_fill_1 FILLER_40_779 ();
 sg13g2_fill_2 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_790 ();
 sg13g2_decap_8 FILLER_40_797 ();
 sg13g2_decap_8 FILLER_40_804 ();
 sg13g2_decap_8 FILLER_40_841 ();
 sg13g2_decap_8 FILLER_40_848 ();
 sg13g2_decap_8 FILLER_40_855 ();
 sg13g2_decap_8 FILLER_40_862 ();
 sg13g2_fill_1 FILLER_40_869 ();
 sg13g2_decap_4 FILLER_40_878 ();
 sg13g2_fill_2 FILLER_40_882 ();
 sg13g2_decap_8 FILLER_40_892 ();
 sg13g2_decap_4 FILLER_40_899 ();
 sg13g2_fill_1 FILLER_40_903 ();
 sg13g2_fill_2 FILLER_40_934 ();
 sg13g2_fill_1 FILLER_40_936 ();
 sg13g2_decap_8 FILLER_40_946 ();
 sg13g2_decap_8 FILLER_40_953 ();
 sg13g2_decap_8 FILLER_40_960 ();
 sg13g2_decap_8 FILLER_40_967 ();
 sg13g2_decap_8 FILLER_40_974 ();
 sg13g2_decap_8 FILLER_40_981 ();
 sg13g2_decap_4 FILLER_40_988 ();
 sg13g2_fill_1 FILLER_40_992 ();
 sg13g2_fill_2 FILLER_40_997 ();
 sg13g2_decap_8 FILLER_40_1027 ();
 sg13g2_decap_8 FILLER_40_1034 ();
 sg13g2_fill_2 FILLER_40_1046 ();
 sg13g2_fill_1 FILLER_40_1048 ();
 sg13g2_decap_4 FILLER_40_1054 ();
 sg13g2_decap_8 FILLER_40_1065 ();
 sg13g2_decap_8 FILLER_40_1072 ();
 sg13g2_decap_4 FILLER_40_1079 ();
 sg13g2_fill_1 FILLER_40_1083 ();
 sg13g2_decap_8 FILLER_40_1088 ();
 sg13g2_decap_8 FILLER_40_1095 ();
 sg13g2_decap_4 FILLER_40_1102 ();
 sg13g2_fill_2 FILLER_40_1106 ();
 sg13g2_decap_8 FILLER_40_1113 ();
 sg13g2_decap_8 FILLER_40_1120 ();
 sg13g2_fill_2 FILLER_40_1127 ();
 sg13g2_fill_1 FILLER_40_1129 ();
 sg13g2_decap_8 FILLER_40_1134 ();
 sg13g2_decap_8 FILLER_40_1141 ();
 sg13g2_decap_8 FILLER_40_1148 ();
 sg13g2_decap_8 FILLER_40_1155 ();
 sg13g2_decap_8 FILLER_40_1166 ();
 sg13g2_decap_8 FILLER_40_1173 ();
 sg13g2_decap_8 FILLER_40_1180 ();
 sg13g2_fill_2 FILLER_40_1187 ();
 sg13g2_fill_1 FILLER_40_1189 ();
 sg13g2_decap_8 FILLER_40_1195 ();
 sg13g2_decap_8 FILLER_40_1202 ();
 sg13g2_decap_8 FILLER_40_1209 ();
 sg13g2_decap_4 FILLER_40_1216 ();
 sg13g2_decap_4 FILLER_40_1224 ();
 sg13g2_fill_2 FILLER_40_1228 ();
 sg13g2_decap_4 FILLER_40_1234 ();
 sg13g2_decap_4 FILLER_40_1251 ();
 sg13g2_decap_8 FILLER_40_1259 ();
 sg13g2_decap_8 FILLER_40_1266 ();
 sg13g2_decap_8 FILLER_40_1273 ();
 sg13g2_decap_8 FILLER_40_1280 ();
 sg13g2_fill_2 FILLER_40_1287 ();
 sg13g2_fill_1 FILLER_40_1289 ();
 sg13g2_decap_8 FILLER_40_1299 ();
 sg13g2_fill_2 FILLER_40_1306 ();
 sg13g2_fill_1 FILLER_40_1308 ();
 sg13g2_fill_2 FILLER_40_1314 ();
 sg13g2_fill_1 FILLER_40_1316 ();
 sg13g2_decap_8 FILLER_40_1332 ();
 sg13g2_decap_8 FILLER_40_1339 ();
 sg13g2_decap_4 FILLER_40_1346 ();
 sg13g2_fill_2 FILLER_40_1357 ();
 sg13g2_fill_2 FILLER_40_1367 ();
 sg13g2_decap_4 FILLER_40_1372 ();
 sg13g2_fill_1 FILLER_40_1376 ();
 sg13g2_fill_1 FILLER_40_1384 ();
 sg13g2_fill_2 FILLER_40_1395 ();
 sg13g2_decap_4 FILLER_40_1401 ();
 sg13g2_fill_2 FILLER_40_1405 ();
 sg13g2_fill_1 FILLER_40_1415 ();
 sg13g2_decap_8 FILLER_40_1424 ();
 sg13g2_fill_2 FILLER_40_1431 ();
 sg13g2_decap_8 FILLER_40_1446 ();
 sg13g2_decap_8 FILLER_40_1453 ();
 sg13g2_decap_8 FILLER_40_1460 ();
 sg13g2_decap_8 FILLER_40_1467 ();
 sg13g2_decap_8 FILLER_40_1474 ();
 sg13g2_decap_4 FILLER_40_1481 ();
 sg13g2_decap_8 FILLER_40_1489 ();
 sg13g2_decap_4 FILLER_40_1496 ();
 sg13g2_fill_2 FILLER_40_1500 ();
 sg13g2_decap_8 FILLER_40_1508 ();
 sg13g2_decap_8 FILLER_40_1515 ();
 sg13g2_decap_8 FILLER_40_1522 ();
 sg13g2_decap_8 FILLER_40_1529 ();
 sg13g2_decap_4 FILLER_40_1536 ();
 sg13g2_fill_2 FILLER_40_1540 ();
 sg13g2_decap_8 FILLER_40_1552 ();
 sg13g2_decap_8 FILLER_40_1559 ();
 sg13g2_fill_2 FILLER_40_1595 ();
 sg13g2_fill_1 FILLER_40_1597 ();
 sg13g2_decap_8 FILLER_40_1602 ();
 sg13g2_decap_8 FILLER_40_1609 ();
 sg13g2_decap_8 FILLER_40_1616 ();
 sg13g2_decap_4 FILLER_40_1623 ();
 sg13g2_fill_2 FILLER_40_1627 ();
 sg13g2_fill_1 FILLER_40_1635 ();
 sg13g2_fill_1 FILLER_40_1662 ();
 sg13g2_fill_1 FILLER_40_1689 ();
 sg13g2_fill_1 FILLER_40_1703 ();
 sg13g2_decap_8 FILLER_40_1712 ();
 sg13g2_decap_8 FILLER_40_1719 ();
 sg13g2_decap_8 FILLER_40_1726 ();
 sg13g2_fill_1 FILLER_40_1753 ();
 sg13g2_decap_8 FILLER_40_1761 ();
 sg13g2_decap_4 FILLER_40_1768 ();
 sg13g2_fill_2 FILLER_40_1772 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_4 FILLER_41_26 ();
 sg13g2_decap_4 FILLER_41_46 ();
 sg13g2_fill_1 FILLER_41_54 ();
 sg13g2_fill_1 FILLER_41_68 ();
 sg13g2_decap_8 FILLER_41_73 ();
 sg13g2_fill_2 FILLER_41_80 ();
 sg13g2_fill_1 FILLER_41_82 ();
 sg13g2_fill_1 FILLER_41_92 ();
 sg13g2_decap_4 FILLER_41_102 ();
 sg13g2_decap_8 FILLER_41_118 ();
 sg13g2_decap_8 FILLER_41_125 ();
 sg13g2_fill_2 FILLER_41_132 ();
 sg13g2_fill_2 FILLER_41_143 ();
 sg13g2_fill_1 FILLER_41_155 ();
 sg13g2_decap_8 FILLER_41_160 ();
 sg13g2_decap_4 FILLER_41_167 ();
 sg13g2_fill_2 FILLER_41_185 ();
 sg13g2_fill_1 FILLER_41_191 ();
 sg13g2_fill_1 FILLER_41_198 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_fill_2 FILLER_41_214 ();
 sg13g2_decap_4 FILLER_41_220 ();
 sg13g2_decap_8 FILLER_41_234 ();
 sg13g2_decap_8 FILLER_41_241 ();
 sg13g2_fill_2 FILLER_41_248 ();
 sg13g2_decap_8 FILLER_41_254 ();
 sg13g2_decap_8 FILLER_41_261 ();
 sg13g2_fill_1 FILLER_41_268 ();
 sg13g2_fill_1 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_295 ();
 sg13g2_fill_2 FILLER_41_302 ();
 sg13g2_decap_8 FILLER_41_310 ();
 sg13g2_decap_8 FILLER_41_317 ();
 sg13g2_decap_8 FILLER_41_324 ();
 sg13g2_fill_2 FILLER_41_331 ();
 sg13g2_decap_8 FILLER_41_340 ();
 sg13g2_decap_8 FILLER_41_365 ();
 sg13g2_fill_1 FILLER_41_372 ();
 sg13g2_fill_2 FILLER_41_382 ();
 sg13g2_fill_1 FILLER_41_384 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_fill_2 FILLER_41_404 ();
 sg13g2_decap_8 FILLER_41_416 ();
 sg13g2_decap_8 FILLER_41_423 ();
 sg13g2_decap_8 FILLER_41_430 ();
 sg13g2_fill_2 FILLER_41_437 ();
 sg13g2_decap_8 FILLER_41_470 ();
 sg13g2_decap_8 FILLER_41_477 ();
 sg13g2_fill_1 FILLER_41_484 ();
 sg13g2_fill_2 FILLER_41_520 ();
 sg13g2_decap_8 FILLER_41_532 ();
 sg13g2_fill_2 FILLER_41_539 ();
 sg13g2_decap_4 FILLER_41_545 ();
 sg13g2_fill_1 FILLER_41_549 ();
 sg13g2_fill_1 FILLER_41_555 ();
 sg13g2_decap_8 FILLER_41_560 ();
 sg13g2_decap_4 FILLER_41_567 ();
 sg13g2_decap_8 FILLER_41_576 ();
 sg13g2_decap_8 FILLER_41_591 ();
 sg13g2_decap_8 FILLER_41_598 ();
 sg13g2_fill_2 FILLER_41_605 ();
 sg13g2_decap_4 FILLER_41_612 ();
 sg13g2_fill_2 FILLER_41_616 ();
 sg13g2_decap_8 FILLER_41_652 ();
 sg13g2_decap_4 FILLER_41_659 ();
 sg13g2_fill_2 FILLER_41_663 ();
 sg13g2_decap_8 FILLER_41_679 ();
 sg13g2_fill_1 FILLER_41_691 ();
 sg13g2_fill_1 FILLER_41_697 ();
 sg13g2_decap_4 FILLER_41_737 ();
 sg13g2_fill_1 FILLER_41_741 ();
 sg13g2_fill_2 FILLER_41_750 ();
 sg13g2_fill_1 FILLER_41_752 ();
 sg13g2_decap_4 FILLER_41_759 ();
 sg13g2_fill_2 FILLER_41_763 ();
 sg13g2_fill_2 FILLER_41_786 ();
 sg13g2_fill_1 FILLER_41_788 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_8 FILLER_41_800 ();
 sg13g2_decap_8 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_fill_1 FILLER_41_821 ();
 sg13g2_decap_8 FILLER_41_827 ();
 sg13g2_decap_4 FILLER_41_834 ();
 sg13g2_decap_4 FILLER_41_846 ();
 sg13g2_fill_1 FILLER_41_850 ();
 sg13g2_fill_1 FILLER_41_858 ();
 sg13g2_decap_4 FILLER_41_877 ();
 sg13g2_decap_8 FILLER_41_885 ();
 sg13g2_decap_8 FILLER_41_892 ();
 sg13g2_decap_8 FILLER_41_899 ();
 sg13g2_decap_8 FILLER_41_906 ();
 sg13g2_decap_8 FILLER_41_913 ();
 sg13g2_decap_8 FILLER_41_920 ();
 sg13g2_decap_8 FILLER_41_927 ();
 sg13g2_fill_2 FILLER_41_934 ();
 sg13g2_decap_8 FILLER_41_939 ();
 sg13g2_decap_4 FILLER_41_946 ();
 sg13g2_fill_1 FILLER_41_950 ();
 sg13g2_decap_4 FILLER_41_957 ();
 sg13g2_decap_4 FILLER_41_965 ();
 sg13g2_fill_2 FILLER_41_987 ();
 sg13g2_fill_1 FILLER_41_989 ();
 sg13g2_decap_8 FILLER_41_999 ();
 sg13g2_decap_4 FILLER_41_1006 ();
 sg13g2_decap_8 FILLER_41_1018 ();
 sg13g2_decap_8 FILLER_41_1025 ();
 sg13g2_decap_8 FILLER_41_1032 ();
 sg13g2_fill_2 FILLER_41_1039 ();
 sg13g2_decap_4 FILLER_41_1049 ();
 sg13g2_fill_1 FILLER_41_1053 ();
 sg13g2_decap_4 FILLER_41_1064 ();
 sg13g2_fill_1 FILLER_41_1068 ();
 sg13g2_decap_4 FILLER_41_1074 ();
 sg13g2_fill_1 FILLER_41_1078 ();
 sg13g2_decap_8 FILLER_41_1087 ();
 sg13g2_decap_8 FILLER_41_1094 ();
 sg13g2_decap_8 FILLER_41_1101 ();
 sg13g2_decap_4 FILLER_41_1108 ();
 sg13g2_fill_2 FILLER_41_1112 ();
 sg13g2_fill_1 FILLER_41_1117 ();
 sg13g2_decap_4 FILLER_41_1149 ();
 sg13g2_fill_2 FILLER_41_1153 ();
 sg13g2_decap_4 FILLER_41_1181 ();
 sg13g2_fill_1 FILLER_41_1185 ();
 sg13g2_decap_8 FILLER_41_1227 ();
 sg13g2_decap_8 FILLER_41_1234 ();
 sg13g2_decap_8 FILLER_41_1241 ();
 sg13g2_decap_8 FILLER_41_1248 ();
 sg13g2_decap_8 FILLER_41_1255 ();
 sg13g2_decap_8 FILLER_41_1262 ();
 sg13g2_fill_1 FILLER_41_1281 ();
 sg13g2_fill_1 FILLER_41_1286 ();
 sg13g2_decap_4 FILLER_41_1313 ();
 sg13g2_fill_1 FILLER_41_1317 ();
 sg13g2_decap_8 FILLER_41_1326 ();
 sg13g2_fill_2 FILLER_41_1338 ();
 sg13g2_fill_2 FILLER_41_1343 ();
 sg13g2_fill_1 FILLER_41_1345 ();
 sg13g2_decap_4 FILLER_41_1350 ();
 sg13g2_fill_1 FILLER_41_1354 ();
 sg13g2_decap_8 FILLER_41_1385 ();
 sg13g2_decap_8 FILLER_41_1395 ();
 sg13g2_decap_8 FILLER_41_1402 ();
 sg13g2_decap_8 FILLER_41_1409 ();
 sg13g2_fill_1 FILLER_41_1416 ();
 sg13g2_decap_4 FILLER_41_1425 ();
 sg13g2_fill_1 FILLER_41_1429 ();
 sg13g2_decap_8 FILLER_41_1438 ();
 sg13g2_fill_2 FILLER_41_1479 ();
 sg13g2_fill_1 FILLER_41_1489 ();
 sg13g2_fill_1 FILLER_41_1494 ();
 sg13g2_fill_1 FILLER_41_1502 ();
 sg13g2_fill_1 FILLER_41_1529 ();
 sg13g2_decap_8 FILLER_41_1541 ();
 sg13g2_decap_8 FILLER_41_1548 ();
 sg13g2_decap_8 FILLER_41_1555 ();
 sg13g2_fill_2 FILLER_41_1562 ();
 sg13g2_fill_1 FILLER_41_1564 ();
 sg13g2_decap_4 FILLER_41_1571 ();
 sg13g2_fill_1 FILLER_41_1575 ();
 sg13g2_decap_8 FILLER_41_1580 ();
 sg13g2_decap_8 FILLER_41_1621 ();
 sg13g2_decap_8 FILLER_41_1628 ();
 sg13g2_decap_8 FILLER_41_1635 ();
 sg13g2_fill_1 FILLER_41_1642 ();
 sg13g2_decap_8 FILLER_41_1647 ();
 sg13g2_decap_8 FILLER_41_1654 ();
 sg13g2_decap_8 FILLER_41_1661 ();
 sg13g2_fill_2 FILLER_41_1668 ();
 sg13g2_fill_1 FILLER_41_1670 ();
 sg13g2_decap_8 FILLER_41_1675 ();
 sg13g2_decap_8 FILLER_41_1682 ();
 sg13g2_decap_8 FILLER_41_1689 ();
 sg13g2_decap_8 FILLER_41_1696 ();
 sg13g2_fill_2 FILLER_41_1703 ();
 sg13g2_fill_1 FILLER_41_1718 ();
 sg13g2_decap_4 FILLER_41_1724 ();
 sg13g2_fill_1 FILLER_41_1728 ();
 sg13g2_fill_1 FILLER_41_1741 ();
 sg13g2_fill_1 FILLER_41_1773 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_4 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_39 ();
 sg13g2_decap_8 FILLER_42_54 ();
 sg13g2_fill_1 FILLER_42_61 ();
 sg13g2_decap_4 FILLER_42_71 ();
 sg13g2_fill_1 FILLER_42_75 ();
 sg13g2_decap_4 FILLER_42_81 ();
 sg13g2_fill_2 FILLER_42_85 ();
 sg13g2_fill_1 FILLER_42_91 ();
 sg13g2_fill_1 FILLER_42_105 ();
 sg13g2_fill_2 FILLER_42_110 ();
 sg13g2_fill_1 FILLER_42_112 ();
 sg13g2_fill_2 FILLER_42_117 ();
 sg13g2_decap_4 FILLER_42_123 ();
 sg13g2_fill_1 FILLER_42_132 ();
 sg13g2_fill_1 FILLER_42_141 ();
 sg13g2_decap_8 FILLER_42_151 ();
 sg13g2_decap_4 FILLER_42_158 ();
 sg13g2_fill_2 FILLER_42_162 ();
 sg13g2_fill_1 FILLER_42_174 ();
 sg13g2_fill_1 FILLER_42_179 ();
 sg13g2_fill_1 FILLER_42_184 ();
 sg13g2_fill_1 FILLER_42_190 ();
 sg13g2_decap_8 FILLER_42_195 ();
 sg13g2_decap_8 FILLER_42_202 ();
 sg13g2_decap_4 FILLER_42_233 ();
 sg13g2_fill_2 FILLER_42_237 ();
 sg13g2_fill_2 FILLER_42_243 ();
 sg13g2_fill_1 FILLER_42_245 ();
 sg13g2_fill_2 FILLER_42_250 ();
 sg13g2_fill_1 FILLER_42_252 ();
 sg13g2_fill_2 FILLER_42_259 ();
 sg13g2_fill_2 FILLER_42_282 ();
 sg13g2_fill_1 FILLER_42_289 ();
 sg13g2_decap_4 FILLER_42_300 ();
 sg13g2_fill_1 FILLER_42_304 ();
 sg13g2_decap_8 FILLER_42_317 ();
 sg13g2_decap_4 FILLER_42_324 ();
 sg13g2_decap_8 FILLER_42_333 ();
 sg13g2_fill_2 FILLER_42_340 ();
 sg13g2_fill_1 FILLER_42_342 ();
 sg13g2_fill_2 FILLER_42_347 ();
 sg13g2_fill_1 FILLER_42_349 ();
 sg13g2_decap_8 FILLER_42_360 ();
 sg13g2_fill_2 FILLER_42_367 ();
 sg13g2_fill_1 FILLER_42_369 ();
 sg13g2_fill_2 FILLER_42_376 ();
 sg13g2_decap_8 FILLER_42_382 ();
 sg13g2_fill_1 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_395 ();
 sg13g2_decap_4 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_42_429 ();
 sg13g2_decap_8 FILLER_42_436 ();
 sg13g2_decap_8 FILLER_42_443 ();
 sg13g2_decap_8 FILLER_42_450 ();
 sg13g2_decap_8 FILLER_42_457 ();
 sg13g2_fill_2 FILLER_42_464 ();
 sg13g2_fill_1 FILLER_42_466 ();
 sg13g2_decap_8 FILLER_42_470 ();
 sg13g2_decap_8 FILLER_42_477 ();
 sg13g2_decap_8 FILLER_42_484 ();
 sg13g2_fill_2 FILLER_42_491 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_decap_4 FILLER_42_516 ();
 sg13g2_decap_4 FILLER_42_524 ();
 sg13g2_decap_8 FILLER_42_532 ();
 sg13g2_decap_8 FILLER_42_539 ();
 sg13g2_decap_8 FILLER_42_546 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_564 ();
 sg13g2_decap_8 FILLER_42_571 ();
 sg13g2_decap_8 FILLER_42_578 ();
 sg13g2_fill_2 FILLER_42_585 ();
 sg13g2_fill_1 FILLER_42_587 ();
 sg13g2_decap_8 FILLER_42_614 ();
 sg13g2_decap_8 FILLER_42_629 ();
 sg13g2_decap_8 FILLER_42_636 ();
 sg13g2_fill_2 FILLER_42_643 ();
 sg13g2_fill_2 FILLER_42_649 ();
 sg13g2_fill_1 FILLER_42_651 ();
 sg13g2_decap_8 FILLER_42_655 ();
 sg13g2_decap_8 FILLER_42_662 ();
 sg13g2_decap_8 FILLER_42_682 ();
 sg13g2_decap_8 FILLER_42_689 ();
 sg13g2_decap_8 FILLER_42_696 ();
 sg13g2_fill_1 FILLER_42_703 ();
 sg13g2_decap_8 FILLER_42_708 ();
 sg13g2_decap_4 FILLER_42_715 ();
 sg13g2_fill_1 FILLER_42_719 ();
 sg13g2_fill_1 FILLER_42_739 ();
 sg13g2_decap_8 FILLER_42_757 ();
 sg13g2_decap_4 FILLER_42_764 ();
 sg13g2_fill_1 FILLER_42_768 ();
 sg13g2_decap_8 FILLER_42_795 ();
 sg13g2_decap_8 FILLER_42_802 ();
 sg13g2_fill_2 FILLER_42_809 ();
 sg13g2_fill_1 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_816 ();
 sg13g2_fill_2 FILLER_42_827 ();
 sg13g2_decap_8 FILLER_42_834 ();
 sg13g2_fill_2 FILLER_42_844 ();
 sg13g2_fill_1 FILLER_42_846 ();
 sg13g2_fill_1 FILLER_42_857 ();
 sg13g2_fill_2 FILLER_42_863 ();
 sg13g2_fill_2 FILLER_42_870 ();
 sg13g2_fill_1 FILLER_42_872 ();
 sg13g2_decap_4 FILLER_42_877 ();
 sg13g2_fill_1 FILLER_42_886 ();
 sg13g2_fill_2 FILLER_42_905 ();
 sg13g2_decap_8 FILLER_42_912 ();
 sg13g2_decap_8 FILLER_42_924 ();
 sg13g2_fill_1 FILLER_42_931 ();
 sg13g2_decap_4 FILLER_42_950 ();
 sg13g2_fill_1 FILLER_42_959 ();
 sg13g2_decap_8 FILLER_42_976 ();
 sg13g2_decap_8 FILLER_42_983 ();
 sg13g2_decap_4 FILLER_42_990 ();
 sg13g2_fill_2 FILLER_42_994 ();
 sg13g2_decap_8 FILLER_42_1016 ();
 sg13g2_fill_2 FILLER_42_1023 ();
 sg13g2_fill_1 FILLER_42_1025 ();
 sg13g2_decap_4 FILLER_42_1033 ();
 sg13g2_fill_2 FILLER_42_1037 ();
 sg13g2_decap_4 FILLER_42_1042 ();
 sg13g2_fill_2 FILLER_42_1059 ();
 sg13g2_fill_1 FILLER_42_1061 ();
 sg13g2_fill_2 FILLER_42_1068 ();
 sg13g2_fill_1 FILLER_42_1080 ();
 sg13g2_decap_8 FILLER_42_1100 ();
 sg13g2_fill_2 FILLER_42_1107 ();
 sg13g2_fill_1 FILLER_42_1109 ();
 sg13g2_decap_8 FILLER_42_1123 ();
 sg13g2_decap_8 FILLER_42_1130 ();
 sg13g2_decap_8 FILLER_42_1137 ();
 sg13g2_decap_8 FILLER_42_1144 ();
 sg13g2_fill_1 FILLER_42_1151 ();
 sg13g2_decap_8 FILLER_42_1157 ();
 sg13g2_decap_8 FILLER_42_1164 ();
 sg13g2_decap_4 FILLER_42_1171 ();
 sg13g2_fill_2 FILLER_42_1175 ();
 sg13g2_fill_1 FILLER_42_1181 ();
 sg13g2_fill_1 FILLER_42_1187 ();
 sg13g2_decap_4 FILLER_42_1193 ();
 sg13g2_decap_4 FILLER_42_1202 ();
 sg13g2_fill_1 FILLER_42_1206 ();
 sg13g2_decap_8 FILLER_42_1211 ();
 sg13g2_decap_8 FILLER_42_1218 ();
 sg13g2_decap_4 FILLER_42_1225 ();
 sg13g2_fill_1 FILLER_42_1229 ();
 sg13g2_decap_4 FILLER_42_1237 ();
 sg13g2_decap_8 FILLER_42_1250 ();
 sg13g2_decap_8 FILLER_42_1257 ();
 sg13g2_fill_2 FILLER_42_1264 ();
 sg13g2_decap_4 FILLER_42_1273 ();
 sg13g2_fill_1 FILLER_42_1277 ();
 sg13g2_decap_8 FILLER_42_1282 ();
 sg13g2_decap_8 FILLER_42_1289 ();
 sg13g2_decap_4 FILLER_42_1296 ();
 sg13g2_fill_1 FILLER_42_1300 ();
 sg13g2_decap_8 FILLER_42_1305 ();
 sg13g2_decap_8 FILLER_42_1312 ();
 sg13g2_decap_4 FILLER_42_1319 ();
 sg13g2_fill_1 FILLER_42_1323 ();
 sg13g2_decap_4 FILLER_42_1336 ();
 sg13g2_fill_2 FILLER_42_1340 ();
 sg13g2_decap_8 FILLER_42_1353 ();
 sg13g2_fill_2 FILLER_42_1360 ();
 sg13g2_fill_2 FILLER_42_1386 ();
 sg13g2_fill_1 FILLER_42_1388 ();
 sg13g2_decap_8 FILLER_42_1419 ();
 sg13g2_decap_4 FILLER_42_1426 ();
 sg13g2_fill_1 FILLER_42_1430 ();
 sg13g2_decap_8 FILLER_42_1435 ();
 sg13g2_decap_4 FILLER_42_1442 ();
 sg13g2_fill_2 FILLER_42_1446 ();
 sg13g2_fill_1 FILLER_42_1454 ();
 sg13g2_decap_8 FILLER_42_1459 ();
 sg13g2_decap_8 FILLER_42_1466 ();
 sg13g2_decap_8 FILLER_42_1473 ();
 sg13g2_decap_4 FILLER_42_1480 ();
 sg13g2_decap_8 FILLER_42_1490 ();
 sg13g2_decap_8 FILLER_42_1497 ();
 sg13g2_decap_4 FILLER_42_1504 ();
 sg13g2_fill_1 FILLER_42_1508 ();
 sg13g2_decap_8 FILLER_42_1513 ();
 sg13g2_decap_8 FILLER_42_1520 ();
 sg13g2_decap_8 FILLER_42_1527 ();
 sg13g2_decap_8 FILLER_42_1542 ();
 sg13g2_decap_8 FILLER_42_1549 ();
 sg13g2_decap_4 FILLER_42_1556 ();
 sg13g2_fill_2 FILLER_42_1560 ();
 sg13g2_decap_8 FILLER_42_1566 ();
 sg13g2_decap_8 FILLER_42_1573 ();
 sg13g2_decap_4 FILLER_42_1580 ();
 sg13g2_fill_1 FILLER_42_1584 ();
 sg13g2_decap_8 FILLER_42_1595 ();
 sg13g2_fill_2 FILLER_42_1602 ();
 sg13g2_fill_1 FILLER_42_1604 ();
 sg13g2_decap_8 FILLER_42_1634 ();
 sg13g2_decap_4 FILLER_42_1641 ();
 sg13g2_decap_8 FILLER_42_1649 ();
 sg13g2_fill_1 FILLER_42_1656 ();
 sg13g2_decap_4 FILLER_42_1670 ();
 sg13g2_fill_2 FILLER_42_1674 ();
 sg13g2_decap_8 FILLER_42_1680 ();
 sg13g2_decap_8 FILLER_42_1687 ();
 sg13g2_decap_4 FILLER_42_1694 ();
 sg13g2_fill_2 FILLER_42_1698 ();
 sg13g2_fill_2 FILLER_42_1708 ();
 sg13g2_fill_2 FILLER_42_1723 ();
 sg13g2_decap_8 FILLER_42_1730 ();
 sg13g2_decap_8 FILLER_42_1737 ();
 sg13g2_decap_8 FILLER_42_1744 ();
 sg13g2_fill_2 FILLER_42_1751 ();
 sg13g2_fill_1 FILLER_42_1753 ();
 sg13g2_decap_4 FILLER_42_1758 ();
 sg13g2_decap_8 FILLER_42_1766 ();
 sg13g2_fill_1 FILLER_42_1773 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_4 FILLER_43_35 ();
 sg13g2_fill_1 FILLER_43_39 ();
 sg13g2_fill_2 FILLER_43_44 ();
 sg13g2_fill_2 FILLER_43_51 ();
 sg13g2_decap_8 FILLER_43_62 ();
 sg13g2_decap_8 FILLER_43_69 ();
 sg13g2_decap_4 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_80 ();
 sg13g2_fill_2 FILLER_43_86 ();
 sg13g2_decap_4 FILLER_43_100 ();
 sg13g2_decap_4 FILLER_43_109 ();
 sg13g2_decap_4 FILLER_43_121 ();
 sg13g2_fill_1 FILLER_43_125 ();
 sg13g2_fill_1 FILLER_43_131 ();
 sg13g2_decap_8 FILLER_43_137 ();
 sg13g2_fill_1 FILLER_43_144 ();
 sg13g2_decap_8 FILLER_43_150 ();
 sg13g2_decap_4 FILLER_43_157 ();
 sg13g2_decap_8 FILLER_43_173 ();
 sg13g2_fill_2 FILLER_43_180 ();
 sg13g2_fill_1 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_187 ();
 sg13g2_fill_2 FILLER_43_194 ();
 sg13g2_fill_1 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_201 ();
 sg13g2_decap_8 FILLER_43_208 ();
 sg13g2_decap_8 FILLER_43_215 ();
 sg13g2_decap_8 FILLER_43_222 ();
 sg13g2_decap_4 FILLER_43_237 ();
 sg13g2_decap_8 FILLER_43_246 ();
 sg13g2_decap_8 FILLER_43_253 ();
 sg13g2_decap_8 FILLER_43_260 ();
 sg13g2_fill_2 FILLER_43_267 ();
 sg13g2_fill_1 FILLER_43_269 ();
 sg13g2_decap_4 FILLER_43_284 ();
 sg13g2_fill_1 FILLER_43_288 ();
 sg13g2_fill_2 FILLER_43_295 ();
 sg13g2_fill_1 FILLER_43_297 ();
 sg13g2_decap_8 FILLER_43_303 ();
 sg13g2_decap_8 FILLER_43_310 ();
 sg13g2_decap_8 FILLER_43_317 ();
 sg13g2_decap_8 FILLER_43_324 ();
 sg13g2_fill_2 FILLER_43_331 ();
 sg13g2_fill_1 FILLER_43_333 ();
 sg13g2_fill_2 FILLER_43_348 ();
 sg13g2_fill_1 FILLER_43_350 ();
 sg13g2_fill_1 FILLER_43_362 ();
 sg13g2_decap_4 FILLER_43_373 ();
 sg13g2_decap_8 FILLER_43_381 ();
 sg13g2_fill_1 FILLER_43_388 ();
 sg13g2_decap_4 FILLER_43_394 ();
 sg13g2_fill_2 FILLER_43_398 ();
 sg13g2_decap_4 FILLER_43_404 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_43_440 ();
 sg13g2_decap_4 FILLER_43_447 ();
 sg13g2_decap_8 FILLER_43_457 ();
 sg13g2_decap_8 FILLER_43_464 ();
 sg13g2_decap_8 FILLER_43_471 ();
 sg13g2_decap_4 FILLER_43_478 ();
 sg13g2_fill_2 FILLER_43_482 ();
 sg13g2_fill_2 FILLER_43_513 ();
 sg13g2_fill_1 FILLER_43_515 ();
 sg13g2_fill_2 FILLER_43_547 ();
 sg13g2_fill_2 FILLER_43_584 ();
 sg13g2_fill_1 FILLER_43_586 ();
 sg13g2_decap_4 FILLER_43_592 ();
 sg13g2_fill_2 FILLER_43_600 ();
 sg13g2_fill_1 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_606 ();
 sg13g2_decap_8 FILLER_43_613 ();
 sg13g2_decap_8 FILLER_43_633 ();
 sg13g2_decap_4 FILLER_43_640 ();
 sg13g2_fill_2 FILLER_43_666 ();
 sg13g2_fill_1 FILLER_43_668 ();
 sg13g2_decap_4 FILLER_43_678 ();
 sg13g2_decap_8 FILLER_43_687 ();
 sg13g2_decap_8 FILLER_43_694 ();
 sg13g2_decap_8 FILLER_43_701 ();
 sg13g2_decap_8 FILLER_43_708 ();
 sg13g2_decap_8 FILLER_43_715 ();
 sg13g2_decap_4 FILLER_43_722 ();
 sg13g2_fill_2 FILLER_43_726 ();
 sg13g2_fill_2 FILLER_43_732 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_4 FILLER_43_777 ();
 sg13g2_fill_2 FILLER_43_781 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_fill_2 FILLER_43_847 ();
 sg13g2_fill_1 FILLER_43_849 ();
 sg13g2_fill_1 FILLER_43_854 ();
 sg13g2_fill_1 FILLER_43_858 ();
 sg13g2_decap_8 FILLER_43_863 ();
 sg13g2_decap_8 FILLER_43_870 ();
 sg13g2_decap_8 FILLER_43_885 ();
 sg13g2_decap_4 FILLER_43_892 ();
 sg13g2_fill_2 FILLER_43_896 ();
 sg13g2_decap_4 FILLER_43_905 ();
 sg13g2_fill_1 FILLER_43_909 ();
 sg13g2_decap_8 FILLER_43_923 ();
 sg13g2_decap_4 FILLER_43_930 ();
 sg13g2_fill_2 FILLER_43_934 ();
 sg13g2_fill_1 FILLER_43_944 ();
 sg13g2_decap_8 FILLER_43_958 ();
 sg13g2_fill_1 FILLER_43_965 ();
 sg13g2_fill_1 FILLER_43_981 ();
 sg13g2_decap_8 FILLER_43_987 ();
 sg13g2_decap_4 FILLER_43_994 ();
 sg13g2_fill_2 FILLER_43_998 ();
 sg13g2_fill_1 FILLER_43_1030 ();
 sg13g2_fill_2 FILLER_43_1035 ();
 sg13g2_decap_4 FILLER_43_1044 ();
 sg13g2_decap_8 FILLER_43_1062 ();
 sg13g2_decap_8 FILLER_43_1069 ();
 sg13g2_decap_8 FILLER_43_1086 ();
 sg13g2_decap_8 FILLER_43_1093 ();
 sg13g2_fill_2 FILLER_43_1100 ();
 sg13g2_decap_8 FILLER_43_1111 ();
 sg13g2_decap_8 FILLER_43_1123 ();
 sg13g2_decap_8 FILLER_43_1130 ();
 sg13g2_fill_1 FILLER_43_1137 ();
 sg13g2_fill_2 FILLER_43_1146 ();
 sg13g2_decap_8 FILLER_43_1187 ();
 sg13g2_fill_2 FILLER_43_1194 ();
 sg13g2_fill_1 FILLER_43_1196 ();
 sg13g2_decap_8 FILLER_43_1219 ();
 sg13g2_fill_1 FILLER_43_1226 ();
 sg13g2_decap_4 FILLER_43_1235 ();
 sg13g2_fill_1 FILLER_43_1239 ();
 sg13g2_fill_2 FILLER_43_1266 ();
 sg13g2_decap_4 FILLER_43_1272 ();
 sg13g2_fill_2 FILLER_43_1276 ();
 sg13g2_decap_8 FILLER_43_1283 ();
 sg13g2_decap_4 FILLER_43_1290 ();
 sg13g2_decap_8 FILLER_43_1320 ();
 sg13g2_decap_8 FILLER_43_1327 ();
 sg13g2_fill_2 FILLER_43_1334 ();
 sg13g2_fill_1 FILLER_43_1336 ();
 sg13g2_decap_8 FILLER_43_1344 ();
 sg13g2_decap_8 FILLER_43_1351 ();
 sg13g2_decap_8 FILLER_43_1358 ();
 sg13g2_decap_8 FILLER_43_1384 ();
 sg13g2_fill_1 FILLER_43_1391 ();
 sg13g2_decap_8 FILLER_43_1398 ();
 sg13g2_decap_8 FILLER_43_1405 ();
 sg13g2_decap_8 FILLER_43_1412 ();
 sg13g2_decap_8 FILLER_43_1419 ();
 sg13g2_fill_2 FILLER_43_1426 ();
 sg13g2_decap_8 FILLER_43_1445 ();
 sg13g2_decap_8 FILLER_43_1452 ();
 sg13g2_decap_8 FILLER_43_1459 ();
 sg13g2_fill_2 FILLER_43_1466 ();
 sg13g2_decap_8 FILLER_43_1472 ();
 sg13g2_decap_8 FILLER_43_1479 ();
 sg13g2_decap_8 FILLER_43_1486 ();
 sg13g2_decap_8 FILLER_43_1493 ();
 sg13g2_fill_2 FILLER_43_1500 ();
 sg13g2_decap_8 FILLER_43_1507 ();
 sg13g2_decap_8 FILLER_43_1514 ();
 sg13g2_decap_8 FILLER_43_1521 ();
 sg13g2_decap_8 FILLER_43_1534 ();
 sg13g2_decap_8 FILLER_43_1541 ();
 sg13g2_decap_4 FILLER_43_1548 ();
 sg13g2_decap_8 FILLER_43_1581 ();
 sg13g2_decap_8 FILLER_43_1588 ();
 sg13g2_decap_8 FILLER_43_1595 ();
 sg13g2_decap_8 FILLER_43_1602 ();
 sg13g2_decap_4 FILLER_43_1609 ();
 sg13g2_decap_8 FILLER_43_1617 ();
 sg13g2_decap_8 FILLER_43_1624 ();
 sg13g2_decap_4 FILLER_43_1631 ();
 sg13g2_fill_1 FILLER_43_1635 ();
 sg13g2_decap_8 FILLER_43_1662 ();
 sg13g2_decap_8 FILLER_43_1698 ();
 sg13g2_decap_8 FILLER_43_1705 ();
 sg13g2_fill_1 FILLER_43_1712 ();
 sg13g2_decap_8 FILLER_43_1730 ();
 sg13g2_fill_2 FILLER_43_1737 ();
 sg13g2_fill_1 FILLER_43_1739 ();
 sg13g2_decap_8 FILLER_43_1748 ();
 sg13g2_decap_8 FILLER_43_1755 ();
 sg13g2_decap_8 FILLER_43_1762 ();
 sg13g2_decap_4 FILLER_43_1769 ();
 sg13g2_fill_1 FILLER_43_1773 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_fill_2 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_44 ();
 sg13g2_fill_2 FILLER_44_50 ();
 sg13g2_decap_8 FILLER_44_57 ();
 sg13g2_decap_8 FILLER_44_64 ();
 sg13g2_decap_8 FILLER_44_71 ();
 sg13g2_decap_8 FILLER_44_78 ();
 sg13g2_fill_2 FILLER_44_85 ();
 sg13g2_decap_4 FILLER_44_95 ();
 sg13g2_decap_4 FILLER_44_103 ();
 sg13g2_fill_2 FILLER_44_107 ();
 sg13g2_decap_4 FILLER_44_113 ();
 sg13g2_decap_8 FILLER_44_127 ();
 sg13g2_decap_4 FILLER_44_134 ();
 sg13g2_fill_1 FILLER_44_138 ();
 sg13g2_decap_8 FILLER_44_143 ();
 sg13g2_fill_1 FILLER_44_150 ();
 sg13g2_decap_4 FILLER_44_155 ();
 sg13g2_fill_1 FILLER_44_159 ();
 sg13g2_fill_2 FILLER_44_164 ();
 sg13g2_fill_2 FILLER_44_185 ();
 sg13g2_fill_2 FILLER_44_193 ();
 sg13g2_fill_1 FILLER_44_200 ();
 sg13g2_fill_2 FILLER_44_216 ();
 sg13g2_fill_1 FILLER_44_222 ();
 sg13g2_fill_2 FILLER_44_227 ();
 sg13g2_fill_1 FILLER_44_239 ();
 sg13g2_fill_1 FILLER_44_250 ();
 sg13g2_fill_1 FILLER_44_255 ();
 sg13g2_fill_2 FILLER_44_280 ();
 sg13g2_fill_1 FILLER_44_282 ();
 sg13g2_fill_1 FILLER_44_292 ();
 sg13g2_fill_1 FILLER_44_297 ();
 sg13g2_fill_2 FILLER_44_302 ();
 sg13g2_decap_8 FILLER_44_316 ();
 sg13g2_decap_8 FILLER_44_323 ();
 sg13g2_fill_2 FILLER_44_330 ();
 sg13g2_fill_1 FILLER_44_332 ();
 sg13g2_decap_4 FILLER_44_341 ();
 sg13g2_fill_2 FILLER_44_345 ();
 sg13g2_decap_8 FILLER_44_351 ();
 sg13g2_decap_4 FILLER_44_358 ();
 sg13g2_fill_2 FILLER_44_372 ();
 sg13g2_decap_8 FILLER_44_379 ();
 sg13g2_decap_8 FILLER_44_386 ();
 sg13g2_fill_2 FILLER_44_393 ();
 sg13g2_fill_2 FILLER_44_400 ();
 sg13g2_fill_1 FILLER_44_402 ();
 sg13g2_fill_1 FILLER_44_410 ();
 sg13g2_fill_1 FILLER_44_428 ();
 sg13g2_decap_4 FILLER_44_435 ();
 sg13g2_decap_8 FILLER_44_447 ();
 sg13g2_decap_8 FILLER_44_454 ();
 sg13g2_decap_8 FILLER_44_461 ();
 sg13g2_decap_8 FILLER_44_468 ();
 sg13g2_decap_8 FILLER_44_492 ();
 sg13g2_decap_8 FILLER_44_499 ();
 sg13g2_decap_4 FILLER_44_506 ();
 sg13g2_fill_2 FILLER_44_513 ();
 sg13g2_fill_1 FILLER_44_515 ();
 sg13g2_decap_8 FILLER_44_533 ();
 sg13g2_decap_8 FILLER_44_540 ();
 sg13g2_decap_8 FILLER_44_547 ();
 sg13g2_decap_8 FILLER_44_554 ();
 sg13g2_decap_8 FILLER_44_561 ();
 sg13g2_decap_8 FILLER_44_568 ();
 sg13g2_decap_8 FILLER_44_575 ();
 sg13g2_decap_8 FILLER_44_582 ();
 sg13g2_decap_8 FILLER_44_589 ();
 sg13g2_decap_8 FILLER_44_596 ();
 sg13g2_decap_8 FILLER_44_607 ();
 sg13g2_decap_8 FILLER_44_614 ();
 sg13g2_decap_8 FILLER_44_621 ();
 sg13g2_decap_8 FILLER_44_628 ();
 sg13g2_fill_2 FILLER_44_635 ();
 sg13g2_fill_1 FILLER_44_637 ();
 sg13g2_decap_8 FILLER_44_643 ();
 sg13g2_fill_2 FILLER_44_650 ();
 sg13g2_decap_8 FILLER_44_659 ();
 sg13g2_decap_8 FILLER_44_666 ();
 sg13g2_fill_1 FILLER_44_673 ();
 sg13g2_fill_1 FILLER_44_679 ();
 sg13g2_fill_2 FILLER_44_685 ();
 sg13g2_decap_8 FILLER_44_695 ();
 sg13g2_decap_8 FILLER_44_702 ();
 sg13g2_decap_8 FILLER_44_709 ();
 sg13g2_decap_8 FILLER_44_716 ();
 sg13g2_decap_8 FILLER_44_723 ();
 sg13g2_decap_8 FILLER_44_730 ();
 sg13g2_fill_2 FILLER_44_737 ();
 sg13g2_decap_8 FILLER_44_743 ();
 sg13g2_fill_1 FILLER_44_750 ();
 sg13g2_decap_4 FILLER_44_754 ();
 sg13g2_fill_1 FILLER_44_758 ();
 sg13g2_decap_8 FILLER_44_774 ();
 sg13g2_decap_4 FILLER_44_781 ();
 sg13g2_decap_4 FILLER_44_789 ();
 sg13g2_fill_2 FILLER_44_793 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_fill_2 FILLER_44_833 ();
 sg13g2_fill_1 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_853 ();
 sg13g2_decap_8 FILLER_44_860 ();
 sg13g2_decap_4 FILLER_44_867 ();
 sg13g2_fill_1 FILLER_44_876 ();
 sg13g2_decap_8 FILLER_44_881 ();
 sg13g2_decap_4 FILLER_44_888 ();
 sg13g2_decap_8 FILLER_44_908 ();
 sg13g2_decap_8 FILLER_44_915 ();
 sg13g2_decap_8 FILLER_44_922 ();
 sg13g2_decap_8 FILLER_44_929 ();
 sg13g2_fill_2 FILLER_44_936 ();
 sg13g2_fill_2 FILLER_44_957 ();
 sg13g2_fill_2 FILLER_44_974 ();
 sg13g2_fill_1 FILLER_44_976 ();
 sg13g2_decap_4 FILLER_44_981 ();
 sg13g2_decap_4 FILLER_44_995 ();
 sg13g2_fill_2 FILLER_44_999 ();
 sg13g2_decap_4 FILLER_44_1006 ();
 sg13g2_fill_1 FILLER_44_1010 ();
 sg13g2_decap_8 FILLER_44_1020 ();
 sg13g2_fill_2 FILLER_44_1027 ();
 sg13g2_fill_2 FILLER_44_1050 ();
 sg13g2_fill_1 FILLER_44_1052 ();
 sg13g2_decap_8 FILLER_44_1058 ();
 sg13g2_decap_8 FILLER_44_1065 ();
 sg13g2_decap_8 FILLER_44_1072 ();
 sg13g2_decap_8 FILLER_44_1079 ();
 sg13g2_decap_4 FILLER_44_1086 ();
 sg13g2_fill_1 FILLER_44_1090 ();
 sg13g2_decap_8 FILLER_44_1103 ();
 sg13g2_decap_8 FILLER_44_1110 ();
 sg13g2_decap_4 FILLER_44_1117 ();
 sg13g2_fill_1 FILLER_44_1121 ();
 sg13g2_decap_8 FILLER_44_1132 ();
 sg13g2_decap_8 FILLER_44_1139 ();
 sg13g2_decap_8 FILLER_44_1146 ();
 sg13g2_fill_2 FILLER_44_1161 ();
 sg13g2_decap_8 FILLER_44_1168 ();
 sg13g2_decap_8 FILLER_44_1179 ();
 sg13g2_decap_8 FILLER_44_1186 ();
 sg13g2_fill_2 FILLER_44_1193 ();
 sg13g2_decap_8 FILLER_44_1226 ();
 sg13g2_decap_8 FILLER_44_1233 ();
 sg13g2_fill_2 FILLER_44_1240 ();
 sg13g2_fill_1 FILLER_44_1242 ();
 sg13g2_decap_8 FILLER_44_1247 ();
 sg13g2_decap_8 FILLER_44_1254 ();
 sg13g2_decap_8 FILLER_44_1261 ();
 sg13g2_decap_4 FILLER_44_1268 ();
 sg13g2_decap_4 FILLER_44_1283 ();
 sg13g2_fill_2 FILLER_44_1287 ();
 sg13g2_decap_8 FILLER_44_1294 ();
 sg13g2_decap_8 FILLER_44_1301 ();
 sg13g2_fill_2 FILLER_44_1308 ();
 sg13g2_decap_8 FILLER_44_1313 ();
 sg13g2_decap_8 FILLER_44_1320 ();
 sg13g2_decap_8 FILLER_44_1327 ();
 sg13g2_decap_8 FILLER_44_1334 ();
 sg13g2_decap_8 FILLER_44_1341 ();
 sg13g2_decap_4 FILLER_44_1348 ();
 sg13g2_decap_8 FILLER_44_1384 ();
 sg13g2_decap_8 FILLER_44_1391 ();
 sg13g2_decap_8 FILLER_44_1402 ();
 sg13g2_decap_8 FILLER_44_1409 ();
 sg13g2_decap_8 FILLER_44_1416 ();
 sg13g2_fill_2 FILLER_44_1423 ();
 sg13g2_decap_4 FILLER_44_1456 ();
 sg13g2_fill_1 FILLER_44_1460 ();
 sg13g2_fill_2 FILLER_44_1487 ();
 sg13g2_fill_2 FILLER_44_1497 ();
 sg13g2_fill_1 FILLER_44_1523 ();
 sg13g2_fill_1 FILLER_44_1539 ();
 sg13g2_fill_1 FILLER_44_1545 ();
 sg13g2_decap_4 FILLER_44_1552 ();
 sg13g2_decap_8 FILLER_44_1585 ();
 sg13g2_decap_8 FILLER_44_1592 ();
 sg13g2_decap_8 FILLER_44_1605 ();
 sg13g2_fill_2 FILLER_44_1612 ();
 sg13g2_decap_8 FILLER_44_1620 ();
 sg13g2_decap_4 FILLER_44_1627 ();
 sg13g2_fill_2 FILLER_44_1631 ();
 sg13g2_decap_8 FILLER_44_1636 ();
 sg13g2_decap_8 FILLER_44_1643 ();
 sg13g2_decap_4 FILLER_44_1650 ();
 sg13g2_fill_1 FILLER_44_1654 ();
 sg13g2_decap_8 FILLER_44_1658 ();
 sg13g2_decap_8 FILLER_44_1665 ();
 sg13g2_decap_8 FILLER_44_1672 ();
 sg13g2_decap_8 FILLER_44_1679 ();
 sg13g2_decap_8 FILLER_44_1686 ();
 sg13g2_decap_8 FILLER_44_1693 ();
 sg13g2_decap_8 FILLER_44_1700 ();
 sg13g2_decap_8 FILLER_44_1707 ();
 sg13g2_decap_8 FILLER_44_1714 ();
 sg13g2_fill_2 FILLER_44_1721 ();
 sg13g2_decap_8 FILLER_44_1732 ();
 sg13g2_decap_8 FILLER_44_1751 ();
 sg13g2_decap_8 FILLER_44_1758 ();
 sg13g2_decap_8 FILLER_44_1765 ();
 sg13g2_fill_2 FILLER_44_1772 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_fill_2 FILLER_45_42 ();
 sg13g2_fill_2 FILLER_45_49 ();
 sg13g2_fill_2 FILLER_45_67 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_fill_2 FILLER_45_84 ();
 sg13g2_fill_2 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_119 ();
 sg13g2_fill_1 FILLER_45_121 ();
 sg13g2_decap_8 FILLER_45_130 ();
 sg13g2_decap_4 FILLER_45_137 ();
 sg13g2_fill_1 FILLER_45_156 ();
 sg13g2_fill_1 FILLER_45_176 ();
 sg13g2_decap_8 FILLER_45_192 ();
 sg13g2_fill_2 FILLER_45_199 ();
 sg13g2_decap_8 FILLER_45_205 ();
 sg13g2_decap_8 FILLER_45_212 ();
 sg13g2_fill_2 FILLER_45_219 ();
 sg13g2_decap_4 FILLER_45_231 ();
 sg13g2_decap_4 FILLER_45_240 ();
 sg13g2_fill_1 FILLER_45_244 ();
 sg13g2_decap_8 FILLER_45_250 ();
 sg13g2_decap_4 FILLER_45_257 ();
 sg13g2_fill_2 FILLER_45_261 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_decap_4 FILLER_45_278 ();
 sg13g2_fill_2 FILLER_45_282 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_fill_2 FILLER_45_301 ();
 sg13g2_decap_4 FILLER_45_308 ();
 sg13g2_fill_2 FILLER_45_317 ();
 sg13g2_fill_1 FILLER_45_319 ();
 sg13g2_decap_8 FILLER_45_339 ();
 sg13g2_decap_8 FILLER_45_346 ();
 sg13g2_fill_2 FILLER_45_353 ();
 sg13g2_fill_2 FILLER_45_360 ();
 sg13g2_fill_2 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_377 ();
 sg13g2_fill_2 FILLER_45_384 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_fill_1 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_404 ();
 sg13g2_fill_1 FILLER_45_411 ();
 sg13g2_fill_1 FILLER_45_417 ();
 sg13g2_decap_8 FILLER_45_428 ();
 sg13g2_fill_2 FILLER_45_445 ();
 sg13g2_decap_8 FILLER_45_452 ();
 sg13g2_decap_8 FILLER_45_459 ();
 sg13g2_decap_8 FILLER_45_466 ();
 sg13g2_decap_8 FILLER_45_473 ();
 sg13g2_decap_8 FILLER_45_480 ();
 sg13g2_decap_8 FILLER_45_487 ();
 sg13g2_decap_8 FILLER_45_494 ();
 sg13g2_decap_8 FILLER_45_501 ();
 sg13g2_decap_8 FILLER_45_508 ();
 sg13g2_fill_1 FILLER_45_515 ();
 sg13g2_decap_4 FILLER_45_545 ();
 sg13g2_fill_2 FILLER_45_549 ();
 sg13g2_fill_1 FILLER_45_556 ();
 sg13g2_decap_8 FILLER_45_587 ();
 sg13g2_fill_2 FILLER_45_594 ();
 sg13g2_decap_8 FILLER_45_625 ();
 sg13g2_decap_4 FILLER_45_632 ();
 sg13g2_fill_2 FILLER_45_636 ();
 sg13g2_fill_1 FILLER_45_642 ();
 sg13g2_decap_4 FILLER_45_651 ();
 sg13g2_decap_4 FILLER_45_659 ();
 sg13g2_fill_1 FILLER_45_663 ();
 sg13g2_fill_2 FILLER_45_668 ();
 sg13g2_fill_1 FILLER_45_670 ();
 sg13g2_fill_1 FILLER_45_675 ();
 sg13g2_decap_4 FILLER_45_686 ();
 sg13g2_decap_8 FILLER_45_698 ();
 sg13g2_decap_8 FILLER_45_705 ();
 sg13g2_fill_2 FILLER_45_712 ();
 sg13g2_fill_1 FILLER_45_714 ();
 sg13g2_decap_8 FILLER_45_719 ();
 sg13g2_decap_8 FILLER_45_726 ();
 sg13g2_decap_8 FILLER_45_733 ();
 sg13g2_decap_8 FILLER_45_740 ();
 sg13g2_decap_4 FILLER_45_747 ();
 sg13g2_decap_4 FILLER_45_755 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_774 ();
 sg13g2_decap_8 FILLER_45_793 ();
 sg13g2_decap_8 FILLER_45_800 ();
 sg13g2_decap_8 FILLER_45_811 ();
 sg13g2_decap_8 FILLER_45_818 ();
 sg13g2_decap_4 FILLER_45_830 ();
 sg13g2_fill_1 FILLER_45_834 ();
 sg13g2_decap_4 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_45_897 ();
 sg13g2_fill_1 FILLER_45_904 ();
 sg13g2_decap_8 FILLER_45_913 ();
 sg13g2_decap_8 FILLER_45_920 ();
 sg13g2_decap_8 FILLER_45_927 ();
 sg13g2_fill_1 FILLER_45_934 ();
 sg13g2_decap_8 FILLER_45_943 ();
 sg13g2_fill_1 FILLER_45_950 ();
 sg13g2_decap_8 FILLER_45_966 ();
 sg13g2_decap_4 FILLER_45_973 ();
 sg13g2_decap_8 FILLER_45_994 ();
 sg13g2_decap_8 FILLER_45_1001 ();
 sg13g2_decap_8 FILLER_45_1008 ();
 sg13g2_decap_8 FILLER_45_1015 ();
 sg13g2_decap_8 FILLER_45_1022 ();
 sg13g2_decap_4 FILLER_45_1029 ();
 sg13g2_fill_1 FILLER_45_1033 ();
 sg13g2_fill_1 FILLER_45_1037 ();
 sg13g2_decap_8 FILLER_45_1042 ();
 sg13g2_decap_8 FILLER_45_1049 ();
 sg13g2_decap_8 FILLER_45_1056 ();
 sg13g2_decap_8 FILLER_45_1063 ();
 sg13g2_decap_8 FILLER_45_1070 ();
 sg13g2_fill_1 FILLER_45_1077 ();
 sg13g2_fill_2 FILLER_45_1099 ();
 sg13g2_fill_1 FILLER_45_1101 ();
 sg13g2_fill_2 FILLER_45_1111 ();
 sg13g2_fill_1 FILLER_45_1113 ();
 sg13g2_decap_8 FILLER_45_1140 ();
 sg13g2_decap_4 FILLER_45_1147 ();
 sg13g2_decap_4 FILLER_45_1156 ();
 sg13g2_decap_8 FILLER_45_1164 ();
 sg13g2_decap_8 FILLER_45_1171 ();
 sg13g2_decap_8 FILLER_45_1178 ();
 sg13g2_fill_1 FILLER_45_1185 ();
 sg13g2_decap_4 FILLER_45_1205 ();
 sg13g2_fill_1 FILLER_45_1209 ();
 sg13g2_decap_8 FILLER_45_1219 ();
 sg13g2_decap_8 FILLER_45_1226 ();
 sg13g2_fill_2 FILLER_45_1233 ();
 sg13g2_fill_1 FILLER_45_1235 ();
 sg13g2_decap_8 FILLER_45_1266 ();
 sg13g2_fill_1 FILLER_45_1273 ();
 sg13g2_decap_4 FILLER_45_1282 ();
 sg13g2_fill_2 FILLER_45_1286 ();
 sg13g2_decap_8 FILLER_45_1292 ();
 sg13g2_decap_8 FILLER_45_1299 ();
 sg13g2_fill_1 FILLER_45_1306 ();
 sg13g2_decap_4 FILLER_45_1315 ();
 sg13g2_fill_1 FILLER_45_1319 ();
 sg13g2_decap_8 FILLER_45_1331 ();
 sg13g2_decap_8 FILLER_45_1338 ();
 sg13g2_decap_4 FILLER_45_1345 ();
 sg13g2_fill_2 FILLER_45_1349 ();
 sg13g2_fill_2 FILLER_45_1355 ();
 sg13g2_fill_1 FILLER_45_1357 ();
 sg13g2_decap_8 FILLER_45_1362 ();
 sg13g2_decap_8 FILLER_45_1369 ();
 sg13g2_decap_4 FILLER_45_1376 ();
 sg13g2_fill_1 FILLER_45_1380 ();
 sg13g2_decap_4 FILLER_45_1386 ();
 sg13g2_fill_1 FILLER_45_1390 ();
 sg13g2_fill_2 FILLER_45_1417 ();
 sg13g2_fill_1 FILLER_45_1419 ();
 sg13g2_decap_8 FILLER_45_1423 ();
 sg13g2_fill_2 FILLER_45_1430 ();
 sg13g2_fill_1 FILLER_45_1432 ();
 sg13g2_decap_4 FILLER_45_1437 ();
 sg13g2_fill_2 FILLER_45_1441 ();
 sg13g2_decap_8 FILLER_45_1450 ();
 sg13g2_decap_8 FILLER_45_1457 ();
 sg13g2_decap_4 FILLER_45_1464 ();
 sg13g2_decap_8 FILLER_45_1473 ();
 sg13g2_decap_8 FILLER_45_1480 ();
 sg13g2_decap_8 FILLER_45_1487 ();
 sg13g2_decap_8 FILLER_45_1494 ();
 sg13g2_decap_8 FILLER_45_1501 ();
 sg13g2_decap_8 FILLER_45_1508 ();
 sg13g2_decap_8 FILLER_45_1515 ();
 sg13g2_decap_8 FILLER_45_1522 ();
 sg13g2_fill_1 FILLER_45_1529 ();
 sg13g2_decap_8 FILLER_45_1535 ();
 sg13g2_decap_8 FILLER_45_1542 ();
 sg13g2_decap_8 FILLER_45_1549 ();
 sg13g2_fill_1 FILLER_45_1556 ();
 sg13g2_decap_4 FILLER_45_1563 ();
 sg13g2_fill_1 FILLER_45_1567 ();
 sg13g2_decap_8 FILLER_45_1572 ();
 sg13g2_decap_8 FILLER_45_1579 ();
 sg13g2_decap_4 FILLER_45_1586 ();
 sg13g2_fill_1 FILLER_45_1590 ();
 sg13g2_fill_1 FILLER_45_1600 ();
 sg13g2_fill_2 FILLER_45_1606 ();
 sg13g2_fill_1 FILLER_45_1608 ();
 sg13g2_fill_2 FILLER_45_1618 ();
 sg13g2_fill_1 FILLER_45_1620 ();
 sg13g2_decap_4 FILLER_45_1653 ();
 sg13g2_fill_1 FILLER_45_1657 ();
 sg13g2_decap_8 FILLER_45_1662 ();
 sg13g2_decap_4 FILLER_45_1669 ();
 sg13g2_decap_8 FILLER_45_1706 ();
 sg13g2_decap_8 FILLER_45_1713 ();
 sg13g2_decap_4 FILLER_45_1720 ();
 sg13g2_decap_8 FILLER_45_1729 ();
 sg13g2_decap_8 FILLER_45_1766 ();
 sg13g2_fill_1 FILLER_45_1773 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_fill_2 FILLER_46_28 ();
 sg13g2_fill_1 FILLER_46_30 ();
 sg13g2_decap_4 FILLER_46_52 ();
 sg13g2_fill_2 FILLER_46_56 ();
 sg13g2_decap_4 FILLER_46_76 ();
 sg13g2_fill_2 FILLER_46_84 ();
 sg13g2_fill_1 FILLER_46_86 ();
 sg13g2_fill_2 FILLER_46_97 ();
 sg13g2_fill_2 FILLER_46_103 ();
 sg13g2_fill_1 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_115 ();
 sg13g2_decap_8 FILLER_46_122 ();
 sg13g2_fill_1 FILLER_46_129 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_fill_2 FILLER_46_147 ();
 sg13g2_decap_4 FILLER_46_158 ();
 sg13g2_fill_1 FILLER_46_162 ();
 sg13g2_decap_8 FILLER_46_174 ();
 sg13g2_decap_4 FILLER_46_181 ();
 sg13g2_fill_1 FILLER_46_185 ();
 sg13g2_fill_2 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_204 ();
 sg13g2_fill_1 FILLER_46_206 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_228 ();
 sg13g2_fill_2 FILLER_46_235 ();
 sg13g2_fill_1 FILLER_46_237 ();
 sg13g2_decap_4 FILLER_46_242 ();
 sg13g2_fill_2 FILLER_46_256 ();
 sg13g2_fill_1 FILLER_46_258 ();
 sg13g2_decap_8 FILLER_46_264 ();
 sg13g2_decap_8 FILLER_46_271 ();
 sg13g2_decap_4 FILLER_46_278 ();
 sg13g2_decap_8 FILLER_46_302 ();
 sg13g2_decap_8 FILLER_46_309 ();
 sg13g2_decap_8 FILLER_46_316 ();
 sg13g2_decap_8 FILLER_46_323 ();
 sg13g2_decap_8 FILLER_46_330 ();
 sg13g2_fill_2 FILLER_46_337 ();
 sg13g2_decap_8 FILLER_46_347 ();
 sg13g2_decap_4 FILLER_46_354 ();
 sg13g2_fill_1 FILLER_46_358 ();
 sg13g2_decap_8 FILLER_46_370 ();
 sg13g2_decap_8 FILLER_46_377 ();
 sg13g2_decap_8 FILLER_46_384 ();
 sg13g2_fill_1 FILLER_46_391 ();
 sg13g2_fill_1 FILLER_46_398 ();
 sg13g2_decap_8 FILLER_46_404 ();
 sg13g2_fill_2 FILLER_46_411 ();
 sg13g2_fill_1 FILLER_46_413 ();
 sg13g2_fill_1 FILLER_46_432 ();
 sg13g2_decap_4 FILLER_46_438 ();
 sg13g2_fill_1 FILLER_46_442 ();
 sg13g2_decap_4 FILLER_46_450 ();
 sg13g2_fill_1 FILLER_46_454 ();
 sg13g2_fill_1 FILLER_46_460 ();
 sg13g2_decap_8 FILLER_46_466 ();
 sg13g2_decap_8 FILLER_46_473 ();
 sg13g2_decap_8 FILLER_46_480 ();
 sg13g2_decap_8 FILLER_46_487 ();
 sg13g2_fill_2 FILLER_46_494 ();
 sg13g2_fill_1 FILLER_46_496 ();
 sg13g2_decap_8 FILLER_46_501 ();
 sg13g2_fill_2 FILLER_46_508 ();
 sg13g2_decap_8 FILLER_46_519 ();
 sg13g2_decap_8 FILLER_46_526 ();
 sg13g2_decap_4 FILLER_46_533 ();
 sg13g2_fill_2 FILLER_46_537 ();
 sg13g2_decap_8 FILLER_46_544 ();
 sg13g2_decap_8 FILLER_46_551 ();
 sg13g2_decap_8 FILLER_46_558 ();
 sg13g2_fill_2 FILLER_46_565 ();
 sg13g2_fill_1 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_572 ();
 sg13g2_decap_8 FILLER_46_579 ();
 sg13g2_decap_4 FILLER_46_586 ();
 sg13g2_fill_1 FILLER_46_590 ();
 sg13g2_decap_8 FILLER_46_597 ();
 sg13g2_decap_8 FILLER_46_604 ();
 sg13g2_decap_8 FILLER_46_611 ();
 sg13g2_decap_8 FILLER_46_618 ();
 sg13g2_decap_8 FILLER_46_625 ();
 sg13g2_fill_2 FILLER_46_632 ();
 sg13g2_fill_1 FILLER_46_634 ();
 sg13g2_decap_8 FILLER_46_674 ();
 sg13g2_fill_2 FILLER_46_681 ();
 sg13g2_fill_1 FILLER_46_683 ();
 sg13g2_decap_8 FILLER_46_692 ();
 sg13g2_decap_4 FILLER_46_699 ();
 sg13g2_fill_2 FILLER_46_706 ();
 sg13g2_fill_1 FILLER_46_708 ();
 sg13g2_decap_4 FILLER_46_739 ();
 sg13g2_fill_1 FILLER_46_743 ();
 sg13g2_decap_4 FILLER_46_749 ();
 sg13g2_fill_1 FILLER_46_753 ();
 sg13g2_decap_8 FILLER_46_758 ();
 sg13g2_decap_8 FILLER_46_765 ();
 sg13g2_decap_8 FILLER_46_772 ();
 sg13g2_decap_8 FILLER_46_779 ();
 sg13g2_decap_8 FILLER_46_796 ();
 sg13g2_fill_2 FILLER_46_803 ();
 sg13g2_fill_1 FILLER_46_805 ();
 sg13g2_decap_4 FILLER_46_810 ();
 sg13g2_decap_8 FILLER_46_818 ();
 sg13g2_fill_1 FILLER_46_825 ();
 sg13g2_decap_4 FILLER_46_830 ();
 sg13g2_fill_1 FILLER_46_834 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_decap_8 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_46_871 ();
 sg13g2_decap_8 FILLER_46_878 ();
 sg13g2_fill_2 FILLER_46_885 ();
 sg13g2_decap_8 FILLER_46_891 ();
 sg13g2_decap_8 FILLER_46_898 ();
 sg13g2_decap_8 FILLER_46_905 ();
 sg13g2_decap_8 FILLER_46_912 ();
 sg13g2_decap_8 FILLER_46_919 ();
 sg13g2_decap_8 FILLER_46_926 ();
 sg13g2_decap_4 FILLER_46_933 ();
 sg13g2_fill_2 FILLER_46_937 ();
 sg13g2_decap_8 FILLER_46_944 ();
 sg13g2_decap_8 FILLER_46_951 ();
 sg13g2_fill_2 FILLER_46_958 ();
 sg13g2_fill_1 FILLER_46_960 ();
 sg13g2_decap_4 FILLER_46_965 ();
 sg13g2_fill_1 FILLER_46_969 ();
 sg13g2_decap_4 FILLER_46_975 ();
 sg13g2_fill_2 FILLER_46_979 ();
 sg13g2_fill_2 FILLER_46_989 ();
 sg13g2_fill_1 FILLER_46_991 ();
 sg13g2_decap_8 FILLER_46_995 ();
 sg13g2_decap_4 FILLER_46_1032 ();
 sg13g2_decap_4 FILLER_46_1045 ();
 sg13g2_decap_8 FILLER_46_1075 ();
 sg13g2_fill_2 FILLER_46_1082 ();
 sg13g2_fill_2 FILLER_46_1094 ();
 sg13g2_decap_8 FILLER_46_1109 ();
 sg13g2_decap_4 FILLER_46_1116 ();
 sg13g2_decap_8 FILLER_46_1124 ();
 sg13g2_decap_8 FILLER_46_1131 ();
 sg13g2_decap_8 FILLER_46_1138 ();
 sg13g2_decap_8 FILLER_46_1145 ();
 sg13g2_fill_2 FILLER_46_1152 ();
 sg13g2_decap_8 FILLER_46_1180 ();
 sg13g2_decap_8 FILLER_46_1187 ();
 sg13g2_fill_2 FILLER_46_1194 ();
 sg13g2_decap_4 FILLER_46_1205 ();
 sg13g2_fill_1 FILLER_46_1209 ();
 sg13g2_decap_8 FILLER_46_1214 ();
 sg13g2_decap_4 FILLER_46_1221 ();
 sg13g2_fill_1 FILLER_46_1225 ();
 sg13g2_fill_2 FILLER_46_1234 ();
 sg13g2_decap_8 FILLER_46_1241 ();
 sg13g2_decap_8 FILLER_46_1248 ();
 sg13g2_fill_2 FILLER_46_1255 ();
 sg13g2_fill_1 FILLER_46_1257 ();
 sg13g2_decap_8 FILLER_46_1262 ();
 sg13g2_decap_4 FILLER_46_1269 ();
 sg13g2_fill_2 FILLER_46_1273 ();
 sg13g2_decap_8 FILLER_46_1283 ();
 sg13g2_decap_8 FILLER_46_1290 ();
 sg13g2_decap_8 FILLER_46_1297 ();
 sg13g2_decap_8 FILLER_46_1304 ();
 sg13g2_decap_8 FILLER_46_1311 ();
 sg13g2_decap_8 FILLER_46_1318 ();
 sg13g2_fill_1 FILLER_46_1325 ();
 sg13g2_decap_8 FILLER_46_1334 ();
 sg13g2_decap_4 FILLER_46_1345 ();
 sg13g2_decap_8 FILLER_46_1357 ();
 sg13g2_decap_4 FILLER_46_1364 ();
 sg13g2_fill_1 FILLER_46_1368 ();
 sg13g2_decap_8 FILLER_46_1384 ();
 sg13g2_decap_8 FILLER_46_1391 ();
 sg13g2_decap_4 FILLER_46_1398 ();
 sg13g2_fill_1 FILLER_46_1402 ();
 sg13g2_fill_2 FILLER_46_1429 ();
 sg13g2_fill_1 FILLER_46_1431 ();
 sg13g2_decap_8 FILLER_46_1435 ();
 sg13g2_decap_4 FILLER_46_1442 ();
 sg13g2_fill_2 FILLER_46_1446 ();
 sg13g2_decap_8 FILLER_46_1474 ();
 sg13g2_decap_8 FILLER_46_1481 ();
 sg13g2_fill_2 FILLER_46_1488 ();
 sg13g2_decap_8 FILLER_46_1494 ();
 sg13g2_decap_8 FILLER_46_1501 ();
 sg13g2_decap_8 FILLER_46_1508 ();
 sg13g2_decap_8 FILLER_46_1515 ();
 sg13g2_fill_2 FILLER_46_1528 ();
 sg13g2_decap_8 FILLER_46_1561 ();
 sg13g2_decap_8 FILLER_46_1568 ();
 sg13g2_decap_8 FILLER_46_1575 ();
 sg13g2_decap_8 FILLER_46_1582 ();
 sg13g2_fill_2 FILLER_46_1589 ();
 sg13g2_fill_1 FILLER_46_1591 ();
 sg13g2_decap_8 FILLER_46_1605 ();
 sg13g2_decap_8 FILLER_46_1612 ();
 sg13g2_decap_8 FILLER_46_1619 ();
 sg13g2_fill_2 FILLER_46_1626 ();
 sg13g2_fill_2 FILLER_46_1632 ();
 sg13g2_fill_1 FILLER_46_1634 ();
 sg13g2_decap_8 FILLER_46_1645 ();
 sg13g2_decap_4 FILLER_46_1652 ();
 sg13g2_fill_1 FILLER_46_1656 ();
 sg13g2_decap_8 FILLER_46_1663 ();
 sg13g2_fill_1 FILLER_46_1670 ();
 sg13g2_decap_4 FILLER_46_1677 ();
 sg13g2_fill_2 FILLER_46_1681 ();
 sg13g2_decap_8 FILLER_46_1687 ();
 sg13g2_decap_8 FILLER_46_1694 ();
 sg13g2_fill_1 FILLER_46_1701 ();
 sg13g2_fill_2 FILLER_46_1708 ();
 sg13g2_decap_4 FILLER_46_1713 ();
 sg13g2_fill_2 FILLER_46_1717 ();
 sg13g2_decap_4 FILLER_46_1731 ();
 sg13g2_fill_2 FILLER_46_1739 ();
 sg13g2_fill_1 FILLER_46_1741 ();
 sg13g2_decap_8 FILLER_46_1746 ();
 sg13g2_decap_8 FILLER_46_1753 ();
 sg13g2_decap_8 FILLER_46_1760 ();
 sg13g2_decap_8 FILLER_46_1767 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_4 FILLER_47_28 ();
 sg13g2_fill_2 FILLER_47_32 ();
 sg13g2_fill_1 FILLER_47_43 ();
 sg13g2_decap_4 FILLER_47_48 ();
 sg13g2_fill_2 FILLER_47_75 ();
 sg13g2_fill_1 FILLER_47_77 ();
 sg13g2_fill_2 FILLER_47_92 ();
 sg13g2_fill_1 FILLER_47_94 ();
 sg13g2_fill_2 FILLER_47_106 ();
 sg13g2_fill_1 FILLER_47_108 ();
 sg13g2_decap_8 FILLER_47_113 ();
 sg13g2_decap_8 FILLER_47_120 ();
 sg13g2_fill_2 FILLER_47_127 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_4 FILLER_47_147 ();
 sg13g2_fill_2 FILLER_47_151 ();
 sg13g2_decap_8 FILLER_47_163 ();
 sg13g2_decap_8 FILLER_47_178 ();
 sg13g2_decap_8 FILLER_47_185 ();
 sg13g2_decap_8 FILLER_47_192 ();
 sg13g2_fill_1 FILLER_47_199 ();
 sg13g2_decap_4 FILLER_47_205 ();
 sg13g2_fill_1 FILLER_47_209 ();
 sg13g2_fill_2 FILLER_47_218 ();
 sg13g2_fill_1 FILLER_47_220 ();
 sg13g2_fill_2 FILLER_47_225 ();
 sg13g2_fill_1 FILLER_47_227 ();
 sg13g2_fill_1 FILLER_47_239 ();
 sg13g2_decap_4 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_255 ();
 sg13g2_decap_4 FILLER_47_262 ();
 sg13g2_fill_1 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_277 ();
 sg13g2_decap_4 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_288 ();
 sg13g2_fill_2 FILLER_47_294 ();
 sg13g2_fill_1 FILLER_47_296 ();
 sg13g2_fill_2 FILLER_47_305 ();
 sg13g2_fill_1 FILLER_47_307 ();
 sg13g2_fill_2 FILLER_47_318 ();
 sg13g2_fill_1 FILLER_47_320 ();
 sg13g2_decap_8 FILLER_47_326 ();
 sg13g2_decap_4 FILLER_47_333 ();
 sg13g2_fill_2 FILLER_47_337 ();
 sg13g2_decap_8 FILLER_47_344 ();
 sg13g2_fill_2 FILLER_47_351 ();
 sg13g2_decap_8 FILLER_47_367 ();
 sg13g2_decap_8 FILLER_47_374 ();
 sg13g2_decap_4 FILLER_47_381 ();
 sg13g2_decap_4 FILLER_47_389 ();
 sg13g2_fill_2 FILLER_47_403 ();
 sg13g2_decap_8 FILLER_47_425 ();
 sg13g2_decap_4 FILLER_47_432 ();
 sg13g2_fill_2 FILLER_47_436 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_fill_2 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_517 ();
 sg13g2_fill_2 FILLER_47_524 ();
 sg13g2_fill_1 FILLER_47_564 ();
 sg13g2_decap_4 FILLER_47_591 ();
 sg13g2_fill_2 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_633 ();
 sg13g2_fill_2 FILLER_47_640 ();
 sg13g2_fill_1 FILLER_47_642 ();
 sg13g2_decap_8 FILLER_47_648 ();
 sg13g2_decap_8 FILLER_47_655 ();
 sg13g2_decap_8 FILLER_47_662 ();
 sg13g2_decap_8 FILLER_47_669 ();
 sg13g2_decap_8 FILLER_47_676 ();
 sg13g2_decap_8 FILLER_47_683 ();
 sg13g2_fill_2 FILLER_47_690 ();
 sg13g2_fill_1 FILLER_47_692 ();
 sg13g2_fill_2 FILLER_47_702 ();
 sg13g2_decap_8 FILLER_47_709 ();
 sg13g2_decap_8 FILLER_47_716 ();
 sg13g2_decap_8 FILLER_47_723 ();
 sg13g2_decap_8 FILLER_47_730 ();
 sg13g2_decap_8 FILLER_47_737 ();
 sg13g2_fill_1 FILLER_47_744 ();
 sg13g2_decap_8 FILLER_47_771 ();
 sg13g2_decap_8 FILLER_47_778 ();
 sg13g2_decap_8 FILLER_47_785 ();
 sg13g2_decap_4 FILLER_47_792 ();
 sg13g2_fill_2 FILLER_47_796 ();
 sg13g2_decap_8 FILLER_47_811 ();
 sg13g2_decap_8 FILLER_47_818 ();
 sg13g2_decap_8 FILLER_47_825 ();
 sg13g2_decap_4 FILLER_47_832 ();
 sg13g2_fill_2 FILLER_47_866 ();
 sg13g2_decap_4 FILLER_47_886 ();
 sg13g2_decap_8 FILLER_47_898 ();
 sg13g2_decap_4 FILLER_47_905 ();
 sg13g2_decap_8 FILLER_47_913 ();
 sg13g2_fill_2 FILLER_47_920 ();
 sg13g2_decap_8 FILLER_47_927 ();
 sg13g2_decap_4 FILLER_47_934 ();
 sg13g2_decap_8 FILLER_47_964 ();
 sg13g2_decap_8 FILLER_47_975 ();
 sg13g2_decap_8 FILLER_47_982 ();
 sg13g2_fill_2 FILLER_47_989 ();
 sg13g2_decap_8 FILLER_47_996 ();
 sg13g2_decap_8 FILLER_47_1003 ();
 sg13g2_decap_8 FILLER_47_1014 ();
 sg13g2_decap_8 FILLER_47_1021 ();
 sg13g2_decap_8 FILLER_47_1028 ();
 sg13g2_fill_2 FILLER_47_1035 ();
 sg13g2_fill_1 FILLER_47_1037 ();
 sg13g2_decap_8 FILLER_47_1047 ();
 sg13g2_decap_8 FILLER_47_1058 ();
 sg13g2_decap_8 FILLER_47_1065 ();
 sg13g2_decap_8 FILLER_47_1072 ();
 sg13g2_fill_1 FILLER_47_1079 ();
 sg13g2_fill_2 FILLER_47_1089 ();
 sg13g2_decap_8 FILLER_47_1125 ();
 sg13g2_decap_8 FILLER_47_1132 ();
 sg13g2_decap_8 FILLER_47_1139 ();
 sg13g2_fill_2 FILLER_47_1146 ();
 sg13g2_decap_4 FILLER_47_1158 ();
 sg13g2_fill_2 FILLER_47_1162 ();
 sg13g2_decap_8 FILLER_47_1168 ();
 sg13g2_decap_8 FILLER_47_1175 ();
 sg13g2_decap_8 FILLER_47_1182 ();
 sg13g2_decap_8 FILLER_47_1189 ();
 sg13g2_decap_8 FILLER_47_1196 ();
 sg13g2_decap_8 FILLER_47_1203 ();
 sg13g2_decap_8 FILLER_47_1210 ();
 sg13g2_decap_8 FILLER_47_1217 ();
 sg13g2_fill_2 FILLER_47_1240 ();
 sg13g2_decap_8 FILLER_47_1247 ();
 sg13g2_decap_8 FILLER_47_1254 ();
 sg13g2_fill_2 FILLER_47_1261 ();
 sg13g2_fill_1 FILLER_47_1263 ();
 sg13g2_decap_8 FILLER_47_1279 ();
 sg13g2_decap_8 FILLER_47_1286 ();
 sg13g2_decap_4 FILLER_47_1293 ();
 sg13g2_fill_2 FILLER_47_1297 ();
 sg13g2_fill_2 FILLER_47_1325 ();
 sg13g2_decap_4 FILLER_47_1336 ();
 sg13g2_fill_1 FILLER_47_1340 ();
 sg13g2_fill_2 FILLER_47_1346 ();
 sg13g2_fill_1 FILLER_47_1360 ();
 sg13g2_fill_1 FILLER_47_1365 ();
 sg13g2_decap_8 FILLER_47_1382 ();
 sg13g2_decap_8 FILLER_47_1389 ();
 sg13g2_decap_8 FILLER_47_1396 ();
 sg13g2_decap_4 FILLER_47_1403 ();
 sg13g2_decap_8 FILLER_47_1411 ();
 sg13g2_decap_8 FILLER_47_1418 ();
 sg13g2_decap_4 FILLER_47_1437 ();
 sg13g2_fill_2 FILLER_47_1441 ();
 sg13g2_decap_4 FILLER_47_1449 ();
 sg13g2_fill_1 FILLER_47_1453 ();
 sg13g2_decap_8 FILLER_47_1458 ();
 sg13g2_decap_8 FILLER_47_1465 ();
 sg13g2_fill_2 FILLER_47_1472 ();
 sg13g2_decap_8 FILLER_47_1509 ();
 sg13g2_fill_1 FILLER_47_1516 ();
 sg13g2_fill_2 FILLER_47_1529 ();
 sg13g2_fill_1 FILLER_47_1531 ();
 sg13g2_decap_8 FILLER_47_1561 ();
 sg13g2_decap_4 FILLER_47_1568 ();
 sg13g2_fill_1 FILLER_47_1572 ();
 sg13g2_decap_4 FILLER_47_1577 ();
 sg13g2_fill_1 FILLER_47_1581 ();
 sg13g2_fill_2 FILLER_47_1585 ();
 sg13g2_fill_1 FILLER_47_1587 ();
 sg13g2_decap_8 FILLER_47_1614 ();
 sg13g2_decap_8 FILLER_47_1621 ();
 sg13g2_decap_8 FILLER_47_1628 ();
 sg13g2_decap_4 FILLER_47_1635 ();
 sg13g2_fill_2 FILLER_47_1639 ();
 sg13g2_decap_8 FILLER_47_1645 ();
 sg13g2_decap_4 FILLER_47_1652 ();
 sg13g2_decap_8 FILLER_47_1669 ();
 sg13g2_decap_8 FILLER_47_1676 ();
 sg13g2_decap_4 FILLER_47_1683 ();
 sg13g2_fill_1 FILLER_47_1687 ();
 sg13g2_decap_8 FILLER_47_1692 ();
 sg13g2_decap_8 FILLER_47_1699 ();
 sg13g2_decap_8 FILLER_47_1706 ();
 sg13g2_decap_4 FILLER_47_1713 ();
 sg13g2_fill_2 FILLER_47_1717 ();
 sg13g2_decap_4 FILLER_47_1722 ();
 sg13g2_fill_1 FILLER_47_1733 ();
 sg13g2_fill_1 FILLER_47_1741 ();
 sg13g2_fill_1 FILLER_47_1752 ();
 sg13g2_decap_8 FILLER_47_1758 ();
 sg13g2_decap_8 FILLER_47_1765 ();
 sg13g2_fill_2 FILLER_47_1772 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_fill_1 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_37 ();
 sg13g2_decap_4 FILLER_48_44 ();
 sg13g2_fill_2 FILLER_48_48 ();
 sg13g2_decap_4 FILLER_48_60 ();
 sg13g2_decap_8 FILLER_48_73 ();
 sg13g2_fill_1 FILLER_48_80 ();
 sg13g2_decap_4 FILLER_48_86 ();
 sg13g2_fill_2 FILLER_48_90 ();
 sg13g2_fill_2 FILLER_48_97 ();
 sg13g2_decap_8 FILLER_48_109 ();
 sg13g2_decap_8 FILLER_48_124 ();
 sg13g2_fill_2 FILLER_48_131 ();
 sg13g2_fill_1 FILLER_48_133 ();
 sg13g2_fill_2 FILLER_48_139 ();
 sg13g2_fill_1 FILLER_48_141 ();
 sg13g2_decap_8 FILLER_48_152 ();
 sg13g2_decap_8 FILLER_48_159 ();
 sg13g2_decap_8 FILLER_48_180 ();
 sg13g2_fill_1 FILLER_48_192 ();
 sg13g2_decap_8 FILLER_48_198 ();
 sg13g2_decap_4 FILLER_48_205 ();
 sg13g2_decap_8 FILLER_48_223 ();
 sg13g2_decap_8 FILLER_48_230 ();
 sg13g2_decap_8 FILLER_48_246 ();
 sg13g2_decap_4 FILLER_48_253 ();
 sg13g2_fill_2 FILLER_48_257 ();
 sg13g2_fill_2 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_273 ();
 sg13g2_fill_1 FILLER_48_279 ();
 sg13g2_fill_2 FILLER_48_285 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_decap_8 FILLER_48_298 ();
 sg13g2_fill_2 FILLER_48_305 ();
 sg13g2_fill_1 FILLER_48_307 ();
 sg13g2_decap_4 FILLER_48_326 ();
 sg13g2_decap_8 FILLER_48_352 ();
 sg13g2_decap_8 FILLER_48_373 ();
 sg13g2_decap_8 FILLER_48_380 ();
 sg13g2_fill_1 FILLER_48_387 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_4 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_403 ();
 sg13g2_decap_4 FILLER_48_410 ();
 sg13g2_fill_2 FILLER_48_414 ();
 sg13g2_decap_4 FILLER_48_424 ();
 sg13g2_fill_1 FILLER_48_428 ();
 sg13g2_decap_4 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_454 ();
 sg13g2_decap_8 FILLER_48_461 ();
 sg13g2_decap_8 FILLER_48_468 ();
 sg13g2_decap_8 FILLER_48_479 ();
 sg13g2_decap_8 FILLER_48_486 ();
 sg13g2_decap_8 FILLER_48_493 ();
 sg13g2_decap_8 FILLER_48_500 ();
 sg13g2_decap_8 FILLER_48_507 ();
 sg13g2_decap_8 FILLER_48_514 ();
 sg13g2_decap_4 FILLER_48_521 ();
 sg13g2_decap_8 FILLER_48_530 ();
 sg13g2_decap_8 FILLER_48_541 ();
 sg13g2_decap_8 FILLER_48_548 ();
 sg13g2_decap_8 FILLER_48_555 ();
 sg13g2_decap_8 FILLER_48_562 ();
 sg13g2_fill_1 FILLER_48_569 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_4 FILLER_48_609 ();
 sg13g2_fill_1 FILLER_48_613 ();
 sg13g2_decap_8 FILLER_48_618 ();
 sg13g2_decap_8 FILLER_48_625 ();
 sg13g2_decap_8 FILLER_48_632 ();
 sg13g2_fill_2 FILLER_48_639 ();
 sg13g2_decap_8 FILLER_48_667 ();
 sg13g2_fill_1 FILLER_48_674 ();
 sg13g2_fill_2 FILLER_48_680 ();
 sg13g2_fill_1 FILLER_48_682 ();
 sg13g2_fill_2 FILLER_48_687 ();
 sg13g2_fill_1 FILLER_48_689 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_4 FILLER_48_700 ();
 sg13g2_fill_2 FILLER_48_704 ();
 sg13g2_decap_4 FILLER_48_710 ();
 sg13g2_decap_8 FILLER_48_718 ();
 sg13g2_decap_8 FILLER_48_725 ();
 sg13g2_decap_4 FILLER_48_732 ();
 sg13g2_fill_2 FILLER_48_736 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_786 ();
 sg13g2_decap_8 FILLER_48_793 ();
 sg13g2_fill_2 FILLER_48_800 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_4 FILLER_48_847 ();
 sg13g2_fill_1 FILLER_48_851 ();
 sg13g2_decap_8 FILLER_48_856 ();
 sg13g2_decap_8 FILLER_48_863 ();
 sg13g2_decap_8 FILLER_48_870 ();
 sg13g2_decap_8 FILLER_48_877 ();
 sg13g2_decap_4 FILLER_48_884 ();
 sg13g2_fill_2 FILLER_48_888 ();
 sg13g2_fill_1 FILLER_48_894 ();
 sg13g2_fill_2 FILLER_48_900 ();
 sg13g2_decap_4 FILLER_48_928 ();
 sg13g2_fill_1 FILLER_48_932 ();
 sg13g2_decap_8 FILLER_48_938 ();
 sg13g2_decap_8 FILLER_48_949 ();
 sg13g2_decap_8 FILLER_48_956 ();
 sg13g2_decap_8 FILLER_48_963 ();
 sg13g2_decap_8 FILLER_48_970 ();
 sg13g2_decap_8 FILLER_48_977 ();
 sg13g2_decap_4 FILLER_48_984 ();
 sg13g2_fill_1 FILLER_48_988 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_4 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1009 ();
 sg13g2_decap_8 FILLER_48_1016 ();
 sg13g2_decap_8 FILLER_48_1023 ();
 sg13g2_decap_8 FILLER_48_1030 ();
 sg13g2_fill_1 FILLER_48_1037 ();
 sg13g2_fill_1 FILLER_48_1090 ();
 sg13g2_fill_2 FILLER_48_1096 ();
 sg13g2_fill_1 FILLER_48_1098 ();
 sg13g2_fill_2 FILLER_48_1108 ();
 sg13g2_fill_1 FILLER_48_1110 ();
 sg13g2_decap_8 FILLER_48_1137 ();
 sg13g2_decap_8 FILLER_48_1144 ();
 sg13g2_fill_1 FILLER_48_1151 ();
 sg13g2_decap_8 FILLER_48_1182 ();
 sg13g2_fill_2 FILLER_48_1189 ();
 sg13g2_decap_4 FILLER_48_1195 ();
 sg13g2_fill_1 FILLER_48_1199 ();
 sg13g2_decap_8 FILLER_48_1204 ();
 sg13g2_decap_8 FILLER_48_1211 ();
 sg13g2_decap_8 FILLER_48_1218 ();
 sg13g2_decap_4 FILLER_48_1242 ();
 sg13g2_fill_1 FILLER_48_1246 ();
 sg13g2_decap_8 FILLER_48_1251 ();
 sg13g2_decap_4 FILLER_48_1258 ();
 sg13g2_fill_1 FILLER_48_1262 ();
 sg13g2_decap_8 FILLER_48_1266 ();
 sg13g2_fill_2 FILLER_48_1277 ();
 sg13g2_fill_1 FILLER_48_1283 ();
 sg13g2_decap_8 FILLER_48_1289 ();
 sg13g2_decap_8 FILLER_48_1296 ();
 sg13g2_decap_8 FILLER_48_1307 ();
 sg13g2_decap_8 FILLER_48_1314 ();
 sg13g2_decap_8 FILLER_48_1321 ();
 sg13g2_fill_1 FILLER_48_1328 ();
 sg13g2_decap_8 FILLER_48_1332 ();
 sg13g2_decap_4 FILLER_48_1339 ();
 sg13g2_fill_1 FILLER_48_1343 ();
 sg13g2_decap_8 FILLER_48_1349 ();
 sg13g2_decap_8 FILLER_48_1356 ();
 sg13g2_decap_8 FILLER_48_1363 ();
 sg13g2_fill_1 FILLER_48_1370 ();
 sg13g2_decap_8 FILLER_48_1375 ();
 sg13g2_decap_8 FILLER_48_1382 ();
 sg13g2_decap_8 FILLER_48_1389 ();
 sg13g2_decap_4 FILLER_48_1396 ();
 sg13g2_fill_1 FILLER_48_1400 ();
 sg13g2_decap_8 FILLER_48_1405 ();
 sg13g2_decap_8 FILLER_48_1412 ();
 sg13g2_fill_2 FILLER_48_1419 ();
 sg13g2_decap_8 FILLER_48_1434 ();
 sg13g2_fill_2 FILLER_48_1441 ();
 sg13g2_fill_1 FILLER_48_1443 ();
 sg13g2_decap_8 FILLER_48_1448 ();
 sg13g2_decap_4 FILLER_48_1455 ();
 sg13g2_decap_8 FILLER_48_1464 ();
 sg13g2_decap_8 FILLER_48_1471 ();
 sg13g2_decap_8 FILLER_48_1478 ();
 sg13g2_decap_8 FILLER_48_1512 ();
 sg13g2_decap_4 FILLER_48_1519 ();
 sg13g2_fill_2 FILLER_48_1523 ();
 sg13g2_fill_2 FILLER_48_1542 ();
 sg13g2_fill_1 FILLER_48_1544 ();
 sg13g2_decap_8 FILLER_48_1548 ();
 sg13g2_decap_4 FILLER_48_1555 ();
 sg13g2_fill_2 FILLER_48_1559 ();
 sg13g2_decap_8 FILLER_48_1597 ();
 sg13g2_decap_8 FILLER_48_1604 ();
 sg13g2_decap_8 FILLER_48_1611 ();
 sg13g2_decap_8 FILLER_48_1618 ();
 sg13g2_decap_8 FILLER_48_1625 ();
 sg13g2_fill_2 FILLER_48_1632 ();
 sg13g2_decap_8 FILLER_48_1666 ();
 sg13g2_decap_8 FILLER_48_1673 ();
 sg13g2_fill_2 FILLER_48_1680 ();
 sg13g2_decap_8 FILLER_48_1708 ();
 sg13g2_decap_8 FILLER_48_1715 ();
 sg13g2_decap_8 FILLER_48_1722 ();
 sg13g2_fill_1 FILLER_48_1729 ();
 sg13g2_fill_2 FILLER_48_1740 ();
 sg13g2_fill_1 FILLER_48_1742 ();
 sg13g2_decap_8 FILLER_48_1751 ();
 sg13g2_decap_8 FILLER_48_1758 ();
 sg13g2_decap_8 FILLER_48_1765 ();
 sg13g2_fill_2 FILLER_48_1772 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_23 ();
 sg13g2_fill_2 FILLER_49_28 ();
 sg13g2_fill_1 FILLER_49_30 ();
 sg13g2_decap_4 FILLER_49_43 ();
 sg13g2_fill_2 FILLER_49_47 ();
 sg13g2_decap_4 FILLER_49_59 ();
 sg13g2_fill_2 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_fill_2 FILLER_49_81 ();
 sg13g2_fill_2 FILLER_49_88 ();
 sg13g2_fill_1 FILLER_49_95 ();
 sg13g2_fill_1 FILLER_49_101 ();
 sg13g2_fill_2 FILLER_49_122 ();
 sg13g2_fill_1 FILLER_49_124 ();
 sg13g2_fill_1 FILLER_49_130 ();
 sg13g2_decap_4 FILLER_49_155 ();
 sg13g2_fill_1 FILLER_49_159 ();
 sg13g2_decap_4 FILLER_49_165 ();
 sg13g2_fill_1 FILLER_49_169 ();
 sg13g2_fill_1 FILLER_49_199 ();
 sg13g2_fill_1 FILLER_49_219 ();
 sg13g2_decap_8 FILLER_49_226 ();
 sg13g2_decap_8 FILLER_49_233 ();
 sg13g2_decap_8 FILLER_49_240 ();
 sg13g2_fill_1 FILLER_49_247 ();
 sg13g2_decap_4 FILLER_49_264 ();
 sg13g2_fill_1 FILLER_49_272 ();
 sg13g2_decap_4 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_293 ();
 sg13g2_decap_8 FILLER_49_300 ();
 sg13g2_decap_8 FILLER_49_307 ();
 sg13g2_fill_2 FILLER_49_314 ();
 sg13g2_fill_1 FILLER_49_316 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_4 FILLER_49_334 ();
 sg13g2_fill_1 FILLER_49_338 ();
 sg13g2_fill_1 FILLER_49_356 ();
 sg13g2_decap_4 FILLER_49_362 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_decap_8 FILLER_49_372 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_fill_2 FILLER_49_386 ();
 sg13g2_fill_2 FILLER_49_393 ();
 sg13g2_fill_1 FILLER_49_395 ();
 sg13g2_decap_8 FILLER_49_402 ();
 sg13g2_decap_8 FILLER_49_409 ();
 sg13g2_decap_4 FILLER_49_416 ();
 sg13g2_decap_4 FILLER_49_432 ();
 sg13g2_fill_1 FILLER_49_436 ();
 sg13g2_fill_1 FILLER_49_447 ();
 sg13g2_decap_8 FILLER_49_457 ();
 sg13g2_decap_8 FILLER_49_464 ();
 sg13g2_decap_8 FILLER_49_471 ();
 sg13g2_decap_8 FILLER_49_478 ();
 sg13g2_decap_8 FILLER_49_485 ();
 sg13g2_fill_2 FILLER_49_492 ();
 sg13g2_decap_8 FILLER_49_534 ();
 sg13g2_decap_8 FILLER_49_541 ();
 sg13g2_fill_2 FILLER_49_548 ();
 sg13g2_decap_8 FILLER_49_554 ();
 sg13g2_decap_8 FILLER_49_561 ();
 sg13g2_decap_8 FILLER_49_568 ();
 sg13g2_decap_8 FILLER_49_575 ();
 sg13g2_decap_8 FILLER_49_582 ();
 sg13g2_fill_2 FILLER_49_589 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_fill_2 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_655 ();
 sg13g2_decap_8 FILLER_49_662 ();
 sg13g2_decap_8 FILLER_49_669 ();
 sg13g2_decap_4 FILLER_49_702 ();
 sg13g2_fill_1 FILLER_49_706 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_4 FILLER_49_779 ();
 sg13g2_fill_2 FILLER_49_795 ();
 sg13g2_fill_1 FILLER_49_797 ();
 sg13g2_decap_8 FILLER_49_802 ();
 sg13g2_fill_2 FILLER_49_809 ();
 sg13g2_fill_1 FILLER_49_811 ();
 sg13g2_decap_8 FILLER_49_816 ();
 sg13g2_fill_2 FILLER_49_823 ();
 sg13g2_fill_1 FILLER_49_825 ();
 sg13g2_decap_8 FILLER_49_830 ();
 sg13g2_decap_4 FILLER_49_837 ();
 sg13g2_fill_2 FILLER_49_841 ();
 sg13g2_fill_1 FILLER_49_851 ();
 sg13g2_decap_8 FILLER_49_857 ();
 sg13g2_decap_8 FILLER_49_864 ();
 sg13g2_decap_8 FILLER_49_871 ();
 sg13g2_fill_2 FILLER_49_878 ();
 sg13g2_fill_1 FILLER_49_880 ();
 sg13g2_decap_8 FILLER_49_885 ();
 sg13g2_decap_8 FILLER_49_892 ();
 sg13g2_decap_8 FILLER_49_899 ();
 sg13g2_decap_8 FILLER_49_906 ();
 sg13g2_decap_8 FILLER_49_913 ();
 sg13g2_decap_8 FILLER_49_920 ();
 sg13g2_decap_8 FILLER_49_927 ();
 sg13g2_decap_8 FILLER_49_934 ();
 sg13g2_decap_8 FILLER_49_941 ();
 sg13g2_decap_4 FILLER_49_948 ();
 sg13g2_fill_1 FILLER_49_952 ();
 sg13g2_decap_4 FILLER_49_957 ();
 sg13g2_decap_8 FILLER_49_974 ();
 sg13g2_decap_4 FILLER_49_981 ();
 sg13g2_fill_1 FILLER_49_985 ();
 sg13g2_decap_4 FILLER_49_1028 ();
 sg13g2_fill_2 FILLER_49_1032 ();
 sg13g2_decap_8 FILLER_49_1047 ();
 sg13g2_decap_4 FILLER_49_1054 ();
 sg13g2_decap_4 FILLER_49_1062 ();
 sg13g2_decap_8 FILLER_49_1070 ();
 sg13g2_decap_4 FILLER_49_1096 ();
 sg13g2_decap_8 FILLER_49_1104 ();
 sg13g2_decap_8 FILLER_49_1111 ();
 sg13g2_decap_8 FILLER_49_1118 ();
 sg13g2_decap_8 FILLER_49_1125 ();
 sg13g2_decap_8 FILLER_49_1132 ();
 sg13g2_decap_4 FILLER_49_1139 ();
 sg13g2_decap_8 FILLER_49_1154 ();
 sg13g2_decap_8 FILLER_49_1161 ();
 sg13g2_decap_8 FILLER_49_1173 ();
 sg13g2_decap_8 FILLER_49_1180 ();
 sg13g2_decap_4 FILLER_49_1187 ();
 sg13g2_fill_2 FILLER_49_1191 ();
 sg13g2_decap_8 FILLER_49_1219 ();
 sg13g2_fill_1 FILLER_49_1226 ();
 sg13g2_fill_1 FILLER_49_1241 ();
 sg13g2_fill_1 FILLER_49_1247 ();
 sg13g2_decap_4 FILLER_49_1257 ();
 sg13g2_fill_2 FILLER_49_1266 ();
 sg13g2_fill_1 FILLER_49_1268 ();
 sg13g2_decap_4 FILLER_49_1274 ();
 sg13g2_fill_2 FILLER_49_1283 ();
 sg13g2_decap_8 FILLER_49_1298 ();
 sg13g2_decap_8 FILLER_49_1305 ();
 sg13g2_decap_8 FILLER_49_1312 ();
 sg13g2_decap_8 FILLER_49_1322 ();
 sg13g2_decap_8 FILLER_49_1329 ();
 sg13g2_fill_2 FILLER_49_1336 ();
 sg13g2_fill_1 FILLER_49_1338 ();
 sg13g2_decap_8 FILLER_49_1349 ();
 sg13g2_fill_2 FILLER_49_1356 ();
 sg13g2_fill_1 FILLER_49_1358 ();
 sg13g2_decap_4 FILLER_49_1390 ();
 sg13g2_fill_1 FILLER_49_1394 ();
 sg13g2_fill_2 FILLER_49_1421 ();
 sg13g2_fill_1 FILLER_49_1423 ();
 sg13g2_decap_8 FILLER_49_1463 ();
 sg13g2_decap_4 FILLER_49_1470 ();
 sg13g2_fill_2 FILLER_49_1474 ();
 sg13g2_decap_8 FILLER_49_1504 ();
 sg13g2_decap_8 FILLER_49_1511 ();
 sg13g2_decap_8 FILLER_49_1518 ();
 sg13g2_fill_2 FILLER_49_1525 ();
 sg13g2_fill_1 FILLER_49_1531 ();
 sg13g2_fill_2 FILLER_49_1561 ();
 sg13g2_decap_8 FILLER_49_1573 ();
 sg13g2_decap_8 FILLER_49_1580 ();
 sg13g2_decap_8 FILLER_49_1587 ();
 sg13g2_decap_8 FILLER_49_1594 ();
 sg13g2_decap_8 FILLER_49_1601 ();
 sg13g2_decap_8 FILLER_49_1608 ();
 sg13g2_decap_4 FILLER_49_1615 ();
 sg13g2_decap_4 FILLER_49_1622 ();
 sg13g2_fill_1 FILLER_49_1626 ();
 sg13g2_decap_8 FILLER_49_1630 ();
 sg13g2_decap_4 FILLER_49_1637 ();
 sg13g2_decap_8 FILLER_49_1679 ();
 sg13g2_decap_8 FILLER_49_1686 ();
 sg13g2_decap_8 FILLER_49_1693 ();
 sg13g2_decap_8 FILLER_49_1700 ();
 sg13g2_decap_8 FILLER_49_1707 ();
 sg13g2_fill_2 FILLER_49_1714 ();
 sg13g2_decap_4 FILLER_49_1725 ();
 sg13g2_decap_4 FILLER_49_1738 ();
 sg13g2_fill_1 FILLER_49_1742 ();
 sg13g2_decap_8 FILLER_49_1747 ();
 sg13g2_decap_8 FILLER_49_1754 ();
 sg13g2_decap_8 FILLER_49_1761 ();
 sg13g2_decap_4 FILLER_49_1768 ();
 sg13g2_fill_2 FILLER_49_1772 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_fill_1 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_30 ();
 sg13g2_decap_8 FILLER_50_37 ();
 sg13g2_fill_1 FILLER_50_44 ();
 sg13g2_fill_2 FILLER_50_49 ();
 sg13g2_fill_1 FILLER_50_51 ();
 sg13g2_fill_1 FILLER_50_56 ();
 sg13g2_decap_4 FILLER_50_76 ();
 sg13g2_fill_1 FILLER_50_80 ();
 sg13g2_fill_2 FILLER_50_93 ();
 sg13g2_fill_1 FILLER_50_95 ();
 sg13g2_fill_2 FILLER_50_102 ();
 sg13g2_fill_1 FILLER_50_104 ();
 sg13g2_fill_2 FILLER_50_109 ();
 sg13g2_decap_4 FILLER_50_121 ();
 sg13g2_fill_1 FILLER_50_125 ();
 sg13g2_decap_8 FILLER_50_130 ();
 sg13g2_fill_1 FILLER_50_137 ();
 sg13g2_fill_1 FILLER_50_146 ();
 sg13g2_fill_2 FILLER_50_157 ();
 sg13g2_decap_4 FILLER_50_169 ();
 sg13g2_fill_2 FILLER_50_173 ();
 sg13g2_fill_1 FILLER_50_185 ();
 sg13g2_decap_4 FILLER_50_196 ();
 sg13g2_decap_8 FILLER_50_208 ();
 sg13g2_fill_2 FILLER_50_219 ();
 sg13g2_fill_2 FILLER_50_226 ();
 sg13g2_fill_1 FILLER_50_228 ();
 sg13g2_decap_4 FILLER_50_235 ();
 sg13g2_fill_2 FILLER_50_251 ();
 sg13g2_decap_4 FILLER_50_258 ();
 sg13g2_decap_8 FILLER_50_267 ();
 sg13g2_decap_4 FILLER_50_274 ();
 sg13g2_decap_4 FILLER_50_291 ();
 sg13g2_fill_1 FILLER_50_295 ();
 sg13g2_decap_4 FILLER_50_301 ();
 sg13g2_fill_1 FILLER_50_305 ();
 sg13g2_fill_2 FILLER_50_310 ();
 sg13g2_decap_8 FILLER_50_318 ();
 sg13g2_decap_4 FILLER_50_325 ();
 sg13g2_decap_8 FILLER_50_334 ();
 sg13g2_decap_8 FILLER_50_341 ();
 sg13g2_decap_8 FILLER_50_353 ();
 sg13g2_decap_8 FILLER_50_360 ();
 sg13g2_fill_2 FILLER_50_367 ();
 sg13g2_fill_1 FILLER_50_369 ();
 sg13g2_decap_8 FILLER_50_375 ();
 sg13g2_decap_4 FILLER_50_382 ();
 sg13g2_fill_2 FILLER_50_386 ();
 sg13g2_decap_4 FILLER_50_398 ();
 sg13g2_fill_1 FILLER_50_402 ();
 sg13g2_fill_2 FILLER_50_413 ();
 sg13g2_fill_1 FILLER_50_415 ();
 sg13g2_decap_8 FILLER_50_421 ();
 sg13g2_decap_8 FILLER_50_428 ();
 sg13g2_decap_8 FILLER_50_435 ();
 sg13g2_fill_2 FILLER_50_446 ();
 sg13g2_fill_1 FILLER_50_448 ();
 sg13g2_decap_8 FILLER_50_454 ();
 sg13g2_decap_8 FILLER_50_461 ();
 sg13g2_decap_8 FILLER_50_468 ();
 sg13g2_decap_8 FILLER_50_475 ();
 sg13g2_decap_8 FILLER_50_482 ();
 sg13g2_decap_8 FILLER_50_489 ();
 sg13g2_decap_8 FILLER_50_496 ();
 sg13g2_decap_8 FILLER_50_503 ();
 sg13g2_decap_8 FILLER_50_514 ();
 sg13g2_decap_4 FILLER_50_521 ();
 sg13g2_fill_1 FILLER_50_525 ();
 sg13g2_decap_8 FILLER_50_535 ();
 sg13g2_fill_1 FILLER_50_542 ();
 sg13g2_fill_2 FILLER_50_569 ();
 sg13g2_fill_1 FILLER_50_571 ();
 sg13g2_fill_1 FILLER_50_582 ();
 sg13g2_decap_8 FILLER_50_614 ();
 sg13g2_decap_8 FILLER_50_621 ();
 sg13g2_decap_8 FILLER_50_628 ();
 sg13g2_fill_2 FILLER_50_643 ();
 sg13g2_decap_8 FILLER_50_650 ();
 sg13g2_decap_8 FILLER_50_657 ();
 sg13g2_fill_2 FILLER_50_664 ();
 sg13g2_fill_1 FILLER_50_666 ();
 sg13g2_fill_2 FILLER_50_679 ();
 sg13g2_fill_1 FILLER_50_681 ();
 sg13g2_decap_8 FILLER_50_685 ();
 sg13g2_decap_8 FILLER_50_692 ();
 sg13g2_decap_8 FILLER_50_699 ();
 sg13g2_decap_8 FILLER_50_706 ();
 sg13g2_decap_8 FILLER_50_713 ();
 sg13g2_fill_2 FILLER_50_720 ();
 sg13g2_decap_8 FILLER_50_730 ();
 sg13g2_decap_8 FILLER_50_737 ();
 sg13g2_decap_8 FILLER_50_744 ();
 sg13g2_decap_4 FILLER_50_751 ();
 sg13g2_fill_1 FILLER_50_755 ();
 sg13g2_decap_8 FILLER_50_760 ();
 sg13g2_decap_8 FILLER_50_767 ();
 sg13g2_decap_8 FILLER_50_774 ();
 sg13g2_decap_8 FILLER_50_781 ();
 sg13g2_decap_8 FILLER_50_802 ();
 sg13g2_fill_2 FILLER_50_809 ();
 sg13g2_decap_8 FILLER_50_821 ();
 sg13g2_fill_2 FILLER_50_828 ();
 sg13g2_fill_2 FILLER_50_838 ();
 sg13g2_decap_8 FILLER_50_866 ();
 sg13g2_fill_2 FILLER_50_873 ();
 sg13g2_fill_2 FILLER_50_883 ();
 sg13g2_decap_4 FILLER_50_898 ();
 sg13g2_fill_1 FILLER_50_902 ();
 sg13g2_decap_8 FILLER_50_907 ();
 sg13g2_decap_8 FILLER_50_914 ();
 sg13g2_decap_8 FILLER_50_921 ();
 sg13g2_decap_8 FILLER_50_928 ();
 sg13g2_decap_4 FILLER_50_935 ();
 sg13g2_fill_2 FILLER_50_974 ();
 sg13g2_decap_4 FILLER_50_984 ();
 sg13g2_decap_8 FILLER_50_997 ();
 sg13g2_decap_8 FILLER_50_1004 ();
 sg13g2_decap_8 FILLER_50_1011 ();
 sg13g2_decap_8 FILLER_50_1018 ();
 sg13g2_decap_8 FILLER_50_1025 ();
 sg13g2_decap_8 FILLER_50_1032 ();
 sg13g2_fill_2 FILLER_50_1039 ();
 sg13g2_fill_1 FILLER_50_1041 ();
 sg13g2_fill_2 FILLER_50_1053 ();
 sg13g2_fill_1 FILLER_50_1055 ();
 sg13g2_decap_8 FILLER_50_1066 ();
 sg13g2_decap_8 FILLER_50_1073 ();
 sg13g2_decap_4 FILLER_50_1088 ();
 sg13g2_decap_8 FILLER_50_1100 ();
 sg13g2_fill_2 FILLER_50_1107 ();
 sg13g2_fill_2 FILLER_50_1129 ();
 sg13g2_fill_1 FILLER_50_1131 ();
 sg13g2_fill_2 FILLER_50_1136 ();
 sg13g2_fill_1 FILLER_50_1138 ();
 sg13g2_decap_4 FILLER_50_1149 ();
 sg13g2_fill_1 FILLER_50_1153 ();
 sg13g2_decap_8 FILLER_50_1158 ();
 sg13g2_decap_4 FILLER_50_1165 ();
 sg13g2_fill_2 FILLER_50_1169 ();
 sg13g2_decap_8 FILLER_50_1175 ();
 sg13g2_decap_8 FILLER_50_1182 ();
 sg13g2_decap_4 FILLER_50_1189 ();
 sg13g2_fill_2 FILLER_50_1193 ();
 sg13g2_fill_2 FILLER_50_1201 ();
 sg13g2_decap_8 FILLER_50_1211 ();
 sg13g2_decap_8 FILLER_50_1218 ();
 sg13g2_decap_8 FILLER_50_1225 ();
 sg13g2_fill_2 FILLER_50_1232 ();
 sg13g2_fill_1 FILLER_50_1234 ();
 sg13g2_decap_8 FILLER_50_1240 ();
 sg13g2_fill_1 FILLER_50_1247 ();
 sg13g2_decap_8 FILLER_50_1262 ();
 sg13g2_fill_1 FILLER_50_1269 ();
 sg13g2_decap_4 FILLER_50_1280 ();
 sg13g2_fill_2 FILLER_50_1284 ();
 sg13g2_decap_4 FILLER_50_1303 ();
 sg13g2_fill_1 FILLER_50_1307 ();
 sg13g2_decap_8 FILLER_50_1312 ();
 sg13g2_fill_2 FILLER_50_1319 ();
 sg13g2_fill_1 FILLER_50_1321 ();
 sg13g2_fill_2 FILLER_50_1330 ();
 sg13g2_decap_4 FILLER_50_1344 ();
 sg13g2_decap_8 FILLER_50_1352 ();
 sg13g2_decap_4 FILLER_50_1359 ();
 sg13g2_fill_1 FILLER_50_1363 ();
 sg13g2_decap_8 FILLER_50_1369 ();
 sg13g2_decap_8 FILLER_50_1376 ();
 sg13g2_decap_8 FILLER_50_1383 ();
 sg13g2_decap_8 FILLER_50_1390 ();
 sg13g2_decap_8 FILLER_50_1397 ();
 sg13g2_decap_8 FILLER_50_1404 ();
 sg13g2_decap_8 FILLER_50_1411 ();
 sg13g2_decap_8 FILLER_50_1418 ();
 sg13g2_decap_8 FILLER_50_1425 ();
 sg13g2_decap_8 FILLER_50_1432 ();
 sg13g2_decap_8 FILLER_50_1442 ();
 sg13g2_fill_2 FILLER_50_1449 ();
 sg13g2_decap_8 FILLER_50_1462 ();
 sg13g2_decap_4 FILLER_50_1469 ();
 sg13g2_fill_1 FILLER_50_1473 ();
 sg13g2_decap_4 FILLER_50_1479 ();
 sg13g2_fill_2 FILLER_50_1503 ();
 sg13g2_fill_1 FILLER_50_1505 ();
 sg13g2_decap_8 FILLER_50_1510 ();
 sg13g2_decap_4 FILLER_50_1517 ();
 sg13g2_fill_1 FILLER_50_1521 ();
 sg13g2_fill_2 FILLER_50_1526 ();
 sg13g2_fill_1 FILLER_50_1536 ();
 sg13g2_fill_1 FILLER_50_1540 ();
 sg13g2_fill_1 FILLER_50_1552 ();
 sg13g2_fill_1 FILLER_50_1566 ();
 sg13g2_decap_8 FILLER_50_1582 ();
 sg13g2_decap_8 FILLER_50_1589 ();
 sg13g2_decap_8 FILLER_50_1596 ();
 sg13g2_decap_8 FILLER_50_1603 ();
 sg13g2_decap_8 FILLER_50_1610 ();
 sg13g2_fill_1 FILLER_50_1617 ();
 sg13g2_decap_8 FILLER_50_1635 ();
 sg13g2_fill_1 FILLER_50_1647 ();
 sg13g2_decap_8 FILLER_50_1673 ();
 sg13g2_decap_8 FILLER_50_1680 ();
 sg13g2_decap_8 FILLER_50_1687 ();
 sg13g2_decap_8 FILLER_50_1694 ();
 sg13g2_fill_2 FILLER_50_1701 ();
 sg13g2_decap_8 FILLER_50_1707 ();
 sg13g2_decap_4 FILLER_50_1714 ();
 sg13g2_decap_8 FILLER_50_1721 ();
 sg13g2_decap_4 FILLER_50_1728 ();
 sg13g2_decap_8 FILLER_50_1759 ();
 sg13g2_decap_8 FILLER_50_1766 ();
 sg13g2_fill_1 FILLER_50_1773 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_fill_2 FILLER_51_32 ();
 sg13g2_fill_1 FILLER_51_34 ();
 sg13g2_decap_4 FILLER_51_44 ();
 sg13g2_fill_1 FILLER_51_53 ();
 sg13g2_decap_8 FILLER_51_68 ();
 sg13g2_decap_8 FILLER_51_75 ();
 sg13g2_decap_4 FILLER_51_82 ();
 sg13g2_fill_2 FILLER_51_86 ();
 sg13g2_decap_4 FILLER_51_98 ();
 sg13g2_decap_4 FILLER_51_106 ();
 sg13g2_fill_1 FILLER_51_110 ();
 sg13g2_fill_2 FILLER_51_117 ();
 sg13g2_decap_8 FILLER_51_123 ();
 sg13g2_decap_4 FILLER_51_130 ();
 sg13g2_fill_1 FILLER_51_134 ();
 sg13g2_decap_4 FILLER_51_145 ();
 sg13g2_fill_2 FILLER_51_149 ();
 sg13g2_decap_4 FILLER_51_156 ();
 sg13g2_fill_2 FILLER_51_160 ();
 sg13g2_fill_2 FILLER_51_172 ();
 sg13g2_decap_4 FILLER_51_184 ();
 sg13g2_fill_1 FILLER_51_188 ();
 sg13g2_fill_1 FILLER_51_194 ();
 sg13g2_decap_4 FILLER_51_199 ();
 sg13g2_fill_2 FILLER_51_203 ();
 sg13g2_decap_4 FILLER_51_210 ();
 sg13g2_decap_8 FILLER_51_225 ();
 sg13g2_decap_8 FILLER_51_232 ();
 sg13g2_decap_4 FILLER_51_248 ();
 sg13g2_fill_1 FILLER_51_252 ();
 sg13g2_fill_1 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_264 ();
 sg13g2_decap_8 FILLER_51_271 ();
 sg13g2_decap_4 FILLER_51_278 ();
 sg13g2_decap_4 FILLER_51_292 ();
 sg13g2_fill_2 FILLER_51_296 ();
 sg13g2_fill_2 FILLER_51_303 ();
 sg13g2_fill_2 FILLER_51_310 ();
 sg13g2_decap_8 FILLER_51_317 ();
 sg13g2_fill_1 FILLER_51_324 ();
 sg13g2_decap_8 FILLER_51_335 ();
 sg13g2_decap_8 FILLER_51_347 ();
 sg13g2_decap_4 FILLER_51_354 ();
 sg13g2_fill_2 FILLER_51_358 ();
 sg13g2_decap_8 FILLER_51_365 ();
 sg13g2_decap_8 FILLER_51_372 ();
 sg13g2_decap_8 FILLER_51_379 ();
 sg13g2_decap_4 FILLER_51_390 ();
 sg13g2_fill_2 FILLER_51_394 ();
 sg13g2_fill_2 FILLER_51_408 ();
 sg13g2_fill_2 FILLER_51_433 ();
 sg13g2_fill_1 FILLER_51_439 ();
 sg13g2_decap_4 FILLER_51_450 ();
 sg13g2_decap_8 FILLER_51_459 ();
 sg13g2_decap_8 FILLER_51_466 ();
 sg13g2_decap_8 FILLER_51_473 ();
 sg13g2_decap_8 FILLER_51_486 ();
 sg13g2_fill_2 FILLER_51_493 ();
 sg13g2_fill_1 FILLER_51_495 ();
 sg13g2_decap_8 FILLER_51_500 ();
 sg13g2_decap_8 FILLER_51_507 ();
 sg13g2_fill_1 FILLER_51_514 ();
 sg13g2_decap_8 FILLER_51_527 ();
 sg13g2_decap_8 FILLER_51_534 ();
 sg13g2_decap_8 FILLER_51_541 ();
 sg13g2_decap_8 FILLER_51_548 ();
 sg13g2_fill_2 FILLER_51_555 ();
 sg13g2_decap_4 FILLER_51_579 ();
 sg13g2_fill_2 FILLER_51_583 ();
 sg13g2_decap_8 FILLER_51_589 ();
 sg13g2_decap_8 FILLER_51_596 ();
 sg13g2_decap_8 FILLER_51_603 ();
 sg13g2_decap_4 FILLER_51_610 ();
 sg13g2_fill_1 FILLER_51_614 ();
 sg13g2_decap_8 FILLER_51_619 ();
 sg13g2_decap_8 FILLER_51_626 ();
 sg13g2_decap_8 FILLER_51_633 ();
 sg13g2_fill_2 FILLER_51_640 ();
 sg13g2_fill_1 FILLER_51_642 ();
 sg13g2_fill_1 FILLER_51_653 ();
 sg13g2_decap_8 FILLER_51_670 ();
 sg13g2_fill_2 FILLER_51_677 ();
 sg13g2_fill_1 FILLER_51_679 ();
 sg13g2_decap_4 FILLER_51_683 ();
 sg13g2_fill_2 FILLER_51_687 ();
 sg13g2_decap_8 FILLER_51_704 ();
 sg13g2_decap_8 FILLER_51_711 ();
 sg13g2_fill_1 FILLER_51_718 ();
 sg13g2_fill_1 FILLER_51_728 ();
 sg13g2_fill_2 FILLER_51_745 ();
 sg13g2_decap_8 FILLER_51_751 ();
 sg13g2_decap_8 FILLER_51_758 ();
 sg13g2_decap_8 FILLER_51_765 ();
 sg13g2_decap_8 FILLER_51_772 ();
 sg13g2_decap_8 FILLER_51_779 ();
 sg13g2_decap_4 FILLER_51_786 ();
 sg13g2_fill_2 FILLER_51_790 ();
 sg13g2_decap_8 FILLER_51_800 ();
 sg13g2_decap_8 FILLER_51_807 ();
 sg13g2_decap_8 FILLER_51_814 ();
 sg13g2_decap_8 FILLER_51_821 ();
 sg13g2_decap_4 FILLER_51_828 ();
 sg13g2_fill_2 FILLER_51_837 ();
 sg13g2_decap_8 FILLER_51_847 ();
 sg13g2_fill_1 FILLER_51_854 ();
 sg13g2_fill_2 FILLER_51_859 ();
 sg13g2_decap_4 FILLER_51_866 ();
 sg13g2_fill_1 FILLER_51_870 ();
 sg13g2_decap_8 FILLER_51_879 ();
 sg13g2_decap_8 FILLER_51_886 ();
 sg13g2_fill_1 FILLER_51_893 ();
 sg13g2_decap_8 FILLER_51_924 ();
 sg13g2_decap_8 FILLER_51_935 ();
 sg13g2_decap_8 FILLER_51_942 ();
 sg13g2_fill_1 FILLER_51_949 ();
 sg13g2_decap_8 FILLER_51_954 ();
 sg13g2_decap_8 FILLER_51_961 ();
 sg13g2_decap_4 FILLER_51_968 ();
 sg13g2_decap_8 FILLER_51_977 ();
 sg13g2_fill_2 FILLER_51_984 ();
 sg13g2_fill_1 FILLER_51_986 ();
 sg13g2_decap_8 FILLER_51_995 ();
 sg13g2_decap_8 FILLER_51_1006 ();
 sg13g2_decap_8 FILLER_51_1013 ();
 sg13g2_decap_8 FILLER_51_1020 ();
 sg13g2_decap_8 FILLER_51_1062 ();
 sg13g2_decap_8 FILLER_51_1069 ();
 sg13g2_decap_8 FILLER_51_1076 ();
 sg13g2_decap_4 FILLER_51_1083 ();
 sg13g2_fill_1 FILLER_51_1087 ();
 sg13g2_decap_8 FILLER_51_1102 ();
 sg13g2_decap_8 FILLER_51_1109 ();
 sg13g2_decap_8 FILLER_51_1116 ();
 sg13g2_decap_8 FILLER_51_1123 ();
 sg13g2_decap_8 FILLER_51_1130 ();
 sg13g2_decap_4 FILLER_51_1137 ();
 sg13g2_fill_2 FILLER_51_1141 ();
 sg13g2_decap_8 FILLER_51_1152 ();
 sg13g2_decap_4 FILLER_51_1159 ();
 sg13g2_fill_1 FILLER_51_1163 ();
 sg13g2_fill_1 FILLER_51_1193 ();
 sg13g2_decap_8 FILLER_51_1204 ();
 sg13g2_decap_8 FILLER_51_1211 ();
 sg13g2_decap_8 FILLER_51_1222 ();
 sg13g2_decap_8 FILLER_51_1229 ();
 sg13g2_decap_8 FILLER_51_1236 ();
 sg13g2_decap_8 FILLER_51_1243 ();
 sg13g2_decap_8 FILLER_51_1250 ();
 sg13g2_decap_8 FILLER_51_1257 ();
 sg13g2_decap_8 FILLER_51_1269 ();
 sg13g2_decap_8 FILLER_51_1276 ();
 sg13g2_decap_4 FILLER_51_1283 ();
 sg13g2_fill_2 FILLER_51_1287 ();
 sg13g2_decap_8 FILLER_51_1297 ();
 sg13g2_decap_8 FILLER_51_1304 ();
 sg13g2_decap_4 FILLER_51_1311 ();
 sg13g2_fill_1 FILLER_51_1315 ();
 sg13g2_decap_8 FILLER_51_1320 ();
 sg13g2_decap_8 FILLER_51_1327 ();
 sg13g2_fill_1 FILLER_51_1334 ();
 sg13g2_decap_8 FILLER_51_1347 ();
 sg13g2_decap_8 FILLER_51_1354 ();
 sg13g2_fill_2 FILLER_51_1387 ();
 sg13g2_decap_8 FILLER_51_1397 ();
 sg13g2_decap_4 FILLER_51_1404 ();
 sg13g2_fill_2 FILLER_51_1408 ();
 sg13g2_decap_8 FILLER_51_1414 ();
 sg13g2_fill_2 FILLER_51_1421 ();
 sg13g2_decap_8 FILLER_51_1430 ();
 sg13g2_decap_4 FILLER_51_1437 ();
 sg13g2_fill_2 FILLER_51_1441 ();
 sg13g2_fill_1 FILLER_51_1461 ();
 sg13g2_decap_4 FILLER_51_1467 ();
 sg13g2_fill_2 FILLER_51_1474 ();
 sg13g2_decap_4 FILLER_51_1511 ();
 sg13g2_fill_1 FILLER_51_1515 ();
 sg13g2_fill_2 FILLER_51_1525 ();
 sg13g2_fill_1 FILLER_51_1527 ();
 sg13g2_decap_4 FILLER_51_1533 ();
 sg13g2_decap_8 FILLER_51_1556 ();
 sg13g2_decap_4 FILLER_51_1563 ();
 sg13g2_fill_1 FILLER_51_1567 ();
 sg13g2_decap_8 FILLER_51_1600 ();
 sg13g2_decap_4 FILLER_51_1607 ();
 sg13g2_fill_2 FILLER_51_1616 ();
 sg13g2_fill_1 FILLER_51_1618 ();
 sg13g2_decap_8 FILLER_51_1634 ();
 sg13g2_fill_2 FILLER_51_1641 ();
 sg13g2_fill_1 FILLER_51_1643 ();
 sg13g2_fill_1 FILLER_51_1652 ();
 sg13g2_decap_8 FILLER_51_1658 ();
 sg13g2_fill_2 FILLER_51_1665 ();
 sg13g2_fill_1 FILLER_51_1667 ();
 sg13g2_decap_8 FILLER_51_1683 ();
 sg13g2_decap_4 FILLER_51_1690 ();
 sg13g2_fill_2 FILLER_51_1736 ();
 sg13g2_fill_2 FILLER_51_1772 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_4 FILLER_52_28 ();
 sg13g2_fill_2 FILLER_52_32 ();
 sg13g2_fill_1 FILLER_52_44 ();
 sg13g2_fill_2 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_51 ();
 sg13g2_fill_1 FILLER_52_62 ();
 sg13g2_decap_4 FILLER_52_68 ();
 sg13g2_fill_1 FILLER_52_81 ();
 sg13g2_fill_2 FILLER_52_87 ();
 sg13g2_decap_4 FILLER_52_99 ();
 sg13g2_fill_2 FILLER_52_111 ();
 sg13g2_decap_4 FILLER_52_119 ();
 sg13g2_decap_4 FILLER_52_134 ();
 sg13g2_fill_1 FILLER_52_138 ();
 sg13g2_fill_2 FILLER_52_144 ();
 sg13g2_decap_8 FILLER_52_151 ();
 sg13g2_fill_1 FILLER_52_158 ();
 sg13g2_fill_2 FILLER_52_163 ();
 sg13g2_fill_1 FILLER_52_165 ();
 sg13g2_decap_8 FILLER_52_183 ();
 sg13g2_fill_2 FILLER_52_190 ();
 sg13g2_fill_1 FILLER_52_192 ();
 sg13g2_decap_4 FILLER_52_203 ();
 sg13g2_fill_2 FILLER_52_218 ();
 sg13g2_decap_8 FILLER_52_234 ();
 sg13g2_decap_4 FILLER_52_241 ();
 sg13g2_decap_8 FILLER_52_249 ();
 sg13g2_decap_4 FILLER_52_256 ();
 sg13g2_decap_8 FILLER_52_264 ();
 sg13g2_fill_2 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_284 ();
 sg13g2_fill_1 FILLER_52_296 ();
 sg13g2_fill_1 FILLER_52_307 ();
 sg13g2_fill_2 FILLER_52_320 ();
 sg13g2_fill_1 FILLER_52_322 ();
 sg13g2_fill_2 FILLER_52_329 ();
 sg13g2_decap_4 FILLER_52_336 ();
 sg13g2_decap_4 FILLER_52_345 ();
 sg13g2_fill_2 FILLER_52_366 ();
 sg13g2_fill_1 FILLER_52_368 ();
 sg13g2_fill_1 FILLER_52_374 ();
 sg13g2_decap_8 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_388 ();
 sg13g2_fill_1 FILLER_52_395 ();
 sg13g2_fill_1 FILLER_52_401 ();
 sg13g2_decap_4 FILLER_52_412 ();
 sg13g2_fill_1 FILLER_52_416 ();
 sg13g2_fill_2 FILLER_52_422 ();
 sg13g2_fill_1 FILLER_52_424 ();
 sg13g2_decap_8 FILLER_52_430 ();
 sg13g2_decap_8 FILLER_52_437 ();
 sg13g2_fill_2 FILLER_52_444 ();
 sg13g2_fill_1 FILLER_52_446 ();
 sg13g2_fill_2 FILLER_52_452 ();
 sg13g2_decap_8 FILLER_52_459 ();
 sg13g2_decap_8 FILLER_52_466 ();
 sg13g2_decap_8 FILLER_52_473 ();
 sg13g2_decap_8 FILLER_52_480 ();
 sg13g2_fill_2 FILLER_52_487 ();
 sg13g2_fill_2 FILLER_52_558 ();
 sg13g2_fill_1 FILLER_52_560 ();
 sg13g2_fill_1 FILLER_52_566 ();
 sg13g2_decap_4 FILLER_52_593 ();
 sg13g2_fill_1 FILLER_52_597 ();
 sg13g2_decap_8 FILLER_52_634 ();
 sg13g2_decap_8 FILLER_52_641 ();
 sg13g2_decap_8 FILLER_52_648 ();
 sg13g2_fill_2 FILLER_52_655 ();
 sg13g2_decap_8 FILLER_52_660 ();
 sg13g2_decap_8 FILLER_52_667 ();
 sg13g2_fill_1 FILLER_52_674 ();
 sg13g2_fill_2 FILLER_52_680 ();
 sg13g2_decap_8 FILLER_52_690 ();
 sg13g2_fill_2 FILLER_52_697 ();
 sg13g2_decap_4 FILLER_52_704 ();
 sg13g2_fill_2 FILLER_52_708 ();
 sg13g2_decap_4 FILLER_52_714 ();
 sg13g2_decap_4 FILLER_52_729 ();
 sg13g2_fill_1 FILLER_52_733 ();
 sg13g2_fill_2 FILLER_52_739 ();
 sg13g2_decap_8 FILLER_52_745 ();
 sg13g2_decap_4 FILLER_52_752 ();
 sg13g2_fill_2 FILLER_52_756 ();
 sg13g2_decap_4 FILLER_52_778 ();
 sg13g2_fill_2 FILLER_52_782 ();
 sg13g2_decap_8 FILLER_52_787 ();
 sg13g2_decap_8 FILLER_52_794 ();
 sg13g2_fill_2 FILLER_52_801 ();
 sg13g2_fill_1 FILLER_52_803 ();
 sg13g2_decap_8 FILLER_52_808 ();
 sg13g2_decap_8 FILLER_52_815 ();
 sg13g2_decap_8 FILLER_52_822 ();
 sg13g2_decap_8 FILLER_52_829 ();
 sg13g2_decap_8 FILLER_52_836 ();
 sg13g2_fill_1 FILLER_52_843 ();
 sg13g2_fill_2 FILLER_52_849 ();
 sg13g2_decap_8 FILLER_52_855 ();
 sg13g2_decap_8 FILLER_52_862 ();
 sg13g2_decap_4 FILLER_52_869 ();
 sg13g2_fill_1 FILLER_52_884 ();
 sg13g2_fill_2 FILLER_52_890 ();
 sg13g2_fill_1 FILLER_52_892 ();
 sg13g2_decap_8 FILLER_52_910 ();
 sg13g2_decap_8 FILLER_52_917 ();
 sg13g2_fill_1 FILLER_52_950 ();
 sg13g2_decap_8 FILLER_52_955 ();
 sg13g2_fill_1 FILLER_52_962 ();
 sg13g2_decap_8 FILLER_52_971 ();
 sg13g2_fill_2 FILLER_52_978 ();
 sg13g2_fill_1 FILLER_52_980 ();
 sg13g2_decap_4 FILLER_52_1014 ();
 sg13g2_fill_2 FILLER_52_1018 ();
 sg13g2_fill_2 FILLER_52_1025 ();
 sg13g2_decap_8 FILLER_52_1038 ();
 sg13g2_decap_4 FILLER_52_1045 ();
 sg13g2_fill_2 FILLER_52_1049 ();
 sg13g2_decap_8 FILLER_52_1062 ();
 sg13g2_decap_8 FILLER_52_1069 ();
 sg13g2_decap_8 FILLER_52_1076 ();
 sg13g2_decap_4 FILLER_52_1083 ();
 sg13g2_fill_1 FILLER_52_1097 ();
 sg13g2_fill_2 FILLER_52_1102 ();
 sg13g2_fill_1 FILLER_52_1104 ();
 sg13g2_decap_4 FILLER_52_1110 ();
 sg13g2_fill_2 FILLER_52_1114 ();
 sg13g2_decap_4 FILLER_52_1125 ();
 sg13g2_decap_4 FILLER_52_1132 ();
 sg13g2_fill_1 FILLER_52_1136 ();
 sg13g2_decap_4 FILLER_52_1142 ();
 sg13g2_fill_2 FILLER_52_1146 ();
 sg13g2_decap_8 FILLER_52_1152 ();
 sg13g2_decap_8 FILLER_52_1159 ();
 sg13g2_decap_8 FILLER_52_1166 ();
 sg13g2_decap_8 FILLER_52_1173 ();
 sg13g2_decap_8 FILLER_52_1180 ();
 sg13g2_decap_4 FILLER_52_1187 ();
 sg13g2_fill_2 FILLER_52_1191 ();
 sg13g2_fill_2 FILLER_52_1201 ();
 sg13g2_fill_1 FILLER_52_1203 ();
 sg13g2_fill_1 FILLER_52_1236 ();
 sg13g2_decap_8 FILLER_52_1256 ();
 sg13g2_fill_2 FILLER_52_1263 ();
 sg13g2_decap_8 FILLER_52_1274 ();
 sg13g2_decap_8 FILLER_52_1281 ();
 sg13g2_fill_1 FILLER_52_1288 ();
 sg13g2_decap_8 FILLER_52_1320 ();
 sg13g2_fill_1 FILLER_52_1327 ();
 sg13g2_decap_8 FILLER_52_1348 ();
 sg13g2_decap_8 FILLER_52_1355 ();
 sg13g2_decap_4 FILLER_52_1362 ();
 sg13g2_fill_1 FILLER_52_1366 ();
 sg13g2_decap_8 FILLER_52_1371 ();
 sg13g2_decap_8 FILLER_52_1378 ();
 sg13g2_decap_8 FILLER_52_1385 ();
 sg13g2_decap_8 FILLER_52_1392 ();
 sg13g2_decap_4 FILLER_52_1399 ();
 sg13g2_fill_2 FILLER_52_1435 ();
 sg13g2_decap_8 FILLER_52_1455 ();
 sg13g2_fill_1 FILLER_52_1462 ();
 sg13g2_fill_2 FILLER_52_1507 ();
 sg13g2_fill_2 FILLER_52_1535 ();
 sg13g2_fill_1 FILLER_52_1537 ();
 sg13g2_decap_8 FILLER_52_1556 ();
 sg13g2_fill_2 FILLER_52_1563 ();
 sg13g2_fill_1 FILLER_52_1565 ();
 sg13g2_decap_8 FILLER_52_1571 ();
 sg13g2_fill_2 FILLER_52_1578 ();
 sg13g2_decap_8 FILLER_52_1584 ();
 sg13g2_decap_4 FILLER_52_1591 ();
 sg13g2_decap_8 FILLER_52_1598 ();
 sg13g2_fill_2 FILLER_52_1605 ();
 sg13g2_fill_1 FILLER_52_1607 ();
 sg13g2_fill_1 FILLER_52_1624 ();
 sg13g2_fill_2 FILLER_52_1633 ();
 sg13g2_fill_1 FILLER_52_1635 ();
 sg13g2_decap_4 FILLER_52_1662 ();
 sg13g2_fill_2 FILLER_52_1666 ();
 sg13g2_decap_8 FILLER_52_1677 ();
 sg13g2_fill_2 FILLER_52_1684 ();
 sg13g2_fill_1 FILLER_52_1686 ();
 sg13g2_fill_2 FILLER_52_1713 ();
 sg13g2_fill_1 FILLER_52_1715 ();
 sg13g2_decap_8 FILLER_52_1724 ();
 sg13g2_decap_8 FILLER_52_1731 ();
 sg13g2_fill_2 FILLER_52_1750 ();
 sg13g2_fill_1 FILLER_52_1752 ();
 sg13g2_decap_8 FILLER_52_1757 ();
 sg13g2_decap_8 FILLER_52_1764 ();
 sg13g2_fill_2 FILLER_52_1771 ();
 sg13g2_fill_1 FILLER_52_1773 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_4 FILLER_53_28 ();
 sg13g2_fill_1 FILLER_53_32 ();
 sg13g2_fill_1 FILLER_53_38 ();
 sg13g2_decap_8 FILLER_53_55 ();
 sg13g2_decap_8 FILLER_53_62 ();
 sg13g2_fill_2 FILLER_53_74 ();
 sg13g2_decap_4 FILLER_53_81 ();
 sg13g2_fill_1 FILLER_53_85 ();
 sg13g2_decap_8 FILLER_53_90 ();
 sg13g2_fill_2 FILLER_53_97 ();
 sg13g2_decap_8 FILLER_53_104 ();
 sg13g2_decap_8 FILLER_53_111 ();
 sg13g2_decap_4 FILLER_53_118 ();
 sg13g2_decap_4 FILLER_53_127 ();
 sg13g2_fill_2 FILLER_53_131 ();
 sg13g2_fill_2 FILLER_53_137 ();
 sg13g2_fill_2 FILLER_53_147 ();
 sg13g2_fill_1 FILLER_53_153 ();
 sg13g2_fill_1 FILLER_53_165 ();
 sg13g2_fill_2 FILLER_53_170 ();
 sg13g2_decap_8 FILLER_53_180 ();
 sg13g2_decap_8 FILLER_53_187 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_decap_4 FILLER_53_224 ();
 sg13g2_decap_4 FILLER_53_232 ();
 sg13g2_fill_1 FILLER_53_236 ();
 sg13g2_decap_8 FILLER_53_242 ();
 sg13g2_decap_4 FILLER_53_249 ();
 sg13g2_decap_4 FILLER_53_257 ();
 sg13g2_decap_8 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_273 ();
 sg13g2_decap_8 FILLER_53_280 ();
 sg13g2_decap_8 FILLER_53_287 ();
 sg13g2_decap_8 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_301 ();
 sg13g2_fill_2 FILLER_53_308 ();
 sg13g2_fill_1 FILLER_53_310 ();
 sg13g2_fill_2 FILLER_53_324 ();
 sg13g2_fill_1 FILLER_53_326 ();
 sg13g2_decap_8 FILLER_53_332 ();
 sg13g2_decap_4 FILLER_53_339 ();
 sg13g2_fill_1 FILLER_53_343 ();
 sg13g2_decap_4 FILLER_53_349 ();
 sg13g2_fill_1 FILLER_53_353 ();
 sg13g2_decap_4 FILLER_53_370 ();
 sg13g2_decap_8 FILLER_53_379 ();
 sg13g2_decap_8 FILLER_53_386 ();
 sg13g2_fill_1 FILLER_53_393 ();
 sg13g2_decap_8 FILLER_53_398 ();
 sg13g2_decap_8 FILLER_53_405 ();
 sg13g2_decap_8 FILLER_53_412 ();
 sg13g2_fill_2 FILLER_53_419 ();
 sg13g2_fill_1 FILLER_53_421 ();
 sg13g2_decap_8 FILLER_53_433 ();
 sg13g2_decap_8 FILLER_53_440 ();
 sg13g2_fill_1 FILLER_53_447 ();
 sg13g2_decap_4 FILLER_53_453 ();
 sg13g2_fill_1 FILLER_53_463 ();
 sg13g2_decap_8 FILLER_53_467 ();
 sg13g2_decap_8 FILLER_53_474 ();
 sg13g2_decap_8 FILLER_53_481 ();
 sg13g2_decap_8 FILLER_53_488 ();
 sg13g2_decap_8 FILLER_53_495 ();
 sg13g2_decap_8 FILLER_53_502 ();
 sg13g2_decap_4 FILLER_53_509 ();
 sg13g2_decap_8 FILLER_53_542 ();
 sg13g2_decap_8 FILLER_53_549 ();
 sg13g2_decap_8 FILLER_53_556 ();
 sg13g2_decap_8 FILLER_53_563 ();
 sg13g2_decap_8 FILLER_53_570 ();
 sg13g2_decap_8 FILLER_53_577 ();
 sg13g2_decap_8 FILLER_53_596 ();
 sg13g2_decap_8 FILLER_53_603 ();
 sg13g2_decap_8 FILLER_53_610 ();
 sg13g2_decap_8 FILLER_53_617 ();
 sg13g2_decap_4 FILLER_53_624 ();
 sg13g2_fill_1 FILLER_53_628 ();
 sg13g2_decap_8 FILLER_53_655 ();
 sg13g2_decap_8 FILLER_53_662 ();
 sg13g2_fill_2 FILLER_53_669 ();
 sg13g2_decap_4 FILLER_53_692 ();
 sg13g2_decap_8 FILLER_53_708 ();
 sg13g2_decap_8 FILLER_53_715 ();
 sg13g2_decap_8 FILLER_53_727 ();
 sg13g2_decap_8 FILLER_53_734 ();
 sg13g2_decap_8 FILLER_53_741 ();
 sg13g2_decap_4 FILLER_53_748 ();
 sg13g2_decap_8 FILLER_53_756 ();
 sg13g2_decap_8 FILLER_53_763 ();
 sg13g2_decap_4 FILLER_53_770 ();
 sg13g2_fill_1 FILLER_53_774 ();
 sg13g2_decap_8 FILLER_53_778 ();
 sg13g2_fill_2 FILLER_53_823 ();
 sg13g2_fill_1 FILLER_53_825 ();
 sg13g2_decap_8 FILLER_53_830 ();
 sg13g2_decap_4 FILLER_53_837 ();
 sg13g2_fill_1 FILLER_53_841 ();
 sg13g2_decap_4 FILLER_53_846 ();
 sg13g2_fill_1 FILLER_53_850 ();
 sg13g2_fill_2 FILLER_53_859 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_fill_2 FILLER_53_867 ();
 sg13g2_fill_1 FILLER_53_869 ();
 sg13g2_decap_8 FILLER_53_878 ();
 sg13g2_decap_8 FILLER_53_885 ();
 sg13g2_decap_4 FILLER_53_892 ();
 sg13g2_fill_1 FILLER_53_896 ();
 sg13g2_fill_2 FILLER_53_911 ();
 sg13g2_fill_2 FILLER_53_929 ();
 sg13g2_decap_8 FILLER_53_944 ();
 sg13g2_decap_8 FILLER_53_951 ();
 sg13g2_decap_4 FILLER_53_958 ();
 sg13g2_fill_2 FILLER_53_962 ();
 sg13g2_decap_8 FILLER_53_970 ();
 sg13g2_decap_4 FILLER_53_977 ();
 sg13g2_fill_2 FILLER_53_981 ();
 sg13g2_decap_8 FILLER_53_988 ();
 sg13g2_fill_2 FILLER_53_999 ();
 sg13g2_fill_1 FILLER_53_1001 ();
 sg13g2_fill_2 FILLER_53_1011 ();
 sg13g2_fill_2 FILLER_53_1018 ();
 sg13g2_fill_1 FILLER_53_1020 ();
 sg13g2_fill_1 FILLER_53_1036 ();
 sg13g2_fill_2 FILLER_53_1041 ();
 sg13g2_fill_1 FILLER_53_1043 ();
 sg13g2_fill_2 FILLER_53_1055 ();
 sg13g2_fill_1 FILLER_53_1057 ();
 sg13g2_decap_8 FILLER_53_1073 ();
 sg13g2_decap_8 FILLER_53_1080 ();
 sg13g2_decap_8 FILLER_53_1087 ();
 sg13g2_decap_8 FILLER_53_1094 ();
 sg13g2_decap_8 FILLER_53_1101 ();
 sg13g2_decap_4 FILLER_53_1108 ();
 sg13g2_fill_2 FILLER_53_1112 ();
 sg13g2_fill_2 FILLER_53_1121 ();
 sg13g2_fill_2 FILLER_53_1128 ();
 sg13g2_fill_2 FILLER_53_1135 ();
 sg13g2_fill_1 FILLER_53_1137 ();
 sg13g2_decap_8 FILLER_53_1142 ();
 sg13g2_fill_1 FILLER_53_1149 ();
 sg13g2_decap_8 FILLER_53_1155 ();
 sg13g2_decap_8 FILLER_53_1162 ();
 sg13g2_fill_2 FILLER_53_1169 ();
 sg13g2_decap_8 FILLER_53_1175 ();
 sg13g2_decap_8 FILLER_53_1182 ();
 sg13g2_decap_8 FILLER_53_1189 ();
 sg13g2_decap_8 FILLER_53_1196 ();
 sg13g2_fill_1 FILLER_53_1203 ();
 sg13g2_decap_8 FILLER_53_1209 ();
 sg13g2_fill_1 FILLER_53_1216 ();
 sg13g2_fill_1 FILLER_53_1221 ();
 sg13g2_fill_2 FILLER_53_1235 ();
 sg13g2_fill_2 FILLER_53_1241 ();
 sg13g2_fill_1 FILLER_53_1243 ();
 sg13g2_fill_1 FILLER_53_1249 ();
 sg13g2_decap_8 FILLER_53_1289 ();
 sg13g2_decap_4 FILLER_53_1296 ();
 sg13g2_fill_1 FILLER_53_1300 ();
 sg13g2_decap_4 FILLER_53_1305 ();
 sg13g2_fill_1 FILLER_53_1309 ();
 sg13g2_decap_8 FILLER_53_1315 ();
 sg13g2_decap_8 FILLER_53_1322 ();
 sg13g2_decap_4 FILLER_53_1329 ();
 sg13g2_fill_2 FILLER_53_1333 ();
 sg13g2_fill_2 FILLER_53_1341 ();
 sg13g2_decap_4 FILLER_53_1352 ();
 sg13g2_fill_1 FILLER_53_1385 ();
 sg13g2_decap_4 FILLER_53_1396 ();
 sg13g2_fill_1 FILLER_53_1400 ();
 sg13g2_fill_1 FILLER_53_1423 ();
 sg13g2_decap_8 FILLER_53_1429 ();
 sg13g2_fill_1 FILLER_53_1436 ();
 sg13g2_decap_8 FILLER_53_1461 ();
 sg13g2_fill_1 FILLER_53_1468 ();
 sg13g2_fill_1 FILLER_53_1476 ();
 sg13g2_fill_1 FILLER_53_1481 ();
 sg13g2_fill_1 FILLER_53_1491 ();
 sg13g2_fill_1 FILLER_53_1495 ();
 sg13g2_fill_2 FILLER_53_1503 ();
 sg13g2_fill_2 FILLER_53_1517 ();
 sg13g2_fill_1 FILLER_53_1554 ();
 sg13g2_fill_2 FILLER_53_1564 ();
 sg13g2_fill_2 FILLER_53_1614 ();
 sg13g2_decap_8 FILLER_53_1622 ();
 sg13g2_decap_4 FILLER_53_1629 ();
 sg13g2_fill_1 FILLER_53_1633 ();
 sg13g2_decap_4 FILLER_53_1637 ();
 sg13g2_fill_2 FILLER_53_1641 ();
 sg13g2_decap_8 FILLER_53_1658 ();
 sg13g2_decap_8 FILLER_53_1665 ();
 sg13g2_decap_8 FILLER_53_1672 ();
 sg13g2_decap_8 FILLER_53_1679 ();
 sg13g2_decap_8 FILLER_53_1686 ();
 sg13g2_fill_2 FILLER_53_1693 ();
 sg13g2_fill_2 FILLER_53_1699 ();
 sg13g2_decap_8 FILLER_53_1716 ();
 sg13g2_decap_8 FILLER_53_1723 ();
 sg13g2_decap_8 FILLER_53_1730 ();
 sg13g2_decap_8 FILLER_53_1737 ();
 sg13g2_decap_4 FILLER_53_1744 ();
 sg13g2_fill_1 FILLER_53_1748 ();
 sg13g2_decap_8 FILLER_53_1753 ();
 sg13g2_decap_8 FILLER_53_1760 ();
 sg13g2_decap_8 FILLER_53_1767 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_fill_2 FILLER_54_28 ();
 sg13g2_fill_1 FILLER_54_30 ();
 sg13g2_fill_2 FILLER_54_41 ();
 sg13g2_fill_2 FILLER_54_55 ();
 sg13g2_fill_2 FILLER_54_61 ();
 sg13g2_fill_1 FILLER_54_63 ();
 sg13g2_fill_2 FILLER_54_69 ();
 sg13g2_fill_1 FILLER_54_71 ();
 sg13g2_decap_4 FILLER_54_82 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_106 ();
 sg13g2_decap_8 FILLER_54_113 ();
 sg13g2_decap_8 FILLER_54_120 ();
 sg13g2_decap_8 FILLER_54_127 ();
 sg13g2_decap_8 FILLER_54_134 ();
 sg13g2_decap_8 FILLER_54_141 ();
 sg13g2_fill_1 FILLER_54_148 ();
 sg13g2_fill_2 FILLER_54_159 ();
 sg13g2_decap_8 FILLER_54_174 ();
 sg13g2_decap_4 FILLER_54_181 ();
 sg13g2_fill_1 FILLER_54_185 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_fill_2 FILLER_54_219 ();
 sg13g2_decap_8 FILLER_54_226 ();
 sg13g2_fill_2 FILLER_54_233 ();
 sg13g2_decap_8 FILLER_54_250 ();
 sg13g2_decap_8 FILLER_54_257 ();
 sg13g2_decap_8 FILLER_54_264 ();
 sg13g2_decap_8 FILLER_54_271 ();
 sg13g2_fill_1 FILLER_54_278 ();
 sg13g2_fill_2 FILLER_54_299 ();
 sg13g2_fill_2 FILLER_54_306 ();
 sg13g2_decap_8 FILLER_54_313 ();
 sg13g2_decap_8 FILLER_54_337 ();
 sg13g2_decap_8 FILLER_54_349 ();
 sg13g2_decap_4 FILLER_54_356 ();
 sg13g2_fill_2 FILLER_54_360 ();
 sg13g2_fill_2 FILLER_54_395 ();
 sg13g2_fill_1 FILLER_54_397 ();
 sg13g2_decap_4 FILLER_54_403 ();
 sg13g2_decap_4 FILLER_54_411 ();
 sg13g2_decap_4 FILLER_54_420 ();
 sg13g2_decap_8 FILLER_54_428 ();
 sg13g2_decap_4 FILLER_54_435 ();
 sg13g2_decap_8 FILLER_54_453 ();
 sg13g2_decap_8 FILLER_54_460 ();
 sg13g2_fill_2 FILLER_54_467 ();
 sg13g2_decap_8 FILLER_54_475 ();
 sg13g2_decap_8 FILLER_54_497 ();
 sg13g2_decap_4 FILLER_54_504 ();
 sg13g2_fill_2 FILLER_54_534 ();
 sg13g2_fill_1 FILLER_54_536 ();
 sg13g2_decap_8 FILLER_54_541 ();
 sg13g2_decap_8 FILLER_54_624 ();
 sg13g2_fill_2 FILLER_54_631 ();
 sg13g2_fill_1 FILLER_54_633 ();
 sg13g2_decap_8 FILLER_54_638 ();
 sg13g2_decap_8 FILLER_54_645 ();
 sg13g2_decap_8 FILLER_54_652 ();
 sg13g2_decap_8 FILLER_54_659 ();
 sg13g2_decap_8 FILLER_54_666 ();
 sg13g2_decap_8 FILLER_54_673 ();
 sg13g2_decap_8 FILLER_54_680 ();
 sg13g2_decap_8 FILLER_54_687 ();
 sg13g2_fill_2 FILLER_54_694 ();
 sg13g2_fill_2 FILLER_54_704 ();
 sg13g2_fill_2 FILLER_54_710 ();
 sg13g2_fill_1 FILLER_54_712 ();
 sg13g2_decap_8 FILLER_54_721 ();
 sg13g2_fill_2 FILLER_54_728 ();
 sg13g2_fill_1 FILLER_54_734 ();
 sg13g2_fill_1 FILLER_54_774 ();
 sg13g2_decap_8 FILLER_54_788 ();
 sg13g2_decap_4 FILLER_54_795 ();
 sg13g2_fill_1 FILLER_54_803 ();
 sg13g2_decap_8 FILLER_54_808 ();
 sg13g2_fill_1 FILLER_54_818 ();
 sg13g2_decap_8 FILLER_54_845 ();
 sg13g2_fill_2 FILLER_54_852 ();
 sg13g2_fill_1 FILLER_54_869 ();
 sg13g2_decap_8 FILLER_54_875 ();
 sg13g2_decap_8 FILLER_54_882 ();
 sg13g2_decap_8 FILLER_54_889 ();
 sg13g2_decap_8 FILLER_54_896 ();
 sg13g2_decap_8 FILLER_54_912 ();
 sg13g2_decap_8 FILLER_54_919 ();
 sg13g2_decap_8 FILLER_54_926 ();
 sg13g2_fill_1 FILLER_54_933 ();
 sg13g2_decap_8 FILLER_54_938 ();
 sg13g2_decap_8 FILLER_54_945 ();
 sg13g2_decap_8 FILLER_54_961 ();
 sg13g2_fill_1 FILLER_54_968 ();
 sg13g2_fill_2 FILLER_54_973 ();
 sg13g2_fill_1 FILLER_54_975 ();
 sg13g2_decap_4 FILLER_54_1008 ();
 sg13g2_decap_4 FILLER_54_1017 ();
 sg13g2_fill_1 FILLER_54_1021 ();
 sg13g2_decap_8 FILLER_54_1027 ();
 sg13g2_decap_8 FILLER_54_1034 ();
 sg13g2_decap_8 FILLER_54_1041 ();
 sg13g2_decap_8 FILLER_54_1048 ();
 sg13g2_decap_8 FILLER_54_1055 ();
 sg13g2_decap_8 FILLER_54_1062 ();
 sg13g2_decap_8 FILLER_54_1069 ();
 sg13g2_decap_8 FILLER_54_1076 ();
 sg13g2_decap_4 FILLER_54_1083 ();
 sg13g2_fill_1 FILLER_54_1087 ();
 sg13g2_decap_8 FILLER_54_1118 ();
 sg13g2_decap_4 FILLER_54_1125 ();
 sg13g2_fill_2 FILLER_54_1129 ();
 sg13g2_decap_8 FILLER_54_1157 ();
 sg13g2_decap_8 FILLER_54_1190 ();
 sg13g2_decap_4 FILLER_54_1197 ();
 sg13g2_decap_8 FILLER_54_1207 ();
 sg13g2_decap_8 FILLER_54_1214 ();
 sg13g2_decap_8 FILLER_54_1221 ();
 sg13g2_decap_4 FILLER_54_1228 ();
 sg13g2_fill_2 FILLER_54_1232 ();
 sg13g2_decap_8 FILLER_54_1260 ();
 sg13g2_decap_8 FILLER_54_1267 ();
 sg13g2_decap_8 FILLER_54_1274 ();
 sg13g2_fill_1 FILLER_54_1281 ();
 sg13g2_decap_8 FILLER_54_1286 ();
 sg13g2_decap_8 FILLER_54_1293 ();
 sg13g2_decap_4 FILLER_54_1300 ();
 sg13g2_fill_2 FILLER_54_1304 ();
 sg13g2_decap_8 FILLER_54_1319 ();
 sg13g2_decap_8 FILLER_54_1326 ();
 sg13g2_fill_1 FILLER_54_1333 ();
 sg13g2_decap_8 FILLER_54_1346 ();
 sg13g2_decap_8 FILLER_54_1353 ();
 sg13g2_fill_2 FILLER_54_1360 ();
 sg13g2_fill_1 FILLER_54_1362 ();
 sg13g2_decap_8 FILLER_54_1367 ();
 sg13g2_fill_2 FILLER_54_1374 ();
 sg13g2_decap_8 FILLER_54_1381 ();
 sg13g2_fill_2 FILLER_54_1388 ();
 sg13g2_fill_1 FILLER_54_1390 ();
 sg13g2_decap_8 FILLER_54_1435 ();
 sg13g2_fill_1 FILLER_54_1442 ();
 sg13g2_fill_1 FILLER_54_1446 ();
 sg13g2_fill_2 FILLER_54_1478 ();
 sg13g2_fill_2 FILLER_54_1512 ();
 sg13g2_decap_4 FILLER_54_1547 ();
 sg13g2_fill_1 FILLER_54_1551 ();
 sg13g2_decap_4 FILLER_54_1557 ();
 sg13g2_fill_1 FILLER_54_1561 ();
 sg13g2_decap_8 FILLER_54_1574 ();
 sg13g2_decap_8 FILLER_54_1581 ();
 sg13g2_decap_4 FILLER_54_1588 ();
 sg13g2_decap_8 FILLER_54_1596 ();
 sg13g2_fill_1 FILLER_54_1603 ();
 sg13g2_fill_1 FILLER_54_1622 ();
 sg13g2_fill_2 FILLER_54_1628 ();
 sg13g2_decap_4 FILLER_54_1638 ();
 sg13g2_fill_1 FILLER_54_1642 ();
 sg13g2_decap_8 FILLER_54_1648 ();
 sg13g2_decap_4 FILLER_54_1655 ();
 sg13g2_fill_1 FILLER_54_1659 ();
 sg13g2_decap_4 FILLER_54_1668 ();
 sg13g2_fill_2 FILLER_54_1698 ();
 sg13g2_fill_1 FILLER_54_1700 ();
 sg13g2_decap_8 FILLER_54_1706 ();
 sg13g2_decap_8 FILLER_54_1713 ();
 sg13g2_decap_8 FILLER_54_1720 ();
 sg13g2_decap_8 FILLER_54_1727 ();
 sg13g2_decap_4 FILLER_54_1768 ();
 sg13g2_fill_2 FILLER_54_1772 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_4 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_25 ();
 sg13g2_fill_1 FILLER_55_30 ();
 sg13g2_fill_1 FILLER_55_41 ();
 sg13g2_fill_2 FILLER_55_47 ();
 sg13g2_fill_1 FILLER_55_49 ();
 sg13g2_decap_4 FILLER_55_55 ();
 sg13g2_fill_1 FILLER_55_59 ();
 sg13g2_decap_4 FILLER_55_65 ();
 sg13g2_fill_1 FILLER_55_69 ();
 sg13g2_fill_1 FILLER_55_75 ();
 sg13g2_decap_8 FILLER_55_82 ();
 sg13g2_fill_1 FILLER_55_89 ();
 sg13g2_decap_4 FILLER_55_97 ();
 sg13g2_fill_1 FILLER_55_101 ();
 sg13g2_decap_8 FILLER_55_107 ();
 sg13g2_decap_8 FILLER_55_114 ();
 sg13g2_decap_4 FILLER_55_121 ();
 sg13g2_decap_8 FILLER_55_130 ();
 sg13g2_fill_2 FILLER_55_137 ();
 sg13g2_fill_1 FILLER_55_139 ();
 sg13g2_decap_8 FILLER_55_145 ();
 sg13g2_fill_2 FILLER_55_152 ();
 sg13g2_fill_1 FILLER_55_154 ();
 sg13g2_fill_2 FILLER_55_164 ();
 sg13g2_fill_1 FILLER_55_166 ();
 sg13g2_decap_8 FILLER_55_172 ();
 sg13g2_decap_8 FILLER_55_179 ();
 sg13g2_decap_8 FILLER_55_186 ();
 sg13g2_decap_8 FILLER_55_193 ();
 sg13g2_decap_4 FILLER_55_200 ();
 sg13g2_decap_8 FILLER_55_208 ();
 sg13g2_decap_8 FILLER_55_215 ();
 sg13g2_decap_8 FILLER_55_222 ();
 sg13g2_decap_8 FILLER_55_229 ();
 sg13g2_decap_4 FILLER_55_236 ();
 sg13g2_fill_2 FILLER_55_240 ();
 sg13g2_decap_8 FILLER_55_268 ();
 sg13g2_decap_8 FILLER_55_275 ();
 sg13g2_decap_4 FILLER_55_282 ();
 sg13g2_fill_1 FILLER_55_286 ();
 sg13g2_fill_2 FILLER_55_296 ();
 sg13g2_fill_1 FILLER_55_298 ();
 sg13g2_decap_4 FILLER_55_304 ();
 sg13g2_decap_8 FILLER_55_317 ();
 sg13g2_decap_8 FILLER_55_324 ();
 sg13g2_fill_2 FILLER_55_331 ();
 sg13g2_decap_8 FILLER_55_338 ();
 sg13g2_decap_8 FILLER_55_345 ();
 sg13g2_decap_8 FILLER_55_352 ();
 sg13g2_decap_4 FILLER_55_359 ();
 sg13g2_decap_4 FILLER_55_369 ();
 sg13g2_decap_4 FILLER_55_381 ();
 sg13g2_decap_4 FILLER_55_389 ();
 sg13g2_fill_1 FILLER_55_402 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_55_430 ();
 sg13g2_decap_8 FILLER_55_437 ();
 sg13g2_decap_8 FILLER_55_444 ();
 sg13g2_decap_8 FILLER_55_451 ();
 sg13g2_decap_8 FILLER_55_458 ();
 sg13g2_fill_2 FILLER_55_465 ();
 sg13g2_fill_1 FILLER_55_472 ();
 sg13g2_decap_8 FILLER_55_492 ();
 sg13g2_decap_4 FILLER_55_499 ();
 sg13g2_fill_1 FILLER_55_503 ();
 sg13g2_decap_4 FILLER_55_509 ();
 sg13g2_fill_2 FILLER_55_517 ();
 sg13g2_decap_8 FILLER_55_524 ();
 sg13g2_decap_8 FILLER_55_531 ();
 sg13g2_fill_1 FILLER_55_538 ();
 sg13g2_decap_8 FILLER_55_543 ();
 sg13g2_decap_8 FILLER_55_550 ();
 sg13g2_decap_8 FILLER_55_557 ();
 sg13g2_fill_2 FILLER_55_564 ();
 sg13g2_decap_8 FILLER_55_570 ();
 sg13g2_decap_8 FILLER_55_577 ();
 sg13g2_decap_8 FILLER_55_587 ();
 sg13g2_decap_4 FILLER_55_594 ();
 sg13g2_fill_2 FILLER_55_598 ();
 sg13g2_decap_4 FILLER_55_604 ();
 sg13g2_fill_1 FILLER_55_608 ();
 sg13g2_decap_4 FILLER_55_612 ();
 sg13g2_fill_2 FILLER_55_616 ();
 sg13g2_decap_8 FILLER_55_624 ();
 sg13g2_decap_8 FILLER_55_631 ();
 sg13g2_decap_8 FILLER_55_638 ();
 sg13g2_fill_1 FILLER_55_645 ();
 sg13g2_decap_8 FILLER_55_651 ();
 sg13g2_fill_2 FILLER_55_658 ();
 sg13g2_decap_8 FILLER_55_689 ();
 sg13g2_decap_4 FILLER_55_696 ();
 sg13g2_fill_1 FILLER_55_700 ();
 sg13g2_decap_8 FILLER_55_706 ();
 sg13g2_decap_4 FILLER_55_718 ();
 sg13g2_fill_2 FILLER_55_722 ();
 sg13g2_decap_8 FILLER_55_728 ();
 sg13g2_decap_8 FILLER_55_735 ();
 sg13g2_decap_8 FILLER_55_747 ();
 sg13g2_fill_1 FILLER_55_754 ();
 sg13g2_fill_1 FILLER_55_763 ();
 sg13g2_fill_2 FILLER_55_772 ();
 sg13g2_fill_1 FILLER_55_774 ();
 sg13g2_decap_8 FILLER_55_779 ();
 sg13g2_fill_2 FILLER_55_786 ();
 sg13g2_fill_1 FILLER_55_788 ();
 sg13g2_decap_8 FILLER_55_829 ();
 sg13g2_decap_8 FILLER_55_836 ();
 sg13g2_decap_8 FILLER_55_843 ();
 sg13g2_decap_8 FILLER_55_850 ();
 sg13g2_decap_4 FILLER_55_857 ();
 sg13g2_decap_4 FILLER_55_866 ();
 sg13g2_decap_8 FILLER_55_877 ();
 sg13g2_fill_2 FILLER_55_884 ();
 sg13g2_fill_1 FILLER_55_886 ();
 sg13g2_fill_2 FILLER_55_892 ();
 sg13g2_fill_1 FILLER_55_894 ();
 sg13g2_decap_8 FILLER_55_908 ();
 sg13g2_decap_8 FILLER_55_915 ();
 sg13g2_decap_8 FILLER_55_922 ();
 sg13g2_decap_8 FILLER_55_929 ();
 sg13g2_decap_8 FILLER_55_936 ();
 sg13g2_decap_8 FILLER_55_943 ();
 sg13g2_decap_8 FILLER_55_950 ();
 sg13g2_decap_4 FILLER_55_957 ();
 sg13g2_fill_2 FILLER_55_961 ();
 sg13g2_fill_2 FILLER_55_973 ();
 sg13g2_fill_1 FILLER_55_975 ();
 sg13g2_fill_2 FILLER_55_979 ();
 sg13g2_fill_1 FILLER_55_981 ();
 sg13g2_fill_2 FILLER_55_995 ();
 sg13g2_decap_8 FILLER_55_1009 ();
 sg13g2_decap_4 FILLER_55_1016 ();
 sg13g2_fill_1 FILLER_55_1020 ();
 sg13g2_decap_8 FILLER_55_1029 ();
 sg13g2_decap_4 FILLER_55_1036 ();
 sg13g2_decap_4 FILLER_55_1045 ();
 sg13g2_fill_1 FILLER_55_1049 ();
 sg13g2_decap_8 FILLER_55_1054 ();
 sg13g2_decap_8 FILLER_55_1061 ();
 sg13g2_decap_8 FILLER_55_1068 ();
 sg13g2_decap_8 FILLER_55_1075 ();
 sg13g2_decap_8 FILLER_55_1082 ();
 sg13g2_decap_4 FILLER_55_1089 ();
 sg13g2_fill_1 FILLER_55_1093 ();
 sg13g2_decap_8 FILLER_55_1098 ();
 sg13g2_decap_8 FILLER_55_1105 ();
 sg13g2_decap_8 FILLER_55_1112 ();
 sg13g2_decap_8 FILLER_55_1119 ();
 sg13g2_decap_8 FILLER_55_1126 ();
 sg13g2_decap_8 FILLER_55_1133 ();
 sg13g2_decap_8 FILLER_55_1140 ();
 sg13g2_decap_8 FILLER_55_1147 ();
 sg13g2_decap_8 FILLER_55_1154 ();
 sg13g2_decap_8 FILLER_55_1165 ();
 sg13g2_decap_8 FILLER_55_1172 ();
 sg13g2_fill_2 FILLER_55_1179 ();
 sg13g2_decap_8 FILLER_55_1195 ();
 sg13g2_decap_4 FILLER_55_1207 ();
 sg13g2_fill_2 FILLER_55_1211 ();
 sg13g2_decap_8 FILLER_55_1221 ();
 sg13g2_decap_8 FILLER_55_1228 ();
 sg13g2_decap_4 FILLER_55_1235 ();
 sg13g2_fill_2 FILLER_55_1239 ();
 sg13g2_decap_8 FILLER_55_1245 ();
 sg13g2_decap_4 FILLER_55_1252 ();
 sg13g2_fill_1 FILLER_55_1256 ();
 sg13g2_decap_4 FILLER_55_1260 ();
 sg13g2_fill_1 FILLER_55_1264 ();
 sg13g2_decap_8 FILLER_55_1303 ();
 sg13g2_fill_1 FILLER_55_1310 ();
 sg13g2_fill_1 FILLER_55_1319 ();
 sg13g2_decap_4 FILLER_55_1323 ();
 sg13g2_decap_8 FILLER_55_1338 ();
 sg13g2_decap_8 FILLER_55_1345 ();
 sg13g2_decap_8 FILLER_55_1352 ();
 sg13g2_decap_8 FILLER_55_1359 ();
 sg13g2_decap_4 FILLER_55_1366 ();
 sg13g2_decap_8 FILLER_55_1374 ();
 sg13g2_decap_4 FILLER_55_1381 ();
 sg13g2_fill_1 FILLER_55_1389 ();
 sg13g2_decap_8 FILLER_55_1399 ();
 sg13g2_decap_8 FILLER_55_1406 ();
 sg13g2_decap_8 FILLER_55_1413 ();
 sg13g2_decap_8 FILLER_55_1420 ();
 sg13g2_decap_8 FILLER_55_1427 ();
 sg13g2_fill_1 FILLER_55_1434 ();
 sg13g2_decap_8 FILLER_55_1440 ();
 sg13g2_decap_8 FILLER_55_1447 ();
 sg13g2_decap_4 FILLER_55_1454 ();
 sg13g2_fill_2 FILLER_55_1458 ();
 sg13g2_decap_8 FILLER_55_1465 ();
 sg13g2_fill_2 FILLER_55_1472 ();
 sg13g2_decap_8 FILLER_55_1478 ();
 sg13g2_fill_1 FILLER_55_1485 ();
 sg13g2_decap_4 FILLER_55_1512 ();
 sg13g2_decap_8 FILLER_55_1521 ();
 sg13g2_decap_4 FILLER_55_1528 ();
 sg13g2_fill_1 FILLER_55_1539 ();
 sg13g2_fill_1 FILLER_55_1546 ();
 sg13g2_fill_2 FILLER_55_1556 ();
 sg13g2_fill_2 FILLER_55_1563 ();
 sg13g2_decap_4 FILLER_55_1579 ();
 sg13g2_fill_1 FILLER_55_1583 ();
 sg13g2_decap_8 FILLER_55_1589 ();
 sg13g2_decap_8 FILLER_55_1596 ();
 sg13g2_decap_8 FILLER_55_1603 ();
 sg13g2_fill_2 FILLER_55_1610 ();
 sg13g2_fill_1 FILLER_55_1612 ();
 sg13g2_decap_4 FILLER_55_1621 ();
 sg13g2_fill_1 FILLER_55_1625 ();
 sg13g2_decap_8 FILLER_55_1633 ();
 sg13g2_decap_8 FILLER_55_1640 ();
 sg13g2_decap_8 FILLER_55_1647 ();
 sg13g2_decap_8 FILLER_55_1654 ();
 sg13g2_decap_4 FILLER_55_1661 ();
 sg13g2_fill_2 FILLER_55_1665 ();
 sg13g2_decap_4 FILLER_55_1672 ();
 sg13g2_fill_1 FILLER_55_1676 ();
 sg13g2_decap_8 FILLER_55_1681 ();
 sg13g2_fill_1 FILLER_55_1688 ();
 sg13g2_decap_8 FILLER_55_1694 ();
 sg13g2_decap_8 FILLER_55_1701 ();
 sg13g2_decap_4 FILLER_55_1732 ();
 sg13g2_fill_1 FILLER_55_1736 ();
 sg13g2_decap_4 FILLER_55_1742 ();
 sg13g2_fill_1 FILLER_55_1746 ();
 sg13g2_decap_8 FILLER_55_1751 ();
 sg13g2_decap_8 FILLER_55_1758 ();
 sg13g2_decap_8 FILLER_55_1765 ();
 sg13g2_fill_2 FILLER_55_1772 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_fill_2 FILLER_56_28 ();
 sg13g2_fill_1 FILLER_56_30 ();
 sg13g2_fill_2 FILLER_56_36 ();
 sg13g2_fill_1 FILLER_56_38 ();
 sg13g2_decap_4 FILLER_56_43 ();
 sg13g2_fill_1 FILLER_56_47 ();
 sg13g2_decap_8 FILLER_56_62 ();
 sg13g2_decap_8 FILLER_56_69 ();
 sg13g2_fill_1 FILLER_56_76 ();
 sg13g2_fill_2 FILLER_56_86 ();
 sg13g2_fill_1 FILLER_56_88 ();
 sg13g2_fill_1 FILLER_56_100 ();
 sg13g2_fill_1 FILLER_56_106 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_fill_1 FILLER_56_125 ();
 sg13g2_fill_2 FILLER_56_131 ();
 sg13g2_fill_1 FILLER_56_146 ();
 sg13g2_fill_2 FILLER_56_152 ();
 sg13g2_decap_8 FILLER_56_178 ();
 sg13g2_decap_8 FILLER_56_190 ();
 sg13g2_fill_2 FILLER_56_197 ();
 sg13g2_decap_8 FILLER_56_209 ();
 sg13g2_fill_1 FILLER_56_216 ();
 sg13g2_decap_8 FILLER_56_230 ();
 sg13g2_decap_8 FILLER_56_237 ();
 sg13g2_fill_2 FILLER_56_244 ();
 sg13g2_fill_1 FILLER_56_246 ();
 sg13g2_fill_1 FILLER_56_250 ();
 sg13g2_decap_8 FILLER_56_255 ();
 sg13g2_fill_2 FILLER_56_262 ();
 sg13g2_decap_8 FILLER_56_274 ();
 sg13g2_decap_8 FILLER_56_286 ();
 sg13g2_decap_8 FILLER_56_293 ();
 sg13g2_decap_8 FILLER_56_300 ();
 sg13g2_decap_4 FILLER_56_307 ();
 sg13g2_fill_1 FILLER_56_311 ();
 sg13g2_fill_1 FILLER_56_320 ();
 sg13g2_decap_8 FILLER_56_325 ();
 sg13g2_fill_1 FILLER_56_332 ();
 sg13g2_decap_4 FILLER_56_338 ();
 sg13g2_fill_1 FILLER_56_342 ();
 sg13g2_decap_8 FILLER_56_366 ();
 sg13g2_decap_4 FILLER_56_373 ();
 sg13g2_fill_2 FILLER_56_377 ();
 sg13g2_decap_8 FILLER_56_383 ();
 sg13g2_decap_8 FILLER_56_390 ();
 sg13g2_decap_8 FILLER_56_397 ();
 sg13g2_decap_8 FILLER_56_404 ();
 sg13g2_decap_8 FILLER_56_411 ();
 sg13g2_decap_8 FILLER_56_418 ();
 sg13g2_fill_2 FILLER_56_425 ();
 sg13g2_decap_4 FILLER_56_440 ();
 sg13g2_fill_1 FILLER_56_444 ();
 sg13g2_decap_8 FILLER_56_451 ();
 sg13g2_fill_2 FILLER_56_467 ();
 sg13g2_fill_1 FILLER_56_469 ();
 sg13g2_decap_4 FILLER_56_477 ();
 sg13g2_fill_1 FILLER_56_481 ();
 sg13g2_decap_8 FILLER_56_497 ();
 sg13g2_decap_8 FILLER_56_504 ();
 sg13g2_decap_8 FILLER_56_511 ();
 sg13g2_decap_8 FILLER_56_518 ();
 sg13g2_fill_2 FILLER_56_525 ();
 sg13g2_fill_1 FILLER_56_527 ();
 sg13g2_decap_8 FILLER_56_532 ();
 sg13g2_decap_8 FILLER_56_539 ();
 sg13g2_fill_1 FILLER_56_546 ();
 sg13g2_decap_8 FILLER_56_551 ();
 sg13g2_fill_2 FILLER_56_566 ();
 sg13g2_decap_8 FILLER_56_576 ();
 sg13g2_decap_8 FILLER_56_583 ();
 sg13g2_decap_8 FILLER_56_590 ();
 sg13g2_fill_1 FILLER_56_597 ();
 sg13g2_fill_2 FILLER_56_603 ();
 sg13g2_decap_8 FILLER_56_656 ();
 sg13g2_fill_2 FILLER_56_663 ();
 sg13g2_fill_1 FILLER_56_665 ();
 sg13g2_decap_8 FILLER_56_670 ();
 sg13g2_decap_8 FILLER_56_677 ();
 sg13g2_decap_8 FILLER_56_684 ();
 sg13g2_fill_1 FILLER_56_691 ();
 sg13g2_decap_8 FILLER_56_696 ();
 sg13g2_fill_2 FILLER_56_703 ();
 sg13g2_decap_4 FILLER_56_710 ();
 sg13g2_fill_2 FILLER_56_714 ();
 sg13g2_decap_8 FILLER_56_731 ();
 sg13g2_decap_8 FILLER_56_738 ();
 sg13g2_decap_8 FILLER_56_745 ();
 sg13g2_decap_4 FILLER_56_752 ();
 sg13g2_decap_8 FILLER_56_769 ();
 sg13g2_decap_8 FILLER_56_776 ();
 sg13g2_decap_8 FILLER_56_783 ();
 sg13g2_decap_4 FILLER_56_790 ();
 sg13g2_fill_1 FILLER_56_794 ();
 sg13g2_fill_1 FILLER_56_802 ();
 sg13g2_decap_4 FILLER_56_826 ();
 sg13g2_fill_2 FILLER_56_830 ();
 sg13g2_decap_8 FILLER_56_845 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_decap_8 FILLER_56_859 ();
 sg13g2_fill_1 FILLER_56_866 ();
 sg13g2_decap_8 FILLER_56_872 ();
 sg13g2_decap_8 FILLER_56_879 ();
 sg13g2_decap_4 FILLER_56_886 ();
 sg13g2_fill_1 FILLER_56_898 ();
 sg13g2_decap_8 FILLER_56_903 ();
 sg13g2_fill_2 FILLER_56_910 ();
 sg13g2_fill_1 FILLER_56_912 ();
 sg13g2_decap_8 FILLER_56_917 ();
 sg13g2_decap_8 FILLER_56_924 ();
 sg13g2_decap_8 FILLER_56_931 ();
 sg13g2_fill_1 FILLER_56_943 ();
 sg13g2_decap_8 FILLER_56_949 ();
 sg13g2_decap_8 FILLER_56_956 ();
 sg13g2_decap_8 FILLER_56_963 ();
 sg13g2_decap_8 FILLER_56_970 ();
 sg13g2_decap_8 FILLER_56_977 ();
 sg13g2_decap_8 FILLER_56_984 ();
 sg13g2_decap_4 FILLER_56_991 ();
 sg13g2_fill_1 FILLER_56_995 ();
 sg13g2_decap_8 FILLER_56_1006 ();
 sg13g2_decap_4 FILLER_56_1013 ();
 sg13g2_fill_1 FILLER_56_1017 ();
 sg13g2_fill_1 FILLER_56_1027 ();
 sg13g2_decap_8 FILLER_56_1032 ();
 sg13g2_fill_2 FILLER_56_1069 ();
 sg13g2_fill_1 FILLER_56_1071 ();
 sg13g2_decap_8 FILLER_56_1077 ();
 sg13g2_decap_4 FILLER_56_1084 ();
 sg13g2_fill_1 FILLER_56_1088 ();
 sg13g2_decap_8 FILLER_56_1115 ();
 sg13g2_decap_8 FILLER_56_1122 ();
 sg13g2_decap_4 FILLER_56_1129 ();
 sg13g2_fill_1 FILLER_56_1133 ();
 sg13g2_decap_8 FILLER_56_1137 ();
 sg13g2_decap_8 FILLER_56_1148 ();
 sg13g2_fill_1 FILLER_56_1155 ();
 sg13g2_decap_8 FILLER_56_1211 ();
 sg13g2_decap_8 FILLER_56_1226 ();
 sg13g2_decap_4 FILLER_56_1237 ();
 sg13g2_fill_1 FILLER_56_1247 ();
 sg13g2_fill_1 FILLER_56_1254 ();
 sg13g2_decap_8 FILLER_56_1259 ();
 sg13g2_decap_8 FILLER_56_1266 ();
 sg13g2_decap_8 FILLER_56_1273 ();
 sg13g2_fill_1 FILLER_56_1280 ();
 sg13g2_decap_4 FILLER_56_1285 ();
 sg13g2_fill_2 FILLER_56_1289 ();
 sg13g2_decap_4 FILLER_56_1295 ();
 sg13g2_fill_2 FILLER_56_1299 ();
 sg13g2_decap_8 FILLER_56_1316 ();
 sg13g2_decap_4 FILLER_56_1323 ();
 sg13g2_decap_8 FILLER_56_1348 ();
 sg13g2_decap_8 FILLER_56_1355 ();
 sg13g2_decap_4 FILLER_56_1362 ();
 sg13g2_decap_8 FILLER_56_1395 ();
 sg13g2_decap_8 FILLER_56_1402 ();
 sg13g2_decap_4 FILLER_56_1409 ();
 sg13g2_fill_2 FILLER_56_1413 ();
 sg13g2_decap_8 FILLER_56_1419 ();
 sg13g2_decap_8 FILLER_56_1426 ();
 sg13g2_decap_8 FILLER_56_1433 ();
 sg13g2_decap_8 FILLER_56_1440 ();
 sg13g2_decap_8 FILLER_56_1447 ();
 sg13g2_fill_2 FILLER_56_1454 ();
 sg13g2_fill_1 FILLER_56_1456 ();
 sg13g2_decap_4 FILLER_56_1461 ();
 sg13g2_decap_8 FILLER_56_1469 ();
 sg13g2_decap_8 FILLER_56_1476 ();
 sg13g2_decap_4 FILLER_56_1495 ();
 sg13g2_fill_1 FILLER_56_1499 ();
 sg13g2_decap_8 FILLER_56_1503 ();
 sg13g2_decap_8 FILLER_56_1510 ();
 sg13g2_decap_8 FILLER_56_1517 ();
 sg13g2_decap_4 FILLER_56_1524 ();
 sg13g2_fill_1 FILLER_56_1545 ();
 sg13g2_fill_1 FILLER_56_1556 ();
 sg13g2_fill_2 FILLER_56_1565 ();
 sg13g2_decap_8 FILLER_56_1572 ();
 sg13g2_fill_2 FILLER_56_1579 ();
 sg13g2_decap_8 FILLER_56_1600 ();
 sg13g2_fill_2 FILLER_56_1607 ();
 sg13g2_decap_8 FILLER_56_1621 ();
 sg13g2_decap_8 FILLER_56_1628 ();
 sg13g2_decap_8 FILLER_56_1635 ();
 sg13g2_decap_8 FILLER_56_1642 ();
 sg13g2_decap_8 FILLER_56_1649 ();
 sg13g2_decap_8 FILLER_56_1656 ();
 sg13g2_fill_2 FILLER_56_1663 ();
 sg13g2_fill_1 FILLER_56_1665 ();
 sg13g2_decap_8 FILLER_56_1670 ();
 sg13g2_decap_4 FILLER_56_1677 ();
 sg13g2_fill_1 FILLER_56_1681 ();
 sg13g2_fill_1 FILLER_56_1687 ();
 sg13g2_decap_8 FILLER_56_1694 ();
 sg13g2_decap_4 FILLER_56_1701 ();
 sg13g2_fill_1 FILLER_56_1705 ();
 sg13g2_decap_8 FILLER_56_1709 ();
 sg13g2_fill_2 FILLER_56_1716 ();
 sg13g2_fill_1 FILLER_56_1718 ();
 sg13g2_fill_2 FILLER_56_1737 ();
 sg13g2_fill_1 FILLER_56_1739 ();
 sg13g2_decap_8 FILLER_56_1766 ();
 sg13g2_fill_1 FILLER_56_1773 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_37 ();
 sg13g2_decap_4 FILLER_57_44 ();
 sg13g2_fill_2 FILLER_57_48 ();
 sg13g2_decap_4 FILLER_57_55 ();
 sg13g2_fill_1 FILLER_57_64 ();
 sg13g2_fill_1 FILLER_57_69 ();
 sg13g2_decap_4 FILLER_57_90 ();
 sg13g2_fill_2 FILLER_57_94 ();
 sg13g2_fill_2 FILLER_57_101 ();
 sg13g2_fill_1 FILLER_57_103 ();
 sg13g2_decap_8 FILLER_57_109 ();
 sg13g2_decap_8 FILLER_57_116 ();
 sg13g2_fill_2 FILLER_57_123 ();
 sg13g2_decap_8 FILLER_57_129 ();
 sg13g2_decap_4 FILLER_57_136 ();
 sg13g2_decap_8 FILLER_57_146 ();
 sg13g2_decap_4 FILLER_57_159 ();
 sg13g2_fill_1 FILLER_57_163 ();
 sg13g2_fill_2 FILLER_57_176 ();
 sg13g2_decap_8 FILLER_57_187 ();
 sg13g2_fill_2 FILLER_57_194 ();
 sg13g2_decap_8 FILLER_57_201 ();
 sg13g2_decap_4 FILLER_57_208 ();
 sg13g2_decap_4 FILLER_57_216 ();
 sg13g2_fill_2 FILLER_57_229 ();
 sg13g2_fill_1 FILLER_57_231 ();
 sg13g2_decap_4 FILLER_57_237 ();
 sg13g2_fill_2 FILLER_57_241 ();
 sg13g2_decap_8 FILLER_57_249 ();
 sg13g2_fill_2 FILLER_57_256 ();
 sg13g2_decap_8 FILLER_57_269 ();
 sg13g2_fill_1 FILLER_57_276 ();
 sg13g2_fill_2 FILLER_57_281 ();
 sg13g2_fill_1 FILLER_57_283 ();
 sg13g2_fill_2 FILLER_57_302 ();
 sg13g2_decap_4 FILLER_57_316 ();
 sg13g2_decap_4 FILLER_57_331 ();
 sg13g2_fill_2 FILLER_57_335 ();
 sg13g2_fill_1 FILLER_57_342 ();
 sg13g2_decap_8 FILLER_57_355 ();
 sg13g2_decap_8 FILLER_57_362 ();
 sg13g2_fill_2 FILLER_57_374 ();
 sg13g2_fill_2 FILLER_57_381 ();
 sg13g2_fill_2 FILLER_57_387 ();
 sg13g2_fill_1 FILLER_57_389 ();
 sg13g2_fill_2 FILLER_57_395 ();
 sg13g2_fill_2 FILLER_57_403 ();
 sg13g2_fill_1 FILLER_57_405 ();
 sg13g2_decap_8 FILLER_57_417 ();
 sg13g2_decap_8 FILLER_57_424 ();
 sg13g2_decap_8 FILLER_57_431 ();
 sg13g2_decap_4 FILLER_57_438 ();
 sg13g2_fill_1 FILLER_57_442 ();
 sg13g2_decap_8 FILLER_57_448 ();
 sg13g2_decap_8 FILLER_57_455 ();
 sg13g2_decap_8 FILLER_57_462 ();
 sg13g2_decap_8 FILLER_57_469 ();
 sg13g2_decap_8 FILLER_57_476 ();
 sg13g2_decap_8 FILLER_57_483 ();
 sg13g2_fill_2 FILLER_57_490 ();
 sg13g2_fill_1 FILLER_57_492 ();
 sg13g2_fill_1 FILLER_57_516 ();
 sg13g2_fill_1 FILLER_57_520 ();
 sg13g2_decap_4 FILLER_57_547 ();
 sg13g2_fill_1 FILLER_57_591 ();
 sg13g2_decap_8 FILLER_57_641 ();
 sg13g2_decap_4 FILLER_57_648 ();
 sg13g2_fill_2 FILLER_57_652 ();
 sg13g2_decap_8 FILLER_57_671 ();
 sg13g2_decap_8 FILLER_57_678 ();
 sg13g2_decap_8 FILLER_57_685 ();
 sg13g2_decap_4 FILLER_57_692 ();
 sg13g2_fill_1 FILLER_57_696 ();
 sg13g2_fill_2 FILLER_57_721 ();
 sg13g2_fill_2 FILLER_57_729 ();
 sg13g2_fill_1 FILLER_57_731 ();
 sg13g2_fill_2 FILLER_57_740 ();
 sg13g2_fill_1 FILLER_57_742 ();
 sg13g2_decap_8 FILLER_57_751 ();
 sg13g2_decap_8 FILLER_57_758 ();
 sg13g2_decap_8 FILLER_57_765 ();
 sg13g2_fill_1 FILLER_57_772 ();
 sg13g2_decap_4 FILLER_57_777 ();
 sg13g2_fill_1 FILLER_57_784 ();
 sg13g2_decap_4 FILLER_57_820 ();
 sg13g2_fill_1 FILLER_57_824 ();
 sg13g2_fill_1 FILLER_57_830 ();
 sg13g2_decap_4 FILLER_57_860 ();
 sg13g2_fill_2 FILLER_57_864 ();
 sg13g2_fill_1 FILLER_57_892 ();
 sg13g2_fill_2 FILLER_57_919 ();
 sg13g2_fill_1 FILLER_57_921 ();
 sg13g2_decap_8 FILLER_57_926 ();
 sg13g2_fill_1 FILLER_57_933 ();
 sg13g2_decap_8 FILLER_57_956 ();
 sg13g2_fill_2 FILLER_57_963 ();
 sg13g2_fill_1 FILLER_57_965 ();
 sg13g2_decap_8 FILLER_57_974 ();
 sg13g2_decap_8 FILLER_57_981 ();
 sg13g2_decap_8 FILLER_57_988 ();
 sg13g2_decap_4 FILLER_57_995 ();
 sg13g2_fill_1 FILLER_57_1004 ();
 sg13g2_decap_8 FILLER_57_1009 ();
 sg13g2_decap_8 FILLER_57_1016 ();
 sg13g2_decap_4 FILLER_57_1023 ();
 sg13g2_decap_8 FILLER_57_1032 ();
 sg13g2_decap_8 FILLER_57_1039 ();
 sg13g2_decap_4 FILLER_57_1046 ();
 sg13g2_fill_2 FILLER_57_1050 ();
 sg13g2_decap_4 FILLER_57_1056 ();
 sg13g2_fill_1 FILLER_57_1060 ();
 sg13g2_decap_8 FILLER_57_1066 ();
 sg13g2_decap_4 FILLER_57_1073 ();
 sg13g2_fill_2 FILLER_57_1077 ();
 sg13g2_fill_2 FILLER_57_1096 ();
 sg13g2_fill_1 FILLER_57_1098 ();
 sg13g2_decap_4 FILLER_57_1103 ();
 sg13g2_fill_2 FILLER_57_1107 ();
 sg13g2_decap_8 FILLER_57_1113 ();
 sg13g2_decap_8 FILLER_57_1120 ();
 sg13g2_fill_1 FILLER_57_1127 ();
 sg13g2_fill_1 FILLER_57_1137 ();
 sg13g2_fill_1 FILLER_57_1164 ();
 sg13g2_fill_1 FILLER_57_1187 ();
 sg13g2_decap_4 FILLER_57_1193 ();
 sg13g2_fill_1 FILLER_57_1201 ();
 sg13g2_decap_4 FILLER_57_1206 ();
 sg13g2_decap_8 FILLER_57_1223 ();
 sg13g2_decap_8 FILLER_57_1230 ();
 sg13g2_decap_8 FILLER_57_1237 ();
 sg13g2_decap_8 FILLER_57_1244 ();
 sg13g2_decap_8 FILLER_57_1251 ();
 sg13g2_decap_8 FILLER_57_1258 ();
 sg13g2_fill_2 FILLER_57_1265 ();
 sg13g2_fill_1 FILLER_57_1267 ();
 sg13g2_decap_8 FILLER_57_1273 ();
 sg13g2_decap_8 FILLER_57_1280 ();
 sg13g2_decap_4 FILLER_57_1287 ();
 sg13g2_decap_8 FILLER_57_1301 ();
 sg13g2_decap_8 FILLER_57_1308 ();
 sg13g2_decap_8 FILLER_57_1315 ();
 sg13g2_decap_8 FILLER_57_1322 ();
 sg13g2_decap_8 FILLER_57_1329 ();
 sg13g2_decap_8 FILLER_57_1336 ();
 sg13g2_decap_8 FILLER_57_1343 ();
 sg13g2_decap_8 FILLER_57_1350 ();
 sg13g2_decap_8 FILLER_57_1357 ();
 sg13g2_decap_8 FILLER_57_1364 ();
 sg13g2_decap_8 FILLER_57_1379 ();
 sg13g2_decap_8 FILLER_57_1386 ();
 sg13g2_decap_8 FILLER_57_1393 ();
 sg13g2_decap_8 FILLER_57_1400 ();
 sg13g2_fill_2 FILLER_57_1407 ();
 sg13g2_fill_2 FILLER_57_1435 ();
 sg13g2_fill_1 FILLER_57_1437 ();
 sg13g2_decap_8 FILLER_57_1441 ();
 sg13g2_fill_1 FILLER_57_1448 ();
 sg13g2_fill_1 FILLER_57_1465 ();
 sg13g2_decap_4 FILLER_57_1491 ();
 sg13g2_fill_1 FILLER_57_1495 ();
 sg13g2_decap_4 FILLER_57_1506 ();
 sg13g2_fill_1 FILLER_57_1510 ();
 sg13g2_decap_8 FILLER_57_1515 ();
 sg13g2_decap_4 FILLER_57_1528 ();
 sg13g2_fill_1 FILLER_57_1532 ();
 sg13g2_decap_8 FILLER_57_1537 ();
 sg13g2_fill_1 FILLER_57_1560 ();
 sg13g2_fill_2 FILLER_57_1575 ();
 sg13g2_fill_1 FILLER_57_1577 ();
 sg13g2_decap_8 FILLER_57_1583 ();
 sg13g2_decap_8 FILLER_57_1590 ();
 sg13g2_fill_2 FILLER_57_1597 ();
 sg13g2_decap_4 FILLER_57_1605 ();
 sg13g2_fill_1 FILLER_57_1616 ();
 sg13g2_decap_4 FILLER_57_1623 ();
 sg13g2_fill_2 FILLER_57_1627 ();
 sg13g2_decap_8 FILLER_57_1632 ();
 sg13g2_fill_2 FILLER_57_1639 ();
 sg13g2_fill_1 FILLER_57_1641 ();
 sg13g2_decap_4 FILLER_57_1668 ();
 sg13g2_fill_1 FILLER_57_1672 ();
 sg13g2_fill_2 FILLER_57_1686 ();
 sg13g2_decap_8 FILLER_57_1696 ();
 sg13g2_fill_2 FILLER_57_1703 ();
 sg13g2_decap_4 FILLER_57_1717 ();
 sg13g2_fill_2 FILLER_57_1721 ();
 sg13g2_fill_2 FILLER_57_1732 ();
 sg13g2_fill_1 FILLER_57_1734 ();
 sg13g2_decap_8 FILLER_57_1740 ();
 sg13g2_decap_8 FILLER_57_1747 ();
 sg13g2_decap_8 FILLER_57_1754 ();
 sg13g2_decap_8 FILLER_57_1761 ();
 sg13g2_decap_4 FILLER_57_1768 ();
 sg13g2_fill_2 FILLER_57_1772 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_fill_2 FILLER_58_35 ();
 sg13g2_fill_1 FILLER_58_37 ();
 sg13g2_fill_2 FILLER_58_42 ();
 sg13g2_fill_1 FILLER_58_44 ();
 sg13g2_decap_4 FILLER_58_58 ();
 sg13g2_fill_1 FILLER_58_62 ();
 sg13g2_decap_4 FILLER_58_68 ();
 sg13g2_fill_2 FILLER_58_81 ();
 sg13g2_fill_1 FILLER_58_83 ();
 sg13g2_decap_8 FILLER_58_102 ();
 sg13g2_decap_8 FILLER_58_109 ();
 sg13g2_decap_8 FILLER_58_116 ();
 sg13g2_fill_1 FILLER_58_123 ();
 sg13g2_decap_4 FILLER_58_134 ();
 sg13g2_fill_1 FILLER_58_143 ();
 sg13g2_decap_8 FILLER_58_148 ();
 sg13g2_fill_2 FILLER_58_155 ();
 sg13g2_fill_1 FILLER_58_157 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_fill_2 FILLER_58_182 ();
 sg13g2_fill_1 FILLER_58_194 ();
 sg13g2_decap_4 FILLER_58_200 ();
 sg13g2_fill_1 FILLER_58_220 ();
 sg13g2_decap_8 FILLER_58_229 ();
 sg13g2_fill_2 FILLER_58_236 ();
 sg13g2_fill_1 FILLER_58_238 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_decap_8 FILLER_58_252 ();
 sg13g2_fill_2 FILLER_58_259 ();
 sg13g2_fill_1 FILLER_58_261 ();
 sg13g2_decap_4 FILLER_58_280 ();
 sg13g2_fill_2 FILLER_58_284 ();
 sg13g2_decap_4 FILLER_58_290 ();
 sg13g2_decap_8 FILLER_58_299 ();
 sg13g2_decap_8 FILLER_58_319 ();
 sg13g2_decap_8 FILLER_58_326 ();
 sg13g2_fill_1 FILLER_58_333 ();
 sg13g2_decap_8 FILLER_58_339 ();
 sg13g2_decap_4 FILLER_58_346 ();
 sg13g2_decap_8 FILLER_58_355 ();
 sg13g2_decap_4 FILLER_58_367 ();
 sg13g2_decap_8 FILLER_58_375 ();
 sg13g2_fill_2 FILLER_58_382 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_58_406 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_fill_2 FILLER_58_417 ();
 sg13g2_decap_4 FILLER_58_424 ();
 sg13g2_fill_2 FILLER_58_428 ();
 sg13g2_decap_8 FILLER_58_440 ();
 sg13g2_decap_4 FILLER_58_447 ();
 sg13g2_fill_1 FILLER_58_451 ();
 sg13g2_decap_8 FILLER_58_458 ();
 sg13g2_decap_8 FILLER_58_465 ();
 sg13g2_decap_8 FILLER_58_472 ();
 sg13g2_decap_8 FILLER_58_479 ();
 sg13g2_fill_2 FILLER_58_486 ();
 sg13g2_decap_8 FILLER_58_521 ();
 sg13g2_decap_8 FILLER_58_528 ();
 sg13g2_decap_8 FILLER_58_535 ();
 sg13g2_decap_4 FILLER_58_542 ();
 sg13g2_decap_4 FILLER_58_550 ();
 sg13g2_fill_2 FILLER_58_554 ();
 sg13g2_decap_8 FILLER_58_560 ();
 sg13g2_decap_8 FILLER_58_567 ();
 sg13g2_decap_8 FILLER_58_574 ();
 sg13g2_decap_8 FILLER_58_581 ();
 sg13g2_decap_8 FILLER_58_588 ();
 sg13g2_fill_2 FILLER_58_595 ();
 sg13g2_decap_8 FILLER_58_638 ();
 sg13g2_fill_2 FILLER_58_645 ();
 sg13g2_fill_1 FILLER_58_647 ();
 sg13g2_decap_8 FILLER_58_683 ();
 sg13g2_decap_4 FILLER_58_690 ();
 sg13g2_fill_2 FILLER_58_694 ();
 sg13g2_fill_1 FILLER_58_712 ();
 sg13g2_fill_2 FILLER_58_721 ();
 sg13g2_fill_2 FILLER_58_729 ();
 sg13g2_fill_1 FILLER_58_731 ();
 sg13g2_decap_8 FILLER_58_737 ();
 sg13g2_decap_8 FILLER_58_744 ();
 sg13g2_decap_8 FILLER_58_751 ();
 sg13g2_decap_8 FILLER_58_758 ();
 sg13g2_decap_8 FILLER_58_765 ();
 sg13g2_decap_8 FILLER_58_772 ();
 sg13g2_decap_8 FILLER_58_779 ();
 sg13g2_decap_8 FILLER_58_786 ();
 sg13g2_decap_4 FILLER_58_793 ();
 sg13g2_fill_1 FILLER_58_797 ();
 sg13g2_decap_8 FILLER_58_802 ();
 sg13g2_decap_8 FILLER_58_809 ();
 sg13g2_decap_8 FILLER_58_816 ();
 sg13g2_decap_8 FILLER_58_823 ();
 sg13g2_decap_8 FILLER_58_833 ();
 sg13g2_fill_1 FILLER_58_840 ();
 sg13g2_decap_8 FILLER_58_845 ();
 sg13g2_decap_8 FILLER_58_852 ();
 sg13g2_decap_8 FILLER_58_859 ();
 sg13g2_decap_8 FILLER_58_866 ();
 sg13g2_fill_2 FILLER_58_873 ();
 sg13g2_decap_8 FILLER_58_879 ();
 sg13g2_decap_8 FILLER_58_886 ();
 sg13g2_decap_8 FILLER_58_893 ();
 sg13g2_decap_8 FILLER_58_900 ();
 sg13g2_decap_8 FILLER_58_907 ();
 sg13g2_decap_8 FILLER_58_914 ();
 sg13g2_decap_8 FILLER_58_921 ();
 sg13g2_decap_8 FILLER_58_928 ();
 sg13g2_decap_8 FILLER_58_935 ();
 sg13g2_decap_8 FILLER_58_942 ();
 sg13g2_decap_8 FILLER_58_949 ();
 sg13g2_decap_4 FILLER_58_956 ();
 sg13g2_decap_4 FILLER_58_964 ();
 sg13g2_fill_1 FILLER_58_979 ();
 sg13g2_fill_2 FILLER_58_1006 ();
 sg13g2_fill_2 FILLER_58_1012 ();
 sg13g2_fill_1 FILLER_58_1014 ();
 sg13g2_decap_8 FILLER_58_1033 ();
 sg13g2_decap_8 FILLER_58_1040 ();
 sg13g2_decap_8 FILLER_58_1047 ();
 sg13g2_decap_8 FILLER_58_1054 ();
 sg13g2_decap_8 FILLER_58_1061 ();
 sg13g2_decap_8 FILLER_58_1068 ();
 sg13g2_decap_8 FILLER_58_1075 ();
 sg13g2_decap_8 FILLER_58_1082 ();
 sg13g2_fill_1 FILLER_58_1097 ();
 sg13g2_fill_2 FILLER_58_1129 ();
 sg13g2_decap_8 FILLER_58_1148 ();
 sg13g2_decap_8 FILLER_58_1155 ();
 sg13g2_fill_2 FILLER_58_1162 ();
 sg13g2_fill_1 FILLER_58_1164 ();
 sg13g2_fill_2 FILLER_58_1168 ();
 sg13g2_fill_1 FILLER_58_1170 ();
 sg13g2_fill_1 FILLER_58_1184 ();
 sg13g2_decap_4 FILLER_58_1199 ();
 sg13g2_fill_2 FILLER_58_1203 ();
 sg13g2_fill_2 FILLER_58_1209 ();
 sg13g2_decap_8 FILLER_58_1223 ();
 sg13g2_fill_2 FILLER_58_1230 ();
 sg13g2_decap_8 FILLER_58_1245 ();
 sg13g2_decap_8 FILLER_58_1260 ();
 sg13g2_fill_1 FILLER_58_1267 ();
 sg13g2_fill_1 FILLER_58_1272 ();
 sg13g2_fill_2 FILLER_58_1281 ();
 sg13g2_fill_1 FILLER_58_1293 ();
 sg13g2_fill_2 FILLER_58_1301 ();
 sg13g2_fill_1 FILLER_58_1307 ();
 sg13g2_fill_1 FILLER_58_1313 ();
 sg13g2_decap_8 FILLER_58_1323 ();
 sg13g2_fill_2 FILLER_58_1330 ();
 sg13g2_fill_2 FILLER_58_1348 ();
 sg13g2_decap_8 FILLER_58_1354 ();
 sg13g2_fill_1 FILLER_58_1370 ();
 sg13g2_decap_8 FILLER_58_1375 ();
 sg13g2_decap_8 FILLER_58_1417 ();
 sg13g2_decap_8 FILLER_58_1424 ();
 sg13g2_decap_8 FILLER_58_1431 ();
 sg13g2_decap_4 FILLER_58_1438 ();
 sg13g2_fill_1 FILLER_58_1442 ();
 sg13g2_decap_8 FILLER_58_1450 ();
 sg13g2_decap_8 FILLER_58_1457 ();
 sg13g2_decap_4 FILLER_58_1464 ();
 sg13g2_fill_2 FILLER_58_1468 ();
 sg13g2_decap_8 FILLER_58_1480 ();
 sg13g2_fill_1 FILLER_58_1504 ();
 sg13g2_decap_4 FILLER_58_1510 ();
 sg13g2_decap_4 FILLER_58_1534 ();
 sg13g2_fill_2 FILLER_58_1541 ();
 sg13g2_decap_4 FILLER_58_1563 ();
 sg13g2_decap_4 FILLER_58_1576 ();
 sg13g2_decap_8 FILLER_58_1585 ();
 sg13g2_decap_8 FILLER_58_1592 ();
 sg13g2_decap_4 FILLER_58_1599 ();
 sg13g2_fill_2 FILLER_58_1606 ();
 sg13g2_fill_1 FILLER_58_1608 ();
 sg13g2_decap_8 FILLER_58_1618 ();
 sg13g2_fill_1 FILLER_58_1625 ();
 sg13g2_decap_8 FILLER_58_1631 ();
 sg13g2_decap_8 FILLER_58_1638 ();
 sg13g2_decap_4 FILLER_58_1645 ();
 sg13g2_fill_1 FILLER_58_1653 ();
 sg13g2_decap_8 FILLER_58_1660 ();
 sg13g2_decap_4 FILLER_58_1667 ();
 sg13g2_fill_2 FILLER_58_1671 ();
 sg13g2_decap_8 FILLER_58_1679 ();
 sg13g2_decap_4 FILLER_58_1686 ();
 sg13g2_decap_8 FILLER_58_1693 ();
 sg13g2_decap_8 FILLER_58_1700 ();
 sg13g2_fill_2 FILLER_58_1707 ();
 sg13g2_fill_1 FILLER_58_1717 ();
 sg13g2_decap_4 FILLER_58_1733 ();
 sg13g2_decap_8 FILLER_58_1741 ();
 sg13g2_decap_4 FILLER_58_1748 ();
 sg13g2_decap_8 FILLER_58_1756 ();
 sg13g2_decap_8 FILLER_58_1763 ();
 sg13g2_decap_4 FILLER_58_1770 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_4 FILLER_59_21 ();
 sg13g2_fill_2 FILLER_59_35 ();
 sg13g2_fill_1 FILLER_59_37 ();
 sg13g2_fill_2 FILLER_59_50 ();
 sg13g2_decap_8 FILLER_59_57 ();
 sg13g2_decap_4 FILLER_59_64 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_decap_4 FILLER_59_92 ();
 sg13g2_decap_8 FILLER_59_104 ();
 sg13g2_fill_2 FILLER_59_116 ();
 sg13g2_decap_8 FILLER_59_127 ();
 sg13g2_fill_1 FILLER_59_134 ();
 sg13g2_decap_8 FILLER_59_145 ();
 sg13g2_decap_4 FILLER_59_152 ();
 sg13g2_fill_2 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_163 ();
 sg13g2_decap_8 FILLER_59_173 ();
 sg13g2_decap_4 FILLER_59_186 ();
 sg13g2_decap_8 FILLER_59_195 ();
 sg13g2_decap_8 FILLER_59_202 ();
 sg13g2_decap_4 FILLER_59_209 ();
 sg13g2_fill_1 FILLER_59_232 ();
 sg13g2_decap_4 FILLER_59_238 ();
 sg13g2_fill_1 FILLER_59_242 ();
 sg13g2_decap_8 FILLER_59_248 ();
 sg13g2_decap_4 FILLER_59_255 ();
 sg13g2_fill_1 FILLER_59_259 ();
 sg13g2_fill_2 FILLER_59_264 ();
 sg13g2_fill_1 FILLER_59_266 ();
 sg13g2_decap_4 FILLER_59_275 ();
 sg13g2_decap_8 FILLER_59_283 ();
 sg13g2_fill_2 FILLER_59_290 ();
 sg13g2_decap_4 FILLER_59_301 ();
 sg13g2_fill_1 FILLER_59_305 ();
 sg13g2_fill_1 FILLER_59_311 ();
 sg13g2_decap_8 FILLER_59_317 ();
 sg13g2_decap_4 FILLER_59_324 ();
 sg13g2_decap_8 FILLER_59_333 ();
 sg13g2_fill_2 FILLER_59_340 ();
 sg13g2_decap_4 FILLER_59_360 ();
 sg13g2_decap_8 FILLER_59_389 ();
 sg13g2_decap_8 FILLER_59_396 ();
 sg13g2_decap_4 FILLER_59_403 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_4 FILLER_59_414 ();
 sg13g2_fill_1 FILLER_59_418 ();
 sg13g2_fill_1 FILLER_59_423 ();
 sg13g2_decap_8 FILLER_59_434 ();
 sg13g2_fill_2 FILLER_59_441 ();
 sg13g2_decap_4 FILLER_59_453 ();
 sg13g2_decap_8 FILLER_59_462 ();
 sg13g2_decap_8 FILLER_59_469 ();
 sg13g2_decap_8 FILLER_59_476 ();
 sg13g2_decap_8 FILLER_59_483 ();
 sg13g2_decap_8 FILLER_59_490 ();
 sg13g2_decap_8 FILLER_59_497 ();
 sg13g2_fill_1 FILLER_59_504 ();
 sg13g2_decap_8 FILLER_59_510 ();
 sg13g2_decap_8 FILLER_59_517 ();
 sg13g2_decap_8 FILLER_59_524 ();
 sg13g2_decap_8 FILLER_59_531 ();
 sg13g2_decap_8 FILLER_59_538 ();
 sg13g2_fill_1 FILLER_59_550 ();
 sg13g2_decap_8 FILLER_59_612 ();
 sg13g2_decap_8 FILLER_59_649 ();
 sg13g2_decap_8 FILLER_59_656 ();
 sg13g2_decap_8 FILLER_59_663 ();
 sg13g2_decap_8 FILLER_59_670 ();
 sg13g2_decap_8 FILLER_59_677 ();
 sg13g2_fill_1 FILLER_59_684 ();
 sg13g2_decap_8 FILLER_59_719 ();
 sg13g2_fill_2 FILLER_59_726 ();
 sg13g2_fill_1 FILLER_59_728 ();
 sg13g2_decap_8 FILLER_59_738 ();
 sg13g2_fill_2 FILLER_59_745 ();
 sg13g2_fill_1 FILLER_59_747 ();
 sg13g2_fill_2 FILLER_59_753 ();
 sg13g2_fill_1 FILLER_59_755 ();
 sg13g2_decap_8 FILLER_59_786 ();
 sg13g2_decap_8 FILLER_59_793 ();
 sg13g2_fill_2 FILLER_59_805 ();
 sg13g2_fill_1 FILLER_59_807 ();
 sg13g2_decap_8 FILLER_59_834 ();
 sg13g2_decap_4 FILLER_59_841 ();
 sg13g2_decap_8 FILLER_59_849 ();
 sg13g2_decap_8 FILLER_59_856 ();
 sg13g2_decap_8 FILLER_59_863 ();
 sg13g2_decap_8 FILLER_59_870 ();
 sg13g2_fill_2 FILLER_59_877 ();
 sg13g2_fill_1 FILLER_59_879 ();
 sg13g2_decap_8 FILLER_59_883 ();
 sg13g2_decap_4 FILLER_59_890 ();
 sg13g2_fill_2 FILLER_59_894 ();
 sg13g2_decap_8 FILLER_59_901 ();
 sg13g2_decap_4 FILLER_59_908 ();
 sg13g2_fill_2 FILLER_59_912 ();
 sg13g2_decap_8 FILLER_59_926 ();
 sg13g2_decap_4 FILLER_59_933 ();
 sg13g2_decap_8 FILLER_59_963 ();
 sg13g2_fill_2 FILLER_59_970 ();
 sg13g2_fill_1 FILLER_59_972 ();
 sg13g2_decap_4 FILLER_59_976 ();
 sg13g2_fill_2 FILLER_59_980 ();
 sg13g2_fill_1 FILLER_59_986 ();
 sg13g2_decap_8 FILLER_59_991 ();
 sg13g2_decap_4 FILLER_59_998 ();
 sg13g2_fill_2 FILLER_59_1002 ();
 sg13g2_decap_8 FILLER_59_1035 ();
 sg13g2_decap_8 FILLER_59_1042 ();
 sg13g2_decap_4 FILLER_59_1049 ();
 sg13g2_decap_8 FILLER_59_1062 ();
 sg13g2_decap_8 FILLER_59_1069 ();
 sg13g2_decap_8 FILLER_59_1076 ();
 sg13g2_fill_2 FILLER_59_1083 ();
 sg13g2_fill_1 FILLER_59_1085 ();
 sg13g2_decap_8 FILLER_59_1096 ();
 sg13g2_decap_8 FILLER_59_1103 ();
 sg13g2_decap_8 FILLER_59_1110 ();
 sg13g2_fill_1 FILLER_59_1117 ();
 sg13g2_fill_2 FILLER_59_1127 ();
 sg13g2_decap_8 FILLER_59_1150 ();
 sg13g2_fill_2 FILLER_59_1157 ();
 sg13g2_fill_1 FILLER_59_1159 ();
 sg13g2_decap_8 FILLER_59_1186 ();
 sg13g2_fill_2 FILLER_59_1193 ();
 sg13g2_fill_1 FILLER_59_1195 ();
 sg13g2_decap_8 FILLER_59_1200 ();
 sg13g2_decap_8 FILLER_59_1207 ();
 sg13g2_decap_8 FILLER_59_1214 ();
 sg13g2_decap_8 FILLER_59_1221 ();
 sg13g2_fill_2 FILLER_59_1228 ();
 sg13g2_decap_8 FILLER_59_1250 ();
 sg13g2_decap_8 FILLER_59_1257 ();
 sg13g2_decap_8 FILLER_59_1264 ();
 sg13g2_decap_8 FILLER_59_1271 ();
 sg13g2_decap_8 FILLER_59_1278 ();
 sg13g2_decap_8 FILLER_59_1285 ();
 sg13g2_decap_4 FILLER_59_1292 ();
 sg13g2_fill_1 FILLER_59_1296 ();
 sg13g2_decap_8 FILLER_59_1302 ();
 sg13g2_decap_8 FILLER_59_1309 ();
 sg13g2_decap_8 FILLER_59_1316 ();
 sg13g2_decap_4 FILLER_59_1323 ();
 sg13g2_fill_2 FILLER_59_1327 ();
 sg13g2_fill_1 FILLER_59_1337 ();
 sg13g2_fill_2 FILLER_59_1342 ();
 sg13g2_decap_8 FILLER_59_1349 ();
 sg13g2_decap_8 FILLER_59_1356 ();
 sg13g2_decap_8 FILLER_59_1363 ();
 sg13g2_decap_8 FILLER_59_1370 ();
 sg13g2_decap_8 FILLER_59_1377 ();
 sg13g2_decap_8 FILLER_59_1384 ();
 sg13g2_decap_4 FILLER_59_1391 ();
 sg13g2_fill_1 FILLER_59_1395 ();
 sg13g2_decap_8 FILLER_59_1406 ();
 sg13g2_decap_8 FILLER_59_1413 ();
 sg13g2_decap_8 FILLER_59_1420 ();
 sg13g2_decap_4 FILLER_59_1427 ();
 sg13g2_fill_1 FILLER_59_1431 ();
 sg13g2_decap_4 FILLER_59_1444 ();
 sg13g2_fill_1 FILLER_59_1448 ();
 sg13g2_decap_8 FILLER_59_1453 ();
 sg13g2_decap_8 FILLER_59_1460 ();
 sg13g2_decap_8 FILLER_59_1467 ();
 sg13g2_fill_2 FILLER_59_1474 ();
 sg13g2_fill_1 FILLER_59_1476 ();
 sg13g2_fill_2 FILLER_59_1482 ();
 sg13g2_fill_2 FILLER_59_1487 ();
 sg13g2_fill_1 FILLER_59_1489 ();
 sg13g2_fill_2 FILLER_59_1499 ();
 sg13g2_fill_1 FILLER_59_1501 ();
 sg13g2_fill_2 FILLER_59_1524 ();
 sg13g2_fill_1 FILLER_59_1532 ();
 sg13g2_fill_2 FILLER_59_1541 ();
 sg13g2_decap_4 FILLER_59_1555 ();
 sg13g2_decap_8 FILLER_59_1578 ();
 sg13g2_decap_8 FILLER_59_1585 ();
 sg13g2_decap_8 FILLER_59_1592 ();
 sg13g2_fill_2 FILLER_59_1599 ();
 sg13g2_fill_1 FILLER_59_1601 ();
 sg13g2_decap_8 FILLER_59_1632 ();
 sg13g2_decap_8 FILLER_59_1639 ();
 sg13g2_decap_8 FILLER_59_1646 ();
 sg13g2_decap_8 FILLER_59_1653 ();
 sg13g2_decap_4 FILLER_59_1660 ();
 sg13g2_fill_1 FILLER_59_1664 ();
 sg13g2_decap_4 FILLER_59_1669 ();
 sg13g2_fill_2 FILLER_59_1673 ();
 sg13g2_fill_2 FILLER_59_1678 ();
 sg13g2_fill_1 FILLER_59_1680 ();
 sg13g2_decap_8 FILLER_59_1686 ();
 sg13g2_decap_8 FILLER_59_1693 ();
 sg13g2_decap_8 FILLER_59_1700 ();
 sg13g2_decap_8 FILLER_59_1707 ();
 sg13g2_fill_2 FILLER_59_1718 ();
 sg13g2_decap_4 FILLER_59_1725 ();
 sg13g2_fill_2 FILLER_59_1729 ();
 sg13g2_decap_4 FILLER_59_1770 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_fill_2 FILLER_60_21 ();
 sg13g2_fill_1 FILLER_60_23 ();
 sg13g2_fill_2 FILLER_60_36 ();
 sg13g2_fill_1 FILLER_60_38 ();
 sg13g2_decap_4 FILLER_60_57 ();
 sg13g2_fill_2 FILLER_60_61 ();
 sg13g2_decap_8 FILLER_60_68 ();
 sg13g2_decap_4 FILLER_60_75 ();
 sg13g2_fill_1 FILLER_60_89 ();
 sg13g2_fill_2 FILLER_60_99 ();
 sg13g2_fill_1 FILLER_60_101 ();
 sg13g2_fill_1 FILLER_60_107 ();
 sg13g2_fill_2 FILLER_60_113 ();
 sg13g2_decap_4 FILLER_60_134 ();
 sg13g2_fill_2 FILLER_60_138 ();
 sg13g2_fill_2 FILLER_60_148 ();
 sg13g2_fill_1 FILLER_60_150 ();
 sg13g2_decap_8 FILLER_60_157 ();
 sg13g2_fill_2 FILLER_60_164 ();
 sg13g2_fill_1 FILLER_60_166 ();
 sg13g2_fill_2 FILLER_60_177 ();
 sg13g2_fill_1 FILLER_60_179 ();
 sg13g2_fill_2 FILLER_60_186 ();
 sg13g2_fill_2 FILLER_60_194 ();
 sg13g2_decap_8 FILLER_60_201 ();
 sg13g2_decap_4 FILLER_60_208 ();
 sg13g2_fill_1 FILLER_60_212 ();
 sg13g2_fill_1 FILLER_60_220 ();
 sg13g2_decap_8 FILLER_60_226 ();
 sg13g2_decap_8 FILLER_60_233 ();
 sg13g2_decap_8 FILLER_60_240 ();
 sg13g2_decap_8 FILLER_60_247 ();
 sg13g2_fill_1 FILLER_60_254 ();
 sg13g2_decap_4 FILLER_60_259 ();
 sg13g2_decap_8 FILLER_60_268 ();
 sg13g2_decap_8 FILLER_60_275 ();
 sg13g2_decap_8 FILLER_60_282 ();
 sg13g2_decap_8 FILLER_60_289 ();
 sg13g2_decap_4 FILLER_60_311 ();
 sg13g2_decap_8 FILLER_60_333 ();
 sg13g2_decap_4 FILLER_60_340 ();
 sg13g2_decap_4 FILLER_60_354 ();
 sg13g2_fill_1 FILLER_60_358 ();
 sg13g2_decap_8 FILLER_60_364 ();
 sg13g2_decap_8 FILLER_60_371 ();
 sg13g2_decap_8 FILLER_60_392 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_fill_2 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_408 ();
 sg13g2_decap_8 FILLER_60_414 ();
 sg13g2_fill_2 FILLER_60_421 ();
 sg13g2_decap_4 FILLER_60_427 ();
 sg13g2_fill_1 FILLER_60_431 ();
 sg13g2_decap_8 FILLER_60_442 ();
 sg13g2_fill_2 FILLER_60_449 ();
 sg13g2_decap_8 FILLER_60_461 ();
 sg13g2_decap_8 FILLER_60_468 ();
 sg13g2_decap_8 FILLER_60_475 ();
 sg13g2_decap_8 FILLER_60_482 ();
 sg13g2_decap_8 FILLER_60_489 ();
 sg13g2_fill_2 FILLER_60_496 ();
 sg13g2_decap_4 FILLER_60_507 ();
 sg13g2_fill_1 FILLER_60_511 ();
 sg13g2_decap_4 FILLER_60_542 ();
 sg13g2_decap_8 FILLER_60_551 ();
 sg13g2_decap_8 FILLER_60_562 ();
 sg13g2_decap_8 FILLER_60_569 ();
 sg13g2_decap_8 FILLER_60_576 ();
 sg13g2_decap_8 FILLER_60_583 ();
 sg13g2_decap_4 FILLER_60_590 ();
 sg13g2_fill_1 FILLER_60_594 ();
 sg13g2_decap_8 FILLER_60_599 ();
 sg13g2_decap_8 FILLER_60_606 ();
 sg13g2_decap_8 FILLER_60_613 ();
 sg13g2_decap_8 FILLER_60_620 ();
 sg13g2_fill_1 FILLER_60_627 ();
 sg13g2_decap_8 FILLER_60_680 ();
 sg13g2_decap_4 FILLER_60_687 ();
 sg13g2_fill_1 FILLER_60_691 ();
 sg13g2_decap_8 FILLER_60_696 ();
 sg13g2_decap_8 FILLER_60_703 ();
 sg13g2_decap_8 FILLER_60_710 ();
 sg13g2_decap_8 FILLER_60_717 ();
 sg13g2_decap_8 FILLER_60_724 ();
 sg13g2_fill_1 FILLER_60_731 ();
 sg13g2_decap_8 FILLER_60_736 ();
 sg13g2_fill_2 FILLER_60_743 ();
 sg13g2_fill_1 FILLER_60_745 ();
 sg13g2_decap_8 FILLER_60_754 ();
 sg13g2_fill_1 FILLER_60_761 ();
 sg13g2_decap_8 FILLER_60_766 ();
 sg13g2_decap_8 FILLER_60_773 ();
 sg13g2_decap_8 FILLER_60_780 ();
 sg13g2_decap_8 FILLER_60_787 ();
 sg13g2_decap_4 FILLER_60_794 ();
 sg13g2_fill_2 FILLER_60_798 ();
 sg13g2_fill_2 FILLER_60_808 ();
 sg13g2_fill_1 FILLER_60_810 ();
 sg13g2_decap_4 FILLER_60_815 ();
 sg13g2_decap_8 FILLER_60_823 ();
 sg13g2_decap_8 FILLER_60_830 ();
 sg13g2_fill_2 FILLER_60_837 ();
 sg13g2_decap_4 FILLER_60_890 ();
 sg13g2_fill_2 FILLER_60_894 ();
 sg13g2_decap_8 FILLER_60_903 ();
 sg13g2_fill_2 FILLER_60_910 ();
 sg13g2_fill_1 FILLER_60_920 ();
 sg13g2_fill_1 FILLER_60_926 ();
 sg13g2_fill_2 FILLER_60_938 ();
 sg13g2_fill_1 FILLER_60_940 ();
 sg13g2_decap_4 FILLER_60_945 ();
 sg13g2_fill_2 FILLER_60_949 ();
 sg13g2_decap_8 FILLER_60_955 ();
 sg13g2_decap_8 FILLER_60_962 ();
 sg13g2_decap_4 FILLER_60_969 ();
 sg13g2_decap_8 FILLER_60_978 ();
 sg13g2_decap_4 FILLER_60_985 ();
 sg13g2_fill_1 FILLER_60_989 ();
 sg13g2_fill_1 FILLER_60_995 ();
 sg13g2_decap_8 FILLER_60_1010 ();
 sg13g2_fill_2 FILLER_60_1017 ();
 sg13g2_fill_1 FILLER_60_1019 ();
 sg13g2_fill_2 FILLER_60_1024 ();
 sg13g2_fill_1 FILLER_60_1026 ();
 sg13g2_decap_8 FILLER_60_1031 ();
 sg13g2_decap_8 FILLER_60_1038 ();
 sg13g2_decap_8 FILLER_60_1045 ();
 sg13g2_decap_8 FILLER_60_1052 ();
 sg13g2_decap_8 FILLER_60_1059 ();
 sg13g2_decap_8 FILLER_60_1066 ();
 sg13g2_decap_8 FILLER_60_1073 ();
 sg13g2_fill_2 FILLER_60_1080 ();
 sg13g2_fill_1 FILLER_60_1112 ();
 sg13g2_fill_1 FILLER_60_1124 ();
 sg13g2_decap_8 FILLER_60_1138 ();
 sg13g2_fill_2 FILLER_60_1145 ();
 sg13g2_decap_8 FILLER_60_1152 ();
 sg13g2_decap_8 FILLER_60_1159 ();
 sg13g2_decap_8 FILLER_60_1166 ();
 sg13g2_fill_1 FILLER_60_1177 ();
 sg13g2_decap_4 FILLER_60_1187 ();
 sg13g2_fill_2 FILLER_60_1191 ();
 sg13g2_fill_2 FILLER_60_1197 ();
 sg13g2_decap_8 FILLER_60_1208 ();
 sg13g2_decap_8 FILLER_60_1215 ();
 sg13g2_decap_4 FILLER_60_1222 ();
 sg13g2_fill_1 FILLER_60_1226 ();
 sg13g2_decap_8 FILLER_60_1247 ();
 sg13g2_decap_8 FILLER_60_1254 ();
 sg13g2_fill_1 FILLER_60_1265 ();
 sg13g2_decap_8 FILLER_60_1292 ();
 sg13g2_decap_4 FILLER_60_1308 ();
 sg13g2_fill_1 FILLER_60_1312 ();
 sg13g2_decap_4 FILLER_60_1318 ();
 sg13g2_fill_1 FILLER_60_1322 ();
 sg13g2_decap_8 FILLER_60_1328 ();
 sg13g2_decap_8 FILLER_60_1340 ();
 sg13g2_decap_8 FILLER_60_1347 ();
 sg13g2_decap_8 FILLER_60_1354 ();
 sg13g2_decap_8 FILLER_60_1361 ();
 sg13g2_decap_8 FILLER_60_1368 ();
 sg13g2_fill_2 FILLER_60_1404 ();
 sg13g2_decap_4 FILLER_60_1422 ();
 sg13g2_fill_1 FILLER_60_1426 ();
 sg13g2_fill_1 FILLER_60_1447 ();
 sg13g2_decap_8 FILLER_60_1452 ();
 sg13g2_decap_8 FILLER_60_1459 ();
 sg13g2_decap_4 FILLER_60_1466 ();
 sg13g2_fill_1 FILLER_60_1470 ();
 sg13g2_decap_8 FILLER_60_1475 ();
 sg13g2_fill_1 FILLER_60_1482 ();
 sg13g2_fill_1 FILLER_60_1513 ();
 sg13g2_fill_1 FILLER_60_1531 ();
 sg13g2_fill_2 FILLER_60_1549 ();
 sg13g2_fill_2 FILLER_60_1573 ();
 sg13g2_decap_8 FILLER_60_1579 ();
 sg13g2_fill_1 FILLER_60_1586 ();
 sg13g2_decap_8 FILLER_60_1592 ();
 sg13g2_decap_8 FILLER_60_1599 ();
 sg13g2_decap_8 FILLER_60_1606 ();
 sg13g2_decap_8 FILLER_60_1613 ();
 sg13g2_decap_8 FILLER_60_1620 ();
 sg13g2_fill_2 FILLER_60_1627 ();
 sg13g2_fill_2 FILLER_60_1634 ();
 sg13g2_fill_2 FILLER_60_1644 ();
 sg13g2_fill_1 FILLER_60_1652 ();
 sg13g2_decap_8 FILLER_60_1686 ();
 sg13g2_decap_8 FILLER_60_1693 ();
 sg13g2_decap_8 FILLER_60_1700 ();
 sg13g2_decap_8 FILLER_60_1707 ();
 sg13g2_decap_8 FILLER_60_1714 ();
 sg13g2_decap_8 FILLER_60_1721 ();
 sg13g2_fill_2 FILLER_60_1728 ();
 sg13g2_fill_2 FILLER_60_1733 ();
 sg13g2_decap_8 FILLER_60_1761 ();
 sg13g2_decap_4 FILLER_60_1768 ();
 sg13g2_fill_2 FILLER_60_1772 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_4 FILLER_61_54 ();
 sg13g2_fill_2 FILLER_61_62 ();
 sg13g2_fill_1 FILLER_61_64 ();
 sg13g2_fill_2 FILLER_61_83 ();
 sg13g2_fill_1 FILLER_61_85 ();
 sg13g2_decap_8 FILLER_61_95 ();
 sg13g2_decap_4 FILLER_61_102 ();
 sg13g2_fill_1 FILLER_61_122 ();
 sg13g2_decap_4 FILLER_61_127 ();
 sg13g2_decap_8 FILLER_61_136 ();
 sg13g2_fill_2 FILLER_61_150 ();
 sg13g2_fill_1 FILLER_61_152 ();
 sg13g2_decap_8 FILLER_61_158 ();
 sg13g2_fill_2 FILLER_61_165 ();
 sg13g2_decap_4 FILLER_61_182 ();
 sg13g2_decap_4 FILLER_61_191 ();
 sg13g2_fill_2 FILLER_61_195 ();
 sg13g2_decap_8 FILLER_61_202 ();
 sg13g2_decap_4 FILLER_61_209 ();
 sg13g2_fill_2 FILLER_61_213 ();
 sg13g2_fill_2 FILLER_61_219 ();
 sg13g2_fill_1 FILLER_61_221 ();
 sg13g2_fill_2 FILLER_61_227 ();
 sg13g2_decap_8 FILLER_61_241 ();
 sg13g2_decap_8 FILLER_61_248 ();
 sg13g2_fill_1 FILLER_61_255 ();
 sg13g2_decap_4 FILLER_61_271 ();
 sg13g2_fill_1 FILLER_61_275 ();
 sg13g2_decap_4 FILLER_61_281 ();
 sg13g2_decap_8 FILLER_61_295 ();
 sg13g2_decap_8 FILLER_61_302 ();
 sg13g2_fill_2 FILLER_61_309 ();
 sg13g2_decap_4 FILLER_61_316 ();
 sg13g2_fill_2 FILLER_61_320 ();
 sg13g2_decap_8 FILLER_61_326 ();
 sg13g2_fill_2 FILLER_61_333 ();
 sg13g2_fill_1 FILLER_61_335 ();
 sg13g2_fill_2 FILLER_61_341 ();
 sg13g2_fill_1 FILLER_61_343 ();
 sg13g2_decap_4 FILLER_61_349 ();
 sg13g2_decap_4 FILLER_61_358 ();
 sg13g2_fill_1 FILLER_61_362 ();
 sg13g2_decap_4 FILLER_61_368 ();
 sg13g2_fill_2 FILLER_61_372 ();
 sg13g2_decap_8 FILLER_61_383 ();
 sg13g2_decap_8 FILLER_61_390 ();
 sg13g2_fill_1 FILLER_61_397 ();
 sg13g2_fill_2 FILLER_61_402 ();
 sg13g2_fill_1 FILLER_61_404 ();
 sg13g2_fill_1 FILLER_61_409 ();
 sg13g2_fill_1 FILLER_61_415 ();
 sg13g2_fill_1 FILLER_61_424 ();
 sg13g2_fill_1 FILLER_61_430 ();
 sg13g2_decap_8 FILLER_61_441 ();
 sg13g2_decap_4 FILLER_61_448 ();
 sg13g2_fill_1 FILLER_61_452 ();
 sg13g2_decap_8 FILLER_61_457 ();
 sg13g2_decap_8 FILLER_61_464 ();
 sg13g2_decap_8 FILLER_61_471 ();
 sg13g2_decap_8 FILLER_61_478 ();
 sg13g2_decap_8 FILLER_61_485 ();
 sg13g2_decap_8 FILLER_61_492 ();
 sg13g2_decap_8 FILLER_61_499 ();
 sg13g2_decap_8 FILLER_61_506 ();
 sg13g2_decap_4 FILLER_61_513 ();
 sg13g2_fill_1 FILLER_61_517 ();
 sg13g2_decap_8 FILLER_61_526 ();
 sg13g2_decap_8 FILLER_61_533 ();
 sg13g2_fill_1 FILLER_61_540 ();
 sg13g2_decap_8 FILLER_61_566 ();
 sg13g2_decap_8 FILLER_61_573 ();
 sg13g2_decap_8 FILLER_61_580 ();
 sg13g2_fill_1 FILLER_61_587 ();
 sg13g2_decap_8 FILLER_61_592 ();
 sg13g2_decap_4 FILLER_61_599 ();
 sg13g2_fill_1 FILLER_61_603 ();
 sg13g2_decap_4 FILLER_61_614 ();
 sg13g2_decap_8 FILLER_61_644 ();
 sg13g2_fill_1 FILLER_61_651 ();
 sg13g2_decap_4 FILLER_61_655 ();
 sg13g2_fill_1 FILLER_61_659 ();
 sg13g2_decap_8 FILLER_61_664 ();
 sg13g2_decap_8 FILLER_61_671 ();
 sg13g2_decap_8 FILLER_61_678 ();
 sg13g2_decap_8 FILLER_61_685 ();
 sg13g2_decap_8 FILLER_61_692 ();
 sg13g2_decap_8 FILLER_61_699 ();
 sg13g2_decap_8 FILLER_61_706 ();
 sg13g2_decap_4 FILLER_61_713 ();
 sg13g2_fill_1 FILLER_61_717 ();
 sg13g2_decap_8 FILLER_61_722 ();
 sg13g2_fill_2 FILLER_61_729 ();
 sg13g2_decap_8 FILLER_61_735 ();
 sg13g2_fill_2 FILLER_61_742 ();
 sg13g2_decap_8 FILLER_61_751 ();
 sg13g2_decap_8 FILLER_61_758 ();
 sg13g2_fill_2 FILLER_61_765 ();
 sg13g2_fill_2 FILLER_61_777 ();
 sg13g2_fill_1 FILLER_61_790 ();
 sg13g2_decap_8 FILLER_61_805 ();
 sg13g2_decap_8 FILLER_61_812 ();
 sg13g2_decap_8 FILLER_61_819 ();
 sg13g2_decap_8 FILLER_61_826 ();
 sg13g2_decap_8 FILLER_61_833 ();
 sg13g2_fill_1 FILLER_61_840 ();
 sg13g2_decap_8 FILLER_61_846 ();
 sg13g2_decap_4 FILLER_61_853 ();
 sg13g2_fill_1 FILLER_61_857 ();
 sg13g2_decap_8 FILLER_61_862 ();
 sg13g2_decap_8 FILLER_61_869 ();
 sg13g2_decap_8 FILLER_61_876 ();
 sg13g2_decap_8 FILLER_61_883 ();
 sg13g2_fill_1 FILLER_61_890 ();
 sg13g2_decap_8 FILLER_61_894 ();
 sg13g2_decap_8 FILLER_61_901 ();
 sg13g2_decap_8 FILLER_61_908 ();
 sg13g2_decap_8 FILLER_61_915 ();
 sg13g2_decap_8 FILLER_61_922 ();
 sg13g2_decap_8 FILLER_61_929 ();
 sg13g2_decap_8 FILLER_61_936 ();
 sg13g2_fill_2 FILLER_61_943 ();
 sg13g2_fill_2 FILLER_61_950 ();
 sg13g2_decap_8 FILLER_61_955 ();
 sg13g2_decap_8 FILLER_61_962 ();
 sg13g2_decap_8 FILLER_61_969 ();
 sg13g2_decap_8 FILLER_61_976 ();
 sg13g2_decap_8 FILLER_61_983 ();
 sg13g2_fill_2 FILLER_61_990 ();
 sg13g2_fill_1 FILLER_61_992 ();
 sg13g2_decap_8 FILLER_61_1001 ();
 sg13g2_decap_8 FILLER_61_1008 ();
 sg13g2_decap_4 FILLER_61_1015 ();
 sg13g2_fill_2 FILLER_61_1019 ();
 sg13g2_fill_1 FILLER_61_1047 ();
 sg13g2_decap_8 FILLER_61_1053 ();
 sg13g2_decap_8 FILLER_61_1060 ();
 sg13g2_decap_8 FILLER_61_1067 ();
 sg13g2_decap_8 FILLER_61_1074 ();
 sg13g2_decap_8 FILLER_61_1081 ();
 sg13g2_decap_8 FILLER_61_1105 ();
 sg13g2_decap_8 FILLER_61_1115 ();
 sg13g2_decap_8 FILLER_61_1122 ();
 sg13g2_decap_8 FILLER_61_1129 ();
 sg13g2_decap_8 FILLER_61_1136 ();
 sg13g2_decap_4 FILLER_61_1143 ();
 sg13g2_fill_1 FILLER_61_1147 ();
 sg13g2_decap_8 FILLER_61_1156 ();
 sg13g2_decap_8 FILLER_61_1163 ();
 sg13g2_fill_2 FILLER_61_1170 ();
 sg13g2_decap_8 FILLER_61_1177 ();
 sg13g2_fill_2 FILLER_61_1184 ();
 sg13g2_decap_8 FILLER_61_1204 ();
 sg13g2_decap_8 FILLER_61_1211 ();
 sg13g2_decap_8 FILLER_61_1218 ();
 sg13g2_decap_4 FILLER_61_1225 ();
 sg13g2_fill_1 FILLER_61_1229 ();
 sg13g2_decap_8 FILLER_61_1248 ();
 sg13g2_decap_8 FILLER_61_1255 ();
 sg13g2_decap_8 FILLER_61_1262 ();
 sg13g2_fill_2 FILLER_61_1269 ();
 sg13g2_decap_8 FILLER_61_1309 ();
 sg13g2_decap_4 FILLER_61_1316 ();
 sg13g2_fill_1 FILLER_61_1320 ();
 sg13g2_decap_8 FILLER_61_1336 ();
 sg13g2_decap_8 FILLER_61_1343 ();
 sg13g2_decap_8 FILLER_61_1350 ();
 sg13g2_decap_8 FILLER_61_1357 ();
 sg13g2_decap_8 FILLER_61_1364 ();
 sg13g2_decap_8 FILLER_61_1371 ();
 sg13g2_decap_8 FILLER_61_1378 ();
 sg13g2_fill_2 FILLER_61_1385 ();
 sg13g2_fill_1 FILLER_61_1387 ();
 sg13g2_decap_4 FILLER_61_1392 ();
 sg13g2_decap_8 FILLER_61_1414 ();
 sg13g2_decap_8 FILLER_61_1421 ();
 sg13g2_decap_8 FILLER_61_1428 ();
 sg13g2_decap_8 FILLER_61_1435 ();
 sg13g2_decap_8 FILLER_61_1442 ();
 sg13g2_decap_4 FILLER_61_1449 ();
 sg13g2_fill_2 FILLER_61_1466 ();
 sg13g2_fill_1 FILLER_61_1473 ();
 sg13g2_decap_8 FILLER_61_1478 ();
 sg13g2_decap_4 FILLER_61_1485 ();
 sg13g2_fill_2 FILLER_61_1489 ();
 sg13g2_decap_8 FILLER_61_1495 ();
 sg13g2_fill_1 FILLER_61_1502 ();
 sg13g2_fill_2 FILLER_61_1507 ();
 sg13g2_fill_1 FILLER_61_1516 ();
 sg13g2_fill_1 FILLER_61_1534 ();
 sg13g2_fill_1 FILLER_61_1564 ();
 sg13g2_fill_1 FILLER_61_1574 ();
 sg13g2_decap_8 FILLER_61_1580 ();
 sg13g2_decap_8 FILLER_61_1587 ();
 sg13g2_decap_8 FILLER_61_1594 ();
 sg13g2_decap_8 FILLER_61_1601 ();
 sg13g2_decap_8 FILLER_61_1608 ();
 sg13g2_decap_8 FILLER_61_1615 ();
 sg13g2_decap_8 FILLER_61_1622 ();
 sg13g2_fill_1 FILLER_61_1629 ();
 sg13g2_decap_8 FILLER_61_1650 ();
 sg13g2_fill_2 FILLER_61_1657 ();
 sg13g2_decap_8 FILLER_61_1677 ();
 sg13g2_decap_8 FILLER_61_1684 ();
 sg13g2_fill_1 FILLER_61_1691 ();
 sg13g2_fill_1 FILLER_61_1718 ();
 sg13g2_decap_8 FILLER_61_1723 ();
 sg13g2_decap_8 FILLER_61_1730 ();
 sg13g2_decap_4 FILLER_61_1737 ();
 sg13g2_fill_1 FILLER_61_1741 ();
 sg13g2_decap_8 FILLER_61_1746 ();
 sg13g2_decap_8 FILLER_61_1753 ();
 sg13g2_decap_8 FILLER_61_1760 ();
 sg13g2_decap_8 FILLER_61_1767 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_21 ();
 sg13g2_fill_1 FILLER_62_25 ();
 sg13g2_fill_2 FILLER_62_35 ();
 sg13g2_fill_1 FILLER_62_37 ();
 sg13g2_fill_2 FILLER_62_46 ();
 sg13g2_fill_1 FILLER_62_48 ();
 sg13g2_fill_2 FILLER_62_58 ();
 sg13g2_decap_4 FILLER_62_68 ();
 sg13g2_fill_2 FILLER_62_72 ();
 sg13g2_fill_2 FILLER_62_79 ();
 sg13g2_decap_4 FILLER_62_87 ();
 sg13g2_fill_2 FILLER_62_91 ();
 sg13g2_decap_4 FILLER_62_97 ();
 sg13g2_fill_2 FILLER_62_101 ();
 sg13g2_decap_8 FILLER_62_107 ();
 sg13g2_fill_1 FILLER_62_114 ();
 sg13g2_fill_2 FILLER_62_125 ();
 sg13g2_fill_1 FILLER_62_127 ();
 sg13g2_decap_8 FILLER_62_132 ();
 sg13g2_fill_2 FILLER_62_139 ();
 sg13g2_fill_2 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_190 ();
 sg13g2_fill_1 FILLER_62_197 ();
 sg13g2_decap_8 FILLER_62_208 ();
 sg13g2_fill_2 FILLER_62_215 ();
 sg13g2_decap_8 FILLER_62_225 ();
 sg13g2_decap_8 FILLER_62_232 ();
 sg13g2_fill_2 FILLER_62_239 ();
 sg13g2_fill_1 FILLER_62_241 ();
 sg13g2_decap_8 FILLER_62_247 ();
 sg13g2_decap_8 FILLER_62_254 ();
 sg13g2_decap_8 FILLER_62_261 ();
 sg13g2_decap_8 FILLER_62_268 ();
 sg13g2_decap_4 FILLER_62_275 ();
 sg13g2_fill_2 FILLER_62_279 ();
 sg13g2_fill_2 FILLER_62_286 ();
 sg13g2_fill_1 FILLER_62_288 ();
 sg13g2_fill_1 FILLER_62_305 ();
 sg13g2_decap_4 FILLER_62_311 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_320 ();
 sg13g2_decap_4 FILLER_62_327 ();
 sg13g2_fill_1 FILLER_62_346 ();
 sg13g2_decap_8 FILLER_62_352 ();
 sg13g2_decap_4 FILLER_62_359 ();
 sg13g2_decap_8 FILLER_62_368 ();
 sg13g2_decap_4 FILLER_62_375 ();
 sg13g2_fill_1 FILLER_62_379 ();
 sg13g2_decap_8 FILLER_62_384 ();
 sg13g2_decap_4 FILLER_62_391 ();
 sg13g2_fill_2 FILLER_62_401 ();
 sg13g2_fill_1 FILLER_62_412 ();
 sg13g2_fill_1 FILLER_62_441 ();
 sg13g2_decap_8 FILLER_62_447 ();
 sg13g2_decap_8 FILLER_62_454 ();
 sg13g2_decap_8 FILLER_62_461 ();
 sg13g2_decap_8 FILLER_62_468 ();
 sg13g2_decap_8 FILLER_62_475 ();
 sg13g2_decap_8 FILLER_62_482 ();
 sg13g2_decap_8 FILLER_62_489 ();
 sg13g2_decap_4 FILLER_62_496 ();
 sg13g2_decap_8 FILLER_62_513 ();
 sg13g2_decap_8 FILLER_62_520 ();
 sg13g2_decap_8 FILLER_62_527 ();
 sg13g2_fill_2 FILLER_62_534 ();
 sg13g2_fill_1 FILLER_62_536 ();
 sg13g2_fill_2 FILLER_62_573 ();
 sg13g2_decap_8 FILLER_62_606 ();
 sg13g2_decap_8 FILLER_62_613 ();
 sg13g2_decap_4 FILLER_62_620 ();
 sg13g2_decap_8 FILLER_62_628 ();
 sg13g2_decap_8 FILLER_62_635 ();
 sg13g2_decap_8 FILLER_62_642 ();
 sg13g2_fill_1 FILLER_62_656 ();
 sg13g2_fill_2 FILLER_62_669 ();
 sg13g2_fill_1 FILLER_62_678 ();
 sg13g2_decap_8 FILLER_62_683 ();
 sg13g2_decap_8 FILLER_62_690 ();
 sg13g2_decap_8 FILLER_62_697 ();
 sg13g2_fill_2 FILLER_62_704 ();
 sg13g2_decap_8 FILLER_62_737 ();
 sg13g2_decap_8 FILLER_62_756 ();
 sg13g2_decap_8 FILLER_62_763 ();
 sg13g2_fill_2 FILLER_62_770 ();
 sg13g2_decap_4 FILLER_62_777 ();
 sg13g2_decap_8 FILLER_62_803 ();
 sg13g2_decap_8 FILLER_62_810 ();
 sg13g2_decap_8 FILLER_62_817 ();
 sg13g2_decap_8 FILLER_62_824 ();
 sg13g2_decap_4 FILLER_62_831 ();
 sg13g2_fill_1 FILLER_62_835 ();
 sg13g2_fill_1 FILLER_62_844 ();
 sg13g2_fill_2 FILLER_62_849 ();
 sg13g2_fill_2 FILLER_62_855 ();
 sg13g2_fill_1 FILLER_62_857 ();
 sg13g2_fill_1 FILLER_62_862 ();
 sg13g2_fill_1 FILLER_62_873 ();
 sg13g2_fill_1 FILLER_62_889 ();
 sg13g2_fill_1 FILLER_62_895 ();
 sg13g2_decap_4 FILLER_62_906 ();
 sg13g2_fill_1 FILLER_62_910 ();
 sg13g2_decap_8 FILLER_62_920 ();
 sg13g2_decap_8 FILLER_62_927 ();
 sg13g2_decap_8 FILLER_62_934 ();
 sg13g2_decap_4 FILLER_62_941 ();
 sg13g2_fill_2 FILLER_62_949 ();
 sg13g2_decap_4 FILLER_62_956 ();
 sg13g2_decap_8 FILLER_62_979 ();
 sg13g2_decap_8 FILLER_62_986 ();
 sg13g2_fill_2 FILLER_62_993 ();
 sg13g2_fill_1 FILLER_62_1003 ();
 sg13g2_decap_8 FILLER_62_1009 ();
 sg13g2_fill_2 FILLER_62_1016 ();
 sg13g2_fill_1 FILLER_62_1018 ();
 sg13g2_fill_2 FILLER_62_1031 ();
 sg13g2_decap_8 FILLER_62_1055 ();
 sg13g2_decap_8 FILLER_62_1062 ();
 sg13g2_decap_4 FILLER_62_1069 ();
 sg13g2_fill_2 FILLER_62_1073 ();
 sg13g2_fill_1 FILLER_62_1092 ();
 sg13g2_decap_4 FILLER_62_1098 ();
 sg13g2_fill_1 FILLER_62_1102 ();
 sg13g2_fill_2 FILLER_62_1115 ();
 sg13g2_decap_8 FILLER_62_1122 ();
 sg13g2_decap_8 FILLER_62_1129 ();
 sg13g2_decap_8 FILLER_62_1136 ();
 sg13g2_fill_1 FILLER_62_1143 ();
 sg13g2_fill_2 FILLER_62_1148 ();
 sg13g2_decap_8 FILLER_62_1155 ();
 sg13g2_fill_2 FILLER_62_1162 ();
 sg13g2_decap_8 FILLER_62_1168 ();
 sg13g2_decap_8 FILLER_62_1175 ();
 sg13g2_decap_8 FILLER_62_1182 ();
 sg13g2_decap_8 FILLER_62_1189 ();
 sg13g2_decap_8 FILLER_62_1196 ();
 sg13g2_decap_4 FILLER_62_1203 ();
 sg13g2_fill_2 FILLER_62_1207 ();
 sg13g2_decap_8 FILLER_62_1217 ();
 sg13g2_decap_8 FILLER_62_1224 ();
 sg13g2_decap_8 FILLER_62_1231 ();
 sg13g2_fill_2 FILLER_62_1238 ();
 sg13g2_decap_8 FILLER_62_1246 ();
 sg13g2_decap_8 FILLER_62_1253 ();
 sg13g2_decap_8 FILLER_62_1260 ();
 sg13g2_fill_2 FILLER_62_1267 ();
 sg13g2_fill_1 FILLER_62_1269 ();
 sg13g2_decap_8 FILLER_62_1279 ();
 sg13g2_decap_4 FILLER_62_1286 ();
 sg13g2_fill_2 FILLER_62_1294 ();
 sg13g2_decap_8 FILLER_62_1300 ();
 sg13g2_decap_8 FILLER_62_1307 ();
 sg13g2_fill_1 FILLER_62_1314 ();
 sg13g2_decap_4 FILLER_62_1318 ();
 sg13g2_fill_2 FILLER_62_1322 ();
 sg13g2_fill_2 FILLER_62_1332 ();
 sg13g2_decap_8 FILLER_62_1339 ();
 sg13g2_fill_2 FILLER_62_1346 ();
 sg13g2_fill_1 FILLER_62_1352 ();
 sg13g2_fill_1 FILLER_62_1382 ();
 sg13g2_decap_8 FILLER_62_1388 ();
 sg13g2_fill_2 FILLER_62_1395 ();
 sg13g2_fill_1 FILLER_62_1397 ();
 sg13g2_decap_8 FILLER_62_1431 ();
 sg13g2_decap_8 FILLER_62_1438 ();
 sg13g2_decap_8 FILLER_62_1445 ();
 sg13g2_fill_2 FILLER_62_1452 ();
 sg13g2_fill_1 FILLER_62_1454 ();
 sg13g2_fill_2 FILLER_62_1477 ();
 sg13g2_decap_4 FILLER_62_1485 ();
 sg13g2_fill_2 FILLER_62_1489 ();
 sg13g2_decap_8 FILLER_62_1495 ();
 sg13g2_decap_8 FILLER_62_1502 ();
 sg13g2_fill_1 FILLER_62_1528 ();
 sg13g2_fill_2 FILLER_62_1537 ();
 sg13g2_fill_1 FILLER_62_1543 ();
 sg13g2_decap_4 FILLER_62_1558 ();
 sg13g2_fill_2 FILLER_62_1562 ();
 sg13g2_decap_8 FILLER_62_1577 ();
 sg13g2_decap_8 FILLER_62_1584 ();
 sg13g2_decap_8 FILLER_62_1591 ();
 sg13g2_decap_8 FILLER_62_1598 ();
 sg13g2_fill_2 FILLER_62_1605 ();
 sg13g2_fill_2 FILLER_62_1637 ();
 sg13g2_decap_8 FILLER_62_1644 ();
 sg13g2_decap_8 FILLER_62_1651 ();
 sg13g2_fill_1 FILLER_62_1658 ();
 sg13g2_decap_4 FILLER_62_1667 ();
 sg13g2_decap_8 FILLER_62_1679 ();
 sg13g2_decap_8 FILLER_62_1686 ();
 sg13g2_decap_4 FILLER_62_1693 ();
 sg13g2_fill_1 FILLER_62_1697 ();
 sg13g2_fill_2 FILLER_62_1708 ();
 sg13g2_fill_1 FILLER_62_1710 ();
 sg13g2_decap_8 FILLER_62_1714 ();
 sg13g2_decap_8 FILLER_62_1764 ();
 sg13g2_fill_2 FILLER_62_1771 ();
 sg13g2_fill_1 FILLER_62_1773 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_fill_2 FILLER_63_35 ();
 sg13g2_fill_1 FILLER_63_37 ();
 sg13g2_decap_4 FILLER_63_43 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_fill_1 FILLER_63_77 ();
 sg13g2_decap_4 FILLER_63_82 ();
 sg13g2_fill_1 FILLER_63_91 ();
 sg13g2_fill_2 FILLER_63_101 ();
 sg13g2_fill_1 FILLER_63_103 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_fill_2 FILLER_63_133 ();
 sg13g2_decap_4 FILLER_63_158 ();
 sg13g2_fill_2 FILLER_63_162 ();
 sg13g2_decap_8 FILLER_63_173 ();
 sg13g2_decap_8 FILLER_63_180 ();
 sg13g2_decap_8 FILLER_63_187 ();
 sg13g2_decap_8 FILLER_63_194 ();
 sg13g2_decap_4 FILLER_63_201 ();
 sg13g2_fill_2 FILLER_63_210 ();
 sg13g2_decap_4 FILLER_63_219 ();
 sg13g2_decap_4 FILLER_63_233 ();
 sg13g2_fill_2 FILLER_63_254 ();
 sg13g2_fill_1 FILLER_63_256 ();
 sg13g2_fill_2 FILLER_63_262 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_fill_1 FILLER_63_284 ();
 sg13g2_decap_8 FILLER_63_301 ();
 sg13g2_decap_8 FILLER_63_308 ();
 sg13g2_fill_2 FILLER_63_315 ();
 sg13g2_decap_4 FILLER_63_322 ();
 sg13g2_fill_1 FILLER_63_326 ();
 sg13g2_fill_1 FILLER_63_332 ();
 sg13g2_fill_1 FILLER_63_340 ();
 sg13g2_decap_8 FILLER_63_346 ();
 sg13g2_decap_8 FILLER_63_363 ();
 sg13g2_decap_8 FILLER_63_370 ();
 sg13g2_decap_8 FILLER_63_377 ();
 sg13g2_decap_8 FILLER_63_384 ();
 sg13g2_fill_1 FILLER_63_391 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_decap_4 FILLER_63_409 ();
 sg13g2_fill_1 FILLER_63_423 ();
 sg13g2_decap_8 FILLER_63_433 ();
 sg13g2_decap_8 FILLER_63_440 ();
 sg13g2_decap_8 FILLER_63_447 ();
 sg13g2_decap_8 FILLER_63_454 ();
 sg13g2_decap_8 FILLER_63_461 ();
 sg13g2_decap_8 FILLER_63_468 ();
 sg13g2_fill_2 FILLER_63_510 ();
 sg13g2_fill_1 FILLER_63_512 ();
 sg13g2_decap_4 FILLER_63_518 ();
 sg13g2_fill_2 FILLER_63_522 ();
 sg13g2_decap_8 FILLER_63_529 ();
 sg13g2_decap_8 FILLER_63_536 ();
 sg13g2_decap_8 FILLER_63_543 ();
 sg13g2_fill_1 FILLER_63_550 ();
 sg13g2_decap_8 FILLER_63_555 ();
 sg13g2_decap_8 FILLER_63_562 ();
 sg13g2_fill_2 FILLER_63_569 ();
 sg13g2_fill_1 FILLER_63_571 ();
 sg13g2_decap_8 FILLER_63_586 ();
 sg13g2_decap_8 FILLER_63_593 ();
 sg13g2_decap_8 FILLER_63_600 ();
 sg13g2_decap_8 FILLER_63_607 ();
 sg13g2_decap_8 FILLER_63_614 ();
 sg13g2_decap_8 FILLER_63_621 ();
 sg13g2_decap_8 FILLER_63_628 ();
 sg13g2_decap_4 FILLER_63_635 ();
 sg13g2_fill_2 FILLER_63_644 ();
 sg13g2_fill_1 FILLER_63_646 ();
 sg13g2_fill_2 FILLER_63_655 ();
 sg13g2_decap_8 FILLER_63_661 ();
 sg13g2_fill_2 FILLER_63_668 ();
 sg13g2_fill_1 FILLER_63_670 ();
 sg13g2_decap_8 FILLER_63_697 ();
 sg13g2_decap_8 FILLER_63_704 ();
 sg13g2_decap_8 FILLER_63_711 ();
 sg13g2_decap_8 FILLER_63_718 ();
 sg13g2_decap_8 FILLER_63_725 ();
 sg13g2_fill_1 FILLER_63_732 ();
 sg13g2_decap_4 FILLER_63_751 ();
 sg13g2_fill_1 FILLER_63_755 ();
 sg13g2_decap_8 FILLER_63_769 ();
 sg13g2_decap_8 FILLER_63_776 ();
 sg13g2_fill_1 FILLER_63_783 ();
 sg13g2_decap_8 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_decap_8 FILLER_63_812 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_decap_8 FILLER_63_840 ();
 sg13g2_fill_2 FILLER_63_847 ();
 sg13g2_fill_1 FILLER_63_849 ();
 sg13g2_decap_8 FILLER_63_855 ();
 sg13g2_decap_8 FILLER_63_862 ();
 sg13g2_decap_8 FILLER_63_869 ();
 sg13g2_decap_8 FILLER_63_876 ();
 sg13g2_fill_1 FILLER_63_898 ();
 sg13g2_decap_8 FILLER_63_917 ();
 sg13g2_decap_4 FILLER_63_924 ();
 sg13g2_fill_2 FILLER_63_928 ();
 sg13g2_decap_4 FILLER_63_934 ();
 sg13g2_decap_8 FILLER_63_950 ();
 sg13g2_decap_8 FILLER_63_962 ();
 sg13g2_fill_1 FILLER_63_972 ();
 sg13g2_decap_8 FILLER_63_982 ();
 sg13g2_fill_2 FILLER_63_989 ();
 sg13g2_fill_1 FILLER_63_991 ();
 sg13g2_decap_8 FILLER_63_996 ();
 sg13g2_decap_8 FILLER_63_1003 ();
 sg13g2_decap_8 FILLER_63_1010 ();
 sg13g2_decap_4 FILLER_63_1017 ();
 sg13g2_fill_1 FILLER_63_1021 ();
 sg13g2_fill_2 FILLER_63_1030 ();
 sg13g2_fill_1 FILLER_63_1032 ();
 sg13g2_decap_8 FILLER_63_1052 ();
 sg13g2_decap_8 FILLER_63_1059 ();
 sg13g2_decap_8 FILLER_63_1066 ();
 sg13g2_decap_8 FILLER_63_1073 ();
 sg13g2_fill_1 FILLER_63_1094 ();
 sg13g2_fill_2 FILLER_63_1109 ();
 sg13g2_fill_1 FILLER_63_1111 ();
 sg13g2_decap_4 FILLER_63_1129 ();
 sg13g2_fill_2 FILLER_63_1140 ();
 sg13g2_fill_1 FILLER_63_1142 ();
 sg13g2_fill_1 FILLER_63_1152 ();
 sg13g2_fill_1 FILLER_63_1156 ();
 sg13g2_decap_4 FILLER_63_1188 ();
 sg13g2_fill_2 FILLER_63_1192 ();
 sg13g2_decap_8 FILLER_63_1198 ();
 sg13g2_fill_2 FILLER_63_1205 ();
 sg13g2_fill_1 FILLER_63_1207 ();
 sg13g2_decap_8 FILLER_63_1212 ();
 sg13g2_decap_8 FILLER_63_1219 ();
 sg13g2_decap_8 FILLER_63_1226 ();
 sg13g2_decap_8 FILLER_63_1255 ();
 sg13g2_decap_8 FILLER_63_1262 ();
 sg13g2_decap_8 FILLER_63_1269 ();
 sg13g2_decap_4 FILLER_63_1276 ();
 sg13g2_decap_8 FILLER_63_1300 ();
 sg13g2_fill_1 FILLER_63_1307 ();
 sg13g2_fill_2 FILLER_63_1313 ();
 sg13g2_decap_8 FILLER_63_1319 ();
 sg13g2_fill_1 FILLER_63_1326 ();
 sg13g2_decap_8 FILLER_63_1335 ();
 sg13g2_decap_8 FILLER_63_1342 ();
 sg13g2_decap_8 FILLER_63_1349 ();
 sg13g2_fill_2 FILLER_63_1356 ();
 sg13g2_fill_1 FILLER_63_1358 ();
 sg13g2_decap_8 FILLER_63_1363 ();
 sg13g2_fill_1 FILLER_63_1370 ();
 sg13g2_decap_8 FILLER_63_1375 ();
 sg13g2_decap_8 FILLER_63_1382 ();
 sg13g2_decap_8 FILLER_63_1389 ();
 sg13g2_decap_4 FILLER_63_1396 ();
 sg13g2_decap_8 FILLER_63_1408 ();
 sg13g2_decap_8 FILLER_63_1415 ();
 sg13g2_decap_8 FILLER_63_1422 ();
 sg13g2_decap_8 FILLER_63_1429 ();
 sg13g2_decap_8 FILLER_63_1436 ();
 sg13g2_decap_4 FILLER_63_1443 ();
 sg13g2_fill_1 FILLER_63_1459 ();
 sg13g2_fill_2 FILLER_63_1471 ();
 sg13g2_fill_1 FILLER_63_1485 ();
 sg13g2_fill_2 FILLER_63_1493 ();
 sg13g2_fill_1 FILLER_63_1495 ();
 sg13g2_decap_4 FILLER_63_1501 ();
 sg13g2_fill_2 FILLER_63_1509 ();
 sg13g2_decap_4 FILLER_63_1516 ();
 sg13g2_fill_2 FILLER_63_1520 ();
 sg13g2_decap_8 FILLER_63_1525 ();
 sg13g2_fill_2 FILLER_63_1532 ();
 sg13g2_decap_8 FILLER_63_1540 ();
 sg13g2_fill_1 FILLER_63_1553 ();
 sg13g2_fill_1 FILLER_63_1558 ();
 sg13g2_fill_2 FILLER_63_1571 ();
 sg13g2_fill_1 FILLER_63_1573 ();
 sg13g2_decap_8 FILLER_63_1579 ();
 sg13g2_decap_8 FILLER_63_1586 ();
 sg13g2_decap_8 FILLER_63_1593 ();
 sg13g2_decap_8 FILLER_63_1600 ();
 sg13g2_decap_8 FILLER_63_1607 ();
 sg13g2_fill_1 FILLER_63_1614 ();
 sg13g2_decap_8 FILLER_63_1619 ();
 sg13g2_decap_8 FILLER_63_1626 ();
 sg13g2_fill_2 FILLER_63_1633 ();
 sg13g2_decap_8 FILLER_63_1638 ();
 sg13g2_decap_8 FILLER_63_1645 ();
 sg13g2_decap_8 FILLER_63_1652 ();
 sg13g2_decap_8 FILLER_63_1659 ();
 sg13g2_decap_8 FILLER_63_1666 ();
 sg13g2_decap_8 FILLER_63_1673 ();
 sg13g2_decap_8 FILLER_63_1680 ();
 sg13g2_decap_8 FILLER_63_1687 ();
 sg13g2_decap_8 FILLER_63_1694 ();
 sg13g2_decap_8 FILLER_63_1701 ();
 sg13g2_decap_8 FILLER_63_1708 ();
 sg13g2_decap_8 FILLER_63_1724 ();
 sg13g2_fill_2 FILLER_63_1731 ();
 sg13g2_decap_8 FILLER_63_1737 ();
 sg13g2_decap_8 FILLER_63_1744 ();
 sg13g2_decap_8 FILLER_63_1751 ();
 sg13g2_decap_8 FILLER_63_1758 ();
 sg13g2_decap_8 FILLER_63_1765 ();
 sg13g2_fill_2 FILLER_63_1772 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_4 FILLER_64_35 ();
 sg13g2_fill_1 FILLER_64_44 ();
 sg13g2_decap_4 FILLER_64_49 ();
 sg13g2_decap_4 FILLER_64_68 ();
 sg13g2_fill_1 FILLER_64_77 ();
 sg13g2_fill_1 FILLER_64_83 ();
 sg13g2_decap_4 FILLER_64_102 ();
 sg13g2_fill_1 FILLER_64_106 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_fill_2 FILLER_64_147 ();
 sg13g2_fill_1 FILLER_64_149 ();
 sg13g2_decap_4 FILLER_64_161 ();
 sg13g2_fill_2 FILLER_64_165 ();
 sg13g2_fill_2 FILLER_64_172 ();
 sg13g2_decap_4 FILLER_64_184 ();
 sg13g2_fill_1 FILLER_64_188 ();
 sg13g2_fill_2 FILLER_64_195 ();
 sg13g2_decap_4 FILLER_64_202 ();
 sg13g2_fill_2 FILLER_64_206 ();
 sg13g2_decap_8 FILLER_64_218 ();
 sg13g2_decap_8 FILLER_64_225 ();
 sg13g2_decap_8 FILLER_64_232 ();
 sg13g2_decap_4 FILLER_64_239 ();
 sg13g2_decap_8 FILLER_64_256 ();
 sg13g2_decap_8 FILLER_64_263 ();
 sg13g2_decap_8 FILLER_64_270 ();
 sg13g2_decap_8 FILLER_64_277 ();
 sg13g2_decap_8 FILLER_64_292 ();
 sg13g2_decap_8 FILLER_64_299 ();
 sg13g2_decap_8 FILLER_64_306 ();
 sg13g2_decap_4 FILLER_64_313 ();
 sg13g2_fill_2 FILLER_64_326 ();
 sg13g2_fill_1 FILLER_64_328 ();
 sg13g2_decap_8 FILLER_64_342 ();
 sg13g2_decap_8 FILLER_64_349 ();
 sg13g2_fill_2 FILLER_64_356 ();
 sg13g2_decap_8 FILLER_64_370 ();
 sg13g2_decap_8 FILLER_64_377 ();
 sg13g2_decap_4 FILLER_64_384 ();
 sg13g2_decap_4 FILLER_64_393 ();
 sg13g2_decap_4 FILLER_64_407 ();
 sg13g2_fill_2 FILLER_64_411 ();
 sg13g2_decap_8 FILLER_64_421 ();
 sg13g2_decap_4 FILLER_64_436 ();
 sg13g2_fill_2 FILLER_64_440 ();
 sg13g2_decap_8 FILLER_64_447 ();
 sg13g2_decap_8 FILLER_64_454 ();
 sg13g2_decap_4 FILLER_64_461 ();
 sg13g2_decap_8 FILLER_64_473 ();
 sg13g2_decap_8 FILLER_64_480 ();
 sg13g2_fill_1 FILLER_64_487 ();
 sg13g2_decap_4 FILLER_64_492 ();
 sg13g2_fill_1 FILLER_64_496 ();
 sg13g2_fill_2 FILLER_64_502 ();
 sg13g2_fill_1 FILLER_64_504 ();
 sg13g2_decap_8 FILLER_64_516 ();
 sg13g2_fill_2 FILLER_64_523 ();
 sg13g2_fill_1 FILLER_64_525 ();
 sg13g2_decap_4 FILLER_64_556 ();
 sg13g2_decap_8 FILLER_64_591 ();
 sg13g2_decap_4 FILLER_64_598 ();
 sg13g2_decap_8 FILLER_64_642 ();
 sg13g2_decap_8 FILLER_64_649 ();
 sg13g2_decap_8 FILLER_64_656 ();
 sg13g2_decap_4 FILLER_64_663 ();
 sg13g2_decap_8 FILLER_64_680 ();
 sg13g2_decap_8 FILLER_64_687 ();
 sg13g2_decap_8 FILLER_64_694 ();
 sg13g2_fill_2 FILLER_64_701 ();
 sg13g2_decap_8 FILLER_64_749 ();
 sg13g2_decap_4 FILLER_64_787 ();
 sg13g2_fill_2 FILLER_64_791 ();
 sg13g2_fill_2 FILLER_64_796 ();
 sg13g2_decap_8 FILLER_64_828 ();
 sg13g2_fill_1 FILLER_64_835 ();
 sg13g2_fill_1 FILLER_64_846 ();
 sg13g2_decap_8 FILLER_64_877 ();
 sg13g2_decap_8 FILLER_64_884 ();
 sg13g2_decap_4 FILLER_64_891 ();
 sg13g2_fill_1 FILLER_64_895 ();
 sg13g2_decap_8 FILLER_64_908 ();
 sg13g2_decap_8 FILLER_64_915 ();
 sg13g2_decap_4 FILLER_64_922 ();
 sg13g2_fill_2 FILLER_64_926 ();
 sg13g2_fill_2 FILLER_64_933 ();
 sg13g2_fill_1 FILLER_64_935 ();
 sg13g2_decap_8 FILLER_64_943 ();
 sg13g2_decap_8 FILLER_64_950 ();
 sg13g2_decap_8 FILLER_64_957 ();
 sg13g2_decap_8 FILLER_64_964 ();
 sg13g2_fill_1 FILLER_64_971 ();
 sg13g2_decap_8 FILLER_64_976 ();
 sg13g2_decap_4 FILLER_64_983 ();
 sg13g2_decap_4 FILLER_64_997 ();
 sg13g2_fill_1 FILLER_64_1001 ();
 sg13g2_decap_8 FILLER_64_1007 ();
 sg13g2_fill_2 FILLER_64_1014 ();
 sg13g2_decap_4 FILLER_64_1029 ();
 sg13g2_fill_1 FILLER_64_1033 ();
 sg13g2_decap_8 FILLER_64_1044 ();
 sg13g2_fill_1 FILLER_64_1051 ();
 sg13g2_decap_4 FILLER_64_1065 ();
 sg13g2_decap_8 FILLER_64_1074 ();
 sg13g2_decap_4 FILLER_64_1081 ();
 sg13g2_fill_2 FILLER_64_1085 ();
 sg13g2_decap_8 FILLER_64_1096 ();
 sg13g2_decap_4 FILLER_64_1103 ();
 sg13g2_fill_1 FILLER_64_1107 ();
 sg13g2_fill_2 FILLER_64_1120 ();
 sg13g2_decap_8 FILLER_64_1132 ();
 sg13g2_decap_4 FILLER_64_1139 ();
 sg13g2_fill_1 FILLER_64_1143 ();
 sg13g2_fill_2 FILLER_64_1147 ();
 sg13g2_decap_8 FILLER_64_1157 ();
 sg13g2_decap_8 FILLER_64_1164 ();
 sg13g2_fill_1 FILLER_64_1171 ();
 sg13g2_decap_8 FILLER_64_1176 ();
 sg13g2_decap_4 FILLER_64_1183 ();
 sg13g2_decap_8 FILLER_64_1218 ();
 sg13g2_decap_8 FILLER_64_1225 ();
 sg13g2_fill_1 FILLER_64_1232 ();
 sg13g2_decap_8 FILLER_64_1243 ();
 sg13g2_decap_8 FILLER_64_1250 ();
 sg13g2_fill_2 FILLER_64_1257 ();
 sg13g2_fill_1 FILLER_64_1259 ();
 sg13g2_decap_8 FILLER_64_1264 ();
 sg13g2_decap_8 FILLER_64_1271 ();
 sg13g2_decap_8 FILLER_64_1278 ();
 sg13g2_fill_1 FILLER_64_1285 ();
 sg13g2_fill_1 FILLER_64_1291 ();
 sg13g2_decap_8 FILLER_64_1318 ();
 sg13g2_decap_4 FILLER_64_1325 ();
 sg13g2_fill_2 FILLER_64_1329 ();
 sg13g2_fill_1 FILLER_64_1345 ();
 sg13g2_decap_8 FILLER_64_1351 ();
 sg13g2_fill_2 FILLER_64_1358 ();
 sg13g2_fill_1 FILLER_64_1360 ();
 sg13g2_decap_4 FILLER_64_1393 ();
 sg13g2_fill_2 FILLER_64_1397 ();
 sg13g2_fill_2 FILLER_64_1436 ();
 sg13g2_fill_1 FILLER_64_1438 ();
 sg13g2_fill_1 FILLER_64_1463 ();
 sg13g2_fill_2 FILLER_64_1486 ();
 sg13g2_decap_8 FILLER_64_1501 ();
 sg13g2_decap_4 FILLER_64_1508 ();
 sg13g2_fill_1 FILLER_64_1512 ();
 sg13g2_fill_1 FILLER_64_1536 ();
 sg13g2_fill_2 FILLER_64_1550 ();
 sg13g2_fill_2 FILLER_64_1557 ();
 sg13g2_decap_8 FILLER_64_1564 ();
 sg13g2_decap_8 FILLER_64_1571 ();
 sg13g2_decap_8 FILLER_64_1578 ();
 sg13g2_decap_8 FILLER_64_1585 ();
 sg13g2_decap_8 FILLER_64_1592 ();
 sg13g2_decap_4 FILLER_64_1599 ();
 sg13g2_fill_1 FILLER_64_1603 ();
 sg13g2_fill_2 FILLER_64_1609 ();
 sg13g2_fill_1 FILLER_64_1611 ();
 sg13g2_fill_2 FILLER_64_1623 ();
 sg13g2_fill_1 FILLER_64_1625 ();
 sg13g2_fill_1 FILLER_64_1634 ();
 sg13g2_decap_4 FILLER_64_1645 ();
 sg13g2_fill_1 FILLER_64_1649 ();
 sg13g2_decap_4 FILLER_64_1656 ();
 sg13g2_fill_1 FILLER_64_1660 ();
 sg13g2_decap_4 FILLER_64_1664 ();
 sg13g2_fill_1 FILLER_64_1668 ();
 sg13g2_decap_8 FILLER_64_1699 ();
 sg13g2_decap_8 FILLER_64_1724 ();
 sg13g2_decap_8 FILLER_64_1731 ();
 sg13g2_fill_2 FILLER_64_1738 ();
 sg13g2_fill_1 FILLER_64_1740 ();
 sg13g2_decap_8 FILLER_64_1754 ();
 sg13g2_decap_8 FILLER_64_1761 ();
 sg13g2_decap_4 FILLER_64_1768 ();
 sg13g2_fill_2 FILLER_64_1772 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_4 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_43 ();
 sg13g2_decap_4 FILLER_65_54 ();
 sg13g2_fill_2 FILLER_65_58 ();
 sg13g2_fill_2 FILLER_65_65 ();
 sg13g2_fill_2 FILLER_65_78 ();
 sg13g2_fill_1 FILLER_65_90 ();
 sg13g2_fill_2 FILLER_65_96 ();
 sg13g2_decap_4 FILLER_65_103 ();
 sg13g2_fill_2 FILLER_65_122 ();
 sg13g2_decap_8 FILLER_65_128 ();
 sg13g2_fill_2 FILLER_65_135 ();
 sg13g2_decap_4 FILLER_65_150 ();
 sg13g2_decap_8 FILLER_65_159 ();
 sg13g2_decap_8 FILLER_65_166 ();
 sg13g2_fill_1 FILLER_65_177 ();
 sg13g2_fill_2 FILLER_65_186 ();
 sg13g2_fill_1 FILLER_65_188 ();
 sg13g2_fill_2 FILLER_65_194 ();
 sg13g2_decap_8 FILLER_65_200 ();
 sg13g2_decap_4 FILLER_65_207 ();
 sg13g2_fill_2 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_236 ();
 sg13g2_decap_4 FILLER_65_243 ();
 sg13g2_fill_2 FILLER_65_247 ();
 sg13g2_fill_2 FILLER_65_253 ();
 sg13g2_fill_1 FILLER_65_255 ();
 sg13g2_fill_2 FILLER_65_264 ();
 sg13g2_fill_2 FILLER_65_274 ();
 sg13g2_fill_1 FILLER_65_276 ();
 sg13g2_fill_2 FILLER_65_293 ();
 sg13g2_decap_8 FILLER_65_300 ();
 sg13g2_decap_4 FILLER_65_307 ();
 sg13g2_decap_8 FILLER_65_316 ();
 sg13g2_fill_2 FILLER_65_355 ();
 sg13g2_fill_1 FILLER_65_357 ();
 sg13g2_fill_1 FILLER_65_368 ();
 sg13g2_fill_1 FILLER_65_381 ();
 sg13g2_decap_4 FILLER_65_392 ();
 sg13g2_fill_1 FILLER_65_396 ();
 sg13g2_decap_8 FILLER_65_409 ();
 sg13g2_decap_8 FILLER_65_416 ();
 sg13g2_decap_4 FILLER_65_423 ();
 sg13g2_fill_1 FILLER_65_427 ();
 sg13g2_decap_8 FILLER_65_451 ();
 sg13g2_decap_8 FILLER_65_458 ();
 sg13g2_decap_8 FILLER_65_465 ();
 sg13g2_decap_4 FILLER_65_472 ();
 sg13g2_decap_4 FILLER_65_482 ();
 sg13g2_decap_4 FILLER_65_490 ();
 sg13g2_fill_1 FILLER_65_494 ();
 sg13g2_decap_8 FILLER_65_498 ();
 sg13g2_decap_8 FILLER_65_505 ();
 sg13g2_decap_8 FILLER_65_512 ();
 sg13g2_decap_8 FILLER_65_519 ();
 sg13g2_decap_8 FILLER_65_526 ();
 sg13g2_fill_2 FILLER_65_533 ();
 sg13g2_decap_8 FILLER_65_539 ();
 sg13g2_decap_8 FILLER_65_551 ();
 sg13g2_decap_8 FILLER_65_558 ();
 sg13g2_fill_1 FILLER_65_565 ();
 sg13g2_fill_2 FILLER_65_569 ();
 sg13g2_fill_1 FILLER_65_571 ();
 sg13g2_decap_8 FILLER_65_576 ();
 sg13g2_decap_4 FILLER_65_583 ();
 sg13g2_fill_1 FILLER_65_587 ();
 sg13g2_fill_2 FILLER_65_601 ();
 sg13g2_decap_8 FILLER_65_607 ();
 sg13g2_fill_2 FILLER_65_614 ();
 sg13g2_decap_8 FILLER_65_620 ();
 sg13g2_decap_8 FILLER_65_627 ();
 sg13g2_fill_1 FILLER_65_634 ();
 sg13g2_fill_1 FILLER_65_646 ();
 sg13g2_decap_8 FILLER_65_685 ();
 sg13g2_decap_8 FILLER_65_692 ();
 sg13g2_decap_8 FILLER_65_699 ();
 sg13g2_decap_8 FILLER_65_706 ();
 sg13g2_decap_8 FILLER_65_713 ();
 sg13g2_fill_2 FILLER_65_724 ();
 sg13g2_fill_1 FILLER_65_726 ();
 sg13g2_fill_2 FILLER_65_751 ();
 sg13g2_decap_4 FILLER_65_761 ();
 sg13g2_fill_2 FILLER_65_765 ();
 sg13g2_decap_8 FILLER_65_771 ();
 sg13g2_decap_8 FILLER_65_778 ();
 sg13g2_decap_8 FILLER_65_785 ();
 sg13g2_decap_8 FILLER_65_792 ();
 sg13g2_decap_8 FILLER_65_799 ();
 sg13g2_decap_8 FILLER_65_810 ();
 sg13g2_decap_8 FILLER_65_817 ();
 sg13g2_decap_8 FILLER_65_824 ();
 sg13g2_decap_8 FILLER_65_831 ();
 sg13g2_decap_8 FILLER_65_838 ();
 sg13g2_decap_8 FILLER_65_845 ();
 sg13g2_fill_2 FILLER_65_852 ();
 sg13g2_decap_8 FILLER_65_858 ();
 sg13g2_decap_8 FILLER_65_865 ();
 sg13g2_decap_8 FILLER_65_872 ();
 sg13g2_decap_8 FILLER_65_883 ();
 sg13g2_decap_8 FILLER_65_890 ();
 sg13g2_decap_4 FILLER_65_897 ();
 sg13g2_decap_8 FILLER_65_904 ();
 sg13g2_decap_4 FILLER_65_911 ();
 sg13g2_fill_2 FILLER_65_915 ();
 sg13g2_fill_1 FILLER_65_936 ();
 sg13g2_decap_8 FILLER_65_943 ();
 sg13g2_fill_2 FILLER_65_950 ();
 sg13g2_fill_1 FILLER_65_952 ();
 sg13g2_fill_2 FILLER_65_962 ();
 sg13g2_decap_8 FILLER_65_986 ();
 sg13g2_decap_4 FILLER_65_993 ();
 sg13g2_fill_1 FILLER_65_997 ();
 sg13g2_decap_4 FILLER_65_1009 ();
 sg13g2_fill_2 FILLER_65_1013 ();
 sg13g2_decap_8 FILLER_65_1040 ();
 sg13g2_decap_4 FILLER_65_1047 ();
 sg13g2_fill_1 FILLER_65_1051 ();
 sg13g2_fill_1 FILLER_65_1065 ();
 sg13g2_decap_4 FILLER_65_1084 ();
 sg13g2_fill_2 FILLER_65_1088 ();
 sg13g2_decap_8 FILLER_65_1099 ();
 sg13g2_fill_2 FILLER_65_1106 ();
 sg13g2_decap_8 FILLER_65_1123 ();
 sg13g2_decap_8 FILLER_65_1130 ();
 sg13g2_decap_8 FILLER_65_1137 ();
 sg13g2_fill_2 FILLER_65_1144 ();
 sg13g2_fill_1 FILLER_65_1146 ();
 sg13g2_decap_8 FILLER_65_1157 ();
 sg13g2_fill_2 FILLER_65_1170 ();
 sg13g2_fill_1 FILLER_65_1172 ();
 sg13g2_decap_8 FILLER_65_1177 ();
 sg13g2_fill_2 FILLER_65_1184 ();
 sg13g2_fill_1 FILLER_65_1186 ();
 sg13g2_decap_8 FILLER_65_1203 ();
 sg13g2_decap_8 FILLER_65_1210 ();
 sg13g2_decap_4 FILLER_65_1217 ();
 sg13g2_fill_2 FILLER_65_1221 ();
 sg13g2_fill_1 FILLER_65_1238 ();
 sg13g2_fill_2 FILLER_65_1252 ();
 sg13g2_fill_2 FILLER_65_1258 ();
 sg13g2_fill_1 FILLER_65_1260 ();
 sg13g2_decap_8 FILLER_65_1270 ();
 sg13g2_decap_8 FILLER_65_1277 ();
 sg13g2_decap_8 FILLER_65_1284 ();
 sg13g2_decap_8 FILLER_65_1291 ();
 sg13g2_fill_1 FILLER_65_1298 ();
 sg13g2_decap_8 FILLER_65_1311 ();
 sg13g2_decap_8 FILLER_65_1318 ();
 sg13g2_decap_8 FILLER_65_1325 ();
 sg13g2_decap_8 FILLER_65_1332 ();
 sg13g2_decap_8 FILLER_65_1339 ();
 sg13g2_fill_1 FILLER_65_1346 ();
 sg13g2_decap_8 FILLER_65_1351 ();
 sg13g2_decap_4 FILLER_65_1358 ();
 sg13g2_fill_2 FILLER_65_1362 ();
 sg13g2_decap_8 FILLER_65_1368 ();
 sg13g2_decap_8 FILLER_65_1375 ();
 sg13g2_decap_8 FILLER_65_1382 ();
 sg13g2_fill_1 FILLER_65_1389 ();
 sg13g2_fill_2 FILLER_65_1393 ();
 sg13g2_decap_8 FILLER_65_1411 ();
 sg13g2_decap_8 FILLER_65_1418 ();
 sg13g2_fill_2 FILLER_65_1425 ();
 sg13g2_fill_2 FILLER_65_1448 ();
 sg13g2_fill_2 FILLER_65_1454 ();
 sg13g2_fill_2 FILLER_65_1467 ();
 sg13g2_fill_2 FILLER_65_1503 ();
 sg13g2_fill_1 FILLER_65_1505 ();
 sg13g2_fill_1 FILLER_65_1514 ();
 sg13g2_decap_8 FILLER_65_1525 ();
 sg13g2_decap_8 FILLER_65_1564 ();
 sg13g2_decap_8 FILLER_65_1571 ();
 sg13g2_decap_8 FILLER_65_1578 ();
 sg13g2_decap_8 FILLER_65_1585 ();
 sg13g2_decap_8 FILLER_65_1592 ();
 sg13g2_decap_4 FILLER_65_1608 ();
 sg13g2_decap_8 FILLER_65_1620 ();
 sg13g2_fill_1 FILLER_65_1631 ();
 sg13g2_decap_4 FILLER_65_1636 ();
 sg13g2_fill_1 FILLER_65_1674 ();
 sg13g2_decap_8 FILLER_65_1692 ();
 sg13g2_fill_2 FILLER_65_1699 ();
 sg13g2_fill_1 FILLER_65_1701 ();
 sg13g2_decap_4 FILLER_65_1705 ();
 sg13g2_decap_8 FILLER_65_1717 ();
 sg13g2_decap_8 FILLER_65_1724 ();
 sg13g2_fill_1 FILLER_65_1731 ();
 sg13g2_fill_1 FILLER_65_1735 ();
 sg13g2_decap_8 FILLER_65_1762 ();
 sg13g2_decap_4 FILLER_65_1769 ();
 sg13g2_fill_1 FILLER_65_1773 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_fill_1 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_39 ();
 sg13g2_decap_8 FILLER_66_46 ();
 sg13g2_decap_8 FILLER_66_53 ();
 sg13g2_decap_8 FILLER_66_60 ();
 sg13g2_decap_8 FILLER_66_67 ();
 sg13g2_decap_8 FILLER_66_74 ();
 sg13g2_fill_1 FILLER_66_81 ();
 sg13g2_fill_1 FILLER_66_90 ();
 sg13g2_fill_2 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_fill_2 FILLER_66_124 ();
 sg13g2_fill_1 FILLER_66_130 ();
 sg13g2_fill_1 FILLER_66_136 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_4 FILLER_66_182 ();
 sg13g2_fill_1 FILLER_66_186 ();
 sg13g2_fill_1 FILLER_66_191 ();
 sg13g2_fill_2 FILLER_66_202 ();
 sg13g2_fill_2 FILLER_66_209 ();
 sg13g2_fill_2 FILLER_66_220 ();
 sg13g2_decap_4 FILLER_66_226 ();
 sg13g2_fill_2 FILLER_66_230 ();
 sg13g2_decap_8 FILLER_66_237 ();
 sg13g2_decap_8 FILLER_66_244 ();
 sg13g2_decap_8 FILLER_66_251 ();
 sg13g2_decap_8 FILLER_66_258 ();
 sg13g2_fill_2 FILLER_66_265 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_decap_4 FILLER_66_272 ();
 sg13g2_fill_2 FILLER_66_276 ();
 sg13g2_decap_4 FILLER_66_282 ();
 sg13g2_decap_8 FILLER_66_299 ();
 sg13g2_fill_1 FILLER_66_306 ();
 sg13g2_decap_4 FILLER_66_311 ();
 sg13g2_decap_8 FILLER_66_319 ();
 sg13g2_fill_1 FILLER_66_326 ();
 sg13g2_fill_1 FILLER_66_345 ();
 sg13g2_fill_2 FILLER_66_354 ();
 sg13g2_fill_1 FILLER_66_361 ();
 sg13g2_decap_4 FILLER_66_366 ();
 sg13g2_fill_1 FILLER_66_382 ();
 sg13g2_fill_2 FILLER_66_386 ();
 sg13g2_fill_2 FILLER_66_393 ();
 sg13g2_fill_2 FILLER_66_403 ();
 sg13g2_decap_8 FILLER_66_426 ();
 sg13g2_decap_8 FILLER_66_433 ();
 sg13g2_decap_8 FILLER_66_440 ();
 sg13g2_decap_8 FILLER_66_447 ();
 sg13g2_decap_8 FILLER_66_454 ();
 sg13g2_decap_8 FILLER_66_461 ();
 sg13g2_decap_8 FILLER_66_468 ();
 sg13g2_fill_2 FILLER_66_475 ();
 sg13g2_fill_1 FILLER_66_477 ();
 sg13g2_decap_8 FILLER_66_509 ();
 sg13g2_fill_1 FILLER_66_516 ();
 sg13g2_decap_8 FILLER_66_543 ();
 sg13g2_decap_4 FILLER_66_550 ();
 sg13g2_decap_4 FILLER_66_564 ();
 sg13g2_fill_1 FILLER_66_568 ();
 sg13g2_decap_8 FILLER_66_573 ();
 sg13g2_fill_1 FILLER_66_580 ();
 sg13g2_decap_4 FILLER_66_590 ();
 sg13g2_fill_1 FILLER_66_594 ();
 sg13g2_decap_8 FILLER_66_621 ();
 sg13g2_decap_8 FILLER_66_628 ();
 sg13g2_fill_1 FILLER_66_635 ();
 sg13g2_fill_1 FILLER_66_662 ();
 sg13g2_decap_8 FILLER_66_676 ();
 sg13g2_decap_8 FILLER_66_683 ();
 sg13g2_decap_8 FILLER_66_690 ();
 sg13g2_decap_8 FILLER_66_697 ();
 sg13g2_decap_8 FILLER_66_704 ();
 sg13g2_fill_1 FILLER_66_711 ();
 sg13g2_decap_8 FILLER_66_716 ();
 sg13g2_decap_8 FILLER_66_723 ();
 sg13g2_decap_8 FILLER_66_730 ();
 sg13g2_fill_2 FILLER_66_737 ();
 sg13g2_fill_1 FILLER_66_739 ();
 sg13g2_decap_8 FILLER_66_756 ();
 sg13g2_decap_8 FILLER_66_763 ();
 sg13g2_fill_2 FILLER_66_770 ();
 sg13g2_fill_1 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_777 ();
 sg13g2_decap_8 FILLER_66_784 ();
 sg13g2_fill_1 FILLER_66_795 ();
 sg13g2_decap_8 FILLER_66_804 ();
 sg13g2_decap_4 FILLER_66_811 ();
 sg13g2_fill_1 FILLER_66_826 ();
 sg13g2_decap_8 FILLER_66_832 ();
 sg13g2_fill_1 FILLER_66_839 ();
 sg13g2_fill_1 FILLER_66_845 ();
 sg13g2_decap_8 FILLER_66_855 ();
 sg13g2_decap_8 FILLER_66_862 ();
 sg13g2_fill_1 FILLER_66_869 ();
 sg13g2_decap_4 FILLER_66_900 ();
 sg13g2_fill_1 FILLER_66_904 ();
 sg13g2_fill_1 FILLER_66_911 ();
 sg13g2_decap_8 FILLER_66_930 ();
 sg13g2_fill_1 FILLER_66_937 ();
 sg13g2_decap_8 FILLER_66_952 ();
 sg13g2_decap_4 FILLER_66_959 ();
 sg13g2_fill_1 FILLER_66_963 ();
 sg13g2_decap_8 FILLER_66_978 ();
 sg13g2_decap_8 FILLER_66_985 ();
 sg13g2_decap_4 FILLER_66_992 ();
 sg13g2_fill_2 FILLER_66_996 ();
 sg13g2_fill_2 FILLER_66_1014 ();
 sg13g2_decap_8 FILLER_66_1042 ();
 sg13g2_decap_8 FILLER_66_1049 ();
 sg13g2_decap_4 FILLER_66_1056 ();
 sg13g2_decap_8 FILLER_66_1065 ();
 sg13g2_decap_8 FILLER_66_1072 ();
 sg13g2_fill_1 FILLER_66_1079 ();
 sg13g2_decap_8 FILLER_66_1085 ();
 sg13g2_fill_2 FILLER_66_1092 ();
 sg13g2_decap_8 FILLER_66_1103 ();
 sg13g2_decap_8 FILLER_66_1110 ();
 sg13g2_decap_8 FILLER_66_1117 ();
 sg13g2_decap_8 FILLER_66_1124 ();
 sg13g2_decap_4 FILLER_66_1131 ();
 sg13g2_decap_8 FILLER_66_1141 ();
 sg13g2_decap_8 FILLER_66_1148 ();
 sg13g2_fill_1 FILLER_66_1155 ();
 sg13g2_decap_4 FILLER_66_1161 ();
 sg13g2_fill_1 FILLER_66_1165 ();
 sg13g2_decap_8 FILLER_66_1192 ();
 sg13g2_decap_8 FILLER_66_1225 ();
 sg13g2_fill_2 FILLER_66_1232 ();
 sg13g2_decap_8 FILLER_66_1239 ();
 sg13g2_decap_8 FILLER_66_1246 ();
 sg13g2_fill_1 FILLER_66_1253 ();
 sg13g2_decap_8 FILLER_66_1259 ();
 sg13g2_decap_8 FILLER_66_1266 ();
 sg13g2_decap_8 FILLER_66_1273 ();
 sg13g2_decap_8 FILLER_66_1280 ();
 sg13g2_decap_8 FILLER_66_1287 ();
 sg13g2_decap_8 FILLER_66_1294 ();
 sg13g2_decap_8 FILLER_66_1301 ();
 sg13g2_fill_1 FILLER_66_1318 ();
 sg13g2_fill_1 FILLER_66_1340 ();
 sg13g2_decap_8 FILLER_66_1349 ();
 sg13g2_decap_8 FILLER_66_1356 ();
 sg13g2_decap_8 FILLER_66_1363 ();
 sg13g2_decap_8 FILLER_66_1370 ();
 sg13g2_decap_4 FILLER_66_1377 ();
 sg13g2_fill_1 FILLER_66_1381 ();
 sg13g2_decap_8 FILLER_66_1408 ();
 sg13g2_decap_4 FILLER_66_1415 ();
 sg13g2_fill_2 FILLER_66_1419 ();
 sg13g2_fill_1 FILLER_66_1451 ();
 sg13g2_fill_2 FILLER_66_1457 ();
 sg13g2_decap_8 FILLER_66_1488 ();
 sg13g2_decap_8 FILLER_66_1495 ();
 sg13g2_fill_2 FILLER_66_1502 ();
 sg13g2_fill_2 FILLER_66_1513 ();
 sg13g2_fill_1 FILLER_66_1515 ();
 sg13g2_fill_2 FILLER_66_1534 ();
 sg13g2_fill_1 FILLER_66_1541 ();
 sg13g2_fill_2 FILLER_66_1549 ();
 sg13g2_decap_4 FILLER_66_1556 ();
 sg13g2_fill_2 FILLER_66_1560 ();
 sg13g2_fill_2 FILLER_66_1568 ();
 sg13g2_decap_8 FILLER_66_1605 ();
 sg13g2_decap_4 FILLER_66_1612 ();
 sg13g2_fill_2 FILLER_66_1616 ();
 sg13g2_decap_8 FILLER_66_1636 ();
 sg13g2_decap_4 FILLER_66_1643 ();
 sg13g2_decap_8 FILLER_66_1651 ();
 sg13g2_decap_8 FILLER_66_1658 ();
 sg13g2_fill_1 FILLER_66_1665 ();
 sg13g2_decap_8 FILLER_66_1670 ();
 sg13g2_decap_8 FILLER_66_1677 ();
 sg13g2_decap_8 FILLER_66_1684 ();
 sg13g2_decap_8 FILLER_66_1691 ();
 sg13g2_decap_4 FILLER_66_1698 ();
 sg13g2_decap_8 FILLER_66_1707 ();
 sg13g2_decap_8 FILLER_66_1714 ();
 sg13g2_decap_8 FILLER_66_1721 ();
 sg13g2_decap_4 FILLER_66_1728 ();
 sg13g2_decap_4 FILLER_66_1737 ();
 sg13g2_decap_8 FILLER_66_1745 ();
 sg13g2_decap_8 FILLER_66_1752 ();
 sg13g2_decap_8 FILLER_66_1759 ();
 sg13g2_decap_8 FILLER_66_1766 ();
 sg13g2_fill_1 FILLER_66_1773 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_54 ();
 sg13g2_decap_8 FILLER_67_61 ();
 sg13g2_decap_8 FILLER_67_68 ();
 sg13g2_decap_8 FILLER_67_75 ();
 sg13g2_decap_8 FILLER_67_82 ();
 sg13g2_fill_2 FILLER_67_89 ();
 sg13g2_decap_4 FILLER_67_96 ();
 sg13g2_fill_1 FILLER_67_100 ();
 sg13g2_decap_8 FILLER_67_106 ();
 sg13g2_decap_8 FILLER_67_113 ();
 sg13g2_decap_8 FILLER_67_120 ();
 sg13g2_decap_8 FILLER_67_127 ();
 sg13g2_decap_8 FILLER_67_134 ();
 sg13g2_fill_2 FILLER_67_141 ();
 sg13g2_decap_8 FILLER_67_148 ();
 sg13g2_decap_4 FILLER_67_155 ();
 sg13g2_fill_2 FILLER_67_159 ();
 sg13g2_decap_8 FILLER_67_164 ();
 sg13g2_decap_4 FILLER_67_176 ();
 sg13g2_decap_8 FILLER_67_184 ();
 sg13g2_fill_2 FILLER_67_191 ();
 sg13g2_fill_1 FILLER_67_193 ();
 sg13g2_decap_8 FILLER_67_198 ();
 sg13g2_fill_1 FILLER_67_205 ();
 sg13g2_fill_1 FILLER_67_211 ();
 sg13g2_decap_8 FILLER_67_221 ();
 sg13g2_decap_4 FILLER_67_228 ();
 sg13g2_fill_2 FILLER_67_232 ();
 sg13g2_fill_1 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_274 ();
 sg13g2_fill_1 FILLER_67_289 ();
 sg13g2_fill_2 FILLER_67_293 ();
 sg13g2_fill_2 FILLER_67_305 ();
 sg13g2_fill_1 FILLER_67_307 ();
 sg13g2_decap_4 FILLER_67_320 ();
 sg13g2_fill_2 FILLER_67_324 ();
 sg13g2_fill_2 FILLER_67_335 ();
 sg13g2_fill_2 FILLER_67_341 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_fill_1 FILLER_67_371 ();
 sg13g2_fill_2 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_394 ();
 sg13g2_fill_2 FILLER_67_401 ();
 sg13g2_fill_1 FILLER_67_403 ();
 sg13g2_decap_4 FILLER_67_409 ();
 sg13g2_fill_2 FILLER_67_413 ();
 sg13g2_decap_8 FILLER_67_419 ();
 sg13g2_decap_8 FILLER_67_426 ();
 sg13g2_decap_8 FILLER_67_439 ();
 sg13g2_decap_8 FILLER_67_446 ();
 sg13g2_decap_8 FILLER_67_453 ();
 sg13g2_decap_8 FILLER_67_460 ();
 sg13g2_decap_8 FILLER_67_467 ();
 sg13g2_decap_4 FILLER_67_474 ();
 sg13g2_fill_2 FILLER_67_478 ();
 sg13g2_decap_8 FILLER_67_485 ();
 sg13g2_decap_8 FILLER_67_492 ();
 sg13g2_decap_4 FILLER_67_499 ();
 sg13g2_fill_2 FILLER_67_521 ();
 sg13g2_fill_1 FILLER_67_523 ();
 sg13g2_decap_8 FILLER_67_550 ();
 sg13g2_decap_4 FILLER_67_557 ();
 sg13g2_fill_1 FILLER_67_561 ();
 sg13g2_decap_8 FILLER_67_588 ();
 sg13g2_decap_8 FILLER_67_595 ();
 sg13g2_decap_8 FILLER_67_602 ();
 sg13g2_decap_8 FILLER_67_609 ();
 sg13g2_decap_8 FILLER_67_616 ();
 sg13g2_decap_8 FILLER_67_623 ();
 sg13g2_decap_4 FILLER_67_630 ();
 sg13g2_fill_2 FILLER_67_639 ();
 sg13g2_decap_8 FILLER_67_644 ();
 sg13g2_decap_8 FILLER_67_651 ();
 sg13g2_decap_8 FILLER_67_658 ();
 sg13g2_decap_8 FILLER_67_665 ();
 sg13g2_decap_8 FILLER_67_672 ();
 sg13g2_decap_4 FILLER_67_679 ();
 sg13g2_fill_2 FILLER_67_683 ();
 sg13g2_fill_2 FILLER_67_689 ();
 sg13g2_fill_1 FILLER_67_691 ();
 sg13g2_fill_2 FILLER_67_702 ();
 sg13g2_fill_1 FILLER_67_704 ();
 sg13g2_decap_8 FILLER_67_731 ();
 sg13g2_fill_1 FILLER_67_738 ();
 sg13g2_decap_8 FILLER_67_742 ();
 sg13g2_fill_2 FILLER_67_749 ();
 sg13g2_fill_1 FILLER_67_751 ();
 sg13g2_decap_4 FILLER_67_755 ();
 sg13g2_fill_2 FILLER_67_759 ();
 sg13g2_fill_2 FILLER_67_792 ();
 sg13g2_decap_8 FILLER_67_801 ();
 sg13g2_decap_8 FILLER_67_808 ();
 sg13g2_decap_8 FILLER_67_840 ();
 sg13g2_decap_4 FILLER_67_847 ();
 sg13g2_decap_8 FILLER_67_856 ();
 sg13g2_decap_8 FILLER_67_871 ();
 sg13g2_decap_8 FILLER_67_878 ();
 sg13g2_decap_8 FILLER_67_885 ();
 sg13g2_decap_8 FILLER_67_892 ();
 sg13g2_decap_8 FILLER_67_899 ();
 sg13g2_decap_8 FILLER_67_906 ();
 sg13g2_decap_8 FILLER_67_918 ();
 sg13g2_decap_8 FILLER_67_925 ();
 sg13g2_decap_8 FILLER_67_932 ();
 sg13g2_decap_8 FILLER_67_939 ();
 sg13g2_fill_1 FILLER_67_946 ();
 sg13g2_decap_4 FILLER_67_958 ();
 sg13g2_decap_8 FILLER_67_965 ();
 sg13g2_fill_2 FILLER_67_972 ();
 sg13g2_decap_8 FILLER_67_978 ();
 sg13g2_decap_8 FILLER_67_985 ();
 sg13g2_decap_8 FILLER_67_992 ();
 sg13g2_decap_8 FILLER_67_999 ();
 sg13g2_decap_8 FILLER_67_1006 ();
 sg13g2_decap_8 FILLER_67_1013 ();
 sg13g2_decap_8 FILLER_67_1020 ();
 sg13g2_decap_8 FILLER_67_1027 ();
 sg13g2_decap_8 FILLER_67_1034 ();
 sg13g2_decap_8 FILLER_67_1041 ();
 sg13g2_decap_8 FILLER_67_1048 ();
 sg13g2_decap_4 FILLER_67_1055 ();
 sg13g2_fill_1 FILLER_67_1059 ();
 sg13g2_fill_1 FILLER_67_1068 ();
 sg13g2_fill_1 FILLER_67_1073 ();
 sg13g2_fill_2 FILLER_67_1083 ();
 sg13g2_fill_1 FILLER_67_1098 ();
 sg13g2_fill_2 FILLER_67_1108 ();
 sg13g2_fill_1 FILLER_67_1110 ();
 sg13g2_decap_8 FILLER_67_1115 ();
 sg13g2_fill_1 FILLER_67_1122 ();
 sg13g2_decap_8 FILLER_67_1128 ();
 sg13g2_decap_8 FILLER_67_1135 ();
 sg13g2_decap_8 FILLER_67_1142 ();
 sg13g2_fill_1 FILLER_67_1149 ();
 sg13g2_decap_8 FILLER_67_1154 ();
 sg13g2_decap_4 FILLER_67_1161 ();
 sg13g2_decap_8 FILLER_67_1170 ();
 sg13g2_decap_8 FILLER_67_1177 ();
 sg13g2_decap_4 FILLER_67_1184 ();
 sg13g2_fill_2 FILLER_67_1188 ();
 sg13g2_decap_8 FILLER_67_1194 ();
 sg13g2_decap_4 FILLER_67_1201 ();
 sg13g2_fill_2 FILLER_67_1205 ();
 sg13g2_decap_8 FILLER_67_1211 ();
 sg13g2_fill_2 FILLER_67_1218 ();
 sg13g2_fill_1 FILLER_67_1220 ();
 sg13g2_decap_8 FILLER_67_1225 ();
 sg13g2_decap_8 FILLER_67_1252 ();
 sg13g2_fill_2 FILLER_67_1259 ();
 sg13g2_fill_2 FILLER_67_1266 ();
 sg13g2_fill_1 FILLER_67_1268 ();
 sg13g2_decap_8 FILLER_67_1273 ();
 sg13g2_decap_8 FILLER_67_1288 ();
 sg13g2_decap_4 FILLER_67_1295 ();
 sg13g2_fill_2 FILLER_67_1326 ();
 sg13g2_decap_8 FILLER_67_1341 ();
 sg13g2_decap_8 FILLER_67_1348 ();
 sg13g2_decap_8 FILLER_67_1355 ();
 sg13g2_fill_2 FILLER_67_1362 ();
 sg13g2_decap_8 FILLER_67_1368 ();
 sg13g2_fill_1 FILLER_67_1384 ();
 sg13g2_decap_8 FILLER_67_1406 ();
 sg13g2_decap_8 FILLER_67_1413 ();
 sg13g2_fill_1 FILLER_67_1420 ();
 sg13g2_fill_1 FILLER_67_1424 ();
 sg13g2_fill_1 FILLER_67_1450 ();
 sg13g2_fill_1 FILLER_67_1455 ();
 sg13g2_fill_1 FILLER_67_1462 ();
 sg13g2_decap_8 FILLER_67_1489 ();
 sg13g2_decap_8 FILLER_67_1496 ();
 sg13g2_fill_1 FILLER_67_1512 ();
 sg13g2_fill_1 FILLER_67_1524 ();
 sg13g2_decap_4 FILLER_67_1556 ();
 sg13g2_fill_2 FILLER_67_1560 ();
 sg13g2_decap_8 FILLER_67_1568 ();
 sg13g2_decap_8 FILLER_67_1575 ();
 sg13g2_decap_8 FILLER_67_1586 ();
 sg13g2_decap_8 FILLER_67_1593 ();
 sg13g2_decap_8 FILLER_67_1600 ();
 sg13g2_decap_8 FILLER_67_1607 ();
 sg13g2_decap_8 FILLER_67_1614 ();
 sg13g2_decap_8 FILLER_67_1621 ();
 sg13g2_decap_4 FILLER_67_1628 ();
 sg13g2_fill_2 FILLER_67_1632 ();
 sg13g2_decap_8 FILLER_67_1637 ();
 sg13g2_decap_4 FILLER_67_1644 ();
 sg13g2_fill_1 FILLER_67_1648 ();
 sg13g2_decap_8 FILLER_67_1655 ();
 sg13g2_decap_8 FILLER_67_1670 ();
 sg13g2_decap_8 FILLER_67_1677 ();
 sg13g2_fill_1 FILLER_67_1684 ();
 sg13g2_fill_1 FILLER_67_1711 ();
 sg13g2_decap_8 FILLER_67_1715 ();
 sg13g2_fill_2 FILLER_67_1722 ();
 sg13g2_fill_1 FILLER_67_1724 ();
 sg13g2_fill_1 FILLER_67_1731 ();
 sg13g2_decap_8 FILLER_67_1747 ();
 sg13g2_decap_8 FILLER_67_1754 ();
 sg13g2_decap_8 FILLER_67_1761 ();
 sg13g2_decap_4 FILLER_67_1768 ();
 sg13g2_fill_2 FILLER_67_1772 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_20 ();
 sg13g2_fill_2 FILLER_68_28 ();
 sg13g2_decap_4 FILLER_68_50 ();
 sg13g2_fill_1 FILLER_68_54 ();
 sg13g2_decap_8 FILLER_68_59 ();
 sg13g2_decap_8 FILLER_68_66 ();
 sg13g2_decap_8 FILLER_68_73 ();
 sg13g2_decap_8 FILLER_68_80 ();
 sg13g2_decap_8 FILLER_68_87 ();
 sg13g2_decap_8 FILLER_68_94 ();
 sg13g2_decap_8 FILLER_68_101 ();
 sg13g2_decap_4 FILLER_68_108 ();
 sg13g2_fill_1 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_117 ();
 sg13g2_fill_2 FILLER_68_124 ();
 sg13g2_fill_1 FILLER_68_126 ();
 sg13g2_fill_2 FILLER_68_156 ();
 sg13g2_decap_8 FILLER_68_170 ();
 sg13g2_decap_8 FILLER_68_177 ();
 sg13g2_decap_8 FILLER_68_184 ();
 sg13g2_decap_8 FILLER_68_191 ();
 sg13g2_fill_2 FILLER_68_198 ();
 sg13g2_fill_1 FILLER_68_200 ();
 sg13g2_fill_1 FILLER_68_211 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_fill_1 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_231 ();
 sg13g2_decap_4 FILLER_68_238 ();
 sg13g2_fill_1 FILLER_68_242 ();
 sg13g2_decap_8 FILLER_68_246 ();
 sg13g2_decap_8 FILLER_68_253 ();
 sg13g2_decap_8 FILLER_68_260 ();
 sg13g2_decap_8 FILLER_68_267 ();
 sg13g2_fill_1 FILLER_68_299 ();
 sg13g2_fill_1 FILLER_68_305 ();
 sg13g2_decap_4 FILLER_68_310 ();
 sg13g2_fill_2 FILLER_68_314 ();
 sg13g2_fill_2 FILLER_68_324 ();
 sg13g2_decap_8 FILLER_68_331 ();
 sg13g2_decap_8 FILLER_68_338 ();
 sg13g2_decap_8 FILLER_68_345 ();
 sg13g2_decap_8 FILLER_68_352 ();
 sg13g2_decap_4 FILLER_68_359 ();
 sg13g2_fill_1 FILLER_68_368 ();
 sg13g2_fill_1 FILLER_68_379 ();
 sg13g2_fill_2 FILLER_68_383 ();
 sg13g2_fill_1 FILLER_68_395 ();
 sg13g2_decap_8 FILLER_68_400 ();
 sg13g2_decap_8 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_68_414 ();
 sg13g2_decap_8 FILLER_68_421 ();
 sg13g2_decap_8 FILLER_68_428 ();
 sg13g2_decap_4 FILLER_68_435 ();
 sg13g2_fill_1 FILLER_68_439 ();
 sg13g2_fill_1 FILLER_68_473 ();
 sg13g2_fill_2 FILLER_68_512 ();
 sg13g2_decap_8 FILLER_68_520 ();
 sg13g2_fill_1 FILLER_68_527 ();
 sg13g2_decap_8 FILLER_68_532 ();
 sg13g2_decap_8 FILLER_68_539 ();
 sg13g2_decap_8 FILLER_68_546 ();
 sg13g2_decap_4 FILLER_68_553 ();
 sg13g2_fill_1 FILLER_68_557 ();
 sg13g2_fill_2 FILLER_68_563 ();
 sg13g2_fill_1 FILLER_68_565 ();
 sg13g2_decap_8 FILLER_68_569 ();
 sg13g2_fill_2 FILLER_68_576 ();
 sg13g2_decap_8 FILLER_68_584 ();
 sg13g2_decap_8 FILLER_68_591 ();
 sg13g2_decap_8 FILLER_68_598 ();
 sg13g2_decap_8 FILLER_68_605 ();
 sg13g2_decap_8 FILLER_68_612 ();
 sg13g2_fill_2 FILLER_68_619 ();
 sg13g2_fill_1 FILLER_68_621 ();
 sg13g2_decap_4 FILLER_68_626 ();
 sg13g2_fill_1 FILLER_68_630 ();
 sg13g2_decap_8 FILLER_68_636 ();
 sg13g2_fill_2 FILLER_68_643 ();
 sg13g2_fill_1 FILLER_68_645 ();
 sg13g2_fill_1 FILLER_68_659 ();
 sg13g2_fill_1 FILLER_68_669 ();
 sg13g2_decap_8 FILLER_68_679 ();
 sg13g2_decap_8 FILLER_68_686 ();
 sg13g2_decap_8 FILLER_68_693 ();
 sg13g2_decap_8 FILLER_68_705 ();
 sg13g2_decap_8 FILLER_68_712 ();
 sg13g2_decap_8 FILLER_68_719 ();
 sg13g2_decap_8 FILLER_68_731 ();
 sg13g2_fill_2 FILLER_68_738 ();
 sg13g2_decap_4 FILLER_68_748 ();
 sg13g2_fill_1 FILLER_68_752 ();
 sg13g2_decap_8 FILLER_68_763 ();
 sg13g2_decap_8 FILLER_68_770 ();
 sg13g2_decap_8 FILLER_68_777 ();
 sg13g2_decap_8 FILLER_68_784 ();
 sg13g2_decap_8 FILLER_68_791 ();
 sg13g2_decap_8 FILLER_68_798 ();
 sg13g2_decap_8 FILLER_68_805 ();
 sg13g2_decap_8 FILLER_68_812 ();
 sg13g2_fill_1 FILLER_68_819 ();
 sg13g2_fill_2 FILLER_68_829 ();
 sg13g2_fill_1 FILLER_68_831 ();
 sg13g2_decap_8 FILLER_68_837 ();
 sg13g2_decap_4 FILLER_68_844 ();
 sg13g2_fill_2 FILLER_68_848 ();
 sg13g2_decap_4 FILLER_68_854 ();
 sg13g2_decap_8 FILLER_68_873 ();
 sg13g2_fill_1 FILLER_68_880 ();
 sg13g2_fill_1 FILLER_68_893 ();
 sg13g2_decap_8 FILLER_68_898 ();
 sg13g2_decap_8 FILLER_68_905 ();
 sg13g2_decap_4 FILLER_68_912 ();
 sg13g2_fill_1 FILLER_68_916 ();
 sg13g2_decap_8 FILLER_68_921 ();
 sg13g2_decap_8 FILLER_68_928 ();
 sg13g2_decap_4 FILLER_68_935 ();
 sg13g2_fill_2 FILLER_68_951 ();
 sg13g2_fill_2 FILLER_68_965 ();
 sg13g2_decap_8 FILLER_68_993 ();
 sg13g2_decap_4 FILLER_68_1000 ();
 sg13g2_fill_2 FILLER_68_1009 ();
 sg13g2_fill_1 FILLER_68_1011 ();
 sg13g2_decap_8 FILLER_68_1016 ();
 sg13g2_decap_8 FILLER_68_1023 ();
 sg13g2_decap_8 FILLER_68_1030 ();
 sg13g2_decap_8 FILLER_68_1037 ();
 sg13g2_decap_8 FILLER_68_1044 ();
 sg13g2_decap_8 FILLER_68_1051 ();
 sg13g2_decap_8 FILLER_68_1058 ();
 sg13g2_decap_8 FILLER_68_1065 ();
 sg13g2_fill_2 FILLER_68_1072 ();
 sg13g2_fill_2 FILLER_68_1089 ();
 sg13g2_fill_2 FILLER_68_1102 ();
 sg13g2_decap_8 FILLER_68_1130 ();
 sg13g2_decap_4 FILLER_68_1137 ();
 sg13g2_fill_2 FILLER_68_1141 ();
 sg13g2_decap_8 FILLER_68_1169 ();
 sg13g2_decap_8 FILLER_68_1176 ();
 sg13g2_fill_1 FILLER_68_1183 ();
 sg13g2_decap_8 FILLER_68_1194 ();
 sg13g2_decap_8 FILLER_68_1201 ();
 sg13g2_decap_8 FILLER_68_1208 ();
 sg13g2_decap_4 FILLER_68_1215 ();
 sg13g2_decap_8 FILLER_68_1250 ();
 sg13g2_decap_4 FILLER_68_1257 ();
 sg13g2_fill_1 FILLER_68_1261 ();
 sg13g2_fill_2 FILLER_68_1318 ();
 sg13g2_fill_1 FILLER_68_1320 ();
 sg13g2_fill_1 FILLER_68_1329 ();
 sg13g2_decap_8 FILLER_68_1339 ();
 sg13g2_decap_8 FILLER_68_1346 ();
 sg13g2_decap_8 FILLER_68_1353 ();
 sg13g2_decap_8 FILLER_68_1360 ();
 sg13g2_fill_2 FILLER_68_1367 ();
 sg13g2_fill_1 FILLER_68_1395 ();
 sg13g2_decap_8 FILLER_68_1422 ();
 sg13g2_fill_1 FILLER_68_1429 ();
 sg13g2_decap_8 FILLER_68_1442 ();
 sg13g2_fill_2 FILLER_68_1449 ();
 sg13g2_fill_1 FILLER_68_1451 ();
 sg13g2_decap_8 FILLER_68_1458 ();
 sg13g2_fill_2 FILLER_68_1465 ();
 sg13g2_fill_1 FILLER_68_1467 ();
 sg13g2_decap_8 FILLER_68_1472 ();
 sg13g2_decap_8 FILLER_68_1479 ();
 sg13g2_decap_8 FILLER_68_1486 ();
 sg13g2_decap_8 FILLER_68_1493 ();
 sg13g2_decap_8 FILLER_68_1500 ();
 sg13g2_decap_8 FILLER_68_1507 ();
 sg13g2_decap_4 FILLER_68_1514 ();
 sg13g2_fill_2 FILLER_68_1518 ();
 sg13g2_fill_1 FILLER_68_1523 ();
 sg13g2_decap_8 FILLER_68_1572 ();
 sg13g2_decap_8 FILLER_68_1579 ();
 sg13g2_decap_4 FILLER_68_1586 ();
 sg13g2_fill_2 FILLER_68_1590 ();
 sg13g2_decap_8 FILLER_68_1596 ();
 sg13g2_decap_8 FILLER_68_1603 ();
 sg13g2_decap_4 FILLER_68_1610 ();
 sg13g2_fill_2 FILLER_68_1618 ();
 sg13g2_fill_1 FILLER_68_1620 ();
 sg13g2_fill_1 FILLER_68_1628 ();
 sg13g2_fill_2 FILLER_68_1632 ();
 sg13g2_fill_1 FILLER_68_1639 ();
 sg13g2_decap_8 FILLER_68_1645 ();
 sg13g2_decap_8 FILLER_68_1652 ();
 sg13g2_fill_2 FILLER_68_1659 ();
 sg13g2_fill_1 FILLER_68_1661 ();
 sg13g2_fill_1 FILLER_68_1692 ();
 sg13g2_decap_8 FILLER_68_1697 ();
 sg13g2_decap_8 FILLER_68_1704 ();
 sg13g2_decap_4 FILLER_68_1711 ();
 sg13g2_fill_1 FILLER_68_1727 ();
 sg13g2_decap_8 FILLER_68_1737 ();
 sg13g2_decap_4 FILLER_68_1744 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_14 ();
 sg13g2_fill_2 FILLER_69_41 ();
 sg13g2_fill_1 FILLER_69_43 ();
 sg13g2_decap_8 FILLER_69_74 ();
 sg13g2_decap_8 FILLER_69_81 ();
 sg13g2_decap_8 FILLER_69_88 ();
 sg13g2_decap_8 FILLER_69_95 ();
 sg13g2_decap_4 FILLER_69_102 ();
 sg13g2_fill_2 FILLER_69_106 ();
 sg13g2_decap_4 FILLER_69_134 ();
 sg13g2_decap_8 FILLER_69_142 ();
 sg13g2_fill_1 FILLER_69_149 ();
 sg13g2_decap_8 FILLER_69_162 ();
 sg13g2_decap_8 FILLER_69_169 ();
 sg13g2_decap_8 FILLER_69_176 ();
 sg13g2_decap_4 FILLER_69_183 ();
 sg13g2_fill_1 FILLER_69_187 ();
 sg13g2_decap_4 FILLER_69_196 ();
 sg13g2_fill_1 FILLER_69_200 ();
 sg13g2_decap_8 FILLER_69_206 ();
 sg13g2_decap_4 FILLER_69_213 ();
 sg13g2_decap_8 FILLER_69_222 ();
 sg13g2_fill_2 FILLER_69_229 ();
 sg13g2_decap_8 FILLER_69_257 ();
 sg13g2_decap_8 FILLER_69_264 ();
 sg13g2_decap_4 FILLER_69_271 ();
 sg13g2_fill_1 FILLER_69_275 ();
 sg13g2_decap_4 FILLER_69_281 ();
 sg13g2_fill_2 FILLER_69_285 ();
 sg13g2_decap_4 FILLER_69_290 ();
 sg13g2_fill_2 FILLER_69_294 ();
 sg13g2_decap_8 FILLER_69_303 ();
 sg13g2_decap_8 FILLER_69_310 ();
 sg13g2_decap_8 FILLER_69_317 ();
 sg13g2_decap_8 FILLER_69_324 ();
 sg13g2_decap_8 FILLER_69_331 ();
 sg13g2_fill_2 FILLER_69_338 ();
 sg13g2_decap_4 FILLER_69_345 ();
 sg13g2_fill_2 FILLER_69_349 ();
 sg13g2_decap_8 FILLER_69_362 ();
 sg13g2_fill_2 FILLER_69_369 ();
 sg13g2_fill_1 FILLER_69_371 ();
 sg13g2_decap_4 FILLER_69_375 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_decap_8 FILLER_69_406 ();
 sg13g2_fill_2 FILLER_69_413 ();
 sg13g2_decap_4 FILLER_69_421 ();
 sg13g2_decap_8 FILLER_69_434 ();
 sg13g2_decap_8 FILLER_69_441 ();
 sg13g2_fill_2 FILLER_69_448 ();
 sg13g2_fill_1 FILLER_69_450 ();
 sg13g2_decap_8 FILLER_69_455 ();
 sg13g2_decap_8 FILLER_69_462 ();
 sg13g2_decap_8 FILLER_69_469 ();
 sg13g2_decap_4 FILLER_69_476 ();
 sg13g2_fill_2 FILLER_69_480 ();
 sg13g2_fill_2 FILLER_69_486 ();
 sg13g2_fill_1 FILLER_69_488 ();
 sg13g2_decap_8 FILLER_69_493 ();
 sg13g2_fill_2 FILLER_69_504 ();
 sg13g2_decap_8 FILLER_69_509 ();
 sg13g2_fill_2 FILLER_69_519 ();
 sg13g2_decap_8 FILLER_69_547 ();
 sg13g2_decap_8 FILLER_69_554 ();
 sg13g2_fill_2 FILLER_69_561 ();
 sg13g2_decap_8 FILLER_69_593 ();
 sg13g2_fill_1 FILLER_69_600 ();
 sg13g2_decap_8 FILLER_69_635 ();
 sg13g2_decap_4 FILLER_69_664 ();
 sg13g2_decap_8 FILLER_69_676 ();
 sg13g2_decap_8 FILLER_69_683 ();
 sg13g2_decap_8 FILLER_69_690 ();
 sg13g2_fill_2 FILLER_69_697 ();
 sg13g2_decap_8 FILLER_69_704 ();
 sg13g2_decap_8 FILLER_69_711 ();
 sg13g2_decap_8 FILLER_69_718 ();
 sg13g2_fill_2 FILLER_69_725 ();
 sg13g2_decap_8 FILLER_69_732 ();
 sg13g2_fill_2 FILLER_69_739 ();
 sg13g2_fill_1 FILLER_69_746 ();
 sg13g2_fill_2 FILLER_69_752 ();
 sg13g2_fill_2 FILLER_69_760 ();
 sg13g2_fill_1 FILLER_69_766 ();
 sg13g2_decap_8 FILLER_69_775 ();
 sg13g2_decap_8 FILLER_69_782 ();
 sg13g2_decap_4 FILLER_69_806 ();
 sg13g2_fill_2 FILLER_69_810 ();
 sg13g2_decap_4 FILLER_69_817 ();
 sg13g2_fill_1 FILLER_69_826 ();
 sg13g2_decap_4 FILLER_69_853 ();
 sg13g2_fill_1 FILLER_69_857 ();
 sg13g2_decap_4 FILLER_69_869 ();
 sg13g2_fill_1 FILLER_69_873 ();
 sg13g2_decap_4 FILLER_69_879 ();
 sg13g2_decap_8 FILLER_69_895 ();
 sg13g2_decap_8 FILLER_69_902 ();
 sg13g2_fill_2 FILLER_69_909 ();
 sg13g2_fill_1 FILLER_69_911 ();
 sg13g2_decap_8 FILLER_69_917 ();
 sg13g2_decap_8 FILLER_69_924 ();
 sg13g2_decap_8 FILLER_69_934 ();
 sg13g2_decap_4 FILLER_69_941 ();
 sg13g2_fill_2 FILLER_69_945 ();
 sg13g2_decap_4 FILLER_69_970 ();
 sg13g2_decap_8 FILLER_69_978 ();
 sg13g2_fill_2 FILLER_69_985 ();
 sg13g2_decap_8 FILLER_69_992 ();
 sg13g2_decap_4 FILLER_69_999 ();
 sg13g2_fill_2 FILLER_69_1003 ();
 sg13g2_decap_4 FILLER_69_1031 ();
 sg13g2_fill_2 FILLER_69_1035 ();
 sg13g2_decap_4 FILLER_69_1040 ();
 sg13g2_fill_2 FILLER_69_1044 ();
 sg13g2_decap_4 FILLER_69_1061 ();
 sg13g2_fill_1 FILLER_69_1090 ();
 sg13g2_decap_8 FILLER_69_1113 ();
 sg13g2_decap_4 FILLER_69_1120 ();
 sg13g2_fill_1 FILLER_69_1124 ();
 sg13g2_decap_8 FILLER_69_1135 ();
 sg13g2_decap_8 FILLER_69_1142 ();
 sg13g2_decap_4 FILLER_69_1149 ();
 sg13g2_fill_1 FILLER_69_1153 ();
 sg13g2_decap_8 FILLER_69_1166 ();
 sg13g2_decap_8 FILLER_69_1173 ();
 sg13g2_fill_2 FILLER_69_1180 ();
 sg13g2_decap_8 FILLER_69_1187 ();
 sg13g2_decap_8 FILLER_69_1194 ();
 sg13g2_decap_8 FILLER_69_1201 ();
 sg13g2_decap_8 FILLER_69_1208 ();
 sg13g2_decap_8 FILLER_69_1215 ();
 sg13g2_decap_4 FILLER_69_1222 ();
 sg13g2_fill_2 FILLER_69_1226 ();
 sg13g2_decap_4 FILLER_69_1246 ();
 sg13g2_fill_1 FILLER_69_1250 ();
 sg13g2_decap_8 FILLER_69_1256 ();
 sg13g2_decap_8 FILLER_69_1263 ();
 sg13g2_decap_8 FILLER_69_1270 ();
 sg13g2_decap_8 FILLER_69_1277 ();
 sg13g2_decap_8 FILLER_69_1284 ();
 sg13g2_decap_8 FILLER_69_1291 ();
 sg13g2_decap_8 FILLER_69_1298 ();
 sg13g2_decap_8 FILLER_69_1305 ();
 sg13g2_decap_8 FILLER_69_1312 ();
 sg13g2_decap_8 FILLER_69_1319 ();
 sg13g2_decap_8 FILLER_69_1331 ();
 sg13g2_decap_8 FILLER_69_1338 ();
 sg13g2_decap_8 FILLER_69_1345 ();
 sg13g2_decap_8 FILLER_69_1352 ();
 sg13g2_decap_8 FILLER_69_1359 ();
 sg13g2_decap_8 FILLER_69_1366 ();
 sg13g2_decap_4 FILLER_69_1373 ();
 sg13g2_decap_8 FILLER_69_1381 ();
 sg13g2_decap_8 FILLER_69_1394 ();
 sg13g2_decap_4 FILLER_69_1401 ();
 sg13g2_fill_1 FILLER_69_1405 ();
 sg13g2_decap_8 FILLER_69_1410 ();
 sg13g2_fill_2 FILLER_69_1417 ();
 sg13g2_fill_1 FILLER_69_1419 ();
 sg13g2_fill_2 FILLER_69_1441 ();
 sg13g2_fill_2 FILLER_69_1450 ();
 sg13g2_decap_8 FILLER_69_1485 ();
 sg13g2_decap_8 FILLER_69_1492 ();
 sg13g2_decap_4 FILLER_69_1499 ();
 sg13g2_fill_2 FILLER_69_1508 ();
 sg13g2_decap_8 FILLER_69_1515 ();
 sg13g2_fill_2 FILLER_69_1522 ();
 sg13g2_fill_1 FILLER_69_1528 ();
 sg13g2_fill_1 FILLER_69_1535 ();
 sg13g2_decap_4 FILLER_69_1548 ();
 sg13g2_fill_2 FILLER_69_1552 ();
 sg13g2_decap_8 FILLER_69_1558 ();
 sg13g2_decap_8 FILLER_69_1565 ();
 sg13g2_decap_8 FILLER_69_1572 ();
 sg13g2_decap_4 FILLER_69_1579 ();
 sg13g2_fill_2 FILLER_69_1583 ();
 sg13g2_fill_1 FILLER_69_1611 ();
 sg13g2_decap_8 FILLER_69_1616 ();
 sg13g2_decap_4 FILLER_69_1623 ();
 sg13g2_fill_2 FILLER_69_1627 ();
 sg13g2_decap_4 FILLER_69_1664 ();
 sg13g2_fill_2 FILLER_69_1668 ();
 sg13g2_decap_8 FILLER_69_1674 ();
 sg13g2_decap_8 FILLER_69_1681 ();
 sg13g2_decap_8 FILLER_69_1688 ();
 sg13g2_decap_8 FILLER_69_1695 ();
 sg13g2_decap_8 FILLER_69_1702 ();
 sg13g2_decap_4 FILLER_69_1709 ();
 sg13g2_fill_1 FILLER_69_1713 ();
 sg13g2_decap_8 FILLER_69_1745 ();
 sg13g2_fill_2 FILLER_69_1752 ();
 sg13g2_fill_1 FILLER_69_1754 ();
 sg13g2_decap_8 FILLER_69_1759 ();
 sg13g2_decap_8 FILLER_69_1766 ();
 sg13g2_fill_1 FILLER_69_1773 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_4 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_32 ();
 sg13g2_fill_1 FILLER_70_39 ();
 sg13g2_decap_4 FILLER_70_64 ();
 sg13g2_decap_8 FILLER_70_72 ();
 sg13g2_decap_8 FILLER_70_79 ();
 sg13g2_decap_8 FILLER_70_86 ();
 sg13g2_decap_8 FILLER_70_93 ();
 sg13g2_decap_8 FILLER_70_113 ();
 sg13g2_decap_8 FILLER_70_120 ();
 sg13g2_decap_8 FILLER_70_127 ();
 sg13g2_decap_8 FILLER_70_134 ();
 sg13g2_decap_8 FILLER_70_141 ();
 sg13g2_decap_8 FILLER_70_148 ();
 sg13g2_decap_8 FILLER_70_155 ();
 sg13g2_fill_2 FILLER_70_162 ();
 sg13g2_fill_1 FILLER_70_164 ();
 sg13g2_fill_2 FILLER_70_180 ();
 sg13g2_decap_8 FILLER_70_187 ();
 sg13g2_fill_2 FILLER_70_194 ();
 sg13g2_fill_1 FILLER_70_200 ();
 sg13g2_fill_1 FILLER_70_206 ();
 sg13g2_decap_8 FILLER_70_212 ();
 sg13g2_decap_8 FILLER_70_219 ();
 sg13g2_decap_8 FILLER_70_226 ();
 sg13g2_decap_4 FILLER_70_233 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_decap_8 FILLER_70_242 ();
 sg13g2_decap_8 FILLER_70_249 ();
 sg13g2_decap_8 FILLER_70_256 ();
 sg13g2_decap_8 FILLER_70_263 ();
 sg13g2_decap_4 FILLER_70_270 ();
 sg13g2_fill_1 FILLER_70_274 ();
 sg13g2_fill_1 FILLER_70_293 ();
 sg13g2_decap_8 FILLER_70_297 ();
 sg13g2_decap_8 FILLER_70_304 ();
 sg13g2_decap_8 FILLER_70_311 ();
 sg13g2_fill_2 FILLER_70_318 ();
 sg13g2_fill_1 FILLER_70_320 ();
 sg13g2_decap_8 FILLER_70_324 ();
 sg13g2_decap_8 FILLER_70_331 ();
 sg13g2_decap_8 FILLER_70_338 ();
 sg13g2_decap_8 FILLER_70_349 ();
 sg13g2_decap_4 FILLER_70_356 ();
 sg13g2_decap_8 FILLER_70_373 ();
 sg13g2_decap_8 FILLER_70_380 ();
 sg13g2_decap_8 FILLER_70_387 ();
 sg13g2_fill_2 FILLER_70_394 ();
 sg13g2_fill_1 FILLER_70_396 ();
 sg13g2_decap_8 FILLER_70_410 ();
 sg13g2_decap_8 FILLER_70_417 ();
 sg13g2_fill_1 FILLER_70_424 ();
 sg13g2_decap_4 FILLER_70_429 ();
 sg13g2_fill_1 FILLER_70_433 ();
 sg13g2_decap_8 FILLER_70_467 ();
 sg13g2_decap_4 FILLER_70_474 ();
 sg13g2_decap_4 FILLER_70_484 ();
 sg13g2_fill_2 FILLER_70_488 ();
 sg13g2_fill_2 FILLER_70_495 ();
 sg13g2_fill_1 FILLER_70_497 ();
 sg13g2_decap_4 FILLER_70_509 ();
 sg13g2_decap_8 FILLER_70_519 ();
 sg13g2_decap_8 FILLER_70_526 ();
 sg13g2_fill_1 FILLER_70_533 ();
 sg13g2_decap_8 FILLER_70_538 ();
 sg13g2_decap_8 FILLER_70_545 ();
 sg13g2_decap_8 FILLER_70_552 ();
 sg13g2_decap_8 FILLER_70_559 ();
 sg13g2_decap_8 FILLER_70_566 ();
 sg13g2_decap_8 FILLER_70_580 ();
 sg13g2_decap_8 FILLER_70_587 ();
 sg13g2_fill_1 FILLER_70_594 ();
 sg13g2_fill_2 FILLER_70_602 ();
 sg13g2_fill_1 FILLER_70_604 ();
 sg13g2_decap_4 FILLER_70_613 ();
 sg13g2_fill_1 FILLER_70_617 ();
 sg13g2_decap_8 FILLER_70_623 ();
 sg13g2_decap_8 FILLER_70_630 ();
 sg13g2_decap_8 FILLER_70_637 ();
 sg13g2_decap_4 FILLER_70_644 ();
 sg13g2_fill_2 FILLER_70_648 ();
 sg13g2_fill_1 FILLER_70_666 ();
 sg13g2_fill_1 FILLER_70_675 ();
 sg13g2_fill_1 FILLER_70_681 ();
 sg13g2_fill_1 FILLER_70_691 ();
 sg13g2_fill_2 FILLER_70_696 ();
 sg13g2_decap_4 FILLER_70_711 ();
 sg13g2_fill_2 FILLER_70_715 ();
 sg13g2_fill_1 FILLER_70_721 ();
 sg13g2_decap_8 FILLER_70_727 ();
 sg13g2_decap_4 FILLER_70_743 ();
 sg13g2_fill_2 FILLER_70_752 ();
 sg13g2_fill_1 FILLER_70_754 ();
 sg13g2_decap_4 FILLER_70_769 ();
 sg13g2_fill_2 FILLER_70_773 ();
 sg13g2_decap_8 FILLER_70_783 ();
 sg13g2_decap_8 FILLER_70_790 ();
 sg13g2_decap_4 FILLER_70_806 ();
 sg13g2_decap_8 FILLER_70_815 ();
 sg13g2_decap_8 FILLER_70_822 ();
 sg13g2_decap_8 FILLER_70_829 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_847 ();
 sg13g2_decap_8 FILLER_70_854 ();
 sg13g2_fill_2 FILLER_70_887 ();
 sg13g2_fill_1 FILLER_70_889 ();
 sg13g2_decap_8 FILLER_70_901 ();
 sg13g2_decap_8 FILLER_70_934 ();
 sg13g2_decap_4 FILLER_70_941 ();
 sg13g2_fill_2 FILLER_70_945 ();
 sg13g2_decap_8 FILLER_70_979 ();
 sg13g2_decap_8 FILLER_70_986 ();
 sg13g2_decap_8 FILLER_70_1007 ();
 sg13g2_fill_2 FILLER_70_1018 ();
 sg13g2_fill_1 FILLER_70_1020 ();
 sg13g2_decap_8 FILLER_70_1026 ();
 sg13g2_decap_8 FILLER_70_1033 ();
 sg13g2_fill_2 FILLER_70_1051 ();
 sg13g2_decap_4 FILLER_70_1058 ();
 sg13g2_decap_8 FILLER_70_1097 ();
 sg13g2_decap_8 FILLER_70_1104 ();
 sg13g2_decap_8 FILLER_70_1111 ();
 sg13g2_decap_4 FILLER_70_1118 ();
 sg13g2_fill_2 FILLER_70_1122 ();
 sg13g2_fill_2 FILLER_70_1150 ();
 sg13g2_fill_1 FILLER_70_1152 ();
 sg13g2_decap_8 FILLER_70_1157 ();
 sg13g2_fill_1 FILLER_70_1164 ();
 sg13g2_decap_8 FILLER_70_1201 ();
 sg13g2_decap_8 FILLER_70_1208 ();
 sg13g2_decap_8 FILLER_70_1215 ();
 sg13g2_decap_8 FILLER_70_1222 ();
 sg13g2_fill_2 FILLER_70_1259 ();
 sg13g2_fill_1 FILLER_70_1261 ();
 sg13g2_decap_4 FILLER_70_1282 ();
 sg13g2_fill_1 FILLER_70_1286 ();
 sg13g2_decap_8 FILLER_70_1313 ();
 sg13g2_decap_4 FILLER_70_1365 ();
 sg13g2_fill_1 FILLER_70_1369 ();
 sg13g2_decap_8 FILLER_70_1374 ();
 sg13g2_decap_8 FILLER_70_1381 ();
 sg13g2_decap_4 FILLER_70_1388 ();
 sg13g2_decap_4 FILLER_70_1423 ();
 sg13g2_fill_2 FILLER_70_1434 ();
 sg13g2_fill_1 FILLER_70_1436 ();
 sg13g2_decap_8 FILLER_70_1442 ();
 sg13g2_fill_2 FILLER_70_1449 ();
 sg13g2_fill_1 FILLER_70_1451 ();
 sg13g2_fill_1 FILLER_70_1459 ();
 sg13g2_decap_8 FILLER_70_1467 ();
 sg13g2_fill_2 FILLER_70_1474 ();
 sg13g2_decap_8 FILLER_70_1482 ();
 sg13g2_fill_2 FILLER_70_1494 ();
 sg13g2_fill_1 FILLER_70_1513 ();
 sg13g2_decap_8 FILLER_70_1558 ();
 sg13g2_decap_4 FILLER_70_1565 ();
 sg13g2_decap_8 FILLER_70_1573 ();
 sg13g2_decap_8 FILLER_70_1580 ();
 sg13g2_decap_8 FILLER_70_1587 ();
 sg13g2_decap_8 FILLER_70_1594 ();
 sg13g2_decap_8 FILLER_70_1601 ();
 sg13g2_decap_4 FILLER_70_1608 ();
 sg13g2_fill_2 FILLER_70_1616 ();
 sg13g2_fill_2 FILLER_70_1626 ();
 sg13g2_fill_1 FILLER_70_1636 ();
 sg13g2_fill_1 FILLER_70_1642 ();
 sg13g2_decap_8 FILLER_70_1647 ();
 sg13g2_decap_4 FILLER_70_1654 ();
 sg13g2_decap_8 FILLER_70_1671 ();
 sg13g2_decap_8 FILLER_70_1678 ();
 sg13g2_decap_8 FILLER_70_1685 ();
 sg13g2_decap_8 FILLER_70_1692 ();
 sg13g2_decap_8 FILLER_70_1699 ();
 sg13g2_decap_4 FILLER_70_1706 ();
 sg13g2_fill_1 FILLER_70_1710 ();
 sg13g2_fill_2 FILLER_70_1721 ();
 sg13g2_decap_8 FILLER_70_1758 ();
 sg13g2_decap_8 FILLER_70_1765 ();
 sg13g2_fill_2 FILLER_70_1772 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_4 FILLER_71_14 ();
 sg13g2_fill_1 FILLER_71_18 ();
 sg13g2_decap_8 FILLER_71_23 ();
 sg13g2_decap_8 FILLER_71_30 ();
 sg13g2_decap_8 FILLER_71_37 ();
 sg13g2_decap_8 FILLER_71_44 ();
 sg13g2_decap_8 FILLER_71_51 ();
 sg13g2_decap_8 FILLER_71_58 ();
 sg13g2_decap_8 FILLER_71_65 ();
 sg13g2_decap_8 FILLER_71_72 ();
 sg13g2_fill_1 FILLER_71_79 ();
 sg13g2_fill_2 FILLER_71_85 ();
 sg13g2_decap_8 FILLER_71_113 ();
 sg13g2_fill_1 FILLER_71_120 ();
 sg13g2_decap_8 FILLER_71_132 ();
 sg13g2_decap_8 FILLER_71_139 ();
 sg13g2_decap_8 FILLER_71_146 ();
 sg13g2_decap_8 FILLER_71_153 ();
 sg13g2_decap_8 FILLER_71_160 ();
 sg13g2_decap_4 FILLER_71_167 ();
 sg13g2_fill_2 FILLER_71_171 ();
 sg13g2_fill_1 FILLER_71_177 ();
 sg13g2_decap_4 FILLER_71_186 ();
 sg13g2_fill_1 FILLER_71_190 ();
 sg13g2_decap_8 FILLER_71_199 ();
 sg13g2_fill_2 FILLER_71_206 ();
 sg13g2_fill_1 FILLER_71_208 ();
 sg13g2_decap_8 FILLER_71_214 ();
 sg13g2_decap_8 FILLER_71_221 ();
 sg13g2_decap_4 FILLER_71_228 ();
 sg13g2_decap_8 FILLER_71_236 ();
 sg13g2_decap_8 FILLER_71_243 ();
 sg13g2_decap_8 FILLER_71_250 ();
 sg13g2_decap_4 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_261 ();
 sg13g2_decap_4 FILLER_71_289 ();
 sg13g2_fill_2 FILLER_71_293 ();
 sg13g2_decap_4 FILLER_71_333 ();
 sg13g2_fill_1 FILLER_71_337 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_fill_2 FILLER_71_378 ();
 sg13g2_fill_1 FILLER_71_380 ();
 sg13g2_decap_4 FILLER_71_410 ();
 sg13g2_decap_8 FILLER_71_444 ();
 sg13g2_decap_8 FILLER_71_451 ();
 sg13g2_decap_8 FILLER_71_458 ();
 sg13g2_decap_8 FILLER_71_465 ();
 sg13g2_decap_8 FILLER_71_472 ();
 sg13g2_decap_8 FILLER_71_479 ();
 sg13g2_decap_8 FILLER_71_486 ();
 sg13g2_decap_8 FILLER_71_493 ();
 sg13g2_fill_2 FILLER_71_500 ();
 sg13g2_fill_1 FILLER_71_502 ();
 sg13g2_decap_4 FILLER_71_506 ();
 sg13g2_fill_1 FILLER_71_510 ();
 sg13g2_decap_8 FILLER_71_515 ();
 sg13g2_decap_8 FILLER_71_522 ();
 sg13g2_decap_4 FILLER_71_529 ();
 sg13g2_fill_1 FILLER_71_533 ();
 sg13g2_decap_8 FILLER_71_537 ();
 sg13g2_fill_1 FILLER_71_544 ();
 sg13g2_decap_8 FILLER_71_549 ();
 sg13g2_decap_4 FILLER_71_556 ();
 sg13g2_decap_4 FILLER_71_565 ();
 sg13g2_fill_2 FILLER_71_569 ();
 sg13g2_decap_8 FILLER_71_623 ();
 sg13g2_decap_8 FILLER_71_630 ();
 sg13g2_decap_8 FILLER_71_637 ();
 sg13g2_decap_4 FILLER_71_648 ();
 sg13g2_decap_8 FILLER_71_657 ();
 sg13g2_decap_8 FILLER_71_664 ();
 sg13g2_decap_8 FILLER_71_671 ();
 sg13g2_decap_4 FILLER_71_678 ();
 sg13g2_fill_2 FILLER_71_682 ();
 sg13g2_fill_1 FILLER_71_694 ();
 sg13g2_fill_2 FILLER_71_703 ();
 sg13g2_decap_8 FILLER_71_713 ();
 sg13g2_fill_2 FILLER_71_737 ();
 sg13g2_fill_1 FILLER_71_739 ();
 sg13g2_fill_2 FILLER_71_748 ();
 sg13g2_fill_2 FILLER_71_760 ();
 sg13g2_decap_8 FILLER_71_774 ();
 sg13g2_decap_8 FILLER_71_781 ();
 sg13g2_decap_8 FILLER_71_788 ();
 sg13g2_fill_2 FILLER_71_795 ();
 sg13g2_decap_8 FILLER_71_823 ();
 sg13g2_decap_8 FILLER_71_830 ();
 sg13g2_decap_8 FILLER_71_837 ();
 sg13g2_decap_8 FILLER_71_848 ();
 sg13g2_decap_8 FILLER_71_855 ();
 sg13g2_decap_4 FILLER_71_862 ();
 sg13g2_fill_1 FILLER_71_870 ();
 sg13g2_decap_8 FILLER_71_883 ();
 sg13g2_decap_8 FILLER_71_890 ();
 sg13g2_decap_8 FILLER_71_897 ();
 sg13g2_decap_8 FILLER_71_904 ();
 sg13g2_fill_2 FILLER_71_911 ();
 sg13g2_fill_1 FILLER_71_913 ();
 sg13g2_decap_8 FILLER_71_918 ();
 sg13g2_decap_8 FILLER_71_925 ();
 sg13g2_decap_8 FILLER_71_932 ();
 sg13g2_decap_8 FILLER_71_939 ();
 sg13g2_decap_8 FILLER_71_946 ();
 sg13g2_decap_8 FILLER_71_953 ();
 sg13g2_decap_4 FILLER_71_964 ();
 sg13g2_fill_1 FILLER_71_968 ();
 sg13g2_decap_8 FILLER_71_982 ();
 sg13g2_fill_1 FILLER_71_989 ();
 sg13g2_decap_4 FILLER_71_1032 ();
 sg13g2_decap_8 FILLER_71_1046 ();
 sg13g2_decap_8 FILLER_71_1053 ();
 sg13g2_decap_8 FILLER_71_1060 ();
 sg13g2_decap_8 FILLER_71_1067 ();
 sg13g2_decap_8 FILLER_71_1074 ();
 sg13g2_decap_8 FILLER_71_1081 ();
 sg13g2_decap_8 FILLER_71_1088 ();
 sg13g2_decap_8 FILLER_71_1113 ();
 sg13g2_decap_4 FILLER_71_1120 ();
 sg13g2_fill_1 FILLER_71_1124 ();
 sg13g2_decap_8 FILLER_71_1137 ();
 sg13g2_decap_8 FILLER_71_1144 ();
 sg13g2_decap_4 FILLER_71_1151 ();
 sg13g2_fill_1 FILLER_71_1155 ();
 sg13g2_decap_4 FILLER_71_1169 ();
 sg13g2_decap_8 FILLER_71_1210 ();
 sg13g2_fill_2 FILLER_71_1217 ();
 sg13g2_decap_8 FILLER_71_1224 ();
 sg13g2_decap_8 FILLER_71_1231 ();
 sg13g2_decap_8 FILLER_71_1238 ();
 sg13g2_decap_8 FILLER_71_1245 ();
 sg13g2_decap_8 FILLER_71_1252 ();
 sg13g2_fill_1 FILLER_71_1259 ();
 sg13g2_fill_1 FILLER_71_1263 ();
 sg13g2_decap_8 FILLER_71_1278 ();
 sg13g2_decap_8 FILLER_71_1285 ();
 sg13g2_decap_4 FILLER_71_1292 ();
 sg13g2_decap_8 FILLER_71_1300 ();
 sg13g2_decap_8 FILLER_71_1307 ();
 sg13g2_decap_4 FILLER_71_1314 ();
 sg13g2_fill_1 FILLER_71_1322 ();
 sg13g2_fill_1 FILLER_71_1328 ();
 sg13g2_decap_8 FILLER_71_1333 ();
 sg13g2_fill_1 FILLER_71_1340 ();
 sg13g2_decap_8 FILLER_71_1392 ();
 sg13g2_decap_8 FILLER_71_1399 ();
 sg13g2_decap_8 FILLER_71_1406 ();
 sg13g2_decap_8 FILLER_71_1413 ();
 sg13g2_decap_8 FILLER_71_1420 ();
 sg13g2_decap_8 FILLER_71_1427 ();
 sg13g2_decap_8 FILLER_71_1434 ();
 sg13g2_decap_4 FILLER_71_1441 ();
 sg13g2_decap_4 FILLER_71_1456 ();
 sg13g2_fill_1 FILLER_71_1460 ();
 sg13g2_decap_4 FILLER_71_1465 ();
 sg13g2_fill_1 FILLER_71_1469 ();
 sg13g2_decap_8 FILLER_71_1473 ();
 sg13g2_decap_8 FILLER_71_1480 ();
 sg13g2_fill_2 FILLER_71_1487 ();
 sg13g2_fill_1 FILLER_71_1489 ();
 sg13g2_decap_4 FILLER_71_1520 ();
 sg13g2_fill_1 FILLER_71_1529 ();
 sg13g2_decap_8 FILLER_71_1534 ();
 sg13g2_decap_8 FILLER_71_1541 ();
 sg13g2_decap_8 FILLER_71_1548 ();
 sg13g2_decap_8 FILLER_71_1555 ();
 sg13g2_fill_1 FILLER_71_1588 ();
 sg13g2_decap_8 FILLER_71_1599 ();
 sg13g2_fill_1 FILLER_71_1606 ();
 sg13g2_decap_8 FILLER_71_1619 ();
 sg13g2_decap_8 FILLER_71_1626 ();
 sg13g2_decap_8 FILLER_71_1633 ();
 sg13g2_decap_8 FILLER_71_1640 ();
 sg13g2_decap_8 FILLER_71_1647 ();
 sg13g2_decap_4 FILLER_71_1654 ();
 sg13g2_decap_8 FILLER_71_1663 ();
 sg13g2_fill_2 FILLER_71_1670 ();
 sg13g2_decap_8 FILLER_71_1676 ();
 sg13g2_decap_8 FILLER_71_1683 ();
 sg13g2_decap_8 FILLER_71_1690 ();
 sg13g2_decap_8 FILLER_71_1697 ();
 sg13g2_decap_8 FILLER_71_1704 ();
 sg13g2_decap_4 FILLER_71_1711 ();
 sg13g2_fill_2 FILLER_71_1727 ();
 sg13g2_decap_8 FILLER_71_1742 ();
 sg13g2_decap_8 FILLER_71_1749 ();
 sg13g2_decap_8 FILLER_71_1756 ();
 sg13g2_decap_8 FILLER_71_1763 ();
 sg13g2_decap_4 FILLER_71_1770 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_14 ();
 sg13g2_decap_4 FILLER_72_46 ();
 sg13g2_decap_4 FILLER_72_61 ();
 sg13g2_fill_2 FILLER_72_65 ();
 sg13g2_decap_8 FILLER_72_72 ();
 sg13g2_decap_8 FILLER_72_79 ();
 sg13g2_decap_8 FILLER_72_86 ();
 sg13g2_fill_2 FILLER_72_93 ();
 sg13g2_decap_8 FILLER_72_99 ();
 sg13g2_decap_8 FILLER_72_106 ();
 sg13g2_decap_8 FILLER_72_113 ();
 sg13g2_fill_1 FILLER_72_120 ();
 sg13g2_decap_4 FILLER_72_155 ();
 sg13g2_decap_8 FILLER_72_162 ();
 sg13g2_fill_2 FILLER_72_169 ();
 sg13g2_fill_1 FILLER_72_171 ();
 sg13g2_fill_2 FILLER_72_183 ();
 sg13g2_fill_1 FILLER_72_190 ();
 sg13g2_fill_2 FILLER_72_209 ();
 sg13g2_fill_2 FILLER_72_223 ();
 sg13g2_fill_2 FILLER_72_251 ();
 sg13g2_fill_2 FILLER_72_257 ();
 sg13g2_decap_8 FILLER_72_285 ();
 sg13g2_decap_8 FILLER_72_292 ();
 sg13g2_decap_8 FILLER_72_299 ();
 sg13g2_fill_2 FILLER_72_306 ();
 sg13g2_decap_8 FILLER_72_331 ();
 sg13g2_decap_8 FILLER_72_338 ();
 sg13g2_decap_8 FILLER_72_345 ();
 sg13g2_decap_8 FILLER_72_352 ();
 sg13g2_decap_8 FILLER_72_359 ();
 sg13g2_decap_8 FILLER_72_366 ();
 sg13g2_decap_8 FILLER_72_373 ();
 sg13g2_decap_4 FILLER_72_380 ();
 sg13g2_fill_2 FILLER_72_384 ();
 sg13g2_decap_8 FILLER_72_390 ();
 sg13g2_decap_8 FILLER_72_400 ();
 sg13g2_decap_8 FILLER_72_407 ();
 sg13g2_decap_8 FILLER_72_414 ();
 sg13g2_decap_4 FILLER_72_421 ();
 sg13g2_fill_2 FILLER_72_425 ();
 sg13g2_decap_8 FILLER_72_432 ();
 sg13g2_decap_8 FILLER_72_439 ();
 sg13g2_fill_1 FILLER_72_446 ();
 sg13g2_decap_8 FILLER_72_451 ();
 sg13g2_decap_8 FILLER_72_462 ();
 sg13g2_decap_8 FILLER_72_469 ();
 sg13g2_decap_8 FILLER_72_476 ();
 sg13g2_decap_8 FILLER_72_483 ();
 sg13g2_decap_8 FILLER_72_490 ();
 sg13g2_decap_8 FILLER_72_497 ();
 sg13g2_decap_8 FILLER_72_530 ();
 sg13g2_fill_1 FILLER_72_537 ();
 sg13g2_decap_8 FILLER_72_564 ();
 sg13g2_decap_4 FILLER_72_571 ();
 sg13g2_fill_2 FILLER_72_575 ();
 sg13g2_decap_8 FILLER_72_581 ();
 sg13g2_fill_2 FILLER_72_588 ();
 sg13g2_fill_1 FILLER_72_590 ();
 sg13g2_decap_8 FILLER_72_596 ();
 sg13g2_decap_8 FILLER_72_603 ();
 sg13g2_decap_8 FILLER_72_610 ();
 sg13g2_decap_8 FILLER_72_617 ();
 sg13g2_decap_8 FILLER_72_624 ();
 sg13g2_decap_8 FILLER_72_631 ();
 sg13g2_decap_8 FILLER_72_638 ();
 sg13g2_fill_2 FILLER_72_645 ();
 sg13g2_decap_4 FILLER_72_651 ();
 sg13g2_fill_2 FILLER_72_655 ();
 sg13g2_decap_8 FILLER_72_665 ();
 sg13g2_decap_4 FILLER_72_672 ();
 sg13g2_fill_2 FILLER_72_676 ();
 sg13g2_decap_4 FILLER_72_683 ();
 sg13g2_fill_1 FILLER_72_687 ();
 sg13g2_decap_8 FILLER_72_692 ();
 sg13g2_decap_8 FILLER_72_699 ();
 sg13g2_decap_8 FILLER_72_706 ();
 sg13g2_decap_8 FILLER_72_713 ();
 sg13g2_fill_2 FILLER_72_720 ();
 sg13g2_fill_1 FILLER_72_722 ();
 sg13g2_decap_8 FILLER_72_727 ();
 sg13g2_decap_8 FILLER_72_734 ();
 sg13g2_fill_1 FILLER_72_741 ();
 sg13g2_decap_8 FILLER_72_782 ();
 sg13g2_decap_8 FILLER_72_789 ();
 sg13g2_decap_8 FILLER_72_796 ();
 sg13g2_fill_1 FILLER_72_803 ();
 sg13g2_decap_8 FILLER_72_808 ();
 sg13g2_decap_8 FILLER_72_815 ();
 sg13g2_decap_4 FILLER_72_822 ();
 sg13g2_fill_1 FILLER_72_826 ();
 sg13g2_decap_4 FILLER_72_832 ();
 sg13g2_fill_1 FILLER_72_836 ();
 sg13g2_fill_2 FILLER_72_863 ();
 sg13g2_fill_2 FILLER_72_879 ();
 sg13g2_decap_4 FILLER_72_886 ();
 sg13g2_decap_8 FILLER_72_894 ();
 sg13g2_decap_8 FILLER_72_901 ();
 sg13g2_decap_8 FILLER_72_908 ();
 sg13g2_decap_4 FILLER_72_915 ();
 sg13g2_fill_2 FILLER_72_919 ();
 sg13g2_decap_8 FILLER_72_952 ();
 sg13g2_decap_8 FILLER_72_959 ();
 sg13g2_decap_8 FILLER_72_966 ();
 sg13g2_decap_8 FILLER_72_973 ();
 sg13g2_decap_8 FILLER_72_980 ();
 sg13g2_decap_4 FILLER_72_987 ();
 sg13g2_fill_2 FILLER_72_991 ();
 sg13g2_decap_4 FILLER_72_998 ();
 sg13g2_decap_8 FILLER_72_1007 ();
 sg13g2_decap_8 FILLER_72_1014 ();
 sg13g2_decap_4 FILLER_72_1021 ();
 sg13g2_fill_1 FILLER_72_1025 ();
 sg13g2_decap_8 FILLER_72_1044 ();
 sg13g2_decap_8 FILLER_72_1061 ();
 sg13g2_decap_8 FILLER_72_1068 ();
 sg13g2_decap_8 FILLER_72_1075 ();
 sg13g2_decap_8 FILLER_72_1082 ();
 sg13g2_decap_8 FILLER_72_1089 ();
 sg13g2_decap_8 FILLER_72_1096 ();
 sg13g2_decap_8 FILLER_72_1112 ();
 sg13g2_decap_8 FILLER_72_1119 ();
 sg13g2_fill_2 FILLER_72_1126 ();
 sg13g2_decap_4 FILLER_72_1132 ();
 sg13g2_fill_2 FILLER_72_1136 ();
 sg13g2_fill_2 FILLER_72_1142 ();
 sg13g2_fill_1 FILLER_72_1144 ();
 sg13g2_decap_8 FILLER_72_1153 ();
 sg13g2_fill_1 FILLER_72_1160 ();
 sg13g2_fill_2 FILLER_72_1165 ();
 sg13g2_fill_1 FILLER_72_1167 ();
 sg13g2_fill_2 FILLER_72_1173 ();
 sg13g2_fill_1 FILLER_72_1175 ();
 sg13g2_decap_8 FILLER_72_1185 ();
 sg13g2_fill_1 FILLER_72_1192 ();
 sg13g2_decap_4 FILLER_72_1207 ();
 sg13g2_fill_2 FILLER_72_1211 ();
 sg13g2_decap_8 FILLER_72_1218 ();
 sg13g2_decap_8 FILLER_72_1225 ();
 sg13g2_decap_8 FILLER_72_1232 ();
 sg13g2_decap_8 FILLER_72_1239 ();
 sg13g2_decap_8 FILLER_72_1246 ();
 sg13g2_fill_1 FILLER_72_1253 ();
 sg13g2_fill_2 FILLER_72_1263 ();
 sg13g2_decap_8 FILLER_72_1279 ();
 sg13g2_decap_8 FILLER_72_1286 ();
 sg13g2_decap_8 FILLER_72_1293 ();
 sg13g2_decap_8 FILLER_72_1300 ();
 sg13g2_decap_8 FILLER_72_1307 ();
 sg13g2_fill_2 FILLER_72_1314 ();
 sg13g2_fill_2 FILLER_72_1320 ();
 sg13g2_fill_1 FILLER_72_1322 ();
 sg13g2_decap_8 FILLER_72_1327 ();
 sg13g2_decap_8 FILLER_72_1334 ();
 sg13g2_fill_2 FILLER_72_1341 ();
 sg13g2_fill_1 FILLER_72_1343 ();
 sg13g2_fill_1 FILLER_72_1359 ();
 sg13g2_decap_8 FILLER_72_1372 ();
 sg13g2_fill_2 FILLER_72_1379 ();
 sg13g2_fill_1 FILLER_72_1381 ();
 sg13g2_decap_8 FILLER_72_1388 ();
 sg13g2_decap_8 FILLER_72_1395 ();
 sg13g2_decap_8 FILLER_72_1402 ();
 sg13g2_decap_8 FILLER_72_1409 ();
 sg13g2_decap_8 FILLER_72_1416 ();
 sg13g2_decap_4 FILLER_72_1423 ();
 sg13g2_decap_8 FILLER_72_1430 ();
 sg13g2_decap_4 FILLER_72_1437 ();
 sg13g2_decap_8 FILLER_72_1480 ();
 sg13g2_decap_4 FILLER_72_1491 ();
 sg13g2_fill_1 FILLER_72_1495 ();
 sg13g2_decap_8 FILLER_72_1500 ();
 sg13g2_decap_4 FILLER_72_1507 ();
 sg13g2_fill_2 FILLER_72_1511 ();
 sg13g2_fill_2 FILLER_72_1522 ();
 sg13g2_fill_1 FILLER_72_1524 ();
 sg13g2_decap_8 FILLER_72_1529 ();
 sg13g2_decap_8 FILLER_72_1536 ();
 sg13g2_decap_8 FILLER_72_1543 ();
 sg13g2_decap_8 FILLER_72_1550 ();
 sg13g2_decap_4 FILLER_72_1557 ();
 sg13g2_fill_2 FILLER_72_1567 ();
 sg13g2_decap_8 FILLER_72_1577 ();
 sg13g2_decap_8 FILLER_72_1584 ();
 sg13g2_decap_8 FILLER_72_1591 ();
 sg13g2_decap_8 FILLER_72_1601 ();
 sg13g2_decap_4 FILLER_72_1608 ();
 sg13g2_fill_2 FILLER_72_1612 ();
 sg13g2_decap_8 FILLER_72_1618 ();
 sg13g2_decap_8 FILLER_72_1625 ();
 sg13g2_decap_8 FILLER_72_1632 ();
 sg13g2_fill_2 FILLER_72_1639 ();
 sg13g2_fill_1 FILLER_72_1641 ();
 sg13g2_decap_4 FILLER_72_1668 ();
 sg13g2_fill_1 FILLER_72_1684 ();
 sg13g2_decap_8 FILLER_72_1693 ();
 sg13g2_fill_1 FILLER_72_1700 ();
 sg13g2_decap_8 FILLER_72_1715 ();
 sg13g2_fill_2 FILLER_72_1722 ();
 sg13g2_decap_8 FILLER_72_1732 ();
 sg13g2_decap_8 FILLER_72_1739 ();
 sg13g2_decap_8 FILLER_72_1746 ();
 sg13g2_decap_8 FILLER_72_1753 ();
 sg13g2_decap_8 FILLER_72_1760 ();
 sg13g2_decap_8 FILLER_72_1767 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_fill_1 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_19 ();
 sg13g2_decap_8 FILLER_73_26 ();
 sg13g2_decap_8 FILLER_73_33 ();
 sg13g2_fill_2 FILLER_73_40 ();
 sg13g2_fill_1 FILLER_73_42 ();
 sg13g2_fill_2 FILLER_73_51 ();
 sg13g2_fill_1 FILLER_73_53 ();
 sg13g2_fill_1 FILLER_73_58 ();
 sg13g2_decap_4 FILLER_73_89 ();
 sg13g2_fill_1 FILLER_73_93 ();
 sg13g2_decap_8 FILLER_73_103 ();
 sg13g2_decap_8 FILLER_73_110 ();
 sg13g2_decap_8 FILLER_73_117 ();
 sg13g2_decap_8 FILLER_73_124 ();
 sg13g2_decap_8 FILLER_73_131 ();
 sg13g2_fill_2 FILLER_73_138 ();
 sg13g2_decap_4 FILLER_73_146 ();
 sg13g2_fill_1 FILLER_73_150 ();
 sg13g2_fill_2 FILLER_73_195 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_223 ();
 sg13g2_fill_1 FILLER_73_230 ();
 sg13g2_decap_8 FILLER_73_234 ();
 sg13g2_decap_4 FILLER_73_245 ();
 sg13g2_fill_1 FILLER_73_249 ();
 sg13g2_fill_2 FILLER_73_274 ();
 sg13g2_fill_2 FILLER_73_286 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_fill_1 FILLER_73_308 ();
 sg13g2_decap_8 FILLER_73_314 ();
 sg13g2_fill_1 FILLER_73_331 ();
 sg13g2_fill_2 FILLER_73_344 ();
 sg13g2_fill_1 FILLER_73_346 ();
 sg13g2_decap_8 FILLER_73_359 ();
 sg13g2_decap_8 FILLER_73_366 ();
 sg13g2_decap_8 FILLER_73_373 ();
 sg13g2_fill_2 FILLER_73_380 ();
 sg13g2_fill_1 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_73_389 ();
 sg13g2_decap_8 FILLER_73_396 ();
 sg13g2_decap_8 FILLER_73_403 ();
 sg13g2_decap_8 FILLER_73_410 ();
 sg13g2_fill_1 FILLER_73_417 ();
 sg13g2_fill_1 FILLER_73_450 ();
 sg13g2_decap_4 FILLER_73_477 ();
 sg13g2_fill_1 FILLER_73_481 ();
 sg13g2_decap_8 FILLER_73_501 ();
 sg13g2_decap_8 FILLER_73_508 ();
 sg13g2_decap_8 FILLER_73_515 ();
 sg13g2_fill_2 FILLER_73_522 ();
 sg13g2_decap_8 FILLER_73_529 ();
 sg13g2_decap_8 FILLER_73_536 ();
 sg13g2_decap_8 FILLER_73_561 ();
 sg13g2_decap_8 FILLER_73_568 ();
 sg13g2_decap_4 FILLER_73_575 ();
 sg13g2_fill_2 FILLER_73_579 ();
 sg13g2_decap_8 FILLER_73_607 ();
 sg13g2_fill_2 FILLER_73_614 ();
 sg13g2_fill_1 FILLER_73_616 ();
 sg13g2_decap_8 FILLER_73_629 ();
 sg13g2_decap_8 FILLER_73_636 ();
 sg13g2_decap_8 FILLER_73_643 ();
 sg13g2_decap_4 FILLER_73_650 ();
 sg13g2_fill_1 FILLER_73_654 ();
 sg13g2_decap_8 FILLER_73_681 ();
 sg13g2_decap_8 FILLER_73_688 ();
 sg13g2_fill_1 FILLER_73_695 ();
 sg13g2_decap_8 FILLER_73_699 ();
 sg13g2_decap_8 FILLER_73_706 ();
 sg13g2_decap_8 FILLER_73_713 ();
 sg13g2_decap_8 FILLER_73_724 ();
 sg13g2_fill_2 FILLER_73_731 ();
 sg13g2_fill_1 FILLER_73_733 ();
 sg13g2_decap_4 FILLER_73_739 ();
 sg13g2_decap_8 FILLER_73_746 ();
 sg13g2_decap_4 FILLER_73_753 ();
 sg13g2_fill_1 FILLER_73_762 ();
 sg13g2_decap_8 FILLER_73_789 ();
 sg13g2_fill_1 FILLER_73_796 ();
 sg13g2_decap_8 FILLER_73_806 ();
 sg13g2_decap_8 FILLER_73_813 ();
 sg13g2_decap_4 FILLER_73_820 ();
 sg13g2_decap_8 FILLER_73_833 ();
 sg13g2_decap_8 FILLER_73_840 ();
 sg13g2_decap_8 FILLER_73_847 ();
 sg13g2_decap_8 FILLER_73_854 ();
 sg13g2_fill_2 FILLER_73_861 ();
 sg13g2_fill_1 FILLER_73_863 ();
 sg13g2_fill_1 FILLER_73_883 ();
 sg13g2_decap_8 FILLER_73_910 ();
 sg13g2_decap_8 FILLER_73_917 ();
 sg13g2_decap_8 FILLER_73_924 ();
 sg13g2_fill_2 FILLER_73_931 ();
 sg13g2_decap_8 FILLER_73_937 ();
 sg13g2_decap_8 FILLER_73_944 ();
 sg13g2_fill_1 FILLER_73_951 ();
 sg13g2_decap_8 FILLER_73_960 ();
 sg13g2_fill_1 FILLER_73_982 ();
 sg13g2_fill_2 FILLER_73_989 ();
 sg13g2_fill_1 FILLER_73_996 ();
 sg13g2_fill_2 FILLER_73_1002 ();
 sg13g2_decap_8 FILLER_73_1010 ();
 sg13g2_decap_8 FILLER_73_1017 ();
 sg13g2_decap_8 FILLER_73_1024 ();
 sg13g2_decap_8 FILLER_73_1031 ();
 sg13g2_decap_8 FILLER_73_1038 ();
 sg13g2_decap_4 FILLER_73_1045 ();
 sg13g2_fill_2 FILLER_73_1049 ();
 sg13g2_fill_2 FILLER_73_1054 ();
 sg13g2_decap_8 FILLER_73_1087 ();
 sg13g2_decap_4 FILLER_73_1094 ();
 sg13g2_fill_2 FILLER_73_1098 ();
 sg13g2_decap_8 FILLER_73_1126 ();
 sg13g2_fill_2 FILLER_73_1133 ();
 sg13g2_fill_1 FILLER_73_1135 ();
 sg13g2_decap_8 FILLER_73_1166 ();
 sg13g2_decap_8 FILLER_73_1173 ();
 sg13g2_fill_1 FILLER_73_1180 ();
 sg13g2_fill_2 FILLER_73_1193 ();
 sg13g2_decap_8 FILLER_73_1199 ();
 sg13g2_decap_8 FILLER_73_1206 ();
 sg13g2_decap_4 FILLER_73_1213 ();
 sg13g2_fill_2 FILLER_73_1217 ();
 sg13g2_decap_8 FILLER_73_1245 ();
 sg13g2_fill_2 FILLER_73_1252 ();
 sg13g2_fill_2 FILLER_73_1258 ();
 sg13g2_fill_2 FILLER_73_1263 ();
 sg13g2_fill_1 FILLER_73_1265 ();
 sg13g2_decap_8 FILLER_73_1272 ();
 sg13g2_decap_8 FILLER_73_1279 ();
 sg13g2_decap_4 FILLER_73_1286 ();
 sg13g2_fill_2 FILLER_73_1290 ();
 sg13g2_decap_8 FILLER_73_1297 ();
 sg13g2_decap_8 FILLER_73_1304 ();
 sg13g2_fill_2 FILLER_73_1311 ();
 sg13g2_fill_1 FILLER_73_1321 ();
 sg13g2_fill_1 FILLER_73_1330 ();
 sg13g2_fill_1 FILLER_73_1337 ();
 sg13g2_fill_2 FILLER_73_1342 ();
 sg13g2_fill_1 FILLER_73_1353 ();
 sg13g2_decap_8 FILLER_73_1359 ();
 sg13g2_decap_8 FILLER_73_1395 ();
 sg13g2_fill_2 FILLER_73_1402 ();
 sg13g2_decap_8 FILLER_73_1408 ();
 sg13g2_decap_8 FILLER_73_1415 ();
 sg13g2_decap_4 FILLER_73_1422 ();
 sg13g2_fill_2 FILLER_73_1426 ();
 sg13g2_decap_8 FILLER_73_1454 ();
 sg13g2_decap_8 FILLER_73_1461 ();
 sg13g2_fill_2 FILLER_73_1468 ();
 sg13g2_decap_4 FILLER_73_1475 ();
 sg13g2_fill_1 FILLER_73_1479 ();
 sg13g2_decap_8 FILLER_73_1489 ();
 sg13g2_decap_4 FILLER_73_1496 ();
 sg13g2_fill_2 FILLER_73_1500 ();
 sg13g2_decap_8 FILLER_73_1517 ();
 sg13g2_decap_8 FILLER_73_1524 ();
 sg13g2_decap_8 FILLER_73_1531 ();
 sg13g2_decap_8 FILLER_73_1538 ();
 sg13g2_fill_2 FILLER_73_1545 ();
 sg13g2_fill_2 FILLER_73_1559 ();
 sg13g2_decap_8 FILLER_73_1564 ();
 sg13g2_decap_8 FILLER_73_1571 ();
 sg13g2_decap_8 FILLER_73_1578 ();
 sg13g2_decap_8 FILLER_73_1599 ();
 sg13g2_decap_8 FILLER_73_1614 ();
 sg13g2_fill_1 FILLER_73_1621 ();
 sg13g2_decap_8 FILLER_73_1627 ();
 sg13g2_decap_8 FILLER_73_1634 ();
 sg13g2_fill_1 FILLER_73_1641 ();
 sg13g2_decap_8 FILLER_73_1645 ();
 sg13g2_decap_8 FILLER_73_1656 ();
 sg13g2_decap_8 FILLER_73_1663 ();
 sg13g2_decap_8 FILLER_73_1670 ();
 sg13g2_decap_8 FILLER_73_1677 ();
 sg13g2_decap_8 FILLER_73_1684 ();
 sg13g2_decap_8 FILLER_73_1691 ();
 sg13g2_decap_8 FILLER_73_1698 ();
 sg13g2_decap_8 FILLER_73_1705 ();
 sg13g2_decap_8 FILLER_73_1712 ();
 sg13g2_decap_8 FILLER_73_1719 ();
 sg13g2_fill_2 FILLER_73_1726 ();
 sg13g2_decap_8 FILLER_73_1741 ();
 sg13g2_decap_8 FILLER_73_1748 ();
 sg13g2_decap_8 FILLER_73_1755 ();
 sg13g2_decap_8 FILLER_73_1762 ();
 sg13g2_decap_4 FILLER_73_1769 ();
 sg13g2_fill_1 FILLER_73_1773 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_4 ();
 sg13g2_fill_1 FILLER_74_32 ();
 sg13g2_fill_1 FILLER_74_46 ();
 sg13g2_fill_2 FILLER_74_59 ();
 sg13g2_fill_1 FILLER_74_61 ();
 sg13g2_decap_4 FILLER_74_66 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_decap_4 FILLER_74_79 ();
 sg13g2_fill_2 FILLER_74_83 ();
 sg13g2_decap_8 FILLER_74_88 ();
 sg13g2_decap_8 FILLER_74_95 ();
 sg13g2_decap_8 FILLER_74_102 ();
 sg13g2_decap_8 FILLER_74_109 ();
 sg13g2_decap_8 FILLER_74_116 ();
 sg13g2_decap_8 FILLER_74_123 ();
 sg13g2_decap_4 FILLER_74_130 ();
 sg13g2_fill_2 FILLER_74_134 ();
 sg13g2_decap_4 FILLER_74_162 ();
 sg13g2_fill_2 FILLER_74_166 ();
 sg13g2_fill_2 FILLER_74_172 ();
 sg13g2_fill_1 FILLER_74_177 ();
 sg13g2_decap_8 FILLER_74_195 ();
 sg13g2_decap_4 FILLER_74_202 ();
 sg13g2_fill_2 FILLER_74_206 ();
 sg13g2_decap_8 FILLER_74_219 ();
 sg13g2_fill_2 FILLER_74_226 ();
 sg13g2_fill_2 FILLER_74_294 ();
 sg13g2_fill_1 FILLER_74_302 ();
 sg13g2_decap_4 FILLER_74_308 ();
 sg13g2_fill_1 FILLER_74_318 ();
 sg13g2_decap_8 FILLER_74_323 ();
 sg13g2_decap_8 FILLER_74_330 ();
 sg13g2_decap_8 FILLER_74_337 ();
 sg13g2_decap_8 FILLER_74_344 ();
 sg13g2_decap_4 FILLER_74_351 ();
 sg13g2_fill_1 FILLER_74_355 ();
 sg13g2_decap_8 FILLER_74_397 ();
 sg13g2_decap_8 FILLER_74_404 ();
 sg13g2_decap_4 FILLER_74_411 ();
 sg13g2_decap_4 FILLER_74_427 ();
 sg13g2_decap_4 FILLER_74_435 ();
 sg13g2_fill_1 FILLER_74_439 ();
 sg13g2_decap_8 FILLER_74_444 ();
 sg13g2_decap_8 FILLER_74_451 ();
 sg13g2_decap_4 FILLER_74_458 ();
 sg13g2_fill_1 FILLER_74_462 ();
 sg13g2_fill_1 FILLER_74_479 ();
 sg13g2_fill_1 FILLER_74_485 ();
 sg13g2_fill_2 FILLER_74_503 ();
 sg13g2_decap_8 FILLER_74_509 ();
 sg13g2_decap_8 FILLER_74_516 ();
 sg13g2_decap_8 FILLER_74_523 ();
 sg13g2_decap_8 FILLER_74_530 ();
 sg13g2_decap_4 FILLER_74_537 ();
 sg13g2_fill_2 FILLER_74_541 ();
 sg13g2_decap_4 FILLER_74_572 ();
 sg13g2_fill_2 FILLER_74_576 ();
 sg13g2_fill_1 FILLER_74_608 ();
 sg13g2_decap_4 FILLER_74_612 ();
 sg13g2_fill_2 FILLER_74_616 ();
 sg13g2_decap_4 FILLER_74_624 ();
 sg13g2_fill_1 FILLER_74_628 ();
 sg13g2_decap_8 FILLER_74_633 ();
 sg13g2_decap_8 FILLER_74_640 ();
 sg13g2_fill_1 FILLER_74_647 ();
 sg13g2_decap_8 FILLER_74_651 ();
 sg13g2_decap_8 FILLER_74_658 ();
 sg13g2_fill_1 FILLER_74_665 ();
 sg13g2_decap_8 FILLER_74_670 ();
 sg13g2_decap_8 FILLER_74_677 ();
 sg13g2_decap_8 FILLER_74_684 ();
 sg13g2_decap_4 FILLER_74_691 ();
 sg13g2_decap_8 FILLER_74_726 ();
 sg13g2_decap_4 FILLER_74_733 ();
 sg13g2_decap_8 FILLER_74_763 ();
 sg13g2_fill_2 FILLER_74_782 ();
 sg13g2_decap_4 FILLER_74_787 ();
 sg13g2_fill_1 FILLER_74_791 ();
 sg13g2_decap_8 FILLER_74_804 ();
 sg13g2_decap_8 FILLER_74_811 ();
 sg13g2_decap_8 FILLER_74_818 ();
 sg13g2_decap_8 FILLER_74_837 ();
 sg13g2_decap_8 FILLER_74_844 ();
 sg13g2_decap_4 FILLER_74_851 ();
 sg13g2_fill_1 FILLER_74_855 ();
 sg13g2_decap_8 FILLER_74_861 ();
 sg13g2_fill_2 FILLER_74_873 ();
 sg13g2_fill_1 FILLER_74_875 ();
 sg13g2_decap_8 FILLER_74_887 ();
 sg13g2_decap_8 FILLER_74_894 ();
 sg13g2_decap_8 FILLER_74_901 ();
 sg13g2_fill_1 FILLER_74_908 ();
 sg13g2_decap_8 FILLER_74_915 ();
 sg13g2_decap_8 FILLER_74_922 ();
 sg13g2_decap_4 FILLER_74_929 ();
 sg13g2_fill_1 FILLER_74_933 ();
 sg13g2_decap_8 FILLER_74_939 ();
 sg13g2_fill_2 FILLER_74_946 ();
 sg13g2_decap_4 FILLER_74_954 ();
 sg13g2_decap_8 FILLER_74_963 ();
 sg13g2_fill_1 FILLER_74_970 ();
 sg13g2_fill_2 FILLER_74_986 ();
 sg13g2_fill_2 FILLER_74_993 ();
 sg13g2_fill_1 FILLER_74_1005 ();
 sg13g2_decap_8 FILLER_74_1011 ();
 sg13g2_decap_8 FILLER_74_1018 ();
 sg13g2_decap_8 FILLER_74_1025 ();
 sg13g2_decap_8 FILLER_74_1032 ();
 sg13g2_decap_4 FILLER_74_1050 ();
 sg13g2_fill_2 FILLER_74_1054 ();
 sg13g2_fill_1 FILLER_74_1060 ();
 sg13g2_fill_2 FILLER_74_1066 ();
 sg13g2_decap_8 FILLER_74_1072 ();
 sg13g2_fill_1 FILLER_74_1079 ();
 sg13g2_decap_8 FILLER_74_1087 ();
 sg13g2_decap_8 FILLER_74_1094 ();
 sg13g2_fill_2 FILLER_74_1101 ();
 sg13g2_fill_1 FILLER_74_1103 ();
 sg13g2_decap_8 FILLER_74_1108 ();
 sg13g2_decap_8 FILLER_74_1115 ();
 sg13g2_decap_8 FILLER_74_1122 ();
 sg13g2_decap_4 FILLER_74_1129 ();
 sg13g2_fill_2 FILLER_74_1146 ();
 sg13g2_decap_8 FILLER_74_1172 ();
 sg13g2_decap_8 FILLER_74_1179 ();
 sg13g2_fill_2 FILLER_74_1186 ();
 sg13g2_fill_1 FILLER_74_1188 ();
 sg13g2_fill_2 FILLER_74_1194 ();
 sg13g2_decap_8 FILLER_74_1200 ();
 sg13g2_decap_8 FILLER_74_1207 ();
 sg13g2_decap_8 FILLER_74_1214 ();
 sg13g2_fill_2 FILLER_74_1221 ();
 sg13g2_fill_1 FILLER_74_1223 ();
 sg13g2_decap_8 FILLER_74_1228 ();
 sg13g2_decap_8 FILLER_74_1235 ();
 sg13g2_decap_8 FILLER_74_1242 ();
 sg13g2_decap_8 FILLER_74_1249 ();
 sg13g2_fill_2 FILLER_74_1269 ();
 sg13g2_decap_8 FILLER_74_1297 ();
 sg13g2_decap_8 FILLER_74_1304 ();
 sg13g2_decap_8 FILLER_74_1311 ();
 sg13g2_decap_4 FILLER_74_1318 ();
 sg13g2_fill_2 FILLER_74_1322 ();
 sg13g2_decap_8 FILLER_74_1332 ();
 sg13g2_decap_4 FILLER_74_1339 ();
 sg13g2_fill_1 FILLER_74_1343 ();
 sg13g2_fill_1 FILLER_74_1348 ();
 sg13g2_decap_8 FILLER_74_1362 ();
 sg13g2_decap_4 FILLER_74_1369 ();
 sg13g2_fill_2 FILLER_74_1373 ();
 sg13g2_decap_8 FILLER_74_1383 ();
 sg13g2_decap_4 FILLER_74_1390 ();
 sg13g2_fill_2 FILLER_74_1394 ();
 sg13g2_fill_2 FILLER_74_1425 ();
 sg13g2_fill_1 FILLER_74_1427 ();
 sg13g2_fill_2 FILLER_74_1434 ();
 sg13g2_decap_8 FILLER_74_1440 ();
 sg13g2_decap_8 FILLER_74_1447 ();
 sg13g2_decap_8 FILLER_74_1454 ();
 sg13g2_decap_8 FILLER_74_1461 ();
 sg13g2_fill_1 FILLER_74_1468 ();
 sg13g2_decap_8 FILLER_74_1478 ();
 sg13g2_decap_8 FILLER_74_1485 ();
 sg13g2_decap_8 FILLER_74_1492 ();
 sg13g2_fill_2 FILLER_74_1499 ();
 sg13g2_fill_1 FILLER_74_1501 ();
 sg13g2_decap_4 FILLER_74_1520 ();
 sg13g2_fill_2 FILLER_74_1529 ();
 sg13g2_decap_8 FILLER_74_1536 ();
 sg13g2_decap_8 FILLER_74_1543 ();
 sg13g2_decap_8 FILLER_74_1592 ();
 sg13g2_decap_4 FILLER_74_1599 ();
 sg13g2_decap_8 FILLER_74_1629 ();
 sg13g2_fill_2 FILLER_74_1636 ();
 sg13g2_fill_1 FILLER_74_1638 ();
 sg13g2_decap_8 FILLER_74_1651 ();
 sg13g2_decap_8 FILLER_74_1662 ();
 sg13g2_fill_2 FILLER_74_1669 ();
 sg13g2_decap_8 FILLER_74_1710 ();
 sg13g2_decap_8 FILLER_74_1717 ();
 sg13g2_fill_2 FILLER_74_1724 ();
 sg13g2_fill_1 FILLER_74_1726 ();
 sg13g2_decap_8 FILLER_74_1757 ();
 sg13g2_decap_8 FILLER_74_1764 ();
 sg13g2_fill_2 FILLER_74_1771 ();
 sg13g2_fill_1 FILLER_74_1773 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_4 FILLER_75_7 ();
 sg13g2_fill_1 FILLER_75_11 ();
 sg13g2_decap_8 FILLER_75_16 ();
 sg13g2_decap_8 FILLER_75_23 ();
 sg13g2_fill_2 FILLER_75_30 ();
 sg13g2_fill_1 FILLER_75_32 ();
 sg13g2_decap_8 FILLER_75_37 ();
 sg13g2_decap_4 FILLER_75_44 ();
 sg13g2_fill_1 FILLER_75_48 ();
 sg13g2_decap_8 FILLER_75_54 ();
 sg13g2_fill_2 FILLER_75_61 ();
 sg13g2_fill_1 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_68 ();
 sg13g2_fill_2 FILLER_75_75 ();
 sg13g2_decap_8 FILLER_75_128 ();
 sg13g2_decap_8 FILLER_75_135 ();
 sg13g2_decap_4 FILLER_75_142 ();
 sg13g2_fill_2 FILLER_75_146 ();
 sg13g2_decap_4 FILLER_75_152 ();
 sg13g2_fill_1 FILLER_75_160 ();
 sg13g2_decap_4 FILLER_75_191 ();
 sg13g2_decap_4 FILLER_75_199 ();
 sg13g2_decap_8 FILLER_75_227 ();
 sg13g2_decap_8 FILLER_75_234 ();
 sg13g2_decap_8 FILLER_75_241 ();
 sg13g2_fill_2 FILLER_75_248 ();
 sg13g2_fill_1 FILLER_75_250 ();
 sg13g2_decap_8 FILLER_75_255 ();
 sg13g2_decap_8 FILLER_75_262 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_4 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_317 ();
 sg13g2_decap_8 FILLER_75_324 ();
 sg13g2_decap_8 FILLER_75_331 ();
 sg13g2_decap_4 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_342 ();
 sg13g2_decap_8 FILLER_75_347 ();
 sg13g2_decap_8 FILLER_75_354 ();
 sg13g2_decap_8 FILLER_75_361 ();
 sg13g2_decap_4 FILLER_75_368 ();
 sg13g2_decap_8 FILLER_75_377 ();
 sg13g2_fill_1 FILLER_75_384 ();
 sg13g2_fill_2 FILLER_75_400 ();
 sg13g2_decap_4 FILLER_75_406 ();
 sg13g2_fill_2 FILLER_75_414 ();
 sg13g2_fill_1 FILLER_75_416 ();
 sg13g2_fill_1 FILLER_75_434 ();
 sg13g2_decap_4 FILLER_75_440 ();
 sg13g2_fill_1 FILLER_75_444 ();
 sg13g2_decap_8 FILLER_75_451 ();
 sg13g2_decap_4 FILLER_75_458 ();
 sg13g2_fill_1 FILLER_75_462 ();
 sg13g2_decap_8 FILLER_75_468 ();
 sg13g2_decap_8 FILLER_75_475 ();
 sg13g2_fill_2 FILLER_75_482 ();
 sg13g2_fill_1 FILLER_75_484 ();
 sg13g2_decap_8 FILLER_75_489 ();
 sg13g2_fill_2 FILLER_75_496 ();
 sg13g2_fill_1 FILLER_75_498 ();
 sg13g2_decap_4 FILLER_75_503 ();
 sg13g2_fill_1 FILLER_75_507 ();
 sg13g2_decap_4 FILLER_75_548 ();
 sg13g2_decap_8 FILLER_75_556 ();
 sg13g2_fill_2 FILLER_75_563 ();
 sg13g2_fill_1 FILLER_75_565 ();
 sg13g2_decap_8 FILLER_75_571 ();
 sg13g2_decap_8 FILLER_75_578 ();
 sg13g2_fill_2 FILLER_75_585 ();
 sg13g2_fill_1 FILLER_75_587 ();
 sg13g2_decap_4 FILLER_75_592 ();
 sg13g2_fill_1 FILLER_75_607 ();
 sg13g2_decap_8 FILLER_75_612 ();
 sg13g2_fill_2 FILLER_75_619 ();
 sg13g2_fill_1 FILLER_75_621 ();
 sg13g2_fill_2 FILLER_75_626 ();
 sg13g2_decap_8 FILLER_75_641 ();
 sg13g2_decap_4 FILLER_75_653 ();
 sg13g2_fill_2 FILLER_75_657 ();
 sg13g2_decap_4 FILLER_75_663 ();
 sg13g2_fill_1 FILLER_75_667 ();
 sg13g2_decap_8 FILLER_75_687 ();
 sg13g2_decap_8 FILLER_75_694 ();
 sg13g2_decap_4 FILLER_75_701 ();
 sg13g2_fill_2 FILLER_75_705 ();
 sg13g2_decap_4 FILLER_75_711 ();
 sg13g2_fill_1 FILLER_75_715 ();
 sg13g2_decap_8 FILLER_75_719 ();
 sg13g2_decap_8 FILLER_75_726 ();
 sg13g2_decap_8 FILLER_75_733 ();
 sg13g2_decap_4 FILLER_75_740 ();
 sg13g2_decap_8 FILLER_75_748 ();
 sg13g2_decap_8 FILLER_75_755 ();
 sg13g2_decap_8 FILLER_75_762 ();
 sg13g2_decap_8 FILLER_75_769 ();
 sg13g2_fill_1 FILLER_75_776 ();
 sg13g2_fill_2 FILLER_75_780 ();
 sg13g2_fill_1 FILLER_75_782 ();
 sg13g2_decap_8 FILLER_75_792 ();
 sg13g2_fill_2 FILLER_75_799 ();
 sg13g2_fill_1 FILLER_75_801 ();
 sg13g2_decap_8 FILLER_75_812 ();
 sg13g2_fill_2 FILLER_75_819 ();
 sg13g2_fill_1 FILLER_75_821 ();
 sg13g2_fill_2 FILLER_75_826 ();
 sg13g2_fill_1 FILLER_75_828 ();
 sg13g2_decap_8 FILLER_75_837 ();
 sg13g2_decap_8 FILLER_75_844 ();
 sg13g2_fill_2 FILLER_75_851 ();
 sg13g2_decap_4 FILLER_75_861 ();
 sg13g2_fill_2 FILLER_75_865 ();
 sg13g2_decap_8 FILLER_75_872 ();
 sg13g2_decap_8 FILLER_75_879 ();
 sg13g2_decap_8 FILLER_75_886 ();
 sg13g2_decap_8 FILLER_75_893 ();
 sg13g2_decap_8 FILLER_75_900 ();
 sg13g2_fill_1 FILLER_75_907 ();
 sg13g2_decap_8 FILLER_75_924 ();
 sg13g2_fill_2 FILLER_75_931 ();
 sg13g2_fill_1 FILLER_75_933 ();
 sg13g2_decap_8 FILLER_75_938 ();
 sg13g2_fill_2 FILLER_75_945 ();
 sg13g2_decap_8 FILLER_75_952 ();
 sg13g2_decap_8 FILLER_75_959 ();
 sg13g2_decap_4 FILLER_75_966 ();
 sg13g2_fill_2 FILLER_75_970 ();
 sg13g2_decap_4 FILLER_75_977 ();
 sg13g2_fill_1 FILLER_75_981 ();
 sg13g2_fill_1 FILLER_75_995 ();
 sg13g2_decap_8 FILLER_75_999 ();
 sg13g2_decap_8 FILLER_75_1006 ();
 sg13g2_decap_8 FILLER_75_1013 ();
 sg13g2_decap_4 FILLER_75_1020 ();
 sg13g2_fill_1 FILLER_75_1024 ();
 sg13g2_decap_8 FILLER_75_1051 ();
 sg13g2_fill_2 FILLER_75_1058 ();
 sg13g2_fill_1 FILLER_75_1060 ();
 sg13g2_decap_8 FILLER_75_1065 ();
 sg13g2_decap_8 FILLER_75_1072 ();
 sg13g2_decap_8 FILLER_75_1079 ();
 sg13g2_decap_8 FILLER_75_1086 ();
 sg13g2_fill_2 FILLER_75_1093 ();
 sg13g2_fill_1 FILLER_75_1095 ();
 sg13g2_decap_4 FILLER_75_1106 ();
 sg13g2_fill_1 FILLER_75_1110 ();
 sg13g2_decap_8 FILLER_75_1124 ();
 sg13g2_decap_8 FILLER_75_1131 ();
 sg13g2_fill_1 FILLER_75_1138 ();
 sg13g2_fill_2 FILLER_75_1152 ();
 sg13g2_fill_2 FILLER_75_1175 ();
 sg13g2_decap_4 FILLER_75_1181 ();
 sg13g2_fill_1 FILLER_75_1193 ();
 sg13g2_fill_2 FILLER_75_1199 ();
 sg13g2_fill_2 FILLER_75_1209 ();
 sg13g2_fill_1 FILLER_75_1215 ();
 sg13g2_decap_8 FILLER_75_1220 ();
 sg13g2_decap_8 FILLER_75_1227 ();
 sg13g2_decap_8 FILLER_75_1234 ();
 sg13g2_decap_8 FILLER_75_1241 ();
 sg13g2_decap_8 FILLER_75_1252 ();
 sg13g2_decap_8 FILLER_75_1259 ();
 sg13g2_decap_8 FILLER_75_1283 ();
 sg13g2_decap_8 FILLER_75_1290 ();
 sg13g2_decap_8 FILLER_75_1297 ();
 sg13g2_decap_8 FILLER_75_1304 ();
 sg13g2_decap_8 FILLER_75_1311 ();
 sg13g2_fill_2 FILLER_75_1318 ();
 sg13g2_fill_1 FILLER_75_1320 ();
 sg13g2_decap_8 FILLER_75_1325 ();
 sg13g2_decap_4 FILLER_75_1332 ();
 sg13g2_decap_8 FILLER_75_1341 ();
 sg13g2_decap_8 FILLER_75_1352 ();
 sg13g2_decap_4 FILLER_75_1359 ();
 sg13g2_fill_1 FILLER_75_1363 ();
 sg13g2_decap_8 FILLER_75_1395 ();
 sg13g2_decap_8 FILLER_75_1402 ();
 sg13g2_decap_8 FILLER_75_1409 ();
 sg13g2_decap_4 FILLER_75_1416 ();
 sg13g2_fill_1 FILLER_75_1432 ();
 sg13g2_decap_8 FILLER_75_1439 ();
 sg13g2_decap_8 FILLER_75_1446 ();
 sg13g2_decap_8 FILLER_75_1453 ();
 sg13g2_decap_8 FILLER_75_1460 ();
 sg13g2_decap_4 FILLER_75_1467 ();
 sg13g2_fill_1 FILLER_75_1471 ();
 sg13g2_fill_1 FILLER_75_1477 ();
 sg13g2_decap_8 FILLER_75_1481 ();
 sg13g2_decap_8 FILLER_75_1488 ();
 sg13g2_decap_4 FILLER_75_1495 ();
 sg13g2_fill_1 FILLER_75_1499 ();
 sg13g2_fill_2 FILLER_75_1507 ();
 sg13g2_fill_1 FILLER_75_1513 ();
 sg13g2_fill_2 FILLER_75_1520 ();
 sg13g2_fill_2 FILLER_75_1525 ();
 sg13g2_fill_2 FILLER_75_1532 ();
 sg13g2_fill_1 FILLER_75_1534 ();
 sg13g2_decap_4 FILLER_75_1540 ();
 sg13g2_fill_2 FILLER_75_1544 ();
 sg13g2_decap_8 FILLER_75_1553 ();
 sg13g2_decap_4 FILLER_75_1560 ();
 sg13g2_decap_8 FILLER_75_1568 ();
 sg13g2_decap_4 FILLER_75_1575 ();
 sg13g2_fill_2 FILLER_75_1579 ();
 sg13g2_decap_8 FILLER_75_1599 ();
 sg13g2_decap_8 FILLER_75_1611 ();
 sg13g2_decap_8 FILLER_75_1618 ();
 sg13g2_fill_2 FILLER_75_1625 ();
 sg13g2_fill_1 FILLER_75_1627 ();
 sg13g2_fill_2 FILLER_75_1633 ();
 sg13g2_fill_1 FILLER_75_1635 ();
 sg13g2_decap_8 FILLER_75_1640 ();
 sg13g2_fill_1 FILLER_75_1647 ();
 sg13g2_decap_8 FILLER_75_1669 ();
 sg13g2_decap_8 FILLER_75_1680 ();
 sg13g2_decap_8 FILLER_75_1687 ();
 sg13g2_decap_8 FILLER_75_1694 ();
 sg13g2_decap_8 FILLER_75_1701 ();
 sg13g2_decap_8 FILLER_75_1708 ();
 sg13g2_decap_8 FILLER_75_1715 ();
 sg13g2_decap_8 FILLER_75_1722 ();
 sg13g2_decap_8 FILLER_75_1729 ();
 sg13g2_decap_8 FILLER_75_1736 ();
 sg13g2_decap_8 FILLER_75_1743 ();
 sg13g2_decap_8 FILLER_75_1750 ();
 sg13g2_decap_8 FILLER_75_1757 ();
 sg13g2_decap_8 FILLER_75_1764 ();
 sg13g2_fill_2 FILLER_75_1771 ();
 sg13g2_fill_1 FILLER_75_1773 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_4 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_11 ();
 sg13g2_decap_8 FILLER_76_16 ();
 sg13g2_decap_8 FILLER_76_23 ();
 sg13g2_decap_8 FILLER_76_30 ();
 sg13g2_fill_2 FILLER_76_37 ();
 sg13g2_fill_1 FILLER_76_39 ();
 sg13g2_decap_8 FILLER_76_66 ();
 sg13g2_decap_8 FILLER_76_73 ();
 sg13g2_fill_2 FILLER_76_80 ();
 sg13g2_decap_8 FILLER_76_87 ();
 sg13g2_decap_8 FILLER_76_94 ();
 sg13g2_decap_8 FILLER_76_101 ();
 sg13g2_fill_1 FILLER_76_108 ();
 sg13g2_decap_8 FILLER_76_113 ();
 sg13g2_decap_8 FILLER_76_120 ();
 sg13g2_decap_8 FILLER_76_127 ();
 sg13g2_fill_2 FILLER_76_149 ();
 sg13g2_decap_8 FILLER_76_155 ();
 sg13g2_decap_4 FILLER_76_162 ();
 sg13g2_decap_8 FILLER_76_170 ();
 sg13g2_decap_8 FILLER_76_177 ();
 sg13g2_decap_8 FILLER_76_184 ();
 sg13g2_decap_8 FILLER_76_191 ();
 sg13g2_decap_4 FILLER_76_198 ();
 sg13g2_fill_1 FILLER_76_202 ();
 sg13g2_fill_2 FILLER_76_224 ();
 sg13g2_fill_1 FILLER_76_226 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_fill_1 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_257 ();
 sg13g2_decap_8 FILLER_76_264 ();
 sg13g2_decap_8 FILLER_76_271 ();
 sg13g2_decap_8 FILLER_76_278 ();
 sg13g2_decap_8 FILLER_76_285 ();
 sg13g2_fill_2 FILLER_76_292 ();
 sg13g2_fill_1 FILLER_76_294 ();
 sg13g2_fill_1 FILLER_76_305 ();
 sg13g2_decap_8 FILLER_76_319 ();
 sg13g2_decap_4 FILLER_76_326 ();
 sg13g2_fill_2 FILLER_76_330 ();
 sg13g2_fill_1 FILLER_76_336 ();
 sg13g2_fill_1 FILLER_76_363 ();
 sg13g2_fill_1 FILLER_76_367 ();
 sg13g2_fill_2 FILLER_76_375 ();
 sg13g2_decap_8 FILLER_76_383 ();
 sg13g2_decap_4 FILLER_76_390 ();
 sg13g2_fill_2 FILLER_76_394 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_413 ();
 sg13g2_decap_8 FILLER_76_420 ();
 sg13g2_decap_8 FILLER_76_427 ();
 sg13g2_decap_8 FILLER_76_434 ();
 sg13g2_fill_2 FILLER_76_449 ();
 sg13g2_fill_2 FILLER_76_455 ();
 sg13g2_fill_1 FILLER_76_487 ();
 sg13g2_fill_2 FILLER_76_498 ();
 sg13g2_decap_8 FILLER_76_505 ();
 sg13g2_decap_8 FILLER_76_512 ();
 sg13g2_decap_8 FILLER_76_519 ();
 sg13g2_decap_4 FILLER_76_526 ();
 sg13g2_decap_8 FILLER_76_534 ();
 sg13g2_decap_8 FILLER_76_541 ();
 sg13g2_decap_8 FILLER_76_548 ();
 sg13g2_decap_8 FILLER_76_555 ();
 sg13g2_fill_2 FILLER_76_562 ();
 sg13g2_fill_1 FILLER_76_564 ();
 sg13g2_decap_8 FILLER_76_569 ();
 sg13g2_decap_8 FILLER_76_576 ();
 sg13g2_decap_8 FILLER_76_583 ();
 sg13g2_decap_8 FILLER_76_590 ();
 sg13g2_decap_4 FILLER_76_597 ();
 sg13g2_fill_1 FILLER_76_601 ();
 sg13g2_decap_8 FILLER_76_632 ();
 sg13g2_decap_8 FILLER_76_639 ();
 sg13g2_fill_2 FILLER_76_646 ();
 sg13g2_fill_1 FILLER_76_648 ();
 sg13g2_fill_1 FILLER_76_678 ();
 sg13g2_fill_2 FILLER_76_695 ();
 sg13g2_decap_8 FILLER_76_706 ();
 sg13g2_decap_8 FILLER_76_742 ();
 sg13g2_decap_8 FILLER_76_749 ();
 sg13g2_decap_4 FILLER_76_756 ();
 sg13g2_fill_1 FILLER_76_760 ();
 sg13g2_decap_4 FILLER_76_764 ();
 sg13g2_decap_8 FILLER_76_793 ();
 sg13g2_decap_4 FILLER_76_800 ();
 sg13g2_fill_2 FILLER_76_804 ();
 sg13g2_fill_1 FILLER_76_811 ();
 sg13g2_decap_4 FILLER_76_828 ();
 sg13g2_fill_1 FILLER_76_832 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_fill_2 FILLER_76_856 ();
 sg13g2_decap_4 FILLER_76_866 ();
 sg13g2_fill_2 FILLER_76_870 ();
 sg13g2_fill_1 FILLER_76_878 ();
 sg13g2_fill_1 FILLER_76_890 ();
 sg13g2_decap_4 FILLER_76_896 ();
 sg13g2_fill_2 FILLER_76_900 ();
 sg13g2_decap_4 FILLER_76_932 ();
 sg13g2_fill_1 FILLER_76_936 ();
 sg13g2_fill_2 FILLER_76_941 ();
 sg13g2_fill_1 FILLER_76_943 ();
 sg13g2_fill_1 FILLER_76_957 ();
 sg13g2_fill_1 FILLER_76_967 ();
 sg13g2_decap_4 FILLER_76_973 ();
 sg13g2_fill_2 FILLER_76_977 ();
 sg13g2_fill_2 FILLER_76_999 ();
 sg13g2_fill_1 FILLER_76_1001 ();
 sg13g2_decap_8 FILLER_76_1012 ();
 sg13g2_decap_8 FILLER_76_1019 ();
 sg13g2_decap_8 FILLER_76_1026 ();
 sg13g2_fill_1 FILLER_76_1033 ();
 sg13g2_decap_4 FILLER_76_1043 ();
 sg13g2_fill_2 FILLER_76_1047 ();
 sg13g2_decap_4 FILLER_76_1089 ();
 sg13g2_fill_1 FILLER_76_1093 ();
 sg13g2_decap_8 FILLER_76_1103 ();
 sg13g2_decap_4 FILLER_76_1110 ();
 sg13g2_fill_1 FILLER_76_1114 ();
 sg13g2_decap_8 FILLER_76_1120 ();
 sg13g2_decap_8 FILLER_76_1127 ();
 sg13g2_decap_8 FILLER_76_1134 ();
 sg13g2_decap_4 FILLER_76_1141 ();
 sg13g2_fill_2 FILLER_76_1161 ();
 sg13g2_fill_1 FILLER_76_1173 ();
 sg13g2_decap_8 FILLER_76_1178 ();
 sg13g2_decap_8 FILLER_76_1185 ();
 sg13g2_decap_4 FILLER_76_1192 ();
 sg13g2_fill_2 FILLER_76_1207 ();
 sg13g2_fill_1 FILLER_76_1209 ();
 sg13g2_decap_4 FILLER_76_1215 ();
 sg13g2_fill_2 FILLER_76_1219 ();
 sg13g2_fill_1 FILLER_76_1240 ();
 sg13g2_fill_2 FILLER_76_1271 ();
 sg13g2_fill_1 FILLER_76_1273 ();
 sg13g2_decap_8 FILLER_76_1305 ();
 sg13g2_fill_2 FILLER_76_1312 ();
 sg13g2_fill_1 FILLER_76_1314 ();
 sg13g2_fill_1 FILLER_76_1341 ();
 sg13g2_decap_8 FILLER_76_1351 ();
 sg13g2_decap_8 FILLER_76_1358 ();
 sg13g2_decap_8 FILLER_76_1365 ();
 sg13g2_decap_8 FILLER_76_1372 ();
 sg13g2_decap_8 FILLER_76_1388 ();
 sg13g2_decap_8 FILLER_76_1395 ();
 sg13g2_fill_2 FILLER_76_1402 ();
 sg13g2_fill_1 FILLER_76_1404 ();
 sg13g2_fill_1 FILLER_76_1436 ();
 sg13g2_decap_8 FILLER_76_1446 ();
 sg13g2_decap_8 FILLER_76_1453 ();
 sg13g2_decap_4 FILLER_76_1464 ();
 sg13g2_fill_1 FILLER_76_1468 ();
 sg13g2_decap_8 FILLER_76_1495 ();
 sg13g2_fill_2 FILLER_76_1502 ();
 sg13g2_fill_2 FILLER_76_1535 ();
 sg13g2_fill_1 FILLER_76_1537 ();
 sg13g2_decap_8 FILLER_76_1545 ();
 sg13g2_fill_1 FILLER_76_1552 ();
 sg13g2_decap_8 FILLER_76_1613 ();
 sg13g2_decap_8 FILLER_76_1620 ();
 sg13g2_fill_2 FILLER_76_1627 ();
 sg13g2_decap_8 FILLER_76_1655 ();
 sg13g2_decap_8 FILLER_76_1662 ();
 sg13g2_decap_8 FILLER_76_1669 ();
 sg13g2_decap_8 FILLER_76_1676 ();
 sg13g2_decap_8 FILLER_76_1683 ();
 sg13g2_decap_8 FILLER_76_1690 ();
 sg13g2_decap_8 FILLER_76_1697 ();
 sg13g2_decap_8 FILLER_76_1704 ();
 sg13g2_decap_8 FILLER_76_1711 ();
 sg13g2_decap_8 FILLER_76_1718 ();
 sg13g2_decap_8 FILLER_76_1725 ();
 sg13g2_decap_8 FILLER_76_1732 ();
 sg13g2_decap_8 FILLER_76_1739 ();
 sg13g2_decap_8 FILLER_76_1746 ();
 sg13g2_decap_8 FILLER_76_1753 ();
 sg13g2_decap_8 FILLER_76_1760 ();
 sg13g2_decap_8 FILLER_76_1767 ();
 sg13g2_decap_4 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_4 ();
 sg13g2_decap_4 FILLER_77_35 ();
 sg13g2_fill_1 FILLER_77_39 ();
 sg13g2_decap_4 FILLER_77_44 ();
 sg13g2_fill_2 FILLER_77_48 ();
 sg13g2_decap_8 FILLER_77_54 ();
 sg13g2_decap_8 FILLER_77_61 ();
 sg13g2_decap_8 FILLER_77_68 ();
 sg13g2_decap_4 FILLER_77_75 ();
 sg13g2_fill_2 FILLER_77_79 ();
 sg13g2_decap_8 FILLER_77_88 ();
 sg13g2_decap_8 FILLER_77_95 ();
 sg13g2_decap_8 FILLER_77_102 ();
 sg13g2_decap_8 FILLER_77_109 ();
 sg13g2_decap_4 FILLER_77_116 ();
 sg13g2_fill_2 FILLER_77_120 ();
 sg13g2_decap_8 FILLER_77_170 ();
 sg13g2_decap_8 FILLER_77_177 ();
 sg13g2_decap_8 FILLER_77_184 ();
 sg13g2_decap_8 FILLER_77_246 ();
 sg13g2_fill_1 FILLER_77_253 ();
 sg13g2_decap_4 FILLER_77_284 ();
 sg13g2_fill_2 FILLER_77_312 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_4 FILLER_77_336 ();
 sg13g2_fill_2 FILLER_77_340 ();
 sg13g2_decap_4 FILLER_77_355 ();
 sg13g2_decap_4 FILLER_77_368 ();
 sg13g2_fill_1 FILLER_77_376 ();
 sg13g2_fill_1 FILLER_77_383 ();
 sg13g2_fill_1 FILLER_77_389 ();
 sg13g2_fill_2 FILLER_77_408 ();
 sg13g2_fill_2 FILLER_77_416 ();
 sg13g2_fill_1 FILLER_77_418 ();
 sg13g2_decap_8 FILLER_77_424 ();
 sg13g2_decap_8 FILLER_77_431 ();
 sg13g2_decap_8 FILLER_77_438 ();
 sg13g2_decap_8 FILLER_77_445 ();
 sg13g2_decap_8 FILLER_77_452 ();
 sg13g2_decap_8 FILLER_77_469 ();
 sg13g2_decap_8 FILLER_77_485 ();
 sg13g2_decap_4 FILLER_77_492 ();
 sg13g2_decap_4 FILLER_77_501 ();
 sg13g2_decap_8 FILLER_77_509 ();
 sg13g2_decap_4 FILLER_77_516 ();
 sg13g2_decap_4 FILLER_77_524 ();
 sg13g2_decap_4 FILLER_77_532 ();
 sg13g2_fill_1 FILLER_77_536 ();
 sg13g2_fill_2 FILLER_77_545 ();
 sg13g2_fill_1 FILLER_77_547 ();
 sg13g2_fill_1 FILLER_77_552 ();
 sg13g2_decap_8 FILLER_77_584 ();
 sg13g2_decap_8 FILLER_77_591 ();
 sg13g2_decap_8 FILLER_77_598 ();
 sg13g2_decap_8 FILLER_77_605 ();
 sg13g2_decap_8 FILLER_77_612 ();
 sg13g2_fill_2 FILLER_77_619 ();
 sg13g2_fill_1 FILLER_77_621 ();
 sg13g2_decap_8 FILLER_77_645 ();
 sg13g2_decap_4 FILLER_77_652 ();
 sg13g2_decap_8 FILLER_77_660 ();
 sg13g2_decap_4 FILLER_77_667 ();
 sg13g2_fill_1 FILLER_77_671 ();
 sg13g2_fill_2 FILLER_77_690 ();
 sg13g2_fill_2 FILLER_77_700 ();
 sg13g2_decap_8 FILLER_77_714 ();
 sg13g2_fill_1 FILLER_77_721 ();
 sg13g2_decap_8 FILLER_77_726 ();
 sg13g2_decap_8 FILLER_77_733 ();
 sg13g2_decap_8 FILLER_77_740 ();
 sg13g2_fill_1 FILLER_77_747 ();
 sg13g2_decap_8 FILLER_77_752 ();
 sg13g2_decap_4 FILLER_77_759 ();
 sg13g2_fill_2 FILLER_77_763 ();
 sg13g2_decap_4 FILLER_77_778 ();
 sg13g2_fill_2 FILLER_77_787 ();
 sg13g2_fill_1 FILLER_77_792 ();
 sg13g2_fill_1 FILLER_77_801 ();
 sg13g2_decap_8 FILLER_77_817 ();
 sg13g2_decap_8 FILLER_77_824 ();
 sg13g2_decap_8 FILLER_77_846 ();
 sg13g2_fill_2 FILLER_77_853 ();
 sg13g2_fill_1 FILLER_77_860 ();
 sg13g2_fill_1 FILLER_77_866 ();
 sg13g2_fill_1 FILLER_77_879 ();
 sg13g2_fill_1 FILLER_77_885 ();
 sg13g2_fill_2 FILLER_77_894 ();
 sg13g2_fill_1 FILLER_77_896 ();
 sg13g2_fill_1 FILLER_77_902 ();
 sg13g2_decap_8 FILLER_77_917 ();
 sg13g2_decap_8 FILLER_77_924 ();
 sg13g2_decap_8 FILLER_77_931 ();
 sg13g2_decap_4 FILLER_77_938 ();
 sg13g2_fill_2 FILLER_77_957 ();
 sg13g2_fill_1 FILLER_77_959 ();
 sg13g2_fill_2 FILLER_77_965 ();
 sg13g2_decap_4 FILLER_77_971 ();
 sg13g2_decap_8 FILLER_77_992 ();
 sg13g2_decap_8 FILLER_77_999 ();
 sg13g2_decap_8 FILLER_77_1006 ();
 sg13g2_decap_8 FILLER_77_1013 ();
 sg13g2_decap_8 FILLER_77_1020 ();
 sg13g2_decap_8 FILLER_77_1027 ();
 sg13g2_fill_1 FILLER_77_1034 ();
 sg13g2_decap_8 FILLER_77_1048 ();
 sg13g2_decap_8 FILLER_77_1055 ();
 sg13g2_decap_8 FILLER_77_1062 ();
 sg13g2_decap_8 FILLER_77_1069 ();
 sg13g2_decap_8 FILLER_77_1076 ();
 sg13g2_decap_8 FILLER_77_1083 ();
 sg13g2_fill_1 FILLER_77_1090 ();
 sg13g2_decap_4 FILLER_77_1107 ();
 sg13g2_decap_8 FILLER_77_1119 ();
 sg13g2_decap_8 FILLER_77_1126 ();
 sg13g2_decap_8 FILLER_77_1133 ();
 sg13g2_fill_2 FILLER_77_1140 ();
 sg13g2_fill_1 FILLER_77_1142 ();
 sg13g2_decap_4 FILLER_77_1156 ();
 sg13g2_fill_1 FILLER_77_1160 ();
 sg13g2_decap_8 FILLER_77_1205 ();
 sg13g2_decap_4 FILLER_77_1217 ();
 sg13g2_fill_2 FILLER_77_1221 ();
 sg13g2_fill_1 FILLER_77_1241 ();
 sg13g2_decap_8 FILLER_77_1246 ();
 sg13g2_decap_8 FILLER_77_1253 ();
 sg13g2_decap_8 FILLER_77_1260 ();
 sg13g2_decap_8 FILLER_77_1267 ();
 sg13g2_decap_4 FILLER_77_1274 ();
 sg13g2_fill_2 FILLER_77_1278 ();
 sg13g2_decap_8 FILLER_77_1284 ();
 sg13g2_decap_8 FILLER_77_1291 ();
 sg13g2_decap_8 FILLER_77_1298 ();
 sg13g2_decap_8 FILLER_77_1305 ();
 sg13g2_decap_8 FILLER_77_1312 ();
 sg13g2_decap_8 FILLER_77_1319 ();
 sg13g2_fill_1 FILLER_77_1326 ();
 sg13g2_decap_8 FILLER_77_1331 ();
 sg13g2_decap_4 FILLER_77_1338 ();
 sg13g2_fill_1 FILLER_77_1342 ();
 sg13g2_decap_4 FILLER_77_1347 ();
 sg13g2_fill_2 FILLER_77_1351 ();
 sg13g2_decap_8 FILLER_77_1361 ();
 sg13g2_decap_8 FILLER_77_1368 ();
 sg13g2_decap_4 FILLER_77_1375 ();
 sg13g2_decap_8 FILLER_77_1385 ();
 sg13g2_decap_8 FILLER_77_1392 ();
 sg13g2_decap_8 FILLER_77_1399 ();
 sg13g2_decap_8 FILLER_77_1406 ();
 sg13g2_decap_4 FILLER_77_1413 ();
 sg13g2_fill_2 FILLER_77_1417 ();
 sg13g2_fill_2 FILLER_77_1442 ();
 sg13g2_fill_1 FILLER_77_1444 ();
 sg13g2_fill_1 FILLER_77_1449 ();
 sg13g2_decap_8 FILLER_77_1455 ();
 sg13g2_decap_8 FILLER_77_1462 ();
 sg13g2_decap_8 FILLER_77_1469 ();
 sg13g2_decap_8 FILLER_77_1480 ();
 sg13g2_decap_8 FILLER_77_1487 ();
 sg13g2_decap_8 FILLER_77_1494 ();
 sg13g2_decap_8 FILLER_77_1501 ();
 sg13g2_decap_8 FILLER_77_1508 ();
 sg13g2_decap_4 FILLER_77_1515 ();
 sg13g2_fill_2 FILLER_77_1519 ();
 sg13g2_decap_8 FILLER_77_1551 ();
 sg13g2_fill_2 FILLER_77_1558 ();
 sg13g2_fill_1 FILLER_77_1560 ();
 sg13g2_decap_8 FILLER_77_1565 ();
 sg13g2_decap_8 FILLER_77_1572 ();
 sg13g2_decap_8 FILLER_77_1579 ();
 sg13g2_decap_4 FILLER_77_1586 ();
 sg13g2_fill_2 FILLER_77_1590 ();
 sg13g2_decap_8 FILLER_77_1596 ();
 sg13g2_decap_8 FILLER_77_1603 ();
 sg13g2_decap_8 FILLER_77_1610 ();
 sg13g2_decap_8 FILLER_77_1617 ();
 sg13g2_decap_8 FILLER_77_1624 ();
 sg13g2_decap_8 FILLER_77_1631 ();
 sg13g2_decap_8 FILLER_77_1638 ();
 sg13g2_decap_8 FILLER_77_1645 ();
 sg13g2_decap_8 FILLER_77_1652 ();
 sg13g2_decap_8 FILLER_77_1659 ();
 sg13g2_decap_8 FILLER_77_1666 ();
 sg13g2_decap_8 FILLER_77_1673 ();
 sg13g2_decap_8 FILLER_77_1680 ();
 sg13g2_decap_8 FILLER_77_1687 ();
 sg13g2_decap_8 FILLER_77_1694 ();
 sg13g2_decap_8 FILLER_77_1701 ();
 sg13g2_decap_8 FILLER_77_1708 ();
 sg13g2_decap_8 FILLER_77_1715 ();
 sg13g2_decap_8 FILLER_77_1722 ();
 sg13g2_decap_8 FILLER_77_1729 ();
 sg13g2_decap_8 FILLER_77_1736 ();
 sg13g2_decap_8 FILLER_77_1743 ();
 sg13g2_decap_8 FILLER_77_1750 ();
 sg13g2_decap_8 FILLER_77_1757 ();
 sg13g2_decap_8 FILLER_77_1764 ();
 sg13g2_fill_2 FILLER_77_1771 ();
 sg13g2_fill_1 FILLER_77_1773 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_4 FILLER_78_7 ();
 sg13g2_fill_2 FILLER_78_11 ();
 sg13g2_decap_8 FILLER_78_17 ();
 sg13g2_decap_8 FILLER_78_24 ();
 sg13g2_decap_8 FILLER_78_31 ();
 sg13g2_fill_2 FILLER_78_38 ();
 sg13g2_decap_8 FILLER_78_53 ();
 sg13g2_fill_1 FILLER_78_60 ();
 sg13g2_decap_4 FILLER_78_65 ();
 sg13g2_decap_4 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_81 ();
 sg13g2_decap_8 FILLER_78_134 ();
 sg13g2_fill_1 FILLER_78_141 ();
 sg13g2_decap_8 FILLER_78_146 ();
 sg13g2_decap_8 FILLER_78_153 ();
 sg13g2_decap_8 FILLER_78_160 ();
 sg13g2_fill_1 FILLER_78_167 ();
 sg13g2_decap_8 FILLER_78_173 ();
 sg13g2_decap_4 FILLER_78_180 ();
 sg13g2_fill_2 FILLER_78_184 ();
 sg13g2_fill_1 FILLER_78_199 ();
 sg13g2_decap_8 FILLER_78_208 ();
 sg13g2_decap_8 FILLER_78_215 ();
 sg13g2_decap_8 FILLER_78_222 ();
 sg13g2_decap_8 FILLER_78_229 ();
 sg13g2_decap_8 FILLER_78_236 ();
 sg13g2_decap_8 FILLER_78_243 ();
 sg13g2_decap_8 FILLER_78_250 ();
 sg13g2_fill_2 FILLER_78_257 ();
 sg13g2_decap_4 FILLER_78_263 ();
 sg13g2_fill_2 FILLER_78_267 ();
 sg13g2_fill_1 FILLER_78_295 ();
 sg13g2_decap_4 FILLER_78_346 ();
 sg13g2_fill_1 FILLER_78_350 ();
 sg13g2_fill_1 FILLER_78_356 ();
 sg13g2_decap_8 FILLER_78_369 ();
 sg13g2_fill_1 FILLER_78_376 ();
 sg13g2_decap_8 FILLER_78_386 ();
 sg13g2_decap_8 FILLER_78_393 ();
 sg13g2_decap_8 FILLER_78_400 ();
 sg13g2_decap_8 FILLER_78_407 ();
 sg13g2_fill_2 FILLER_78_414 ();
 sg13g2_fill_1 FILLER_78_416 ();
 sg13g2_decap_4 FILLER_78_429 ();
 sg13g2_decap_4 FILLER_78_437 ();
 sg13g2_decap_4 FILLER_78_449 ();
 sg13g2_fill_1 FILLER_78_453 ();
 sg13g2_decap_8 FILLER_78_459 ();
 sg13g2_decap_8 FILLER_78_466 ();
 sg13g2_decap_4 FILLER_78_473 ();
 sg13g2_fill_2 FILLER_78_477 ();
 sg13g2_decap_8 FILLER_78_487 ();
 sg13g2_decap_8 FILLER_78_494 ();
 sg13g2_fill_1 FILLER_78_501 ();
 sg13g2_decap_8 FILLER_78_506 ();
 sg13g2_decap_4 FILLER_78_513 ();
 sg13g2_fill_2 FILLER_78_517 ();
 sg13g2_decap_4 FILLER_78_527 ();
 sg13g2_decap_8 FILLER_78_557 ();
 sg13g2_decap_8 FILLER_78_564 ();
 sg13g2_decap_8 FILLER_78_571 ();
 sg13g2_decap_8 FILLER_78_578 ();
 sg13g2_decap_8 FILLER_78_585 ();
 sg13g2_decap_8 FILLER_78_592 ();
 sg13g2_decap_4 FILLER_78_599 ();
 sg13g2_fill_1 FILLER_78_603 ();
 sg13g2_decap_8 FILLER_78_647 ();
 sg13g2_decap_8 FILLER_78_654 ();
 sg13g2_fill_2 FILLER_78_661 ();
 sg13g2_fill_1 FILLER_78_663 ();
 sg13g2_decap_4 FILLER_78_706 ();
 sg13g2_decap_8 FILLER_78_722 ();
 sg13g2_decap_8 FILLER_78_734 ();
 sg13g2_decap_8 FILLER_78_741 ();
 sg13g2_decap_8 FILLER_78_748 ();
 sg13g2_decap_8 FILLER_78_755 ();
 sg13g2_decap_4 FILLER_78_762 ();
 sg13g2_fill_1 FILLER_78_766 ();
 sg13g2_fill_2 FILLER_78_793 ();
 sg13g2_fill_1 FILLER_78_799 ();
 sg13g2_decap_8 FILLER_78_860 ();
 sg13g2_decap_4 FILLER_78_867 ();
 sg13g2_fill_1 FILLER_78_871 ();
 sg13g2_decap_8 FILLER_78_877 ();
 sg13g2_decap_8 FILLER_78_884 ();
 sg13g2_decap_8 FILLER_78_891 ();
 sg13g2_decap_4 FILLER_78_898 ();
 sg13g2_decap_4 FILLER_78_906 ();
 sg13g2_fill_2 FILLER_78_910 ();
 sg13g2_decap_8 FILLER_78_916 ();
 sg13g2_decap_8 FILLER_78_923 ();
 sg13g2_decap_4 FILLER_78_930 ();
 sg13g2_decap_4 FILLER_78_938 ();
 sg13g2_fill_1 FILLER_78_942 ();
 sg13g2_decap_8 FILLER_78_955 ();
 sg13g2_decap_8 FILLER_78_962 ();
 sg13g2_decap_8 FILLER_78_969 ();
 sg13g2_decap_8 FILLER_78_976 ();
 sg13g2_decap_8 FILLER_78_983 ();
 sg13g2_decap_8 FILLER_78_990 ();
 sg13g2_decap_8 FILLER_78_997 ();
 sg13g2_fill_2 FILLER_78_1004 ();
 sg13g2_fill_1 FILLER_78_1006 ();
 sg13g2_decap_4 FILLER_78_1029 ();
 sg13g2_fill_1 FILLER_78_1033 ();
 sg13g2_decap_8 FILLER_78_1052 ();
 sg13g2_decap_8 FILLER_78_1059 ();
 sg13g2_decap_4 FILLER_78_1066 ();
 sg13g2_decap_4 FILLER_78_1076 ();
 sg13g2_fill_1 FILLER_78_1080 ();
 sg13g2_fill_1 FILLER_78_1094 ();
 sg13g2_fill_1 FILLER_78_1109 ();
 sg13g2_decap_8 FILLER_78_1121 ();
 sg13g2_fill_2 FILLER_78_1154 ();
 sg13g2_decap_8 FILLER_78_1164 ();
 sg13g2_decap_8 FILLER_78_1171 ();
 sg13g2_decap_8 FILLER_78_1178 ();
 sg13g2_fill_2 FILLER_78_1185 ();
 sg13g2_decap_4 FILLER_78_1205 ();
 sg13g2_decap_8 FILLER_78_1213 ();
 sg13g2_decap_8 FILLER_78_1220 ();
 sg13g2_decap_8 FILLER_78_1227 ();
 sg13g2_decap_8 FILLER_78_1234 ();
 sg13g2_decap_4 FILLER_78_1241 ();
 sg13g2_fill_1 FILLER_78_1245 ();
 sg13g2_decap_8 FILLER_78_1272 ();
 sg13g2_decap_8 FILLER_78_1279 ();
 sg13g2_decap_8 FILLER_78_1286 ();
 sg13g2_decap_8 FILLER_78_1293 ();
 sg13g2_decap_8 FILLER_78_1300 ();
 sg13g2_decap_8 FILLER_78_1307 ();
 sg13g2_decap_4 FILLER_78_1314 ();
 sg13g2_fill_2 FILLER_78_1318 ();
 sg13g2_decap_8 FILLER_78_1346 ();
 sg13g2_decap_8 FILLER_78_1353 ();
 sg13g2_decap_8 FILLER_78_1360 ();
 sg13g2_decap_8 FILLER_78_1367 ();
 sg13g2_decap_8 FILLER_78_1374 ();
 sg13g2_fill_1 FILLER_78_1381 ();
 sg13g2_fill_2 FILLER_78_1385 ();
 sg13g2_decap_8 FILLER_78_1413 ();
 sg13g2_decap_8 FILLER_78_1420 ();
 sg13g2_decap_8 FILLER_78_1427 ();
 sg13g2_decap_8 FILLER_78_1434 ();
 sg13g2_decap_4 FILLER_78_1458 ();
 sg13g2_decap_8 FILLER_78_1540 ();
 sg13g2_decap_8 FILLER_78_1547 ();
 sg13g2_decap_8 FILLER_78_1554 ();
 sg13g2_decap_8 FILLER_78_1561 ();
 sg13g2_decap_8 FILLER_78_1568 ();
 sg13g2_decap_8 FILLER_78_1575 ();
 sg13g2_decap_8 FILLER_78_1582 ();
 sg13g2_decap_8 FILLER_78_1589 ();
 sg13g2_decap_8 FILLER_78_1596 ();
 sg13g2_decap_8 FILLER_78_1603 ();
 sg13g2_decap_8 FILLER_78_1610 ();
 sg13g2_decap_8 FILLER_78_1617 ();
 sg13g2_decap_8 FILLER_78_1624 ();
 sg13g2_decap_8 FILLER_78_1631 ();
 sg13g2_decap_8 FILLER_78_1638 ();
 sg13g2_decap_8 FILLER_78_1645 ();
 sg13g2_decap_8 FILLER_78_1652 ();
 sg13g2_decap_8 FILLER_78_1659 ();
 sg13g2_decap_8 FILLER_78_1666 ();
 sg13g2_decap_8 FILLER_78_1673 ();
 sg13g2_decap_8 FILLER_78_1680 ();
 sg13g2_decap_8 FILLER_78_1687 ();
 sg13g2_decap_8 FILLER_78_1694 ();
 sg13g2_decap_8 FILLER_78_1701 ();
 sg13g2_decap_8 FILLER_78_1708 ();
 sg13g2_decap_8 FILLER_78_1715 ();
 sg13g2_decap_8 FILLER_78_1722 ();
 sg13g2_decap_8 FILLER_78_1729 ();
 sg13g2_decap_8 FILLER_78_1736 ();
 sg13g2_decap_8 FILLER_78_1743 ();
 sg13g2_decap_8 FILLER_78_1750 ();
 sg13g2_decap_8 FILLER_78_1757 ();
 sg13g2_decap_8 FILLER_78_1764 ();
 sg13g2_fill_2 FILLER_78_1771 ();
 sg13g2_fill_1 FILLER_78_1773 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_34 ();
 sg13g2_decap_4 FILLER_79_41 ();
 sg13g2_fill_1 FILLER_79_45 ();
 sg13g2_decap_4 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_85 ();
 sg13g2_decap_8 FILLER_79_92 ();
 sg13g2_decap_8 FILLER_79_99 ();
 sg13g2_decap_8 FILLER_79_106 ();
 sg13g2_fill_1 FILLER_79_113 ();
 sg13g2_decap_8 FILLER_79_118 ();
 sg13g2_decap_8 FILLER_79_125 ();
 sg13g2_decap_8 FILLER_79_132 ();
 sg13g2_decap_4 FILLER_79_139 ();
 sg13g2_fill_2 FILLER_79_143 ();
 sg13g2_decap_4 FILLER_79_171 ();
 sg13g2_decap_4 FILLER_79_179 ();
 sg13g2_fill_2 FILLER_79_183 ();
 sg13g2_fill_2 FILLER_79_189 ();
 sg13g2_fill_1 FILLER_79_191 ();
 sg13g2_fill_2 FILLER_79_196 ();
 sg13g2_fill_2 FILLER_79_208 ();
 sg13g2_fill_1 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_241 ();
 sg13g2_fill_2 FILLER_79_248 ();
 sg13g2_fill_1 FILLER_79_276 ();
 sg13g2_decap_8 FILLER_79_281 ();
 sg13g2_decap_8 FILLER_79_288 ();
 sg13g2_fill_1 FILLER_79_295 ();
 sg13g2_decap_8 FILLER_79_302 ();
 sg13g2_fill_1 FILLER_79_309 ();
 sg13g2_decap_8 FILLER_79_346 ();
 sg13g2_decap_8 FILLER_79_383 ();
 sg13g2_decap_8 FILLER_79_390 ();
 sg13g2_decap_8 FILLER_79_397 ();
 sg13g2_decap_8 FILLER_79_404 ();
 sg13g2_decap_8 FILLER_79_411 ();
 sg13g2_decap_8 FILLER_79_426 ();
 sg13g2_decap_8 FILLER_79_433 ();
 sg13g2_decap_4 FILLER_79_440 ();
 sg13g2_decap_8 FILLER_79_474 ();
 sg13g2_decap_8 FILLER_79_511 ();
 sg13g2_decap_4 FILLER_79_518 ();
 sg13g2_decap_8 FILLER_79_556 ();
 sg13g2_decap_8 FILLER_79_563 ();
 sg13g2_fill_2 FILLER_79_570 ();
 sg13g2_decap_8 FILLER_79_577 ();
 sg13g2_decap_8 FILLER_79_584 ();
 sg13g2_decap_8 FILLER_79_591 ();
 sg13g2_decap_8 FILLER_79_598 ();
 sg13g2_decap_4 FILLER_79_605 ();
 sg13g2_fill_2 FILLER_79_609 ();
 sg13g2_decap_8 FILLER_79_615 ();
 sg13g2_decap_8 FILLER_79_622 ();
 sg13g2_decap_8 FILLER_79_629 ();
 sg13g2_decap_8 FILLER_79_636 ();
 sg13g2_fill_2 FILLER_79_643 ();
 sg13g2_fill_1 FILLER_79_645 ();
 sg13g2_fill_2 FILLER_79_672 ();
 sg13g2_fill_1 FILLER_79_674 ();
 sg13g2_fill_2 FILLER_79_680 ();
 sg13g2_fill_2 FILLER_79_695 ();
 sg13g2_fill_1 FILLER_79_701 ();
 sg13g2_fill_2 FILLER_79_706 ();
 sg13g2_decap_8 FILLER_79_712 ();
 sg13g2_decap_8 FILLER_79_719 ();
 sg13g2_decap_8 FILLER_79_726 ();
 sg13g2_decap_8 FILLER_79_764 ();
 sg13g2_fill_2 FILLER_79_771 ();
 sg13g2_fill_1 FILLER_79_773 ();
 sg13g2_decap_8 FILLER_79_778 ();
 sg13g2_decap_8 FILLER_79_785 ();
 sg13g2_decap_8 FILLER_79_792 ();
 sg13g2_decap_8 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_806 ();
 sg13g2_fill_1 FILLER_79_813 ();
 sg13g2_decap_8 FILLER_79_818 ();
 sg13g2_decap_8 FILLER_79_825 ();
 sg13g2_decap_4 FILLER_79_832 ();
 sg13g2_fill_1 FILLER_79_836 ();
 sg13g2_decap_8 FILLER_79_841 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_decap_8 FILLER_79_855 ();
 sg13g2_decap_8 FILLER_79_862 ();
 sg13g2_decap_4 FILLER_79_869 ();
 sg13g2_fill_1 FILLER_79_873 ();
 sg13g2_fill_1 FILLER_79_900 ();
 sg13g2_decap_4 FILLER_79_905 ();
 sg13g2_fill_2 FILLER_79_909 ();
 sg13g2_decap_8 FILLER_79_937 ();
 sg13g2_decap_8 FILLER_79_944 ();
 sg13g2_decap_4 FILLER_79_951 ();
 sg13g2_fill_1 FILLER_79_955 ();
 sg13g2_decap_8 FILLER_79_986 ();
 sg13g2_decap_8 FILLER_79_993 ();
 sg13g2_decap_8 FILLER_79_1000 ();
 sg13g2_decap_8 FILLER_79_1007 ();
 sg13g2_decap_8 FILLER_79_1014 ();
 sg13g2_decap_8 FILLER_79_1021 ();
 sg13g2_decap_8 FILLER_79_1054 ();
 sg13g2_fill_2 FILLER_79_1061 ();
 sg13g2_decap_4 FILLER_79_1089 ();
 sg13g2_fill_1 FILLER_79_1097 ();
 sg13g2_decap_8 FILLER_79_1113 ();
 sg13g2_decap_8 FILLER_79_1120 ();
 sg13g2_decap_4 FILLER_79_1127 ();
 sg13g2_fill_2 FILLER_79_1131 ();
 sg13g2_decap_8 FILLER_79_1137 ();
 sg13g2_decap_8 FILLER_79_1144 ();
 sg13g2_decap_8 FILLER_79_1151 ();
 sg13g2_decap_4 FILLER_79_1158 ();
 sg13g2_fill_2 FILLER_79_1162 ();
 sg13g2_decap_8 FILLER_79_1178 ();
 sg13g2_decap_8 FILLER_79_1185 ();
 sg13g2_decap_8 FILLER_79_1192 ();
 sg13g2_fill_2 FILLER_79_1199 ();
 sg13g2_fill_1 FILLER_79_1201 ();
 sg13g2_decap_8 FILLER_79_1228 ();
 sg13g2_decap_8 FILLER_79_1235 ();
 sg13g2_decap_8 FILLER_79_1242 ();
 sg13g2_decap_4 FILLER_79_1249 ();
 sg13g2_fill_1 FILLER_79_1253 ();
 sg13g2_decap_8 FILLER_79_1258 ();
 sg13g2_decap_8 FILLER_79_1265 ();
 sg13g2_decap_8 FILLER_79_1272 ();
 sg13g2_decap_8 FILLER_79_1279 ();
 sg13g2_decap_8 FILLER_79_1286 ();
 sg13g2_decap_8 FILLER_79_1293 ();
 sg13g2_decap_8 FILLER_79_1300 ();
 sg13g2_decap_8 FILLER_79_1307 ();
 sg13g2_decap_8 FILLER_79_1314 ();
 sg13g2_decap_8 FILLER_79_1321 ();
 sg13g2_decap_8 FILLER_79_1328 ();
 sg13g2_decap_8 FILLER_79_1335 ();
 sg13g2_decap_8 FILLER_79_1342 ();
 sg13g2_decap_8 FILLER_79_1349 ();
 sg13g2_decap_8 FILLER_79_1356 ();
 sg13g2_decap_8 FILLER_79_1363 ();
 sg13g2_decap_8 FILLER_79_1370 ();
 sg13g2_decap_8 FILLER_79_1377 ();
 sg13g2_decap_8 FILLER_79_1384 ();
 sg13g2_fill_2 FILLER_79_1391 ();
 sg13g2_fill_1 FILLER_79_1393 ();
 sg13g2_decap_8 FILLER_79_1398 ();
 sg13g2_decap_8 FILLER_79_1405 ();
 sg13g2_decap_8 FILLER_79_1412 ();
 sg13g2_decap_8 FILLER_79_1419 ();
 sg13g2_decap_8 FILLER_79_1426 ();
 sg13g2_fill_1 FILLER_79_1433 ();
 sg13g2_decap_8 FILLER_79_1460 ();
 sg13g2_decap_4 FILLER_79_1467 ();
 sg13g2_fill_2 FILLER_79_1471 ();
 sg13g2_decap_8 FILLER_79_1477 ();
 sg13g2_decap_8 FILLER_79_1484 ();
 sg13g2_decap_8 FILLER_79_1491 ();
 sg13g2_decap_8 FILLER_79_1498 ();
 sg13g2_fill_2 FILLER_79_1505 ();
 sg13g2_fill_1 FILLER_79_1507 ();
 sg13g2_decap_8 FILLER_79_1512 ();
 sg13g2_decap_8 FILLER_79_1519 ();
 sg13g2_decap_8 FILLER_79_1526 ();
 sg13g2_decap_8 FILLER_79_1533 ();
 sg13g2_decap_8 FILLER_79_1540 ();
 sg13g2_decap_8 FILLER_79_1547 ();
 sg13g2_decap_8 FILLER_79_1554 ();
 sg13g2_decap_8 FILLER_79_1561 ();
 sg13g2_decap_8 FILLER_79_1568 ();
 sg13g2_decap_8 FILLER_79_1575 ();
 sg13g2_decap_8 FILLER_79_1582 ();
 sg13g2_decap_8 FILLER_79_1589 ();
 sg13g2_decap_8 FILLER_79_1596 ();
 sg13g2_decap_8 FILLER_79_1603 ();
 sg13g2_decap_8 FILLER_79_1610 ();
 sg13g2_decap_8 FILLER_79_1617 ();
 sg13g2_decap_8 FILLER_79_1624 ();
 sg13g2_decap_8 FILLER_79_1631 ();
 sg13g2_decap_8 FILLER_79_1638 ();
 sg13g2_decap_8 FILLER_79_1645 ();
 sg13g2_decap_8 FILLER_79_1652 ();
 sg13g2_decap_8 FILLER_79_1659 ();
 sg13g2_decap_8 FILLER_79_1666 ();
 sg13g2_decap_8 FILLER_79_1673 ();
 sg13g2_decap_8 FILLER_79_1680 ();
 sg13g2_decap_8 FILLER_79_1687 ();
 sg13g2_decap_8 FILLER_79_1694 ();
 sg13g2_decap_8 FILLER_79_1701 ();
 sg13g2_decap_8 FILLER_79_1708 ();
 sg13g2_decap_8 FILLER_79_1715 ();
 sg13g2_decap_8 FILLER_79_1722 ();
 sg13g2_decap_8 FILLER_79_1729 ();
 sg13g2_decap_8 FILLER_79_1736 ();
 sg13g2_decap_8 FILLER_79_1743 ();
 sg13g2_decap_8 FILLER_79_1750 ();
 sg13g2_decap_8 FILLER_79_1757 ();
 sg13g2_decap_8 FILLER_79_1764 ();
 sg13g2_fill_2 FILLER_79_1771 ();
 sg13g2_fill_1 FILLER_79_1773 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_fill_1 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_19 ();
 sg13g2_decap_8 FILLER_80_26 ();
 sg13g2_decap_8 FILLER_80_33 ();
 sg13g2_decap_8 FILLER_80_40 ();
 sg13g2_decap_4 FILLER_80_47 ();
 sg13g2_fill_2 FILLER_80_51 ();
 sg13g2_decap_8 FILLER_80_57 ();
 sg13g2_decap_8 FILLER_80_64 ();
 sg13g2_decap_4 FILLER_80_71 ();
 sg13g2_fill_1 FILLER_80_111 ();
 sg13g2_fill_1 FILLER_80_120 ();
 sg13g2_decap_4 FILLER_80_137 ();
 sg13g2_fill_2 FILLER_80_141 ();
 sg13g2_decap_8 FILLER_80_147 ();
 sg13g2_decap_8 FILLER_80_162 ();
 sg13g2_fill_2 FILLER_80_169 ();
 sg13g2_fill_1 FILLER_80_171 ();
 sg13g2_fill_2 FILLER_80_192 ();
 sg13g2_fill_1 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_203 ();
 sg13g2_fill_2 FILLER_80_210 ();
 sg13g2_decap_4 FILLER_80_217 ();
 sg13g2_fill_1 FILLER_80_221 ();
 sg13g2_fill_1 FILLER_80_226 ();
 sg13g2_fill_1 FILLER_80_239 ();
 sg13g2_fill_1 FILLER_80_244 ();
 sg13g2_fill_2 FILLER_80_261 ();
 sg13g2_decap_8 FILLER_80_271 ();
 sg13g2_decap_8 FILLER_80_278 ();
 sg13g2_decap_8 FILLER_80_285 ();
 sg13g2_decap_8 FILLER_80_292 ();
 sg13g2_decap_8 FILLER_80_299 ();
 sg13g2_decap_8 FILLER_80_306 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_332 ();
 sg13g2_decap_8 FILLER_80_339 ();
 sg13g2_decap_8 FILLER_80_346 ();
 sg13g2_decap_8 FILLER_80_353 ();
 sg13g2_decap_4 FILLER_80_360 ();
 sg13g2_decap_4 FILLER_80_376 ();
 sg13g2_fill_2 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_fill_1 FILLER_80_398 ();
 sg13g2_decap_8 FILLER_80_403 ();
 sg13g2_fill_1 FILLER_80_410 ();
 sg13g2_decap_8 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_444 ();
 sg13g2_fill_2 FILLER_80_451 ();
 sg13g2_fill_1 FILLER_80_453 ();
 sg13g2_decap_8 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_decap_8 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_479 ();
 sg13g2_decap_4 FILLER_80_486 ();
 sg13g2_fill_2 FILLER_80_490 ();
 sg13g2_decap_8 FILLER_80_496 ();
 sg13g2_decap_8 FILLER_80_503 ();
 sg13g2_decap_8 FILLER_80_510 ();
 sg13g2_decap_8 FILLER_80_517 ();
 sg13g2_decap_8 FILLER_80_524 ();
 sg13g2_fill_2 FILLER_80_531 ();
 sg13g2_decap_8 FILLER_80_537 ();
 sg13g2_decap_8 FILLER_80_544 ();
 sg13g2_fill_2 FILLER_80_551 ();
 sg13g2_decap_8 FILLER_80_583 ();
 sg13g2_decap_8 FILLER_80_590 ();
 sg13g2_decap_8 FILLER_80_597 ();
 sg13g2_decap_8 FILLER_80_604 ();
 sg13g2_decap_8 FILLER_80_611 ();
 sg13g2_decap_8 FILLER_80_618 ();
 sg13g2_decap_8 FILLER_80_625 ();
 sg13g2_decap_8 FILLER_80_632 ();
 sg13g2_decap_8 FILLER_80_639 ();
 sg13g2_decap_8 FILLER_80_646 ();
 sg13g2_fill_1 FILLER_80_653 ();
 sg13g2_decap_8 FILLER_80_658 ();
 sg13g2_decap_8 FILLER_80_665 ();
 sg13g2_decap_8 FILLER_80_672 ();
 sg13g2_decap_8 FILLER_80_679 ();
 sg13g2_fill_2 FILLER_80_692 ();
 sg13g2_decap_8 FILLER_80_713 ();
 sg13g2_decap_8 FILLER_80_720 ();
 sg13g2_decap_8 FILLER_80_727 ();
 sg13g2_decap_8 FILLER_80_734 ();
 sg13g2_decap_8 FILLER_80_745 ();
 sg13g2_decap_8 FILLER_80_752 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_decap_8 FILLER_80_766 ();
 sg13g2_decap_8 FILLER_80_773 ();
 sg13g2_decap_8 FILLER_80_780 ();
 sg13g2_decap_8 FILLER_80_787 ();
 sg13g2_decap_8 FILLER_80_794 ();
 sg13g2_decap_8 FILLER_80_801 ();
 sg13g2_decap_8 FILLER_80_808 ();
 sg13g2_decap_8 FILLER_80_815 ();
 sg13g2_decap_8 FILLER_80_822 ();
 sg13g2_decap_8 FILLER_80_829 ();
 sg13g2_decap_8 FILLER_80_836 ();
 sg13g2_decap_8 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_850 ();
 sg13g2_decap_8 FILLER_80_857 ();
 sg13g2_decap_8 FILLER_80_864 ();
 sg13g2_decap_8 FILLER_80_871 ();
 sg13g2_fill_2 FILLER_80_878 ();
 sg13g2_decap_8 FILLER_80_884 ();
 sg13g2_decap_8 FILLER_80_891 ();
 sg13g2_decap_8 FILLER_80_898 ();
 sg13g2_decap_8 FILLER_80_905 ();
 sg13g2_decap_8 FILLER_80_912 ();
 sg13g2_fill_1 FILLER_80_919 ();
 sg13g2_decap_8 FILLER_80_924 ();
 sg13g2_decap_8 FILLER_80_931 ();
 sg13g2_decap_8 FILLER_80_938 ();
 sg13g2_decap_8 FILLER_80_945 ();
 sg13g2_decap_8 FILLER_80_952 ();
 sg13g2_decap_4 FILLER_80_959 ();
 sg13g2_fill_2 FILLER_80_963 ();
 sg13g2_decap_8 FILLER_80_969 ();
 sg13g2_decap_8 FILLER_80_976 ();
 sg13g2_decap_8 FILLER_80_983 ();
 sg13g2_decap_8 FILLER_80_990 ();
 sg13g2_decap_8 FILLER_80_997 ();
 sg13g2_decap_8 FILLER_80_1004 ();
 sg13g2_decap_8 FILLER_80_1011 ();
 sg13g2_decap_8 FILLER_80_1018 ();
 sg13g2_decap_8 FILLER_80_1025 ();
 sg13g2_decap_8 FILLER_80_1032 ();
 sg13g2_decap_8 FILLER_80_1039 ();
 sg13g2_decap_8 FILLER_80_1046 ();
 sg13g2_decap_8 FILLER_80_1053 ();
 sg13g2_decap_8 FILLER_80_1060 ();
 sg13g2_decap_4 FILLER_80_1067 ();
 sg13g2_decap_8 FILLER_80_1075 ();
 sg13g2_decap_8 FILLER_80_1082 ();
 sg13g2_decap_8 FILLER_80_1089 ();
 sg13g2_decap_8 FILLER_80_1096 ();
 sg13g2_decap_8 FILLER_80_1103 ();
 sg13g2_decap_8 FILLER_80_1110 ();
 sg13g2_decap_8 FILLER_80_1117 ();
 sg13g2_decap_8 FILLER_80_1124 ();
 sg13g2_decap_8 FILLER_80_1131 ();
 sg13g2_decap_8 FILLER_80_1138 ();
 sg13g2_decap_8 FILLER_80_1145 ();
 sg13g2_fill_1 FILLER_80_1152 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_decap_8 FILLER_80_1186 ();
 sg13g2_decap_8 FILLER_80_1193 ();
 sg13g2_decap_8 FILLER_80_1200 ();
 sg13g2_decap_8 FILLER_80_1207 ();
 sg13g2_decap_8 FILLER_80_1214 ();
 sg13g2_decap_8 FILLER_80_1221 ();
 sg13g2_decap_8 FILLER_80_1228 ();
 sg13g2_decap_8 FILLER_80_1235 ();
 sg13g2_decap_8 FILLER_80_1242 ();
 sg13g2_decap_8 FILLER_80_1249 ();
 sg13g2_decap_8 FILLER_80_1256 ();
 sg13g2_decap_8 FILLER_80_1263 ();
 sg13g2_decap_8 FILLER_80_1270 ();
 sg13g2_decap_8 FILLER_80_1277 ();
 sg13g2_decap_8 FILLER_80_1284 ();
 sg13g2_decap_8 FILLER_80_1291 ();
 sg13g2_decap_8 FILLER_80_1298 ();
 sg13g2_decap_8 FILLER_80_1305 ();
 sg13g2_decap_8 FILLER_80_1312 ();
 sg13g2_decap_8 FILLER_80_1319 ();
 sg13g2_decap_8 FILLER_80_1326 ();
 sg13g2_decap_8 FILLER_80_1333 ();
 sg13g2_decap_8 FILLER_80_1340 ();
 sg13g2_decap_8 FILLER_80_1347 ();
 sg13g2_decap_8 FILLER_80_1354 ();
 sg13g2_decap_8 FILLER_80_1361 ();
 sg13g2_decap_8 FILLER_80_1368 ();
 sg13g2_decap_8 FILLER_80_1375 ();
 sg13g2_decap_8 FILLER_80_1382 ();
 sg13g2_decap_8 FILLER_80_1389 ();
 sg13g2_decap_8 FILLER_80_1396 ();
 sg13g2_decap_8 FILLER_80_1403 ();
 sg13g2_decap_8 FILLER_80_1410 ();
 sg13g2_decap_8 FILLER_80_1417 ();
 sg13g2_decap_8 FILLER_80_1424 ();
 sg13g2_decap_8 FILLER_80_1431 ();
 sg13g2_decap_8 FILLER_80_1438 ();
 sg13g2_decap_8 FILLER_80_1445 ();
 sg13g2_decap_8 FILLER_80_1452 ();
 sg13g2_decap_8 FILLER_80_1459 ();
 sg13g2_decap_8 FILLER_80_1466 ();
 sg13g2_decap_8 FILLER_80_1473 ();
 sg13g2_decap_8 FILLER_80_1480 ();
 sg13g2_decap_8 FILLER_80_1487 ();
 sg13g2_decap_8 FILLER_80_1494 ();
 sg13g2_decap_8 FILLER_80_1501 ();
 sg13g2_decap_8 FILLER_80_1508 ();
 sg13g2_decap_8 FILLER_80_1515 ();
 sg13g2_decap_8 FILLER_80_1522 ();
 sg13g2_decap_8 FILLER_80_1529 ();
 sg13g2_decap_8 FILLER_80_1536 ();
 sg13g2_decap_8 FILLER_80_1543 ();
 sg13g2_decap_8 FILLER_80_1550 ();
 sg13g2_decap_8 FILLER_80_1557 ();
 sg13g2_decap_8 FILLER_80_1564 ();
 sg13g2_decap_8 FILLER_80_1571 ();
 sg13g2_decap_8 FILLER_80_1578 ();
 sg13g2_decap_8 FILLER_80_1585 ();
 sg13g2_decap_8 FILLER_80_1592 ();
 sg13g2_decap_8 FILLER_80_1599 ();
 sg13g2_decap_8 FILLER_80_1606 ();
 sg13g2_decap_8 FILLER_80_1613 ();
 sg13g2_decap_8 FILLER_80_1620 ();
 sg13g2_decap_8 FILLER_80_1627 ();
 sg13g2_decap_8 FILLER_80_1634 ();
 sg13g2_decap_8 FILLER_80_1641 ();
 sg13g2_decap_8 FILLER_80_1648 ();
 sg13g2_decap_8 FILLER_80_1655 ();
 sg13g2_decap_8 FILLER_80_1662 ();
 sg13g2_decap_8 FILLER_80_1669 ();
 sg13g2_decap_8 FILLER_80_1676 ();
 sg13g2_decap_8 FILLER_80_1683 ();
 sg13g2_decap_8 FILLER_80_1690 ();
 sg13g2_decap_8 FILLER_80_1697 ();
 sg13g2_decap_8 FILLER_80_1704 ();
 sg13g2_decap_8 FILLER_80_1711 ();
 sg13g2_decap_8 FILLER_80_1718 ();
 sg13g2_decap_8 FILLER_80_1725 ();
 sg13g2_decap_8 FILLER_80_1732 ();
 sg13g2_decap_8 FILLER_80_1739 ();
 sg13g2_decap_8 FILLER_80_1746 ();
 sg13g2_decap_8 FILLER_80_1753 ();
 sg13g2_decap_8 FILLER_80_1760 ();
 sg13g2_decap_8 FILLER_80_1767 ();
endmodule
