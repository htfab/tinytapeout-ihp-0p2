module tt_um_htfab_rotfpga2 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire clknet_0_clk;
 wire net133;
 wire \g.cfg_d ;
 wire \g.cfg_h ;
 wire \g.cfg_v ;
 wire \g.g_y[0].g_x[0].t.in_lb ;
 wire \g.g_y[0].g_x[0].t.out_sc ;
 wire \g.g_y[0].g_x[0].t.r_d ;
 wire \g.g_y[0].g_x[0].t.r_ghl ;
 wire \g.g_y[0].g_x[0].t.r_gnl ;
 wire \g.g_y[0].g_x[0].t.r_h ;
 wire \g.g_y[0].g_x[0].t.r_v ;
 wire \g.g_y[0].g_x[0].t.w_dh ;
 wire \g.g_y[0].g_x[0].t.w_na ;
 wire \g.g_y[0].g_x[0].t.w_si ;
 wire \g.g_y[0].g_x[1].t.out_sc ;
 wire \g.g_y[0].g_x[1].t.r_d ;
 wire \g.g_y[0].g_x[1].t.r_h ;
 wire \g.g_y[0].g_x[1].t.r_v ;
 wire \g.g_y[0].g_x[1].t.w_si ;
 wire \g.g_y[0].g_x[2].t.in_lb ;
 wire \g.g_y[0].g_x[2].t.out_sc ;
 wire \g.g_y[0].g_x[2].t.r_d ;
 wire \g.g_y[0].g_x[2].t.r_ghl ;
 wire \g.g_y[0].g_x[2].t.r_gnl ;
 wire \g.g_y[0].g_x[2].t.r_h ;
 wire \g.g_y[0].g_x[2].t.r_v ;
 wire \g.g_y[0].g_x[2].t.w_dh ;
 wire \g.g_y[0].g_x[2].t.w_na ;
 wire \g.g_y[0].g_x[2].t.w_si ;
 wire \g.g_y[0].g_x[3].t.out_sc ;
 wire \g.g_y[0].g_x[3].t.r_d ;
 wire \g.g_y[0].g_x[3].t.r_h ;
 wire \g.g_y[0].g_x[3].t.r_v ;
 wire \g.g_y[0].g_x[3].t.w_si ;
 wire \g.g_y[0].g_x[4].t.out_sc ;
 wire \g.g_y[0].g_x[4].t.r_d ;
 wire \g.g_y[0].g_x[4].t.r_ghl ;
 wire \g.g_y[0].g_x[4].t.r_gnl ;
 wire \g.g_y[0].g_x[4].t.r_h ;
 wire \g.g_y[0].g_x[4].t.r_v ;
 wire \g.g_y[0].g_x[4].t.w_dh ;
 wire \g.g_y[0].g_x[4].t.w_na ;
 wire \g.g_y[0].g_x[4].t.w_si ;
 wire \g.g_y[0].g_x[5].t.out_sc ;
 wire \g.g_y[0].g_x[5].t.r_d ;
 wire \g.g_y[0].g_x[5].t.r_h ;
 wire \g.g_y[0].g_x[5].t.r_v ;
 wire \g.g_y[0].g_x[5].t.w_si ;
 wire \g.g_y[0].g_x[6].t.out_sc ;
 wire \g.g_y[0].g_x[6].t.r_d ;
 wire \g.g_y[0].g_x[6].t.r_ghl ;
 wire \g.g_y[0].g_x[6].t.r_gnl ;
 wire \g.g_y[0].g_x[6].t.r_h ;
 wire \g.g_y[0].g_x[6].t.r_v ;
 wire \g.g_y[0].g_x[6].t.w_dh ;
 wire \g.g_y[0].g_x[6].t.w_na ;
 wire \g.g_y[0].g_x[6].t.w_si ;
 wire \g.g_y[0].g_x[7].t.out_r ;
 wire \g.g_y[0].g_x[7].t.out_sc ;
 wire \g.g_y[0].g_x[7].t.r_d ;
 wire \g.g_y[0].g_x[7].t.r_h ;
 wire \g.g_y[0].g_x[7].t.r_v ;
 wire \g.g_y[0].g_x[7].t.w_si ;
 wire \g.g_y[1].g_x[0].t.out_sc ;
 wire \g.g_y[1].g_x[0].t.r_d ;
 wire \g.g_y[1].g_x[0].t.r_h ;
 wire \g.g_y[1].g_x[0].t.r_v ;
 wire \g.g_y[1].g_x[0].t.w_si ;
 wire \g.g_y[1].g_x[1].t.in_lb ;
 wire \g.g_y[1].g_x[1].t.out_sc ;
 wire \g.g_y[1].g_x[1].t.r_d ;
 wire \g.g_y[1].g_x[1].t.r_ghl ;
 wire \g.g_y[1].g_x[1].t.r_gnl ;
 wire \g.g_y[1].g_x[1].t.r_h ;
 wire \g.g_y[1].g_x[1].t.r_v ;
 wire \g.g_y[1].g_x[1].t.w_dh ;
 wire \g.g_y[1].g_x[1].t.w_na ;
 wire \g.g_y[1].g_x[1].t.w_si ;
 wire \g.g_y[1].g_x[2].t.out_sc ;
 wire \g.g_y[1].g_x[2].t.r_d ;
 wire \g.g_y[1].g_x[2].t.r_h ;
 wire \g.g_y[1].g_x[2].t.r_v ;
 wire \g.g_y[1].g_x[2].t.w_si ;
 wire \g.g_y[1].g_x[3].t.in_lb ;
 wire \g.g_y[1].g_x[3].t.out_sc ;
 wire \g.g_y[1].g_x[3].t.r_d ;
 wire \g.g_y[1].g_x[3].t.r_ghl ;
 wire \g.g_y[1].g_x[3].t.r_gnl ;
 wire \g.g_y[1].g_x[3].t.r_h ;
 wire \g.g_y[1].g_x[3].t.r_v ;
 wire \g.g_y[1].g_x[3].t.w_dh ;
 wire \g.g_y[1].g_x[3].t.w_na ;
 wire \g.g_y[1].g_x[3].t.w_si ;
 wire \g.g_y[1].g_x[4].t.out_sc ;
 wire \g.g_y[1].g_x[4].t.r_d ;
 wire \g.g_y[1].g_x[4].t.r_h ;
 wire \g.g_y[1].g_x[4].t.r_v ;
 wire \g.g_y[1].g_x[4].t.w_si ;
 wire \g.g_y[1].g_x[5].t.out_sc ;
 wire \g.g_y[1].g_x[5].t.r_d ;
 wire \g.g_y[1].g_x[5].t.r_ghl ;
 wire \g.g_y[1].g_x[5].t.r_gnl ;
 wire \g.g_y[1].g_x[5].t.r_h ;
 wire \g.g_y[1].g_x[5].t.r_v ;
 wire \g.g_y[1].g_x[5].t.w_dh ;
 wire \g.g_y[1].g_x[5].t.w_na ;
 wire \g.g_y[1].g_x[5].t.w_si ;
 wire \g.g_y[1].g_x[6].t.out_sc ;
 wire \g.g_y[1].g_x[6].t.r_d ;
 wire \g.g_y[1].g_x[6].t.r_h ;
 wire \g.g_y[1].g_x[6].t.r_v ;
 wire \g.g_y[1].g_x[6].t.w_si ;
 wire \g.g_y[1].g_x[7].t.out_r ;
 wire \g.g_y[1].g_x[7].t.out_sc ;
 wire \g.g_y[1].g_x[7].t.r_d ;
 wire \g.g_y[1].g_x[7].t.r_ghl ;
 wire \g.g_y[1].g_x[7].t.r_gnl ;
 wire \g.g_y[1].g_x[7].t.r_h ;
 wire \g.g_y[1].g_x[7].t.r_v ;
 wire \g.g_y[1].g_x[7].t.w_dh ;
 wire \g.g_y[1].g_x[7].t.w_na ;
 wire \g.g_y[1].g_x[7].t.w_si ;
 wire \g.g_y[2].g_x[0].t.out_sc ;
 wire \g.g_y[2].g_x[0].t.r_d ;
 wire \g.g_y[2].g_x[0].t.r_ghl ;
 wire \g.g_y[2].g_x[0].t.r_gnl ;
 wire \g.g_y[2].g_x[0].t.r_h ;
 wire \g.g_y[2].g_x[0].t.r_v ;
 wire \g.g_y[2].g_x[0].t.w_dh ;
 wire \g.g_y[2].g_x[0].t.w_na ;
 wire \g.g_y[2].g_x[0].t.w_si ;
 wire \g.g_y[2].g_x[1].t.out_sc ;
 wire \g.g_y[2].g_x[1].t.r_d ;
 wire \g.g_y[2].g_x[1].t.r_h ;
 wire \g.g_y[2].g_x[1].t.r_v ;
 wire \g.g_y[2].g_x[1].t.w_si ;
 wire \g.g_y[2].g_x[2].t.out_sc ;
 wire \g.g_y[2].g_x[2].t.r_d ;
 wire \g.g_y[2].g_x[2].t.r_ghl ;
 wire \g.g_y[2].g_x[2].t.r_gnl ;
 wire \g.g_y[2].g_x[2].t.r_h ;
 wire \g.g_y[2].g_x[2].t.r_v ;
 wire \g.g_y[2].g_x[2].t.w_dh ;
 wire \g.g_y[2].g_x[2].t.w_na ;
 wire \g.g_y[2].g_x[2].t.w_si ;
 wire \g.g_y[2].g_x[3].t.out_sc ;
 wire \g.g_y[2].g_x[3].t.r_d ;
 wire \g.g_y[2].g_x[3].t.r_h ;
 wire \g.g_y[2].g_x[3].t.r_v ;
 wire \g.g_y[2].g_x[3].t.w_si ;
 wire \g.g_y[2].g_x[4].t.out_sc ;
 wire \g.g_y[2].g_x[4].t.r_d ;
 wire \g.g_y[2].g_x[4].t.r_ghl ;
 wire \g.g_y[2].g_x[4].t.r_gnl ;
 wire \g.g_y[2].g_x[4].t.r_h ;
 wire \g.g_y[2].g_x[4].t.r_v ;
 wire \g.g_y[2].g_x[4].t.w_dh ;
 wire \g.g_y[2].g_x[4].t.w_na ;
 wire \g.g_y[2].g_x[4].t.w_si ;
 wire \g.g_y[2].g_x[5].t.out_sc ;
 wire \g.g_y[2].g_x[5].t.r_d ;
 wire \g.g_y[2].g_x[5].t.r_h ;
 wire \g.g_y[2].g_x[5].t.r_v ;
 wire \g.g_y[2].g_x[5].t.w_si ;
 wire \g.g_y[2].g_x[6].t.out_sc ;
 wire \g.g_y[2].g_x[6].t.r_d ;
 wire \g.g_y[2].g_x[6].t.r_ghl ;
 wire \g.g_y[2].g_x[6].t.r_gnl ;
 wire \g.g_y[2].g_x[6].t.r_h ;
 wire \g.g_y[2].g_x[6].t.r_v ;
 wire \g.g_y[2].g_x[6].t.w_dh ;
 wire \g.g_y[2].g_x[6].t.w_na ;
 wire \g.g_y[2].g_x[6].t.w_si ;
 wire \g.g_y[2].g_x[7].t.out_r ;
 wire \g.g_y[2].g_x[7].t.out_sc ;
 wire \g.g_y[2].g_x[7].t.r_d ;
 wire \g.g_y[2].g_x[7].t.r_h ;
 wire \g.g_y[2].g_x[7].t.r_v ;
 wire \g.g_y[2].g_x[7].t.w_si ;
 wire \g.g_y[3].g_x[0].t.out_sc ;
 wire \g.g_y[3].g_x[0].t.r_d ;
 wire \g.g_y[3].g_x[0].t.r_h ;
 wire \g.g_y[3].g_x[0].t.r_v ;
 wire \g.g_y[3].g_x[0].t.w_si ;
 wire \g.g_y[3].g_x[1].t.out_sc ;
 wire \g.g_y[3].g_x[1].t.r_d ;
 wire \g.g_y[3].g_x[1].t.r_ghl ;
 wire \g.g_y[3].g_x[1].t.r_gnl ;
 wire \g.g_y[3].g_x[1].t.r_h ;
 wire \g.g_y[3].g_x[1].t.r_v ;
 wire \g.g_y[3].g_x[1].t.w_dh ;
 wire \g.g_y[3].g_x[1].t.w_na ;
 wire \g.g_y[3].g_x[1].t.w_si ;
 wire \g.g_y[3].g_x[2].t.out_sc ;
 wire \g.g_y[3].g_x[2].t.r_d ;
 wire \g.g_y[3].g_x[2].t.r_h ;
 wire \g.g_y[3].g_x[2].t.r_v ;
 wire \g.g_y[3].g_x[2].t.w_si ;
 wire \g.g_y[3].g_x[3].t.out_sc ;
 wire \g.g_y[3].g_x[3].t.r_d ;
 wire \g.g_y[3].g_x[3].t.r_ghl ;
 wire \g.g_y[3].g_x[3].t.r_gnl ;
 wire \g.g_y[3].g_x[3].t.r_h ;
 wire \g.g_y[3].g_x[3].t.r_v ;
 wire \g.g_y[3].g_x[3].t.w_dh ;
 wire \g.g_y[3].g_x[3].t.w_na ;
 wire \g.g_y[3].g_x[3].t.w_si ;
 wire \g.g_y[3].g_x[4].t.out_sc ;
 wire \g.g_y[3].g_x[4].t.r_d ;
 wire \g.g_y[3].g_x[4].t.r_h ;
 wire \g.g_y[3].g_x[4].t.r_v ;
 wire \g.g_y[3].g_x[4].t.w_si ;
 wire \g.g_y[3].g_x[5].t.out_sc ;
 wire \g.g_y[3].g_x[5].t.r_d ;
 wire \g.g_y[3].g_x[5].t.r_ghl ;
 wire \g.g_y[3].g_x[5].t.r_gnl ;
 wire \g.g_y[3].g_x[5].t.r_h ;
 wire \g.g_y[3].g_x[5].t.r_v ;
 wire \g.g_y[3].g_x[5].t.w_dh ;
 wire \g.g_y[3].g_x[5].t.w_na ;
 wire \g.g_y[3].g_x[5].t.w_si ;
 wire \g.g_y[3].g_x[6].t.out_sc ;
 wire \g.g_y[3].g_x[6].t.r_d ;
 wire \g.g_y[3].g_x[6].t.r_h ;
 wire \g.g_y[3].g_x[6].t.r_v ;
 wire \g.g_y[3].g_x[6].t.w_si ;
 wire \g.g_y[3].g_x[7].t.out_r ;
 wire \g.g_y[3].g_x[7].t.out_sc ;
 wire \g.g_y[3].g_x[7].t.r_d ;
 wire \g.g_y[3].g_x[7].t.r_ghl ;
 wire \g.g_y[3].g_x[7].t.r_gnl ;
 wire \g.g_y[3].g_x[7].t.r_h ;
 wire \g.g_y[3].g_x[7].t.r_v ;
 wire \g.g_y[3].g_x[7].t.w_dh ;
 wire \g.g_y[3].g_x[7].t.w_na ;
 wire \g.g_y[3].g_x[7].t.w_si ;
 wire \g.g_y[4].g_x[0].t.out_sc ;
 wire \g.g_y[4].g_x[0].t.r_d ;
 wire \g.g_y[4].g_x[0].t.r_ghl ;
 wire \g.g_y[4].g_x[0].t.r_gnl ;
 wire \g.g_y[4].g_x[0].t.r_h ;
 wire \g.g_y[4].g_x[0].t.r_v ;
 wire \g.g_y[4].g_x[0].t.w_dh ;
 wire \g.g_y[4].g_x[0].t.w_na ;
 wire \g.g_y[4].g_x[0].t.w_si ;
 wire \g.g_y[4].g_x[1].t.out_sc ;
 wire \g.g_y[4].g_x[1].t.r_d ;
 wire \g.g_y[4].g_x[1].t.r_h ;
 wire \g.g_y[4].g_x[1].t.r_v ;
 wire \g.g_y[4].g_x[1].t.w_si ;
 wire \g.g_y[4].g_x[2].t.out_sc ;
 wire \g.g_y[4].g_x[2].t.r_d ;
 wire \g.g_y[4].g_x[2].t.r_ghl ;
 wire \g.g_y[4].g_x[2].t.r_gnl ;
 wire \g.g_y[4].g_x[2].t.r_h ;
 wire \g.g_y[4].g_x[2].t.r_v ;
 wire \g.g_y[4].g_x[2].t.w_dh ;
 wire \g.g_y[4].g_x[2].t.w_na ;
 wire \g.g_y[4].g_x[2].t.w_si ;
 wire \g.g_y[4].g_x[3].t.out_sc ;
 wire \g.g_y[4].g_x[3].t.r_d ;
 wire \g.g_y[4].g_x[3].t.r_h ;
 wire \g.g_y[4].g_x[3].t.r_v ;
 wire \g.g_y[4].g_x[3].t.w_si ;
 wire \g.g_y[4].g_x[4].t.out_sc ;
 wire \g.g_y[4].g_x[4].t.r_d ;
 wire \g.g_y[4].g_x[4].t.r_ghl ;
 wire \g.g_y[4].g_x[4].t.r_gnl ;
 wire \g.g_y[4].g_x[4].t.r_h ;
 wire \g.g_y[4].g_x[4].t.r_v ;
 wire \g.g_y[4].g_x[4].t.w_dh ;
 wire \g.g_y[4].g_x[4].t.w_na ;
 wire \g.g_y[4].g_x[4].t.w_si ;
 wire \g.g_y[4].g_x[5].t.out_sc ;
 wire \g.g_y[4].g_x[5].t.r_d ;
 wire \g.g_y[4].g_x[5].t.r_h ;
 wire \g.g_y[4].g_x[5].t.r_v ;
 wire \g.g_y[4].g_x[5].t.w_si ;
 wire \g.g_y[4].g_x[6].t.out_sc ;
 wire \g.g_y[4].g_x[6].t.r_d ;
 wire \g.g_y[4].g_x[6].t.r_ghl ;
 wire \g.g_y[4].g_x[6].t.r_gnl ;
 wire \g.g_y[4].g_x[6].t.r_h ;
 wire \g.g_y[4].g_x[6].t.r_v ;
 wire \g.g_y[4].g_x[6].t.w_dh ;
 wire \g.g_y[4].g_x[6].t.w_na ;
 wire \g.g_y[4].g_x[6].t.w_si ;
 wire \g.g_y[4].g_x[7].t.out_r ;
 wire \g.g_y[4].g_x[7].t.out_sc ;
 wire \g.g_y[4].g_x[7].t.r_d ;
 wire \g.g_y[4].g_x[7].t.r_h ;
 wire \g.g_y[4].g_x[7].t.r_v ;
 wire \g.g_y[4].g_x[7].t.w_si ;
 wire \g.g_y[5].g_x[0].t.out_sc ;
 wire \g.g_y[5].g_x[0].t.r_d ;
 wire \g.g_y[5].g_x[0].t.r_h ;
 wire \g.g_y[5].g_x[0].t.r_v ;
 wire \g.g_y[5].g_x[0].t.w_si ;
 wire \g.g_y[5].g_x[1].t.out_sc ;
 wire \g.g_y[5].g_x[1].t.r_d ;
 wire \g.g_y[5].g_x[1].t.r_ghl ;
 wire \g.g_y[5].g_x[1].t.r_gnl ;
 wire \g.g_y[5].g_x[1].t.r_h ;
 wire \g.g_y[5].g_x[1].t.r_v ;
 wire \g.g_y[5].g_x[1].t.w_dh ;
 wire \g.g_y[5].g_x[1].t.w_na ;
 wire \g.g_y[5].g_x[1].t.w_si ;
 wire \g.g_y[5].g_x[2].t.out_sc ;
 wire \g.g_y[5].g_x[2].t.r_d ;
 wire \g.g_y[5].g_x[2].t.r_h ;
 wire \g.g_y[5].g_x[2].t.r_v ;
 wire \g.g_y[5].g_x[2].t.w_si ;
 wire \g.g_y[5].g_x[3].t.out_sc ;
 wire \g.g_y[5].g_x[3].t.r_d ;
 wire \g.g_y[5].g_x[3].t.r_ghl ;
 wire \g.g_y[5].g_x[3].t.r_gnl ;
 wire \g.g_y[5].g_x[3].t.r_h ;
 wire \g.g_y[5].g_x[3].t.r_v ;
 wire \g.g_y[5].g_x[3].t.w_dh ;
 wire \g.g_y[5].g_x[3].t.w_na ;
 wire \g.g_y[5].g_x[3].t.w_si ;
 wire \g.g_y[5].g_x[4].t.out_sc ;
 wire \g.g_y[5].g_x[4].t.r_d ;
 wire \g.g_y[5].g_x[4].t.r_h ;
 wire \g.g_y[5].g_x[4].t.r_v ;
 wire \g.g_y[5].g_x[4].t.w_si ;
 wire \g.g_y[5].g_x[5].t.out_sc ;
 wire \g.g_y[5].g_x[5].t.r_d ;
 wire \g.g_y[5].g_x[5].t.r_ghl ;
 wire \g.g_y[5].g_x[5].t.r_gnl ;
 wire \g.g_y[5].g_x[5].t.r_h ;
 wire \g.g_y[5].g_x[5].t.r_v ;
 wire \g.g_y[5].g_x[5].t.w_dh ;
 wire \g.g_y[5].g_x[5].t.w_na ;
 wire \g.g_y[5].g_x[5].t.w_si ;
 wire \g.g_y[5].g_x[6].t.out_sc ;
 wire \g.g_y[5].g_x[6].t.r_d ;
 wire \g.g_y[5].g_x[6].t.r_h ;
 wire \g.g_y[5].g_x[6].t.r_v ;
 wire \g.g_y[5].g_x[6].t.w_si ;
 wire \g.g_y[5].g_x[7].t.out_r ;
 wire \g.g_y[5].g_x[7].t.out_sc ;
 wire \g.g_y[5].g_x[7].t.r_d ;
 wire \g.g_y[5].g_x[7].t.r_ghl ;
 wire \g.g_y[5].g_x[7].t.r_gnl ;
 wire \g.g_y[5].g_x[7].t.r_h ;
 wire \g.g_y[5].g_x[7].t.r_v ;
 wire \g.g_y[5].g_x[7].t.w_dh ;
 wire \g.g_y[5].g_x[7].t.w_na ;
 wire \g.g_y[5].g_x[7].t.w_si ;
 wire \g.g_y[6].g_x[0].t.out_sc ;
 wire \g.g_y[6].g_x[0].t.r_d ;
 wire \g.g_y[6].g_x[0].t.r_ghl ;
 wire \g.g_y[6].g_x[0].t.r_gnl ;
 wire \g.g_y[6].g_x[0].t.r_h ;
 wire \g.g_y[6].g_x[0].t.r_v ;
 wire \g.g_y[6].g_x[0].t.w_dh ;
 wire \g.g_y[6].g_x[0].t.w_na ;
 wire \g.g_y[6].g_x[0].t.w_si ;
 wire \g.g_y[6].g_x[1].t.out_sc ;
 wire \g.g_y[6].g_x[1].t.r_d ;
 wire \g.g_y[6].g_x[1].t.r_h ;
 wire \g.g_y[6].g_x[1].t.r_v ;
 wire \g.g_y[6].g_x[1].t.w_si ;
 wire \g.g_y[6].g_x[2].t.out_sc ;
 wire \g.g_y[6].g_x[2].t.r_d ;
 wire \g.g_y[6].g_x[2].t.r_ghl ;
 wire \g.g_y[6].g_x[2].t.r_gnl ;
 wire \g.g_y[6].g_x[2].t.r_h ;
 wire \g.g_y[6].g_x[2].t.r_v ;
 wire \g.g_y[6].g_x[2].t.w_dh ;
 wire \g.g_y[6].g_x[2].t.w_na ;
 wire \g.g_y[6].g_x[2].t.w_si ;
 wire \g.g_y[6].g_x[3].t.out_sc ;
 wire \g.g_y[6].g_x[3].t.r_d ;
 wire \g.g_y[6].g_x[3].t.r_h ;
 wire \g.g_y[6].g_x[3].t.r_v ;
 wire \g.g_y[6].g_x[3].t.w_si ;
 wire \g.g_y[6].g_x[4].t.out_sc ;
 wire \g.g_y[6].g_x[4].t.r_d ;
 wire \g.g_y[6].g_x[4].t.r_ghl ;
 wire \g.g_y[6].g_x[4].t.r_gnl ;
 wire \g.g_y[6].g_x[4].t.r_h ;
 wire \g.g_y[6].g_x[4].t.r_v ;
 wire \g.g_y[6].g_x[4].t.w_dh ;
 wire \g.g_y[6].g_x[4].t.w_na ;
 wire \g.g_y[6].g_x[4].t.w_si ;
 wire \g.g_y[6].g_x[5].t.out_sc ;
 wire \g.g_y[6].g_x[5].t.r_d ;
 wire \g.g_y[6].g_x[5].t.r_h ;
 wire \g.g_y[6].g_x[5].t.r_v ;
 wire \g.g_y[6].g_x[5].t.w_si ;
 wire \g.g_y[6].g_x[6].t.out_sc ;
 wire \g.g_y[6].g_x[6].t.r_d ;
 wire \g.g_y[6].g_x[6].t.r_ghl ;
 wire \g.g_y[6].g_x[6].t.r_gnl ;
 wire \g.g_y[6].g_x[6].t.r_h ;
 wire \g.g_y[6].g_x[6].t.r_v ;
 wire \g.g_y[6].g_x[6].t.w_dh ;
 wire \g.g_y[6].g_x[6].t.w_na ;
 wire \g.g_y[6].g_x[6].t.w_si ;
 wire \g.g_y[6].g_x[7].t.out_r ;
 wire \g.g_y[6].g_x[7].t.out_sc ;
 wire \g.g_y[6].g_x[7].t.r_d ;
 wire \g.g_y[6].g_x[7].t.r_h ;
 wire \g.g_y[6].g_x[7].t.r_v ;
 wire \g.g_y[6].g_x[7].t.w_si ;
 wire \g.g_y[7].g_x[0].t.out_sc ;
 wire \g.g_y[7].g_x[0].t.r_d ;
 wire \g.g_y[7].g_x[0].t.r_h ;
 wire \g.g_y[7].g_x[0].t.r_v ;
 wire \g.g_y[7].g_x[0].t.w_si ;
 wire \g.g_y[7].g_x[1].t.out_sc ;
 wire \g.g_y[7].g_x[1].t.r_d ;
 wire \g.g_y[7].g_x[1].t.r_ghl ;
 wire \g.g_y[7].g_x[1].t.r_gnl ;
 wire \g.g_y[7].g_x[1].t.r_h ;
 wire \g.g_y[7].g_x[1].t.r_v ;
 wire \g.g_y[7].g_x[1].t.w_dh ;
 wire \g.g_y[7].g_x[1].t.w_na ;
 wire \g.g_y[7].g_x[1].t.w_si ;
 wire \g.g_y[7].g_x[2].t.out_sc ;
 wire \g.g_y[7].g_x[2].t.r_d ;
 wire \g.g_y[7].g_x[2].t.r_h ;
 wire \g.g_y[7].g_x[2].t.r_v ;
 wire \g.g_y[7].g_x[2].t.w_si ;
 wire \g.g_y[7].g_x[3].t.out_sc ;
 wire \g.g_y[7].g_x[3].t.r_d ;
 wire \g.g_y[7].g_x[3].t.r_ghl ;
 wire \g.g_y[7].g_x[3].t.r_gnl ;
 wire \g.g_y[7].g_x[3].t.r_h ;
 wire \g.g_y[7].g_x[3].t.r_v ;
 wire \g.g_y[7].g_x[3].t.w_dh ;
 wire \g.g_y[7].g_x[3].t.w_na ;
 wire \g.g_y[7].g_x[3].t.w_si ;
 wire \g.g_y[7].g_x[4].t.out_sc ;
 wire \g.g_y[7].g_x[4].t.r_d ;
 wire \g.g_y[7].g_x[4].t.r_h ;
 wire \g.g_y[7].g_x[4].t.r_v ;
 wire \g.g_y[7].g_x[4].t.w_si ;
 wire \g.g_y[7].g_x[5].t.out_sc ;
 wire \g.g_y[7].g_x[5].t.r_d ;
 wire \g.g_y[7].g_x[5].t.r_ghl ;
 wire \g.g_y[7].g_x[5].t.r_gnl ;
 wire \g.g_y[7].g_x[5].t.r_h ;
 wire \g.g_y[7].g_x[5].t.r_v ;
 wire \g.g_y[7].g_x[5].t.w_dh ;
 wire \g.g_y[7].g_x[5].t.w_na ;
 wire \g.g_y[7].g_x[5].t.w_si ;
 wire \g.g_y[7].g_x[6].t.out_sc ;
 wire \g.g_y[7].g_x[6].t.r_d ;
 wire \g.g_y[7].g_x[6].t.r_h ;
 wire \g.g_y[7].g_x[6].t.r_v ;
 wire \g.g_y[7].g_x[6].t.w_si ;
 wire \g.g_y[7].g_x[7].t.out_r ;
 wire \g.g_y[7].g_x[7].t.out_sc ;
 wire \g.g_y[7].g_x[7].t.r_d ;
 wire \g.g_y[7].g_x[7].t.r_ghl ;
 wire \g.g_y[7].g_x[7].t.r_gnl ;
 wire \g.g_y[7].g_x[7].t.r_h ;
 wire \g.g_y[7].g_x[7].t.r_v ;
 wire \g.g_y[7].g_x[7].t.w_dh ;
 wire \g.g_y[7].g_x[7].t.w_na ;
 wire \g.g_y[7].g_x[7].t.w_si ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _2346_ (.A(rst_n),
    .X(_1777_));
 sg13g2_inv_1 _2347_ (.Y(_1778_),
    .A(_1777_));
 sg13g2_a21o_1 _2348_ (.A2(net11),
    .A1(net12),
    .B1(_1778_),
    .X(\g.cfg_d ));
 sg13g2_inv_1 _2349_ (.Y(_1779_),
    .A(net12));
 sg13g2_o21ai_1 _2350_ (.B1(_1777_),
    .Y(\g.cfg_h ),
    .A1(_1779_),
    .A2(net11));
 sg13g2_inv_1 _2351_ (.Y(_1780_),
    .A(net15));
 sg13g2_inv_1 _2352_ (.Y(_1781_),
    .A(net14));
 sg13g2_nand3_1 _2353_ (.B(_1780_),
    .C(_1781_),
    .A(_1777_),
    .Y(\g.g_y[0].g_x[0].t.in_lb ));
 sg13g2_a21o_1 _2354_ (.A2(net11),
    .A1(_1779_),
    .B1(_1778_),
    .X(\g.cfg_v ));
 sg13g2_buf_1 _2355_ (.A(\g.g_y[0].g_x[1].t.r_d ),
    .X(_1782_));
 sg13g2_buf_1 _2356_ (.A(\g.g_y[0].g_x[2].t.r_ghl ),
    .X(_1783_));
 sg13g2_buf_2 _2357_ (.A(\g.g_y[0].g_x[2].t.r_d ),
    .X(_1784_));
 sg13g2_mux2_1 _2358_ (.A0(\g.g_y[0].g_x[2].t.out_sc ),
    .A1(\g.g_y[0].g_x[2].t.r_gnl ),
    .S(_1784_),
    .X(_1785_));
 sg13g2_inv_1 _2359_ (.Y(_1786_),
    .A(\g.g_y[0].g_x[2].t.r_h ));
 sg13g2_mux2_1 _2360_ (.A0(_1783_),
    .A1(_1785_),
    .S(_1786_),
    .X(_1787_));
 sg13g2_buf_1 _2361_ (.A(\g.g_y[0].g_x[0].t.r_ghl ),
    .X(_1788_));
 sg13g2_buf_2 _2362_ (.A(\g.g_y[0].g_x[0].t.r_d ),
    .X(_1789_));
 sg13g2_mux2_1 _2363_ (.A0(\g.g_y[0].g_x[0].t.out_sc ),
    .A1(\g.g_y[0].g_x[0].t.r_gnl ),
    .S(_1789_),
    .X(_1790_));
 sg13g2_buf_2 _2364_ (.A(\g.g_y[0].g_x[0].t.r_h ),
    .X(_1791_));
 sg13g2_mux2_1 _2365_ (.A0(_1788_),
    .A1(_1790_),
    .S(_1791_),
    .X(_1792_));
 sg13g2_buf_1 _2366_ (.A(\g.g_y[0].g_x[1].t.r_h ),
    .X(_1793_));
 sg13g2_mux2_1 _2367_ (.A0(_1787_),
    .A1(_1792_),
    .S(net83),
    .X(_1794_));
 sg13g2_buf_1 _2368_ (.A(\g.g_y[7].g_x[1].t.r_ghl ),
    .X(_1795_));
 sg13g2_buf_2 _2369_ (.A(\g.g_y[7].g_x[1].t.r_d ),
    .X(_1796_));
 sg13g2_mux2_1 _2370_ (.A0(\g.g_y[7].g_x[1].t.r_gnl ),
    .A1(\g.g_y[7].g_x[1].t.out_sc ),
    .S(_1796_),
    .X(_1797_));
 sg13g2_buf_1 _2371_ (.A(_1797_),
    .X(_1798_));
 sg13g2_buf_2 _2372_ (.A(\g.g_y[7].g_x[1].t.r_v ),
    .X(_1799_));
 sg13g2_mux2_1 _2373_ (.A0(_1795_),
    .A1(_1798_),
    .S(_1799_),
    .X(_1800_));
 sg13g2_buf_1 _2374_ (.A(\g.g_y[1].g_x[1].t.r_ghl ),
    .X(_1801_));
 sg13g2_buf_2 _2375_ (.A(\g.g_y[1].g_x[1].t.r_d ),
    .X(_1802_));
 sg13g2_mux2_1 _2376_ (.A0(\g.g_y[1].g_x[1].t.r_gnl ),
    .A1(\g.g_y[1].g_x[1].t.out_sc ),
    .S(_1802_),
    .X(_1803_));
 sg13g2_inv_1 _2377_ (.Y(_1804_),
    .A(\g.g_y[1].g_x[1].t.r_v ));
 sg13g2_mux2_1 _2378_ (.A0(_1801_),
    .A1(_1803_),
    .S(_1804_),
    .X(_1805_));
 sg13g2_buf_1 _2379_ (.A(\g.g_y[0].g_x[1].t.r_v ),
    .X(_1806_));
 sg13g2_inv_1 _2380_ (.Y(_1807_),
    .A(_1806_));
 sg13g2_mux2_1 _2381_ (.A0(_1800_),
    .A1(_1805_),
    .S(_1807_),
    .X(_1808_));
 sg13g2_nand3_1 _2382_ (.B(_1794_),
    .C(_1808_),
    .A(net66),
    .Y(_1809_));
 sg13g2_nor2_1 _2383_ (.A(\g.g_y[0].g_x[1].t.out_sc ),
    .B(net66),
    .Y(_1810_));
 sg13g2_nor2_1 _2384_ (.A(net83),
    .B(_1810_),
    .Y(_1811_));
 sg13g2_mux2_1 _2385_ (.A0(_1792_),
    .A1(_1787_),
    .S(net83),
    .X(_1812_));
 sg13g2_mux2_1 _2386_ (.A0(_1800_),
    .A1(_1805_),
    .S(_1806_),
    .X(_1813_));
 sg13g2_mux2_1 _2387_ (.A0(_1812_),
    .A1(_1813_),
    .S(_1782_),
    .X(_1814_));
 sg13g2_buf_2 _2388_ (.A(_1814_),
    .X(_1815_));
 sg13g2_inv_1 _2389_ (.Y(_1816_),
    .A(_1791_));
 sg13g2_a221oi_1 _2390_ (.B2(net83),
    .C1(_1816_),
    .B1(_1815_),
    .A1(_1809_),
    .Y(_1817_),
    .A2(_1811_));
 sg13g2_nor2_1 _2391_ (.A(_1791_),
    .B(net1),
    .Y(_1818_));
 sg13g2_or2_1 _2392_ (.X(_1819_),
    .B(_1818_),
    .A(_1789_));
 sg13g2_buf_2 _2393_ (.A(\g.g_y[0].g_x[0].t.r_v ),
    .X(_1820_));
 sg13g2_buf_1 _2394_ (.A(\g.g_y[1].g_x[0].t.r_v ),
    .X(_1821_));
 sg13g2_buf_2 _2395_ (.A(\g.g_y[1].g_x[0].t.r_h ),
    .X(_1822_));
 sg13g2_mux2_1 _2396_ (.A0(\g.g_y[1].g_x[1].t.out_sc ),
    .A1(\g.g_y[1].g_x[1].t.r_gnl ),
    .S(_1802_),
    .X(_1823_));
 sg13g2_buf_1 _2397_ (.A(\g.g_y[1].g_x[1].t.r_h ),
    .X(_1824_));
 sg13g2_inv_1 _2398_ (.Y(_1825_),
    .A(_1824_));
 sg13g2_mux2_1 _2399_ (.A0(_1801_),
    .A1(_1823_),
    .S(_1825_),
    .X(_1826_));
 sg13g2_buf_1 _2400_ (.A(_1826_),
    .X(_1827_));
 sg13g2_buf_1 _2401_ (.A(\g.g_y[1].g_x[0].t.r_d ),
    .X(_1828_));
 sg13g2_nor2b_1 _2402_ (.A(_1822_),
    .B_N(net2),
    .Y(_1829_));
 sg13g2_or2_1 _2403_ (.X(_1830_),
    .B(_1829_),
    .A(_1828_));
 sg13g2_a21o_1 _2404_ (.A2(_1827_),
    .A1(_1822_),
    .B1(_1830_),
    .X(_1831_));
 sg13g2_buf_1 _2405_ (.A(_1828_),
    .X(_1832_));
 sg13g2_buf_2 _2406_ (.A(\g.g_y[2].g_x[0].t.r_v ),
    .X(_1833_));
 sg13g2_buf_2 _2407_ (.A(\g.g_y[2].g_x[0].t.r_d ),
    .X(_1834_));
 sg13g2_mux2_1 _2408_ (.A0(\g.g_y[2].g_x[0].t.r_gnl ),
    .A1(\g.g_y[2].g_x[0].t.out_sc ),
    .S(_1834_),
    .X(_1835_));
 sg13g2_buf_1 _2409_ (.A(\g.g_y[2].g_x[0].t.r_ghl ),
    .X(_1836_));
 sg13g2_nand2b_1 _2410_ (.Y(_1837_),
    .B(_1833_),
    .A_N(_1836_));
 sg13g2_o21ai_1 _2411_ (.B1(_1837_),
    .Y(_1838_),
    .A1(_1833_),
    .A2(_1835_));
 sg13g2_nand2_1 _2412_ (.Y(_1839_),
    .A(_1832_),
    .B(_1838_));
 sg13g2_nand3_1 _2413_ (.B(_1831_),
    .C(_1839_),
    .A(_1821_),
    .Y(_1840_));
 sg13g2_nand2b_1 _2414_ (.Y(_1841_),
    .B(_1825_),
    .A_N(_1823_));
 sg13g2_nor2b_1 _2415_ (.A(_1801_),
    .B_N(_1824_),
    .Y(_1842_));
 sg13g2_nor3_1 _2416_ (.A(_1822_),
    .B(_1828_),
    .C(_1842_),
    .Y(_1843_));
 sg13g2_inv_1 _2417_ (.Y(_1844_),
    .A(net2));
 sg13g2_inv_1 _2418_ (.Y(_1845_),
    .A(_1822_));
 sg13g2_nor3_1 _2419_ (.A(_1844_),
    .B(_1845_),
    .C(_1828_),
    .Y(_1846_));
 sg13g2_a21oi_1 _2420_ (.A1(_1841_),
    .A2(_1843_),
    .Y(_1847_),
    .B1(_1846_));
 sg13g2_nand2b_1 _2421_ (.Y(_1848_),
    .B(_1828_),
    .A_N(\g.g_y[1].g_x[0].t.out_sc ));
 sg13g2_nor2b_1 _2422_ (.A(_1821_),
    .B_N(_1848_),
    .Y(_1849_));
 sg13g2_o21ai_1 _2423_ (.B1(_1849_),
    .Y(_1850_),
    .A1(_1838_),
    .A2(_1847_));
 sg13g2_nand3_1 _2424_ (.B(_1840_),
    .C(_1850_),
    .A(_1820_),
    .Y(_1851_));
 sg13g2_inv_1 _2425_ (.Y(_1852_),
    .A(_1820_));
 sg13g2_buf_1 _2426_ (.A(\g.g_y[7].g_x[0].t.r_v ),
    .X(_1853_));
 sg13g2_inv_1 _2427_ (.Y(_1854_),
    .A(_1853_));
 sg13g2_buf_1 _2428_ (.A(\g.g_y[7].g_x[0].t.r_h ),
    .X(_1855_));
 sg13g2_inv_1 _2429_ (.Y(_1856_),
    .A(_1855_));
 sg13g2_buf_1 _2430_ (.A(\g.g_y[7].g_x[1].t.r_h ),
    .X(_1857_));
 sg13g2_mux2_1 _2431_ (.A0(\g.g_y[7].g_x[1].t.out_sc ),
    .A1(\g.g_y[7].g_x[1].t.r_gnl ),
    .S(_1796_),
    .X(_1858_));
 sg13g2_nand2b_1 _2432_ (.Y(_1859_),
    .B(_1857_),
    .A_N(_1795_));
 sg13g2_o21ai_1 _2433_ (.B1(_1859_),
    .Y(_1860_),
    .A1(_1857_),
    .A2(_1858_));
 sg13g2_buf_1 _2434_ (.A(_1860_),
    .X(_1861_));
 sg13g2_buf_1 _2435_ (.A(\g.g_y[7].g_x[0].t.r_d ),
    .X(_1862_));
 sg13g2_nor2b_1 _2436_ (.A(_1855_),
    .B_N(net8),
    .Y(_1863_));
 sg13g2_nor2_1 _2437_ (.A(net65),
    .B(_1863_),
    .Y(_1864_));
 sg13g2_o21ai_1 _2438_ (.B1(_1864_),
    .Y(_1865_),
    .A1(_1856_),
    .A2(_1861_));
 sg13g2_inv_1 _2439_ (.Y(_1866_),
    .A(\g.g_y[6].g_x[0].t.r_v ));
 sg13g2_buf_2 _2440_ (.A(\g.g_y[6].g_x[0].t.r_d ),
    .X(_1867_));
 sg13g2_mux2_1 _2441_ (.A0(\g.g_y[6].g_x[0].t.r_gnl ),
    .A1(\g.g_y[6].g_x[0].t.out_sc ),
    .S(_1867_),
    .X(_1868_));
 sg13g2_buf_1 _2442_ (.A(\g.g_y[6].g_x[0].t.r_ghl ),
    .X(_1869_));
 sg13g2_or2_1 _2443_ (.X(_1870_),
    .B(\g.g_y[6].g_x[0].t.r_v ),
    .A(_1869_));
 sg13g2_o21ai_1 _2444_ (.B1(_1870_),
    .Y(_1871_),
    .A1(_1866_),
    .A2(_1868_));
 sg13g2_buf_1 _2445_ (.A(_1871_),
    .X(_1872_));
 sg13g2_nand2_1 _2446_ (.Y(_1873_),
    .A(_1862_),
    .B(_1872_));
 sg13g2_nand3_1 _2447_ (.B(_1865_),
    .C(_1873_),
    .A(_1854_),
    .Y(_1874_));
 sg13g2_inv_1 _2448_ (.Y(_1875_),
    .A(net65));
 sg13g2_and2_1 _2449_ (.A(net8),
    .B(_1855_),
    .X(_1876_));
 sg13g2_and3_1 _2450_ (.X(_1877_),
    .A(_1856_),
    .B(_1875_),
    .C(_1859_));
 sg13g2_inv_1 _2451_ (.Y(_1878_),
    .A(_1857_));
 sg13g2_nand2b_1 _2452_ (.Y(_1879_),
    .B(_1878_),
    .A_N(_1858_));
 sg13g2_a22oi_1 _2453_ (.Y(_1880_),
    .B1(_1877_),
    .B2(_1879_),
    .A2(_1876_),
    .A1(_1875_));
 sg13g2_nand2b_1 _2454_ (.Y(_1881_),
    .B(net65),
    .A_N(\g.g_y[7].g_x[0].t.out_sc ));
 sg13g2_and2_1 _2455_ (.A(_1853_),
    .B(_1881_),
    .X(_1882_));
 sg13g2_o21ai_1 _2456_ (.B1(_1882_),
    .Y(_1883_),
    .A1(_1872_),
    .A2(_1880_));
 sg13g2_nand3_1 _2457_ (.B(_1874_),
    .C(_1883_),
    .A(_1852_),
    .Y(_1884_));
 sg13g2_nand3_1 _2458_ (.B(_1851_),
    .C(_1884_),
    .A(_1789_),
    .Y(_1885_));
 sg13g2_o21ai_1 _2459_ (.B1(_1885_),
    .Y(\g.g_y[0].g_x[0].t.w_dh ),
    .A1(_1817_),
    .A2(_1819_));
 sg13g2_a21oi_1 _2460_ (.A1(_1874_),
    .A2(_1883_),
    .Y(_1886_),
    .B1(_1852_));
 sg13g2_a21oi_1 _2461_ (.A1(_1840_),
    .A2(_1850_),
    .Y(_1887_),
    .B1(_1820_));
 sg13g2_a22oi_1 _2462_ (.Y(_1888_),
    .B1(_1815_),
    .B2(_1793_),
    .A2(_1811_),
    .A1(_1809_));
 sg13g2_nand2_1 _2463_ (.Y(_1889_),
    .A(_1791_),
    .B(net1));
 sg13g2_o21ai_1 _2464_ (.B1(_1889_),
    .Y(_1890_),
    .A1(_1791_),
    .A2(_1888_));
 sg13g2_o21ai_1 _2465_ (.B1(_1890_),
    .Y(\g.g_y[0].g_x[0].t.w_na ),
    .A1(_1886_),
    .A2(_1887_));
 sg13g2_inv_1 _2466_ (.Y(_1891_),
    .A(_1789_));
 sg13g2_nand2b_1 _2467_ (.Y(_1892_),
    .B(_1777_),
    .A_N(net9));
 sg13g2_buf_1 _2468_ (.A(_1892_),
    .X(_1893_));
 sg13g2_buf_1 _2469_ (.A(_1893_),
    .X(_1894_));
 sg13g2_or4_1 _2470_ (.A(_1891_),
    .B(_1817_),
    .C(_1818_),
    .D(net82),
    .X(_1895_));
 sg13g2_nor3_1 _2471_ (.A(_1778_),
    .B(_1789_),
    .C(net9),
    .Y(_1896_));
 sg13g2_nand3_1 _2472_ (.B(_1884_),
    .C(_1896_),
    .A(_1851_),
    .Y(_1897_));
 sg13g2_nand3_1 _2473_ (.B(net9),
    .C(net10),
    .A(_1777_),
    .Y(_1898_));
 sg13g2_nand3_1 _2474_ (.B(_1897_),
    .C(_1898_),
    .A(_1895_),
    .Y(\g.g_y[0].g_x[0].t.w_si ));
 sg13g2_mux2_1 _2475_ (.A0(_1813_),
    .A1(_1812_),
    .S(net66),
    .X(_1899_));
 sg13g2_nor2_2 _2476_ (.A(_1778_),
    .B(net9),
    .Y(_1900_));
 sg13g2_buf_1 _2477_ (.A(_1900_),
    .X(_1901_));
 sg13g2_buf_2 _2478_ (.A(net81),
    .X(_1902_));
 sg13g2_mux2_1 _2479_ (.A0(\g.g_y[0].g_x[0].t.out_sc ),
    .A1(_1899_),
    .S(_1902_),
    .X(\g.g_y[0].g_x[1].t.w_si ));
 sg13g2_nor2_1 _2480_ (.A(_1778_),
    .B(net13),
    .Y(_1903_));
 sg13g2_a21oi_1 _2481_ (.A1(net15),
    .A2(net14),
    .Y(\g.g_y[0].g_x[2].t.in_lb ),
    .B1(_1903_));
 sg13g2_inv_1 _2482_ (.Y(_1904_),
    .A(_1784_));
 sg13g2_buf_1 _2483_ (.A(\g.g_y[1].g_x[2].t.r_d ),
    .X(_1905_));
 sg13g2_buf_2 _2484_ (.A(\g.g_y[1].g_x[3].t.r_d ),
    .X(_1906_));
 sg13g2_mux2_1 _2485_ (.A0(\g.g_y[1].g_x[3].t.out_sc ),
    .A1(\g.g_y[1].g_x[3].t.r_gnl ),
    .S(_1906_),
    .X(_1907_));
 sg13g2_buf_1 _2486_ (.A(_1907_),
    .X(_1908_));
 sg13g2_buf_2 _2487_ (.A(\g.g_y[1].g_x[3].t.r_h ),
    .X(_1909_));
 sg13g2_inv_1 _2488_ (.Y(_1910_),
    .A(_1909_));
 sg13g2_nand2b_1 _2489_ (.Y(_1911_),
    .B(_1910_),
    .A_N(_1908_));
 sg13g2_buf_2 _2490_ (.A(\g.g_y[1].g_x[3].t.r_ghl ),
    .X(_1912_));
 sg13g2_inv_1 _2491_ (.Y(_1913_),
    .A(_1912_));
 sg13g2_buf_1 _2492_ (.A(\g.g_y[1].g_x[2].t.r_h ),
    .X(_1914_));
 sg13g2_a21oi_1 _2493_ (.A1(_1913_),
    .A2(_1909_),
    .Y(_1915_),
    .B1(_1914_));
 sg13g2_mux2_1 _2494_ (.A0(_1801_),
    .A1(_1823_),
    .S(_1824_),
    .X(_1916_));
 sg13g2_a22oi_1 _2495_ (.Y(_1917_),
    .B1(_1916_),
    .B2(_1914_),
    .A2(_1915_),
    .A1(_1911_));
 sg13g2_buf_2 _2496_ (.A(\g.g_y[2].g_x[2].t.r_d ),
    .X(_1918_));
 sg13g2_mux2_1 _2497_ (.A0(\g.g_y[2].g_x[2].t.r_gnl ),
    .A1(\g.g_y[2].g_x[2].t.out_sc ),
    .S(_1918_),
    .X(_1919_));
 sg13g2_buf_1 _2498_ (.A(\g.g_y[2].g_x[2].t.r_v ),
    .X(_1920_));
 sg13g2_inv_1 _2499_ (.Y(_1921_),
    .A(_1920_));
 sg13g2_nand2b_1 _2500_ (.Y(_1922_),
    .B(_1921_),
    .A_N(_1919_));
 sg13g2_buf_1 _2501_ (.A(\g.g_y[2].g_x[2].t.r_ghl ),
    .X(_1923_));
 sg13g2_inv_1 _2502_ (.Y(_1924_),
    .A(_1923_));
 sg13g2_buf_1 _2503_ (.A(\g.g_y[1].g_x[2].t.r_v ),
    .X(_1925_));
 sg13g2_a21oi_1 _2504_ (.A1(_1924_),
    .A2(_1920_),
    .Y(_1926_),
    .B1(_1925_));
 sg13g2_mux2_1 _2505_ (.A0(\g.g_y[0].g_x[2].t.r_gnl ),
    .A1(\g.g_y[0].g_x[2].t.out_sc ),
    .S(_1784_),
    .X(_1927_));
 sg13g2_buf_1 _2506_ (.A(_1927_),
    .X(_1928_));
 sg13g2_buf_2 _2507_ (.A(\g.g_y[0].g_x[2].t.r_v ),
    .X(_1929_));
 sg13g2_mux2_1 _2508_ (.A0(_1783_),
    .A1(_1928_),
    .S(_1929_),
    .X(_1930_));
 sg13g2_a22oi_1 _2509_ (.Y(_1931_),
    .B1(_1930_),
    .B2(_1925_),
    .A2(_1926_),
    .A1(_1922_));
 sg13g2_or3_1 _2510_ (.A(_1905_),
    .B(_1917_),
    .C(_1931_),
    .X(_1932_));
 sg13g2_buf_1 _2511_ (.A(_1932_),
    .X(_1933_));
 sg13g2_inv_1 _2512_ (.Y(_1934_),
    .A(\g.g_y[1].g_x[2].t.out_sc ));
 sg13g2_a21oi_1 _2513_ (.A1(net63),
    .A2(_1934_),
    .Y(_1935_),
    .B1(_1925_));
 sg13g2_mux2_1 _2514_ (.A0(_1912_),
    .A1(_1908_),
    .S(_1910_),
    .X(_1936_));
 sg13g2_inv_1 _2515_ (.Y(_1937_),
    .A(_1914_));
 sg13g2_mux2_1 _2516_ (.A0(_1936_),
    .A1(_1916_),
    .S(_1937_),
    .X(_1938_));
 sg13g2_mux2_1 _2517_ (.A0(_1923_),
    .A1(_1919_),
    .S(_1921_),
    .X(_1939_));
 sg13g2_inv_1 _2518_ (.Y(_1940_),
    .A(_1925_));
 sg13g2_mux2_1 _2519_ (.A0(_1939_),
    .A1(_1930_),
    .S(_1940_),
    .X(_1941_));
 sg13g2_buf_1 _2520_ (.A(_1941_),
    .X(_1942_));
 sg13g2_mux2_1 _2521_ (.A0(_1938_),
    .A1(_1942_),
    .S(\g.g_y[1].g_x[2].t.r_d ),
    .X(_1943_));
 sg13g2_buf_1 _2522_ (.A(_1943_),
    .X(_1944_));
 sg13g2_inv_1 _2523_ (.Y(_1945_),
    .A(_1929_));
 sg13g2_a221oi_1 _2524_ (.B2(_1925_),
    .C1(_1945_),
    .B1(_1944_),
    .A1(_1933_),
    .Y(_1946_),
    .A2(_1935_));
 sg13g2_buf_2 _2525_ (.A(\g.g_y[7].g_x[2].t.r_v ),
    .X(_1947_));
 sg13g2_inv_1 _2526_ (.Y(_1948_),
    .A(_1947_));
 sg13g2_buf_1 _2527_ (.A(\g.g_y[6].g_x[2].t.r_ghl ),
    .X(_1949_));
 sg13g2_buf_2 _2528_ (.A(\g.g_y[6].g_x[2].t.r_d ),
    .X(_1950_));
 sg13g2_mux2_1 _2529_ (.A0(\g.g_y[6].g_x[2].t.r_gnl ),
    .A1(\g.g_y[6].g_x[2].t.out_sc ),
    .S(_1950_),
    .X(_1951_));
 sg13g2_buf_2 _2530_ (.A(\g.g_y[6].g_x[2].t.r_v ),
    .X(_1952_));
 sg13g2_mux2_1 _2531_ (.A0(_1949_),
    .A1(_1951_),
    .S(_1952_),
    .X(_1953_));
 sg13g2_mux2_1 _2532_ (.A0(_1783_),
    .A1(_1928_),
    .S(_1945_),
    .X(_1954_));
 sg13g2_mux2_1 _2533_ (.A0(_1953_),
    .A1(_1954_),
    .S(_1947_),
    .X(_1955_));
 sg13g2_buf_1 _2534_ (.A(_1955_),
    .X(_1956_));
 sg13g2_mux2_1 _2535_ (.A0(_1795_),
    .A1(_1858_),
    .S(_1857_),
    .X(_1957_));
 sg13g2_buf_2 _2536_ (.A(\g.g_y[7].g_x[3].t.r_ghl ),
    .X(_1958_));
 sg13g2_buf_2 _2537_ (.A(\g.g_y[7].g_x[3].t.r_d ),
    .X(_1959_));
 sg13g2_mux2_1 _2538_ (.A0(\g.g_y[7].g_x[3].t.out_sc ),
    .A1(\g.g_y[7].g_x[3].t.r_gnl ),
    .S(_1959_),
    .X(_1960_));
 sg13g2_buf_2 _2539_ (.A(\g.g_y[7].g_x[3].t.r_h ),
    .X(_1961_));
 sg13g2_inv_1 _2540_ (.Y(_1962_),
    .A(_1961_));
 sg13g2_mux2_1 _2541_ (.A0(_1958_),
    .A1(_1960_),
    .S(_1962_),
    .X(_1963_));
 sg13g2_buf_1 _2542_ (.A(\g.g_y[7].g_x[2].t.r_h ),
    .X(_1964_));
 sg13g2_mux2_1 _2543_ (.A0(_1957_),
    .A1(_1963_),
    .S(_1964_),
    .X(_1965_));
 sg13g2_buf_2 _2544_ (.A(\g.g_y[7].g_x[2].t.r_d ),
    .X(_1966_));
 sg13g2_inv_1 _2545_ (.Y(_1967_),
    .A(_1966_));
 sg13g2_mux2_1 _2546_ (.A0(_1956_),
    .A1(_1965_),
    .S(_1967_),
    .X(_1968_));
 sg13g2_nand2b_1 _2547_ (.Y(_1969_),
    .B(_1962_),
    .A_N(_1960_));
 sg13g2_inv_1 _2548_ (.Y(_1970_),
    .A(_1958_));
 sg13g2_a21oi_1 _2549_ (.A1(_1970_),
    .A2(_1961_),
    .Y(_1971_),
    .B1(_1964_));
 sg13g2_a22oi_1 _2550_ (.Y(_1972_),
    .B1(_1969_),
    .B2(_1971_),
    .A2(_1957_),
    .A1(_1964_));
 sg13g2_buf_1 _2551_ (.A(_1972_),
    .X(_1973_));
 sg13g2_nand2b_1 _2552_ (.Y(_1974_),
    .B(_1945_),
    .A_N(_1928_));
 sg13g2_nand2b_1 _2553_ (.Y(_1975_),
    .B(_1929_),
    .A_N(_1783_));
 sg13g2_and2_1 _2554_ (.A(_1948_),
    .B(_1975_),
    .X(_1976_));
 sg13g2_a22oi_1 _2555_ (.Y(_1977_),
    .B1(_1974_),
    .B2(_1976_),
    .A2(_1953_),
    .A1(_1947_));
 sg13g2_or3_1 _2556_ (.A(_1966_),
    .B(_1973_),
    .C(_1977_),
    .X(_1978_));
 sg13g2_nand2b_1 _2557_ (.Y(_1979_),
    .B(_1966_),
    .A_N(\g.g_y[7].g_x[2].t.out_sc ));
 sg13g2_and2_1 _2558_ (.A(_1947_),
    .B(_1979_),
    .X(_1980_));
 sg13g2_a221oi_1 _2559_ (.B2(_1980_),
    .C1(_1929_),
    .B1(_1978_),
    .A1(_1948_),
    .Y(_1981_),
    .A2(_1968_));
 sg13g2_nor3_1 _2560_ (.A(_1904_),
    .B(_1946_),
    .C(_1981_),
    .Y(_1982_));
 sg13g2_buf_2 _2561_ (.A(\g.g_y[0].g_x[3].t.r_h ),
    .X(_1983_));
 sg13g2_mux2_1 _2562_ (.A0(_1783_),
    .A1(_1785_),
    .S(\g.g_y[0].g_x[2].t.r_h ),
    .X(_1984_));
 sg13g2_buf_2 _2563_ (.A(\g.g_y[0].g_x[4].t.r_d ),
    .X(_1985_));
 sg13g2_mux2_1 _2564_ (.A0(\g.g_y[0].g_x[4].t.out_sc ),
    .A1(\g.g_y[0].g_x[4].t.r_gnl ),
    .S(_1985_),
    .X(_1986_));
 sg13g2_buf_1 _2565_ (.A(_1986_),
    .X(_1987_));
 sg13g2_buf_2 _2566_ (.A(\g.g_y[0].g_x[4].t.r_h ),
    .X(_1988_));
 sg13g2_inv_1 _2567_ (.Y(_1989_),
    .A(_1988_));
 sg13g2_nand2b_1 _2568_ (.Y(_1990_),
    .B(_1989_),
    .A_N(_1987_));
 sg13g2_buf_2 _2569_ (.A(\g.g_y[0].g_x[4].t.r_ghl ),
    .X(_1991_));
 sg13g2_inv_1 _2570_ (.Y(_1992_),
    .A(_1991_));
 sg13g2_a21oi_1 _2571_ (.A1(_1992_),
    .A2(_1988_),
    .Y(_1993_),
    .B1(_1983_));
 sg13g2_a22oi_1 _2572_ (.Y(_1994_),
    .B1(_1990_),
    .B2(_1993_),
    .A2(_1984_),
    .A1(_1983_));
 sg13g2_buf_2 _2573_ (.A(\g.g_y[0].g_x[3].t.r_v ),
    .X(_1995_));
 sg13g2_mux2_1 _2574_ (.A0(\g.g_y[7].g_x[3].t.r_gnl ),
    .A1(\g.g_y[7].g_x[3].t.out_sc ),
    .S(_1959_),
    .X(_1996_));
 sg13g2_buf_2 _2575_ (.A(\g.g_y[7].g_x[3].t.r_v ),
    .X(_1997_));
 sg13g2_mux2_1 _2576_ (.A0(_1958_),
    .A1(_1996_),
    .S(_1997_),
    .X(_1998_));
 sg13g2_mux2_1 _2577_ (.A0(\g.g_y[1].g_x[3].t.r_gnl ),
    .A1(\g.g_y[1].g_x[3].t.out_sc ),
    .S(_1906_),
    .X(_1999_));
 sg13g2_buf_1 _2578_ (.A(_1999_),
    .X(_2000_));
 sg13g2_buf_2 _2579_ (.A(\g.g_y[1].g_x[3].t.r_v ),
    .X(_2001_));
 sg13g2_inv_1 _2580_ (.Y(_2002_),
    .A(_2001_));
 sg13g2_nand2b_1 _2581_ (.Y(_2003_),
    .B(_2002_),
    .A_N(_2000_));
 sg13g2_a21oi_1 _2582_ (.A1(_1913_),
    .A2(_2001_),
    .Y(_2004_),
    .B1(_1995_));
 sg13g2_a22oi_1 _2583_ (.Y(_2005_),
    .B1(_2003_),
    .B2(_2004_),
    .A2(_1998_),
    .A1(_1995_));
 sg13g2_buf_1 _2584_ (.A(\g.g_y[0].g_x[3].t.r_d ),
    .X(_2006_));
 sg13g2_nor2b_1 _2585_ (.A(_1983_),
    .B_N(net62),
    .Y(_2007_));
 sg13g2_o21ai_1 _2586_ (.B1(_2007_),
    .Y(_2008_),
    .A1(_1994_),
    .A2(_2005_));
 sg13g2_mux2_1 _2587_ (.A0(_1912_),
    .A1(_2000_),
    .S(_2002_),
    .X(_2009_));
 sg13g2_mux2_1 _2588_ (.A0(_1998_),
    .A1(_2009_),
    .S(_1995_),
    .X(_2010_));
 sg13g2_buf_1 _2589_ (.A(_2010_),
    .X(_2011_));
 sg13g2_and2_1 _2590_ (.A(_1983_),
    .B(net62),
    .X(_2012_));
 sg13g2_nand2_1 _2591_ (.Y(_2013_),
    .A(_2011_),
    .B(_2012_));
 sg13g2_mux2_1 _2592_ (.A0(_1991_),
    .A1(_1987_),
    .S(_1989_),
    .X(_2014_));
 sg13g2_nor2b_1 _2593_ (.A(_2006_),
    .B_N(_1983_),
    .Y(_2015_));
 sg13g2_nor2_1 _2594_ (.A(_1983_),
    .B(net62),
    .Y(_2016_));
 sg13g2_a22oi_1 _2595_ (.Y(_2017_),
    .B1(_2016_),
    .B2(\g.g_y[0].g_x[3].t.out_sc ),
    .A2(_2015_),
    .A1(_2014_));
 sg13g2_nand4_1 _2596_ (.B(_2008_),
    .C(_2013_),
    .A(\g.g_y[0].g_x[2].t.r_h ),
    .Y(_2018_),
    .D(_2017_));
 sg13g2_nand2_1 _2597_ (.Y(_2019_),
    .A(net83),
    .B(net66));
 sg13g2_a21o_1 _2598_ (.A2(_1808_),
    .A1(_1794_),
    .B1(_2019_),
    .X(_2020_));
 sg13g2_nor2b_1 _2599_ (.A(net83),
    .B_N(net66),
    .Y(_2021_));
 sg13g2_nor2_1 _2600_ (.A(net83),
    .B(net66),
    .Y(_2022_));
 sg13g2_nand2_1 _2601_ (.Y(_2023_),
    .A(net83),
    .B(\g.g_y[0].g_x[1].t.out_sc ));
 sg13g2_nor2_1 _2602_ (.A(_1782_),
    .B(_2023_),
    .Y(_2024_));
 sg13g2_a221oi_1 _2603_ (.B2(_1792_),
    .C1(_2024_),
    .B1(_2022_),
    .A1(_1813_),
    .Y(_2025_),
    .A2(_2021_));
 sg13g2_nand3_1 _2604_ (.B(_2020_),
    .C(_2025_),
    .A(_1786_),
    .Y(_2026_));
 sg13g2_nand3_1 _2605_ (.B(_2018_),
    .C(_2026_),
    .A(_1904_),
    .Y(_2027_));
 sg13g2_nand2b_1 _2606_ (.Y(\g.g_y[0].g_x[2].t.w_dh ),
    .B(_2027_),
    .A_N(_1982_));
 sg13g2_nand3_1 _2607_ (.B(_2013_),
    .C(_2017_),
    .A(_2008_),
    .Y(_2028_));
 sg13g2_a21oi_1 _2608_ (.A1(_2020_),
    .A2(_2025_),
    .Y(_2029_),
    .B1(_1786_));
 sg13g2_a21o_1 _2609_ (.A2(_2028_),
    .A1(_1786_),
    .B1(_2029_),
    .X(_2030_));
 sg13g2_a22oi_1 _2610_ (.Y(_2031_),
    .B1(_1978_),
    .B2(_1980_),
    .A2(_1968_),
    .A1(_1948_));
 sg13g2_a221oi_1 _2611_ (.B2(_1925_),
    .C1(_1929_),
    .B1(_1944_),
    .A1(_1933_),
    .Y(_2032_),
    .A2(_1935_));
 sg13g2_a21oi_1 _2612_ (.A1(_1929_),
    .A2(_2031_),
    .Y(_2033_),
    .B1(_2032_));
 sg13g2_nand2_1 _2613_ (.Y(\g.g_y[0].g_x[2].t.w_na ),
    .A(_2030_),
    .B(_2033_));
 sg13g2_buf_1 _2614_ (.A(_1893_),
    .X(_2034_));
 sg13g2_or4_1 _2615_ (.A(_1784_),
    .B(net78),
    .C(_1946_),
    .D(_1981_),
    .X(_2035_));
 sg13g2_nand4_1 _2616_ (.B(net64),
    .C(_2018_),
    .A(_1784_),
    .Y(_2036_),
    .D(_2026_));
 sg13g2_buf_1 _2617_ (.A(_1893_),
    .X(_2037_));
 sg13g2_buf_1 _2618_ (.A(net77),
    .X(_2038_));
 sg13g2_nand2_1 _2619_ (.Y(_2039_),
    .A(\g.g_y[0].g_x[1].t.out_sc ),
    .B(net61));
 sg13g2_nand3_1 _2620_ (.B(_2036_),
    .C(_2039_),
    .A(_2035_),
    .Y(\g.g_y[0].g_x[2].t.w_si ));
 sg13g2_buf_1 _2621_ (.A(net82),
    .X(_2040_));
 sg13g2_mux2_1 _2622_ (.A0(_1984_),
    .A1(_2014_),
    .S(_1983_),
    .X(_2041_));
 sg13g2_nor2b_1 _2623_ (.A(net62),
    .B_N(_2011_),
    .Y(_2042_));
 sg13g2_a21oi_1 _2624_ (.A1(net62),
    .A2(_2041_),
    .Y(_2043_),
    .B1(_2042_));
 sg13g2_buf_1 _2625_ (.A(net77),
    .X(_2044_));
 sg13g2_nand2_1 _2626_ (.Y(_2045_),
    .A(\g.g_y[0].g_x[2].t.out_sc ),
    .B(net59));
 sg13g2_o21ai_1 _2627_ (.B1(_2045_),
    .Y(\g.g_y[0].g_x[3].t.w_si ),
    .A1(net60),
    .A2(_2043_));
 sg13g2_inv_1 _2628_ (.Y(_2046_),
    .A(_1985_));
 sg13g2_buf_1 _2629_ (.A(\g.g_y[1].g_x[4].t.r_d ),
    .X(_2047_));
 sg13g2_inv_1 _2630_ (.Y(_2048_),
    .A(\g.g_y[1].g_x[4].t.r_h ));
 sg13g2_buf_8 _2631_ (.A(\g.g_y[1].g_x[5].t.r_d ),
    .X(_2049_));
 sg13g2_mux2_1 _2632_ (.A0(\g.g_y[1].g_x[5].t.out_sc ),
    .A1(\g.g_y[1].g_x[5].t.r_gnl ),
    .S(_2049_),
    .X(_2050_));
 sg13g2_inv_1 _2633_ (.Y(_2051_),
    .A(\g.g_y[1].g_x[5].t.r_h ));
 sg13g2_mux2_1 _2634_ (.A0(\g.g_y[1].g_x[5].t.r_ghl ),
    .A1(_2050_),
    .S(_2051_),
    .X(_2052_));
 sg13g2_or2_1 _2635_ (.X(_2053_),
    .B(_1908_),
    .A(_1910_));
 sg13g2_a21oi_1 _2636_ (.A1(_1913_),
    .A2(_1910_),
    .Y(_2054_),
    .B1(_2048_));
 sg13g2_a22oi_1 _2637_ (.Y(_2055_),
    .B1(_2053_),
    .B2(_2054_),
    .A2(_2052_),
    .A1(_2048_));
 sg13g2_buf_1 _2638_ (.A(_2055_),
    .X(_2056_));
 sg13g2_buf_1 _2639_ (.A(\g.g_y[1].g_x[4].t.r_v ),
    .X(_2057_));
 sg13g2_mux2_1 _2640_ (.A0(\g.g_y[0].g_x[4].t.r_gnl ),
    .A1(\g.g_y[0].g_x[4].t.out_sc ),
    .S(_1985_),
    .X(_2058_));
 sg13g2_buf_2 _2641_ (.A(\g.g_y[0].g_x[4].t.r_v ),
    .X(_2059_));
 sg13g2_mux2_1 _2642_ (.A0(_1991_),
    .A1(_2058_),
    .S(_2059_),
    .X(_2060_));
 sg13g2_buf_8 _2643_ (.A(\g.g_y[2].g_x[4].t.r_d ),
    .X(_2061_));
 sg13g2_mux2_1 _2644_ (.A0(\g.g_y[2].g_x[4].t.r_gnl ),
    .A1(\g.g_y[2].g_x[4].t.out_sc ),
    .S(_2061_),
    .X(_2062_));
 sg13g2_buf_1 _2645_ (.A(\g.g_y[2].g_x[4].t.r_v ),
    .X(_2063_));
 sg13g2_inv_1 _2646_ (.Y(_2064_),
    .A(net56));
 sg13g2_nand2b_1 _2647_ (.Y(_2065_),
    .B(_2064_),
    .A_N(_2062_));
 sg13g2_buf_1 _2648_ (.A(\g.g_y[2].g_x[4].t.r_ghl ),
    .X(_2066_));
 sg13g2_inv_1 _2649_ (.Y(_2067_),
    .A(_2066_));
 sg13g2_a21oi_1 _2650_ (.A1(_2067_),
    .A2(net56),
    .Y(_2068_),
    .B1(net57));
 sg13g2_a22oi_1 _2651_ (.Y(_2069_),
    .B1(_2065_),
    .B2(_2068_),
    .A2(_2060_),
    .A1(net57));
 sg13g2_buf_1 _2652_ (.A(_2069_),
    .X(_2070_));
 sg13g2_or3_1 _2653_ (.A(net58),
    .B(_2056_),
    .C(_2070_),
    .X(_2071_));
 sg13g2_buf_1 _2654_ (.A(_2071_),
    .X(_2072_));
 sg13g2_nand2b_1 _2655_ (.Y(_2073_),
    .B(net58),
    .A_N(\g.g_y[1].g_x[4].t.out_sc ));
 sg13g2_nor2b_1 _2656_ (.A(_2057_),
    .B_N(_2073_),
    .Y(_2074_));
 sg13g2_mux2_1 _2657_ (.A0(_1912_),
    .A1(_1908_),
    .S(_1909_),
    .X(_2075_));
 sg13g2_mux2_1 _2658_ (.A0(_2052_),
    .A1(_2075_),
    .S(_2048_),
    .X(_2076_));
 sg13g2_mux2_1 _2659_ (.A0(_2066_),
    .A1(_2062_),
    .S(_2064_),
    .X(_2077_));
 sg13g2_mux2_1 _2660_ (.A0(_2060_),
    .A1(_2077_),
    .S(net57),
    .X(_2078_));
 sg13g2_buf_1 _2661_ (.A(_2078_),
    .X(_2079_));
 sg13g2_mux2_1 _2662_ (.A0(_2076_),
    .A1(_2079_),
    .S(_2047_),
    .X(_2080_));
 sg13g2_buf_1 _2663_ (.A(_2080_),
    .X(_2081_));
 sg13g2_inv_1 _2664_ (.Y(_2082_),
    .A(_2059_));
 sg13g2_a221oi_1 _2665_ (.B2(_2057_),
    .C1(_2082_),
    .B1(_2081_),
    .A1(_2072_),
    .Y(_2083_),
    .A2(_2074_));
 sg13g2_buf_1 _2666_ (.A(\g.g_y[7].g_x[4].t.r_d ),
    .X(_2084_));
 sg13g2_buf_1 _2667_ (.A(\g.g_y[7].g_x[5].t.r_d ),
    .X(_2085_));
 sg13g2_mux2_1 _2668_ (.A0(\g.g_y[7].g_x[5].t.out_sc ),
    .A1(\g.g_y[7].g_x[5].t.r_gnl ),
    .S(_2085_),
    .X(_2086_));
 sg13g2_buf_1 _2669_ (.A(_2086_),
    .X(_2087_));
 sg13g2_buf_2 _2670_ (.A(\g.g_y[7].g_x[5].t.r_h ),
    .X(_2088_));
 sg13g2_inv_2 _2671_ (.Y(_2089_),
    .A(_2088_));
 sg13g2_nand2b_1 _2672_ (.Y(_2090_),
    .B(_2089_),
    .A_N(_2087_));
 sg13g2_buf_2 _2673_ (.A(\g.g_y[7].g_x[4].t.r_h ),
    .X(_2091_));
 sg13g2_inv_2 _2674_ (.Y(_2092_),
    .A(_2091_));
 sg13g2_buf_1 _2675_ (.A(\g.g_y[7].g_x[5].t.r_ghl ),
    .X(_2093_));
 sg13g2_nand2b_1 _2676_ (.Y(_2094_),
    .B(_2088_),
    .A_N(_2093_));
 sg13g2_and2_1 _2677_ (.A(_2092_),
    .B(_2094_),
    .X(_2095_));
 sg13g2_mux2_1 _2678_ (.A0(_1958_),
    .A1(_1960_),
    .S(_1961_),
    .X(_2096_));
 sg13g2_a22oi_1 _2679_ (.Y(_2097_),
    .B1(_2096_),
    .B2(_2091_),
    .A2(_2095_),
    .A1(_2090_));
 sg13g2_buf_1 _2680_ (.A(_2097_),
    .X(_2098_));
 sg13g2_nand2b_1 _2681_ (.Y(_2099_),
    .B(_2082_),
    .A_N(_2058_));
 sg13g2_buf_2 _2682_ (.A(\g.g_y[7].g_x[4].t.r_v ),
    .X(_2100_));
 sg13g2_a21oi_1 _2683_ (.A1(_1992_),
    .A2(_2059_),
    .Y(_2101_),
    .B1(_2100_));
 sg13g2_buf_1 _2684_ (.A(\g.g_y[6].g_x[4].t.r_ghl ),
    .X(_2102_));
 sg13g2_buf_1 _2685_ (.A(\g.g_y[6].g_x[4].t.r_d ),
    .X(_2103_));
 sg13g2_mux2_1 _2686_ (.A0(\g.g_y[6].g_x[4].t.r_gnl ),
    .A1(\g.g_y[6].g_x[4].t.out_sc ),
    .S(_2103_),
    .X(_2104_));
 sg13g2_buf_2 _2687_ (.A(\g.g_y[6].g_x[4].t.r_v ),
    .X(_2105_));
 sg13g2_mux2_1 _2688_ (.A0(_2102_),
    .A1(_2104_),
    .S(_2105_),
    .X(_2106_));
 sg13g2_a22oi_1 _2689_ (.Y(_2107_),
    .B1(_2106_),
    .B2(_2100_),
    .A2(_2101_),
    .A1(_2099_));
 sg13g2_buf_1 _2690_ (.A(_2107_),
    .X(_2108_));
 sg13g2_or3_1 _2691_ (.A(net55),
    .B(_2098_),
    .C(_2108_),
    .X(_2109_));
 sg13g2_buf_1 _2692_ (.A(_2109_),
    .X(_2110_));
 sg13g2_inv_2 _2693_ (.Y(_2111_),
    .A(_2100_));
 sg13g2_inv_1 _2694_ (.Y(_2112_),
    .A(\g.g_y[7].g_x[4].t.r_d ));
 sg13g2_nor2_1 _2695_ (.A(_2112_),
    .B(\g.g_y[7].g_x[4].t.out_sc ),
    .Y(_2113_));
 sg13g2_nor2_1 _2696_ (.A(_2111_),
    .B(_2113_),
    .Y(_2114_));
 sg13g2_mux2_1 _2697_ (.A0(_1991_),
    .A1(_2058_),
    .S(_2082_),
    .X(_2115_));
 sg13g2_mux2_1 _2698_ (.A0(_2115_),
    .A1(_2106_),
    .S(_2111_),
    .X(_2116_));
 sg13g2_buf_2 _2699_ (.A(_2116_),
    .X(_2117_));
 sg13g2_mux2_1 _2700_ (.A0(_2093_),
    .A1(_2087_),
    .S(_2089_),
    .X(_2118_));
 sg13g2_mux2_1 _2701_ (.A0(_2118_),
    .A1(_2096_),
    .S(_2092_),
    .X(_2119_));
 sg13g2_mux2_1 _2702_ (.A0(_2117_),
    .A1(_2119_),
    .S(_2112_),
    .X(_2120_));
 sg13g2_buf_1 _2703_ (.A(_2120_),
    .X(_2121_));
 sg13g2_a221oi_1 _2704_ (.B2(_2111_),
    .C1(_2059_),
    .B1(_2121_),
    .A1(_2110_),
    .Y(_2122_),
    .A2(_2114_));
 sg13g2_nor3_1 _2705_ (.A(_2046_),
    .B(_2083_),
    .C(_2122_),
    .Y(_2123_));
 sg13g2_buf_1 _2706_ (.A(\g.g_y[0].g_x[5].t.r_v ),
    .X(_2124_));
 sg13g2_inv_1 _2707_ (.Y(_2125_),
    .A(net54));
 sg13g2_mux2_1 _2708_ (.A0(\g.g_y[1].g_x[5].t.r_gnl ),
    .A1(\g.g_y[1].g_x[5].t.out_sc ),
    .S(_2049_),
    .X(_2126_));
 sg13g2_buf_2 _2709_ (.A(\g.g_y[1].g_x[5].t.r_v ),
    .X(_2127_));
 sg13g2_inv_1 _2710_ (.Y(_2128_),
    .A(_2127_));
 sg13g2_mux2_1 _2711_ (.A0(\g.g_y[1].g_x[5].t.r_ghl ),
    .A1(_2126_),
    .S(_2128_),
    .X(_2129_));
 sg13g2_buf_1 _2712_ (.A(_2129_),
    .X(_2130_));
 sg13g2_buf_2 _2713_ (.A(\g.g_y[7].g_x[5].t.r_v ),
    .X(_2131_));
 sg13g2_inv_2 _2714_ (.Y(_2132_),
    .A(_2131_));
 sg13g2_mux2_1 _2715_ (.A0(\g.g_y[7].g_x[5].t.r_gnl ),
    .A1(\g.g_y[7].g_x[5].t.out_sc ),
    .S(_2085_),
    .X(_2133_));
 sg13g2_or2_1 _2716_ (.X(_2134_),
    .B(_2133_),
    .A(_2132_));
 sg13g2_buf_1 _2717_ (.A(_2134_),
    .X(_2135_));
 sg13g2_or2_1 _2718_ (.X(_2136_),
    .B(_2131_),
    .A(_2093_));
 sg13g2_and2_1 _2719_ (.A(net54),
    .B(_2136_),
    .X(_2137_));
 sg13g2_a22oi_1 _2720_ (.Y(_2138_),
    .B1(_2135_),
    .B2(_2137_),
    .A2(_2130_),
    .A1(_2125_));
 sg13g2_buf_1 _2721_ (.A(\g.g_y[0].g_x[5].t.r_d ),
    .X(_2139_));
 sg13g2_buf_2 _2722_ (.A(\g.g_y[0].g_x[6].t.r_d ),
    .X(_2140_));
 sg13g2_mux2_1 _2723_ (.A0(\g.g_y[0].g_x[6].t.out_sc ),
    .A1(\g.g_y[0].g_x[6].t.r_gnl ),
    .S(_2140_),
    .X(_2141_));
 sg13g2_inv_1 _2724_ (.Y(_2142_),
    .A(\g.g_y[0].g_x[6].t.r_h ));
 sg13g2_mux2_1 _2725_ (.A0(\g.g_y[0].g_x[6].t.r_ghl ),
    .A1(_2141_),
    .S(_2142_),
    .X(_2143_));
 sg13g2_buf_2 _2726_ (.A(_2143_),
    .X(_2144_));
 sg13g2_nand2_1 _2727_ (.Y(_2145_),
    .A(net53),
    .B(_2144_));
 sg13g2_buf_2 _2728_ (.A(\g.g_y[0].g_x[5].t.r_h ),
    .X(_2146_));
 sg13g2_nor2_1 _2729_ (.A(\g.g_y[0].g_x[5].t.out_sc ),
    .B(net53),
    .Y(_2147_));
 sg13g2_nor2_1 _2730_ (.A(_2146_),
    .B(_2147_),
    .Y(_2148_));
 sg13g2_o21ai_1 _2731_ (.B1(_2148_),
    .Y(_2149_),
    .A1(_2138_),
    .A2(_2145_));
 sg13g2_and2_1 _2732_ (.A(_2125_),
    .B(_2136_),
    .X(_2150_));
 sg13g2_inv_1 _2733_ (.Y(_2151_),
    .A(net53));
 sg13g2_a221oi_1 _2734_ (.B2(_2150_),
    .C1(_2151_),
    .B1(_2135_),
    .A1(net54),
    .Y(_2152_),
    .A2(_2130_));
 sg13g2_buf_1 _2735_ (.A(_2152_),
    .X(_2153_));
 sg13g2_o21ai_1 _2736_ (.B1(_2146_),
    .Y(_2154_),
    .A1(net53),
    .A2(_2144_));
 sg13g2_or2_1 _2737_ (.X(_2155_),
    .B(_2154_),
    .A(_2153_));
 sg13g2_nand3_1 _2738_ (.B(_2149_),
    .C(_2155_),
    .A(_1988_),
    .Y(_2156_));
 sg13g2_o21ai_1 _2739_ (.B1(_2012_),
    .Y(_2157_),
    .A1(_1994_),
    .A2(_2005_));
 sg13g2_and2_1 _2740_ (.A(_1984_),
    .B(_2016_),
    .X(_2158_));
 sg13g2_a221oi_1 _2741_ (.B2(\g.g_y[0].g_x[3].t.out_sc ),
    .C1(_2158_),
    .B1(_2015_),
    .A1(_2007_),
    .Y(_2159_),
    .A2(_2011_));
 sg13g2_nand3_1 _2742_ (.B(_2157_),
    .C(_2159_),
    .A(_1989_),
    .Y(_2160_));
 sg13g2_nand3_1 _2743_ (.B(_2156_),
    .C(_2160_),
    .A(_2046_),
    .Y(_2161_));
 sg13g2_nand2b_1 _2744_ (.Y(\g.g_y[0].g_x[4].t.w_dh ),
    .B(_2161_),
    .A_N(_2123_));
 sg13g2_a21oi_1 _2745_ (.A1(_2157_),
    .A2(_2159_),
    .Y(_2162_),
    .B1(_1989_));
 sg13g2_a21oi_1 _2746_ (.A1(_2149_),
    .A2(_2155_),
    .Y(_2163_),
    .B1(_1988_));
 sg13g2_a22oi_1 _2747_ (.Y(_2164_),
    .B1(_2121_),
    .B2(_2111_),
    .A2(_2114_),
    .A1(_2110_));
 sg13g2_a221oi_1 _2748_ (.B2(net57),
    .C1(_2059_),
    .B1(_2081_),
    .A1(_2072_),
    .Y(_2165_),
    .A2(_2074_));
 sg13g2_a21oi_1 _2749_ (.A1(_2059_),
    .A2(_2164_),
    .Y(_2166_),
    .B1(_2165_));
 sg13g2_o21ai_1 _2750_ (.B1(_2166_),
    .Y(\g.g_y[0].g_x[4].t.w_na ),
    .A1(_2162_),
    .A2(_2163_));
 sg13g2_or4_1 _2751_ (.A(_1985_),
    .B(net78),
    .C(_2083_),
    .D(_2122_),
    .X(_2167_));
 sg13g2_nand4_1 _2752_ (.B(net64),
    .C(_2156_),
    .A(_1985_),
    .Y(_2168_),
    .D(_2160_));
 sg13g2_nand2_1 _2753_ (.Y(_2169_),
    .A(\g.g_y[0].g_x[3].t.out_sc ),
    .B(net61));
 sg13g2_nand3_1 _2754_ (.B(_2168_),
    .C(_2169_),
    .A(_2167_),
    .Y(\g.g_y[0].g_x[4].t.w_si ));
 sg13g2_or2_1 _2755_ (.X(_2170_),
    .B(_1987_),
    .A(_1989_));
 sg13g2_a21oi_1 _2756_ (.A1(_1992_),
    .A2(_1989_),
    .Y(_2171_),
    .B1(_2146_));
 sg13g2_a22oi_1 _2757_ (.Y(_2172_),
    .B1(_2170_),
    .B2(_2171_),
    .A2(_2144_),
    .A1(_2146_));
 sg13g2_a221oi_1 _2758_ (.B2(_2150_),
    .C1(net53),
    .B1(_2135_),
    .A1(net54),
    .Y(_2173_),
    .A2(_2130_));
 sg13g2_a21o_1 _2759_ (.A2(_2172_),
    .A1(net53),
    .B1(_2173_),
    .X(_2174_));
 sg13g2_buf_1 _2760_ (.A(net77),
    .X(_2175_));
 sg13g2_nand2_1 _2761_ (.Y(_2176_),
    .A(\g.g_y[0].g_x[4].t.out_sc ),
    .B(net52));
 sg13g2_o21ai_1 _2762_ (.B1(_2176_),
    .Y(\g.g_y[0].g_x[5].t.w_si ),
    .A1(net60),
    .A2(_2174_));
 sg13g2_buf_2 _2763_ (.A(\g.g_y[0].g_x[7].t.r_h ),
    .X(_2177_));
 sg13g2_mux2_1 _2764_ (.A0(\g.g_y[0].g_x[6].t.r_ghl ),
    .A1(_2141_),
    .S(\g.g_y[0].g_x[6].t.r_h ),
    .X(_2178_));
 sg13g2_nand2b_1 _2765_ (.Y(_2179_),
    .B(_1816_),
    .A_N(_1790_));
 sg13g2_inv_1 _2766_ (.Y(_2180_),
    .A(_1788_));
 sg13g2_a21oi_1 _2767_ (.A1(_2180_),
    .A2(_1791_),
    .Y(_2181_),
    .B1(_2177_));
 sg13g2_a22oi_1 _2768_ (.Y(_2182_),
    .B1(_2179_),
    .B2(_2181_),
    .A2(_2178_),
    .A1(_2177_));
 sg13g2_buf_2 _2769_ (.A(\g.g_y[7].g_x[7].t.r_d ),
    .X(_2183_));
 sg13g2_mux2_1 _2770_ (.A0(\g.g_y[7].g_x[7].t.r_gnl ),
    .A1(\g.g_y[7].g_x[7].t.out_sc ),
    .S(_2183_),
    .X(_2184_));
 sg13g2_buf_1 _2771_ (.A(\g.g_y[7].g_x[7].t.r_v ),
    .X(_2185_));
 sg13g2_mux2_1 _2772_ (.A0(\g.g_y[7].g_x[7].t.r_ghl ),
    .A1(_2184_),
    .S(_2185_),
    .X(_2186_));
 sg13g2_buf_1 _2773_ (.A(_2186_),
    .X(_2187_));
 sg13g2_buf_1 _2774_ (.A(\g.g_y[1].g_x[7].t.r_ghl ),
    .X(_2188_));
 sg13g2_buf_2 _2775_ (.A(\g.g_y[1].g_x[7].t.r_d ),
    .X(_2189_));
 sg13g2_mux2_1 _2776_ (.A0(\g.g_y[1].g_x[7].t.r_gnl ),
    .A1(\g.g_y[1].g_x[7].t.out_sc ),
    .S(_2189_),
    .X(_2190_));
 sg13g2_buf_2 _2777_ (.A(_2190_),
    .X(_2191_));
 sg13g2_buf_2 _2778_ (.A(\g.g_y[1].g_x[7].t.r_v ),
    .X(_2192_));
 sg13g2_inv_1 _2779_ (.Y(_2193_),
    .A(_2192_));
 sg13g2_mux2_1 _2780_ (.A0(_2188_),
    .A1(_2191_),
    .S(_2193_),
    .X(_2194_));
 sg13g2_buf_2 _2781_ (.A(\g.g_y[0].g_x[7].t.r_v ),
    .X(_2195_));
 sg13g2_inv_1 _2782_ (.Y(_2196_),
    .A(_2195_));
 sg13g2_mux2_1 _2783_ (.A0(_2187_),
    .A1(_2194_),
    .S(_2196_),
    .X(_2197_));
 sg13g2_buf_1 _2784_ (.A(\g.g_y[0].g_x[7].t.r_d ),
    .X(_2198_));
 sg13g2_buf_1 _2785_ (.A(_2198_),
    .X(_2199_));
 sg13g2_nand3b_1 _2786_ (.B(_2197_),
    .C(net28),
    .Y(_2200_),
    .A_N(_2182_));
 sg13g2_buf_1 _2787_ (.A(\g.g_y[0].g_x[7].t.out_sc ),
    .X(_2201_));
 sg13g2_nor2_1 _2788_ (.A(_2201_),
    .B(net28),
    .Y(_2202_));
 sg13g2_nor2_1 _2789_ (.A(_2177_),
    .B(_2202_),
    .Y(_2203_));
 sg13g2_mux2_1 _2790_ (.A0(_1788_),
    .A1(_1790_),
    .S(_1816_),
    .X(_2204_));
 sg13g2_mux2_1 _2791_ (.A0(_2178_),
    .A1(_2204_),
    .S(_2177_),
    .X(_2205_));
 sg13g2_buf_1 _2792_ (.A(_2205_),
    .X(_2206_));
 sg13g2_mux2_1 _2793_ (.A0(_2187_),
    .A1(_2194_),
    .S(_2195_),
    .X(_2207_));
 sg13g2_mux2_1 _2794_ (.A0(_2206_),
    .A1(_2207_),
    .S(net28),
    .X(_2208_));
 sg13g2_a221oi_1 _2795_ (.B2(_2177_),
    .C1(_2142_),
    .B1(_2208_),
    .A1(_2200_),
    .Y(_2209_),
    .A2(_2203_));
 sg13g2_mux2_1 _2796_ (.A0(_1991_),
    .A1(_1987_),
    .S(_1988_),
    .X(_2210_));
 sg13g2_nand2_1 _2797_ (.Y(_2211_),
    .A(_2139_),
    .B(_2210_));
 sg13g2_nor2b_1 _2798_ (.A(_2147_),
    .B_N(_2146_),
    .Y(_2212_));
 sg13g2_o21ai_1 _2799_ (.B1(_2212_),
    .Y(_2213_),
    .A1(_2138_),
    .A2(_2211_));
 sg13g2_nor2_1 _2800_ (.A(_2139_),
    .B(_2210_),
    .Y(_2214_));
 sg13g2_or3_1 _2801_ (.A(_2146_),
    .B(_2153_),
    .C(_2214_),
    .X(_2215_));
 sg13g2_nand3_1 _2802_ (.B(_2213_),
    .C(_2215_),
    .A(_2142_),
    .Y(_2216_));
 sg13g2_nand2b_1 _2803_ (.Y(_2217_),
    .B(_2216_),
    .A_N(_2209_));
 sg13g2_buf_1 _2804_ (.A(\g.g_y[1].g_x[6].t.r_v ),
    .X(_2218_));
 sg13g2_buf_1 _2805_ (.A(\g.g_y[1].g_x[6].t.r_d ),
    .X(_2219_));
 sg13g2_buf_1 _2806_ (.A(\g.g_y[1].g_x[6].t.r_h ),
    .X(_2220_));
 sg13g2_mux2_1 _2807_ (.A0(\g.g_y[1].g_x[5].t.r_ghl ),
    .A1(_2050_),
    .S(\g.g_y[1].g_x[5].t.r_h ),
    .X(_2221_));
 sg13g2_buf_1 _2808_ (.A(_2221_),
    .X(_2222_));
 sg13g2_buf_2 _2809_ (.A(\g.g_y[1].g_x[7].t.r_h ),
    .X(_2223_));
 sg13g2_mux2_1 _2810_ (.A0(\g.g_y[1].g_x[7].t.out_sc ),
    .A1(\g.g_y[1].g_x[7].t.r_gnl ),
    .S(_2189_),
    .X(_2224_));
 sg13g2_or2_1 _2811_ (.X(_2225_),
    .B(_2224_),
    .A(_2223_));
 sg13g2_buf_1 _2812_ (.A(_2225_),
    .X(_2226_));
 sg13g2_inv_1 _2813_ (.Y(_2227_),
    .A(_2220_));
 sg13g2_nand2b_1 _2814_ (.Y(_2228_),
    .B(_2223_),
    .A_N(_2188_));
 sg13g2_and2_1 _2815_ (.A(_2227_),
    .B(_2228_),
    .X(_2229_));
 sg13g2_a22oi_1 _2816_ (.Y(_2230_),
    .B1(_2226_),
    .B2(_2229_),
    .A2(_2222_),
    .A1(_2220_));
 sg13g2_buf_1 _2817_ (.A(_2230_),
    .X(_2231_));
 sg13g2_mux2_1 _2818_ (.A0(\g.g_y[0].g_x[6].t.r_gnl ),
    .A1(\g.g_y[0].g_x[6].t.out_sc ),
    .S(_2140_),
    .X(_2232_));
 sg13g2_buf_2 _2819_ (.A(\g.g_y[0].g_x[6].t.r_v ),
    .X(_2233_));
 sg13g2_mux2_1 _2820_ (.A0(\g.g_y[0].g_x[6].t.r_ghl ),
    .A1(_2232_),
    .S(_2233_),
    .X(_2234_));
 sg13g2_buf_8 _2821_ (.A(\g.g_y[2].g_x[6].t.r_d ),
    .X(_2235_));
 sg13g2_mux2_1 _2822_ (.A0(\g.g_y[2].g_x[6].t.r_gnl ),
    .A1(\g.g_y[2].g_x[6].t.out_sc ),
    .S(_2235_),
    .X(_2236_));
 sg13g2_buf_1 _2823_ (.A(_2236_),
    .X(_2237_));
 sg13g2_buf_2 _2824_ (.A(\g.g_y[2].g_x[6].t.r_v ),
    .X(_2238_));
 sg13g2_inv_1 _2825_ (.Y(_2239_),
    .A(_2238_));
 sg13g2_nand2b_1 _2826_ (.Y(_2240_),
    .B(_2239_),
    .A_N(_2237_));
 sg13g2_buf_2 _2827_ (.A(\g.g_y[2].g_x[6].t.r_ghl ),
    .X(_2241_));
 sg13g2_inv_1 _2828_ (.Y(_2242_),
    .A(_2241_));
 sg13g2_a21oi_1 _2829_ (.A1(_2242_),
    .A2(_2238_),
    .Y(_2243_),
    .B1(net51));
 sg13g2_a22oi_1 _2830_ (.Y(_2244_),
    .B1(_2240_),
    .B2(_2243_),
    .A2(_2234_),
    .A1(net51));
 sg13g2_buf_1 _2831_ (.A(_2244_),
    .X(_2245_));
 sg13g2_or4_1 _2832_ (.A(net51),
    .B(_2219_),
    .C(_2231_),
    .D(_2245_),
    .X(_2246_));
 sg13g2_and2_1 _2833_ (.A(_2220_),
    .B(_2228_),
    .X(_2247_));
 sg13g2_a221oi_1 _2834_ (.B2(_2247_),
    .C1(_2219_),
    .B1(_2226_),
    .A1(_2227_),
    .Y(_2248_),
    .A2(_2222_));
 sg13g2_inv_1 _2835_ (.Y(_2249_),
    .A(net51));
 sg13g2_a21oi_1 _2836_ (.A1(_2242_),
    .A2(_2238_),
    .Y(_2250_),
    .B1(_2249_));
 sg13g2_inv_1 _2837_ (.Y(_2251_),
    .A(_2219_));
 sg13g2_a221oi_1 _2838_ (.B2(_2250_),
    .C1(_2251_),
    .B1(_2240_),
    .A1(_2249_),
    .Y(_2252_),
    .A2(_2234_));
 sg13g2_o21ai_1 _2839_ (.B1(net51),
    .Y(_2253_),
    .A1(_2248_),
    .A2(_2252_));
 sg13g2_inv_1 _2840_ (.Y(_2254_),
    .A(_2233_));
 sg13g2_a21o_1 _2841_ (.A2(_2253_),
    .A1(_2246_),
    .B1(_2254_),
    .X(_2255_));
 sg13g2_buf_1 _2842_ (.A(\g.g_y[7].g_x[6].t.r_v ),
    .X(_2256_));
 sg13g2_mux2_1 _2843_ (.A0(\g.g_y[0].g_x[6].t.r_ghl ),
    .A1(_2232_),
    .S(_2254_),
    .X(_2257_));
 sg13g2_buf_1 _2844_ (.A(\g.g_y[6].g_x[6].t.r_v ),
    .X(_2258_));
 sg13g2_inv_1 _2845_ (.Y(_2259_),
    .A(net49));
 sg13g2_buf_2 _2846_ (.A(\g.g_y[6].g_x[6].t.r_d ),
    .X(_2260_));
 sg13g2_mux2_1 _2847_ (.A0(\g.g_y[6].g_x[6].t.r_gnl ),
    .A1(\g.g_y[6].g_x[6].t.out_sc ),
    .S(_2260_),
    .X(_2261_));
 sg13g2_buf_1 _2848_ (.A(_2261_),
    .X(_2262_));
 sg13g2_or2_1 _2849_ (.X(_2263_),
    .B(_2262_),
    .A(_2259_));
 sg13g2_buf_2 _2850_ (.A(\g.g_y[6].g_x[6].t.r_ghl ),
    .X(_2264_));
 sg13g2_nor2_1 _2851_ (.A(_2264_),
    .B(net49),
    .Y(_2265_));
 sg13g2_nor2_1 _2852_ (.A(net50),
    .B(_2265_),
    .Y(_2266_));
 sg13g2_buf_1 _2853_ (.A(\g.g_y[7].g_x[6].t.r_d ),
    .X(_2267_));
 sg13g2_inv_1 _2854_ (.Y(_2268_),
    .A(net48));
 sg13g2_a221oi_1 _2855_ (.B2(_2266_),
    .C1(_2268_),
    .B1(_2263_),
    .A1(net50),
    .Y(_2269_),
    .A2(_2257_));
 sg13g2_buf_2 _2856_ (.A(\g.g_y[7].g_x[7].t.r_h ),
    .X(_2270_));
 sg13g2_mux2_1 _2857_ (.A0(\g.g_y[7].g_x[7].t.out_sc ),
    .A1(\g.g_y[7].g_x[7].t.r_gnl ),
    .S(_2183_),
    .X(_2271_));
 sg13g2_or2_1 _2858_ (.X(_2272_),
    .B(_2271_),
    .A(_2270_));
 sg13g2_buf_1 _2859_ (.A(_2272_),
    .X(_2273_));
 sg13g2_buf_2 _2860_ (.A(\g.g_y[7].g_x[6].t.r_h ),
    .X(_2274_));
 sg13g2_nand2b_1 _2861_ (.Y(_2275_),
    .B(_2270_),
    .A_N(\g.g_y[7].g_x[7].t.r_ghl ));
 sg13g2_and2_1 _2862_ (.A(_2274_),
    .B(_2275_),
    .X(_2276_));
 sg13g2_mux2_1 _2863_ (.A0(_2093_),
    .A1(_2087_),
    .S(_2088_),
    .X(_2277_));
 sg13g2_buf_1 _2864_ (.A(_2277_),
    .X(_2278_));
 sg13g2_inv_1 _2865_ (.Y(_2279_),
    .A(_2274_));
 sg13g2_a221oi_1 _2866_ (.B2(_2279_),
    .C1(net48),
    .B1(_2278_),
    .A1(_2273_),
    .Y(_0000_),
    .A2(_2276_));
 sg13g2_or2_1 _2867_ (.X(_0001_),
    .B(_0000_),
    .A(_2269_));
 sg13g2_nand2b_1 _2868_ (.Y(_0002_),
    .B(_2219_),
    .A_N(\g.g_y[1].g_x[6].t.out_sc ));
 sg13g2_nor3_1 _2869_ (.A(_2254_),
    .B(net51),
    .C(_0002_),
    .Y(_0003_));
 sg13g2_inv_2 _2870_ (.Y(_0004_),
    .A(net50));
 sg13g2_buf_1 _2871_ (.A(\g.g_y[7].g_x[6].t.out_sc ),
    .X(_0005_));
 sg13g2_nor2_1 _2872_ (.A(_2268_),
    .B(_0005_),
    .Y(_0006_));
 sg13g2_o21ai_1 _2873_ (.B1(_2254_),
    .Y(_0007_),
    .A1(_0004_),
    .A2(_0006_));
 sg13g2_nand2b_1 _2874_ (.Y(_0008_),
    .B(_0007_),
    .A_N(_0003_));
 sg13g2_o21ai_1 _2875_ (.B1(_0008_),
    .Y(_0009_),
    .A1(_2233_),
    .A2(_0001_));
 sg13g2_and2_1 _2876_ (.A(_2279_),
    .B(_2275_),
    .X(_0010_));
 sg13g2_a22oi_1 _2877_ (.Y(_0011_),
    .B1(_0010_),
    .B2(_2273_),
    .A2(_2278_),
    .A1(_2274_));
 sg13g2_buf_1 _2878_ (.A(_0011_),
    .X(_0012_));
 sg13g2_nor2_1 _2879_ (.A(_0004_),
    .B(_2265_),
    .Y(_0013_));
 sg13g2_a22oi_1 _2880_ (.Y(_0014_),
    .B1(_2263_),
    .B2(_0013_),
    .A2(_2257_),
    .A1(_0004_));
 sg13g2_buf_1 _2881_ (.A(_0014_),
    .X(_0015_));
 sg13g2_nor3_2 _2882_ (.A(net48),
    .B(_0012_),
    .C(_0015_),
    .Y(_0016_));
 sg13g2_nor2_1 _2883_ (.A(_2233_),
    .B(_0004_),
    .Y(_0017_));
 sg13g2_a22oi_1 _2884_ (.Y(_0018_),
    .B1(_0016_),
    .B2(_0017_),
    .A2(_0008_),
    .A1(_2256_));
 sg13g2_nand4_1 _2885_ (.B(_2255_),
    .C(_0009_),
    .A(_2140_),
    .Y(_0019_),
    .D(_0018_));
 sg13g2_o21ai_1 _2886_ (.B1(_0019_),
    .Y(\g.g_y[0].g_x[6].t.w_dh ),
    .A1(_2140_),
    .A2(_2217_));
 sg13g2_nor2_1 _2887_ (.A(_2248_),
    .B(_2252_),
    .Y(_0020_));
 sg13g2_nor2_1 _2888_ (.A(_2249_),
    .B(_0020_),
    .Y(_0021_));
 sg13g2_or3_1 _2889_ (.A(_2219_),
    .B(_2231_),
    .C(_2245_),
    .X(_0022_));
 sg13g2_buf_1 _2890_ (.A(_0022_),
    .X(_0023_));
 sg13g2_a21oi_1 _2891_ (.A1(_0023_),
    .A2(_0002_),
    .Y(_0024_),
    .B1(net51));
 sg13g2_o21ai_1 _2892_ (.B1(_2254_),
    .Y(_0025_),
    .A1(_0021_),
    .A2(_0024_));
 sg13g2_o21ai_1 _2893_ (.B1(_2256_),
    .Y(_0026_),
    .A1(_0006_),
    .A2(_0016_));
 sg13g2_nand2_1 _2894_ (.Y(_0027_),
    .A(_0004_),
    .B(_0001_));
 sg13g2_a21o_1 _2895_ (.A2(_0027_),
    .A1(_0026_),
    .B1(_2254_),
    .X(_0028_));
 sg13g2_and2_1 _2896_ (.A(_2213_),
    .B(_2215_),
    .X(_0029_));
 sg13g2_a221oi_1 _2897_ (.B2(_2177_),
    .C1(\g.g_y[0].g_x[6].t.r_h ),
    .B1(_2208_),
    .A1(_2200_),
    .Y(_0030_),
    .A2(_2203_));
 sg13g2_a21oi_1 _2898_ (.A1(\g.g_y[0].g_x[6].t.r_h ),
    .A2(_0029_),
    .Y(_0031_),
    .B1(_0030_));
 sg13g2_nand3_1 _2899_ (.B(_0028_),
    .C(_0031_),
    .A(_0025_),
    .Y(\g.g_y[0].g_x[6].t.w_na ));
 sg13g2_and2_1 _2900_ (.A(_2140_),
    .B(net81),
    .X(_0032_));
 sg13g2_nand3b_1 _2901_ (.B(_2216_),
    .C(_0032_),
    .Y(_0033_),
    .A_N(_2209_));
 sg13g2_nor2_1 _2902_ (.A(_2140_),
    .B(net77),
    .Y(_0034_));
 sg13g2_nand4_1 _2903_ (.B(_0009_),
    .C(_0018_),
    .A(_2255_),
    .Y(_0035_),
    .D(_0034_));
 sg13g2_nand2_1 _2904_ (.Y(_0036_),
    .A(\g.g_y[0].g_x[5].t.out_sc ),
    .B(net61));
 sg13g2_nand3_1 _2905_ (.B(_0035_),
    .C(_0036_),
    .A(_0033_),
    .Y(\g.g_y[0].g_x[6].t.w_si ));
 sg13g2_inv_1 _2906_ (.Y(_0037_),
    .A(_2177_));
 sg13g2_o21ai_1 _2907_ (.B1(_2200_),
    .Y(_0038_),
    .A1(_2201_),
    .A2(net28));
 sg13g2_nand2_1 _2908_ (.Y(_0039_),
    .A(_0037_),
    .B(_2208_));
 sg13g2_o21ai_1 _2909_ (.B1(_0039_),
    .Y(\g.g_y[0].g_x[7].t.out_r ),
    .A1(_0037_),
    .A2(_0038_));
 sg13g2_mux2_1 _2910_ (.A0(_2207_),
    .A1(_2206_),
    .S(net28),
    .X(_0040_));
 sg13g2_mux2_1 _2911_ (.A0(\g.g_y[0].g_x[6].t.out_sc ),
    .A1(_0040_),
    .S(net64),
    .X(\g.g_y[0].g_x[7].t.w_si ));
 sg13g2_mux2_1 _2912_ (.A0(\g.g_y[0].g_x[0].t.r_gnl ),
    .A1(\g.g_y[0].g_x[0].t.out_sc ),
    .S(_1789_),
    .X(_0041_));
 sg13g2_or2_1 _2913_ (.X(_0042_),
    .B(_1820_),
    .A(_1788_));
 sg13g2_o21ai_1 _2914_ (.B1(_0042_),
    .Y(_0043_),
    .A1(_1852_),
    .A2(_0041_));
 sg13g2_mux2_1 _2915_ (.A0(_0043_),
    .A1(_1838_),
    .S(_1821_),
    .X(_0044_));
 sg13g2_a21oi_1 _2916_ (.A1(_1822_),
    .A2(_1827_),
    .Y(_0045_),
    .B1(_1829_));
 sg13g2_mux2_1 _2917_ (.A0(_0044_),
    .A1(_0045_),
    .S(net29),
    .X(_0046_));
 sg13g2_nand2_1 _2918_ (.Y(_0047_),
    .A(_2201_),
    .B(net52));
 sg13g2_o21ai_1 _2919_ (.B1(_0047_),
    .Y(\g.g_y[1].g_x[0].t.w_si ),
    .A1(_2040_),
    .A2(_0046_));
 sg13g2_a21oi_1 _2920_ (.A1(net15),
    .A2(_1781_),
    .Y(\g.g_y[1].g_x[1].t.in_lb ),
    .B1(_1903_));
 sg13g2_inv_1 _2921_ (.Y(_0048_),
    .A(_1802_));
 sg13g2_nor2b_1 _2922_ (.A(_1914_),
    .B_N(net63),
    .Y(_0049_));
 sg13g2_o21ai_1 _2923_ (.B1(_0049_),
    .Y(_0050_),
    .A1(_1917_),
    .A2(_1931_));
 sg13g2_and2_1 _2924_ (.A(_1914_),
    .B(net63),
    .X(_0051_));
 sg13g2_nor2_1 _2925_ (.A(_1914_),
    .B(net63),
    .Y(_0052_));
 sg13g2_nor2_1 _2926_ (.A(_1937_),
    .B(net63),
    .Y(_0053_));
 sg13g2_and2_1 _2927_ (.A(_1936_),
    .B(_0053_),
    .X(_0054_));
 sg13g2_a221oi_1 _2928_ (.B2(\g.g_y[1].g_x[2].t.out_sc ),
    .C1(_0054_),
    .B1(_0052_),
    .A1(_1942_),
    .Y(_0055_),
    .A2(_0051_));
 sg13g2_nand3_1 _2929_ (.B(_0050_),
    .C(_0055_),
    .A(_1824_),
    .Y(_0056_));
 sg13g2_inv_1 _2930_ (.Y(_0057_),
    .A(_1833_));
 sg13g2_mux2_1 _2931_ (.A0(_1836_),
    .A1(_1835_),
    .S(_0057_),
    .X(_0058_));
 sg13g2_mux2_1 _2932_ (.A0(_1788_),
    .A1(_0041_),
    .S(_1820_),
    .X(_0059_));
 sg13g2_mux2_1 _2933_ (.A0(_0058_),
    .A1(_0059_),
    .S(_1821_),
    .X(_0060_));
 sg13g2_and2_1 _2934_ (.A(net2),
    .B(net29),
    .X(_0061_));
 sg13g2_o21ai_1 _2935_ (.B1(_1822_),
    .Y(_0062_),
    .A1(net29),
    .A2(\g.g_y[1].g_x[0].t.out_sc ));
 sg13g2_a21oi_1 _2936_ (.A1(_0060_),
    .A2(_0061_),
    .Y(_0063_),
    .B1(_0062_));
 sg13g2_nor2_1 _2937_ (.A(net2),
    .B(_1828_),
    .Y(_0064_));
 sg13g2_nor2_1 _2938_ (.A(_1822_),
    .B(_0064_),
    .Y(_0065_));
 sg13g2_inv_1 _2939_ (.Y(_0066_),
    .A(_0065_));
 sg13g2_a21oi_1 _2940_ (.A1(net29),
    .A2(_0044_),
    .Y(_0067_),
    .B1(_0066_));
 sg13g2_or3_1 _2941_ (.A(_1824_),
    .B(_0063_),
    .C(_0067_),
    .X(_0068_));
 sg13g2_and3_1 _2942_ (.X(_0069_),
    .A(_0048_),
    .B(_0056_),
    .C(_0068_));
 sg13g2_nand3b_1 _2943_ (.B(_1794_),
    .C(_1808_),
    .Y(_0070_),
    .A_N(net66));
 sg13g2_buf_1 _2944_ (.A(_0070_),
    .X(_0071_));
 sg13g2_nand2b_1 _2945_ (.Y(_0072_),
    .B(net66),
    .A_N(\g.g_y[0].g_x[1].t.out_sc ));
 sg13g2_and2_1 _2946_ (.A(_1806_),
    .B(_0072_),
    .X(_0073_));
 sg13g2_a221oi_1 _2947_ (.B2(_0073_),
    .C1(\g.g_y[1].g_x[1].t.r_v ),
    .B1(_0071_),
    .A1(_1807_),
    .Y(_0074_),
    .A2(_1815_));
 sg13g2_mux2_1 _2948_ (.A0(\g.g_y[2].g_x[0].t.out_sc ),
    .A1(\g.g_y[2].g_x[0].t.r_gnl ),
    .S(_1834_),
    .X(_0075_));
 sg13g2_buf_1 _2949_ (.A(\g.g_y[2].g_x[0].t.r_h ),
    .X(_0076_));
 sg13g2_mux2_1 _2950_ (.A0(_1836_),
    .A1(_0075_),
    .S(_0076_),
    .X(_0077_));
 sg13g2_mux2_1 _2951_ (.A0(\g.g_y[2].g_x[2].t.out_sc ),
    .A1(\g.g_y[2].g_x[2].t.r_gnl ),
    .S(_1918_),
    .X(_0078_));
 sg13g2_buf_2 _2952_ (.A(\g.g_y[2].g_x[2].t.r_h ),
    .X(_0079_));
 sg13g2_inv_1 _2953_ (.Y(_0080_),
    .A(_0079_));
 sg13g2_mux2_1 _2954_ (.A0(_1923_),
    .A1(_0078_),
    .S(_0080_),
    .X(_0081_));
 sg13g2_buf_1 _2955_ (.A(\g.g_y[2].g_x[1].t.r_h ),
    .X(_0082_));
 sg13g2_inv_2 _2956_ (.Y(_0083_),
    .A(_0082_));
 sg13g2_mux2_1 _2957_ (.A0(_0077_),
    .A1(_0081_),
    .S(_0083_),
    .X(_0084_));
 sg13g2_buf_1 _2958_ (.A(\g.g_y[2].g_x[1].t.r_d ),
    .X(_0085_));
 sg13g2_buf_1 _2959_ (.A(_0085_),
    .X(_0086_));
 sg13g2_buf_1 _2960_ (.A(\g.g_y[3].g_x[1].t.r_v ),
    .X(_0087_));
 sg13g2_buf_8 _2961_ (.A(\g.g_y[3].g_x[1].t.r_d ),
    .X(_0088_));
 sg13g2_mux2_1 _2962_ (.A0(\g.g_y[3].g_x[1].t.r_gnl ),
    .A1(\g.g_y[3].g_x[1].t.out_sc ),
    .S(_0088_),
    .X(_0089_));
 sg13g2_nand2b_1 _2963_ (.Y(_0090_),
    .B(_0087_),
    .A_N(\g.g_y[3].g_x[1].t.r_ghl ));
 sg13g2_o21ai_1 _2964_ (.B1(_0090_),
    .Y(_0091_),
    .A1(_0087_),
    .A2(_0089_));
 sg13g2_nor2_1 _2965_ (.A(net27),
    .B(_0091_),
    .Y(_0092_));
 sg13g2_nand2_1 _2966_ (.Y(_0093_),
    .A(_0084_),
    .B(_0092_));
 sg13g2_inv_1 _2967_ (.Y(_0094_),
    .A(\g.g_y[2].g_x[1].t.out_sc ));
 sg13g2_buf_1 _2968_ (.A(\g.g_y[2].g_x[1].t.r_v ),
    .X(_0095_));
 sg13g2_a21oi_1 _2969_ (.A1(net27),
    .A2(_0094_),
    .Y(_0096_),
    .B1(_0095_));
 sg13g2_nand2b_1 _2970_ (.Y(_0097_),
    .B(_0080_),
    .A_N(_0078_));
 sg13g2_a21oi_1 _2971_ (.A1(_1924_),
    .A2(_0079_),
    .Y(_0098_),
    .B1(_0083_));
 sg13g2_a221oi_1 _2972_ (.B2(_0098_),
    .C1(_0085_),
    .B1(_0097_),
    .A1(_0083_),
    .Y(_0099_),
    .A2(_0077_));
 sg13g2_a21oi_1 _2973_ (.A1(net27),
    .A2(_0091_),
    .Y(_0100_),
    .B1(_0099_));
 sg13g2_a221oi_1 _2974_ (.B2(_0095_),
    .C1(_1804_),
    .B1(_0100_),
    .A1(_0093_),
    .Y(_0101_),
    .A2(_0096_));
 sg13g2_nor3_1 _2975_ (.A(_0048_),
    .B(_0074_),
    .C(_0101_),
    .Y(_0102_));
 sg13g2_or2_1 _2976_ (.X(\g.g_y[1].g_x[1].t.w_dh ),
    .B(_0102_),
    .A(_0069_));
 sg13g2_nand3_1 _2977_ (.B(_0050_),
    .C(_0055_),
    .A(_1825_),
    .Y(_0103_));
 sg13g2_a22oi_1 _2978_ (.Y(_0104_),
    .B1(_0071_),
    .B2(_0073_),
    .A2(_1815_),
    .A1(_1807_));
 sg13g2_nand2_1 _2979_ (.Y(_0105_),
    .A(\g.g_y[1].g_x[1].t.r_v ),
    .B(_0104_));
 sg13g2_nor2_1 _2980_ (.A(_0063_),
    .B(_0067_),
    .Y(_0106_));
 sg13g2_a22oi_1 _2981_ (.Y(_0107_),
    .B1(_0100_),
    .B2(_0095_),
    .A2(_0096_),
    .A1(_0093_));
 sg13g2_a22oi_1 _2982_ (.Y(_0108_),
    .B1(_0107_),
    .B2(_1804_),
    .A2(_0106_),
    .A1(_1824_));
 sg13g2_nand3_1 _2983_ (.B(_0105_),
    .C(_0108_),
    .A(_0103_),
    .Y(\g.g_y[1].g_x[1].t.w_na ));
 sg13g2_buf_1 _2984_ (.A(net77),
    .X(_0109_));
 sg13g2_nand2_1 _2985_ (.Y(_0110_),
    .A(\g.g_y[1].g_x[0].t.out_sc ),
    .B(net47));
 sg13g2_buf_1 _2986_ (.A(_1893_),
    .X(_0111_));
 sg13g2_or4_1 _2987_ (.A(_1802_),
    .B(net74),
    .C(_0074_),
    .D(_0101_),
    .X(_0112_));
 sg13g2_buf_1 _2988_ (.A(_1900_),
    .X(_0113_));
 sg13g2_nand4_1 _2989_ (.B(net73),
    .C(_0056_),
    .A(_1802_),
    .Y(_0114_),
    .D(_0068_));
 sg13g2_nand3_1 _2990_ (.B(_0112_),
    .C(_0114_),
    .A(_0110_),
    .Y(\g.g_y[1].g_x[1].t.w_si ));
 sg13g2_nor2b_1 _2991_ (.A(net63),
    .B_N(_1942_),
    .Y(_0115_));
 sg13g2_a21oi_1 _2992_ (.A1(net63),
    .A2(_1938_),
    .Y(_0116_),
    .B1(_0115_));
 sg13g2_nand2_1 _2993_ (.Y(_0117_),
    .A(\g.g_y[1].g_x[1].t.out_sc ),
    .B(net52));
 sg13g2_o21ai_1 _2994_ (.B1(_0117_),
    .Y(\g.g_y[1].g_x[2].t.w_si ),
    .A1(net60),
    .A2(_0116_));
 sg13g2_a21oi_1 _2995_ (.A1(_1780_),
    .A2(net14),
    .Y(\g.g_y[1].g_x[3].t.in_lb ),
    .B1(_1903_));
 sg13g2_nor2b_1 _2996_ (.A(\g.g_y[1].g_x[4].t.r_h ),
    .B_N(net58),
    .Y(_0118_));
 sg13g2_o21ai_1 _2997_ (.B1(_0118_),
    .Y(_0119_),
    .A1(_2056_),
    .A2(_2070_));
 sg13g2_and2_1 _2998_ (.A(\g.g_y[1].g_x[4].t.r_h ),
    .B(net58),
    .X(_0120_));
 sg13g2_nand2_1 _2999_ (.Y(_0121_),
    .A(_2079_),
    .B(_0120_));
 sg13g2_nor2_1 _3000_ (.A(_2048_),
    .B(net58),
    .Y(_0122_));
 sg13g2_nor2_1 _3001_ (.A(\g.g_y[1].g_x[4].t.r_h ),
    .B(net58),
    .Y(_0123_));
 sg13g2_a22oi_1 _3002_ (.Y(_0124_),
    .B1(_0123_),
    .B2(\g.g_y[1].g_x[4].t.out_sc ),
    .A2(_0122_),
    .A1(_2052_));
 sg13g2_nand4_1 _3003_ (.B(_0119_),
    .C(_0121_),
    .A(_1909_),
    .Y(_0125_),
    .D(_0124_));
 sg13g2_o21ai_1 _3004_ (.B1(_0051_),
    .Y(_0126_),
    .A1(_1917_),
    .A2(_1931_));
 sg13g2_nor3_1 _3005_ (.A(_1937_),
    .B(net63),
    .C(_1934_),
    .Y(_0127_));
 sg13g2_a221oi_1 _3006_ (.B2(_1916_),
    .C1(_0127_),
    .B1(_0052_),
    .A1(_1942_),
    .Y(_0128_),
    .A2(_0049_));
 sg13g2_nand3_1 _3007_ (.B(_0126_),
    .C(_0128_),
    .A(_1910_),
    .Y(_0129_));
 sg13g2_and2_1 _3008_ (.A(_0125_),
    .B(_0129_),
    .X(_0130_));
 sg13g2_or3_1 _3009_ (.A(net62),
    .B(_1994_),
    .C(_2005_),
    .X(_0131_));
 sg13g2_buf_1 _3010_ (.A(_0131_),
    .X(_0132_));
 sg13g2_nand2b_1 _3011_ (.Y(_0133_),
    .B(net62),
    .A_N(\g.g_y[0].g_x[3].t.out_sc ));
 sg13g2_and2_1 _3012_ (.A(_1995_),
    .B(_0133_),
    .X(_0134_));
 sg13g2_mux2_1 _3013_ (.A0(_2041_),
    .A1(_2011_),
    .S(net62),
    .X(_0135_));
 sg13g2_buf_1 _3014_ (.A(_0135_),
    .X(_0136_));
 sg13g2_inv_1 _3015_ (.Y(_0137_),
    .A(_1995_));
 sg13g2_a221oi_1 _3016_ (.B2(_0137_),
    .C1(_2001_),
    .B1(_0136_),
    .A1(_0132_),
    .Y(_0138_),
    .A2(_0134_));
 sg13g2_buf_2 _3017_ (.A(\g.g_y[2].g_x[3].t.r_d ),
    .X(_0139_));
 sg13g2_buf_2 _3018_ (.A(\g.g_y[2].g_x[4].t.r_h ),
    .X(_0140_));
 sg13g2_mux2_1 _3019_ (.A0(\g.g_y[2].g_x[4].t.out_sc ),
    .A1(\g.g_y[2].g_x[4].t.r_gnl ),
    .S(_2061_),
    .X(_0141_));
 sg13g2_nand2b_1 _3020_ (.Y(_0142_),
    .B(_0140_),
    .A_N(_2066_));
 sg13g2_o21ai_1 _3021_ (.B1(_0142_),
    .Y(_0143_),
    .A1(_0140_),
    .A2(_0141_));
 sg13g2_or2_1 _3022_ (.X(_0144_),
    .B(_0079_),
    .A(_1923_));
 sg13g2_o21ai_1 _3023_ (.B1(_0144_),
    .Y(_0145_),
    .A1(_0080_),
    .A2(_0078_));
 sg13g2_buf_1 _3024_ (.A(\g.g_y[2].g_x[3].t.r_h ),
    .X(_0146_));
 sg13g2_mux2_1 _3025_ (.A0(_0143_),
    .A1(_0145_),
    .S(_0146_),
    .X(_0147_));
 sg13g2_buf_1 _3026_ (.A(_0147_),
    .X(_0148_));
 sg13g2_buf_2 _3027_ (.A(\g.g_y[3].g_x[3].t.r_v ),
    .X(_0149_));
 sg13g2_buf_2 _3028_ (.A(\g.g_y[3].g_x[3].t.r_d ),
    .X(_0150_));
 sg13g2_mux2_1 _3029_ (.A0(\g.g_y[3].g_x[3].t.r_gnl ),
    .A1(\g.g_y[3].g_x[3].t.out_sc ),
    .S(_0150_),
    .X(_0151_));
 sg13g2_buf_1 _3030_ (.A(\g.g_y[3].g_x[3].t.r_ghl ),
    .X(_0152_));
 sg13g2_nand2b_1 _3031_ (.Y(_0153_),
    .B(_0149_),
    .A_N(_0152_));
 sg13g2_o21ai_1 _3032_ (.B1(_0153_),
    .Y(_0154_),
    .A1(_0149_),
    .A2(_0151_));
 sg13g2_or3_1 _3033_ (.A(_0139_),
    .B(_0148_),
    .C(_0154_),
    .X(_0155_));
 sg13g2_buf_1 _3034_ (.A(\g.g_y[2].g_x[3].t.r_v ),
    .X(_0156_));
 sg13g2_inv_1 _3035_ (.Y(_0157_),
    .A(_0139_));
 sg13g2_nor2_1 _3036_ (.A(_0157_),
    .B(\g.g_y[2].g_x[3].t.out_sc ),
    .Y(_0158_));
 sg13g2_nor2_1 _3037_ (.A(_0156_),
    .B(_0158_),
    .Y(_0159_));
 sg13g2_mux2_1 _3038_ (.A0(_0145_),
    .A1(_0143_),
    .S(_0146_),
    .X(_0160_));
 sg13g2_nand2_1 _3039_ (.Y(_0161_),
    .A(_0157_),
    .B(_0160_));
 sg13g2_inv_1 _3040_ (.Y(_0162_),
    .A(_0156_));
 sg13g2_a21oi_1 _3041_ (.A1(_0139_),
    .A2(_0154_),
    .Y(_0163_),
    .B1(_0162_));
 sg13g2_a221oi_1 _3042_ (.B2(_0163_),
    .C1(_2002_),
    .B1(_0161_),
    .A1(_0155_),
    .Y(_0164_),
    .A2(_0159_));
 sg13g2_nor2_1 _3043_ (.A(_0138_),
    .B(_0164_),
    .Y(_0165_));
 sg13g2_mux2_1 _3044_ (.A0(_0130_),
    .A1(_0165_),
    .S(_1906_),
    .X(\g.g_y[1].g_x[3].t.w_dh ));
 sg13g2_nand4_1 _3045_ (.B(_0119_),
    .C(_0121_),
    .A(_1910_),
    .Y(_0166_),
    .D(_0124_));
 sg13g2_nand3_1 _3046_ (.B(_0126_),
    .C(_0128_),
    .A(_1909_),
    .Y(_0167_));
 sg13g2_a22oi_1 _3047_ (.Y(_0168_),
    .B1(_0161_),
    .B2(_0163_),
    .A2(_0159_),
    .A1(_0155_));
 sg13g2_a221oi_1 _3048_ (.B2(_0137_),
    .C1(_2002_),
    .B1(_0136_),
    .A1(_0132_),
    .Y(_0169_),
    .A2(_0134_));
 sg13g2_a21oi_1 _3049_ (.A1(_2002_),
    .A2(_0168_),
    .Y(_0170_),
    .B1(_0169_));
 sg13g2_nand3_1 _3050_ (.B(_0167_),
    .C(_0170_),
    .A(_0166_),
    .Y(\g.g_y[1].g_x[3].t.w_na ));
 sg13g2_nand2_1 _3051_ (.Y(_0171_),
    .A(\g.g_y[1].g_x[2].t.out_sc ),
    .B(net47));
 sg13g2_or4_1 _3052_ (.A(_1906_),
    .B(net74),
    .C(_0138_),
    .D(_0164_),
    .X(_0172_));
 sg13g2_nand4_1 _3053_ (.B(net73),
    .C(_0125_),
    .A(_1906_),
    .Y(_0173_),
    .D(_0129_));
 sg13g2_nand3_1 _3054_ (.B(_0172_),
    .C(_0173_),
    .A(_0171_),
    .Y(\g.g_y[1].g_x[3].t.w_si ));
 sg13g2_nor2b_1 _3055_ (.A(net58),
    .B_N(_2079_),
    .Y(_0174_));
 sg13g2_a21oi_1 _3056_ (.A1(_2047_),
    .A2(_2076_),
    .Y(_0175_),
    .B1(_0174_));
 sg13g2_nand2_1 _3057_ (.Y(_0176_),
    .A(\g.g_y[1].g_x[3].t.out_sc ),
    .B(net52));
 sg13g2_o21ai_1 _3058_ (.B1(_0176_),
    .Y(\g.g_y[1].g_x[4].t.w_si ),
    .A1(net60),
    .A2(_0175_));
 sg13g2_inv_1 _3059_ (.Y(_0177_),
    .A(_2049_));
 sg13g2_buf_2 _3060_ (.A(\g.g_y[2].g_x[5].t.r_d ),
    .X(_0178_));
 sg13g2_buf_2 _3061_ (.A(\g.g_y[2].g_x[5].t.r_h ),
    .X(_0179_));
 sg13g2_mux2_1 _3062_ (.A0(_2066_),
    .A1(_0141_),
    .S(_0140_),
    .X(_0180_));
 sg13g2_buf_1 _3063_ (.A(_0180_),
    .X(_0181_));
 sg13g2_mux2_1 _3064_ (.A0(\g.g_y[2].g_x[6].t.out_sc ),
    .A1(\g.g_y[2].g_x[6].t.r_gnl ),
    .S(_2235_),
    .X(_0182_));
 sg13g2_buf_2 _3065_ (.A(\g.g_y[2].g_x[6].t.r_h ),
    .X(_0183_));
 sg13g2_inv_1 _3066_ (.Y(_0184_),
    .A(_0183_));
 sg13g2_nand2b_1 _3067_ (.Y(_0185_),
    .B(_0184_),
    .A_N(_0182_));
 sg13g2_inv_2 _3068_ (.Y(_0186_),
    .A(_0179_));
 sg13g2_nand2b_1 _3069_ (.Y(_0187_),
    .B(_0183_),
    .A_N(_2241_));
 sg13g2_and2_1 _3070_ (.A(_0186_),
    .B(_0187_),
    .X(_0188_));
 sg13g2_a22oi_1 _3071_ (.Y(_0189_),
    .B1(_0185_),
    .B2(_0188_),
    .A2(_0181_),
    .A1(_0179_));
 sg13g2_buf_1 _3072_ (.A(_0189_),
    .X(_0190_));
 sg13g2_buf_2 _3073_ (.A(\g.g_y[2].g_x[5].t.r_v ),
    .X(_0191_));
 sg13g2_mux2_1 _3074_ (.A0(\g.g_y[1].g_x[5].t.r_ghl ),
    .A1(_2126_),
    .S(_2127_),
    .X(_0192_));
 sg13g2_buf_1 _3075_ (.A(\g.g_y[3].g_x[5].t.r_v ),
    .X(_0193_));
 sg13g2_buf_8 _3076_ (.A(\g.g_y[3].g_x[5].t.r_d ),
    .X(_0194_));
 sg13g2_mux2_1 _3077_ (.A0(\g.g_y[3].g_x[5].t.r_gnl ),
    .A1(\g.g_y[3].g_x[5].t.out_sc ),
    .S(_0194_),
    .X(_0195_));
 sg13g2_or2_1 _3078_ (.X(_0196_),
    .B(_0195_),
    .A(net46));
 sg13g2_inv_1 _3079_ (.Y(_0197_),
    .A(_0191_));
 sg13g2_buf_1 _3080_ (.A(\g.g_y[3].g_x[5].t.r_ghl ),
    .X(_0198_));
 sg13g2_nand2b_1 _3081_ (.Y(_0199_),
    .B(net46),
    .A_N(_0198_));
 sg13g2_and2_1 _3082_ (.A(_0197_),
    .B(_0199_),
    .X(_0200_));
 sg13g2_a22oi_1 _3083_ (.Y(_0201_),
    .B1(_0196_),
    .B2(_0200_),
    .A2(_0192_),
    .A1(_0191_));
 sg13g2_buf_1 _3084_ (.A(_0201_),
    .X(_0202_));
 sg13g2_or3_1 _3085_ (.A(_0178_),
    .B(_0190_),
    .C(_0202_),
    .X(_0203_));
 sg13g2_buf_1 _3086_ (.A(_0203_),
    .X(_0204_));
 sg13g2_inv_1 _3087_ (.Y(_0205_),
    .A(_0178_));
 sg13g2_nor2_1 _3088_ (.A(_0205_),
    .B(\g.g_y[2].g_x[5].t.out_sc ),
    .Y(_0206_));
 sg13g2_nor2_1 _3089_ (.A(_0191_),
    .B(_0206_),
    .Y(_0207_));
 sg13g2_and2_1 _3090_ (.A(_0191_),
    .B(_0199_),
    .X(_0208_));
 sg13g2_a221oi_1 _3091_ (.B2(_0208_),
    .C1(_0205_),
    .B1(_0196_),
    .A1(_0197_),
    .Y(_0209_),
    .A2(_0192_));
 sg13g2_and2_1 _3092_ (.A(_0179_),
    .B(_0187_),
    .X(_0210_));
 sg13g2_a221oi_1 _3093_ (.B2(_0210_),
    .C1(_0178_),
    .B1(_0185_),
    .A1(_0186_),
    .Y(_0211_),
    .A2(_0181_));
 sg13g2_nor2_1 _3094_ (.A(_0209_),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_a221oi_1 _3095_ (.B2(_0191_),
    .C1(_2128_),
    .B1(_0212_),
    .A1(_0204_),
    .Y(_0213_),
    .A2(_0207_));
 sg13g2_mux2_1 _3096_ (.A0(_2093_),
    .A1(_2133_),
    .S(_2131_),
    .X(_0214_));
 sg13g2_mux2_1 _3097_ (.A0(_2130_),
    .A1(_0214_),
    .S(net54),
    .X(_0215_));
 sg13g2_mux2_1 _3098_ (.A0(_2144_),
    .A1(_2210_),
    .S(_2146_),
    .X(_0216_));
 sg13g2_nand3_1 _3099_ (.B(_0215_),
    .C(_0216_),
    .A(_2151_),
    .Y(_0217_));
 sg13g2_nand2b_1 _3100_ (.Y(_0218_),
    .B(net53),
    .A_N(\g.g_y[0].g_x[5].t.out_sc ));
 sg13g2_and2_1 _3101_ (.A(net54),
    .B(_0218_),
    .X(_0219_));
 sg13g2_a221oi_1 _3102_ (.B2(_2171_),
    .C1(net53),
    .B1(_2170_),
    .A1(_2146_),
    .Y(_0220_),
    .A2(_2144_));
 sg13g2_nor2_1 _3103_ (.A(_2153_),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_a221oi_1 _3104_ (.B2(_2125_),
    .C1(_2127_),
    .B1(_0221_),
    .A1(_0217_),
    .Y(_0222_),
    .A2(_0219_));
 sg13g2_nor3_1 _3105_ (.A(_0177_),
    .B(_0213_),
    .C(_0222_),
    .Y(_0223_));
 sg13g2_nor2_1 _3106_ (.A(_2220_),
    .B(_2251_),
    .Y(_0224_));
 sg13g2_o21ai_1 _3107_ (.B1(_0224_),
    .Y(_0225_),
    .A1(_2231_),
    .A2(_2245_));
 sg13g2_mux2_1 _3108_ (.A0(_2241_),
    .A1(_2237_),
    .S(_2239_),
    .X(_0226_));
 sg13g2_mux2_1 _3109_ (.A0(_2234_),
    .A1(_0226_),
    .S(_2218_),
    .X(_0227_));
 sg13g2_nor2_1 _3110_ (.A(_2227_),
    .B(_2251_),
    .Y(_0228_));
 sg13g2_nand2_1 _3111_ (.Y(_0229_),
    .A(_0227_),
    .B(_0228_));
 sg13g2_and2_1 _3112_ (.A(_2226_),
    .B(_2228_),
    .X(_0230_));
 sg13g2_nor2_1 _3113_ (.A(_2227_),
    .B(_2219_),
    .Y(_0231_));
 sg13g2_nor2_1 _3114_ (.A(_2220_),
    .B(_2219_),
    .Y(_0232_));
 sg13g2_a22oi_1 _3115_ (.Y(_0233_),
    .B1(_0232_),
    .B2(\g.g_y[1].g_x[6].t.out_sc ),
    .A2(_0231_),
    .A1(_0230_));
 sg13g2_nand4_1 _3116_ (.B(_0225_),
    .C(_0229_),
    .A(\g.g_y[1].g_x[5].t.r_h ),
    .Y(_0234_),
    .D(_0233_));
 sg13g2_o21ai_1 _3117_ (.B1(_0120_),
    .Y(_0235_),
    .A1(_2056_),
    .A2(_2070_));
 sg13g2_and2_1 _3118_ (.A(_2075_),
    .B(_0123_),
    .X(_0236_));
 sg13g2_a221oi_1 _3119_ (.B2(\g.g_y[1].g_x[4].t.out_sc ),
    .C1(_0236_),
    .B1(_0122_),
    .A1(_2079_),
    .Y(_0237_),
    .A2(_0118_));
 sg13g2_nand3_1 _3120_ (.B(_0235_),
    .C(_0237_),
    .A(_2051_),
    .Y(_0238_));
 sg13g2_nand3_1 _3121_ (.B(_0234_),
    .C(_0238_),
    .A(_0177_),
    .Y(_0239_));
 sg13g2_nand2b_1 _3122_ (.Y(\g.g_y[1].g_x[5].t.w_dh ),
    .B(_0239_),
    .A_N(_0223_));
 sg13g2_nand4_1 _3123_ (.B(_0225_),
    .C(_0229_),
    .A(_2051_),
    .Y(_0240_),
    .D(_0233_));
 sg13g2_nand3_1 _3124_ (.B(_0235_),
    .C(_0237_),
    .A(\g.g_y[1].g_x[5].t.r_h ),
    .Y(_0241_));
 sg13g2_a22oi_1 _3125_ (.Y(_0242_),
    .B1(_0221_),
    .B2(_2125_),
    .A2(_0219_),
    .A1(_0217_));
 sg13g2_a221oi_1 _3126_ (.B2(_0191_),
    .C1(_2127_),
    .B1(_0212_),
    .A1(_0204_),
    .Y(_0243_),
    .A2(_0207_));
 sg13g2_a21oi_1 _3127_ (.A1(_2127_),
    .A2(_0242_),
    .Y(_0244_),
    .B1(_0243_));
 sg13g2_nand3_1 _3128_ (.B(_0241_),
    .C(_0244_),
    .A(_0240_),
    .Y(\g.g_y[1].g_x[5].t.w_na ));
 sg13g2_or4_1 _3129_ (.A(_2049_),
    .B(_2034_),
    .C(_0213_),
    .D(_0222_),
    .X(_0245_));
 sg13g2_buf_1 _3130_ (.A(_1901_),
    .X(_0246_));
 sg13g2_nand4_1 _3131_ (.B(net45),
    .C(_0234_),
    .A(_2049_),
    .Y(_0247_),
    .D(_0238_));
 sg13g2_nand2_1 _3132_ (.Y(_0248_),
    .A(\g.g_y[1].g_x[4].t.out_sc ),
    .B(net61));
 sg13g2_nand3_1 _3133_ (.B(_0247_),
    .C(_0248_),
    .A(_0245_),
    .Y(\g.g_y[1].g_x[5].t.w_si ));
 sg13g2_nand2_1 _3134_ (.Y(_0249_),
    .A(_2227_),
    .B(_2222_));
 sg13g2_nand2_1 _3135_ (.Y(_0250_),
    .A(_2226_),
    .B(_2247_));
 sg13g2_a21oi_1 _3136_ (.A1(_0249_),
    .A2(_0250_),
    .Y(_0251_),
    .B1(_2251_));
 sg13g2_a21oi_1 _3137_ (.A1(_2251_),
    .A2(_0227_),
    .Y(_0252_),
    .B1(_0251_));
 sg13g2_nand2_1 _3138_ (.Y(_0253_),
    .A(\g.g_y[1].g_x[5].t.out_sc ),
    .B(net52));
 sg13g2_o21ai_1 _3139_ (.B1(_0253_),
    .Y(\g.g_y[1].g_x[6].t.w_si ),
    .A1(net60),
    .A2(_0252_));
 sg13g2_mux2_1 _3140_ (.A0(_2188_),
    .A1(_2224_),
    .S(_2223_),
    .X(\g.g_y[1].g_x[7].t.out_r ));
 sg13g2_nand2_1 _3141_ (.Y(_0254_),
    .A(_2195_),
    .B(_2187_));
 sg13g2_nor4_1 _3142_ (.A(_2196_),
    .B(_2199_),
    .C(_2182_),
    .D(_0254_),
    .Y(_0255_));
 sg13g2_nor3_1 _3143_ (.A(_2195_),
    .B(net28),
    .C(_2206_),
    .Y(_0256_));
 sg13g2_nand2_1 _3144_ (.Y(_0257_),
    .A(_2196_),
    .B(_2198_));
 sg13g2_and2_1 _3145_ (.A(_2195_),
    .B(_2198_),
    .X(_0258_));
 sg13g2_nand2b_1 _3146_ (.Y(_0259_),
    .B(_0258_),
    .A_N(_2201_));
 sg13g2_o21ai_1 _3147_ (.B1(_0259_),
    .Y(_0260_),
    .A1(_2187_),
    .A2(_0257_));
 sg13g2_nor4_1 _3148_ (.A(_2192_),
    .B(_0255_),
    .C(_0256_),
    .D(_0260_),
    .Y(_0261_));
 sg13g2_buf_2 _3149_ (.A(\g.g_y[2].g_x[7].t.r_h ),
    .X(_0262_));
 sg13g2_mux2_1 _3150_ (.A0(_2241_),
    .A1(_0182_),
    .S(_0183_),
    .X(_0263_));
 sg13g2_inv_1 _3151_ (.Y(_0264_),
    .A(_0076_));
 sg13g2_nand2b_1 _3152_ (.Y(_0265_),
    .B(_0264_),
    .A_N(_0075_));
 sg13g2_inv_1 _3153_ (.Y(_0266_),
    .A(_0262_));
 sg13g2_nand2b_1 _3154_ (.Y(_0267_),
    .B(_0076_),
    .A_N(_1836_));
 sg13g2_and2_1 _3155_ (.A(_0266_),
    .B(_0267_),
    .X(_0268_));
 sg13g2_a22oi_1 _3156_ (.Y(_0269_),
    .B1(_0265_),
    .B2(_0268_),
    .A2(_0263_),
    .A1(_0262_));
 sg13g2_buf_2 _3157_ (.A(\g.g_y[3].g_x[7].t.r_v ),
    .X(_0270_));
 sg13g2_buf_8 _3158_ (.A(\g.g_y[3].g_x[7].t.r_d ),
    .X(_0271_));
 sg13g2_mux2_1 _3159_ (.A0(\g.g_y[3].g_x[7].t.r_gnl ),
    .A1(\g.g_y[3].g_x[7].t.out_sc ),
    .S(_0271_),
    .X(_0272_));
 sg13g2_buf_1 _3160_ (.A(_0272_),
    .X(_0273_));
 sg13g2_nand2b_1 _3161_ (.Y(_0274_),
    .B(_0270_),
    .A_N(\g.g_y[3].g_x[7].t.r_ghl ));
 sg13g2_o21ai_1 _3162_ (.B1(_0274_),
    .Y(_0275_),
    .A1(_0270_),
    .A2(_0273_));
 sg13g2_buf_1 _3163_ (.A(\g.g_y[2].g_x[7].t.r_d ),
    .X(_0276_));
 sg13g2_inv_1 _3164_ (.Y(_0277_),
    .A(_0276_));
 sg13g2_nand2b_1 _3165_ (.Y(_0278_),
    .B(_0277_),
    .A_N(_0275_));
 sg13g2_buf_1 _3166_ (.A(\g.g_y[2].g_x[7].t.r_v ),
    .X(_0279_));
 sg13g2_inv_1 _3167_ (.Y(_0280_),
    .A(_0279_));
 sg13g2_nand2b_1 _3168_ (.Y(_0281_),
    .B(_0276_),
    .A_N(\g.g_y[2].g_x[7].t.out_sc ));
 sg13g2_and2_1 _3169_ (.A(_0280_),
    .B(_0281_),
    .X(_0282_));
 sg13g2_o21ai_1 _3170_ (.B1(_0282_),
    .Y(_0283_),
    .A1(_0269_),
    .A2(_0278_));
 sg13g2_and2_1 _3171_ (.A(_0262_),
    .B(_0267_),
    .X(_0284_));
 sg13g2_a221oi_1 _3172_ (.B2(_0284_),
    .C1(_0276_),
    .B1(_0265_),
    .A1(_0266_),
    .Y(_0285_),
    .A2(_0263_));
 sg13g2_buf_1 _3173_ (.A(_0285_),
    .X(_0286_));
 sg13g2_a21oi_1 _3174_ (.A1(_0276_),
    .A2(_0275_),
    .Y(_0287_),
    .B1(_0280_));
 sg13g2_nand2b_1 _3175_ (.Y(_0288_),
    .B(_0287_),
    .A_N(_0286_));
 sg13g2_a21oi_1 _3176_ (.A1(_0283_),
    .A2(_0288_),
    .Y(_0289_),
    .B1(_2193_));
 sg13g2_o21ai_1 _3177_ (.B1(_2189_),
    .Y(_0290_),
    .A1(_0261_),
    .A2(_0289_));
 sg13g2_and2_1 _3178_ (.A(net29),
    .B(_1827_),
    .X(_0291_));
 sg13g2_o21ai_1 _3179_ (.B1(_1845_),
    .Y(_0292_),
    .A1(net29),
    .A2(\g.g_y[1].g_x[0].t.out_sc ));
 sg13g2_a21o_1 _3180_ (.A2(_0291_),
    .A1(_0060_),
    .B1(_0292_),
    .X(_0293_));
 sg13g2_o21ai_1 _3181_ (.B1(_1822_),
    .Y(_0294_),
    .A1(net29),
    .A2(_1827_));
 sg13g2_a21o_1 _3182_ (.A2(_0044_),
    .A1(net29),
    .B1(_0294_),
    .X(_0295_));
 sg13g2_nand3_1 _3183_ (.B(_0293_),
    .C(_0295_),
    .A(_2223_),
    .Y(_0296_));
 sg13g2_o21ai_1 _3184_ (.B1(_0228_),
    .Y(_0297_),
    .A1(_2231_),
    .A2(_2245_));
 sg13g2_and2_1 _3185_ (.A(_2222_),
    .B(_0232_),
    .X(_0298_));
 sg13g2_a221oi_1 _3186_ (.B2(\g.g_y[1].g_x[6].t.out_sc ),
    .C1(_0298_),
    .B1(_0231_),
    .A1(_0227_),
    .Y(_0299_),
    .A2(_0224_));
 sg13g2_nand3b_1 _3187_ (.B(_0297_),
    .C(_0299_),
    .Y(_0300_),
    .A_N(_2223_));
 sg13g2_nand3b_1 _3188_ (.B(_0296_),
    .C(_0300_),
    .Y(_0301_),
    .A_N(_2189_));
 sg13g2_nand2_1 _3189_ (.Y(\g.g_y[1].g_x[7].t.w_dh ),
    .A(_0290_),
    .B(_0301_));
 sg13g2_nor4_1 _3190_ (.A(_2193_),
    .B(_0255_),
    .C(_0256_),
    .D(_0260_),
    .Y(_0302_));
 sg13g2_a21oi_1 _3191_ (.A1(_0283_),
    .A2(_0288_),
    .Y(_0303_),
    .B1(_2192_));
 sg13g2_nand2_1 _3192_ (.Y(_0304_),
    .A(_0293_),
    .B(_0295_));
 sg13g2_nand2_1 _3193_ (.Y(_0305_),
    .A(_0297_),
    .B(_0299_));
 sg13g2_mux2_1 _3194_ (.A0(_0304_),
    .A1(_0305_),
    .S(_2223_),
    .X(_0306_));
 sg13g2_o21ai_1 _3195_ (.B1(_0306_),
    .Y(\g.g_y[1].g_x[7].t.w_na ),
    .A1(_0302_),
    .A2(_0303_));
 sg13g2_nand2_1 _3196_ (.Y(_0307_),
    .A(\g.g_y[1].g_x[6].t.out_sc ),
    .B(net47));
 sg13g2_nand4_1 _3197_ (.B(net45),
    .C(_0296_),
    .A(_2189_),
    .Y(_0308_),
    .D(_0300_));
 sg13g2_nor2_1 _3198_ (.A(_2189_),
    .B(net82),
    .Y(_0309_));
 sg13g2_o21ai_1 _3199_ (.B1(_0309_),
    .Y(_0310_),
    .A1(_0261_),
    .A2(_0289_));
 sg13g2_nand3_1 _3200_ (.B(_0308_),
    .C(_0310_),
    .A(_0307_),
    .Y(\g.g_y[1].g_x[7].t.w_si ));
 sg13g2_inv_1 _3201_ (.Y(_0311_),
    .A(\g.g_y[3].g_x[0].t.r_h ));
 sg13g2_buf_2 _3202_ (.A(\g.g_y[3].g_x[1].t.r_h ),
    .X(_0312_));
 sg13g2_mux2_1 _3203_ (.A0(\g.g_y[3].g_x[1].t.out_sc ),
    .A1(\g.g_y[3].g_x[1].t.r_gnl ),
    .S(_0088_),
    .X(_0313_));
 sg13g2_nand2b_1 _3204_ (.Y(_0314_),
    .B(_0312_),
    .A_N(\g.g_y[3].g_x[1].t.r_ghl ));
 sg13g2_o21ai_1 _3205_ (.B1(_0314_),
    .Y(_0315_),
    .A1(_0312_),
    .A2(_0313_));
 sg13g2_buf_1 _3206_ (.A(_0315_),
    .X(_0316_));
 sg13g2_buf_2 _3207_ (.A(\g.g_y[3].g_x[0].t.r_d ),
    .X(_0317_));
 sg13g2_nor2b_1 _3208_ (.A(\g.g_y[3].g_x[0].t.r_h ),
    .B_N(net4),
    .Y(_0318_));
 sg13g2_nor2_1 _3209_ (.A(_0317_),
    .B(_0318_),
    .Y(_0319_));
 sg13g2_o21ai_1 _3210_ (.B1(_0319_),
    .Y(_0320_),
    .A1(_0311_),
    .A2(_0316_));
 sg13g2_buf_2 _3211_ (.A(\g.g_y[4].g_x[0].t.r_v ),
    .X(_0321_));
 sg13g2_buf_8 _3212_ (.A(\g.g_y[4].g_x[0].t.r_d ),
    .X(_0322_));
 sg13g2_mux2_1 _3213_ (.A0(\g.g_y[4].g_x[0].t.r_gnl ),
    .A1(\g.g_y[4].g_x[0].t.out_sc ),
    .S(_0322_),
    .X(_0323_));
 sg13g2_buf_1 _3214_ (.A(_0323_),
    .X(_0324_));
 sg13g2_buf_1 _3215_ (.A(\g.g_y[4].g_x[0].t.r_ghl ),
    .X(_0325_));
 sg13g2_nand2b_1 _3216_ (.Y(_0326_),
    .B(_0321_),
    .A_N(_0325_));
 sg13g2_o21ai_1 _3217_ (.B1(_0326_),
    .Y(_0327_),
    .A1(_0321_),
    .A2(_0324_));
 sg13g2_buf_2 _3218_ (.A(_0327_),
    .X(_0328_));
 sg13g2_buf_1 _3219_ (.A(\g.g_y[3].g_x[0].t.r_v ),
    .X(_0329_));
 sg13g2_inv_1 _3220_ (.Y(_0330_),
    .A(_0329_));
 sg13g2_a21oi_1 _3221_ (.A1(_0317_),
    .A2(_0328_),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_nand2_1 _3222_ (.Y(_0332_),
    .A(_0320_),
    .B(_0331_));
 sg13g2_inv_1 _3223_ (.Y(_0333_),
    .A(net4));
 sg13g2_mux2_1 _3224_ (.A0(_0333_),
    .A1(_0316_),
    .S(_0311_),
    .X(_0334_));
 sg13g2_inv_2 _3225_ (.Y(_0335_),
    .A(_0317_));
 sg13g2_nand2b_1 _3226_ (.Y(_0336_),
    .B(_0335_),
    .A_N(_0328_));
 sg13g2_nand2b_1 _3227_ (.Y(_0337_),
    .B(_0317_),
    .A_N(\g.g_y[3].g_x[0].t.out_sc ));
 sg13g2_and2_1 _3228_ (.A(_0330_),
    .B(_0337_),
    .X(_0338_));
 sg13g2_o21ai_1 _3229_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_0334_),
    .A2(_0336_));
 sg13g2_nand3_1 _3230_ (.B(_0332_),
    .C(_0339_),
    .A(_1833_),
    .Y(_0340_));
 sg13g2_nand2_1 _3231_ (.Y(_0341_),
    .A(_1832_),
    .B(_0043_));
 sg13g2_nand3b_1 _3232_ (.B(_1831_),
    .C(_0341_),
    .Y(_0342_),
    .A_N(_1821_));
 sg13g2_and2_1 _3233_ (.A(_1821_),
    .B(_1848_),
    .X(_0343_));
 sg13g2_o21ai_1 _3234_ (.B1(_0343_),
    .Y(_0344_),
    .A1(_1847_),
    .A2(_0043_));
 sg13g2_nand3_1 _3235_ (.B(_0342_),
    .C(_0344_),
    .A(_0057_),
    .Y(_0345_));
 sg13g2_and3_1 _3236_ (.X(_0346_),
    .A(_1834_),
    .B(_0340_),
    .C(_0345_));
 sg13g2_or2_1 _3237_ (.X(_0347_),
    .B(\g.g_y[1].g_x[1].t.r_v ),
    .A(_1801_));
 sg13g2_o21ai_1 _3238_ (.B1(_0347_),
    .Y(_0348_),
    .A1(_1804_),
    .A2(_1803_));
 sg13g2_buf_1 _3239_ (.A(_0348_),
    .X(_0349_));
 sg13g2_mux2_1 _3240_ (.A0(_0091_),
    .A1(_0349_),
    .S(_0095_),
    .X(_0350_));
 sg13g2_nand3b_1 _3241_ (.B(net27),
    .C(_0084_),
    .Y(_0351_),
    .A_N(_0350_));
 sg13g2_buf_1 _3242_ (.A(_0351_),
    .X(_0352_));
 sg13g2_nor2_1 _3243_ (.A(_0085_),
    .B(\g.g_y[2].g_x[1].t.out_sc ),
    .Y(_0353_));
 sg13g2_nor2_1 _3244_ (.A(_0082_),
    .B(_0353_),
    .Y(_0354_));
 sg13g2_inv_1 _3245_ (.Y(_0355_),
    .A(_0095_));
 sg13g2_mux2_1 _3246_ (.A0(_0091_),
    .A1(_0349_),
    .S(_0355_),
    .X(_0356_));
 sg13g2_a21oi_2 _3247_ (.B1(_0099_),
    .Y(_0357_),
    .A2(_0356_),
    .A1(net27));
 sg13g2_a221oi_1 _3248_ (.B2(_0082_),
    .C1(_0264_),
    .B1(_0357_),
    .A1(_0352_),
    .Y(_0358_),
    .A2(_0354_));
 sg13g2_nor2_1 _3249_ (.A(_0076_),
    .B(net3),
    .Y(_0359_));
 sg13g2_nor3_1 _3250_ (.A(_1834_),
    .B(_0358_),
    .C(_0359_),
    .Y(_0360_));
 sg13g2_or2_1 _3251_ (.X(\g.g_y[2].g_x[0].t.w_dh ),
    .B(_0360_),
    .A(_0346_));
 sg13g2_a21oi_1 _3252_ (.A1(_0342_),
    .A2(_0344_),
    .Y(_0361_),
    .B1(_0057_));
 sg13g2_a21oi_1 _3253_ (.A1(_0332_),
    .A2(_0339_),
    .Y(_0362_),
    .B1(_1833_));
 sg13g2_a22oi_1 _3254_ (.Y(_0363_),
    .B1(_0357_),
    .B2(_0082_),
    .A2(_0354_),
    .A1(_0352_));
 sg13g2_nand2_1 _3255_ (.Y(_0364_),
    .A(_0076_),
    .B(net3));
 sg13g2_o21ai_1 _3256_ (.B1(_0364_),
    .Y(_0365_),
    .A1(_0076_),
    .A2(_0363_));
 sg13g2_o21ai_1 _3257_ (.B1(_0365_),
    .Y(\g.g_y[2].g_x[0].t.w_na ),
    .A1(_0361_),
    .A2(_0362_));
 sg13g2_nand2_1 _3258_ (.Y(_0366_),
    .A(\g.g_y[1].g_x[7].t.out_sc ),
    .B(net47));
 sg13g2_inv_1 _3259_ (.Y(_0367_),
    .A(_1834_));
 sg13g2_or4_1 _3260_ (.A(_0367_),
    .B(net74),
    .C(_0358_),
    .D(_0359_),
    .X(_0368_));
 sg13g2_nand4_1 _3261_ (.B(net73),
    .C(_0340_),
    .A(_0367_),
    .Y(_0369_),
    .D(_0345_));
 sg13g2_nand3_1 _3262_ (.B(_0368_),
    .C(_0369_),
    .A(_0366_),
    .Y(\g.g_y[2].g_x[0].t.w_si ));
 sg13g2_a22oi_1 _3263_ (.Y(_0370_),
    .B1(_0097_),
    .B2(_0098_),
    .A2(_0077_),
    .A1(_0083_));
 sg13g2_mux2_1 _3264_ (.A0(_0356_),
    .A1(_0370_),
    .S(net27),
    .X(_0371_));
 sg13g2_nand2_1 _3265_ (.Y(_0372_),
    .A(\g.g_y[2].g_x[0].t.out_sc ),
    .B(_2175_));
 sg13g2_o21ai_1 _3266_ (.B1(_0372_),
    .Y(\g.g_y[2].g_x[1].t.w_si ),
    .A1(_2040_),
    .A2(_0371_));
 sg13g2_nor2_1 _3267_ (.A(_0083_),
    .B(_0353_),
    .Y(_0373_));
 sg13g2_a221oi_1 _3268_ (.B2(_0352_),
    .C1(_0079_),
    .B1(_0373_),
    .A1(_0083_),
    .Y(_0374_),
    .A2(_0357_));
 sg13g2_or2_1 _3269_ (.X(_0375_),
    .B(_2001_),
    .A(_1912_));
 sg13g2_o21ai_1 _3270_ (.B1(_0375_),
    .Y(_0376_),
    .A1(_2002_),
    .A2(_2000_));
 sg13g2_mux2_1 _3271_ (.A0(_0154_),
    .A1(_0376_),
    .S(_0156_),
    .X(_0377_));
 sg13g2_nor2_1 _3272_ (.A(_0146_),
    .B(_0157_),
    .Y(_0378_));
 sg13g2_o21ai_1 _3273_ (.B1(_0378_),
    .Y(_0379_),
    .A1(_0148_),
    .A2(_0377_));
 sg13g2_inv_1 _3274_ (.Y(_0380_),
    .A(_0149_));
 sg13g2_mux2_1 _3275_ (.A0(_0152_),
    .A1(_0151_),
    .S(_0380_),
    .X(_0381_));
 sg13g2_mux2_1 _3276_ (.A0(_1912_),
    .A1(_2000_),
    .S(_2001_),
    .X(_0382_));
 sg13g2_mux2_1 _3277_ (.A0(_0381_),
    .A1(_0382_),
    .S(_0162_),
    .X(_0383_));
 sg13g2_and2_1 _3278_ (.A(_0146_),
    .B(_0139_),
    .X(_0384_));
 sg13g2_nor2_1 _3279_ (.A(_0146_),
    .B(_0139_),
    .Y(_0385_));
 sg13g2_nor2b_1 _3280_ (.A(_0139_),
    .B_N(_0146_),
    .Y(_0386_));
 sg13g2_nor2b_1 _3281_ (.A(_0143_),
    .B_N(_0386_),
    .Y(_0387_));
 sg13g2_a221oi_1 _3282_ (.B2(\g.g_y[2].g_x[3].t.out_sc ),
    .C1(_0387_),
    .B1(_0385_),
    .A1(_0383_),
    .Y(_0388_),
    .A2(_0384_));
 sg13g2_nand3_1 _3283_ (.B(_0379_),
    .C(_0388_),
    .A(_0079_),
    .Y(_0389_));
 sg13g2_nor2b_1 _3284_ (.A(_0374_),
    .B_N(_0389_),
    .Y(_0390_));
 sg13g2_a21oi_1 _3285_ (.A1(_1905_),
    .A2(_1934_),
    .Y(_0391_),
    .B1(_1940_));
 sg13g2_a221oi_1 _3286_ (.B2(_1933_),
    .C1(_1920_),
    .B1(_0391_),
    .A1(_1940_),
    .Y(_0392_),
    .A2(_1944_));
 sg13g2_buf_1 _3287_ (.A(\g.g_y[3].g_x[2].t.r_d ),
    .X(_0393_));
 sg13g2_buf_1 _3288_ (.A(_0393_),
    .X(_0394_));
 sg13g2_buf_1 _3289_ (.A(\g.g_y[3].g_x[3].t.r_h ),
    .X(_0395_));
 sg13g2_mux2_1 _3290_ (.A0(\g.g_y[3].g_x[3].t.out_sc ),
    .A1(\g.g_y[3].g_x[3].t.r_gnl ),
    .S(_0150_),
    .X(_0396_));
 sg13g2_nand2b_1 _3291_ (.Y(_0397_),
    .B(_0395_),
    .A_N(_0152_));
 sg13g2_o21ai_1 _3292_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_0395_),
    .A2(_0396_));
 sg13g2_inv_1 _3293_ (.Y(_0399_),
    .A(_0312_));
 sg13g2_or2_1 _3294_ (.X(_0400_),
    .B(_0312_),
    .A(\g.g_y[3].g_x[1].t.r_ghl ));
 sg13g2_o21ai_1 _3295_ (.B1(_0400_),
    .Y(_0401_),
    .A1(_0399_),
    .A2(_0313_));
 sg13g2_buf_1 _3296_ (.A(\g.g_y[3].g_x[2].t.r_h ),
    .X(_0402_));
 sg13g2_mux2_1 _3297_ (.A0(_0398_),
    .A1(_0401_),
    .S(_0402_),
    .X(_0403_));
 sg13g2_buf_1 _3298_ (.A(_0403_),
    .X(_0404_));
 sg13g2_buf_1 _3299_ (.A(\g.g_y[4].g_x[2].t.r_d ),
    .X(_0405_));
 sg13g2_mux2_1 _3300_ (.A0(\g.g_y[4].g_x[2].t.r_gnl ),
    .A1(\g.g_y[4].g_x[2].t.out_sc ),
    .S(_0405_),
    .X(_0406_));
 sg13g2_buf_1 _3301_ (.A(_0406_),
    .X(_0407_));
 sg13g2_buf_2 _3302_ (.A(\g.g_y[4].g_x[2].t.r_v ),
    .X(_0408_));
 sg13g2_inv_1 _3303_ (.Y(_0409_),
    .A(_0408_));
 sg13g2_nand2b_1 _3304_ (.Y(_0410_),
    .B(_0409_),
    .A_N(_0407_));
 sg13g2_buf_2 _3305_ (.A(\g.g_y[4].g_x[2].t.r_ghl ),
    .X(_0411_));
 sg13g2_nand2b_1 _3306_ (.Y(_0412_),
    .B(_0408_),
    .A_N(_0411_));
 sg13g2_nand2_1 _3307_ (.Y(_0413_),
    .A(_0410_),
    .B(_0412_));
 sg13g2_or3_1 _3308_ (.A(net26),
    .B(_0404_),
    .C(_0413_),
    .X(_0414_));
 sg13g2_buf_1 _3309_ (.A(\g.g_y[3].g_x[2].t.r_v ),
    .X(_0415_));
 sg13g2_nor2b_1 _3310_ (.A(\g.g_y[3].g_x[2].t.out_sc ),
    .B_N(_0393_),
    .Y(_0416_));
 sg13g2_nor2_1 _3311_ (.A(_0415_),
    .B(_0416_),
    .Y(_0417_));
 sg13g2_mux2_1 _3312_ (.A0(_0401_),
    .A1(_0398_),
    .S(_0402_),
    .X(_0418_));
 sg13g2_nand2b_1 _3313_ (.Y(_0419_),
    .B(_0418_),
    .A_N(net26));
 sg13g2_inv_1 _3314_ (.Y(_0420_),
    .A(_0415_));
 sg13g2_a21oi_1 _3315_ (.A1(net26),
    .A2(_0413_),
    .Y(_0421_),
    .B1(_0420_));
 sg13g2_a221oi_1 _3316_ (.B2(_0421_),
    .C1(_1921_),
    .B1(_0419_),
    .A1(_0414_),
    .Y(_0422_),
    .A2(_0417_));
 sg13g2_nor2_1 _3317_ (.A(_0392_),
    .B(_0422_),
    .Y(_0423_));
 sg13g2_mux2_1 _3318_ (.A0(_0390_),
    .A1(_0423_),
    .S(_1918_),
    .X(\g.g_y[2].g_x[2].t.w_dh ));
 sg13g2_a22oi_1 _3319_ (.Y(_0424_),
    .B1(_0373_),
    .B2(_0352_),
    .A2(_0357_),
    .A1(_0083_));
 sg13g2_nand2_1 _3320_ (.Y(_0425_),
    .A(_0079_),
    .B(_0424_));
 sg13g2_nand3_1 _3321_ (.B(_0379_),
    .C(_0388_),
    .A(_0080_),
    .Y(_0426_));
 sg13g2_a22oi_1 _3322_ (.Y(_0427_),
    .B1(_0419_),
    .B2(_0421_),
    .A2(_0417_),
    .A1(_0414_));
 sg13g2_a221oi_1 _3323_ (.B2(_1933_),
    .C1(_1921_),
    .B1(_0391_),
    .A1(_1940_),
    .Y(_0428_),
    .A2(_1944_));
 sg13g2_a21oi_1 _3324_ (.A1(_1921_),
    .A2(_0427_),
    .Y(_0429_),
    .B1(_0428_));
 sg13g2_nand3_1 _3325_ (.B(_0426_),
    .C(_0429_),
    .A(_0425_),
    .Y(\g.g_y[2].g_x[2].t.w_na ));
 sg13g2_or4_1 _3326_ (.A(_1918_),
    .B(net78),
    .C(_0392_),
    .D(_0422_),
    .X(_0430_));
 sg13g2_and2_1 _3327_ (.A(_1918_),
    .B(net81),
    .X(_0431_));
 sg13g2_nand3b_1 _3328_ (.B(_0389_),
    .C(_0431_),
    .Y(_0432_),
    .A_N(_0374_));
 sg13g2_nand2_1 _3329_ (.Y(_0433_),
    .A(\g.g_y[2].g_x[1].t.out_sc ),
    .B(net61));
 sg13g2_nand3_1 _3330_ (.B(_0432_),
    .C(_0433_),
    .A(_0430_),
    .Y(\g.g_y[2].g_x[2].t.w_si ));
 sg13g2_nor2_1 _3331_ (.A(_0157_),
    .B(_0160_),
    .Y(_0434_));
 sg13g2_a21oi_1 _3332_ (.A1(_0157_),
    .A2(_0383_),
    .Y(_0435_),
    .B1(_0434_));
 sg13g2_nand2_1 _3333_ (.Y(_0436_),
    .A(\g.g_y[2].g_x[2].t.out_sc ),
    .B(net52));
 sg13g2_o21ai_1 _3334_ (.B1(_0436_),
    .Y(\g.g_y[2].g_x[3].t.w_si ),
    .A1(net60),
    .A2(_0435_));
 sg13g2_nor2_1 _3335_ (.A(_0179_),
    .B(_0205_),
    .Y(_0437_));
 sg13g2_o21ai_1 _3336_ (.B1(_0437_),
    .Y(_0438_),
    .A1(_0190_),
    .A2(_0202_));
 sg13g2_mux2_1 _3337_ (.A0(_0195_),
    .A1(_0198_),
    .S(net46),
    .X(_0439_));
 sg13g2_mux2_1 _3338_ (.A0(_0192_),
    .A1(_0439_),
    .S(_0191_),
    .X(_0440_));
 sg13g2_nand3_1 _3339_ (.B(_0178_),
    .C(_0440_),
    .A(_0179_),
    .Y(_0441_));
 sg13g2_and2_1 _3340_ (.A(_0185_),
    .B(_0187_),
    .X(_0442_));
 sg13g2_nor2_1 _3341_ (.A(_0186_),
    .B(_0178_),
    .Y(_0443_));
 sg13g2_nor2_1 _3342_ (.A(_0179_),
    .B(_0178_),
    .Y(_0444_));
 sg13g2_a22oi_1 _3343_ (.Y(_0445_),
    .B1(_0444_),
    .B2(\g.g_y[2].g_x[5].t.out_sc ),
    .A2(_0443_),
    .A1(_0442_));
 sg13g2_nand4_1 _3344_ (.B(_0438_),
    .C(_0441_),
    .A(_0140_),
    .Y(_0446_),
    .D(_0445_));
 sg13g2_inv_1 _3345_ (.Y(_0447_),
    .A(_0140_));
 sg13g2_o21ai_1 _3346_ (.B1(_0384_),
    .Y(_0448_),
    .A1(_0148_),
    .A2(_0377_));
 sg13g2_nand2_1 _3347_ (.Y(_0449_),
    .A(_0378_),
    .B(_0383_));
 sg13g2_nor2b_1 _3348_ (.A(_0145_),
    .B_N(_0385_),
    .Y(_0450_));
 sg13g2_a21oi_1 _3349_ (.A1(\g.g_y[2].g_x[3].t.out_sc ),
    .A2(_0386_),
    .Y(_0451_),
    .B1(_0450_));
 sg13g2_nand4_1 _3350_ (.B(_0448_),
    .C(_0449_),
    .A(_0447_),
    .Y(_0452_),
    .D(_0451_));
 sg13g2_nand2_1 _3351_ (.Y(_0453_),
    .A(_0446_),
    .B(_0452_));
 sg13g2_buf_1 _3352_ (.A(\g.g_y[3].g_x[4].t.r_v ),
    .X(_0454_));
 sg13g2_inv_2 _3353_ (.Y(_0455_),
    .A(net44));
 sg13g2_buf_1 _3354_ (.A(\g.g_y[3].g_x[4].t.r_d ),
    .X(_0456_));
 sg13g2_inv_2 _3355_ (.Y(_0457_),
    .A(_0456_));
 sg13g2_buf_1 _3356_ (.A(\g.g_y[3].g_x[4].t.out_sc ),
    .X(_0458_));
 sg13g2_nor2_1 _3357_ (.A(_0457_),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_nand2_1 _3358_ (.Y(_0460_),
    .A(_0455_),
    .B(_0459_));
 sg13g2_nor2_1 _3359_ (.A(net56),
    .B(net57),
    .Y(_0461_));
 sg13g2_nand2_1 _3360_ (.Y(_0462_),
    .A(net57),
    .B(_2073_));
 sg13g2_nor2_1 _3361_ (.A(net56),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_a221oi_1 _3362_ (.B2(_2081_),
    .C1(_0463_),
    .B1(_0461_),
    .A1(net56),
    .Y(_0464_),
    .A2(_0460_));
 sg13g2_nor2_1 _3363_ (.A(_2064_),
    .B(_0455_),
    .Y(_0465_));
 sg13g2_buf_1 _3364_ (.A(\g.g_y[3].g_x[4].t.r_h ),
    .X(_0466_));
 sg13g2_mux2_1 _3365_ (.A0(\g.g_y[3].g_x[5].t.out_sc ),
    .A1(\g.g_y[3].g_x[5].t.r_gnl ),
    .S(_0194_),
    .X(_0467_));
 sg13g2_buf_2 _3366_ (.A(\g.g_y[3].g_x[5].t.r_h ),
    .X(_0468_));
 sg13g2_inv_1 _3367_ (.Y(_0469_),
    .A(_0468_));
 sg13g2_mux2_1 _3368_ (.A0(_0198_),
    .A1(_0467_),
    .S(_0469_),
    .X(_0470_));
 sg13g2_buf_1 _3369_ (.A(_0470_),
    .X(_0471_));
 sg13g2_inv_1 _3370_ (.Y(_0472_),
    .A(_0395_));
 sg13g2_or2_1 _3371_ (.X(_0473_),
    .B(_0396_),
    .A(_0472_));
 sg13g2_nor2_1 _3372_ (.A(_0152_),
    .B(_0395_),
    .Y(_0474_));
 sg13g2_nor2_1 _3373_ (.A(_0466_),
    .B(_0474_),
    .Y(_0475_));
 sg13g2_a221oi_1 _3374_ (.B2(_0475_),
    .C1(_0456_),
    .B1(_0473_),
    .A1(_0466_),
    .Y(_0476_),
    .A2(_0471_));
 sg13g2_buf_8 _3375_ (.A(\g.g_y[4].g_x[4].t.r_d ),
    .X(_0477_));
 sg13g2_mux2_1 _3376_ (.A0(\g.g_y[4].g_x[4].t.r_gnl ),
    .A1(\g.g_y[4].g_x[4].t.out_sc ),
    .S(_0477_),
    .X(_0478_));
 sg13g2_buf_2 _3377_ (.A(\g.g_y[4].g_x[4].t.r_ghl ),
    .X(_0479_));
 sg13g2_buf_1 _3378_ (.A(\g.g_y[4].g_x[4].t.r_v ),
    .X(_0480_));
 sg13g2_mux2_1 _3379_ (.A0(_0478_),
    .A1(_0479_),
    .S(net43),
    .X(_0481_));
 sg13g2_nor2_1 _3380_ (.A(_0457_),
    .B(_0481_),
    .Y(_0482_));
 sg13g2_or2_1 _3381_ (.X(_0483_),
    .B(_0482_),
    .A(_0476_));
 sg13g2_nor2_1 _3382_ (.A(_2064_),
    .B(net44),
    .Y(_0484_));
 sg13g2_inv_1 _3383_ (.Y(_0485_),
    .A(_0466_));
 sg13g2_nor2_1 _3384_ (.A(_0485_),
    .B(_0474_),
    .Y(_0486_));
 sg13g2_a22oi_1 _3385_ (.Y(_0487_),
    .B1(_0473_),
    .B2(_0486_),
    .A2(_0471_),
    .A1(_0485_));
 sg13g2_buf_1 _3386_ (.A(_0487_),
    .X(_0488_));
 sg13g2_mux2_1 _3387_ (.A0(_2066_),
    .A1(_2062_),
    .S(net56),
    .X(_0489_));
 sg13g2_buf_1 _3388_ (.A(_0489_),
    .X(_0490_));
 sg13g2_nor2b_1 _3389_ (.A(_0479_),
    .B_N(net43),
    .Y(_0491_));
 sg13g2_nor2_1 _3390_ (.A(net44),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_or2_1 _3391_ (.X(_0493_),
    .B(_0478_),
    .A(net43));
 sg13g2_a22oi_1 _3392_ (.Y(_0494_),
    .B1(_0492_),
    .B2(_0493_),
    .A2(_0490_),
    .A1(net44));
 sg13g2_nor3_1 _3393_ (.A(_0456_),
    .B(_0488_),
    .C(_0494_),
    .Y(_0495_));
 sg13g2_nand2b_1 _3394_ (.Y(_0496_),
    .B(net57),
    .A_N(net58));
 sg13g2_nor4_1 _3395_ (.A(net56),
    .B(_2056_),
    .C(_2070_),
    .D(_0496_),
    .Y(_0497_));
 sg13g2_a221oi_1 _3396_ (.B2(_0495_),
    .C1(_0497_),
    .B1(_0484_),
    .A1(_0465_),
    .Y(_0498_),
    .A2(_0483_));
 sg13g2_nand3b_1 _3397_ (.B(_0498_),
    .C(_2061_),
    .Y(_0499_),
    .A_N(_0464_));
 sg13g2_o21ai_1 _3398_ (.B1(_0499_),
    .Y(\g.g_y[2].g_x[4].t.w_dh ),
    .A1(_2061_),
    .A2(_0453_));
 sg13g2_nand4_1 _3399_ (.B(_0438_),
    .C(_0441_),
    .A(_0447_),
    .Y(_0500_),
    .D(_0445_));
 sg13g2_nand4_1 _3400_ (.B(_0448_),
    .C(_0449_),
    .A(_0140_),
    .Y(_0501_),
    .D(_0451_));
 sg13g2_nor2_1 _3401_ (.A(_0455_),
    .B(_0491_),
    .Y(_0502_));
 sg13g2_a221oi_1 _3402_ (.B2(_0493_),
    .C1(_0457_),
    .B1(_0502_),
    .A1(_0455_),
    .Y(_0503_),
    .A2(_0490_));
 sg13g2_nor3_1 _3403_ (.A(_0455_),
    .B(_0476_),
    .C(_0503_),
    .Y(_0504_));
 sg13g2_nor3_1 _3404_ (.A(net44),
    .B(_0495_),
    .C(_0459_),
    .Y(_0505_));
 sg13g2_or3_1 _3405_ (.A(net56),
    .B(_0504_),
    .C(_0505_),
    .X(_0506_));
 sg13g2_nand2b_1 _3406_ (.Y(_0507_),
    .B(_2081_),
    .A_N(net57));
 sg13g2_nand2b_1 _3407_ (.Y(_0508_),
    .B(_2072_),
    .A_N(_0462_));
 sg13g2_nand3_1 _3408_ (.B(_0507_),
    .C(_0508_),
    .A(_2063_),
    .Y(_0509_));
 sg13g2_nand4_1 _3409_ (.B(_0501_),
    .C(_0506_),
    .A(_0500_),
    .Y(\g.g_y[2].g_x[4].t.w_na ),
    .D(_0509_));
 sg13g2_nand2_1 _3410_ (.Y(_0510_),
    .A(\g.g_y[2].g_x[3].t.out_sc ),
    .B(net47));
 sg13g2_nor2_1 _3411_ (.A(_2061_),
    .B(net78),
    .Y(_0511_));
 sg13g2_nand3b_1 _3412_ (.B(_0511_),
    .C(_0498_),
    .Y(_0512_),
    .A_N(_0464_));
 sg13g2_nand4_1 _3413_ (.B(net73),
    .C(_0446_),
    .A(_2061_),
    .Y(_0513_),
    .D(_0452_));
 sg13g2_nand3_1 _3414_ (.B(_0512_),
    .C(_0513_),
    .A(_0510_),
    .Y(\g.g_y[2].g_x[4].t.w_si ));
 sg13g2_nand2_1 _3415_ (.Y(_0514_),
    .A(_0186_),
    .B(_0181_));
 sg13g2_nand2_1 _3416_ (.Y(_0515_),
    .A(_0185_),
    .B(_0210_));
 sg13g2_a21oi_1 _3417_ (.A1(_0514_),
    .A2(_0515_),
    .Y(_0516_),
    .B1(_0205_));
 sg13g2_a21oi_1 _3418_ (.A1(_0205_),
    .A2(_0440_),
    .Y(_0517_),
    .B1(_0516_));
 sg13g2_nand2_1 _3419_ (.Y(_0518_),
    .A(\g.g_y[2].g_x[4].t.out_sc ),
    .B(net52));
 sg13g2_o21ai_1 _3420_ (.B1(_0518_),
    .Y(\g.g_y[2].g_x[5].t.w_si ),
    .A1(net60),
    .A2(_0517_));
 sg13g2_or2_1 _3421_ (.X(_0519_),
    .B(_0202_),
    .A(_0190_));
 sg13g2_mux4_1 _3422_ (.S0(_0186_),
    .A0(\g.g_y[2].g_x[5].t.out_sc ),
    .A1(_0181_),
    .A2(_0519_),
    .A3(_0440_),
    .S1(_0178_),
    .X(_0520_));
 sg13g2_nor2_1 _3423_ (.A(_0184_),
    .B(_0266_),
    .Y(_0521_));
 sg13g2_mux2_1 _3424_ (.A0(_2188_),
    .A1(_2191_),
    .S(_2192_),
    .X(_0522_));
 sg13g2_and2_1 _3425_ (.A(_0279_),
    .B(_0274_),
    .X(_0523_));
 sg13g2_inv_1 _3426_ (.Y(_0524_),
    .A(_0270_));
 sg13g2_nand2b_1 _3427_ (.Y(_0525_),
    .B(_0524_),
    .A_N(_0273_));
 sg13g2_a221oi_1 _3428_ (.B2(_0525_),
    .C1(_0277_),
    .B1(_0523_),
    .A1(_0280_),
    .Y(_0526_),
    .A2(_0522_));
 sg13g2_nor2_1 _3429_ (.A(_0286_),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_or2_1 _3430_ (.X(_0528_),
    .B(_2192_),
    .A(_2188_));
 sg13g2_o21ai_1 _3431_ (.B1(_0528_),
    .Y(_0529_),
    .A1(_2193_),
    .A2(_2191_));
 sg13g2_mux2_1 _3432_ (.A0(_0275_),
    .A1(_0529_),
    .S(_0279_),
    .X(_0530_));
 sg13g2_nor3_1 _3433_ (.A(_0277_),
    .B(_0269_),
    .C(_0530_),
    .Y(_0531_));
 sg13g2_nor2_1 _3434_ (.A(_0276_),
    .B(\g.g_y[2].g_x[7].t.out_sc ),
    .Y(_0532_));
 sg13g2_nor4_1 _3435_ (.A(_0184_),
    .B(_0262_),
    .C(_0531_),
    .D(_0532_),
    .Y(_0533_));
 sg13g2_a221oi_1 _3436_ (.B2(_0527_),
    .C1(_0533_),
    .B1(_0521_),
    .A1(_0184_),
    .Y(_0534_),
    .A2(_0520_));
 sg13g2_inv_1 _3437_ (.Y(_0535_),
    .A(_2235_));
 sg13g2_buf_2 _3438_ (.A(\g.g_y[3].g_x[6].t.r_d ),
    .X(_0536_));
 sg13g2_buf_2 _3439_ (.A(\g.g_y[3].g_x[7].t.r_h ),
    .X(_0537_));
 sg13g2_mux2_1 _3440_ (.A0(\g.g_y[3].g_x[7].t.out_sc ),
    .A1(\g.g_y[3].g_x[7].t.r_gnl ),
    .S(_0271_),
    .X(_0538_));
 sg13g2_or2_1 _3441_ (.X(_0539_),
    .B(_0538_),
    .A(_0537_));
 sg13g2_buf_1 _3442_ (.A(_0539_),
    .X(_0540_));
 sg13g2_buf_1 _3443_ (.A(\g.g_y[3].g_x[6].t.r_h ),
    .X(_0541_));
 sg13g2_inv_1 _3444_ (.Y(_0542_),
    .A(_0541_));
 sg13g2_nand2b_1 _3445_ (.Y(_0543_),
    .B(_0537_),
    .A_N(\g.g_y[3].g_x[7].t.r_ghl ));
 sg13g2_and2_1 _3446_ (.A(_0542_),
    .B(_0543_),
    .X(_0544_));
 sg13g2_mux2_1 _3447_ (.A0(_0198_),
    .A1(_0467_),
    .S(_0468_),
    .X(_0545_));
 sg13g2_buf_1 _3448_ (.A(_0545_),
    .X(_0546_));
 sg13g2_a22oi_1 _3449_ (.Y(_0547_),
    .B1(_0546_),
    .B2(_0541_),
    .A2(_0544_),
    .A1(_0540_));
 sg13g2_buf_2 _3450_ (.A(\g.g_y[4].g_x[6].t.r_v ),
    .X(_0548_));
 sg13g2_buf_8 _3451_ (.A(\g.g_y[4].g_x[6].t.r_d ),
    .X(_0549_));
 sg13g2_mux2_1 _3452_ (.A0(\g.g_y[4].g_x[6].t.r_gnl ),
    .A1(\g.g_y[4].g_x[6].t.out_sc ),
    .S(_0549_),
    .X(_0550_));
 sg13g2_buf_1 _3453_ (.A(\g.g_y[4].g_x[6].t.r_ghl ),
    .X(_0551_));
 sg13g2_nand2b_1 _3454_ (.Y(_0552_),
    .B(_0548_),
    .A_N(_0551_));
 sg13g2_o21ai_1 _3455_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0548_),
    .A2(_0550_));
 sg13g2_or2_1 _3456_ (.X(_0554_),
    .B(_2238_),
    .A(_2241_));
 sg13g2_o21ai_1 _3457_ (.B1(_0554_),
    .Y(_0555_),
    .A1(_2239_),
    .A2(_2237_));
 sg13g2_buf_1 _3458_ (.A(\g.g_y[3].g_x[6].t.r_v ),
    .X(_0556_));
 sg13g2_mux2_1 _3459_ (.A0(_0553_),
    .A1(_0555_),
    .S(_0556_),
    .X(_0557_));
 sg13g2_or3_1 _3460_ (.A(_0536_),
    .B(_0547_),
    .C(_0557_),
    .X(_0558_));
 sg13g2_buf_1 _3461_ (.A(_0558_),
    .X(_0559_));
 sg13g2_inv_1 _3462_ (.Y(_0560_),
    .A(_0556_));
 sg13g2_nand2b_1 _3463_ (.Y(_0561_),
    .B(_0536_),
    .A_N(\g.g_y[3].g_x[6].t.out_sc ));
 sg13g2_and2_1 _3464_ (.A(_0560_),
    .B(_0561_),
    .X(_0562_));
 sg13g2_mux2_1 _3465_ (.A0(_0553_),
    .A1(_0555_),
    .S(_0560_),
    .X(_0563_));
 sg13g2_and2_1 _3466_ (.A(_0541_),
    .B(_0543_),
    .X(_0564_));
 sg13g2_a221oi_1 _3467_ (.B2(_0540_),
    .C1(_0536_),
    .B1(_0564_),
    .A1(_0542_),
    .Y(_0565_),
    .A2(_0546_));
 sg13g2_a21oi_2 _3468_ (.B1(_0565_),
    .Y(_0566_),
    .A2(_0563_),
    .A1(_0536_));
 sg13g2_a221oi_1 _3469_ (.B2(_0556_),
    .C1(_2239_),
    .B1(_0566_),
    .A1(_0559_),
    .Y(_0567_),
    .A2(_0562_));
 sg13g2_and2_1 _3470_ (.A(net51),
    .B(_0002_),
    .X(_0568_));
 sg13g2_a221oi_1 _3471_ (.B2(_0023_),
    .C1(_2238_),
    .B1(_0568_),
    .A1(_2249_),
    .Y(_0569_),
    .A2(_0020_));
 sg13g2_or3_1 _3472_ (.A(_0535_),
    .B(_0567_),
    .C(_0569_),
    .X(_0570_));
 sg13g2_o21ai_1 _3473_ (.B1(_0570_),
    .Y(\g.g_y[2].g_x[6].t.w_dh ),
    .A1(_2235_),
    .A2(_0534_));
 sg13g2_a221oi_1 _3474_ (.B2(_0556_),
    .C1(_2238_),
    .B1(_0566_),
    .A1(_0559_),
    .Y(_0571_),
    .A2(_0562_));
 sg13g2_a221oi_1 _3475_ (.B2(_0023_),
    .C1(_2239_),
    .B1(_0568_),
    .A1(_2249_),
    .Y(_0572_),
    .A2(_0020_));
 sg13g2_nor2_1 _3476_ (.A(_0184_),
    .B(_0520_),
    .Y(_0573_));
 sg13g2_nor3_1 _3477_ (.A(_0262_),
    .B(_0531_),
    .C(_0532_),
    .Y(_0574_));
 sg13g2_nor3_1 _3478_ (.A(_0266_),
    .B(_0286_),
    .C(_0526_),
    .Y(_0575_));
 sg13g2_nor3_1 _3479_ (.A(_0183_),
    .B(_0574_),
    .C(_0575_),
    .Y(_0576_));
 sg13g2_or4_1 _3480_ (.A(_0571_),
    .B(_0572_),
    .C(_0573_),
    .D(_0576_),
    .X(\g.g_y[2].g_x[6].t.w_na ));
 sg13g2_nor2_1 _3481_ (.A(_0535_),
    .B(net82),
    .Y(_0577_));
 sg13g2_nor2_1 _3482_ (.A(_2235_),
    .B(net61),
    .Y(_0578_));
 sg13g2_or2_1 _3483_ (.X(_0579_),
    .B(_0569_),
    .A(_0567_));
 sg13g2_nor2_1 _3484_ (.A(\g.g_y[2].g_x[5].t.out_sc ),
    .B(net64),
    .Y(_0580_));
 sg13g2_a221oi_1 _3485_ (.B2(_0579_),
    .C1(_0580_),
    .B1(_0578_),
    .A1(_0534_),
    .Y(\g.g_y[2].g_x[6].t.w_si ),
    .A2(_0577_));
 sg13g2_nor3_1 _3486_ (.A(_0266_),
    .B(_0531_),
    .C(_0532_),
    .Y(_0581_));
 sg13g2_a21o_1 _3487_ (.A2(_0527_),
    .A1(_0266_),
    .B1(_0581_),
    .X(\g.g_y[2].g_x[7].t.out_r ));
 sg13g2_a221oi_1 _3488_ (.B2(_0284_),
    .C1(_0277_),
    .B1(_0265_),
    .A1(_0266_),
    .Y(_0582_),
    .A2(_0263_));
 sg13g2_a221oi_1 _3489_ (.B2(_0525_),
    .C1(_0276_),
    .B1(_0523_),
    .A1(_0280_),
    .Y(_0583_),
    .A2(_0522_));
 sg13g2_nor3_1 _3490_ (.A(_1894_),
    .B(_0582_),
    .C(_0583_),
    .Y(_0584_));
 sg13g2_a21o_1 _3491_ (.A2(net59),
    .A1(\g.g_y[2].g_x[6].t.out_sc ),
    .B1(_0584_),
    .X(\g.g_y[2].g_x[7].t.w_si ));
 sg13g2_buf_1 _3492_ (.A(net82),
    .X(_0585_));
 sg13g2_or2_1 _3493_ (.X(_0586_),
    .B(_1833_),
    .A(_1836_));
 sg13g2_o21ai_1 _3494_ (.B1(_0586_),
    .Y(_0587_),
    .A1(_0057_),
    .A2(_1835_));
 sg13g2_buf_1 _3495_ (.A(_0587_),
    .X(_0588_));
 sg13g2_nor2_1 _3496_ (.A(_0329_),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_nor2_1 _3497_ (.A(_0330_),
    .B(_0328_),
    .Y(_0590_));
 sg13g2_nor2_1 _3498_ (.A(_0589_),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_nor2_1 _3499_ (.A(_0311_),
    .B(_0316_),
    .Y(_0592_));
 sg13g2_nor3_1 _3500_ (.A(_0335_),
    .B(_0592_),
    .C(_0318_),
    .Y(_0593_));
 sg13g2_a21o_1 _3501_ (.A2(_0591_),
    .A1(_0335_),
    .B1(_0593_),
    .X(_0594_));
 sg13g2_nand2_1 _3502_ (.Y(_0595_),
    .A(\g.g_y[2].g_x[7].t.out_sc ),
    .B(_2175_));
 sg13g2_o21ai_1 _3503_ (.B1(_0595_),
    .Y(\g.g_y[3].g_x[0].t.w_si ),
    .A1(net42),
    .A2(_0594_));
 sg13g2_inv_1 _3504_ (.Y(_0596_),
    .A(_0088_));
 sg13g2_mux2_1 _3505_ (.A0(_1923_),
    .A1(_1919_),
    .S(_1920_),
    .X(_0597_));
 sg13g2_buf_1 _3506_ (.A(_0597_),
    .X(_0598_));
 sg13g2_and2_1 _3507_ (.A(_0420_),
    .B(_0412_),
    .X(_0599_));
 sg13g2_a22oi_1 _3508_ (.Y(_0600_),
    .B1(_0599_),
    .B2(_0410_),
    .A2(_0598_),
    .A1(_0415_));
 sg13g2_nor2b_1 _3509_ (.A(_0402_),
    .B_N(net26),
    .Y(_0601_));
 sg13g2_o21ai_1 _3510_ (.B1(_0601_),
    .Y(_0602_),
    .A1(_0404_),
    .A2(_0600_));
 sg13g2_nor2_1 _3511_ (.A(_0402_),
    .B(_0393_),
    .Y(_0603_));
 sg13g2_mux2_1 _3512_ (.A0(_0411_),
    .A1(_0407_),
    .S(_0409_),
    .X(_0604_));
 sg13g2_mux2_1 _3513_ (.A0(_0604_),
    .A1(_0598_),
    .S(_0420_),
    .X(_0605_));
 sg13g2_and2_1 _3514_ (.A(_0402_),
    .B(net26),
    .X(_0606_));
 sg13g2_nor2b_1 _3515_ (.A(_0393_),
    .B_N(_0402_),
    .Y(_0607_));
 sg13g2_nor2b_1 _3516_ (.A(_0398_),
    .B_N(_0607_),
    .Y(_0608_));
 sg13g2_a221oi_1 _3517_ (.B2(_0606_),
    .C1(_0608_),
    .B1(_0605_),
    .A1(\g.g_y[3].g_x[2].t.out_sc ),
    .Y(_0609_),
    .A2(_0603_));
 sg13g2_nand3_1 _3518_ (.B(_0602_),
    .C(_0609_),
    .A(_0312_),
    .Y(_0610_));
 sg13g2_mux2_1 _3519_ (.A0(_0328_),
    .A1(_0588_),
    .S(_0329_),
    .X(_0611_));
 sg13g2_nand2_1 _3520_ (.Y(_0612_),
    .A(net4),
    .B(_0317_));
 sg13g2_nor2_1 _3521_ (.A(_0317_),
    .B(\g.g_y[3].g_x[0].t.out_sc ),
    .Y(_0613_));
 sg13g2_nor2_1 _3522_ (.A(_0311_),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_o21ai_1 _3523_ (.B1(_0614_),
    .Y(_0615_),
    .A1(_0611_),
    .A2(_0612_));
 sg13g2_o21ai_1 _3524_ (.B1(_0317_),
    .Y(_0616_),
    .A1(_0330_),
    .A2(_0328_));
 sg13g2_a21oi_1 _3525_ (.A1(_0333_),
    .A2(_0335_),
    .Y(_0617_),
    .B1(\g.g_y[3].g_x[0].t.r_h ));
 sg13g2_o21ai_1 _3526_ (.B1(_0617_),
    .Y(_0618_),
    .A1(_0589_),
    .A2(_0616_));
 sg13g2_nand3_1 _3527_ (.B(_0615_),
    .C(_0618_),
    .A(_0399_),
    .Y(_0619_));
 sg13g2_and3_1 _3528_ (.X(_0620_),
    .A(_0596_),
    .B(_0610_),
    .C(_0619_));
 sg13g2_buf_1 _3529_ (.A(\g.g_y[4].g_x[1].t.r_d ),
    .X(_0621_));
 sg13g2_inv_2 _3530_ (.Y(_0622_),
    .A(_0621_));
 sg13g2_mux2_1 _3531_ (.A0(\g.g_y[4].g_x[0].t.out_sc ),
    .A1(\g.g_y[4].g_x[0].t.r_gnl ),
    .S(_0322_),
    .X(_0623_));
 sg13g2_buf_2 _3532_ (.A(\g.g_y[4].g_x[0].t.r_h ),
    .X(_0624_));
 sg13g2_mux2_1 _3533_ (.A0(_0325_),
    .A1(_0623_),
    .S(_0624_),
    .X(_0625_));
 sg13g2_buf_2 _3534_ (.A(_0625_),
    .X(_0626_));
 sg13g2_mux2_1 _3535_ (.A0(\g.g_y[4].g_x[2].t.out_sc ),
    .A1(\g.g_y[4].g_x[2].t.r_gnl ),
    .S(_0405_),
    .X(_0627_));
 sg13g2_buf_2 _3536_ (.A(\g.g_y[4].g_x[2].t.r_h ),
    .X(_0628_));
 sg13g2_inv_1 _3537_ (.Y(_0629_),
    .A(_0628_));
 sg13g2_mux2_1 _3538_ (.A0(_0411_),
    .A1(_0627_),
    .S(_0629_),
    .X(_0630_));
 sg13g2_buf_1 _3539_ (.A(\g.g_y[4].g_x[1].t.r_h ),
    .X(_0631_));
 sg13g2_inv_1 _3540_ (.Y(_0632_),
    .A(_0631_));
 sg13g2_mux2_1 _3541_ (.A0(_0626_),
    .A1(_0630_),
    .S(_0632_),
    .X(_0633_));
 sg13g2_mux2_1 _3542_ (.A0(\g.g_y[3].g_x[1].t.r_ghl ),
    .A1(_0089_),
    .S(_0087_),
    .X(_0634_));
 sg13g2_buf_1 _3543_ (.A(_0634_),
    .X(_0635_));
 sg13g2_buf_1 _3544_ (.A(\g.g_y[5].g_x[1].t.r_ghl ),
    .X(_0636_));
 sg13g2_buf_1 _3545_ (.A(\g.g_y[5].g_x[1].t.r_d ),
    .X(_0637_));
 sg13g2_mux2_1 _3546_ (.A0(\g.g_y[5].g_x[1].t.r_gnl ),
    .A1(\g.g_y[5].g_x[1].t.out_sc ),
    .S(_0637_),
    .X(_0638_));
 sg13g2_buf_1 _3547_ (.A(_0638_),
    .X(_0639_));
 sg13g2_buf_2 _3548_ (.A(\g.g_y[5].g_x[1].t.r_v ),
    .X(_0640_));
 sg13g2_inv_2 _3549_ (.Y(_0641_),
    .A(_0640_));
 sg13g2_mux2_1 _3550_ (.A0(_0636_),
    .A1(_0639_),
    .S(_0641_),
    .X(_0642_));
 sg13g2_buf_2 _3551_ (.A(\g.g_y[4].g_x[1].t.r_v ),
    .X(_0643_));
 sg13g2_inv_1 _3552_ (.Y(_0644_),
    .A(_0643_));
 sg13g2_mux2_1 _3553_ (.A0(_0635_),
    .A1(_0642_),
    .S(_0644_),
    .X(_0645_));
 sg13g2_nand3_1 _3554_ (.B(_0633_),
    .C(_0645_),
    .A(_0622_),
    .Y(_0646_));
 sg13g2_nor2_1 _3555_ (.A(_0622_),
    .B(\g.g_y[4].g_x[1].t.out_sc ),
    .Y(_0647_));
 sg13g2_nor2_1 _3556_ (.A(_0643_),
    .B(_0647_),
    .Y(_0648_));
 sg13g2_nand2b_1 _3557_ (.Y(_0649_),
    .B(_0641_),
    .A_N(_0639_));
 sg13g2_inv_1 _3558_ (.Y(_0650_),
    .A(_0636_));
 sg13g2_a21oi_1 _3559_ (.A1(_0650_),
    .A2(_0640_),
    .Y(_0651_),
    .B1(_0644_));
 sg13g2_a221oi_1 _3560_ (.B2(_0651_),
    .C1(_0622_),
    .B1(_0649_),
    .A1(_0644_),
    .Y(_0652_),
    .A2(_0635_));
 sg13g2_buf_1 _3561_ (.A(_0652_),
    .X(_0653_));
 sg13g2_nand2b_1 _3562_ (.Y(_0654_),
    .B(_0629_),
    .A_N(_0627_));
 sg13g2_inv_1 _3563_ (.Y(_0655_),
    .A(_0411_));
 sg13g2_a21oi_1 _3564_ (.A1(_0655_),
    .A2(_0628_),
    .Y(_0656_),
    .B1(_0632_));
 sg13g2_a221oi_1 _3565_ (.B2(_0656_),
    .C1(_0621_),
    .B1(_0654_),
    .A1(_0632_),
    .Y(_0657_),
    .A2(_0626_));
 sg13g2_nor2_1 _3566_ (.A(_0653_),
    .B(_0657_),
    .Y(_0658_));
 sg13g2_inv_1 _3567_ (.Y(_0659_),
    .A(_0087_));
 sg13g2_a221oi_1 _3568_ (.B2(_0643_),
    .C1(_0659_),
    .B1(_0658_),
    .A1(_0646_),
    .Y(_0660_),
    .A2(_0648_));
 sg13g2_nor2_1 _3569_ (.A(net27),
    .B(_0349_),
    .Y(_0661_));
 sg13g2_nand2_1 _3570_ (.Y(_0662_),
    .A(_0084_),
    .B(_0661_));
 sg13g2_a21oi_1 _3571_ (.A1(_0086_),
    .A2(_0094_),
    .Y(_0663_),
    .B1(_0355_));
 sg13g2_a21oi_1 _3572_ (.A1(_0086_),
    .A2(_0349_),
    .Y(_0664_),
    .B1(_0095_));
 sg13g2_nand2b_1 _3573_ (.Y(_0665_),
    .B(_0370_),
    .A_N(net27));
 sg13g2_a221oi_1 _3574_ (.B2(_0665_),
    .C1(_0087_),
    .B1(_0664_),
    .A1(_0662_),
    .Y(_0666_),
    .A2(_0663_));
 sg13g2_nor3_1 _3575_ (.A(_0596_),
    .B(_0660_),
    .C(_0666_),
    .Y(_0667_));
 sg13g2_or2_1 _3576_ (.X(\g.g_y[3].g_x[1].t.w_dh ),
    .B(_0667_),
    .A(_0620_));
 sg13g2_a21oi_1 _3577_ (.A1(_0615_),
    .A2(_0618_),
    .Y(_0668_),
    .B1(_0399_));
 sg13g2_a21oi_1 _3578_ (.A1(_0602_),
    .A2(_0609_),
    .Y(_0669_),
    .B1(_0312_));
 sg13g2_a22oi_1 _3579_ (.Y(_0670_),
    .B1(_0658_),
    .B2(_0643_),
    .A2(_0648_),
    .A1(_0646_));
 sg13g2_a221oi_1 _3580_ (.B2(_0665_),
    .C1(_0659_),
    .B1(_0664_),
    .A1(_0662_),
    .Y(_0671_),
    .A2(_0663_));
 sg13g2_a21oi_1 _3581_ (.A1(_0659_),
    .A2(_0670_),
    .Y(_0672_),
    .B1(_0671_));
 sg13g2_o21ai_1 _3582_ (.B1(_0672_),
    .Y(\g.g_y[3].g_x[1].t.w_na ),
    .A1(_0668_),
    .A2(_0669_));
 sg13g2_nand2_1 _3583_ (.Y(_0673_),
    .A(\g.g_y[3].g_x[0].t.out_sc ),
    .B(_0109_));
 sg13g2_nand4_1 _3584_ (.B(net45),
    .C(_0610_),
    .A(_0088_),
    .Y(_0674_),
    .D(_0619_));
 sg13g2_or4_1 _3585_ (.A(_0088_),
    .B(net74),
    .C(_0660_),
    .D(_0666_),
    .X(_0675_));
 sg13g2_nand3_1 _3586_ (.B(_0674_),
    .C(_0675_),
    .A(_0673_),
    .Y(\g.g_y[3].g_x[1].t.w_si ));
 sg13g2_nand2_1 _3587_ (.Y(_0676_),
    .A(net26),
    .B(_0418_));
 sg13g2_o21ai_1 _3588_ (.B1(_0676_),
    .Y(_0677_),
    .A1(net26),
    .A2(_0605_));
 sg13g2_nand2_1 _3589_ (.Y(_0678_),
    .A(\g.g_y[3].g_x[1].t.out_sc ),
    .B(net52));
 sg13g2_o21ai_1 _3590_ (.B1(_0678_),
    .Y(\g.g_y[3].g_x[2].t.w_si ),
    .A1(net42),
    .A2(_0677_));
 sg13g2_inv_1 _3591_ (.Y(_0679_),
    .A(_0150_));
 sg13g2_or4_1 _3592_ (.A(_0162_),
    .B(_0139_),
    .C(_0148_),
    .D(_0376_),
    .X(_0680_));
 sg13g2_nor2_1 _3593_ (.A(_0156_),
    .B(_0139_),
    .Y(_0681_));
 sg13g2_nor3_1 _3594_ (.A(_0156_),
    .B(_0157_),
    .C(_0382_),
    .Y(_0682_));
 sg13g2_a221oi_1 _3595_ (.B2(_0681_),
    .C1(_0682_),
    .B1(_0160_),
    .A1(_0156_),
    .Y(_0683_),
    .A2(_0158_));
 sg13g2_a21oi_1 _3596_ (.A1(_0680_),
    .A2(_0683_),
    .Y(_0684_),
    .B1(_0149_));
 sg13g2_buf_2 _3597_ (.A(\g.g_y[4].g_x[3].t.r_d ),
    .X(_0685_));
 sg13g2_mux2_1 _3598_ (.A0(\g.g_y[4].g_x[4].t.out_sc ),
    .A1(\g.g_y[4].g_x[4].t.r_gnl ),
    .S(_0477_),
    .X(_0686_));
 sg13g2_buf_1 _3599_ (.A(_0686_),
    .X(_0687_));
 sg13g2_buf_2 _3600_ (.A(\g.g_y[4].g_x[4].t.r_h ),
    .X(_0688_));
 sg13g2_inv_1 _3601_ (.Y(_0689_),
    .A(_0688_));
 sg13g2_nand2b_1 _3602_ (.Y(_0690_),
    .B(_0689_),
    .A_N(_0687_));
 sg13g2_inv_1 _3603_ (.Y(_0691_),
    .A(_0479_));
 sg13g2_buf_1 _3604_ (.A(\g.g_y[4].g_x[3].t.r_h ),
    .X(_0692_));
 sg13g2_a21oi_1 _3605_ (.A1(_0691_),
    .A2(_0688_),
    .Y(_0693_),
    .B1(_0692_));
 sg13g2_mux2_1 _3606_ (.A0(_0411_),
    .A1(_0627_),
    .S(_0628_),
    .X(_0694_));
 sg13g2_buf_1 _3607_ (.A(_0694_),
    .X(_0695_));
 sg13g2_a22oi_1 _3608_ (.Y(_0696_),
    .B1(_0695_),
    .B2(_0692_),
    .A2(_0693_),
    .A1(_0690_));
 sg13g2_buf_2 _3609_ (.A(\g.g_y[5].g_x[3].t.r_d ),
    .X(_0697_));
 sg13g2_mux2_1 _3610_ (.A0(\g.g_y[5].g_x[3].t.r_gnl ),
    .A1(\g.g_y[5].g_x[3].t.out_sc ),
    .S(_0697_),
    .X(_0698_));
 sg13g2_buf_2 _3611_ (.A(\g.g_y[5].g_x[3].t.r_v ),
    .X(_0699_));
 sg13g2_inv_1 _3612_ (.Y(_0700_),
    .A(_0699_));
 sg13g2_nand2b_1 _3613_ (.Y(_0701_),
    .B(_0700_),
    .A_N(_0698_));
 sg13g2_buf_1 _3614_ (.A(\g.g_y[5].g_x[3].t.r_ghl ),
    .X(_0702_));
 sg13g2_inv_1 _3615_ (.Y(_0703_),
    .A(_0702_));
 sg13g2_buf_2 _3616_ (.A(\g.g_y[4].g_x[3].t.r_v ),
    .X(_0704_));
 sg13g2_a21oi_1 _3617_ (.A1(_0703_),
    .A2(_0699_),
    .Y(_0705_),
    .B1(_0704_));
 sg13g2_mux2_1 _3618_ (.A0(_0152_),
    .A1(_0151_),
    .S(_0149_),
    .X(_0706_));
 sg13g2_a22oi_1 _3619_ (.Y(_0707_),
    .B1(_0706_),
    .B2(_0704_),
    .A2(_0705_),
    .A1(_0701_));
 sg13g2_or3_1 _3620_ (.A(_0685_),
    .B(_0696_),
    .C(_0707_),
    .X(_0708_));
 sg13g2_buf_1 _3621_ (.A(_0708_),
    .X(_0709_));
 sg13g2_inv_1 _3622_ (.Y(_0710_),
    .A(_0704_));
 sg13g2_nand2b_1 _3623_ (.Y(_0711_),
    .B(_0685_),
    .A_N(\g.g_y[4].g_x[3].t.out_sc ));
 sg13g2_and2_1 _3624_ (.A(_0710_),
    .B(_0711_),
    .X(_0712_));
 sg13g2_a21oi_1 _3625_ (.A1(_0703_),
    .A2(_0699_),
    .Y(_0713_),
    .B1(_0710_));
 sg13g2_inv_1 _3626_ (.Y(_0714_),
    .A(_0685_));
 sg13g2_a221oi_1 _3627_ (.B2(_0701_),
    .C1(_0714_),
    .B1(_0713_),
    .A1(_0710_),
    .Y(_0715_),
    .A2(_0706_));
 sg13g2_inv_1 _3628_ (.Y(_0716_),
    .A(_0692_));
 sg13g2_a21oi_1 _3629_ (.A1(_0691_),
    .A2(_0688_),
    .Y(_0717_),
    .B1(_0716_));
 sg13g2_a221oi_1 _3630_ (.B2(_0690_),
    .C1(_0685_),
    .B1(_0717_),
    .A1(_0716_),
    .Y(_0718_),
    .A2(_0695_));
 sg13g2_nor2_1 _3631_ (.A(_0715_),
    .B(_0718_),
    .Y(_0719_));
 sg13g2_a221oi_1 _3632_ (.B2(_0704_),
    .C1(_0380_),
    .B1(_0719_),
    .A1(_0709_),
    .Y(_0720_),
    .A2(_0712_));
 sg13g2_or2_1 _3633_ (.X(_0721_),
    .B(_0720_),
    .A(_0684_));
 sg13g2_nor2_1 _3634_ (.A(_0466_),
    .B(_0457_),
    .Y(_0722_));
 sg13g2_o21ai_1 _3635_ (.B1(_0722_),
    .Y(_0723_),
    .A1(_0488_),
    .A2(_0494_));
 sg13g2_mux2_1 _3636_ (.A0(_0481_),
    .A1(_0490_),
    .S(_0455_),
    .X(_0724_));
 sg13g2_nor2_1 _3637_ (.A(_0485_),
    .B(_0457_),
    .Y(_0725_));
 sg13g2_nand2_1 _3638_ (.Y(_0726_),
    .A(_0724_),
    .B(_0725_));
 sg13g2_nor2_1 _3639_ (.A(_0485_),
    .B(_0456_),
    .Y(_0727_));
 sg13g2_nor2_1 _3640_ (.A(_0466_),
    .B(_0456_),
    .Y(_0728_));
 sg13g2_a22oi_1 _3641_ (.Y(_0729_),
    .B1(_0728_),
    .B2(_0458_),
    .A2(_0727_),
    .A1(_0471_));
 sg13g2_nand4_1 _3642_ (.B(_0723_),
    .C(_0726_),
    .A(_0395_),
    .Y(_0730_),
    .D(_0729_));
 sg13g2_o21ai_1 _3643_ (.B1(_0606_),
    .Y(_0731_),
    .A1(_0404_),
    .A2(_0600_));
 sg13g2_nand2_1 _3644_ (.Y(_0732_),
    .A(_0601_),
    .B(_0605_));
 sg13g2_nor2b_1 _3645_ (.A(_0401_),
    .B_N(_0603_),
    .Y(_0733_));
 sg13g2_a21oi_1 _3646_ (.A1(\g.g_y[3].g_x[2].t.out_sc ),
    .A2(_0607_),
    .Y(_0734_),
    .B1(_0733_));
 sg13g2_nand4_1 _3647_ (.B(_0731_),
    .C(_0732_),
    .A(_0472_),
    .Y(_0735_),
    .D(_0734_));
 sg13g2_nand3_1 _3648_ (.B(_0730_),
    .C(_0735_),
    .A(_0679_),
    .Y(_0736_));
 sg13g2_o21ai_1 _3649_ (.B1(_0736_),
    .Y(\g.g_y[3].g_x[3].t.w_dh ),
    .A1(_0679_),
    .A2(_0721_));
 sg13g2_nand3_1 _3650_ (.B(_0726_),
    .C(_0729_),
    .A(_0723_),
    .Y(_0737_));
 sg13g2_nand3_1 _3651_ (.B(_0732_),
    .C(_0734_),
    .A(_0731_),
    .Y(_0738_));
 sg13g2_mux2_1 _3652_ (.A0(_0737_),
    .A1(_0738_),
    .S(_0395_),
    .X(_0739_));
 sg13g2_a22oi_1 _3653_ (.Y(_0740_),
    .B1(_0719_),
    .B2(_0704_),
    .A2(_0712_),
    .A1(_0709_));
 sg13g2_nand2_1 _3654_ (.Y(_0741_),
    .A(_0380_),
    .B(_0740_));
 sg13g2_a21o_1 _3655_ (.A2(_0683_),
    .A1(_0680_),
    .B1(_0380_),
    .X(_0742_));
 sg13g2_nand3_1 _3656_ (.B(_0741_),
    .C(_0742_),
    .A(_0739_),
    .Y(\g.g_y[3].g_x[3].t.w_na ));
 sg13g2_nand2_1 _3657_ (.Y(_0743_),
    .A(\g.g_y[3].g_x[2].t.out_sc ),
    .B(net47));
 sg13g2_nand4_1 _3658_ (.B(net45),
    .C(_0730_),
    .A(_0150_),
    .Y(_0744_),
    .D(_0735_));
 sg13g2_or4_1 _3659_ (.A(_0150_),
    .B(net74),
    .C(_0684_),
    .D(_0720_),
    .X(_0745_));
 sg13g2_nand3_1 _3660_ (.B(_0744_),
    .C(_0745_),
    .A(_0743_),
    .Y(\g.g_y[3].g_x[3].t.w_si ));
 sg13g2_nor2_1 _3661_ (.A(_0472_),
    .B(_0396_),
    .Y(_0746_));
 sg13g2_nor2_1 _3662_ (.A(_0746_),
    .B(_0474_),
    .Y(_0747_));
 sg13g2_mux2_1 _3663_ (.A0(_0471_),
    .A1(_0747_),
    .S(_0485_),
    .X(_0748_));
 sg13g2_nand2b_1 _3664_ (.Y(_0749_),
    .B(_0457_),
    .A_N(_0724_));
 sg13g2_o21ai_1 _3665_ (.B1(_0749_),
    .Y(_0750_),
    .A1(_0457_),
    .A2(_0748_));
 sg13g2_buf_1 _3666_ (.A(net77),
    .X(_0751_));
 sg13g2_nand2_1 _3667_ (.Y(_0752_),
    .A(\g.g_y[3].g_x[3].t.out_sc ),
    .B(net41));
 sg13g2_o21ai_1 _3668_ (.B1(_0752_),
    .Y(\g.g_y[3].g_x[4].t.w_si ),
    .A1(net42),
    .A2(_0750_));
 sg13g2_buf_1 _3669_ (.A(\g.g_y[4].g_x[5].t.r_v ),
    .X(_0753_));
 sg13g2_inv_2 _3670_ (.Y(_0754_),
    .A(_0753_));
 sg13g2_mux2_1 _3671_ (.A0(_0198_),
    .A1(_0195_),
    .S(_0193_),
    .X(_0755_));
 sg13g2_buf_8 _3672_ (.A(\g.g_y[5].g_x[5].t.r_d ),
    .X(_0756_));
 sg13g2_mux2_1 _3673_ (.A0(\g.g_y[5].g_x[5].t.r_gnl ),
    .A1(\g.g_y[5].g_x[5].t.out_sc ),
    .S(_0756_),
    .X(_0757_));
 sg13g2_buf_1 _3674_ (.A(_0757_),
    .X(_0758_));
 sg13g2_buf_2 _3675_ (.A(\g.g_y[5].g_x[5].t.r_v ),
    .X(_0759_));
 sg13g2_inv_2 _3676_ (.Y(_0760_),
    .A(_0759_));
 sg13g2_nand2b_1 _3677_ (.Y(_0761_),
    .B(_0760_),
    .A_N(_0758_));
 sg13g2_buf_2 _3678_ (.A(\g.g_y[5].g_x[5].t.r_ghl ),
    .X(_0762_));
 sg13g2_inv_1 _3679_ (.Y(_0763_),
    .A(_0762_));
 sg13g2_a21oi_1 _3680_ (.A1(_0763_),
    .A2(_0759_),
    .Y(_0764_),
    .B1(_0754_));
 sg13g2_buf_2 _3681_ (.A(\g.g_y[4].g_x[5].t.r_d ),
    .X(_0765_));
 sg13g2_inv_1 _3682_ (.Y(_0766_),
    .A(_0765_));
 sg13g2_a221oi_1 _3683_ (.B2(_0764_),
    .C1(_0766_),
    .B1(_0761_),
    .A1(_0754_),
    .Y(_0767_),
    .A2(_0755_));
 sg13g2_buf_2 _3684_ (.A(_0767_),
    .X(_0768_));
 sg13g2_or2_1 _3685_ (.X(_0769_),
    .B(_0687_),
    .A(_0689_));
 sg13g2_buf_1 _3686_ (.A(\g.g_y[4].g_x[5].t.r_h ),
    .X(_0770_));
 sg13g2_a21oi_1 _3687_ (.A1(_0691_),
    .A2(_0689_),
    .Y(_0771_),
    .B1(_0770_));
 sg13g2_mux2_1 _3688_ (.A0(\g.g_y[4].g_x[6].t.out_sc ),
    .A1(\g.g_y[4].g_x[6].t.r_gnl ),
    .S(_0549_),
    .X(_0772_));
 sg13g2_buf_2 _3689_ (.A(\g.g_y[4].g_x[6].t.r_h ),
    .X(_0773_));
 sg13g2_inv_1 _3690_ (.Y(_0774_),
    .A(_0773_));
 sg13g2_mux2_1 _3691_ (.A0(_0551_),
    .A1(_0772_),
    .S(_0774_),
    .X(_0775_));
 sg13g2_buf_1 _3692_ (.A(_0775_),
    .X(_0776_));
 sg13g2_a221oi_1 _3693_ (.B2(_0770_),
    .C1(_0765_),
    .B1(_0776_),
    .A1(_0769_),
    .Y(_0777_),
    .A2(_0771_));
 sg13g2_o21ai_1 _3694_ (.B1(_0753_),
    .Y(_0778_),
    .A1(_0768_),
    .A2(_0777_));
 sg13g2_nand2b_1 _3695_ (.Y(_0779_),
    .B(_0765_),
    .A_N(\g.g_y[4].g_x[5].t.out_sc ));
 sg13g2_nand2b_1 _3696_ (.Y(_0780_),
    .B(_0754_),
    .A_N(_0779_));
 sg13g2_mux2_1 _3697_ (.A0(_0762_),
    .A1(_0758_),
    .S(_0760_),
    .X(_0781_));
 sg13g2_mux2_1 _3698_ (.A0(_0479_),
    .A1(_0687_),
    .S(_0688_),
    .X(_0782_));
 sg13g2_inv_1 _3699_ (.Y(_0783_),
    .A(_0770_));
 sg13g2_mux2_1 _3700_ (.A0(_0782_),
    .A1(_0776_),
    .S(_0783_),
    .X(_0784_));
 sg13g2_nand4_1 _3701_ (.B(_0766_),
    .C(_0781_),
    .A(_0754_),
    .Y(_0785_),
    .D(_0784_));
 sg13g2_nand4_1 _3702_ (.B(_0778_),
    .C(_0780_),
    .A(net46),
    .Y(_0786_),
    .D(_0785_));
 sg13g2_or2_1 _3703_ (.X(_0787_),
    .B(_0178_),
    .A(net46));
 sg13g2_or4_1 _3704_ (.A(_0197_),
    .B(_0190_),
    .C(_0202_),
    .D(_0787_),
    .X(_0788_));
 sg13g2_o21ai_1 _3705_ (.B1(_0197_),
    .Y(_0789_),
    .A1(_0209_),
    .A2(_0211_));
 sg13g2_a21oi_1 _3706_ (.A1(_0191_),
    .A2(_0206_),
    .Y(_0790_),
    .B1(net46));
 sg13g2_nand3_1 _3707_ (.B(_0789_),
    .C(_0790_),
    .A(_0788_),
    .Y(_0791_));
 sg13g2_inv_1 _3708_ (.Y(_0792_),
    .A(_0194_));
 sg13g2_a21oi_1 _3709_ (.A1(_0786_),
    .A2(_0791_),
    .Y(_0793_),
    .B1(_0792_));
 sg13g2_inv_1 _3710_ (.Y(_0794_),
    .A(_0536_));
 sg13g2_nor2_1 _3711_ (.A(_0541_),
    .B(_0794_),
    .Y(_0795_));
 sg13g2_o21ai_1 _3712_ (.B1(_0795_),
    .Y(_0796_),
    .A1(_0547_),
    .A2(_0557_));
 sg13g2_inv_1 _3713_ (.Y(_0797_),
    .A(_0548_));
 sg13g2_mux2_1 _3714_ (.A0(_0551_),
    .A1(_0550_),
    .S(_0797_),
    .X(_0798_));
 sg13g2_mux2_1 _3715_ (.A0(_2241_),
    .A1(_2237_),
    .S(_2238_),
    .X(_0799_));
 sg13g2_mux2_1 _3716_ (.A0(_0798_),
    .A1(_0799_),
    .S(_0560_),
    .X(_0800_));
 sg13g2_nor2_1 _3717_ (.A(_0542_),
    .B(_0794_),
    .Y(_0801_));
 sg13g2_nor2_1 _3718_ (.A(_0541_),
    .B(_0536_),
    .Y(_0802_));
 sg13g2_nor2_1 _3719_ (.A(_0542_),
    .B(_0536_),
    .Y(_0803_));
 sg13g2_and3_1 _3720_ (.X(_0804_),
    .A(_0540_),
    .B(_0543_),
    .C(_0803_));
 sg13g2_a221oi_1 _3721_ (.B2(\g.g_y[3].g_x[6].t.out_sc ),
    .C1(_0804_),
    .B1(_0802_),
    .A1(_0800_),
    .Y(_0805_),
    .A2(_0801_));
 sg13g2_nand3_1 _3722_ (.B(_0796_),
    .C(_0805_),
    .A(_0468_),
    .Y(_0806_));
 sg13g2_o21ai_1 _3723_ (.B1(_0725_),
    .Y(_0807_),
    .A1(_0488_),
    .A2(_0494_));
 sg13g2_nand2_1 _3724_ (.Y(_0808_),
    .A(_0724_),
    .B(_0722_));
 sg13g2_a22oi_1 _3725_ (.Y(_0809_),
    .B1(_0728_),
    .B2(_0747_),
    .A2(_0727_),
    .A1(_0458_));
 sg13g2_nand4_1 _3726_ (.B(_0807_),
    .C(_0808_),
    .A(_0469_),
    .Y(_0810_),
    .D(_0809_));
 sg13g2_nand3_1 _3727_ (.B(_0806_),
    .C(_0810_),
    .A(_0792_),
    .Y(_0811_));
 sg13g2_nand2b_1 _3728_ (.Y(\g.g_y[3].g_x[5].t.w_dh ),
    .B(_0811_),
    .A_N(_0793_));
 sg13g2_nand3_1 _3729_ (.B(_0808_),
    .C(_0809_),
    .A(_0807_),
    .Y(_0812_));
 sg13g2_a21oi_1 _3730_ (.A1(_0796_),
    .A2(_0805_),
    .Y(_0813_),
    .B1(_0468_));
 sg13g2_a21oi_1 _3731_ (.A1(_0468_),
    .A2(_0812_),
    .Y(_0814_),
    .B1(_0813_));
 sg13g2_mux2_1 _3732_ (.A0(_0755_),
    .A1(_0781_),
    .S(_0754_),
    .X(_0815_));
 sg13g2_nand3_1 _3733_ (.B(_0784_),
    .C(_0815_),
    .A(_0766_),
    .Y(_0816_));
 sg13g2_a21o_1 _3734_ (.A2(_0816_),
    .A1(_0779_),
    .B1(_0753_),
    .X(_0817_));
 sg13g2_a21o_1 _3735_ (.A2(_0817_),
    .A1(_0778_),
    .B1(net46),
    .X(_0818_));
 sg13g2_inv_1 _3736_ (.Y(_0819_),
    .A(_0789_));
 sg13g2_inv_1 _3737_ (.Y(_0820_),
    .A(_0206_));
 sg13g2_a21oi_1 _3738_ (.A1(_0204_),
    .A2(_0820_),
    .Y(_0821_),
    .B1(_0197_));
 sg13g2_o21ai_1 _3739_ (.B1(net46),
    .Y(_0822_),
    .A1(_0819_),
    .A2(_0821_));
 sg13g2_nand3b_1 _3740_ (.B(_0818_),
    .C(_0822_),
    .Y(\g.g_y[3].g_x[5].t.w_na ),
    .A_N(_0814_));
 sg13g2_and2_1 _3741_ (.A(_0458_),
    .B(net78),
    .X(_0823_));
 sg13g2_nand2_1 _3742_ (.Y(_0824_),
    .A(_0792_),
    .B(net81));
 sg13g2_a21oi_1 _3743_ (.A1(_0786_),
    .A2(_0791_),
    .Y(_0825_),
    .B1(_0824_));
 sg13g2_and4_1 _3744_ (.A(_0194_),
    .B(net73),
    .C(_0806_),
    .D(_0810_),
    .X(_0826_));
 sg13g2_or3_1 _3745_ (.A(_0823_),
    .B(_0825_),
    .C(_0826_),
    .X(\g.g_y[3].g_x[5].t.w_si ));
 sg13g2_a221oi_1 _3746_ (.B2(_0540_),
    .C1(_0794_),
    .B1(_0564_),
    .A1(_0542_),
    .Y(_0827_),
    .A2(_0546_));
 sg13g2_a21o_1 _3747_ (.A2(_0563_),
    .A1(_0794_),
    .B1(_0827_),
    .X(_0828_));
 sg13g2_nand2_1 _3748_ (.Y(_0829_),
    .A(\g.g_y[3].g_x[5].t.out_sc ),
    .B(net41));
 sg13g2_o21ai_1 _3749_ (.B1(_0829_),
    .Y(\g.g_y[3].g_x[6].t.w_si ),
    .A1(net42),
    .A2(_0828_));
 sg13g2_inv_1 _3750_ (.Y(_0830_),
    .A(\g.g_y[3].g_x[7].t.r_ghl ));
 sg13g2_nand2_1 _3751_ (.Y(_0831_),
    .A(_0537_),
    .B(_0538_));
 sg13g2_o21ai_1 _3752_ (.B1(_0831_),
    .Y(\g.g_y[3].g_x[7].t.out_r ),
    .A1(_0830_),
    .A2(_0537_));
 sg13g2_inv_1 _3753_ (.Y(_0832_),
    .A(_0271_));
 sg13g2_inv_1 _3754_ (.Y(_0833_),
    .A(\g.g_y[4].g_x[7].t.r_d ));
 sg13g2_mux2_1 _3755_ (.A0(_0623_),
    .A1(_0325_),
    .S(_0624_),
    .X(_0834_));
 sg13g2_buf_1 _3756_ (.A(_0834_),
    .X(_0835_));
 sg13g2_mux2_1 _3757_ (.A0(_0551_),
    .A1(_0772_),
    .S(_0773_),
    .X(_0836_));
 sg13g2_buf_1 _3758_ (.A(\g.g_y[4].g_x[7].t.r_h ),
    .X(_0837_));
 sg13g2_mux2_1 _3759_ (.A0(_0835_),
    .A1(_0836_),
    .S(net70),
    .X(_0838_));
 sg13g2_buf_1 _3760_ (.A(_0838_),
    .X(_0839_));
 sg13g2_mux2_1 _3761_ (.A0(\g.g_y[3].g_x[7].t.r_ghl ),
    .A1(_0273_),
    .S(_0270_),
    .X(_0840_));
 sg13g2_buf_8 _3762_ (.A(\g.g_y[5].g_x[7].t.r_d ),
    .X(_0841_));
 sg13g2_mux2_1 _3763_ (.A0(\g.g_y[5].g_x[7].t.r_gnl ),
    .A1(\g.g_y[5].g_x[7].t.out_sc ),
    .S(_0841_),
    .X(_0842_));
 sg13g2_buf_2 _3764_ (.A(\g.g_y[5].g_x[7].t.r_v ),
    .X(_0843_));
 sg13g2_mux2_1 _3765_ (.A0(_0842_),
    .A1(\g.g_y[5].g_x[7].t.r_ghl ),
    .S(_0843_),
    .X(_0844_));
 sg13g2_buf_2 _3766_ (.A(\g.g_y[4].g_x[7].t.r_v ),
    .X(_0845_));
 sg13g2_inv_1 _3767_ (.Y(_0846_),
    .A(_0845_));
 sg13g2_mux2_1 _3768_ (.A0(_0840_),
    .A1(_0844_),
    .S(_0846_),
    .X(_0847_));
 sg13g2_buf_1 _3769_ (.A(_0847_),
    .X(_0848_));
 sg13g2_nand3_1 _3770_ (.B(_0839_),
    .C(_0848_),
    .A(_0833_),
    .Y(_0849_));
 sg13g2_nor2_1 _3771_ (.A(_0833_),
    .B(\g.g_y[4].g_x[7].t.out_sc ),
    .Y(_0850_));
 sg13g2_nor2_1 _3772_ (.A(_0845_),
    .B(_0850_),
    .Y(_0851_));
 sg13g2_buf_1 _3773_ (.A(\g.g_y[4].g_x[7].t.r_d ),
    .X(_0852_));
 sg13g2_a21oi_1 _3774_ (.A1(_0830_),
    .A2(_0524_),
    .Y(_0853_),
    .B1(_0845_));
 sg13g2_or2_1 _3775_ (.X(_0854_),
    .B(_0273_),
    .A(_0524_));
 sg13g2_a22oi_1 _3776_ (.Y(_0855_),
    .B1(_0853_),
    .B2(_0854_),
    .A2(_0844_),
    .A1(_0845_));
 sg13g2_buf_1 _3777_ (.A(_0855_),
    .X(_0856_));
 sg13g2_inv_1 _3778_ (.Y(_0857_),
    .A(_0551_));
 sg13g2_a21oi_1 _3779_ (.A1(_0857_),
    .A2(_0774_),
    .Y(_0858_),
    .B1(net70));
 sg13g2_or2_1 _3780_ (.X(_0859_),
    .B(_0772_),
    .A(_0774_));
 sg13g2_a221oi_1 _3781_ (.B2(_0859_),
    .C1(net40),
    .B1(_0858_),
    .A1(net70),
    .Y(_0860_),
    .A2(_0835_));
 sg13g2_a21oi_1 _3782_ (.A1(net40),
    .A2(_0856_),
    .Y(_0861_),
    .B1(_0860_));
 sg13g2_a221oi_1 _3783_ (.B2(_0845_),
    .C1(_0524_),
    .B1(_0861_),
    .A1(_0849_),
    .Y(_0862_),
    .A2(_0851_));
 sg13g2_nand2_1 _3784_ (.Y(_0863_),
    .A(_0277_),
    .B(_0522_));
 sg13g2_and2_1 _3785_ (.A(_0279_),
    .B(_0281_),
    .X(_0864_));
 sg13g2_o21ai_1 _3786_ (.B1(_0864_),
    .Y(_0865_),
    .A1(_0269_),
    .A2(_0863_));
 sg13g2_a21oi_1 _3787_ (.A1(_0276_),
    .A2(_0529_),
    .Y(_0866_),
    .B1(_0279_));
 sg13g2_nand2b_1 _3788_ (.Y(_0867_),
    .B(_0866_),
    .A_N(_0286_));
 sg13g2_nand3_1 _3789_ (.B(_0865_),
    .C(_0867_),
    .A(_0524_),
    .Y(_0868_));
 sg13g2_nand2b_1 _3790_ (.Y(_0869_),
    .B(_0868_),
    .A_N(_0862_));
 sg13g2_or2_1 _3791_ (.X(_0870_),
    .B(_0316_),
    .A(_0335_));
 sg13g2_nor2_1 _3792_ (.A(\g.g_y[3].g_x[0].t.r_h ),
    .B(_0613_),
    .Y(_0871_));
 sg13g2_o21ai_1 _3793_ (.B1(_0871_),
    .Y(_0872_),
    .A1(_0611_),
    .A2(_0870_));
 sg13g2_a21oi_1 _3794_ (.A1(_0335_),
    .A2(_0316_),
    .Y(_0873_),
    .B1(_0311_));
 sg13g2_o21ai_1 _3795_ (.B1(_0873_),
    .Y(_0874_),
    .A1(_0589_),
    .A2(_0616_));
 sg13g2_nand3_1 _3796_ (.B(_0872_),
    .C(_0874_),
    .A(_0537_),
    .Y(_0875_));
 sg13g2_o21ai_1 _3797_ (.B1(_0801_),
    .Y(_0876_),
    .A1(_0547_),
    .A2(_0557_));
 sg13g2_and2_1 _3798_ (.A(_0546_),
    .B(_0802_),
    .X(_0877_));
 sg13g2_a221oi_1 _3799_ (.B2(\g.g_y[3].g_x[6].t.out_sc ),
    .C1(_0877_),
    .B1(_0803_),
    .A1(_0800_),
    .Y(_0878_),
    .A2(_0795_));
 sg13g2_nand3b_1 _3800_ (.B(_0876_),
    .C(_0878_),
    .Y(_0879_),
    .A_N(_0537_));
 sg13g2_nand3_1 _3801_ (.B(_0875_),
    .C(_0879_),
    .A(_0832_),
    .Y(_0880_));
 sg13g2_o21ai_1 _3802_ (.B1(_0880_),
    .Y(\g.g_y[3].g_x[7].t.w_dh ),
    .A1(_0832_),
    .A2(_0869_));
 sg13g2_nand3b_1 _3803_ (.B(_0872_),
    .C(_0874_),
    .Y(_0881_),
    .A_N(_0537_));
 sg13g2_nand3_1 _3804_ (.B(_0876_),
    .C(_0878_),
    .A(_0537_),
    .Y(_0882_));
 sg13g2_a22oi_1 _3805_ (.Y(_0883_),
    .B1(_0861_),
    .B2(_0845_),
    .A2(_0851_),
    .A1(_0849_));
 sg13g2_and3_1 _3806_ (.X(_0884_),
    .A(_0270_),
    .B(_0865_),
    .C(_0867_));
 sg13g2_a21oi_1 _3807_ (.A1(_0524_),
    .A2(_0883_),
    .Y(_0885_),
    .B1(_0884_));
 sg13g2_nand3_1 _3808_ (.B(_0882_),
    .C(_0885_),
    .A(_0881_),
    .Y(\g.g_y[3].g_x[7].t.w_na ));
 sg13g2_nand2_1 _3809_ (.Y(_0886_),
    .A(\g.g_y[3].g_x[6].t.out_sc ),
    .B(net47));
 sg13g2_nor2_1 _3810_ (.A(_0271_),
    .B(net74),
    .Y(_0887_));
 sg13g2_nand3b_1 _3811_ (.B(_0868_),
    .C(_0887_),
    .Y(_0888_),
    .A_N(_0862_));
 sg13g2_nand4_1 _3812_ (.B(_0113_),
    .C(_0875_),
    .A(_0271_),
    .Y(_0889_),
    .D(_0879_));
 sg13g2_nand3_1 _3813_ (.B(_0888_),
    .C(_0889_),
    .A(_0886_),
    .Y(\g.g_y[3].g_x[7].t.w_si ));
 sg13g2_buf_1 _3814_ (.A(\g.g_y[5].g_x[0].t.r_d ),
    .X(_0890_));
 sg13g2_inv_1 _3815_ (.Y(_0891_),
    .A(net39));
 sg13g2_mux2_1 _3816_ (.A0(_1869_),
    .A1(_1868_),
    .S(_1866_),
    .X(_0892_));
 sg13g2_buf_2 _3817_ (.A(_0892_),
    .X(_0893_));
 sg13g2_buf_1 _3818_ (.A(\g.g_y[5].g_x[0].t.r_v ),
    .X(_0894_));
 sg13g2_o21ai_1 _3819_ (.B1(net38),
    .Y(_0895_),
    .A1(_0891_),
    .A2(_0893_));
 sg13g2_buf_1 _3820_ (.A(\g.g_y[5].g_x[0].t.r_h ),
    .X(_0896_));
 sg13g2_inv_1 _3821_ (.Y(_0897_),
    .A(_0896_));
 sg13g2_buf_2 _3822_ (.A(\g.g_y[5].g_x[1].t.r_h ),
    .X(_0898_));
 sg13g2_mux2_1 _3823_ (.A0(\g.g_y[5].g_x[1].t.out_sc ),
    .A1(\g.g_y[5].g_x[1].t.r_gnl ),
    .S(_0637_),
    .X(_0899_));
 sg13g2_nand2b_1 _3824_ (.Y(_0900_),
    .B(_0898_),
    .A_N(_0636_));
 sg13g2_o21ai_1 _3825_ (.B1(_0900_),
    .Y(_0901_),
    .A1(_0898_),
    .A2(_0899_));
 sg13g2_buf_1 _3826_ (.A(_0901_),
    .X(_0902_));
 sg13g2_nor2b_1 _3827_ (.A(_0896_),
    .B_N(net6),
    .Y(_0903_));
 sg13g2_nor2_1 _3828_ (.A(net39),
    .B(_0903_),
    .Y(_0904_));
 sg13g2_o21ai_1 _3829_ (.B1(_0904_),
    .Y(_0905_),
    .A1(_0897_),
    .A2(_0902_));
 sg13g2_nand2b_1 _3830_ (.Y(_0906_),
    .B(_0905_),
    .A_N(_0895_));
 sg13g2_inv_1 _3831_ (.Y(_0907_),
    .A(net6));
 sg13g2_mux2_1 _3832_ (.A0(_0907_),
    .A1(_0902_),
    .S(_0897_),
    .X(_0908_));
 sg13g2_nand2_1 _3833_ (.Y(_0909_),
    .A(_0891_),
    .B(_0893_));
 sg13g2_nand2b_1 _3834_ (.Y(_0910_),
    .B(net39),
    .A_N(\g.g_y[5].g_x[0].t.out_sc ));
 sg13g2_nor2b_1 _3835_ (.A(net38),
    .B_N(_0910_),
    .Y(_0911_));
 sg13g2_o21ai_1 _3836_ (.B1(_0911_),
    .Y(_0912_),
    .A1(_0908_),
    .A2(_0909_));
 sg13g2_nand3_1 _3837_ (.B(_0906_),
    .C(_0912_),
    .A(_0321_),
    .Y(_0913_));
 sg13g2_inv_1 _3838_ (.Y(_0914_),
    .A(_0321_));
 sg13g2_a21oi_1 _3839_ (.A1(_0317_),
    .A2(_0588_),
    .Y(_0915_),
    .B1(_0329_));
 sg13g2_nand2_1 _3840_ (.Y(_0916_),
    .A(_0320_),
    .B(_0915_));
 sg13g2_nand2b_1 _3841_ (.Y(_0917_),
    .B(_0335_),
    .A_N(_0588_));
 sg13g2_and2_1 _3842_ (.A(_0329_),
    .B(_0337_),
    .X(_0918_));
 sg13g2_o21ai_1 _3843_ (.B1(_0918_),
    .Y(_0919_),
    .A1(_0334_),
    .A2(_0917_));
 sg13g2_nand3_1 _3844_ (.B(_0916_),
    .C(_0919_),
    .A(_0914_),
    .Y(_0920_));
 sg13g2_and3_1 _3845_ (.X(_0921_),
    .A(_0322_),
    .B(_0913_),
    .C(_0920_));
 sg13g2_nand3_1 _3846_ (.B(_0633_),
    .C(_0645_),
    .A(_0621_),
    .Y(_0922_));
 sg13g2_nor2_1 _3847_ (.A(_0621_),
    .B(\g.g_y[4].g_x[1].t.out_sc ),
    .Y(_0923_));
 sg13g2_nor2_1 _3848_ (.A(_0631_),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_o21ai_1 _3849_ (.B1(_0631_),
    .Y(_0925_),
    .A1(_0621_),
    .A2(_0630_));
 sg13g2_o21ai_1 _3850_ (.B1(_0624_),
    .Y(_0926_),
    .A1(_0653_),
    .A2(_0925_));
 sg13g2_a21oi_1 _3851_ (.A1(_0922_),
    .A2(_0924_),
    .Y(_0927_),
    .B1(_0926_));
 sg13g2_nor2_1 _3852_ (.A(_0624_),
    .B(net5),
    .Y(_0928_));
 sg13g2_nor3_1 _3853_ (.A(_0322_),
    .B(_0927_),
    .C(_0928_),
    .Y(_0929_));
 sg13g2_or2_1 _3854_ (.X(\g.g_y[4].g_x[0].t.w_dh ),
    .B(_0929_),
    .A(_0921_));
 sg13g2_a21oi_1 _3855_ (.A1(_0916_),
    .A2(_0919_),
    .Y(_0930_),
    .B1(_0914_));
 sg13g2_a21oi_1 _3856_ (.A1(_0906_),
    .A2(_0912_),
    .Y(_0931_),
    .B1(_0321_));
 sg13g2_nor2_1 _3857_ (.A(_0653_),
    .B(_0925_),
    .Y(_0932_));
 sg13g2_a21oi_1 _3858_ (.A1(_0922_),
    .A2(_0924_),
    .Y(_0933_),
    .B1(_0932_));
 sg13g2_nand2_1 _3859_ (.Y(_0934_),
    .A(_0624_),
    .B(net5));
 sg13g2_o21ai_1 _3860_ (.B1(_0934_),
    .Y(_0935_),
    .A1(_0624_),
    .A2(_0933_));
 sg13g2_o21ai_1 _3861_ (.B1(_0935_),
    .Y(\g.g_y[4].g_x[0].t.w_na ),
    .A1(_0930_),
    .A2(_0931_));
 sg13g2_nand2_1 _3862_ (.Y(_0936_),
    .A(\g.g_y[3].g_x[7].t.out_sc ),
    .B(_0109_));
 sg13g2_inv_1 _3863_ (.Y(_0937_),
    .A(_0322_));
 sg13g2_or4_1 _3864_ (.A(_0937_),
    .B(net74),
    .C(_0927_),
    .D(_0928_),
    .X(_0938_));
 sg13g2_nand4_1 _3865_ (.B(_0113_),
    .C(_0913_),
    .A(_0937_),
    .Y(_0939_),
    .D(_0920_));
 sg13g2_nand3_1 _3866_ (.B(_0938_),
    .C(_0939_),
    .A(_0936_),
    .Y(\g.g_y[4].g_x[0].t.w_si ));
 sg13g2_a22oi_1 _3867_ (.Y(_0940_),
    .B1(_0649_),
    .B2(_0651_),
    .A2(_0635_),
    .A1(_0644_));
 sg13g2_a221oi_1 _3868_ (.B2(_0656_),
    .C1(_0622_),
    .B1(_0654_),
    .A1(_0632_),
    .Y(_0941_),
    .A2(_0626_));
 sg13g2_a21oi_1 _3869_ (.A1(_0622_),
    .A2(_0940_),
    .Y(_0942_),
    .B1(_0941_));
 sg13g2_mux2_1 _3870_ (.A0(\g.g_y[4].g_x[0].t.out_sc ),
    .A1(_0942_),
    .S(net64),
    .X(\g.g_y[4].g_x[1].t.w_si ));
 sg13g2_nand2_1 _3871_ (.Y(_0943_),
    .A(_0415_),
    .B(_0598_));
 sg13g2_or3_1 _3872_ (.A(_0394_),
    .B(_0404_),
    .C(_0943_),
    .X(_0944_));
 sg13g2_nand2_1 _3873_ (.Y(_0945_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_a21oi_1 _3874_ (.A1(_0394_),
    .A2(_0598_),
    .Y(_0946_),
    .B1(_0415_));
 sg13g2_o21ai_1 _3875_ (.B1(_0946_),
    .Y(_0947_),
    .A1(net26),
    .A2(_0418_));
 sg13g2_nand4_1 _3876_ (.B(_0944_),
    .C(_0945_),
    .A(_0409_),
    .Y(_0948_),
    .D(_0947_));
 sg13g2_buf_1 _3877_ (.A(\g.g_y[5].g_x[2].t.r_d ),
    .X(_0949_));
 sg13g2_inv_1 _3878_ (.Y(_0950_),
    .A(net37));
 sg13g2_mux2_1 _3879_ (.A0(\g.g_y[5].g_x[3].t.out_sc ),
    .A1(\g.g_y[5].g_x[3].t.r_gnl ),
    .S(_0697_),
    .X(_0951_));
 sg13g2_buf_2 _3880_ (.A(\g.g_y[5].g_x[3].t.r_h ),
    .X(_0952_));
 sg13g2_inv_1 _3881_ (.Y(_0953_),
    .A(_0952_));
 sg13g2_nand2b_1 _3882_ (.Y(_0954_),
    .B(_0953_),
    .A_N(_0951_));
 sg13g2_buf_1 _3883_ (.A(\g.g_y[5].g_x[2].t.r_h ),
    .X(_0955_));
 sg13g2_nand2b_1 _3884_ (.Y(_0956_),
    .B(_0952_),
    .A_N(_0702_));
 sg13g2_and2_1 _3885_ (.A(_0955_),
    .B(_0956_),
    .X(_0957_));
 sg13g2_mux2_1 _3886_ (.A0(_0636_),
    .A1(_0899_),
    .S(_0898_),
    .X(_0958_));
 sg13g2_inv_1 _3887_ (.Y(_0959_),
    .A(_0955_));
 sg13g2_a22oi_1 _3888_ (.Y(_0960_),
    .B1(_0958_),
    .B2(_0959_),
    .A2(_0957_),
    .A1(_0954_));
 sg13g2_mux2_1 _3889_ (.A0(_1951_),
    .A1(_1949_),
    .S(_1952_),
    .X(_0961_));
 sg13g2_buf_1 _3890_ (.A(\g.g_y[5].g_x[2].t.r_v ),
    .X(_0962_));
 sg13g2_o21ai_1 _3891_ (.B1(_0962_),
    .Y(_0963_),
    .A1(_0950_),
    .A2(_0961_));
 sg13g2_a21o_1 _3892_ (.A2(_0960_),
    .A1(_0950_),
    .B1(_0963_),
    .X(_0964_));
 sg13g2_and2_1 _3893_ (.A(_0959_),
    .B(_0956_),
    .X(_0965_));
 sg13g2_a22oi_1 _3894_ (.Y(_0966_),
    .B1(_0965_),
    .B2(_0954_),
    .A2(_0958_),
    .A1(_0955_));
 sg13g2_buf_1 _3895_ (.A(_0966_),
    .X(_0967_));
 sg13g2_inv_1 _3896_ (.Y(_0968_),
    .A(_0962_));
 sg13g2_nand3_1 _3897_ (.B(_0950_),
    .C(_0961_),
    .A(_0968_),
    .Y(_0969_));
 sg13g2_o21ai_1 _3898_ (.B1(_0968_),
    .Y(_0970_),
    .A1(_0967_),
    .A2(_0969_));
 sg13g2_nand2b_1 _3899_ (.Y(_0971_),
    .B(net37),
    .A_N(\g.g_y[5].g_x[2].t.out_sc ));
 sg13g2_o21ai_1 _3900_ (.B1(_0408_),
    .Y(_0972_),
    .A1(_0962_),
    .A2(_0971_));
 sg13g2_a21o_1 _3901_ (.A2(_0970_),
    .A1(_0964_),
    .B1(_0972_),
    .X(_0973_));
 sg13g2_inv_1 _3902_ (.Y(_0974_),
    .A(_0405_));
 sg13g2_a21oi_1 _3903_ (.A1(_0948_),
    .A2(_0973_),
    .Y(_0975_),
    .B1(_0974_));
 sg13g2_nor2_1 _3904_ (.A(_0692_),
    .B(_0714_),
    .Y(_0976_));
 sg13g2_o21ai_1 _3905_ (.B1(_0976_),
    .Y(_0977_),
    .A1(_0696_),
    .A2(_0707_));
 sg13g2_mux2_1 _3906_ (.A0(_0702_),
    .A1(_0698_),
    .S(_0700_),
    .X(_0978_));
 sg13g2_mux2_1 _3907_ (.A0(_0978_),
    .A1(_0706_),
    .S(_0710_),
    .X(_0979_));
 sg13g2_nor2_1 _3908_ (.A(_0716_),
    .B(_0714_),
    .Y(_0980_));
 sg13g2_nand2_1 _3909_ (.Y(_0981_),
    .A(_0979_),
    .B(_0980_));
 sg13g2_nor2_1 _3910_ (.A(_0688_),
    .B(_0687_),
    .Y(_0982_));
 sg13g2_a21oi_1 _3911_ (.A1(_0691_),
    .A2(_0688_),
    .Y(_0983_),
    .B1(_0982_));
 sg13g2_nor2_1 _3912_ (.A(_0716_),
    .B(_0685_),
    .Y(_0984_));
 sg13g2_nor2_1 _3913_ (.A(_0692_),
    .B(_0685_),
    .Y(_0985_));
 sg13g2_a22oi_1 _3914_ (.Y(_0986_),
    .B1(_0985_),
    .B2(\g.g_y[4].g_x[3].t.out_sc ),
    .A2(_0984_),
    .A1(_0983_));
 sg13g2_nand4_1 _3915_ (.B(_0977_),
    .C(_0981_),
    .A(_0628_),
    .Y(_0987_),
    .D(_0986_));
 sg13g2_and4_1 _3916_ (.A(_0631_),
    .B(_0621_),
    .C(_0626_),
    .D(_0645_),
    .X(_0988_));
 sg13g2_nor2_1 _3917_ (.A(_0631_),
    .B(_0622_),
    .Y(_0989_));
 sg13g2_nand2_1 _3918_ (.Y(_0990_),
    .A(_0632_),
    .B(_0622_));
 sg13g2_nand2_1 _3919_ (.Y(_0991_),
    .A(_0631_),
    .B(_0923_));
 sg13g2_o21ai_1 _3920_ (.B1(_0991_),
    .Y(_0992_),
    .A1(_0626_),
    .A2(_0990_));
 sg13g2_a21o_1 _3921_ (.A2(_0989_),
    .A1(_0940_),
    .B1(_0992_),
    .X(_0993_));
 sg13g2_o21ai_1 _3922_ (.B1(_0629_),
    .Y(_0994_),
    .A1(_0988_),
    .A2(_0993_));
 sg13g2_nand3_1 _3923_ (.B(_0987_),
    .C(_0994_),
    .A(_0974_),
    .Y(_0995_));
 sg13g2_nand2b_1 _3924_ (.Y(\g.g_y[4].g_x[2].t.w_dh ),
    .B(_0995_),
    .A_N(_0975_));
 sg13g2_nand4_1 _3925_ (.B(_0977_),
    .C(_0981_),
    .A(_0629_),
    .Y(_0996_),
    .D(_0986_));
 sg13g2_o21ai_1 _3926_ (.B1(_0628_),
    .Y(_0997_),
    .A1(_0988_),
    .A2(_0993_));
 sg13g2_nand3_1 _3927_ (.B(_0945_),
    .C(_0947_),
    .A(_0944_),
    .Y(_0998_));
 sg13g2_nand2_1 _3928_ (.Y(_0999_),
    .A(_0408_),
    .B(_0998_));
 sg13g2_nand2b_1 _3929_ (.Y(_1000_),
    .B(_1952_),
    .A_N(_1949_));
 sg13g2_o21ai_1 _3930_ (.B1(_1000_),
    .Y(_1001_),
    .A1(_1952_),
    .A2(_1951_));
 sg13g2_or2_1 _3931_ (.X(_1002_),
    .B(_0408_),
    .A(_0411_));
 sg13g2_o21ai_1 _3932_ (.B1(_1002_),
    .Y(_1003_),
    .A1(_0409_),
    .A2(_0407_));
 sg13g2_mux2_1 _3933_ (.A0(_1001_),
    .A1(_1003_),
    .S(_0962_),
    .X(_1004_));
 sg13g2_nor3_1 _3934_ (.A(net37),
    .B(_0967_),
    .C(_1004_),
    .Y(_1005_));
 sg13g2_nand2_1 _3935_ (.Y(_1006_),
    .A(_0968_),
    .B(_0971_));
 sg13g2_o21ai_1 _3936_ (.B1(_0964_),
    .Y(_1007_),
    .A1(_1005_),
    .A2(_1006_));
 sg13g2_nand2b_1 _3937_ (.Y(_1008_),
    .B(_0409_),
    .A_N(_1007_));
 sg13g2_nand4_1 _3938_ (.B(_0997_),
    .C(_0999_),
    .A(_0996_),
    .Y(\g.g_y[4].g_x[2].t.w_na ),
    .D(_1008_));
 sg13g2_buf_1 _3939_ (.A(net77),
    .X(_1009_));
 sg13g2_nand2_1 _3940_ (.Y(_1010_),
    .A(\g.g_y[4].g_x[1].t.out_sc ),
    .B(net36));
 sg13g2_nand4_1 _3941_ (.B(net45),
    .C(_0987_),
    .A(_0405_),
    .Y(_1011_),
    .D(_0994_));
 sg13g2_nand2_1 _3942_ (.Y(_1012_),
    .A(_0974_),
    .B(net81));
 sg13g2_a21o_1 _3943_ (.A2(_0973_),
    .A1(_0948_),
    .B1(_1012_),
    .X(_1013_));
 sg13g2_nand3_1 _3944_ (.B(_1011_),
    .C(_1013_),
    .A(_1010_),
    .Y(\g.g_y[4].g_x[2].t.w_si ));
 sg13g2_nand2_1 _3945_ (.Y(_1014_),
    .A(_0690_),
    .B(_0717_));
 sg13g2_nand2_1 _3946_ (.Y(_1015_),
    .A(_0716_),
    .B(_0695_));
 sg13g2_nand3_1 _3947_ (.B(_1014_),
    .C(_1015_),
    .A(_0685_),
    .Y(_1016_));
 sg13g2_o21ai_1 _3948_ (.B1(_1016_),
    .Y(_1017_),
    .A1(_0685_),
    .A2(_0979_));
 sg13g2_nand2_1 _3949_ (.Y(_1018_),
    .A(\g.g_y[4].g_x[2].t.out_sc ),
    .B(net41));
 sg13g2_o21ai_1 _3950_ (.B1(_1018_),
    .Y(\g.g_y[4].g_x[3].t.w_si ),
    .A1(net42),
    .A2(_1017_));
 sg13g2_nand3_1 _3951_ (.B(_0784_),
    .C(_0815_),
    .A(_0765_),
    .Y(_1019_));
 sg13g2_buf_1 _3952_ (.A(_1019_),
    .X(_1020_));
 sg13g2_nor2_1 _3953_ (.A(_0765_),
    .B(\g.g_y[4].g_x[5].t.out_sc ),
    .Y(_1021_));
 sg13g2_nor2_1 _3954_ (.A(_0770_),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_o21ai_1 _3955_ (.B1(_0770_),
    .Y(_1023_),
    .A1(_0765_),
    .A2(_0776_));
 sg13g2_o21ai_1 _3956_ (.B1(_0688_),
    .Y(_1024_),
    .A1(_0768_),
    .A2(_1023_));
 sg13g2_a21o_1 _3957_ (.A2(_1022_),
    .A1(_1020_),
    .B1(_1024_),
    .X(_1025_));
 sg13g2_o21ai_1 _3958_ (.B1(_0980_),
    .Y(_1026_),
    .A1(_0696_),
    .A2(_0707_));
 sg13g2_nand2_1 _3959_ (.Y(_1027_),
    .A(_0979_),
    .B(_0976_));
 sg13g2_a22oi_1 _3960_ (.Y(_1028_),
    .B1(_0985_),
    .B2(_0695_),
    .A2(_0984_),
    .A1(\g.g_y[4].g_x[3].t.out_sc ));
 sg13g2_nand4_1 _3961_ (.B(_1026_),
    .C(_1027_),
    .A(_0689_),
    .Y(_1029_),
    .D(_1028_));
 sg13g2_nand2_1 _3962_ (.Y(_1030_),
    .A(_1025_),
    .B(_1029_));
 sg13g2_or3_1 _3963_ (.A(_0454_),
    .B(_0476_),
    .C(_0503_),
    .X(_1031_));
 sg13g2_nand3_1 _3964_ (.B(_0457_),
    .C(_0490_),
    .A(net44),
    .Y(_1032_));
 sg13g2_o21ai_1 _3965_ (.B1(net44),
    .Y(_1033_),
    .A1(_0488_),
    .A2(_1032_));
 sg13g2_nand3b_1 _3966_ (.B(_1031_),
    .C(_1033_),
    .Y(_1034_),
    .A_N(net43));
 sg13g2_buf_2 _3967_ (.A(\g.g_y[5].g_x[4].t.r_v ),
    .X(_1035_));
 sg13g2_inv_2 _3968_ (.Y(_1036_),
    .A(_1035_));
 sg13g2_buf_2 _3969_ (.A(\g.g_y[5].g_x[4].t.r_d ),
    .X(_1037_));
 sg13g2_buf_1 _3970_ (.A(\g.g_y[5].g_x[4].t.r_h ),
    .X(_1038_));
 sg13g2_inv_1 _3971_ (.Y(_1039_),
    .A(_1038_));
 sg13g2_mux2_1 _3972_ (.A0(\g.g_y[5].g_x[5].t.out_sc ),
    .A1(\g.g_y[5].g_x[5].t.r_gnl ),
    .S(_0756_),
    .X(_1040_));
 sg13g2_buf_2 _3973_ (.A(_1040_),
    .X(_1041_));
 sg13g2_buf_2 _3974_ (.A(\g.g_y[5].g_x[5].t.r_h ),
    .X(_1042_));
 sg13g2_inv_1 _3975_ (.Y(_1043_),
    .A(_1042_));
 sg13g2_mux2_1 _3976_ (.A0(_0762_),
    .A1(_1041_),
    .S(_1043_),
    .X(_1044_));
 sg13g2_or2_1 _3977_ (.X(_1045_),
    .B(_0951_),
    .A(_0953_));
 sg13g2_buf_1 _3978_ (.A(_1045_),
    .X(_1046_));
 sg13g2_nor2_1 _3979_ (.A(_0702_),
    .B(_0952_),
    .Y(_1047_));
 sg13g2_nor2_1 _3980_ (.A(_1039_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_a22oi_1 _3981_ (.Y(_1049_),
    .B1(_1046_),
    .B2(_1048_),
    .A2(_1044_),
    .A1(_1039_));
 sg13g2_mux2_1 _3982_ (.A0(_0479_),
    .A1(_0478_),
    .S(\g.g_y[4].g_x[4].t.r_v ),
    .X(_1050_));
 sg13g2_inv_1 _3983_ (.Y(_1051_),
    .A(_2105_));
 sg13g2_nand2b_1 _3984_ (.Y(_1052_),
    .B(_1051_),
    .A_N(_2104_));
 sg13g2_nand2b_1 _3985_ (.Y(_1053_),
    .B(_2105_),
    .A_N(_2102_));
 sg13g2_and2_1 _3986_ (.A(_1036_),
    .B(_1053_),
    .X(_1054_));
 sg13g2_a22oi_1 _3987_ (.Y(_1055_),
    .B1(_1052_),
    .B2(_1054_),
    .A2(_1050_),
    .A1(_1035_));
 sg13g2_buf_1 _3988_ (.A(_1055_),
    .X(_1056_));
 sg13g2_nor3_2 _3989_ (.A(_1037_),
    .B(_1049_),
    .C(_1056_),
    .Y(_1057_));
 sg13g2_nand3_1 _3990_ (.B(_1036_),
    .C(_1057_),
    .A(net43),
    .Y(_1058_));
 sg13g2_and2_1 _3991_ (.A(net43),
    .B(_1035_),
    .X(_1059_));
 sg13g2_and2_1 _3992_ (.A(_1035_),
    .B(_1053_),
    .X(_1060_));
 sg13g2_inv_1 _3993_ (.Y(_1061_),
    .A(_1037_));
 sg13g2_a221oi_1 _3994_ (.B2(_1060_),
    .C1(_1061_),
    .B1(_1052_),
    .A1(_1036_),
    .Y(_1062_),
    .A2(_1050_));
 sg13g2_buf_1 _3995_ (.A(_1062_),
    .X(_1063_));
 sg13g2_nor2_1 _3996_ (.A(_1038_),
    .B(_1047_),
    .Y(_1064_));
 sg13g2_a221oi_1 _3997_ (.B2(_1064_),
    .C1(_1037_),
    .B1(_1046_),
    .A1(_1038_),
    .Y(_1065_),
    .A2(_1044_));
 sg13g2_or2_1 _3998_ (.X(_1066_),
    .B(_1065_),
    .A(_1063_));
 sg13g2_buf_1 _3999_ (.A(_1066_),
    .X(_1067_));
 sg13g2_nand2_1 _4000_ (.Y(_1068_),
    .A(net44),
    .B(_0459_));
 sg13g2_nor2_2 _4001_ (.A(_1061_),
    .B(\g.g_y[5].g_x[4].t.out_sc ),
    .Y(_1069_));
 sg13g2_nand3_1 _4002_ (.B(_1036_),
    .C(_1069_),
    .A(net43),
    .Y(_1070_));
 sg13g2_o21ai_1 _4003_ (.B1(_1070_),
    .Y(_1071_),
    .A1(_0480_),
    .A2(_1068_));
 sg13g2_a21oi_1 _4004_ (.A1(_1059_),
    .A2(_1067_),
    .Y(_1072_),
    .B1(_1071_));
 sg13g2_nand4_1 _4005_ (.B(_1034_),
    .C(_1058_),
    .A(_0477_),
    .Y(_1073_),
    .D(_1072_));
 sg13g2_o21ai_1 _4006_ (.B1(_1073_),
    .Y(\g.g_y[4].g_x[4].t.w_dh ),
    .A1(_0477_),
    .A2(_1030_));
 sg13g2_nor2_1 _4007_ (.A(_1036_),
    .B(_1067_),
    .Y(_1074_));
 sg13g2_nor3_1 _4008_ (.A(_1035_),
    .B(_1069_),
    .C(_1057_),
    .Y(_1075_));
 sg13g2_or3_1 _4009_ (.A(_0480_),
    .B(_1074_),
    .C(_1075_),
    .X(_1076_));
 sg13g2_nor3_1 _4010_ (.A(_0455_),
    .B(_0495_),
    .C(_0459_),
    .Y(_1077_));
 sg13g2_nand3b_1 _4011_ (.B(net43),
    .C(_1031_),
    .Y(_1078_),
    .A_N(_1077_));
 sg13g2_nor2_1 _4012_ (.A(_0768_),
    .B(_1023_),
    .Y(_1079_));
 sg13g2_a21o_1 _4013_ (.A2(_1022_),
    .A1(_1020_),
    .B1(_1079_),
    .X(_1080_));
 sg13g2_nand3_1 _4014_ (.B(_1027_),
    .C(_1028_),
    .A(_1026_),
    .Y(_1081_));
 sg13g2_mux2_1 _4015_ (.A0(_1080_),
    .A1(_1081_),
    .S(_0688_),
    .X(_1082_));
 sg13g2_nand3_1 _4016_ (.B(_1078_),
    .C(_1082_),
    .A(_1076_),
    .Y(\g.g_y[4].g_x[4].t.w_na ));
 sg13g2_nand2_1 _4017_ (.Y(_1083_),
    .A(\g.g_y[4].g_x[3].t.out_sc ),
    .B(net36));
 sg13g2_nor2_1 _4018_ (.A(_0477_),
    .B(net77),
    .Y(_1084_));
 sg13g2_nand4_1 _4019_ (.B(_1058_),
    .C(_1072_),
    .A(_1034_),
    .Y(_1085_),
    .D(_1084_));
 sg13g2_nand4_1 _4020_ (.B(net73),
    .C(_1025_),
    .A(_0477_),
    .Y(_1086_),
    .D(_1029_));
 sg13g2_nand3_1 _4021_ (.B(_1085_),
    .C(_1086_),
    .A(_1083_),
    .Y(\g.g_y[4].g_x[4].t.w_si ));
 sg13g2_a221oi_1 _4022_ (.B2(_0770_),
    .C1(_0766_),
    .B1(_0776_),
    .A1(_0769_),
    .Y(_1087_),
    .A2(_0771_));
 sg13g2_a221oi_1 _4023_ (.B2(_0764_),
    .C1(_0765_),
    .B1(_0761_),
    .A1(_0754_),
    .Y(_1088_),
    .A2(_0755_));
 sg13g2_nor3_1 _4024_ (.A(net82),
    .B(_1087_),
    .C(_1088_),
    .Y(_1089_));
 sg13g2_a21o_1 _4025_ (.A2(net59),
    .A1(\g.g_y[4].g_x[4].t.out_sc ),
    .B1(_1089_),
    .X(\g.g_y[4].g_x[5].t.w_si ));
 sg13g2_buf_1 _4026_ (.A(\g.g_y[5].g_x[6].t.r_d ),
    .X(_1090_));
 sg13g2_inv_1 _4027_ (.Y(_1091_),
    .A(_1090_));
 sg13g2_mux2_1 _4028_ (.A0(\g.g_y[5].g_x[7].t.out_sc ),
    .A1(\g.g_y[5].g_x[7].t.r_gnl ),
    .S(_0841_),
    .X(_1092_));
 sg13g2_buf_2 _4029_ (.A(\g.g_y[5].g_x[7].t.r_h ),
    .X(_1093_));
 sg13g2_mux2_1 _4030_ (.A0(_1092_),
    .A1(\g.g_y[5].g_x[7].t.r_ghl ),
    .S(_1093_),
    .X(_1094_));
 sg13g2_buf_1 _4031_ (.A(_1094_),
    .X(_1095_));
 sg13g2_mux2_1 _4032_ (.A0(_0762_),
    .A1(_1041_),
    .S(_1042_),
    .X(_1096_));
 sg13g2_buf_1 _4033_ (.A(\g.g_y[5].g_x[6].t.r_h ),
    .X(_1097_));
 sg13g2_mux2_1 _4034_ (.A0(_1095_),
    .A1(_1096_),
    .S(net69),
    .X(_1098_));
 sg13g2_buf_1 _4035_ (.A(_1098_),
    .X(_1099_));
 sg13g2_mux2_1 _4036_ (.A0(_0551_),
    .A1(_0550_),
    .S(_0548_),
    .X(_1100_));
 sg13g2_buf_1 _4037_ (.A(_1100_),
    .X(_1101_));
 sg13g2_mux2_1 _4038_ (.A0(_2264_),
    .A1(_2262_),
    .S(_2259_),
    .X(_1102_));
 sg13g2_buf_2 _4039_ (.A(\g.g_y[5].g_x[6].t.r_v ),
    .X(_1103_));
 sg13g2_inv_2 _4040_ (.Y(_1104_),
    .A(_1103_));
 sg13g2_mux2_1 _4041_ (.A0(_1101_),
    .A1(_1102_),
    .S(_1104_),
    .X(_1105_));
 sg13g2_nand3_1 _4042_ (.B(_1099_),
    .C(_1105_),
    .A(_1091_),
    .Y(_1106_));
 sg13g2_nand2b_1 _4043_ (.Y(_1107_),
    .B(_1090_),
    .A_N(\g.g_y[5].g_x[6].t.out_sc ));
 sg13g2_and2_1 _4044_ (.A(_1104_),
    .B(_1107_),
    .X(_1108_));
 sg13g2_a21oi_1 _4045_ (.A1(_0763_),
    .A2(_1043_),
    .Y(_1109_),
    .B1(net69));
 sg13g2_or2_1 _4046_ (.X(_1110_),
    .B(_1041_),
    .A(_1043_));
 sg13g2_a221oi_1 _4047_ (.B2(_1110_),
    .C1(net35),
    .B1(_1109_),
    .A1(net69),
    .Y(_1111_),
    .A2(_1095_));
 sg13g2_nand2b_1 _4048_ (.Y(_1112_),
    .B(_2259_),
    .A_N(_2262_));
 sg13g2_inv_1 _4049_ (.Y(_1113_),
    .A(_2264_));
 sg13g2_a21oi_1 _4050_ (.A1(_1113_),
    .A2(net49),
    .Y(_1114_),
    .B1(_1104_));
 sg13g2_a221oi_1 _4051_ (.B2(_1114_),
    .C1(_1091_),
    .B1(_1112_),
    .A1(_1104_),
    .Y(_1115_),
    .A2(_1101_));
 sg13g2_buf_1 _4052_ (.A(_1115_),
    .X(_1116_));
 sg13g2_nor2_1 _4053_ (.A(_1111_),
    .B(_1116_),
    .Y(_1117_));
 sg13g2_a221oi_1 _4054_ (.B2(_1103_),
    .C1(_0797_),
    .B1(_1117_),
    .A1(_1106_),
    .Y(_1118_),
    .A2(_1108_));
 sg13g2_and2_1 _4055_ (.A(_0556_),
    .B(_0561_),
    .X(_1119_));
 sg13g2_a221oi_1 _4056_ (.B2(_0559_),
    .C1(_0548_),
    .B1(_1119_),
    .A1(_0560_),
    .Y(_1120_),
    .A2(_0566_));
 sg13g2_o21ai_1 _4057_ (.B1(_0549_),
    .Y(_1121_),
    .A1(_1118_),
    .A2(_1120_));
 sg13g2_nand2b_1 _4058_ (.Y(_1122_),
    .B(net40),
    .A_N(_0837_));
 sg13g2_a21oi_1 _4059_ (.A1(_0839_),
    .A2(_0848_),
    .Y(_1123_),
    .B1(_1122_));
 sg13g2_nand2_1 _4060_ (.Y(_1124_),
    .A(net70),
    .B(net40));
 sg13g2_nor2b_1 _4061_ (.A(net40),
    .B_N(net70),
    .Y(_1125_));
 sg13g2_nor2_1 _4062_ (.A(net70),
    .B(net40),
    .Y(_1126_));
 sg13g2_a22oi_1 _4063_ (.Y(_1127_),
    .B1(_1126_),
    .B2(\g.g_y[4].g_x[7].t.out_sc ),
    .A2(_1125_),
    .A1(_0835_));
 sg13g2_o21ai_1 _4064_ (.B1(_1127_),
    .Y(_1128_),
    .A1(_0856_),
    .A2(_1124_));
 sg13g2_o21ai_1 _4065_ (.B1(_0773_),
    .Y(_1129_),
    .A1(_1123_),
    .A2(_1128_));
 sg13g2_nor3_1 _4066_ (.A(_0773_),
    .B(_0783_),
    .C(_1021_),
    .Y(_1130_));
 sg13g2_nor2_1 _4067_ (.A(_0765_),
    .B(_0782_),
    .Y(_1131_));
 sg13g2_nor4_1 _4068_ (.A(_0773_),
    .B(_0770_),
    .C(_0768_),
    .D(_1131_),
    .Y(_1132_));
 sg13g2_a21oi_1 _4069_ (.A1(_1020_),
    .A2(_1130_),
    .Y(_1133_),
    .B1(_1132_));
 sg13g2_nand3b_1 _4070_ (.B(_1129_),
    .C(_1133_),
    .Y(_1134_),
    .A_N(_0549_));
 sg13g2_and2_1 _4071_ (.A(_1121_),
    .B(_1134_),
    .X(\g.g_y[4].g_x[6].t.w_dh ));
 sg13g2_nor3_1 _4072_ (.A(_0773_),
    .B(_1123_),
    .C(_1128_),
    .Y(_1135_));
 sg13g2_nor2_1 _4073_ (.A(_0768_),
    .B(_0777_),
    .Y(_1136_));
 sg13g2_nor2_1 _4074_ (.A(_0783_),
    .B(_1021_),
    .Y(_1137_));
 sg13g2_a221oi_1 _4075_ (.B2(_1137_),
    .C1(_0774_),
    .B1(_1020_),
    .A1(_0783_),
    .Y(_1138_),
    .A2(_1136_));
 sg13g2_a221oi_1 _4076_ (.B2(_1103_),
    .C1(_0548_),
    .B1(_1117_),
    .A1(_1106_),
    .Y(_1139_),
    .A2(_1108_));
 sg13g2_a221oi_1 _4077_ (.B2(_0559_),
    .C1(_0797_),
    .B1(_1119_),
    .A1(_0560_),
    .Y(_1140_),
    .A2(_0566_));
 sg13g2_or4_1 _4078_ (.A(_1135_),
    .B(_1138_),
    .C(_1139_),
    .D(_1140_),
    .X(\g.g_y[4].g_x[6].t.w_na ));
 sg13g2_and2_1 _4079_ (.A(\g.g_y[4].g_x[5].t.out_sc ),
    .B(_2034_),
    .X(_1141_));
 sg13g2_nor4_1 _4080_ (.A(_0549_),
    .B(net78),
    .C(_1118_),
    .D(_1120_),
    .Y(_1142_));
 sg13g2_nand2_1 _4081_ (.Y(_1143_),
    .A(_0549_),
    .B(net81));
 sg13g2_a21oi_1 _4082_ (.A1(_1129_),
    .A2(_1133_),
    .Y(_1144_),
    .B1(_1143_));
 sg13g2_or3_1 _4083_ (.A(_1141_),
    .B(_1142_),
    .C(_1144_),
    .X(\g.g_y[4].g_x[6].t.w_si ));
 sg13g2_a21o_1 _4084_ (.A2(_0856_),
    .A1(net40),
    .B1(_0860_),
    .X(_1145_));
 sg13g2_nand3_1 _4085_ (.B(_0839_),
    .C(_0848_),
    .A(_0852_),
    .Y(_1146_));
 sg13g2_or2_1 _4086_ (.X(_1147_),
    .B(\g.g_y[4].g_x[7].t.out_sc ),
    .A(_0852_));
 sg13g2_nand3_1 _4087_ (.B(_1146_),
    .C(_1147_),
    .A(net70),
    .Y(_1148_));
 sg13g2_o21ai_1 _4088_ (.B1(_1148_),
    .Y(\g.g_y[4].g_x[7].t.out_r ),
    .A1(_0837_),
    .A2(_1145_));
 sg13g2_a22oi_1 _4089_ (.Y(_1149_),
    .B1(_0858_),
    .B2(_0859_),
    .A2(_0835_),
    .A1(net70));
 sg13g2_mux2_1 _4090_ (.A0(_0856_),
    .A1(_1149_),
    .S(net40),
    .X(_1150_));
 sg13g2_nand2_1 _4091_ (.Y(_1151_),
    .A(\g.g_y[4].g_x[6].t.out_sc ),
    .B(net41));
 sg13g2_o21ai_1 _4092_ (.B1(_1151_),
    .Y(\g.g_y[4].g_x[7].t.w_si ),
    .A1(net42),
    .A2(_1150_));
 sg13g2_inv_1 _4093_ (.Y(_1152_),
    .A(_0902_));
 sg13g2_a21oi_1 _4094_ (.A1(_0896_),
    .A2(_1152_),
    .Y(_1153_),
    .B1(_0903_));
 sg13g2_or2_1 _4095_ (.X(_1154_),
    .B(_0324_),
    .A(_0914_));
 sg13g2_inv_1 _4096_ (.Y(_1155_),
    .A(_0325_));
 sg13g2_a21oi_1 _4097_ (.A1(_1155_),
    .A2(_0914_),
    .Y(_1156_),
    .B1(net38));
 sg13g2_a221oi_1 _4098_ (.B2(_1156_),
    .C1(_0890_),
    .B1(_1154_),
    .A1(_0894_),
    .Y(_1157_),
    .A2(_0893_));
 sg13g2_a21o_1 _4099_ (.A2(_1153_),
    .A1(net39),
    .B1(_1157_),
    .X(_1158_));
 sg13g2_nand2_1 _4100_ (.Y(_1159_),
    .A(\g.g_y[4].g_x[7].t.out_sc ),
    .B(net41));
 sg13g2_o21ai_1 _4101_ (.B1(_1159_),
    .Y(\g.g_y[5].g_x[0].t.w_si ),
    .A1(net42),
    .A2(_1158_));
 sg13g2_inv_1 _4102_ (.Y(_1160_),
    .A(_0637_));
 sg13g2_nor2_1 _4103_ (.A(_0955_),
    .B(_0950_),
    .Y(_1161_));
 sg13g2_o21ai_1 _4104_ (.B1(_1161_),
    .Y(_1162_),
    .A1(_0967_),
    .A2(_1004_));
 sg13g2_mux2_1 _4105_ (.A0(_0411_),
    .A1(_0407_),
    .S(_0408_),
    .X(_1163_));
 sg13g2_mux2_1 _4106_ (.A0(_0961_),
    .A1(_1163_),
    .S(_0968_),
    .X(_1164_));
 sg13g2_nor2_1 _4107_ (.A(_0959_),
    .B(_0950_),
    .Y(_1165_));
 sg13g2_nor2_1 _4108_ (.A(_0955_),
    .B(net37),
    .Y(_1166_));
 sg13g2_nor2_1 _4109_ (.A(_0959_),
    .B(net37),
    .Y(_1167_));
 sg13g2_and3_1 _4110_ (.X(_1168_),
    .A(_0954_),
    .B(_0956_),
    .C(_1167_));
 sg13g2_a221oi_1 _4111_ (.B2(\g.g_y[5].g_x[2].t.out_sc ),
    .C1(_1168_),
    .B1(_1166_),
    .A1(_1164_),
    .Y(_1169_),
    .A2(_1165_));
 sg13g2_nand3_1 _4112_ (.B(_1162_),
    .C(_1169_),
    .A(_0898_),
    .Y(_1170_));
 sg13g2_nor2b_1 _4113_ (.A(_0321_),
    .B_N(_0325_),
    .Y(_1171_));
 sg13g2_a21o_1 _4114_ (.A2(_0324_),
    .A1(_0321_),
    .B1(_1171_),
    .X(_1172_));
 sg13g2_and2_1 _4115_ (.A(net38),
    .B(net39),
    .X(_1173_));
 sg13g2_nor2_1 _4116_ (.A(net38),
    .B(_0891_),
    .Y(_1174_));
 sg13g2_a22oi_1 _4117_ (.Y(_1175_),
    .B1(_1174_),
    .B2(_0893_),
    .A2(_1173_),
    .A1(_1172_));
 sg13g2_nor2_1 _4118_ (.A(net39),
    .B(\g.g_y[5].g_x[0].t.out_sc ),
    .Y(_1176_));
 sg13g2_nor2_1 _4119_ (.A(_0897_),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_o21ai_1 _4120_ (.B1(_1177_),
    .Y(_1178_),
    .A1(_0907_),
    .A2(_1175_));
 sg13g2_a221oi_1 _4121_ (.B2(_1156_),
    .C1(_0891_),
    .B1(_1154_),
    .A1(net38),
    .Y(_1179_),
    .A2(_0893_));
 sg13g2_o21ai_1 _4122_ (.B1(_0897_),
    .Y(_1180_),
    .A1(net6),
    .A2(net39));
 sg13g2_or2_1 _4123_ (.X(_1181_),
    .B(_1180_),
    .A(_1179_));
 sg13g2_nand3b_1 _4124_ (.B(_1178_),
    .C(_1181_),
    .Y(_1182_),
    .A_N(_0898_));
 sg13g2_and3_1 _4125_ (.X(_1183_),
    .A(_1160_),
    .B(_1170_),
    .C(_1182_));
 sg13g2_buf_1 _4126_ (.A(\g.g_y[6].g_x[1].t.r_v ),
    .X(_1184_));
 sg13g2_inv_1 _4127_ (.Y(_1185_),
    .A(net34));
 sg13g2_buf_1 _4128_ (.A(\g.g_y[6].g_x[1].t.r_d ),
    .X(_1186_));
 sg13g2_inv_1 _4129_ (.Y(_1187_),
    .A(_1186_));
 sg13g2_buf_2 _4130_ (.A(\g.g_y[6].g_x[0].t.r_h ),
    .X(_1188_));
 sg13g2_inv_1 _4131_ (.Y(_1189_),
    .A(_1188_));
 sg13g2_mux2_1 _4132_ (.A0(\g.g_y[6].g_x[0].t.out_sc ),
    .A1(\g.g_y[6].g_x[0].t.r_gnl ),
    .S(_1867_),
    .X(_1190_));
 sg13g2_or2_1 _4133_ (.X(_1191_),
    .B(_1188_),
    .A(_1869_));
 sg13g2_o21ai_1 _4134_ (.B1(_1191_),
    .Y(_1192_),
    .A1(_1189_),
    .A2(_1190_));
 sg13g2_buf_1 _4135_ (.A(\g.g_y[6].g_x[2].t.r_h ),
    .X(_1193_));
 sg13g2_mux2_1 _4136_ (.A0(\g.g_y[6].g_x[2].t.out_sc ),
    .A1(\g.g_y[6].g_x[2].t.r_gnl ),
    .S(_1950_),
    .X(_1194_));
 sg13g2_nand2b_1 _4137_ (.Y(_1195_),
    .B(_1193_),
    .A_N(_1949_));
 sg13g2_o21ai_1 _4138_ (.B1(_1195_),
    .Y(_1196_),
    .A1(_1193_),
    .A2(_1194_));
 sg13g2_buf_1 _4139_ (.A(\g.g_y[6].g_x[1].t.r_h ),
    .X(_1197_));
 sg13g2_mux2_1 _4140_ (.A0(_1192_),
    .A1(_1196_),
    .S(net68),
    .X(_1198_));
 sg13g2_buf_1 _4141_ (.A(_1198_),
    .X(_1199_));
 sg13g2_inv_1 _4142_ (.Y(_1200_),
    .A(_1799_));
 sg13g2_mux2_1 _4143_ (.A0(_1795_),
    .A1(_1798_),
    .S(_1200_),
    .X(_1201_));
 sg13g2_nor2_1 _4144_ (.A(net25),
    .B(_1201_),
    .Y(_1202_));
 sg13g2_a21oi_1 _4145_ (.A1(net25),
    .A2(_1199_),
    .Y(_1203_),
    .B1(_1202_));
 sg13g2_nor3_1 _4146_ (.A(_0641_),
    .B(_1185_),
    .C(_1203_),
    .Y(_1204_));
 sg13g2_nand4_1 _4147_ (.B(_0622_),
    .C(_0633_),
    .A(_0643_),
    .Y(_1205_),
    .D(_0635_));
 sg13g2_o21ai_1 _4148_ (.B1(_0644_),
    .Y(_1206_),
    .A1(_0653_),
    .A2(_0657_));
 sg13g2_a21oi_1 _4149_ (.A1(_1205_),
    .A2(_1206_),
    .Y(_1207_),
    .B1(_0640_));
 sg13g2_mux2_1 _4150_ (.A0(_1196_),
    .A1(_1192_),
    .S(net68),
    .X(_1208_));
 sg13g2_buf_1 _4151_ (.A(_1208_),
    .X(_1209_));
 sg13g2_nand2b_1 _4152_ (.Y(_1210_),
    .B(_1799_),
    .A_N(_1795_));
 sg13g2_o21ai_1 _4153_ (.B1(_1210_),
    .Y(_1211_),
    .A1(_1799_),
    .A2(_1798_));
 sg13g2_or2_1 _4154_ (.X(_1212_),
    .B(_0640_),
    .A(_0636_));
 sg13g2_o21ai_1 _4155_ (.B1(_1212_),
    .Y(_1213_),
    .A1(_0641_),
    .A2(_0639_));
 sg13g2_mux2_1 _4156_ (.A0(_1211_),
    .A1(_1213_),
    .S(net34),
    .X(_1214_));
 sg13g2_or3_1 _4157_ (.A(net33),
    .B(_1209_),
    .C(_1214_),
    .X(_1215_));
 sg13g2_nor2_1 _4158_ (.A(net25),
    .B(\g.g_y[6].g_x[1].t.out_sc ),
    .Y(_1216_));
 sg13g2_nor2_1 _4159_ (.A(_0641_),
    .B(_1216_),
    .Y(_1217_));
 sg13g2_a21oi_1 _4160_ (.A1(_0643_),
    .A2(_0647_),
    .Y(_1218_),
    .B1(_0640_));
 sg13g2_a221oi_1 _4161_ (.B2(_1217_),
    .C1(_1218_),
    .B1(_1215_),
    .A1(_0640_),
    .Y(_1219_),
    .A2(net34));
 sg13g2_nor4_1 _4162_ (.A(_1160_),
    .B(_1204_),
    .C(_1207_),
    .D(_1219_),
    .Y(_1220_));
 sg13g2_or2_1 _4163_ (.X(\g.g_y[5].g_x[1].t.w_dh ),
    .B(_1220_),
    .A(_1183_));
 sg13g2_nand2_1 _4164_ (.Y(_1221_),
    .A(_0644_),
    .B(_0658_));
 sg13g2_nand3b_1 _4165_ (.B(_0643_),
    .C(_0646_),
    .Y(_1222_),
    .A_N(_0647_));
 sg13g2_nand3_1 _4166_ (.B(_1221_),
    .C(_1222_),
    .A(_0640_),
    .Y(_1223_));
 sg13g2_mux2_1 _4167_ (.A0(_0636_),
    .A1(_0639_),
    .S(_0640_),
    .X(_1224_));
 sg13g2_and2_1 _4168_ (.A(net34),
    .B(_1210_),
    .X(_1225_));
 sg13g2_nand2b_1 _4169_ (.Y(_1226_),
    .B(_1200_),
    .A_N(_1798_));
 sg13g2_a221oi_1 _4170_ (.B2(_1226_),
    .C1(net25),
    .B1(_1225_),
    .A1(_1185_),
    .Y(_1227_),
    .A2(_1224_));
 sg13g2_a21oi_1 _4171_ (.A1(net25),
    .A2(_1199_),
    .Y(_1228_),
    .B1(_1227_));
 sg13g2_nor2_1 _4172_ (.A(net34),
    .B(_1216_),
    .Y(_1229_));
 sg13g2_a22oi_1 _4173_ (.Y(_1230_),
    .B1(_1229_),
    .B2(_1215_),
    .A2(_1228_),
    .A1(net34));
 sg13g2_nand2_1 _4174_ (.Y(_1231_),
    .A(_0641_),
    .B(_1230_));
 sg13g2_nand3b_1 _4175_ (.B(_1162_),
    .C(_1169_),
    .Y(_1232_),
    .A_N(_0898_));
 sg13g2_nand3_1 _4176_ (.B(_1178_),
    .C(_1181_),
    .A(_0898_),
    .Y(_1233_));
 sg13g2_nand4_1 _4177_ (.B(_1231_),
    .C(_1232_),
    .A(_1223_),
    .Y(\g.g_y[5].g_x[1].t.w_na ),
    .D(_1233_));
 sg13g2_nand2_1 _4178_ (.Y(_1234_),
    .A(\g.g_y[5].g_x[0].t.out_sc ),
    .B(net36));
 sg13g2_nand4_1 _4179_ (.B(net45),
    .C(_1170_),
    .A(_0637_),
    .Y(_1235_),
    .D(_1182_));
 sg13g2_nand2_1 _4180_ (.Y(_1236_),
    .A(_1160_),
    .B(_1900_));
 sg13g2_or4_1 _4181_ (.A(_1204_),
    .B(_1207_),
    .C(_1219_),
    .D(_1236_),
    .X(_1237_));
 sg13g2_nand3_1 _4182_ (.B(_1235_),
    .C(_1237_),
    .A(_1234_),
    .Y(\g.g_y[5].g_x[1].t.w_si ));
 sg13g2_nand2_1 _4183_ (.Y(_1238_),
    .A(net37),
    .B(_0960_));
 sg13g2_o21ai_1 _4184_ (.B1(_1238_),
    .Y(_1239_),
    .A1(net37),
    .A2(_1164_));
 sg13g2_nand2_1 _4185_ (.Y(_1240_),
    .A(\g.g_y[5].g_x[1].t.out_sc ),
    .B(net41));
 sg13g2_o21ai_1 _4186_ (.B1(_1240_),
    .Y(\g.g_y[5].g_x[2].t.w_si ),
    .A1(net42),
    .A2(_1239_));
 sg13g2_buf_2 _4187_ (.A(\g.g_y[6].g_x[3].t.r_d ),
    .X(_1241_));
 sg13g2_inv_1 _4188_ (.Y(_1242_),
    .A(\g.g_y[6].g_x[3].t.out_sc ));
 sg13g2_nand2_1 _4189_ (.Y(_1243_),
    .A(_1241_),
    .B(_1242_));
 sg13g2_mux2_1 _4190_ (.A0(\g.g_y[6].g_x[4].t.out_sc ),
    .A1(\g.g_y[6].g_x[4].t.r_gnl ),
    .S(_2103_),
    .X(_1244_));
 sg13g2_buf_2 _4191_ (.A(\g.g_y[6].g_x[4].t.r_h ),
    .X(_1245_));
 sg13g2_inv_1 _4192_ (.Y(_1246_),
    .A(_1245_));
 sg13g2_nand2b_1 _4193_ (.Y(_1247_),
    .B(_1246_),
    .A_N(_1244_));
 sg13g2_inv_1 _4194_ (.Y(_1248_),
    .A(_2102_));
 sg13g2_buf_1 _4195_ (.A(\g.g_y[6].g_x[3].t.r_h ),
    .X(_1249_));
 sg13g2_a21oi_1 _4196_ (.A1(_1248_),
    .A2(_1245_),
    .Y(_1250_),
    .B1(_1249_));
 sg13g2_mux2_1 _4197_ (.A0(_1949_),
    .A1(_1194_),
    .S(_1193_),
    .X(_1251_));
 sg13g2_a22oi_1 _4198_ (.Y(_1252_),
    .B1(_1251_),
    .B2(_1249_),
    .A2(_1250_),
    .A1(_1247_));
 sg13g2_inv_1 _4199_ (.Y(_1253_),
    .A(_1997_));
 sg13g2_nand2b_1 _4200_ (.Y(_1254_),
    .B(_1253_),
    .A_N(_1996_));
 sg13g2_buf_1 _4201_ (.A(\g.g_y[6].g_x[3].t.r_v ),
    .X(_1255_));
 sg13g2_a21oi_1 _4202_ (.A1(_1970_),
    .A2(_1997_),
    .Y(_1256_),
    .B1(_1255_));
 sg13g2_mux2_1 _4203_ (.A0(_0702_),
    .A1(_0698_),
    .S(_0699_),
    .X(_1257_));
 sg13g2_a22oi_1 _4204_ (.Y(_1258_),
    .B1(_1257_),
    .B2(_1255_),
    .A2(_1256_),
    .A1(_1254_));
 sg13g2_or3_1 _4205_ (.A(_1241_),
    .B(_1252_),
    .C(_1258_),
    .X(_1259_));
 sg13g2_buf_1 _4206_ (.A(_1259_),
    .X(_1260_));
 sg13g2_inv_2 _4207_ (.Y(_1261_),
    .A(_1255_));
 sg13g2_nand2_1 _4208_ (.Y(_1262_),
    .A(_0699_),
    .B(_1261_));
 sg13g2_a21oi_1 _4209_ (.A1(_1243_),
    .A2(_1260_),
    .Y(_1263_),
    .B1(_1262_));
 sg13g2_nand2_1 _4210_ (.Y(_1264_),
    .A(_0700_),
    .B(_0704_));
 sg13g2_a21oi_1 _4211_ (.A1(_0709_),
    .A2(_0711_),
    .Y(_1265_),
    .B1(_1264_));
 sg13g2_mux2_1 _4212_ (.A0(_1958_),
    .A1(_1996_),
    .S(_1253_),
    .X(_1266_));
 sg13g2_mux2_1 _4213_ (.A0(_1266_),
    .A1(_1257_),
    .S(_1261_),
    .X(_1267_));
 sg13g2_mux2_1 _4214_ (.A0(_2102_),
    .A1(_1244_),
    .S(_1246_),
    .X(_1268_));
 sg13g2_inv_1 _4215_ (.Y(_1269_),
    .A(_1249_));
 sg13g2_mux2_1 _4216_ (.A0(_1268_),
    .A1(_1251_),
    .S(_1269_),
    .X(_1270_));
 sg13g2_inv_1 _4217_ (.Y(_1271_),
    .A(_1241_));
 sg13g2_mux2_1 _4218_ (.A0(_1267_),
    .A1(_1270_),
    .S(_1271_),
    .X(_1272_));
 sg13g2_buf_1 _4219_ (.A(_1272_),
    .X(_1273_));
 sg13g2_nand2_1 _4220_ (.Y(_1274_),
    .A(_0699_),
    .B(_1255_));
 sg13g2_nor2_1 _4221_ (.A(_0699_),
    .B(_0704_),
    .Y(_1275_));
 sg13g2_o21ai_1 _4222_ (.B1(_1275_),
    .Y(_1276_),
    .A1(_0715_),
    .A2(_0718_));
 sg13g2_o21ai_1 _4223_ (.B1(_1276_),
    .Y(_1277_),
    .A1(_1273_),
    .A2(_1274_));
 sg13g2_nor3_1 _4224_ (.A(_1263_),
    .B(_1265_),
    .C(_1277_),
    .Y(_1278_));
 sg13g2_inv_1 _4225_ (.Y(_1279_),
    .A(_0697_));
 sg13g2_nand2b_1 _4226_ (.Y(_1280_),
    .B(_1042_),
    .A_N(_0762_));
 sg13g2_o21ai_1 _4227_ (.B1(_1280_),
    .Y(_1281_),
    .A1(_1042_),
    .A2(_1041_));
 sg13g2_nor4_1 _4228_ (.A(_1038_),
    .B(_1061_),
    .C(_1281_),
    .D(_1056_),
    .Y(_1282_));
 sg13g2_mux2_1 _4229_ (.A0(_2102_),
    .A1(_2104_),
    .S(_1051_),
    .X(_1283_));
 sg13g2_mux2_1 _4230_ (.A0(_1050_),
    .A1(_1283_),
    .S(_1035_),
    .X(_1284_));
 sg13g2_nand2_1 _4231_ (.Y(_1285_),
    .A(_1038_),
    .B(_1037_));
 sg13g2_nor2_1 _4232_ (.A(_1037_),
    .B(\g.g_y[5].g_x[4].t.out_sc ),
    .Y(_1286_));
 sg13g2_nor2_1 _4233_ (.A(_1039_),
    .B(_1037_),
    .Y(_1287_));
 sg13g2_a22oi_1 _4234_ (.Y(_1288_),
    .B1(_1287_),
    .B2(_1281_),
    .A2(_1286_),
    .A1(_1039_));
 sg13g2_o21ai_1 _4235_ (.B1(_1288_),
    .Y(_1289_),
    .A1(_1284_),
    .A2(_1285_));
 sg13g2_o21ai_1 _4236_ (.B1(_0952_),
    .Y(_1290_),
    .A1(_1282_),
    .A2(_1289_));
 sg13g2_o21ai_1 _4237_ (.B1(_1165_),
    .Y(_1291_),
    .A1(_0967_),
    .A2(_1004_));
 sg13g2_nand2_1 _4238_ (.Y(_1292_),
    .A(_1161_),
    .B(_1164_));
 sg13g2_a22oi_1 _4239_ (.Y(_1293_),
    .B1(_1166_),
    .B2(_0958_),
    .A2(_1167_),
    .A1(\g.g_y[5].g_x[2].t.out_sc ));
 sg13g2_nand4_1 _4240_ (.B(_1291_),
    .C(_1292_),
    .A(_0953_),
    .Y(_1294_),
    .D(_1293_));
 sg13g2_and3_1 _4241_ (.X(_1295_),
    .A(_1279_),
    .B(_1290_),
    .C(_1294_));
 sg13g2_a21o_1 _4242_ (.A2(_1278_),
    .A1(_0697_),
    .B1(_1295_),
    .X(\g.g_y[5].g_x[3].t.w_dh ));
 sg13g2_nor2_1 _4243_ (.A(_0704_),
    .B(_0719_),
    .Y(_1296_));
 sg13g2_a21oi_1 _4244_ (.A1(_0709_),
    .A2(_0711_),
    .Y(_1297_),
    .B1(_0710_));
 sg13g2_o21ai_1 _4245_ (.B1(_0699_),
    .Y(_1298_),
    .A1(_1296_),
    .A2(_1297_));
 sg13g2_nor2_1 _4246_ (.A(_1261_),
    .B(_1273_),
    .Y(_1299_));
 sg13g2_a21oi_1 _4247_ (.A1(_1243_),
    .A2(_1260_),
    .Y(_1300_),
    .B1(_1255_));
 sg13g2_o21ai_1 _4248_ (.B1(_0700_),
    .Y(_1301_),
    .A1(_1299_),
    .A2(_1300_));
 sg13g2_nand4_1 _4249_ (.B(_1291_),
    .C(_1292_),
    .A(_0952_),
    .Y(_1302_),
    .D(_1293_));
 sg13g2_o21ai_1 _4250_ (.B1(_0953_),
    .Y(_1303_),
    .A1(_1282_),
    .A2(_1289_));
 sg13g2_nand4_1 _4251_ (.B(_1301_),
    .C(_1302_),
    .A(_1298_),
    .Y(\g.g_y[5].g_x[3].t.w_na ),
    .D(_1303_));
 sg13g2_nand2_1 _4252_ (.Y(_1304_),
    .A(\g.g_y[5].g_x[2].t.out_sc ),
    .B(net36));
 sg13g2_nand4_1 _4253_ (.B(net45),
    .C(_1290_),
    .A(_0697_),
    .Y(_1305_),
    .D(_1294_));
 sg13g2_nand2_1 _4254_ (.Y(_1306_),
    .A(_1279_),
    .B(_1900_));
 sg13g2_or4_1 _4255_ (.A(_1263_),
    .B(_1265_),
    .C(_1277_),
    .D(_1306_),
    .X(_1307_));
 sg13g2_nand3_1 _4256_ (.B(_1305_),
    .C(_1307_),
    .A(_1304_),
    .Y(\g.g_y[5].g_x[3].t.w_si ));
 sg13g2_a221oi_1 _4257_ (.B2(_1064_),
    .C1(_1061_),
    .B1(_1046_),
    .A1(_1038_),
    .Y(_1308_),
    .A2(_1044_));
 sg13g2_nor2_1 _4258_ (.A(_1037_),
    .B(_1284_),
    .Y(_1309_));
 sg13g2_nor3_1 _4259_ (.A(net82),
    .B(_1308_),
    .C(_1309_),
    .Y(_1310_));
 sg13g2_a21o_1 _4260_ (.A2(net59),
    .A1(\g.g_y[5].g_x[3].t.out_sc ),
    .B1(_1310_),
    .X(\g.g_y[5].g_x[4].t.w_si ));
 sg13g2_nand2_1 _4261_ (.Y(_1311_),
    .A(_1043_),
    .B(_1038_));
 sg13g2_or4_1 _4262_ (.A(_1061_),
    .B(_1049_),
    .C(_1056_),
    .D(_1311_),
    .X(_1312_));
 sg13g2_o21ai_1 _4263_ (.B1(net69),
    .Y(_1313_),
    .A1(net35),
    .A2(_1095_));
 sg13g2_nor2_1 _4264_ (.A(net35),
    .B(\g.g_y[5].g_x[6].t.out_sc ),
    .Y(_1314_));
 sg13g2_o21ai_1 _4265_ (.B1(_1042_),
    .Y(_1315_),
    .A1(net69),
    .A2(_1314_));
 sg13g2_inv_1 _4266_ (.Y(_1316_),
    .A(_1315_));
 sg13g2_o21ai_1 _4267_ (.B1(_1316_),
    .Y(_1317_),
    .A1(_1116_),
    .A2(_1313_));
 sg13g2_nor2_1 _4268_ (.A(_1043_),
    .B(net69),
    .Y(_1318_));
 sg13g2_nand4_1 _4269_ (.B(_1099_),
    .C(_1105_),
    .A(net35),
    .Y(_1319_),
    .D(_1318_));
 sg13g2_mux2_1 _4270_ (.A0(_0702_),
    .A1(_0951_),
    .S(_0952_),
    .X(_1320_));
 sg13g2_o21ai_1 _4271_ (.B1(_1039_),
    .Y(_1321_),
    .A1(_1037_),
    .A2(_1320_));
 sg13g2_nor2_1 _4272_ (.A(_1039_),
    .B(_1286_),
    .Y(_1322_));
 sg13g2_nor2_1 _4273_ (.A(_1042_),
    .B(_1322_),
    .Y(_1323_));
 sg13g2_o21ai_1 _4274_ (.B1(_1323_),
    .Y(_1324_),
    .A1(_1063_),
    .A2(_1321_));
 sg13g2_and4_1 _4275_ (.A(_1312_),
    .B(_1317_),
    .C(_1319_),
    .D(_1324_),
    .X(_1325_));
 sg13g2_mux2_1 _4276_ (.A0(_2093_),
    .A1(_2133_),
    .S(_2132_),
    .X(_1326_));
 sg13g2_buf_2 _4277_ (.A(_1326_),
    .X(_1327_));
 sg13g2_or2_1 _4278_ (.X(_1328_),
    .B(_0758_),
    .A(_0760_));
 sg13g2_buf_1 _4279_ (.A(_1328_),
    .X(_1329_));
 sg13g2_a21oi_1 _4280_ (.A1(_0763_),
    .A2(_0760_),
    .Y(_1330_),
    .B1(\g.g_y[6].g_x[5].t.r_v ));
 sg13g2_inv_1 _4281_ (.Y(_1331_),
    .A(\g.g_y[6].g_x[5].t.r_d ));
 sg13g2_a221oi_1 _4282_ (.B2(_1330_),
    .C1(_1331_),
    .B1(_1329_),
    .A1(\g.g_y[6].g_x[5].t.r_v ),
    .Y(_1332_),
    .A2(_1327_));
 sg13g2_buf_1 _4283_ (.A(_1332_),
    .X(_1333_));
 sg13g2_mux2_1 _4284_ (.A0(\g.g_y[6].g_x[6].t.out_sc ),
    .A1(\g.g_y[6].g_x[6].t.r_gnl ),
    .S(_2260_),
    .X(_1334_));
 sg13g2_buf_1 _4285_ (.A(_1334_),
    .X(_1335_));
 sg13g2_buf_1 _4286_ (.A(\g.g_y[6].g_x[6].t.r_h ),
    .X(_1336_));
 sg13g2_inv_1 _4287_ (.Y(_1337_),
    .A(net67));
 sg13g2_nand2b_1 _4288_ (.Y(_1338_),
    .B(_1337_),
    .A_N(_1335_));
 sg13g2_buf_2 _4289_ (.A(\g.g_y[6].g_x[5].t.r_h ),
    .X(_1339_));
 sg13g2_inv_1 _4290_ (.Y(_1340_),
    .A(_1339_));
 sg13g2_a21oi_1 _4291_ (.A1(_1113_),
    .A2(net67),
    .Y(_1341_),
    .B1(_1340_));
 sg13g2_mux2_1 _4292_ (.A0(_2102_),
    .A1(_1244_),
    .S(_1245_),
    .X(_1342_));
 sg13g2_buf_2 _4293_ (.A(_1342_),
    .X(_1343_));
 sg13g2_buf_1 _4294_ (.A(\g.g_y[6].g_x[5].t.r_d ),
    .X(_1344_));
 sg13g2_a221oi_1 _4295_ (.B2(_1340_),
    .C1(net32),
    .B1(_1343_),
    .A1(_1338_),
    .Y(_1345_),
    .A2(_1341_));
 sg13g2_buf_1 _4296_ (.A(\g.g_y[6].g_x[5].t.r_v ),
    .X(_1346_));
 sg13g2_o21ai_1 _4297_ (.B1(net31),
    .Y(_1347_),
    .A1(_1333_),
    .A2(_1345_));
 sg13g2_inv_1 _4298_ (.Y(_1348_),
    .A(net31));
 sg13g2_mux2_1 _4299_ (.A0(_2264_),
    .A1(_1335_),
    .S(_1337_),
    .X(_1349_));
 sg13g2_mux2_1 _4300_ (.A0(_1349_),
    .A1(_1343_),
    .S(_1339_),
    .X(_1350_));
 sg13g2_nand4_1 _4301_ (.B(_1331_),
    .C(_1327_),
    .A(_1348_),
    .Y(_1351_),
    .D(_1350_));
 sg13g2_nand2b_1 _4302_ (.Y(_1352_),
    .B(net32),
    .A_N(\g.g_y[6].g_x[5].t.out_sc ));
 sg13g2_nand2b_1 _4303_ (.Y(_1353_),
    .B(_1348_),
    .A_N(_1352_));
 sg13g2_nand3_1 _4304_ (.B(_1351_),
    .C(_1353_),
    .A(_1347_),
    .Y(_1354_));
 sg13g2_and2_1 _4305_ (.A(_0753_),
    .B(_0779_),
    .X(_1355_));
 sg13g2_a221oi_1 _4306_ (.B2(_1355_),
    .C1(_0759_),
    .B1(_0816_),
    .A1(_0754_),
    .Y(_1356_),
    .A2(_1136_));
 sg13g2_a21oi_1 _4307_ (.A1(_0759_),
    .A2(_1354_),
    .Y(_1357_),
    .B1(_1356_));
 sg13g2_mux2_1 _4308_ (.A0(_1325_),
    .A1(_1357_),
    .S(_0756_),
    .X(\g.g_y[5].g_x[5].t.w_dh ));
 sg13g2_or3_1 _4309_ (.A(_1061_),
    .B(_1049_),
    .C(_1056_),
    .X(_1358_));
 sg13g2_o21ai_1 _4310_ (.B1(_1042_),
    .Y(_1359_),
    .A1(_1063_),
    .A2(_1321_));
 sg13g2_a21oi_1 _4311_ (.A1(_1358_),
    .A2(_1322_),
    .Y(_1360_),
    .B1(_1359_));
 sg13g2_nor2_1 _4312_ (.A(_1116_),
    .B(_1313_),
    .Y(_1361_));
 sg13g2_and3_1 _4313_ (.X(_1362_),
    .A(net35),
    .B(_1099_),
    .C(_1105_));
 sg13g2_nor3_1 _4314_ (.A(net69),
    .B(_1314_),
    .C(_1362_),
    .Y(_1363_));
 sg13g2_nor3_1 _4315_ (.A(_1042_),
    .B(_1361_),
    .C(_1363_),
    .Y(_1364_));
 sg13g2_a221oi_1 _4316_ (.B2(_1355_),
    .C1(_0760_),
    .B1(_0816_),
    .A1(_0754_),
    .Y(_1365_),
    .A2(_1136_));
 sg13g2_and2_1 _4317_ (.A(_0760_),
    .B(_1354_),
    .X(_1366_));
 sg13g2_or4_1 _4318_ (.A(_1360_),
    .B(_1364_),
    .C(_1365_),
    .D(_1366_),
    .X(\g.g_y[5].g_x[5].t.w_na ));
 sg13g2_inv_1 _4319_ (.Y(_1367_),
    .A(\g.g_y[5].g_x[4].t.out_sc ));
 sg13g2_nor3_1 _4320_ (.A(_0760_),
    .B(net31),
    .C(_1352_),
    .Y(_1368_));
 sg13g2_a21oi_1 _4321_ (.A1(_1347_),
    .A2(_1351_),
    .Y(_1369_),
    .B1(_0760_));
 sg13g2_or4_1 _4322_ (.A(_0756_),
    .B(_1368_),
    .C(_1369_),
    .D(_1356_),
    .X(_1370_));
 sg13g2_a21oi_1 _4323_ (.A1(_0756_),
    .A2(_1325_),
    .Y(_1371_),
    .B1(net36));
 sg13g2_a22oi_1 _4324_ (.Y(\g.g_y[5].g_x[5].t.w_si ),
    .B1(_1370_),
    .B2(_1371_),
    .A2(net60),
    .A1(_1367_));
 sg13g2_a221oi_1 _4325_ (.B2(_1114_),
    .C1(net35),
    .B1(_1112_),
    .A1(_1104_),
    .Y(_1372_),
    .A2(_1101_));
 sg13g2_a221oi_1 _4326_ (.B2(_1110_),
    .C1(_1091_),
    .B1(_1109_),
    .A1(net69),
    .Y(_1373_),
    .A2(_1095_));
 sg13g2_nor3_1 _4327_ (.A(_1894_),
    .B(_1372_),
    .C(_1373_),
    .Y(_1374_));
 sg13g2_a21o_1 _4328_ (.A2(net59),
    .A1(\g.g_y[5].g_x[5].t.out_sc ),
    .B1(_1374_),
    .X(\g.g_y[5].g_x[6].t.w_si ));
 sg13g2_mux2_1 _4329_ (.A0(\g.g_y[5].g_x[7].t.r_ghl ),
    .A1(_1092_),
    .S(_1093_),
    .X(\g.g_y[5].g_x[7].t.out_r ));
 sg13g2_inv_1 _4330_ (.Y(_1375_),
    .A(_0841_));
 sg13g2_o21ai_1 _4331_ (.B1(_1097_),
    .Y(_1376_),
    .A1(net35),
    .A2(\g.g_y[5].g_x[6].t.out_sc ));
 sg13g2_nor2_1 _4332_ (.A(net35),
    .B(_1096_),
    .Y(_1377_));
 sg13g2_or3_1 _4333_ (.A(_1097_),
    .B(_1116_),
    .C(_1377_),
    .X(_1378_));
 sg13g2_o21ai_1 _4334_ (.B1(_1378_),
    .Y(_1379_),
    .A1(_1362_),
    .A2(_1376_));
 sg13g2_o21ai_1 _4335_ (.B1(_0896_),
    .Y(_1380_),
    .A1(net39),
    .A2(_1152_));
 sg13g2_nor2_1 _4336_ (.A(_0896_),
    .B(_1176_),
    .Y(_1381_));
 sg13g2_o21ai_1 _4337_ (.B1(_1381_),
    .Y(_1382_),
    .A1(_0902_),
    .A2(_1175_));
 sg13g2_o21ai_1 _4338_ (.B1(_1382_),
    .Y(_1383_),
    .A1(_1179_),
    .A2(_1380_));
 sg13g2_mux2_1 _4339_ (.A0(_1379_),
    .A1(_1383_),
    .S(_1093_),
    .X(_1384_));
 sg13g2_buf_2 _4340_ (.A(\g.g_y[6].g_x[7].t.r_d ),
    .X(_1385_));
 sg13g2_inv_1 _4341_ (.Y(_1386_),
    .A(_1385_));
 sg13g2_buf_2 _4342_ (.A(\g.g_y[6].g_x[7].t.r_h ),
    .X(_1387_));
 sg13g2_mux2_1 _4343_ (.A0(_1869_),
    .A1(_1190_),
    .S(_1189_),
    .X(_1388_));
 sg13g2_buf_1 _4344_ (.A(_1388_),
    .X(_1389_));
 sg13g2_or2_1 _4345_ (.X(_1390_),
    .B(_1335_),
    .A(_1337_));
 sg13g2_nor2_1 _4346_ (.A(_2264_),
    .B(net67),
    .Y(_1391_));
 sg13g2_nor2_1 _4347_ (.A(_1387_),
    .B(_1391_),
    .Y(_1392_));
 sg13g2_a22oi_1 _4348_ (.Y(_1393_),
    .B1(_1390_),
    .B2(_1392_),
    .A2(_1389_),
    .A1(_1387_));
 sg13g2_buf_1 _4349_ (.A(\g.g_y[6].g_x[7].t.r_v ),
    .X(_1394_));
 sg13g2_inv_1 _4350_ (.Y(_1395_),
    .A(net30));
 sg13g2_mux2_1 _4351_ (.A0(\g.g_y[5].g_x[7].t.r_ghl ),
    .A1(_0842_),
    .S(_0843_),
    .X(_1396_));
 sg13g2_buf_2 _4352_ (.A(_1396_),
    .X(_1397_));
 sg13g2_inv_1 _4353_ (.Y(_1398_),
    .A(_2185_));
 sg13g2_nand2b_1 _4354_ (.Y(_1399_),
    .B(_1398_),
    .A_N(_2184_));
 sg13g2_nand2b_1 _4355_ (.Y(_1400_),
    .B(_2185_),
    .A_N(\g.g_y[7].g_x[7].t.r_ghl ));
 sg13g2_and2_1 _4356_ (.A(net30),
    .B(_1400_),
    .X(_1401_));
 sg13g2_a221oi_1 _4357_ (.B2(_1401_),
    .C1(_1386_),
    .B1(_1399_),
    .A1(_1395_),
    .Y(_1402_),
    .A2(_1397_));
 sg13g2_a21o_1 _4358_ (.A2(_1393_),
    .A1(_1386_),
    .B1(_1402_),
    .X(_1403_));
 sg13g2_buf_1 _4359_ (.A(_1403_),
    .X(_1404_));
 sg13g2_and2_1 _4360_ (.A(_0843_),
    .B(_1394_),
    .X(_1405_));
 sg13g2_nor2_1 _4361_ (.A(_0843_),
    .B(_0845_),
    .Y(_1406_));
 sg13g2_nor2_1 _4362_ (.A(_0843_),
    .B(_0846_),
    .Y(_1407_));
 sg13g2_and4_1 _4363_ (.A(_0833_),
    .B(_0839_),
    .C(_0848_),
    .D(_1407_),
    .X(_1408_));
 sg13g2_a221oi_1 _4364_ (.B2(_1145_),
    .C1(_1408_),
    .B1(_1406_),
    .A1(_1404_),
    .Y(_1409_),
    .A2(_1405_));
 sg13g2_inv_1 _4365_ (.Y(_1410_),
    .A(_1387_));
 sg13g2_nor2_1 _4366_ (.A(_1410_),
    .B(_1391_),
    .Y(_1411_));
 sg13g2_a22oi_1 _4367_ (.Y(_1412_),
    .B1(_1390_),
    .B2(_1411_),
    .A2(_1389_),
    .A1(_1410_));
 sg13g2_buf_1 _4368_ (.A(_1412_),
    .X(_1413_));
 sg13g2_and2_1 _4369_ (.A(_1395_),
    .B(_1400_),
    .X(_1414_));
 sg13g2_a22oi_1 _4370_ (.Y(_1415_),
    .B1(_1399_),
    .B2(_1414_),
    .A2(_1397_),
    .A1(net30));
 sg13g2_buf_1 _4371_ (.A(_1415_),
    .X(_1416_));
 sg13g2_nor2b_1 _4372_ (.A(_1394_),
    .B_N(_0843_),
    .Y(_1417_));
 sg13g2_nand2_1 _4373_ (.Y(_1418_),
    .A(_1386_),
    .B(_1417_));
 sg13g2_nor3_1 _4374_ (.A(_1413_),
    .B(_1416_),
    .C(_1418_),
    .Y(_1419_));
 sg13g2_nor2_1 _4375_ (.A(_1386_),
    .B(\g.g_y[6].g_x[7].t.out_sc ),
    .Y(_1420_));
 sg13g2_a22oi_1 _4376_ (.Y(_1421_),
    .B1(_1417_),
    .B2(_1420_),
    .A2(_1407_),
    .A1(_0850_));
 sg13g2_inv_1 _4377_ (.Y(_1422_),
    .A(_1421_));
 sg13g2_nor3_1 _4378_ (.A(_1375_),
    .B(_1419_),
    .C(_1422_),
    .Y(_1423_));
 sg13g2_and2_1 _4379_ (.A(_1409_),
    .B(_1423_),
    .X(_1424_));
 sg13g2_a21o_1 _4380_ (.A2(_1384_),
    .A1(_1375_),
    .B1(_1424_),
    .X(\g.g_y[5].g_x[7].t.w_dh ));
 sg13g2_nor2_1 _4381_ (.A(_1395_),
    .B(_1404_),
    .Y(_1425_));
 sg13g2_nor3_1 _4382_ (.A(_1385_),
    .B(_1413_),
    .C(_1416_),
    .Y(_1426_));
 sg13g2_nor3_1 _4383_ (.A(net30),
    .B(_1420_),
    .C(_1426_),
    .Y(_1427_));
 sg13g2_or3_1 _4384_ (.A(_0843_),
    .B(_1425_),
    .C(_1427_),
    .X(_1428_));
 sg13g2_nor2_1 _4385_ (.A(_0846_),
    .B(_0850_),
    .Y(_1429_));
 sg13g2_a22oi_1 _4386_ (.Y(_1430_),
    .B1(_1429_),
    .B2(_0849_),
    .A2(_0861_),
    .A1(_0846_));
 sg13g2_nand2_1 _4387_ (.Y(_1431_),
    .A(_0843_),
    .B(_1430_));
 sg13g2_mux2_1 _4388_ (.A0(_1383_),
    .A1(_1379_),
    .S(_1093_),
    .X(_1432_));
 sg13g2_nand3_1 _4389_ (.B(_1431_),
    .C(_1432_),
    .A(_1428_),
    .Y(\g.g_y[5].g_x[7].t.w_na ));
 sg13g2_and2_1 _4390_ (.A(_0841_),
    .B(_1093_),
    .X(_1433_));
 sg13g2_nor2_1 _4391_ (.A(_1375_),
    .B(_1093_),
    .Y(_1434_));
 sg13g2_a22oi_1 _4392_ (.Y(_1435_),
    .B1(_1434_),
    .B2(_1379_),
    .A2(_1433_),
    .A1(_1383_));
 sg13g2_nor4_1 _4393_ (.A(_0841_),
    .B(_2037_),
    .C(_1419_),
    .D(_1422_),
    .Y(_1436_));
 sg13g2_a22oi_1 _4394_ (.Y(_1437_),
    .B1(_1409_),
    .B2(_1436_),
    .A2(_2038_),
    .A1(\g.g_y[5].g_x[6].t.out_sc ));
 sg13g2_o21ai_1 _4395_ (.B1(_1437_),
    .Y(\g.g_y[5].g_x[7].t.w_si ),
    .A1(_0585_),
    .A2(_1435_));
 sg13g2_nand2b_1 _4396_ (.Y(_1438_),
    .B(_1820_),
    .A_N(_1788_));
 sg13g2_o21ai_1 _4397_ (.B1(_1438_),
    .Y(_1439_),
    .A1(_1820_),
    .A2(_0041_));
 sg13g2_buf_1 _4398_ (.A(_1439_),
    .X(_1440_));
 sg13g2_nand2_1 _4399_ (.Y(_1441_),
    .A(_1862_),
    .B(_1440_));
 sg13g2_nand3_1 _4400_ (.B(_1865_),
    .C(_1441_),
    .A(_1853_),
    .Y(_1442_));
 sg13g2_and2_1 _4401_ (.A(_1854_),
    .B(_1881_),
    .X(_1443_));
 sg13g2_o21ai_1 _4402_ (.B1(_1443_),
    .Y(_1444_),
    .A1(_1880_),
    .A2(_1440_));
 sg13g2_nand3_1 _4403_ (.B(_1442_),
    .C(_1444_),
    .A(\g.g_y[6].g_x[0].t.r_v ),
    .Y(_1445_));
 sg13g2_a21oi_1 _4404_ (.A1(_0321_),
    .A2(_0324_),
    .Y(_1446_),
    .B1(_1171_));
 sg13g2_a21oi_1 _4405_ (.A1(_0890_),
    .A2(_1446_),
    .Y(_1447_),
    .B1(net38));
 sg13g2_nand2_1 _4406_ (.Y(_1448_),
    .A(_0905_),
    .B(_1447_));
 sg13g2_nand2_1 _4407_ (.Y(_1449_),
    .A(_0891_),
    .B(_1172_));
 sg13g2_and2_1 _4408_ (.A(net38),
    .B(_0910_),
    .X(_1450_));
 sg13g2_o21ai_1 _4409_ (.B1(_1450_),
    .Y(_1451_),
    .A1(_0908_),
    .A2(_1449_));
 sg13g2_nand3_1 _4410_ (.B(_1448_),
    .C(_1451_),
    .A(_1866_),
    .Y(_1452_));
 sg13g2_and3_1 _4411_ (.X(_1453_),
    .A(_1867_),
    .B(_1445_),
    .C(_1452_));
 sg13g2_or3_1 _4412_ (.A(net25),
    .B(_1209_),
    .C(_1214_),
    .X(_1454_));
 sg13g2_inv_1 _4413_ (.Y(_1455_),
    .A(\g.g_y[6].g_x[1].t.out_sc ));
 sg13g2_a21oi_1 _4414_ (.A1(_1187_),
    .A2(_1455_),
    .Y(_1456_),
    .B1(net68));
 sg13g2_a221oi_1 _4415_ (.B2(_1456_),
    .C1(_1189_),
    .B1(_1454_),
    .A1(net68),
    .Y(_1457_),
    .A2(_1228_));
 sg13g2_nor2_1 _4416_ (.A(_1188_),
    .B(net7),
    .Y(_1458_));
 sg13g2_nor3_1 _4417_ (.A(_1867_),
    .B(_1457_),
    .C(_1458_),
    .Y(_1459_));
 sg13g2_or2_1 _4418_ (.X(\g.g_y[6].g_x[0].t.w_dh ),
    .B(_1459_),
    .A(_1453_));
 sg13g2_nand3_1 _4419_ (.B(_1442_),
    .C(_1444_),
    .A(_1866_),
    .Y(_1460_));
 sg13g2_nand3_1 _4420_ (.B(_1448_),
    .C(_1451_),
    .A(\g.g_y[6].g_x[0].t.r_v ),
    .Y(_1461_));
 sg13g2_nand2b_1 _4421_ (.Y(_1462_),
    .B(_1188_),
    .A_N(net7));
 sg13g2_a22oi_1 _4422_ (.Y(_1463_),
    .B1(_1454_),
    .B2(_1456_),
    .A2(_1228_),
    .A1(_1197_));
 sg13g2_nand2_1 _4423_ (.Y(_1464_),
    .A(_1189_),
    .B(_1463_));
 sg13g2_nand4_1 _4424_ (.B(_1461_),
    .C(_1462_),
    .A(_1460_),
    .Y(\g.g_y[6].g_x[0].t.w_na ),
    .D(_1464_));
 sg13g2_nand2_1 _4425_ (.Y(_1465_),
    .A(\g.g_y[5].g_x[7].t.out_sc ),
    .B(net36));
 sg13g2_nor2_1 _4426_ (.A(net74),
    .B(_1458_),
    .Y(_1466_));
 sg13g2_nand3b_1 _4427_ (.B(_1466_),
    .C(_1867_),
    .Y(_1467_),
    .A_N(_1457_));
 sg13g2_nor2_1 _4428_ (.A(_1867_),
    .B(_0111_),
    .Y(_1468_));
 sg13g2_nand3_1 _4429_ (.B(_1452_),
    .C(_1468_),
    .A(_1445_),
    .Y(_1469_));
 sg13g2_nand3_1 _4430_ (.B(_1467_),
    .C(_1469_),
    .A(_1465_),
    .Y(\g.g_y[6].g_x[0].t.w_si ));
 sg13g2_mux2_1 _4431_ (.A0(_1201_),
    .A1(_1224_),
    .S(_1185_),
    .X(_1470_));
 sg13g2_nand2_1 _4432_ (.Y(_1471_),
    .A(net33),
    .B(_1199_));
 sg13g2_o21ai_1 _4433_ (.B1(_1471_),
    .Y(_1472_),
    .A1(net33),
    .A2(_1470_));
 sg13g2_nand2_1 _4434_ (.Y(_1473_),
    .A(\g.g_y[6].g_x[0].t.out_sc ),
    .B(net41));
 sg13g2_o21ai_1 _4435_ (.B1(_1473_),
    .Y(\g.g_y[6].g_x[1].t.w_si ),
    .A1(_0585_),
    .A2(_1472_));
 sg13g2_inv_1 _4436_ (.Y(_1474_),
    .A(_1950_));
 sg13g2_nor2_1 _4437_ (.A(_1249_),
    .B(_1271_),
    .Y(_1475_));
 sg13g2_o21ai_1 _4438_ (.B1(_1475_),
    .Y(_1476_),
    .A1(_1252_),
    .A2(_1258_));
 sg13g2_nor2_1 _4439_ (.A(_1269_),
    .B(_1271_),
    .Y(_1477_));
 sg13g2_nor2_1 _4440_ (.A(_1269_),
    .B(_1241_),
    .Y(_1478_));
 sg13g2_nor3_1 _4441_ (.A(_1249_),
    .B(_1241_),
    .C(_1242_),
    .Y(_1479_));
 sg13g2_a221oi_1 _4442_ (.B2(_1268_),
    .C1(_1479_),
    .B1(_1478_),
    .A1(_1267_),
    .Y(_1480_),
    .A2(_1477_));
 sg13g2_nand3_1 _4443_ (.B(_1476_),
    .C(_1480_),
    .A(_1193_),
    .Y(_1481_));
 sg13g2_inv_1 _4444_ (.Y(_1482_),
    .A(_1193_));
 sg13g2_and2_1 _4445_ (.A(net68),
    .B(net33),
    .X(_1483_));
 sg13g2_o21ai_1 _4446_ (.B1(_1483_),
    .Y(_1484_),
    .A1(_1209_),
    .A2(_1214_));
 sg13g2_nor2_1 _4447_ (.A(net68),
    .B(net25),
    .Y(_1485_));
 sg13g2_nor2b_1 _4448_ (.A(net33),
    .B_N(net68),
    .Y(_1486_));
 sg13g2_nor3_1 _4449_ (.A(net68),
    .B(net33),
    .C(_1192_),
    .Y(_1487_));
 sg13g2_a221oi_1 _4450_ (.B2(\g.g_y[6].g_x[1].t.out_sc ),
    .C1(_1487_),
    .B1(_1486_),
    .A1(_1470_),
    .Y(_1488_),
    .A2(_1485_));
 sg13g2_nand3_1 _4451_ (.B(_1484_),
    .C(_1488_),
    .A(_1482_),
    .Y(_1489_));
 sg13g2_and2_1 _4452_ (.A(_1481_),
    .B(_1489_),
    .X(_1490_));
 sg13g2_o21ai_1 _4453_ (.B1(_1975_),
    .Y(_1491_),
    .A1(_1929_),
    .A2(_1928_));
 sg13g2_nor4_1 _4454_ (.A(_1947_),
    .B(_1966_),
    .C(_1491_),
    .D(_1973_),
    .Y(_1492_));
 sg13g2_nand2_1 _4455_ (.Y(_1493_),
    .A(_1947_),
    .B(_1967_));
 sg13g2_nor2_1 _4456_ (.A(_1948_),
    .B(_1967_),
    .Y(_1494_));
 sg13g2_nor2_1 _4457_ (.A(_1947_),
    .B(_1979_),
    .Y(_1495_));
 sg13g2_a21oi_1 _4458_ (.A1(_1491_),
    .A2(_1494_),
    .Y(_1496_),
    .B1(_1495_));
 sg13g2_o21ai_1 _4459_ (.B1(_1496_),
    .Y(_1497_),
    .A1(_1965_),
    .A2(_1493_));
 sg13g2_o21ai_1 _4460_ (.B1(_1952_),
    .Y(_1498_),
    .A1(_1492_),
    .A2(_1497_));
 sg13g2_or4_1 _4461_ (.A(_0968_),
    .B(net37),
    .C(_0967_),
    .D(_1003_),
    .X(_1499_));
 sg13g2_nor2_1 _4462_ (.A(_0962_),
    .B(_0949_),
    .Y(_1500_));
 sg13g2_nor2_1 _4463_ (.A(_0962_),
    .B(_0950_),
    .Y(_1501_));
 sg13g2_nor2_1 _4464_ (.A(_0968_),
    .B(_0971_),
    .Y(_1502_));
 sg13g2_a221oi_1 _4465_ (.B2(_1003_),
    .C1(_1502_),
    .B1(_1501_),
    .A1(_0960_),
    .Y(_1503_),
    .A2(_1500_));
 sg13g2_a21o_1 _4466_ (.A2(_1503_),
    .A1(_1499_),
    .B1(_1952_),
    .X(_1504_));
 sg13g2_and3_1 _4467_ (.X(_1505_),
    .A(_1950_),
    .B(_1498_),
    .C(_1504_));
 sg13g2_a21o_1 _4468_ (.A2(_1490_),
    .A1(_1474_),
    .B1(_1505_),
    .X(\g.g_y[6].g_x[2].t.w_dh ));
 sg13g2_a21oi_1 _4469_ (.A1(_1484_),
    .A2(_1488_),
    .Y(_1506_),
    .B1(_1482_));
 sg13g2_a21oi_1 _4470_ (.A1(_1476_),
    .A2(_1480_),
    .Y(_1507_),
    .B1(_1193_));
 sg13g2_nor2_1 _4471_ (.A(_1492_),
    .B(_1497_),
    .Y(_1508_));
 sg13g2_and2_1 _4472_ (.A(_1499_),
    .B(_1503_),
    .X(_1509_));
 sg13g2_mux2_1 _4473_ (.A0(_1508_),
    .A1(_1509_),
    .S(_1952_),
    .X(_1510_));
 sg13g2_o21ai_1 _4474_ (.B1(_1510_),
    .Y(\g.g_y[6].g_x[2].t.w_na ),
    .A1(_1506_),
    .A2(_1507_));
 sg13g2_nand2_1 _4475_ (.Y(_1511_),
    .A(\g.g_y[6].g_x[1].t.out_sc ),
    .B(net36));
 sg13g2_nand4_1 _4476_ (.B(net45),
    .C(_1481_),
    .A(_1950_),
    .Y(_1512_),
    .D(_1489_));
 sg13g2_nand4_1 _4477_ (.B(net73),
    .C(_1498_),
    .A(_1474_),
    .Y(_1513_),
    .D(_1504_));
 sg13g2_nand3_1 _4478_ (.B(_1512_),
    .C(_1513_),
    .A(_1511_),
    .Y(\g.g_y[6].g_x[2].t.w_si ));
 sg13g2_mux2_1 _4479_ (.A0(_1267_),
    .A1(_1270_),
    .S(_1241_),
    .X(_1514_));
 sg13g2_mux2_1 _4480_ (.A0(\g.g_y[6].g_x[2].t.out_sc ),
    .A1(_1514_),
    .S(net64),
    .X(\g.g_y[6].g_x[3].t.w_si ));
 sg13g2_inv_1 _4481_ (.Y(_1515_),
    .A(_2103_));
 sg13g2_nor2_1 _4482_ (.A(_1063_),
    .B(_1065_),
    .Y(_1516_));
 sg13g2_nand2_1 _4483_ (.Y(_1517_),
    .A(_1051_),
    .B(_1036_));
 sg13g2_nor2_1 _4484_ (.A(_1051_),
    .B(_2100_),
    .Y(_1518_));
 sg13g2_nor2_1 _4485_ (.A(_2105_),
    .B(_1036_),
    .Y(_1519_));
 sg13g2_a22oi_1 _4486_ (.Y(_1520_),
    .B1(_1519_),
    .B2(_1069_),
    .A2(_1518_),
    .A1(_2113_));
 sg13g2_o21ai_1 _4487_ (.B1(_1520_),
    .Y(_1521_),
    .A1(_1516_),
    .A2(_1517_));
 sg13g2_nand2_1 _4488_ (.Y(_1522_),
    .A(_2105_),
    .B(_2111_));
 sg13g2_nor4_1 _4489_ (.A(net55),
    .B(_2098_),
    .C(_2108_),
    .D(_1522_),
    .Y(_1523_));
 sg13g2_a21o_1 _4490_ (.A2(_1519_),
    .A1(_1057_),
    .B1(_1523_),
    .X(_1524_));
 sg13g2_nor3_1 _4491_ (.A(_1051_),
    .B(_2111_),
    .C(_2121_),
    .Y(_1525_));
 sg13g2_nor4_1 _4492_ (.A(_1515_),
    .B(_1521_),
    .C(_1524_),
    .D(_1525_),
    .Y(_1526_));
 sg13g2_or3_1 _4493_ (.A(_1271_),
    .B(_1252_),
    .C(_1258_),
    .X(_1527_));
 sg13g2_a21oi_1 _4494_ (.A1(_1271_),
    .A2(_1242_),
    .Y(_1528_),
    .B1(_1269_));
 sg13g2_a21oi_1 _4495_ (.A1(_1970_),
    .A2(_1997_),
    .Y(_1529_),
    .B1(_1261_));
 sg13g2_a221oi_1 _4496_ (.B2(_1254_),
    .C1(_1271_),
    .B1(_1529_),
    .A1(_1261_),
    .Y(_1530_),
    .A2(_1257_));
 sg13g2_o21ai_1 _4497_ (.B1(_1269_),
    .Y(_1531_),
    .A1(_1241_),
    .A2(_1251_));
 sg13g2_o21ai_1 _4498_ (.B1(_1246_),
    .Y(_1532_),
    .A1(_1530_),
    .A2(_1531_));
 sg13g2_a21o_1 _4499_ (.A2(_1528_),
    .A1(_1527_),
    .B1(_1532_),
    .X(_1533_));
 sg13g2_mux2_1 _4500_ (.A0(_0762_),
    .A1(_0758_),
    .S(_0759_),
    .X(_1534_));
 sg13g2_mux2_1 _4501_ (.A0(_1327_),
    .A1(_1534_),
    .S(net31),
    .X(_1535_));
 sg13g2_nand3_1 _4502_ (.B(_1350_),
    .C(_1535_),
    .A(net32),
    .Y(_1536_));
 sg13g2_nor2_1 _4503_ (.A(net32),
    .B(\g.g_y[6].g_x[5].t.out_sc ),
    .Y(_1537_));
 sg13g2_nor2_1 _4504_ (.A(_1339_),
    .B(_1537_),
    .Y(_1538_));
 sg13g2_o21ai_1 _4505_ (.B1(_1339_),
    .Y(_1539_),
    .A1(_1344_),
    .A2(_1349_));
 sg13g2_o21ai_1 _4506_ (.B1(_1245_),
    .Y(_1540_),
    .A1(_1333_),
    .A2(_1539_));
 sg13g2_a21o_1 _4507_ (.A2(_1538_),
    .A1(_1536_),
    .B1(_1540_),
    .X(_1541_));
 sg13g2_and3_1 _4508_ (.X(_1542_),
    .A(_1515_),
    .B(_1533_),
    .C(_1541_));
 sg13g2_or2_1 _4509_ (.X(\g.g_y[6].g_x[4].t.w_dh ),
    .B(_1542_),
    .A(_1526_));
 sg13g2_nor2_1 _4510_ (.A(_1530_),
    .B(_1531_),
    .Y(_1543_));
 sg13g2_a21oi_1 _4511_ (.A1(_1527_),
    .A2(_1528_),
    .Y(_1544_),
    .B1(_1543_));
 sg13g2_nor2_1 _4512_ (.A(_1333_),
    .B(_1539_),
    .Y(_1545_));
 sg13g2_a21oi_1 _4513_ (.A1(_1536_),
    .A2(_1538_),
    .Y(_1546_),
    .B1(_1545_));
 sg13g2_mux2_1 _4514_ (.A0(_1544_),
    .A1(_1546_),
    .S(_1246_),
    .X(_1547_));
 sg13g2_nor2_1 _4515_ (.A(_1035_),
    .B(_1067_),
    .Y(_1548_));
 sg13g2_nor3_1 _4516_ (.A(_1036_),
    .B(_1069_),
    .C(_1057_),
    .Y(_1549_));
 sg13g2_nor3_1 _4517_ (.A(_1051_),
    .B(_1548_),
    .C(_1549_),
    .Y(_1550_));
 sg13g2_nor2_1 _4518_ (.A(_2100_),
    .B(_2113_),
    .Y(_1551_));
 sg13g2_a221oi_1 _4519_ (.B2(_2110_),
    .C1(_2105_),
    .B1(_1551_),
    .A1(_2100_),
    .Y(_1552_),
    .A2(_2121_));
 sg13g2_or3_1 _4520_ (.A(_1547_),
    .B(_1550_),
    .C(_1552_),
    .X(\g.g_y[6].g_x[4].t.w_na ));
 sg13g2_nand2_1 _4521_ (.Y(_1553_),
    .A(\g.g_y[6].g_x[3].t.out_sc ),
    .B(net36));
 sg13g2_nand2_1 _4522_ (.Y(_1554_),
    .A(_1515_),
    .B(net81));
 sg13g2_or4_1 _4523_ (.A(_1521_),
    .B(_1524_),
    .C(_1525_),
    .D(_1554_),
    .X(_1555_));
 sg13g2_nand4_1 _4524_ (.B(net73),
    .C(_1533_),
    .A(_2103_),
    .Y(_1556_),
    .D(_1541_));
 sg13g2_nand3_1 _4525_ (.B(_1555_),
    .C(_1556_),
    .A(_1553_),
    .Y(\g.g_y[6].g_x[4].t.w_si ));
 sg13g2_a221oi_1 _4526_ (.B2(_1330_),
    .C1(net32),
    .B1(_1329_),
    .A1(net31),
    .Y(_1557_),
    .A2(_1327_));
 sg13g2_a221oi_1 _4527_ (.B2(_1340_),
    .C1(_1331_),
    .B1(_1343_),
    .A1(_1338_),
    .Y(_1558_),
    .A2(_1341_));
 sg13g2_nor3_1 _4528_ (.A(net82),
    .B(_1557_),
    .C(_1558_),
    .Y(_1559_));
 sg13g2_a21o_1 _4529_ (.A2(net59),
    .A1(\g.g_y[6].g_x[4].t.out_sc ),
    .B1(_1559_),
    .X(\g.g_y[6].g_x[5].t.w_si ));
 sg13g2_o21ai_1 _4530_ (.B1(_1104_),
    .Y(_1560_),
    .A1(_1111_),
    .A2(_1116_));
 sg13g2_and3_1 _4531_ (.X(_1561_),
    .A(_1103_),
    .B(_1091_),
    .C(_1101_));
 sg13g2_a21oi_1 _4532_ (.A1(_1099_),
    .A2(_1561_),
    .Y(_1562_),
    .B1(net49));
 sg13g2_or4_1 _4533_ (.A(net50),
    .B(net48),
    .C(_0012_),
    .D(_0015_),
    .X(_1563_));
 sg13g2_a22oi_1 _4534_ (.Y(_1564_),
    .B1(_1563_),
    .B2(net49),
    .A2(_1562_),
    .A1(_1560_));
 sg13g2_nor2_1 _4535_ (.A(_2269_),
    .B(_0000_),
    .Y(_1565_));
 sg13g2_o21ai_1 _4536_ (.B1(net49),
    .Y(_1566_),
    .A1(net50),
    .A2(_0006_));
 sg13g2_a21oi_1 _4537_ (.A1(net50),
    .A2(_1565_),
    .Y(_1567_),
    .B1(_1566_));
 sg13g2_nor3_1 _4538_ (.A(net49),
    .B(_1104_),
    .C(_1107_),
    .Y(_1568_));
 sg13g2_nor3_1 _4539_ (.A(_1564_),
    .B(_1567_),
    .C(_1568_),
    .Y(_1569_));
 sg13g2_nand4_1 _4540_ (.B(net32),
    .C(_1343_),
    .A(_1339_),
    .Y(_1570_),
    .D(_1535_));
 sg13g2_nor3_1 _4541_ (.A(_1339_),
    .B(_1344_),
    .C(_1343_),
    .Y(_1571_));
 sg13g2_nand2_1 _4542_ (.Y(_1572_),
    .A(_1340_),
    .B(net32));
 sg13g2_a221oi_1 _4543_ (.B2(_1330_),
    .C1(_1572_),
    .B1(_1329_),
    .A1(net31),
    .Y(_1573_),
    .A2(_1327_));
 sg13g2_nor3_1 _4544_ (.A(net67),
    .B(_1571_),
    .C(_1573_),
    .Y(_1574_));
 sg13g2_nor2_1 _4545_ (.A(_1385_),
    .B(_1389_),
    .Y(_1575_));
 sg13g2_o21ai_1 _4546_ (.B1(_1387_),
    .Y(_1576_),
    .A1(_1402_),
    .A2(_1575_));
 sg13g2_a22oi_1 _4547_ (.Y(_1577_),
    .B1(_1576_),
    .B2(net67),
    .A2(_1574_),
    .A1(_1570_));
 sg13g2_nor2_1 _4548_ (.A(_1337_),
    .B(_1387_),
    .Y(_1578_));
 sg13g2_nand2_1 _4549_ (.Y(_1579_),
    .A(_1385_),
    .B(_1578_));
 sg13g2_nor3_1 _4550_ (.A(_1413_),
    .B(_1416_),
    .C(_1579_),
    .Y(_1580_));
 sg13g2_nor2_1 _4551_ (.A(net67),
    .B(_1340_),
    .Y(_1581_));
 sg13g2_nor2_1 _4552_ (.A(_1385_),
    .B(\g.g_y[6].g_x[7].t.out_sc ),
    .Y(_1582_));
 sg13g2_a22oi_1 _4553_ (.Y(_1583_),
    .B1(_1578_),
    .B2(_1582_),
    .A2(_1581_),
    .A1(_1537_));
 sg13g2_nand2b_1 _4554_ (.Y(_1584_),
    .B(_1583_),
    .A_N(_1580_));
 sg13g2_nor3_1 _4555_ (.A(_2260_),
    .B(_1577_),
    .C(_1584_),
    .Y(_1585_));
 sg13g2_a21o_1 _4556_ (.A2(_1569_),
    .A1(_2260_),
    .B1(_1585_),
    .X(\g.g_y[6].g_x[6].t.w_dh ));
 sg13g2_nand2_1 _4557_ (.Y(_1586_),
    .A(net50),
    .B(_1565_));
 sg13g2_or3_1 _4558_ (.A(net50),
    .B(_0006_),
    .C(_0016_),
    .X(_1587_));
 sg13g2_nand3_1 _4559_ (.B(_1586_),
    .C(_1587_),
    .A(_2259_),
    .Y(_1588_));
 sg13g2_nand2_1 _4560_ (.Y(_1589_),
    .A(_1104_),
    .B(_1117_));
 sg13g2_nand3_1 _4561_ (.B(_1106_),
    .C(_1107_),
    .A(_1103_),
    .Y(_1590_));
 sg13g2_nand3_1 _4562_ (.B(_1589_),
    .C(_1590_),
    .A(net49),
    .Y(_1591_));
 sg13g2_or2_1 _4563_ (.X(_1592_),
    .B(_1573_),
    .A(_1571_));
 sg13g2_or2_1 _4564_ (.X(_1593_),
    .B(\g.g_y[6].g_x[5].t.out_sc ),
    .A(net32));
 sg13g2_a21oi_1 _4565_ (.A1(_1536_),
    .A2(_1593_),
    .Y(_1594_),
    .B1(_1340_));
 sg13g2_o21ai_1 _4566_ (.B1(net67),
    .Y(_1595_),
    .A1(_1592_),
    .A2(_1594_));
 sg13g2_nor3_1 _4567_ (.A(_1386_),
    .B(_1413_),
    .C(_1416_),
    .Y(_1596_));
 sg13g2_nor2_1 _4568_ (.A(_1582_),
    .B(_1596_),
    .Y(_1597_));
 sg13g2_o21ai_1 _4569_ (.B1(_1337_),
    .Y(_1598_),
    .A1(_1410_),
    .A2(_1404_));
 sg13g2_a21o_1 _4570_ (.A2(_1597_),
    .A1(_1410_),
    .B1(_1598_),
    .X(_1599_));
 sg13g2_nand4_1 _4571_ (.B(_1591_),
    .C(_1595_),
    .A(_1588_),
    .Y(\g.g_y[6].g_x[6].t.w_na ),
    .D(_1599_));
 sg13g2_nand2_1 _4572_ (.Y(_1600_),
    .A(\g.g_y[6].g_x[5].t.out_sc ),
    .B(_1009_));
 sg13g2_or2_1 _4573_ (.X(_1601_),
    .B(_1568_),
    .A(_2260_));
 sg13g2_or4_1 _4574_ (.A(_2037_),
    .B(_1564_),
    .C(_1567_),
    .D(_1601_),
    .X(_1602_));
 sg13g2_nand2_1 _4575_ (.Y(_1603_),
    .A(_2260_),
    .B(net81));
 sg13g2_or3_1 _4576_ (.A(_1577_),
    .B(_1584_),
    .C(_1603_),
    .X(_1604_));
 sg13g2_nand3_1 _4577_ (.B(_1602_),
    .C(_1604_),
    .A(_1600_),
    .Y(\g.g_y[6].g_x[6].t.w_si ));
 sg13g2_nand2_1 _4578_ (.Y(_1605_),
    .A(_1387_),
    .B(_1597_));
 sg13g2_o21ai_1 _4579_ (.B1(_1605_),
    .Y(\g.g_y[6].g_x[7].t.out_r ),
    .A1(_1387_),
    .A2(_1404_));
 sg13g2_a221oi_1 _4580_ (.B2(_1401_),
    .C1(_1385_),
    .B1(_1399_),
    .A1(_1395_),
    .Y(_1606_),
    .A2(_1397_));
 sg13g2_a21o_1 _4581_ (.A2(_1393_),
    .A1(_1385_),
    .B1(_1606_),
    .X(_1607_));
 sg13g2_nand2_1 _4582_ (.Y(_1608_),
    .A(\g.g_y[6].g_x[6].t.out_sc ),
    .B(_0751_));
 sg13g2_o21ai_1 _4583_ (.B1(_1608_),
    .Y(\g.g_y[6].g_x[7].t.w_si ),
    .A1(net59),
    .A2(_1607_));
 sg13g2_inv_1 _4584_ (.Y(_1609_),
    .A(_1861_));
 sg13g2_a21oi_1 _4585_ (.A1(_1855_),
    .A2(_1609_),
    .Y(_1610_),
    .B1(_1863_));
 sg13g2_mux2_1 _4586_ (.A0(_1872_),
    .A1(_1440_),
    .S(_1853_),
    .X(_1611_));
 sg13g2_mux2_1 _4587_ (.A0(_1610_),
    .A1(_1611_),
    .S(_1875_),
    .X(_1612_));
 sg13g2_nand2_1 _4588_ (.Y(_1613_),
    .A(\g.g_y[6].g_x[7].t.out_sc ),
    .B(_0751_));
 sg13g2_o21ai_1 _4589_ (.B1(_1613_),
    .Y(\g.g_y[7].g_x[0].t.w_si ),
    .A1(_2044_),
    .A2(_1612_));
 sg13g2_inv_1 _4590_ (.Y(_1614_),
    .A(_1796_));
 sg13g2_nor2_1 _4591_ (.A(_1964_),
    .B(_1967_),
    .Y(_1615_));
 sg13g2_o21ai_1 _4592_ (.B1(_1615_),
    .Y(_1616_),
    .A1(_1973_),
    .A2(_1977_));
 sg13g2_inv_1 _4593_ (.Y(_1617_),
    .A(_1964_));
 sg13g2_nor2_1 _4594_ (.A(_1617_),
    .B(_1967_),
    .Y(_1618_));
 sg13g2_nand2_1 _4595_ (.Y(_1619_),
    .A(_1956_),
    .B(_1618_));
 sg13g2_nor2_1 _4596_ (.A(_1617_),
    .B(_1966_),
    .Y(_1620_));
 sg13g2_nor2_1 _4597_ (.A(_1964_),
    .B(_1966_),
    .Y(_1621_));
 sg13g2_a22oi_1 _4598_ (.Y(_1622_),
    .B1(_1621_),
    .B2(\g.g_y[7].g_x[2].t.out_sc ),
    .A2(_1620_),
    .A1(_1963_));
 sg13g2_nand4_1 _4599_ (.B(_1616_),
    .C(_1619_),
    .A(_1857_),
    .Y(_1623_),
    .D(_1622_));
 sg13g2_mux2_1 _4600_ (.A0(_1872_),
    .A1(_1440_),
    .S(_1854_),
    .X(_1624_));
 sg13g2_nand2_1 _4601_ (.Y(_1625_),
    .A(net8),
    .B(net65));
 sg13g2_nor2_1 _4602_ (.A(\g.g_y[7].g_x[0].t.out_sc ),
    .B(net65),
    .Y(_1626_));
 sg13g2_nor2_1 _4603_ (.A(_1856_),
    .B(_1626_),
    .Y(_1627_));
 sg13g2_o21ai_1 _4604_ (.B1(_1627_),
    .Y(_1628_),
    .A1(_1624_),
    .A2(_1625_));
 sg13g2_o21ai_1 _4605_ (.B1(_1856_),
    .Y(_1629_),
    .A1(net8),
    .A2(net65));
 sg13g2_a21o_1 _4606_ (.A2(_1611_),
    .A1(net65),
    .B1(_1629_),
    .X(_1630_));
 sg13g2_nand3_1 _4607_ (.B(_1628_),
    .C(_1630_),
    .A(_1878_),
    .Y(_1631_));
 sg13g2_and3_1 _4608_ (.X(_1632_),
    .A(_1614_),
    .B(_1623_),
    .C(_1631_));
 sg13g2_and2_1 _4609_ (.A(_1807_),
    .B(_0072_),
    .X(_1633_));
 sg13g2_a221oi_1 _4610_ (.B2(_1633_),
    .C1(_1200_),
    .B1(_0071_),
    .A1(_1806_),
    .Y(_1634_),
    .A2(_1815_));
 sg13g2_or4_1 _4611_ (.A(_1185_),
    .B(net33),
    .C(_1209_),
    .D(_1213_),
    .X(_1635_));
 sg13g2_nor2_1 _4612_ (.A(net34),
    .B(net33),
    .Y(_1636_));
 sg13g2_nor3_1 _4613_ (.A(net34),
    .B(net25),
    .C(_1224_),
    .Y(_1637_));
 sg13g2_a221oi_1 _4614_ (.B2(_1199_),
    .C1(_1637_),
    .B1(_1636_),
    .A1(_1184_),
    .Y(_1638_),
    .A2(_1216_));
 sg13g2_a21oi_1 _4615_ (.A1(_1635_),
    .A2(_1638_),
    .Y(_1639_),
    .B1(_1799_));
 sg13g2_nor3_1 _4616_ (.A(_1614_),
    .B(_1634_),
    .C(_1639_),
    .Y(_1640_));
 sg13g2_or2_1 _4617_ (.X(\g.g_y[7].g_x[1].t.w_dh ),
    .B(_1640_),
    .A(_1632_));
 sg13g2_nand4_1 _4618_ (.B(_1616_),
    .C(_1619_),
    .A(_1878_),
    .Y(_1641_),
    .D(_1622_));
 sg13g2_nand3_1 _4619_ (.B(_1628_),
    .C(_1630_),
    .A(_1857_),
    .Y(_1642_));
 sg13g2_a22oi_1 _4620_ (.Y(_1643_),
    .B1(_0071_),
    .B2(_1633_),
    .A2(_1815_),
    .A1(_1806_));
 sg13g2_a21oi_1 _4621_ (.A1(_1635_),
    .A2(_1638_),
    .Y(_1644_),
    .B1(_1200_));
 sg13g2_a21oi_1 _4622_ (.A1(_1200_),
    .A2(_1643_),
    .Y(_1645_),
    .B1(_1644_));
 sg13g2_nand3_1 _4623_ (.B(_1642_),
    .C(_1645_),
    .A(_1641_),
    .Y(\g.g_y[7].g_x[1].t.w_na ));
 sg13g2_nand2_1 _4624_ (.Y(_1646_),
    .A(\g.g_y[7].g_x[0].t.out_sc ),
    .B(_1009_));
 sg13g2_nand4_1 _4625_ (.B(_0246_),
    .C(_1623_),
    .A(_1796_),
    .Y(_1647_),
    .D(_1631_));
 sg13g2_or4_1 _4626_ (.A(_1796_),
    .B(_0111_),
    .C(_1634_),
    .D(_1639_),
    .X(_1648_));
 sg13g2_nand3_1 _4627_ (.B(_1647_),
    .C(_1648_),
    .A(_1646_),
    .Y(\g.g_y[7].g_x[1].t.w_si ));
 sg13g2_mux2_1 _4628_ (.A0(_1956_),
    .A1(_1965_),
    .S(_1966_),
    .X(_1649_));
 sg13g2_mux2_1 _4629_ (.A0(\g.g_y[7].g_x[1].t.out_sc ),
    .A1(_1649_),
    .S(net64),
    .X(\g.g_y[7].g_x[2].t.w_si ));
 sg13g2_inv_1 _4630_ (.Y(_1650_),
    .A(_1959_));
 sg13g2_and2_1 _4631_ (.A(_0137_),
    .B(_0133_),
    .X(_1651_));
 sg13g2_a221oi_1 _4632_ (.B2(_0132_),
    .C1(_1253_),
    .B1(_1651_),
    .A1(_1995_),
    .Y(_1652_),
    .A2(_0136_));
 sg13g2_a21oi_1 _4633_ (.A1(_1241_),
    .A2(_1242_),
    .Y(_1653_),
    .B1(_1261_));
 sg13g2_a221oi_1 _4634_ (.B2(_1260_),
    .C1(_1997_),
    .B1(_1653_),
    .A1(_1261_),
    .Y(_1654_),
    .A2(_1273_));
 sg13g2_nor3_1 _4635_ (.A(_1650_),
    .B(_1652_),
    .C(_1654_),
    .Y(_1655_));
 sg13g2_o21ai_1 _4636_ (.B1(_2094_),
    .Y(_1656_),
    .A1(_2088_),
    .A2(_2087_));
 sg13g2_nor4_1 _4637_ (.A(_2091_),
    .B(_2112_),
    .C(_1656_),
    .D(_2108_),
    .Y(_1657_));
 sg13g2_nand2_1 _4638_ (.Y(_1658_),
    .A(_2091_),
    .B(net55));
 sg13g2_nor2_1 _4639_ (.A(net55),
    .B(\g.g_y[7].g_x[4].t.out_sc ),
    .Y(_1659_));
 sg13g2_nor2_1 _4640_ (.A(_2092_),
    .B(net55),
    .Y(_1660_));
 sg13g2_a22oi_1 _4641_ (.Y(_1661_),
    .B1(_1660_),
    .B2(_1656_),
    .A2(_1659_),
    .A1(_2092_));
 sg13g2_o21ai_1 _4642_ (.B1(_1661_),
    .Y(_1662_),
    .A1(_2117_),
    .A2(_1658_));
 sg13g2_o21ai_1 _4643_ (.B1(_1961_),
    .Y(_1663_),
    .A1(_1657_),
    .A2(_1662_));
 sg13g2_o21ai_1 _4644_ (.B1(_1618_),
    .Y(_1664_),
    .A1(_1973_),
    .A2(_1977_));
 sg13g2_and2_1 _4645_ (.A(_1957_),
    .B(_1621_),
    .X(_1665_));
 sg13g2_a221oi_1 _4646_ (.B2(\g.g_y[7].g_x[2].t.out_sc ),
    .C1(_1665_),
    .B1(_1620_),
    .A1(_1956_),
    .Y(_1666_),
    .A2(_1615_));
 sg13g2_nand3_1 _4647_ (.B(_1664_),
    .C(_1666_),
    .A(_1962_),
    .Y(_1667_));
 sg13g2_nand3_1 _4648_ (.B(_1663_),
    .C(_1667_),
    .A(_1650_),
    .Y(_1668_));
 sg13g2_nand2b_1 _4649_ (.Y(\g.g_y[7].g_x[3].t.w_dh ),
    .B(_1668_),
    .A_N(_1655_));
 sg13g2_nand3_1 _4650_ (.B(_1664_),
    .C(_1666_),
    .A(_1961_),
    .Y(_1669_));
 sg13g2_o21ai_1 _4651_ (.B1(_1962_),
    .Y(_1670_),
    .A1(_1657_),
    .A2(_1662_));
 sg13g2_a22oi_1 _4652_ (.Y(_1671_),
    .B1(_1653_),
    .B2(_1260_),
    .A2(_1273_),
    .A1(_1261_));
 sg13g2_a221oi_1 _4653_ (.B2(_0132_),
    .C1(_1997_),
    .B1(_1651_),
    .A1(_1995_),
    .Y(_1672_),
    .A2(_0136_));
 sg13g2_a21oi_1 _4654_ (.A1(_1997_),
    .A2(_1671_),
    .Y(_1673_),
    .B1(_1672_));
 sg13g2_nand3_1 _4655_ (.B(_1670_),
    .C(_1673_),
    .A(_1669_),
    .Y(\g.g_y[7].g_x[3].t.w_na ));
 sg13g2_or4_1 _4656_ (.A(_1959_),
    .B(net78),
    .C(_1652_),
    .D(_1654_),
    .X(_1674_));
 sg13g2_nand4_1 _4657_ (.B(_0246_),
    .C(_1663_),
    .A(_1959_),
    .Y(_1675_),
    .D(_1667_));
 sg13g2_nand2_1 _4658_ (.Y(_1676_),
    .A(\g.g_y[7].g_x[2].t.out_sc ),
    .B(net61));
 sg13g2_nand3_1 _4659_ (.B(_1675_),
    .C(_1676_),
    .A(_1674_),
    .Y(\g.g_y[7].g_x[3].t.w_si ));
 sg13g2_and2_1 _4660_ (.A(net55),
    .B(_2119_),
    .X(_1677_));
 sg13g2_a21oi_1 _4661_ (.A1(_2112_),
    .A2(_2117_),
    .Y(_1678_),
    .B1(_1677_));
 sg13g2_nand2_1 _4662_ (.Y(_1679_),
    .A(\g.g_y[7].g_x[3].t.out_sc ),
    .B(net41));
 sg13g2_o21ai_1 _4663_ (.B1(_1679_),
    .Y(\g.g_y[7].g_x[4].t.w_si ),
    .A1(net59),
    .A2(_1678_));
 sg13g2_inv_1 _4664_ (.Y(_1680_),
    .A(_2085_));
 sg13g2_o21ai_1 _4665_ (.B1(_2124_),
    .Y(_1681_),
    .A1(_2153_),
    .A2(_0220_));
 sg13g2_nand4_1 _4666_ (.B(_2151_),
    .C(_0215_),
    .A(_2125_),
    .Y(_1682_),
    .D(_0216_));
 sg13g2_a21oi_1 _4667_ (.A1(_1681_),
    .A2(_1682_),
    .Y(_1683_),
    .B1(_2132_));
 sg13g2_nand3_1 _4668_ (.B(_1350_),
    .C(_1535_),
    .A(_1331_),
    .Y(_1684_));
 sg13g2_nand2_1 _4669_ (.Y(_1685_),
    .A(_2132_),
    .B(net31));
 sg13g2_a21oi_1 _4670_ (.A1(_1684_),
    .A2(_1352_),
    .Y(_1686_),
    .B1(_1685_));
 sg13g2_nor3_1 _4671_ (.A(_2132_),
    .B(net54),
    .C(_0218_),
    .Y(_1687_));
 sg13g2_nor2_1 _4672_ (.A(_2131_),
    .B(net31),
    .Y(_1688_));
 sg13g2_o21ai_1 _4673_ (.B1(_1688_),
    .Y(_1689_),
    .A1(_1333_),
    .A2(_1345_));
 sg13g2_nand2b_1 _4674_ (.Y(_1690_),
    .B(_1689_),
    .A_N(_1687_));
 sg13g2_nor4_1 _4675_ (.A(_1680_),
    .B(_1683_),
    .C(_1686_),
    .D(_1690_),
    .Y(_1691_));
 sg13g2_and2_1 _4676_ (.A(_2273_),
    .B(_2275_),
    .X(_1692_));
 sg13g2_nor2_1 _4677_ (.A(net48),
    .B(_1692_),
    .Y(_1693_));
 sg13g2_nor2_1 _4678_ (.A(_2089_),
    .B(_2279_),
    .Y(_1694_));
 sg13g2_o21ai_1 _4679_ (.B1(_1694_),
    .Y(_1695_),
    .A1(_2269_),
    .A2(_1693_));
 sg13g2_nand3_1 _4680_ (.B(_2092_),
    .C(net55),
    .A(_2089_),
    .Y(_1696_));
 sg13g2_or4_1 _4681_ (.A(_2088_),
    .B(_2091_),
    .C(net55),
    .D(_2096_),
    .X(_1697_));
 sg13g2_o21ai_1 _4682_ (.B1(_1697_),
    .Y(_1698_),
    .A1(_2117_),
    .A2(_1696_));
 sg13g2_nor2_1 _4683_ (.A(_2088_),
    .B(_2092_),
    .Y(_1699_));
 sg13g2_nand2_1 _4684_ (.Y(_1700_),
    .A(_2084_),
    .B(_1699_));
 sg13g2_nor3_1 _4685_ (.A(_2098_),
    .B(_2108_),
    .C(_1700_),
    .Y(_1701_));
 sg13g2_nor2_1 _4686_ (.A(_2089_),
    .B(_2274_),
    .Y(_1702_));
 sg13g2_nand2_1 _4687_ (.Y(_1703_),
    .A(net48),
    .B(_1702_));
 sg13g2_nor3_1 _4688_ (.A(_0012_),
    .B(_0015_),
    .C(_1703_),
    .Y(_1704_));
 sg13g2_nor2_1 _4689_ (.A(net48),
    .B(_0005_),
    .Y(_1705_));
 sg13g2_a22oi_1 _4690_ (.Y(_1706_),
    .B1(_1699_),
    .B2(_1659_),
    .A2(_1705_),
    .A1(_1702_));
 sg13g2_inv_1 _4691_ (.Y(_1707_),
    .A(_1706_));
 sg13g2_nor4_1 _4692_ (.A(_1698_),
    .B(_1701_),
    .C(_1704_),
    .D(_1707_),
    .Y(_1708_));
 sg13g2_nand3_1 _4693_ (.B(_1695_),
    .C(_1708_),
    .A(_1680_),
    .Y(_1709_));
 sg13g2_nand2b_1 _4694_ (.Y(\g.g_y[7].g_x[5].t.w_dh ),
    .B(_1709_),
    .A_N(_1691_));
 sg13g2_a21o_1 _4695_ (.A2(_0218_),
    .A1(_0217_),
    .B1(net54),
    .X(_1710_));
 sg13g2_a21oi_1 _4696_ (.A1(_1681_),
    .A2(_1710_),
    .Y(_1711_),
    .B1(_2131_));
 sg13g2_nor3_1 _4697_ (.A(_1346_),
    .B(_1333_),
    .C(_1345_),
    .Y(_1712_));
 sg13g2_nand3_1 _4698_ (.B(_1684_),
    .C(_1352_),
    .A(_1346_),
    .Y(_1713_));
 sg13g2_nand3b_1 _4699_ (.B(_1713_),
    .C(_2131_),
    .Y(_1714_),
    .A_N(_1712_));
 sg13g2_or2_1 _4700_ (.X(_1715_),
    .B(_2108_),
    .A(_2098_));
 sg13g2_mux4_1 _4701_ (.S0(_2084_),
    .A0(\g.g_y[7].g_x[4].t.out_sc ),
    .A1(_1715_),
    .A2(_2119_),
    .A3(_2117_),
    .S1(_2092_),
    .X(_1716_));
 sg13g2_or2_1 _4702_ (.X(_1717_),
    .B(_0015_),
    .A(_0012_));
 sg13g2_mux2_1 _4703_ (.A0(_2264_),
    .A1(_2262_),
    .S(_2258_),
    .X(_1718_));
 sg13g2_mux2_1 _4704_ (.A0(_2257_),
    .A1(_1718_),
    .S(_0004_),
    .X(_1719_));
 sg13g2_mux4_1 _4705_ (.S0(_2274_),
    .A0(_0005_),
    .A1(_1692_),
    .A2(_1717_),
    .A3(_1719_),
    .S1(net48),
    .X(_1720_));
 sg13g2_mux2_1 _4706_ (.A0(_1716_),
    .A1(_1720_),
    .S(_2089_),
    .X(_1721_));
 sg13g2_nand3b_1 _4707_ (.B(_1714_),
    .C(_1721_),
    .Y(\g.g_y[7].g_x[5].t.w_na ),
    .A_N(_1711_));
 sg13g2_nand4_1 _4708_ (.B(net64),
    .C(_1695_),
    .A(_2085_),
    .Y(_1722_),
    .D(_1708_));
 sg13g2_nand2_1 _4709_ (.Y(_1723_),
    .A(_1680_),
    .B(_1901_));
 sg13g2_or4_1 _4710_ (.A(_1683_),
    .B(_1686_),
    .C(_1690_),
    .D(_1723_),
    .X(_1724_));
 sg13g2_nand2_1 _4711_ (.Y(_1725_),
    .A(\g.g_y[7].g_x[4].t.out_sc ),
    .B(net61));
 sg13g2_nand3_1 _4712_ (.B(_1724_),
    .C(_1725_),
    .A(_1722_),
    .Y(\g.g_y[7].g_x[5].t.w_si ));
 sg13g2_nand2_1 _4713_ (.Y(_1726_),
    .A(_2273_),
    .B(_2276_));
 sg13g2_nand2_1 _4714_ (.Y(_1727_),
    .A(_2279_),
    .B(_2278_));
 sg13g2_a21oi_1 _4715_ (.A1(_1726_),
    .A2(_1727_),
    .Y(_1728_),
    .B1(_2268_));
 sg13g2_a21oi_1 _4716_ (.A1(_2268_),
    .A2(_1719_),
    .Y(_1729_),
    .B1(_1728_));
 sg13g2_nand2_1 _4717_ (.Y(_1730_),
    .A(\g.g_y[7].g_x[5].t.out_sc ),
    .B(net47));
 sg13g2_o21ai_1 _4718_ (.B1(_1730_),
    .Y(\g.g_y[7].g_x[6].t.w_si ),
    .A1(_2044_),
    .A2(_1729_));
 sg13g2_mux2_1 _4719_ (.A0(\g.g_y[7].g_x[7].t.r_ghl ),
    .A1(_2271_),
    .S(_2270_),
    .X(\g.g_y[7].g_x[7].t.out_r ));
 sg13g2_or2_1 _4720_ (.X(_1731_),
    .B(_1861_),
    .A(_1875_));
 sg13g2_nor2_1 _4721_ (.A(_1855_),
    .B(_1626_),
    .Y(_1732_));
 sg13g2_o21ai_1 _4722_ (.B1(_1732_),
    .Y(_1733_),
    .A1(_1624_),
    .A2(_1731_));
 sg13g2_nor2_1 _4723_ (.A(_1854_),
    .B(_1440_),
    .Y(_1734_));
 sg13g2_o21ai_1 _4724_ (.B1(net65),
    .Y(_1735_),
    .A1(_1853_),
    .A2(_1872_));
 sg13g2_a21oi_1 _4725_ (.A1(_1875_),
    .A2(_1861_),
    .Y(_1736_),
    .B1(_1856_));
 sg13g2_o21ai_1 _4726_ (.B1(_1736_),
    .Y(_1737_),
    .A1(_1734_),
    .A2(_1735_));
 sg13g2_nand3_1 _4727_ (.B(_1733_),
    .C(_1737_),
    .A(_2270_),
    .Y(_1738_));
 sg13g2_nor2_1 _4728_ (.A(_2279_),
    .B(_2268_),
    .Y(_1739_));
 sg13g2_o21ai_1 _4729_ (.B1(_1739_),
    .Y(_1740_),
    .A1(_0012_),
    .A2(_0015_));
 sg13g2_nor2_1 _4730_ (.A(_2274_),
    .B(_2268_),
    .Y(_1741_));
 sg13g2_nor2_1 _4731_ (.A(_2274_),
    .B(_2267_),
    .Y(_1742_));
 sg13g2_and3_1 _4732_ (.X(_1743_),
    .A(_2274_),
    .B(_2268_),
    .C(_0005_));
 sg13g2_a221oi_1 _4733_ (.B2(_2278_),
    .C1(_1743_),
    .B1(_1742_),
    .A1(_1719_),
    .Y(_1744_),
    .A2(_1741_));
 sg13g2_nand3b_1 _4734_ (.B(_1740_),
    .C(_1744_),
    .Y(_1745_),
    .A_N(_2270_));
 sg13g2_nand3b_1 _4735_ (.B(_1738_),
    .C(_1745_),
    .Y(_1746_),
    .A_N(_2183_));
 sg13g2_nand3_1 _4736_ (.B(_1397_),
    .C(_1389_),
    .A(net30),
    .Y(_1747_));
 sg13g2_nor2b_1 _4737_ (.A(net67),
    .B_N(_2264_),
    .Y(_1748_));
 sg13g2_a21oi_1 _4738_ (.A1(_1336_),
    .A2(_1335_),
    .Y(_1749_),
    .B1(_1748_));
 sg13g2_a21oi_1 _4739_ (.A1(_1395_),
    .A2(_1749_),
    .Y(_1750_),
    .B1(_1387_));
 sg13g2_a21o_1 _4740_ (.A2(_1335_),
    .A1(_1336_),
    .B1(_1748_),
    .X(_1751_));
 sg13g2_nand3_1 _4741_ (.B(_1397_),
    .C(_1751_),
    .A(net30),
    .Y(_1752_));
 sg13g2_nand2b_1 _4742_ (.Y(_1753_),
    .B(_1188_),
    .A_N(_1869_));
 sg13g2_o21ai_1 _4743_ (.B1(_1753_),
    .Y(_1754_),
    .A1(_1188_),
    .A2(_1190_));
 sg13g2_a21oi_1 _4744_ (.A1(_1395_),
    .A2(_1754_),
    .Y(_1755_),
    .B1(_1410_));
 sg13g2_a221oi_1 _4745_ (.B2(_1755_),
    .C1(_1385_),
    .B1(_1752_),
    .A1(_1747_),
    .Y(_1756_),
    .A2(_1750_));
 sg13g2_nor3_1 _4746_ (.A(net30),
    .B(_1386_),
    .C(_1397_),
    .Y(_1757_));
 sg13g2_a21o_1 _4747_ (.A2(_1420_),
    .A1(net30),
    .B1(_1757_),
    .X(_1758_));
 sg13g2_o21ai_1 _4748_ (.B1(_1398_),
    .Y(_1759_),
    .A1(_1756_),
    .A2(_1758_));
 sg13g2_nand2b_1 _4749_ (.Y(_1760_),
    .B(_2192_),
    .A_N(_2188_));
 sg13g2_o21ai_1 _4750_ (.B1(_1760_),
    .Y(_1761_),
    .A1(_2192_),
    .A2(_2191_));
 sg13g2_nor4_1 _4751_ (.A(_2195_),
    .B(_2199_),
    .C(_2182_),
    .D(_1761_),
    .Y(_1762_));
 sg13g2_nand2b_1 _4752_ (.Y(_1763_),
    .B(_2195_),
    .A_N(net28));
 sg13g2_nor2_1 _4753_ (.A(_2195_),
    .B(_2201_),
    .Y(_1764_));
 sg13g2_a22oi_1 _4754_ (.Y(_1765_),
    .B1(_1764_),
    .B2(net28),
    .A2(_0258_),
    .A1(_1761_));
 sg13g2_o21ai_1 _4755_ (.B1(_1765_),
    .Y(_1766_),
    .A1(_2206_),
    .A2(_1763_));
 sg13g2_o21ai_1 _4756_ (.B1(_2185_),
    .Y(_1767_),
    .A1(_1762_),
    .A2(_1766_));
 sg13g2_nand3_1 _4757_ (.B(_1759_),
    .C(_1767_),
    .A(_2183_),
    .Y(_1768_));
 sg13g2_nand2_1 _4758_ (.Y(\g.g_y[7].g_x[7].t.w_dh ),
    .A(_1746_),
    .B(_1768_));
 sg13g2_nand3_1 _4759_ (.B(_1740_),
    .C(_1744_),
    .A(_2270_),
    .Y(_1769_));
 sg13g2_nand3b_1 _4760_ (.B(_1733_),
    .C(_1737_),
    .Y(_1770_),
    .A_N(_2270_));
 sg13g2_o21ai_1 _4761_ (.B1(_2185_),
    .Y(_1771_),
    .A1(_1756_),
    .A2(_1758_));
 sg13g2_o21ai_1 _4762_ (.B1(_1398_),
    .Y(_1772_),
    .A1(_1762_),
    .A2(_1766_));
 sg13g2_nand4_1 _4763_ (.B(_1770_),
    .C(_1771_),
    .A(_1769_),
    .Y(\g.g_y[7].g_x[7].t.w_na ),
    .D(_1772_));
 sg13g2_nand4_1 _4764_ (.B(_1902_),
    .C(_1738_),
    .A(_2183_),
    .Y(_1773_),
    .D(_1745_));
 sg13g2_nor2_1 _4765_ (.A(_2183_),
    .B(net78),
    .Y(_1774_));
 sg13g2_nand3_1 _4766_ (.B(_1767_),
    .C(_1774_),
    .A(_1759_),
    .Y(_1775_));
 sg13g2_nand2_1 _4767_ (.Y(_1776_),
    .A(_0005_),
    .B(_2038_));
 sg13g2_nand3_1 _4768_ (.B(_1775_),
    .C(_1776_),
    .A(_1773_),
    .Y(\g.g_y[7].g_x[7].t.w_si ));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _4778__133 (.L_HI(net133));
 sg13g2_buf_1 _4771_ (.A(net119),
    .X(uio_oe[0]));
 sg13g2_buf_1 _4772_ (.A(net120),
    .X(uio_oe[1]));
 sg13g2_buf_1 _4773_ (.A(net121),
    .X(uio_oe[2]));
 sg13g2_buf_1 _4774_ (.A(net122),
    .X(uio_oe[3]));
 sg13g2_buf_1 _4775_ (.A(net123),
    .X(uio_oe[4]));
 sg13g2_buf_1 _4776_ (.A(net124),
    .X(uio_oe[5]));
 sg13g2_buf_1 _4777_ (.A(net125),
    .X(uio_oe[6]));
 sg13g2_buf_1 _4778_ (.A(net133),
    .X(uio_oe[7]));
 sg13g2_buf_1 _4779_ (.A(net126),
    .X(uio_out[0]));
 sg13g2_buf_1 _4780_ (.A(net127),
    .X(uio_out[1]));
 sg13g2_buf_1 _4781_ (.A(net128),
    .X(uio_out[2]));
 sg13g2_buf_1 _4782_ (.A(net129),
    .X(uio_out[3]));
 sg13g2_buf_1 _4783_ (.A(net130),
    .X(uio_out[4]));
 sg13g2_buf_1 _4784_ (.A(net131),
    .X(uio_out[5]));
 sg13g2_buf_1 _4785_ (.A(net132),
    .X(uio_out[6]));
 sg13g2_buf_1 _4786_ (.A(\g.g_y[7].g_x[7].t.out_sc ),
    .X(net16));
 sg13g2_buf_1 _4787_ (.A(\g.g_y[0].g_x[7].t.out_r ),
    .X(net17));
 sg13g2_buf_1 _4788_ (.A(\g.g_y[1].g_x[7].t.out_r ),
    .X(net18));
 sg13g2_buf_1 _4789_ (.A(\g.g_y[2].g_x[7].t.out_r ),
    .X(net19));
 sg13g2_buf_1 _4790_ (.A(\g.g_y[3].g_x[7].t.out_r ),
    .X(net20));
 sg13g2_buf_1 _4791_ (.A(\g.g_y[4].g_x[7].t.out_r ),
    .X(net21));
 sg13g2_buf_1 _4792_ (.A(\g.g_y[5].g_x[7].t.out_r ),
    .X(net22));
 sg13g2_buf_1 _4793_ (.A(\g.g_y[6].g_x[7].t.out_r ),
    .X(net23));
 sg13g2_buf_1 _4794_ (.A(\g.g_y[7].g_x[7].t.out_r ),
    .X(net24));
 sg13g2_dlhq_1 \g.g_y[0].g_x[0].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[0].t.out_sc ),
    .GATE(net104),
    .Q(\g.g_y[0].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[0].g_x[0].t.w_dh ),
    .GATE_N(net107),
    .RESET_B(net134),
    .Q(\g.g_y[0].g_x[0].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[0].g_x[0].t.w_na ),
    .GATE_N(net107),
    .RESET_B(net135),
    .Q(\g.g_y[0].g_x[0].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[0].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[0].t.out_sc ),
    .GATE(net117),
    .Q(\g.g_y[0].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[0].t.r_sc$_DFF_P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net136),
    .D(\g.g_y[0].g_x[0].t.w_si ),
    .Q_N(_2281_),
    .Q(\g.g_y[0].g_x[0].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[0].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[0].t.out_sc ),
    .GATE(net93),
    .Q(\g.g_y[0].g_x[0].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[1].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[1].t.out_sc ),
    .GATE(net104),
    .Q(\g.g_y[0].g_x[1].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[1].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[1].t.out_sc ),
    .GATE(net115),
    .Q(\g.g_y[0].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[1].t.r_sc$_DFF_P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net137),
    .D(\g.g_y[0].g_x[1].t.w_si ),
    .Q_N(_2282_),
    .Q(\g.g_y[0].g_x[1].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[1].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[1].t.out_sc ),
    .GATE(net92),
    .Q(\g.g_y[0].g_x[1].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[2].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[2].t.out_sc ),
    .GATE(net97),
    .Q(\g.g_y[0].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[0].g_x[2].t.w_dh ),
    .GATE_N(net79),
    .RESET_B(net138),
    .Q(\g.g_y[0].g_x[2].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[0].g_x[2].t.w_na ),
    .GATE_N(net79),
    .RESET_B(net139),
    .Q(\g.g_y[0].g_x[2].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[2].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[2].t.out_sc ),
    .GATE(net112),
    .Q(\g.g_y[0].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[2].t.r_sc$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net140),
    .D(\g.g_y[0].g_x[2].t.w_si ),
    .Q_N(_2283_),
    .Q(\g.g_y[0].g_x[2].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[2].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[2].t.out_sc ),
    .GATE(net86),
    .Q(\g.g_y[0].g_x[2].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[3].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[3].t.out_sc ),
    .GATE(net97),
    .Q(\g.g_y[0].g_x[3].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[3].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[3].t.out_sc ),
    .GATE(net109),
    .Q(\g.g_y[0].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[3].t.r_sc$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net141),
    .D(\g.g_y[0].g_x[3].t.w_si ),
    .Q_N(_2284_),
    .Q(\g.g_y[0].g_x[3].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[3].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[3].t.out_sc ),
    .GATE(net87),
    .Q(\g.g_y[0].g_x[3].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[4].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[4].t.out_sc ),
    .GATE(net96),
    .Q(\g.g_y[0].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[0].g_x[4].t.w_dh ),
    .GATE_N(net106),
    .RESET_B(net142),
    .Q(\g.g_y[0].g_x[4].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[0].g_x[4].t.w_na ),
    .GATE_N(net106),
    .RESET_B(net143),
    .Q(\g.g_y[0].g_x[4].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[4].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[4].t.out_sc ),
    .GATE(net109),
    .Q(\g.g_y[0].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[4].t.r_sc$_DFF_P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net144),
    .D(\g.g_y[0].g_x[4].t.w_si ),
    .Q_N(_2285_),
    .Q(\g.g_y[0].g_x[4].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[4].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[4].t.out_sc ),
    .GATE(net85),
    .Q(\g.g_y[0].g_x[4].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[5].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[5].t.out_sc ),
    .GATE(net100),
    .Q(\g.g_y[0].g_x[5].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[5].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[5].t.out_sc ),
    .GATE(net113),
    .Q(\g.g_y[0].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[5].t.r_sc$_DFF_P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net145),
    .D(\g.g_y[0].g_x[5].t.w_si ),
    .Q_N(_2286_),
    .Q(\g.g_y[0].g_x[5].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[5].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[5].t.out_sc ),
    .GATE(net89),
    .Q(\g.g_y[0].g_x[5].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[6].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[6].t.out_sc ),
    .GATE(net100),
    .Q(\g.g_y[0].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[0].g_x[6].t.w_dh ),
    .GATE_N(net80),
    .RESET_B(net146),
    .Q(\g.g_y[0].g_x[6].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[0].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[0].g_x[6].t.w_na ),
    .GATE_N(net80),
    .RESET_B(net147),
    .Q(\g.g_y[0].g_x[6].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[6].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[6].t.out_sc ),
    .GATE(net114),
    .Q(\g.g_y[0].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[6].t.r_sc$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net148),
    .D(\g.g_y[0].g_x[6].t.w_si ),
    .Q_N(_2287_),
    .Q(\g.g_y[0].g_x[6].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[6].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[6].t.out_sc ),
    .GATE(net90),
    .Q(\g.g_y[0].g_x[6].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[7].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[7].t.out_sc ),
    .GATE(net103),
    .Q(\g.g_y[0].g_x[7].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[7].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[7].t.out_sc ),
    .GATE(net115),
    .Q(\g.g_y[0].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[0].g_x[7].t.r_sc$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net149),
    .D(\g.g_y[0].g_x[7].t.w_si ),
    .Q_N(_2288_),
    .Q(\g.g_y[0].g_x[7].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[0].g_x[7].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[0].g_x[7].t.out_sc ),
    .GATE(net91),
    .Q(\g.g_y[0].g_x[7].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[0].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[0].t.out_sc ),
    .GATE(net103),
    .Q(\g.g_y[1].g_x[0].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[0].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[0].t.out_sc ),
    .GATE(net116),
    .Q(\g.g_y[1].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[0].t.r_sc$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net150),
    .D(\g.g_y[1].g_x[0].t.w_si ),
    .Q_N(_2289_),
    .Q(\g.g_y[1].g_x[0].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[0].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[0].t.out_sc ),
    .GATE(net93),
    .Q(\g.g_y[1].g_x[0].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[1].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[1].t.out_sc ),
    .GATE(net102),
    .Q(\g.g_y[1].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[1].g_x[1].t.w_dh ),
    .GATE_N(net75),
    .RESET_B(net151),
    .Q(\g.g_y[1].g_x[1].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[1].g_x[1].t.w_na ),
    .GATE_N(net75),
    .RESET_B(net152),
    .Q(\g.g_y[1].g_x[1].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[1].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[1].t.out_sc ),
    .GATE(net116),
    .Q(\g.g_y[1].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[1].t.r_sc$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net153),
    .D(\g.g_y[1].g_x[1].t.w_si ),
    .Q_N(_2290_),
    .Q(\g.g_y[1].g_x[1].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[1].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[1].t.out_sc ),
    .GATE(net92),
    .Q(\g.g_y[1].g_x[1].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[2].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[2].t.out_sc ),
    .GATE(net98),
    .Q(\g.g_y[1].g_x[2].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[2].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[2].t.out_sc ),
    .GATE(net111),
    .Q(\g.g_y[1].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[2].t.r_sc$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net154),
    .D(\g.g_y[1].g_x[2].t.w_si ),
    .Q_N(_2291_),
    .Q(\g.g_y[1].g_x[2].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[2].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[2].t.out_sc ),
    .GATE(net86),
    .Q(\g.g_y[1].g_x[2].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[3].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[3].t.out_sc ),
    .GATE(net98),
    .Q(\g.g_y[1].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[1].g_x[3].t.w_dh ),
    .GATE_N(net71),
    .RESET_B(net155),
    .Q(\g.g_y[1].g_x[3].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[1].g_x[3].t.w_na ),
    .GATE_N(net71),
    .RESET_B(net156),
    .Q(\g.g_y[1].g_x[3].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[3].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[3].t.out_sc ),
    .GATE(net111),
    .Q(\g.g_y[1].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[3].t.r_sc$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net157),
    .D(\g.g_y[1].g_x[3].t.w_si ),
    .Q_N(_2292_),
    .Q(\g.g_y[1].g_x[3].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[3].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[3].t.out_sc ),
    .GATE(net86),
    .Q(\g.g_y[1].g_x[3].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[4].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[4].t.out_sc ),
    .GATE(net95),
    .Q(\g.g_y[1].g_x[4].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[4].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[4].t.out_sc ),
    .GATE(net108),
    .Q(\g.g_y[1].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[4].t.r_sc$_DFF_P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net158),
    .D(\g.g_y[1].g_x[4].t.w_si ),
    .Q_N(_2293_),
    .Q(\g.g_y[1].g_x[4].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[4].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[4].t.out_sc ),
    .GATE(net84),
    .Q(\g.g_y[1].g_x[4].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[5].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[5].t.out_sc ),
    .GATE(net102),
    .Q(\g.g_y[1].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[1].g_x[5].t.w_dh ),
    .GATE_N(net75),
    .RESET_B(net159),
    .Q(\g.g_y[1].g_x[5].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[1].g_x[5].t.w_na ),
    .GATE_N(net75),
    .RESET_B(net160),
    .Q(\g.g_y[1].g_x[5].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[5].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[5].t.out_sc ),
    .GATE(net116),
    .Q(\g.g_y[1].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[5].t.r_sc$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net161),
    .D(\g.g_y[1].g_x[5].t.w_si ),
    .Q_N(_2294_),
    .Q(\g.g_y[1].g_x[5].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[5].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[5].t.out_sc ),
    .GATE(net89),
    .Q(\g.g_y[1].g_x[5].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[6].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[6].t.out_sc ),
    .GATE(net102),
    .Q(\g.g_y[1].g_x[6].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[6].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[6].t.out_sc ),
    .GATE(net116),
    .Q(\g.g_y[1].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[6].t.r_sc$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net162),
    .D(\g.g_y[1].g_x[6].t.w_si ),
    .Q_N(_2295_),
    .Q(\g.g_y[1].g_x[6].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[6].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[6].t.out_sc ),
    .GATE(net89),
    .Q(\g.g_y[1].g_x[6].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[7].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[7].t.out_sc ),
    .GATE(net103),
    .Q(\g.g_y[1].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[1].g_x[7].t.w_dh ),
    .GATE_N(net72),
    .RESET_B(net163),
    .Q(\g.g_y[1].g_x[7].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[1].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[1].g_x[7].t.w_na ),
    .GATE_N(net72),
    .RESET_B(net164),
    .Q(\g.g_y[1].g_x[7].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[7].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[7].t.out_sc ),
    .GATE(net115),
    .Q(\g.g_y[1].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[1].g_x[7].t.r_sc$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net165),
    .D(\g.g_y[1].g_x[7].t.w_si ),
    .Q_N(_2296_),
    .Q(\g.g_y[1].g_x[7].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[1].g_x[7].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[1].g_x[7].t.out_sc ),
    .GATE(net91),
    .Q(\g.g_y[1].g_x[7].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[0].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[0].t.out_sc ),
    .GATE(net104),
    .Q(\g.g_y[2].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[2].g_x[0].t.w_dh ),
    .GATE_N(net80),
    .RESET_B(net166),
    .Q(\g.g_y[2].g_x[0].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[2].g_x[0].t.w_na ),
    .GATE_N(net80),
    .RESET_B(net167),
    .Q(\g.g_y[2].g_x[0].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[0].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[0].t.out_sc ),
    .GATE(net117),
    .Q(\g.g_y[2].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[0].t.r_sc$_DFF_P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net168),
    .D(\g.g_y[2].g_x[0].t.w_si ),
    .Q_N(_2297_),
    .Q(\g.g_y[2].g_x[0].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[0].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[0].t.out_sc ),
    .GATE(net93),
    .Q(\g.g_y[2].g_x[0].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[1].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[1].t.out_sc ),
    .GATE(net99),
    .Q(\g.g_y[2].g_x[1].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[1].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[1].t.out_sc ),
    .GATE(net110),
    .Q(\g.g_y[2].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[1].t.r_sc$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net169),
    .D(\g.g_y[2].g_x[1].t.w_si ),
    .Q_N(_2298_),
    .Q(\g.g_y[2].g_x[1].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[1].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[1].t.out_sc ),
    .GATE(net87),
    .Q(\g.g_y[2].g_x[1].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[2].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[2].t.out_sc ),
    .GATE(net97),
    .Q(\g.g_y[2].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[2].g_x[2].t.w_dh ),
    .GATE_N(net106),
    .RESET_B(net170),
    .Q(\g.g_y[2].g_x[2].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[2].g_x[2].t.w_na ),
    .GATE_N(net106),
    .RESET_B(net171),
    .Q(\g.g_y[2].g_x[2].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[2].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[2].t.out_sc ),
    .GATE(net110),
    .Q(\g.g_y[2].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[2].t.r_sc$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net172),
    .D(\g.g_y[2].g_x[2].t.w_si ),
    .Q_N(_2299_),
    .Q(\g.g_y[2].g_x[2].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[2].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[2].t.out_sc ),
    .GATE(net86),
    .Q(\g.g_y[2].g_x[2].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[3].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[3].t.out_sc ),
    .GATE(net98),
    .Q(\g.g_y[2].g_x[3].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[3].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[3].t.out_sc ),
    .GATE(net111),
    .Q(\g.g_y[2].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[3].t.r_sc$_DFF_P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net173),
    .D(\g.g_y[2].g_x[3].t.w_si ),
    .Q_N(_2300_),
    .Q(\g.g_y[2].g_x[3].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[3].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[3].t.out_sc ),
    .GATE(net86),
    .Q(\g.g_y[2].g_x[3].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[4].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[4].t.out_sc ),
    .GATE(net95),
    .Q(\g.g_y[2].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[2].g_x[4].t.w_dh ),
    .GATE_N(net79),
    .RESET_B(net174),
    .Q(\g.g_y[2].g_x[4].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[2].g_x[4].t.w_na ),
    .GATE_N(net79),
    .RESET_B(net175),
    .Q(\g.g_y[2].g_x[4].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[4].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[4].t.out_sc ),
    .GATE(net108),
    .Q(\g.g_y[2].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[4].t.r_sc$_DFF_P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net176),
    .D(\g.g_y[2].g_x[4].t.w_si ),
    .Q_N(_2301_),
    .Q(\g.g_y[2].g_x[4].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[4].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[4].t.out_sc ),
    .GATE(net84),
    .Q(\g.g_y[2].g_x[4].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[5].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[5].t.out_sc ),
    .GATE(net97),
    .Q(\g.g_y[2].g_x[5].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[5].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[5].t.out_sc ),
    .GATE(net110),
    .Q(\g.g_y[2].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[5].t.r_sc$_DFF_P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net177),
    .D(\g.g_y[2].g_x[5].t.w_si ),
    .Q_N(_2302_),
    .Q(\g.g_y[2].g_x[5].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[5].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[5].t.out_sc ),
    .GATE(net89),
    .Q(\g.g_y[2].g_x[5].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[6].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[6].t.out_sc ),
    .GATE(net102),
    .Q(\g.g_y[2].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[2].g_x[6].t.w_dh ),
    .GATE_N(net107),
    .RESET_B(net178),
    .Q(\g.g_y[2].g_x[6].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[2].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[2].g_x[6].t.w_na ),
    .GATE_N(net107),
    .RESET_B(net179),
    .Q(\g.g_y[2].g_x[6].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[6].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[6].t.out_sc ),
    .GATE(net115),
    .Q(\g.g_y[2].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[6].t.r_sc$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net180),
    .D(\g.g_y[2].g_x[6].t.w_si ),
    .Q_N(_2303_),
    .Q(\g.g_y[2].g_x[6].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[6].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[6].t.out_sc ),
    .GATE(net92),
    .Q(\g.g_y[2].g_x[6].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[7].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[7].t.out_sc ),
    .GATE(net103),
    .Q(\g.g_y[2].g_x[7].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[7].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[7].t.out_sc ),
    .GATE(net115),
    .Q(\g.g_y[2].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[2].g_x[7].t.r_sc$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net181),
    .D(\g.g_y[2].g_x[7].t.w_si ),
    .Q_N(_2304_),
    .Q(\g.g_y[2].g_x[7].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[2].g_x[7].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[2].g_x[7].t.out_sc ),
    .GATE(net91),
    .Q(\g.g_y[2].g_x[7].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[0].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[0].t.out_sc ),
    .GATE(net103),
    .Q(\g.g_y[3].g_x[0].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[0].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[0].t.out_sc ),
    .GATE(net117),
    .Q(\g.g_y[3].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[0].t.r_sc$_DFF_P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net182),
    .D(\g.g_y[3].g_x[0].t.w_si ),
    .Q_N(_2305_),
    .Q(\g.g_y[3].g_x[0].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[0].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[0].t.out_sc ),
    .GATE(net91),
    .Q(\g.g_y[3].g_x[0].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[1].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[1].t.out_sc ),
    .GATE(net102),
    .Q(\g.g_y[3].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[3].g_x[1].t.w_dh ),
    .GATE_N(net71),
    .RESET_B(net183),
    .Q(\g.g_y[3].g_x[1].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[3].g_x[1].t.w_na ),
    .GATE_N(net71),
    .RESET_B(net184),
    .Q(\g.g_y[3].g_x[1].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[1].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[1].t.out_sc ),
    .GATE(net111),
    .Q(\g.g_y[3].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[1].t.r_sc$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net185),
    .D(\g.g_y[3].g_x[1].t.w_si ),
    .Q_N(_2306_),
    .Q(\g.g_y[3].g_x[1].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[1].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[1].t.out_sc ),
    .GATE(net92),
    .Q(\g.g_y[3].g_x[1].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[2].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[2].t.out_sc ),
    .GATE(net98),
    .Q(\g.g_y[3].g_x[2].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[2].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[2].t.out_sc ),
    .GATE(net111),
    .Q(\g.g_y[3].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[2].t.r_sc$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net186),
    .D(\g.g_y[3].g_x[2].t.w_si ),
    .Q_N(_2307_),
    .Q(\g.g_y[3].g_x[2].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[2].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[2].t.out_sc ),
    .GATE(net86),
    .Q(\g.g_y[3].g_x[2].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[3].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[3].t.out_sc ),
    .GATE(net95),
    .Q(\g.g_y[3].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[3].g_x[3].t.w_dh ),
    .GATE_N(net76),
    .RESET_B(net187),
    .Q(\g.g_y[3].g_x[3].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[3].g_x[3].t.w_na ),
    .GATE_N(net76),
    .RESET_B(net188),
    .Q(\g.g_y[3].g_x[3].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[3].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[3].t.out_sc ),
    .GATE(net108),
    .Q(\g.g_y[3].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[3].t.r_sc$_DFF_P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net189),
    .D(\g.g_y[3].g_x[3].t.w_si ),
    .Q_N(_2308_),
    .Q(\g.g_y[3].g_x[3].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[3].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[3].t.out_sc ),
    .GATE(net84),
    .Q(\g.g_y[3].g_x[3].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[4].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[4].t.out_sc ),
    .GATE(net95),
    .Q(\g.g_y[3].g_x[4].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[4].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[4].t.out_sc ),
    .GATE(net108),
    .Q(\g.g_y[3].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[4].t.r_sc$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net190),
    .D(\g.g_y[3].g_x[4].t.w_si ),
    .Q_N(_2309_),
    .Q(\g.g_y[3].g_x[4].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[4].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[4].t.out_sc ),
    .GATE(net84),
    .Q(\g.g_y[3].g_x[4].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[5].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[5].t.out_sc ),
    .GATE(net95),
    .Q(\g.g_y[3].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[3].g_x[5].t.w_dh ),
    .GATE_N(net71),
    .RESET_B(net191),
    .Q(\g.g_y[3].g_x[5].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[3].g_x[5].t.w_na ),
    .GATE_N(net71),
    .RESET_B(net192),
    .Q(\g.g_y[3].g_x[5].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[5].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[5].t.out_sc ),
    .GATE(net108),
    .Q(\g.g_y[3].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[5].t.r_sc$_DFF_P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net193),
    .D(\g.g_y[3].g_x[5].t.w_si ),
    .Q_N(_2310_),
    .Q(\g.g_y[3].g_x[5].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[5].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[5].t.out_sc ),
    .GATE(net85),
    .Q(\g.g_y[3].g_x[5].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[6].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[6].t.out_sc ),
    .GATE(net100),
    .Q(\g.g_y[3].g_x[6].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[6].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[6].t.out_sc ),
    .GATE(net113),
    .Q(\g.g_y[3].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[6].t.r_sc$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net194),
    .D(\g.g_y[3].g_x[6].t.w_si ),
    .Q_N(_2311_),
    .Q(\g.g_y[3].g_x[6].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[6].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[6].t.out_sc ),
    .GATE(net90),
    .Q(\g.g_y[3].g_x[6].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[7].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[7].t.out_sc ),
    .GATE(net101),
    .Q(\g.g_y[3].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[3].g_x[7].t.w_dh ),
    .GATE_N(net75),
    .RESET_B(net195),
    .Q(\g.g_y[3].g_x[7].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[3].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[3].g_x[7].t.w_na ),
    .GATE_N(net75),
    .RESET_B(net196),
    .Q(\g.g_y[3].g_x[7].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[7].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[7].t.out_sc ),
    .GATE(net114),
    .Q(\g.g_y[3].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[3].g_x[7].t.r_sc$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net197),
    .D(\g.g_y[3].g_x[7].t.w_si ),
    .Q_N(_2312_),
    .Q(\g.g_y[3].g_x[7].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[3].g_x[7].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[3].g_x[7].t.out_sc ),
    .GATE(net94),
    .Q(\g.g_y[3].g_x[7].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[0].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[0].t.out_sc ),
    .GATE(net104),
    .Q(\g.g_y[4].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[4].g_x[0].t.w_dh ),
    .GATE_N(net107),
    .RESET_B(net198),
    .Q(\g.g_y[4].g_x[0].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[4].g_x[0].t.w_na ),
    .GATE_N(net107),
    .RESET_B(net199),
    .Q(\g.g_y[4].g_x[0].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[0].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[0].t.out_sc ),
    .GATE(net116),
    .Q(\g.g_y[4].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[0].t.r_sc$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net200),
    .D(\g.g_y[4].g_x[0].t.w_si ),
    .Q_N(_2313_),
    .Q(\g.g_y[4].g_x[0].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[0].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[0].t.out_sc ),
    .GATE(net91),
    .Q(\g.g_y[4].g_x[0].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[1].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[1].t.out_sc ),
    .GATE(net97),
    .Q(\g.g_y[4].g_x[1].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[1].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[1].t.out_sc ),
    .GATE(net110),
    .Q(\g.g_y[4].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[1].t.r_sc$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net201),
    .D(\g.g_y[4].g_x[1].t.w_si ),
    .Q_N(_2314_),
    .Q(\g.g_y[4].g_x[1].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[1].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[1].t.out_sc ),
    .GATE(net92),
    .Q(\g.g_y[4].g_x[1].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[2].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[2].t.out_sc ),
    .GATE(net98),
    .Q(\g.g_y[4].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[4].g_x[2].t.w_dh ),
    .GATE_N(net79),
    .RESET_B(net202),
    .Q(\g.g_y[4].g_x[2].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[4].g_x[2].t.w_na ),
    .GATE_N(net79),
    .RESET_B(net203),
    .Q(\g.g_y[4].g_x[2].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[2].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[2].t.out_sc ),
    .GATE(net110),
    .Q(\g.g_y[4].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[2].t.r_sc$_DFF_P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net204),
    .D(\g.g_y[4].g_x[2].t.w_si ),
    .Q_N(_2315_),
    .Q(\g.g_y[4].g_x[2].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[2].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[2].t.out_sc ),
    .GATE(net86),
    .Q(\g.g_y[4].g_x[2].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[3].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[3].t.out_sc ),
    .GATE(net95),
    .Q(\g.g_y[4].g_x[3].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[3].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[3].t.out_sc ),
    .GATE(net108),
    .Q(\g.g_y[4].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[3].t.r_sc$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net205),
    .D(\g.g_y[4].g_x[3].t.w_si ),
    .Q_N(_2316_),
    .Q(\g.g_y[4].g_x[3].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[3].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[3].t.out_sc ),
    .GATE(net84),
    .Q(\g.g_y[4].g_x[3].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[4].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[4].t.out_sc ),
    .GATE(net95),
    .Q(\g.g_y[4].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[4].g_x[4].t.w_dh ),
    .GATE_N(net106),
    .RESET_B(net206),
    .Q(\g.g_y[4].g_x[4].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[4].g_x[4].t.w_na ),
    .GATE_N(net106),
    .RESET_B(net207),
    .Q(\g.g_y[4].g_x[4].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[4].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[4].t.out_sc ),
    .GATE(net108),
    .Q(\g.g_y[4].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[4].t.r_sc$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net208),
    .D(\g.g_y[4].g_x[4].t.w_si ),
    .Q_N(_2317_),
    .Q(\g.g_y[4].g_x[4].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[4].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[4].t.out_sc ),
    .GATE(net84),
    .Q(\g.g_y[4].g_x[4].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[5].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[5].t.out_sc ),
    .GATE(net96),
    .Q(\g.g_y[4].g_x[5].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[5].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[5].t.out_sc ),
    .GATE(net109),
    .Q(\g.g_y[4].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[5].t.r_sc$_DFF_P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net209),
    .D(\g.g_y[4].g_x[5].t.w_si ),
    .Q_N(_2318_),
    .Q(\g.g_y[4].g_x[5].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[5].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[5].t.out_sc ),
    .GATE(net85),
    .Q(\g.g_y[4].g_x[5].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[6].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[6].t.out_sc ),
    .GATE(net100),
    .Q(\g.g_y[4].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[4].g_x[6].t.w_dh ),
    .GATE_N(net80),
    .RESET_B(net210),
    .Q(\g.g_y[4].g_x[6].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[4].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[4].g_x[6].t.w_na ),
    .GATE_N(net80),
    .RESET_B(net211),
    .Q(\g.g_y[4].g_x[6].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[6].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[6].t.out_sc ),
    .GATE(net113),
    .Q(\g.g_y[4].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[6].t.r_sc$_DFF_P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net212),
    .D(\g.g_y[4].g_x[6].t.w_si ),
    .Q_N(_2319_),
    .Q(\g.g_y[4].g_x[6].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[6].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[6].t.out_sc ),
    .GATE(net90),
    .Q(\g.g_y[4].g_x[6].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[7].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[7].t.out_sc ),
    .GATE(net101),
    .Q(\g.g_y[4].g_x[7].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[7].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[7].t.out_sc ),
    .GATE(net114),
    .Q(\g.g_y[4].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[4].g_x[7].t.r_sc$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net213),
    .D(\g.g_y[4].g_x[7].t.w_si ),
    .Q_N(_2320_),
    .Q(\g.g_y[4].g_x[7].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[4].g_x[7].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[4].g_x[7].t.out_sc ),
    .GATE(net90),
    .Q(\g.g_y[4].g_x[7].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[0].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[0].t.out_sc ),
    .GATE(net103),
    .Q(\g.g_y[5].g_x[0].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[0].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[0].t.out_sc ),
    .GATE(net115),
    .Q(\g.g_y[5].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[0].t.r_sc$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net214),
    .D(\g.g_y[5].g_x[0].t.w_si ),
    .Q_N(_2321_),
    .Q(\g.g_y[5].g_x[0].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[0].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[0].t.out_sc ),
    .GATE(net91),
    .Q(\g.g_y[5].g_x[0].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[1].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[1].t.out_sc ),
    .GATE(net102),
    .Q(\g.g_y[5].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[5].g_x[1].t.w_dh ),
    .GATE_N(net75),
    .RESET_B(net215),
    .Q(\g.g_y[5].g_x[1].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[5].g_x[1].t.w_na ),
    .GATE_N(net75),
    .RESET_B(net216),
    .Q(\g.g_y[5].g_x[1].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[1].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[1].t.out_sc ),
    .GATE(net116),
    .Q(\g.g_y[5].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[1].t.r_sc$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net217),
    .D(\g.g_y[5].g_x[1].t.w_si ),
    .Q_N(_2322_),
    .Q(\g.g_y[5].g_x[1].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[1].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[1].t.out_sc ),
    .GATE(net92),
    .Q(\g.g_y[5].g_x[1].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[2].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[2].t.out_sc ),
    .GATE(net98),
    .Q(\g.g_y[5].g_x[2].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[2].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[2].t.out_sc ),
    .GATE(net111),
    .Q(\g.g_y[5].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[2].t.r_sc$_DFF_P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net218),
    .D(\g.g_y[5].g_x[2].t.w_si ),
    .Q_N(_2323_),
    .Q(\g.g_y[5].g_x[2].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[2].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[2].t.out_sc ),
    .GATE(net86),
    .Q(\g.g_y[5].g_x[2].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[3].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[3].t.out_sc ),
    .GATE(net98),
    .Q(\g.g_y[5].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[5].g_x[3].t.w_dh ),
    .GATE_N(net71),
    .RESET_B(net219),
    .Q(\g.g_y[5].g_x[3].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[5].g_x[3].t.w_na ),
    .GATE_N(net71),
    .RESET_B(net220),
    .Q(\g.g_y[5].g_x[3].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[3].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[3].t.out_sc ),
    .GATE(net111),
    .Q(\g.g_y[5].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[3].t.r_sc$_DFF_P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net221),
    .D(\g.g_y[5].g_x[3].t.w_si ),
    .Q_N(_2324_),
    .Q(\g.g_y[5].g_x[3].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[3].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[3].t.out_sc ),
    .GATE(net85),
    .Q(\g.g_y[5].g_x[3].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[4].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[4].t.out_sc ),
    .GATE(net95),
    .Q(\g.g_y[5].g_x[4].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[4].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[4].t.out_sc ),
    .GATE(net108),
    .Q(\g.g_y[5].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[4].t.r_sc$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net222),
    .D(\g.g_y[5].g_x[4].t.w_si ),
    .Q_N(_2325_),
    .Q(\g.g_y[5].g_x[4].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[4].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[4].t.out_sc ),
    .GATE(net84),
    .Q(\g.g_y[5].g_x[4].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[5].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[5].t.out_sc ),
    .GATE(net96),
    .Q(\g.g_y[5].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[5].g_x[5].t.w_dh ),
    .GATE_N(net76),
    .RESET_B(net223),
    .Q(\g.g_y[5].g_x[5].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[5].g_x[5].t.w_na ),
    .GATE_N(net76),
    .RESET_B(net224),
    .Q(\g.g_y[5].g_x[5].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[5].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[5].t.out_sc ),
    .GATE(net113),
    .Q(\g.g_y[5].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[5].t.r_sc$_DFF_P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net225),
    .D(\g.g_y[5].g_x[5].t.w_si ),
    .Q_N(_2326_),
    .Q(\g.g_y[5].g_x[5].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[5].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[5].t.out_sc ),
    .GATE(net85),
    .Q(\g.g_y[5].g_x[5].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[6].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[6].t.out_sc ),
    .GATE(net100),
    .Q(\g.g_y[5].g_x[6].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[6].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[6].t.out_sc ),
    .GATE(net113),
    .Q(\g.g_y[5].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[6].t.r_sc$_DFF_P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net226),
    .D(\g.g_y[5].g_x[6].t.w_si ),
    .Q_N(_2327_),
    .Q(\g.g_y[5].g_x[6].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[6].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[6].t.out_sc ),
    .GATE(net89),
    .Q(\g.g_y[5].g_x[6].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[7].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[7].t.out_sc ),
    .GATE(net101),
    .Q(\g.g_y[5].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[5].g_x[7].t.w_dh ),
    .GATE_N(net72),
    .RESET_B(net227),
    .Q(\g.g_y[5].g_x[7].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[5].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[5].g_x[7].t.w_na ),
    .GATE_N(net72),
    .RESET_B(net228),
    .Q(\g.g_y[5].g_x[7].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[7].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[7].t.out_sc ),
    .GATE(net114),
    .Q(\g.g_y[5].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[5].g_x[7].t.r_sc$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net229),
    .D(\g.g_y[5].g_x[7].t.w_si ),
    .Q_N(_2328_),
    .Q(\g.g_y[5].g_x[7].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[5].g_x[7].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[5].g_x[7].t.out_sc ),
    .GATE(net90),
    .Q(\g.g_y[5].g_x[7].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[0].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[0].t.out_sc ),
    .GATE(net103),
    .Q(\g.g_y[6].g_x[0].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[6].g_x[0].t.w_dh ),
    .GATE_N(net80),
    .RESET_B(net230),
    .Q(\g.g_y[6].g_x[0].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[6].g_x[0].t.w_na ),
    .GATE_N(net80),
    .RESET_B(net231),
    .Q(\g.g_y[6].g_x[0].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[0].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[0].t.out_sc ),
    .GATE(net115),
    .Q(\g.g_y[6].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[0].t.r_sc$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net232),
    .D(\g.g_y[6].g_x[0].t.w_si ),
    .Q_N(_2329_),
    .Q(\g.g_y[6].g_x[0].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[0].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[0].t.out_sc ),
    .GATE(net91),
    .Q(\g.g_y[6].g_x[0].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[1].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[1].t.out_sc ),
    .GATE(net102),
    .Q(\g.g_y[6].g_x[1].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[1].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[1].t.out_sc ),
    .GATE(net116),
    .Q(\g.g_y[6].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[1].t.r_sc$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net233),
    .D(\g.g_y[6].g_x[1].t.w_si ),
    .Q_N(_2330_),
    .Q(\g.g_y[6].g_x[1].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[1].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[1].t.out_sc ),
    .GATE(net92),
    .Q(\g.g_y[6].g_x[1].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[2].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[2].t.out_sc ),
    .GATE(net97),
    .Q(\g.g_y[6].g_x[2].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[6].g_x[2].t.w_dh ),
    .GATE_N(net106),
    .RESET_B(net234),
    .Q(\g.g_y[6].g_x[2].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[6].g_x[2].t.w_na ),
    .GATE_N(net106),
    .RESET_B(net235),
    .Q(\g.g_y[6].g_x[2].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[2].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[2].t.out_sc ),
    .GATE(net110),
    .Q(\g.g_y[6].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[2].t.r_sc$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net236),
    .D(\g.g_y[6].g_x[2].t.w_si ),
    .Q_N(_2331_),
    .Q(\g.g_y[6].g_x[2].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[2].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[2].t.out_sc ),
    .GATE(net87),
    .Q(\g.g_y[6].g_x[2].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[3].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[3].t.out_sc ),
    .GATE(net96),
    .Q(\g.g_y[6].g_x[3].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[3].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[3].t.out_sc ),
    .GATE(net109),
    .Q(\g.g_y[6].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[3].t.r_sc$_DFF_P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net237),
    .D(\g.g_y[6].g_x[3].t.w_si ),
    .Q_N(_2332_),
    .Q(\g.g_y[6].g_x[3].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[3].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[3].t.out_sc ),
    .GATE(net85),
    .Q(\g.g_y[6].g_x[3].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[4].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[4].t.out_sc ),
    .GATE(net96),
    .Q(\g.g_y[6].g_x[4].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[6].g_x[4].t.w_dh ),
    .GATE_N(net79),
    .RESET_B(net238),
    .Q(\g.g_y[6].g_x[4].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[6].g_x[4].t.w_na ),
    .GATE_N(net79),
    .RESET_B(net239),
    .Q(\g.g_y[6].g_x[4].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[4].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[4].t.out_sc ),
    .GATE(net109),
    .Q(\g.g_y[6].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[4].t.r_sc$_DFF_P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net240),
    .D(\g.g_y[6].g_x[4].t.w_si ),
    .Q_N(_2333_),
    .Q(\g.g_y[6].g_x[4].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[4].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[4].t.out_sc ),
    .GATE(net84),
    .Q(\g.g_y[6].g_x[4].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[5].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[5].t.out_sc ),
    .GATE(net100),
    .Q(\g.g_y[6].g_x[5].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[5].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[5].t.out_sc ),
    .GATE(net113),
    .Q(\g.g_y[6].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[5].t.r_sc$_DFF_P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net241),
    .D(\g.g_y[6].g_x[5].t.w_si ),
    .Q_N(_2334_),
    .Q(\g.g_y[6].g_x[5].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[5].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[5].t.out_sc ),
    .GATE(net89),
    .Q(\g.g_y[6].g_x[5].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[6].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[6].t.out_sc ),
    .GATE(net100),
    .Q(\g.g_y[6].g_x[6].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[6].g_x[6].t.w_dh ),
    .GATE_N(net107),
    .RESET_B(net242),
    .Q(\g.g_y[6].g_x[6].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[6].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[6].g_x[6].t.w_na ),
    .GATE_N(net107),
    .RESET_B(net243),
    .Q(\g.g_y[6].g_x[6].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[6].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[6].t.out_sc ),
    .GATE(net114),
    .Q(\g.g_y[6].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[6].t.r_sc$_DFF_P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net244),
    .D(\g.g_y[6].g_x[6].t.w_si ),
    .Q_N(_2335_),
    .Q(\g.g_y[6].g_x[6].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[6].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[6].t.out_sc ),
    .GATE(net90),
    .Q(\g.g_y[6].g_x[6].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[7].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[7].t.out_sc ),
    .GATE(net101),
    .Q(\g.g_y[6].g_x[7].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[7].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[7].t.out_sc ),
    .GATE(net114),
    .Q(\g.g_y[6].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[6].g_x[7].t.r_sc$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net245),
    .D(\g.g_y[6].g_x[7].t.w_si ),
    .Q_N(_2336_),
    .Q(\g.g_y[6].g_x[7].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[6].g_x[7].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[6].g_x[7].t.out_sc ),
    .GATE(net90),
    .Q(\g.g_y[6].g_x[7].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[0].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[0].t.out_sc ),
    .GATE(net103),
    .Q(\g.g_y[7].g_x[0].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[0].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[0].t.out_sc ),
    .GATE(net115),
    .Q(\g.g_y[7].g_x[0].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[0].t.r_sc$_DFF_P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net246),
    .D(\g.g_y[7].g_x[0].t.w_si ),
    .Q_N(_2337_),
    .Q(\g.g_y[7].g_x[0].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[0].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[0].t.out_sc ),
    .GATE(net91),
    .Q(\g.g_y[7].g_x[0].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[1].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[1].t.out_sc ),
    .GATE(net102),
    .Q(\g.g_y[7].g_x[1].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[7].g_x[1].t.w_dh ),
    .GATE_N(net72),
    .RESET_B(net247),
    .Q(\g.g_y[7].g_x[1].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[7].g_x[1].t.w_na ),
    .GATE_N(net72),
    .RESET_B(net248),
    .Q(\g.g_y[7].g_x[1].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[1].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[1].t.out_sc ),
    .GATE(net116),
    .Q(\g.g_y[7].g_x[1].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[1].t.r_sc$_DFF_P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net249),
    .D(\g.g_y[7].g_x[1].t.w_si ),
    .Q_N(_2338_),
    .Q(\g.g_y[7].g_x[1].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[1].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[1].t.out_sc ),
    .GATE(net92),
    .Q(\g.g_y[7].g_x[1].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[2].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[2].t.out_sc ),
    .GATE(net97),
    .Q(\g.g_y[7].g_x[2].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[2].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[2].t.out_sc ),
    .GATE(net110),
    .Q(\g.g_y[7].g_x[2].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[2].t.r_sc$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net250),
    .D(\g.g_y[7].g_x[2].t.w_si ),
    .Q_N(_2339_),
    .Q(\g.g_y[7].g_x[2].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[2].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[2].t.out_sc ),
    .GATE(net87),
    .Q(\g.g_y[7].g_x[2].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[3].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[3].t.out_sc ),
    .GATE(net97),
    .Q(\g.g_y[7].g_x[3].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[7].g_x[3].t.w_dh ),
    .GATE_N(net76),
    .RESET_B(net251),
    .Q(\g.g_y[7].g_x[3].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[7].g_x[3].t.w_na ),
    .GATE_N(net76),
    .RESET_B(net252),
    .Q(\g.g_y[7].g_x[3].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[3].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[3].t.out_sc ),
    .GATE(net110),
    .Q(\g.g_y[7].g_x[3].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[3].t.r_sc$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net253),
    .D(\g.g_y[7].g_x[3].t.w_si ),
    .Q_N(_2340_),
    .Q(\g.g_y[7].g_x[3].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[3].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[3].t.out_sc ),
    .GATE(net87),
    .Q(\g.g_y[7].g_x[3].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[4].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[4].t.out_sc ),
    .GATE(net96),
    .Q(\g.g_y[7].g_x[4].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[4].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[4].t.out_sc ),
    .GATE(net109),
    .Q(\g.g_y[7].g_x[4].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[4].t.r_sc$_DFF_P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net254),
    .D(\g.g_y[7].g_x[4].t.w_si ),
    .Q_N(_2341_),
    .Q(\g.g_y[7].g_x[4].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[4].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[4].t.out_sc ),
    .GATE(net85),
    .Q(\g.g_y[7].g_x[4].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[5].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[5].t.out_sc ),
    .GATE(net100),
    .Q(\g.g_y[7].g_x[5].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[7].g_x[5].t.w_dh ),
    .GATE_N(net72),
    .RESET_B(net255),
    .Q(\g.g_y[7].g_x[5].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[7].g_x[5].t.w_na ),
    .GATE_N(net72),
    .RESET_B(net256),
    .Q(\g.g_y[7].g_x[5].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[5].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[5].t.out_sc ),
    .GATE(net113),
    .Q(\g.g_y[7].g_x[5].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[5].t.r_sc$_DFF_P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net257),
    .D(\g.g_y[7].g_x[5].t.w_si ),
    .Q_N(_2342_),
    .Q(\g.g_y[7].g_x[5].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[5].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[5].t.out_sc ),
    .GATE(net89),
    .Q(\g.g_y[7].g_x[5].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[6].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[6].t.out_sc ),
    .GATE(net101),
    .Q(\g.g_y[7].g_x[6].t.r_d ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[6].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[6].t.out_sc ),
    .GATE(net113),
    .Q(\g.g_y[7].g_x[6].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[6].t.r_sc$_DFF_P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net258),
    .D(\g.g_y[7].g_x[6].t.w_si ),
    .Q_N(_2343_),
    .Q(\g.g_y[7].g_x[6].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[6].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[6].t.out_sc ),
    .GATE(net89),
    .Q(\g.g_y[7].g_x[6].t.r_v ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[7].t.r_d$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[7].t.out_sc ),
    .GATE(net101),
    .Q(\g.g_y[7].g_x[7].t.r_d ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[7].g_x[7].t.w_dh ),
    .GATE_N(\g.g_y[1].g_x[1].t.in_lb ),
    .RESET_B(net259),
    .Q(\g.g_y[7].g_x[7].t.r_ghl ));
 sg13g2_dllrq_1 \g.g_y[7].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N  (.D(\g.g_y[7].g_x[7].t.w_na ),
    .GATE_N(net76),
    .RESET_B(net260),
    .Q(\g.g_y[7].g_x[7].t.r_gnl ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[7].t.r_h$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[7].t.out_sc ),
    .GATE(net114),
    .Q(\g.g_y[7].g_x[7].t.r_h ));
 sg13g2_dfrbp_1 \g.g_y[7].g_x[7].t.r_sc$_DFF_P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net261),
    .D(\g.g_y[7].g_x[7].t.w_si ),
    .Q_N(_2280_),
    .Q(\g.g_y[7].g_x[7].t.out_sc ));
 sg13g2_dlhq_1 \g.g_y[7].g_x[7].t.r_v$_DLATCH_P_._TECHMAP_DLATCH_P  (.D(\g.g_y[7].g_x[7].t.out_sc ),
    .GATE(net94),
    .Q(\g.g_y[7].g_x[7].t.r_v ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[7]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout25 (.A(_1187_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0394_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0086_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_2199_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1832_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1394_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1346_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1344_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1186_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1184_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1090_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1009_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0949_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0894_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0890_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0852_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0751_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0585_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0480_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0454_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0246_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0193_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0109_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2267_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_2258_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_2256_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_2218_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_2175_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2139_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2124_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2084_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_2063_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2057_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2047_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_2044_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_2040_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_2038_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_2006_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1905_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1902_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1862_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1782_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1336_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1197_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1097_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0837_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(\g.g_y[1].g_x[3].t.in_lb ),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(\g.g_y[1].g_x[3].t.in_lb ),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0113_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0111_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(net76),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(\g.g_y[1].g_x[1].t.in_lb ),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_2037_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_2034_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(\g.g_y[0].g_x[2].t.in_lb ),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(\g.g_y[0].g_x[2].t.in_lb ),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1901_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1894_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1793_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(net88),
    .X(net84));
 sg13g2_buf_1 fanout85 (.A(net88),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(net88),
    .X(net86));
 sg13g2_buf_1 fanout87 (.A(net88),
    .X(net87));
 sg13g2_buf_1 fanout88 (.A(\g.cfg_v ),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(net90),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(net94),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(net93),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(net94),
    .X(net92));
 sg13g2_buf_1 fanout93 (.A(net94),
    .X(net93));
 sg13g2_buf_1 fanout94 (.A(\g.cfg_v ),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(net99),
    .X(net95));
 sg13g2_buf_1 fanout96 (.A(net99),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(net99),
    .X(net98));
 sg13g2_buf_1 fanout99 (.A(net105),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(net105),
    .X(net100));
 sg13g2_buf_1 fanout101 (.A(net105),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(net104),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_1 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_1 fanout105 (.A(\g.cfg_d ),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(\g.g_y[0].g_x[0].t.in_lb ),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(\g.g_y[0].g_x[0].t.in_lb ),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(net112),
    .X(net108));
 sg13g2_buf_1 fanout109 (.A(net112),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(net111),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(net112),
    .X(net111));
 sg13g2_buf_1 fanout112 (.A(\g.cfg_h ),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(net118),
    .X(net113));
 sg13g2_buf_1 fanout114 (.A(net118),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(net117),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(net118),
    .X(net116));
 sg13g2_buf_1 fanout117 (.A(net118),
    .X(net117));
 sg13g2_buf_1 fanout118 (.A(\g.cfg_h ),
    .X(net118));
 sg13g2_tielo _4771__119 (.L_LO(net119));
 sg13g2_tielo _4772__120 (.L_LO(net120));
 sg13g2_tielo _4773__121 (.L_LO(net121));
 sg13g2_tielo _4774__122 (.L_LO(net122));
 sg13g2_tielo _4775__123 (.L_LO(net123));
 sg13g2_tielo _4776__124 (.L_LO(net124));
 sg13g2_tielo _4777__125 (.L_LO(net125));
 sg13g2_tielo _4779__126 (.L_LO(net126));
 sg13g2_tielo _4780__127 (.L_LO(net127));
 sg13g2_tielo _4781__128 (.L_LO(net128));
 sg13g2_tielo _4782__129 (.L_LO(net129));
 sg13g2_tielo _4783__130 (.L_LO(net130));
 sg13g2_tielo _4784__131 (.L_LO(net131));
 sg13g2_tielo _4785__132 (.L_LO(net132));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_134  (.L_HI(net134));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_135  (.L_HI(net135));
 sg13g2_tiehi \g.g_y[0].g_x[0].t.r_sc$_DFF_P__136  (.L_HI(net136));
 sg13g2_tiehi \g.g_y[0].g_x[1].t.r_sc$_DFF_P__137  (.L_HI(net137));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_138  (.L_HI(net138));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_139  (.L_HI(net139));
 sg13g2_tiehi \g.g_y[0].g_x[2].t.r_sc$_DFF_P__140  (.L_HI(net140));
 sg13g2_tiehi \g.g_y[0].g_x[3].t.r_sc$_DFF_P__141  (.L_HI(net141));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_142  (.L_HI(net142));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_143  (.L_HI(net143));
 sg13g2_tiehi \g.g_y[0].g_x[4].t.r_sc$_DFF_P__144  (.L_HI(net144));
 sg13g2_tiehi \g.g_y[0].g_x[5].t.r_sc$_DFF_P__145  (.L_HI(net145));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_146  (.L_HI(net146));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_147  (.L_HI(net147));
 sg13g2_tiehi \g.g_y[0].g_x[6].t.r_sc$_DFF_P__148  (.L_HI(net148));
 sg13g2_tiehi \g.g_y[0].g_x[7].t.r_sc$_DFF_P__149  (.L_HI(net149));
 sg13g2_tiehi \g.g_y[1].g_x[0].t.r_sc$_DFF_P__150  (.L_HI(net150));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_151  (.L_HI(net151));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_152  (.L_HI(net152));
 sg13g2_tiehi \g.g_y[1].g_x[1].t.r_sc$_DFF_P__153  (.L_HI(net153));
 sg13g2_tiehi \g.g_y[1].g_x[2].t.r_sc$_DFF_P__154  (.L_HI(net154));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_155  (.L_HI(net155));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_156  (.L_HI(net156));
 sg13g2_tiehi \g.g_y[1].g_x[3].t.r_sc$_DFF_P__157  (.L_HI(net157));
 sg13g2_tiehi \g.g_y[1].g_x[4].t.r_sc$_DFF_P__158  (.L_HI(net158));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_159  (.L_HI(net159));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_160  (.L_HI(net160));
 sg13g2_tiehi \g.g_y[1].g_x[5].t.r_sc$_DFF_P__161  (.L_HI(net161));
 sg13g2_tiehi \g.g_y[1].g_x[6].t.r_sc$_DFF_P__162  (.L_HI(net162));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_163  (.L_HI(net163));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_164  (.L_HI(net164));
 sg13g2_tiehi \g.g_y[1].g_x[7].t.r_sc$_DFF_P__165  (.L_HI(net165));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_166  (.L_HI(net166));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_167  (.L_HI(net167));
 sg13g2_tiehi \g.g_y[2].g_x[0].t.r_sc$_DFF_P__168  (.L_HI(net168));
 sg13g2_tiehi \g.g_y[2].g_x[1].t.r_sc$_DFF_P__169  (.L_HI(net169));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_170  (.L_HI(net170));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_171  (.L_HI(net171));
 sg13g2_tiehi \g.g_y[2].g_x[2].t.r_sc$_DFF_P__172  (.L_HI(net172));
 sg13g2_tiehi \g.g_y[2].g_x[3].t.r_sc$_DFF_P__173  (.L_HI(net173));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_174  (.L_HI(net174));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_175  (.L_HI(net175));
 sg13g2_tiehi \g.g_y[2].g_x[4].t.r_sc$_DFF_P__176  (.L_HI(net176));
 sg13g2_tiehi \g.g_y[2].g_x[5].t.r_sc$_DFF_P__177  (.L_HI(net177));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_178  (.L_HI(net178));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_179  (.L_HI(net179));
 sg13g2_tiehi \g.g_y[2].g_x[6].t.r_sc$_DFF_P__180  (.L_HI(net180));
 sg13g2_tiehi \g.g_y[2].g_x[7].t.r_sc$_DFF_P__181  (.L_HI(net181));
 sg13g2_tiehi \g.g_y[3].g_x[0].t.r_sc$_DFF_P__182  (.L_HI(net182));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_183  (.L_HI(net183));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_184  (.L_HI(net184));
 sg13g2_tiehi \g.g_y[3].g_x[1].t.r_sc$_DFF_P__185  (.L_HI(net185));
 sg13g2_tiehi \g.g_y[3].g_x[2].t.r_sc$_DFF_P__186  (.L_HI(net186));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_187  (.L_HI(net187));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_188  (.L_HI(net188));
 sg13g2_tiehi \g.g_y[3].g_x[3].t.r_sc$_DFF_P__189  (.L_HI(net189));
 sg13g2_tiehi \g.g_y[3].g_x[4].t.r_sc$_DFF_P__190  (.L_HI(net190));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_191  (.L_HI(net191));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_192  (.L_HI(net192));
 sg13g2_tiehi \g.g_y[3].g_x[5].t.r_sc$_DFF_P__193  (.L_HI(net193));
 sg13g2_tiehi \g.g_y[3].g_x[6].t.r_sc$_DFF_P__194  (.L_HI(net194));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_195  (.L_HI(net195));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_196  (.L_HI(net196));
 sg13g2_tiehi \g.g_y[3].g_x[7].t.r_sc$_DFF_P__197  (.L_HI(net197));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_198  (.L_HI(net198));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_199  (.L_HI(net199));
 sg13g2_tiehi \g.g_y[4].g_x[0].t.r_sc$_DFF_P__200  (.L_HI(net200));
 sg13g2_tiehi \g.g_y[4].g_x[1].t.r_sc$_DFF_P__201  (.L_HI(net201));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_202  (.L_HI(net202));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_203  (.L_HI(net203));
 sg13g2_tiehi \g.g_y[4].g_x[2].t.r_sc$_DFF_P__204  (.L_HI(net204));
 sg13g2_tiehi \g.g_y[4].g_x[3].t.r_sc$_DFF_P__205  (.L_HI(net205));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_206  (.L_HI(net206));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_207  (.L_HI(net207));
 sg13g2_tiehi \g.g_y[4].g_x[4].t.r_sc$_DFF_P__208  (.L_HI(net208));
 sg13g2_tiehi \g.g_y[4].g_x[5].t.r_sc$_DFF_P__209  (.L_HI(net209));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_210  (.L_HI(net210));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_211  (.L_HI(net211));
 sg13g2_tiehi \g.g_y[4].g_x[6].t.r_sc$_DFF_P__212  (.L_HI(net212));
 sg13g2_tiehi \g.g_y[4].g_x[7].t.r_sc$_DFF_P__213  (.L_HI(net213));
 sg13g2_tiehi \g.g_y[5].g_x[0].t.r_sc$_DFF_P__214  (.L_HI(net214));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_215  (.L_HI(net215));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_216  (.L_HI(net216));
 sg13g2_tiehi \g.g_y[5].g_x[1].t.r_sc$_DFF_P__217  (.L_HI(net217));
 sg13g2_tiehi \g.g_y[5].g_x[2].t.r_sc$_DFF_P__218  (.L_HI(net218));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_219  (.L_HI(net219));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_220  (.L_HI(net220));
 sg13g2_tiehi \g.g_y[5].g_x[3].t.r_sc$_DFF_P__221  (.L_HI(net221));
 sg13g2_tiehi \g.g_y[5].g_x[4].t.r_sc$_DFF_P__222  (.L_HI(net222));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_223  (.L_HI(net223));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_224  (.L_HI(net224));
 sg13g2_tiehi \g.g_y[5].g_x[5].t.r_sc$_DFF_P__225  (.L_HI(net225));
 sg13g2_tiehi \g.g_y[5].g_x[6].t.r_sc$_DFF_P__226  (.L_HI(net226));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_227  (.L_HI(net227));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_228  (.L_HI(net228));
 sg13g2_tiehi \g.g_y[5].g_x[7].t.r_sc$_DFF_P__229  (.L_HI(net229));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_230  (.L_HI(net230));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_231  (.L_HI(net231));
 sg13g2_tiehi \g.g_y[6].g_x[0].t.r_sc$_DFF_P__232  (.L_HI(net232));
 sg13g2_tiehi \g.g_y[6].g_x[1].t.r_sc$_DFF_P__233  (.L_HI(net233));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_234  (.L_HI(net234));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_235  (.L_HI(net235));
 sg13g2_tiehi \g.g_y[6].g_x[2].t.r_sc$_DFF_P__236  (.L_HI(net236));
 sg13g2_tiehi \g.g_y[6].g_x[3].t.r_sc$_DFF_P__237  (.L_HI(net237));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_238  (.L_HI(net238));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_239  (.L_HI(net239));
 sg13g2_tiehi \g.g_y[6].g_x[4].t.r_sc$_DFF_P__240  (.L_HI(net240));
 sg13g2_tiehi \g.g_y[6].g_x[5].t.r_sc$_DFF_P__241  (.L_HI(net241));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_242  (.L_HI(net242));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_243  (.L_HI(net243));
 sg13g2_tiehi \g.g_y[6].g_x[6].t.r_sc$_DFF_P__244  (.L_HI(net244));
 sg13g2_tiehi \g.g_y[6].g_x[7].t.r_sc$_DFF_P__245  (.L_HI(net245));
 sg13g2_tiehi \g.g_y[7].g_x[0].t.r_sc$_DFF_P__246  (.L_HI(net246));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_247  (.L_HI(net247));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_248  (.L_HI(net248));
 sg13g2_tiehi \g.g_y[7].g_x[1].t.r_sc$_DFF_P__249  (.L_HI(net249));
 sg13g2_tiehi \g.g_y[7].g_x[2].t.r_sc$_DFF_P__250  (.L_HI(net250));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_251  (.L_HI(net251));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_252  (.L_HI(net252));
 sg13g2_tiehi \g.g_y[7].g_x[3].t.r_sc$_DFF_P__253  (.L_HI(net253));
 sg13g2_tiehi \g.g_y[7].g_x[4].t.r_sc$_DFF_P__254  (.L_HI(net254));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_255  (.L_HI(net255));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_256  (.L_HI(net256));
 sg13g2_tiehi \g.g_y[7].g_x[5].t.r_sc$_DFF_P__257  (.L_HI(net257));
 sg13g2_tiehi \g.g_y[7].g_x[6].t.r_sc$_DFF_P__258  (.L_HI(net258));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_ghl$_DLATCH_N_._TECHMAP_DLATCH_N_259  (.L_HI(net259));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_gnl$_DLATCH_N_._TECHMAP_DLATCH_N_260  (.L_HI(net260));
 sg13g2_tiehi \g.g_y[7].g_x[7].t.r_sc$_DFF_P__261  (.L_HI(net261));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_4 FILLER_0_224 ();
 sg13g2_fill_2 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_fill_2 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_fill_2 FILLER_1_161 ();
 sg13g2_fill_1 FILLER_1_163 ();
 sg13g2_decap_4 FILLER_1_185 ();
 sg13g2_fill_1 FILLER_1_189 ();
 sg13g2_fill_2 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_248 ();
 sg13g2_decap_4 FILLER_1_255 ();
 sg13g2_fill_1 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_fill_1 FILLER_2_161 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_fill_2 FILLER_2_188 ();
 sg13g2_decap_8 FILLER_2_194 ();
 sg13g2_decap_4 FILLER_2_201 ();
 sg13g2_fill_1 FILLER_2_205 ();
 sg13g2_fill_2 FILLER_2_223 ();
 sg13g2_fill_1 FILLER_2_225 ();
 sg13g2_fill_1 FILLER_2_248 ();
 sg13g2_fill_2 FILLER_2_252 ();
 sg13g2_fill_1 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_260 ();
 sg13g2_decap_8 FILLER_2_267 ();
 sg13g2_fill_1 FILLER_2_274 ();
 sg13g2_decap_4 FILLER_2_279 ();
 sg13g2_fill_1 FILLER_2_283 ();
 sg13g2_decap_4 FILLER_2_289 ();
 sg13g2_decap_8 FILLER_2_297 ();
 sg13g2_decap_8 FILLER_2_304 ();
 sg13g2_decap_8 FILLER_2_311 ();
 sg13g2_decap_8 FILLER_2_318 ();
 sg13g2_decap_8 FILLER_2_325 ();
 sg13g2_decap_8 FILLER_2_332 ();
 sg13g2_decap_8 FILLER_2_339 ();
 sg13g2_decap_8 FILLER_2_346 ();
 sg13g2_decap_8 FILLER_2_353 ();
 sg13g2_decap_8 FILLER_2_360 ();
 sg13g2_decap_8 FILLER_2_367 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_2_409 ();
 sg13g2_decap_8 FILLER_2_416 ();
 sg13g2_decap_8 FILLER_2_423 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_4 FILLER_3_175 ();
 sg13g2_fill_1 FILLER_3_179 ();
 sg13g2_fill_2 FILLER_3_198 ();
 sg13g2_fill_1 FILLER_3_204 ();
 sg13g2_fill_1 FILLER_3_217 ();
 sg13g2_fill_1 FILLER_3_235 ();
 sg13g2_fill_2 FILLER_3_261 ();
 sg13g2_decap_8 FILLER_3_272 ();
 sg13g2_fill_2 FILLER_3_279 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_fill_2 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_170 ();
 sg13g2_fill_2 FILLER_4_175 ();
 sg13g2_fill_1 FILLER_4_177 ();
 sg13g2_fill_1 FILLER_4_182 ();
 sg13g2_fill_2 FILLER_4_216 ();
 sg13g2_fill_1 FILLER_4_267 ();
 sg13g2_decap_8 FILLER_4_306 ();
 sg13g2_decap_8 FILLER_4_313 ();
 sg13g2_decap_8 FILLER_4_320 ();
 sg13g2_decap_8 FILLER_4_327 ();
 sg13g2_decap_8 FILLER_4_334 ();
 sg13g2_decap_8 FILLER_4_341 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_8 FILLER_4_404 ();
 sg13g2_decap_8 FILLER_4_411 ();
 sg13g2_decap_8 FILLER_4_418 ();
 sg13g2_decap_4 FILLER_4_425 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_4 FILLER_5_147 ();
 sg13g2_fill_2 FILLER_5_155 ();
 sg13g2_fill_1 FILLER_5_157 ();
 sg13g2_fill_1 FILLER_5_179 ();
 sg13g2_fill_2 FILLER_5_216 ();
 sg13g2_fill_1 FILLER_5_222 ();
 sg13g2_fill_1 FILLER_5_233 ();
 sg13g2_fill_2 FILLER_5_239 ();
 sg13g2_fill_1 FILLER_5_241 ();
 sg13g2_decap_4 FILLER_5_274 ();
 sg13g2_fill_1 FILLER_5_278 ();
 sg13g2_fill_2 FILLER_5_289 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_decap_8 FILLER_5_332 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_decap_8 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_409 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_4 FILLER_6_140 ();
 sg13g2_fill_1 FILLER_6_144 ();
 sg13g2_fill_2 FILLER_6_175 ();
 sg13g2_fill_1 FILLER_6_177 ();
 sg13g2_fill_1 FILLER_6_196 ();
 sg13g2_fill_2 FILLER_6_202 ();
 sg13g2_fill_2 FILLER_6_208 ();
 sg13g2_fill_2 FILLER_6_236 ();
 sg13g2_fill_1 FILLER_6_241 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_4 FILLER_6_270 ();
 sg13g2_fill_2 FILLER_6_274 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_303 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_4 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_decap_8 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_4 FILLER_7_161 ();
 sg13g2_fill_2 FILLER_7_199 ();
 sg13g2_decap_8 FILLER_7_205 ();
 sg13g2_fill_2 FILLER_7_212 ();
 sg13g2_fill_2 FILLER_7_219 ();
 sg13g2_fill_2 FILLER_7_226 ();
 sg13g2_fill_2 FILLER_7_236 ();
 sg13g2_fill_1 FILLER_7_302 ();
 sg13g2_decap_4 FILLER_7_329 ();
 sg13g2_fill_1 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_8 FILLER_7_403 ();
 sg13g2_decap_8 FILLER_7_410 ();
 sg13g2_decap_8 FILLER_7_417 ();
 sg13g2_decap_4 FILLER_7_424 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_4 FILLER_8_133 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_160 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_1 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_193 ();
 sg13g2_decap_4 FILLER_8_204 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_228 ();
 sg13g2_fill_1 FILLER_8_249 ();
 sg13g2_fill_1 FILLER_8_255 ();
 sg13g2_fill_2 FILLER_8_261 ();
 sg13g2_fill_2 FILLER_8_268 ();
 sg13g2_fill_1 FILLER_8_294 ();
 sg13g2_fill_2 FILLER_8_300 ();
 sg13g2_fill_2 FILLER_8_319 ();
 sg13g2_fill_2 FILLER_8_338 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_8_409 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_4 FILLER_9_126 ();
 sg13g2_fill_2 FILLER_9_151 ();
 sg13g2_fill_1 FILLER_9_183 ();
 sg13g2_fill_2 FILLER_9_270 ();
 sg13g2_fill_2 FILLER_9_292 ();
 sg13g2_fill_1 FILLER_9_294 ();
 sg13g2_fill_2 FILLER_9_300 ();
 sg13g2_fill_2 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_309 ();
 sg13g2_fill_2 FILLER_9_315 ();
 sg13g2_fill_1 FILLER_9_317 ();
 sg13g2_fill_2 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_decap_8 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_9_415 ();
 sg13g2_decap_8 FILLER_9_422 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_4 FILLER_10_112 ();
 sg13g2_fill_1 FILLER_10_116 ();
 sg13g2_fill_1 FILLER_10_181 ();
 sg13g2_fill_1 FILLER_10_197 ();
 sg13g2_fill_2 FILLER_10_224 ();
 sg13g2_fill_2 FILLER_10_237 ();
 sg13g2_fill_2 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_fill_1 FILLER_10_285 ();
 sg13g2_fill_2 FILLER_10_303 ();
 sg13g2_fill_2 FILLER_10_309 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_fill_1 FILLER_10_339 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_decap_8 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_144 ();
 sg13g2_fill_2 FILLER_11_165 ();
 sg13g2_fill_2 FILLER_11_189 ();
 sg13g2_fill_1 FILLER_11_201 ();
 sg13g2_decap_4 FILLER_11_226 ();
 sg13g2_decap_4 FILLER_11_234 ();
 sg13g2_fill_1 FILLER_11_238 ();
 sg13g2_fill_1 FILLER_11_245 ();
 sg13g2_decap_4 FILLER_11_263 ();
 sg13g2_fill_1 FILLER_11_267 ();
 sg13g2_fill_1 FILLER_11_277 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_decap_4 FILLER_11_337 ();
 sg13g2_fill_2 FILLER_11_341 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_8 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_11_412 ();
 sg13g2_decap_8 FILLER_11_419 ();
 sg13g2_decap_4 FILLER_11_426 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_4 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_181 ();
 sg13g2_decap_4 FILLER_12_188 ();
 sg13g2_fill_2 FILLER_12_192 ();
 sg13g2_fill_1 FILLER_12_197 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_252 ();
 sg13g2_fill_1 FILLER_12_263 ();
 sg13g2_decap_4 FILLER_12_341 ();
 sg13g2_fill_2 FILLER_12_345 ();
 sg13g2_fill_1 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_366 ();
 sg13g2_decap_4 FILLER_12_373 ();
 sg13g2_fill_2 FILLER_12_377 ();
 sg13g2_fill_2 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_12_409 ();
 sg13g2_decap_8 FILLER_12_416 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_fill_1 FILLER_13_133 ();
 sg13g2_fill_2 FILLER_13_142 ();
 sg13g2_fill_2 FILLER_13_158 ();
 sg13g2_fill_1 FILLER_13_160 ();
 sg13g2_decap_4 FILLER_13_183 ();
 sg13g2_fill_2 FILLER_13_191 ();
 sg13g2_fill_1 FILLER_13_193 ();
 sg13g2_fill_2 FILLER_13_197 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_226 ();
 sg13g2_fill_1 FILLER_13_233 ();
 sg13g2_fill_2 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_335 ();
 sg13g2_fill_2 FILLER_13_363 ();
 sg13g2_fill_1 FILLER_13_374 ();
 sg13g2_fill_2 FILLER_13_397 ();
 sg13g2_fill_1 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_8 FILLER_13_419 ();
 sg13g2_decap_4 FILLER_13_426 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_4 FILLER_14_123 ();
 sg13g2_fill_1 FILLER_14_127 ();
 sg13g2_fill_2 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_fill_1 FILLER_14_356 ();
 sg13g2_fill_2 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_409 ();
 sg13g2_decap_8 FILLER_14_416 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_154 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_fill_1 FILLER_15_195 ();
 sg13g2_fill_2 FILLER_15_200 ();
 sg13g2_decap_4 FILLER_15_224 ();
 sg13g2_decap_4 FILLER_15_233 ();
 sg13g2_fill_1 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_fill_2 FILLER_15_260 ();
 sg13g2_fill_1 FILLER_15_267 ();
 sg13g2_fill_1 FILLER_15_271 ();
 sg13g2_fill_1 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_285 ();
 sg13g2_decap_8 FILLER_15_292 ();
 sg13g2_fill_1 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_fill_2 FILLER_15_375 ();
 sg13g2_fill_1 FILLER_15_382 ();
 sg13g2_fill_1 FILLER_15_396 ();
 sg13g2_decap_8 FILLER_15_423 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_decap_4 FILLER_16_144 ();
 sg13g2_fill_2 FILLER_16_148 ();
 sg13g2_fill_1 FILLER_16_160 ();
 sg13g2_fill_2 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_203 ();
 sg13g2_decap_4 FILLER_16_253 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_decap_4 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_4 FILLER_16_356 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_fill_2 FILLER_16_404 ();
 sg13g2_decap_8 FILLER_16_410 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_4 FILLER_16_424 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_decap_4 FILLER_17_211 ();
 sg13g2_decap_4 FILLER_17_219 ();
 sg13g2_decap_4 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_328 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_355 ();
 sg13g2_decap_4 FILLER_17_362 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_fill_2 FILLER_17_396 ();
 sg13g2_fill_1 FILLER_17_398 ();
 sg13g2_decap_8 FILLER_17_416 ();
 sg13g2_decap_8 FILLER_17_423 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_141 ();
 sg13g2_fill_2 FILLER_18_151 ();
 sg13g2_decap_4 FILLER_18_160 ();
 sg13g2_fill_2 FILLER_18_164 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_190 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_204 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_decap_4 FILLER_18_212 ();
 sg13g2_fill_2 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_226 ();
 sg13g2_decap_4 FILLER_18_263 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_299 ();
 sg13g2_fill_1 FILLER_18_301 ();
 sg13g2_decap_4 FILLER_18_305 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_372 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_fill_2 FILLER_18_383 ();
 sg13g2_fill_1 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_18_411 ();
 sg13g2_decap_8 FILLER_18_418 ();
 sg13g2_decap_4 FILLER_18_425 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_4 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_143 ();
 sg13g2_fill_1 FILLER_19_148 ();
 sg13g2_fill_1 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_160 ();
 sg13g2_decap_8 FILLER_19_167 ();
 sg13g2_decap_4 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_178 ();
 sg13g2_decap_4 FILLER_19_185 ();
 sg13g2_fill_1 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_4 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_fill_1 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_1 FILLER_19_245 ();
 sg13g2_fill_1 FILLER_19_256 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_fill_1 FILLER_19_269 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_319 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_fill_1 FILLER_19_331 ();
 sg13g2_fill_2 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_349 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_377 ();
 sg13g2_fill_1 FILLER_19_379 ();
 sg13g2_decap_8 FILLER_19_404 ();
 sg13g2_decap_8 FILLER_19_411 ();
 sg13g2_decap_8 FILLER_19_418 ();
 sg13g2_decap_4 FILLER_19_425 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_4 FILLER_20_98 ();
 sg13g2_fill_1 FILLER_20_102 ();
 sg13g2_fill_1 FILLER_20_138 ();
 sg13g2_fill_1 FILLER_20_167 ();
 sg13g2_fill_2 FILLER_20_185 ();
 sg13g2_fill_2 FILLER_20_191 ();
 sg13g2_fill_1 FILLER_20_218 ();
 sg13g2_decap_8 FILLER_20_248 ();
 sg13g2_decap_8 FILLER_20_255 ();
 sg13g2_fill_2 FILLER_20_262 ();
 sg13g2_fill_1 FILLER_20_276 ();
 sg13g2_fill_2 FILLER_20_289 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_fill_1 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_347 ();
 sg13g2_fill_2 FILLER_20_366 ();
 sg13g2_fill_1 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_fill_2 FILLER_20_386 ();
 sg13g2_fill_1 FILLER_20_391 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_decap_4 FILLER_20_425 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_4 FILLER_21_84 ();
 sg13g2_fill_2 FILLER_21_88 ();
 sg13g2_fill_1 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_121 ();
 sg13g2_fill_2 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_fill_2 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_247 ();
 sg13g2_fill_1 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_284 ();
 sg13g2_decap_4 FILLER_21_290 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_2 FILLER_21_315 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_decap_4 FILLER_21_359 ();
 sg13g2_fill_1 FILLER_21_363 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_4 FILLER_21_393 ();
 sg13g2_fill_2 FILLER_21_397 ();
 sg13g2_decap_8 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_416 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_103 ();
 sg13g2_fill_2 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_114 ();
 sg13g2_fill_2 FILLER_22_165 ();
 sg13g2_fill_2 FILLER_22_170 ();
 sg13g2_fill_1 FILLER_22_172 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_fill_2 FILLER_22_249 ();
 sg13g2_fill_2 FILLER_22_344 ();
 sg13g2_fill_1 FILLER_22_352 ();
 sg13g2_fill_2 FILLER_22_370 ();
 sg13g2_fill_1 FILLER_22_372 ();
 sg13g2_fill_1 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_389 ();
 sg13g2_fill_2 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_4 FILLER_22_424 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_110 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_147 ();
 sg13g2_decap_4 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_277 ();
 sg13g2_decap_4 FILLER_23_282 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_fill_1 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_421 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_142 ();
 sg13g2_fill_1 FILLER_24_144 ();
 sg13g2_fill_1 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_decap_4 FILLER_24_223 ();
 sg13g2_fill_2 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_234 ();
 sg13g2_fill_2 FILLER_24_241 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_262 ();
 sg13g2_decap_4 FILLER_24_282 ();
 sg13g2_fill_2 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_4 FILLER_24_424 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_4 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_fill_2 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_131 ();
 sg13g2_decap_4 FILLER_25_177 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_decap_4 FILLER_25_214 ();
 sg13g2_fill_2 FILLER_25_218 ();
 sg13g2_decap_4 FILLER_25_228 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_fill_1 FILLER_25_273 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_fill_1 FILLER_25_294 ();
 sg13g2_decap_4 FILLER_25_299 ();
 sg13g2_decap_4 FILLER_25_308 ();
 sg13g2_fill_1 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_fill_1 FILLER_25_367 ();
 sg13g2_fill_2 FILLER_25_393 ();
 sg13g2_fill_2 FILLER_25_410 ();
 sg13g2_fill_1 FILLER_25_412 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_4 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_105 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_fill_1 FILLER_26_120 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_181 ();
 sg13g2_decap_4 FILLER_26_208 ();
 sg13g2_fill_1 FILLER_26_212 ();
 sg13g2_fill_1 FILLER_26_230 ();
 sg13g2_decap_4 FILLER_26_243 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_4 FILLER_27_113 ();
 sg13g2_fill_2 FILLER_27_131 ();
 sg13g2_fill_1 FILLER_27_133 ();
 sg13g2_fill_1 FILLER_27_138 ();
 sg13g2_decap_4 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_154 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_2 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_195 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_275 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_fill_1 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_329 ();
 sg13g2_fill_2 FILLER_27_340 ();
 sg13g2_fill_1 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_353 ();
 sg13g2_fill_2 FILLER_27_360 ();
 sg13g2_fill_2 FILLER_27_372 ();
 sg13g2_fill_1 FILLER_27_374 ();
 sg13g2_fill_2 FILLER_27_385 ();
 sg13g2_fill_1 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_392 ();
 sg13g2_fill_1 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_412 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_98 ();
 sg13g2_fill_2 FILLER_28_102 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_fill_1 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_180 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_fill_1 FILLER_28_233 ();
 sg13g2_decap_8 FILLER_28_261 ();
 sg13g2_decap_4 FILLER_28_273 ();
 sg13g2_decap_4 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_decap_4 FILLER_28_332 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_341 ();
 sg13g2_fill_2 FILLER_28_355 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_fill_2 FILLER_28_372 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_fill_1 FILLER_28_389 ();
 sg13g2_decap_8 FILLER_28_412 ();
 sg13g2_decap_8 FILLER_28_419 ();
 sg13g2_decap_4 FILLER_28_426 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_4 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_174 ();
 sg13g2_fill_1 FILLER_29_181 ();
 sg13g2_decap_4 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_decap_4 FILLER_29_232 ();
 sg13g2_decap_4 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_252 ();
 sg13g2_decap_4 FILLER_29_280 ();
 sg13g2_fill_2 FILLER_29_284 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_299 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_1 FILLER_29_384 ();
 sg13g2_decap_4 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_29_398 ();
 sg13g2_decap_8 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_29_412 ();
 sg13g2_decap_8 FILLER_29_419 ();
 sg13g2_decap_4 FILLER_29_426 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_131 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_184 ();
 sg13g2_fill_1 FILLER_30_200 ();
 sg13g2_fill_1 FILLER_30_227 ();
 sg13g2_decap_8 FILLER_30_258 ();
 sg13g2_decap_8 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_272 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_344 ();
 sg13g2_decap_4 FILLER_30_359 ();
 sg13g2_fill_1 FILLER_30_371 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_4 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_decap_4 FILLER_31_134 ();
 sg13g2_fill_2 FILLER_31_138 ();
 sg13g2_fill_2 FILLER_31_157 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_fill_2 FILLER_31_170 ();
 sg13g2_fill_2 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_196 ();
 sg13g2_fill_2 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_fill_2 FILLER_31_222 ();
 sg13g2_decap_4 FILLER_31_234 ();
 sg13g2_fill_1 FILLER_31_238 ();
 sg13g2_decap_4 FILLER_31_256 ();
 sg13g2_fill_2 FILLER_31_260 ();
 sg13g2_decap_4 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_358 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_decap_8 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_4 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_111 ();
 sg13g2_fill_1 FILLER_32_113 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_4 FILLER_32_133 ();
 sg13g2_fill_2 FILLER_32_137 ();
 sg13g2_decap_4 FILLER_32_146 ();
 sg13g2_fill_1 FILLER_32_150 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_262 ();
 sg13g2_fill_1 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_346 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_fill_1 FILLER_32_365 ();
 sg13g2_fill_1 FILLER_32_372 ();
 sg13g2_fill_1 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_32_400 ();
 sg13g2_decap_8 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_32_414 ();
 sg13g2_decap_8 FILLER_32_421 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_81 ();
 sg13g2_fill_2 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_101 ();
 sg13g2_decap_4 FILLER_33_107 ();
 sg13g2_fill_2 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_138 ();
 sg13g2_fill_1 FILLER_33_164 ();
 sg13g2_fill_2 FILLER_33_179 ();
 sg13g2_fill_1 FILLER_33_181 ();
 sg13g2_fill_1 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_fill_1 FILLER_33_222 ();
 sg13g2_fill_1 FILLER_33_228 ();
 sg13g2_fill_1 FILLER_33_233 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_fill_2 FILLER_33_318 ();
 sg13g2_fill_1 FILLER_33_342 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_decap_4 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_396 ();
 sg13g2_fill_1 FILLER_33_398 ();
 sg13g2_decap_8 FILLER_33_409 ();
 sg13g2_decap_8 FILLER_33_416 ();
 sg13g2_decap_8 FILLER_33_423 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_108 ();
 sg13g2_fill_1 FILLER_34_193 ();
 sg13g2_fill_2 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_226 ();
 sg13g2_decap_8 FILLER_34_236 ();
 sg13g2_decap_8 FILLER_34_243 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_decap_4 FILLER_34_275 ();
 sg13g2_fill_2 FILLER_34_288 ();
 sg13g2_decap_4 FILLER_34_301 ();
 sg13g2_fill_1 FILLER_34_309 ();
 sg13g2_fill_2 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_fill_2 FILLER_34_356 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_fill_1 FILLER_34_388 ();
 sg13g2_fill_2 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_411 ();
 sg13g2_decap_8 FILLER_34_418 ();
 sg13g2_decap_4 FILLER_34_425 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_4 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_128 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_2 FILLER_35_159 ();
 sg13g2_fill_1 FILLER_35_161 ();
 sg13g2_fill_2 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_fill_1 FILLER_35_267 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_fill_1 FILLER_35_315 ();
 sg13g2_decap_4 FILLER_35_351 ();
 sg13g2_fill_2 FILLER_35_355 ();
 sg13g2_fill_2 FILLER_35_362 ();
 sg13g2_fill_1 FILLER_35_364 ();
 sg13g2_decap_4 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_404 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_4 FILLER_36_84 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_130 ();
 sg13g2_fill_1 FILLER_36_136 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_fill_1 FILLER_36_161 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_2 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_191 ();
 sg13g2_fill_1 FILLER_36_193 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_245 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_fill_1 FILLER_36_257 ();
 sg13g2_fill_1 FILLER_36_300 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_345 ();
 sg13g2_fill_1 FILLER_36_347 ();
 sg13g2_fill_1 FILLER_36_370 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_fill_1 FILLER_36_396 ();
 sg13g2_fill_2 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_419 ();
 sg13g2_decap_4 FILLER_36_426 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_fill_2 FILLER_37_104 ();
 sg13g2_fill_1 FILLER_37_106 ();
 sg13g2_decap_4 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_fill_2 FILLER_37_144 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_162 ();
 sg13g2_fill_2 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_250 ();
 sg13g2_fill_1 FILLER_37_261 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_fill_1 FILLER_37_296 ();
 sg13g2_fill_2 FILLER_37_312 ();
 sg13g2_fill_1 FILLER_37_314 ();
 sg13g2_fill_1 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_fill_2 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_103 ();
 sg13g2_decap_4 FILLER_38_110 ();
 sg13g2_fill_2 FILLER_38_114 ();
 sg13g2_fill_1 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_186 ();
 sg13g2_fill_2 FILLER_38_202 ();
 sg13g2_fill_2 FILLER_38_257 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_fill_2 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_289 ();
 sg13g2_decap_4 FILLER_38_329 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_4 FILLER_38_417 ();
 sg13g2_fill_1 FILLER_38_421 ();
 sg13g2_decap_4 FILLER_38_426 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_4 FILLER_39_98 ();
 sg13g2_fill_1 FILLER_39_102 ();
 sg13g2_fill_2 FILLER_39_124 ();
 sg13g2_fill_2 FILLER_39_132 ();
 sg13g2_fill_1 FILLER_39_134 ();
 sg13g2_decap_4 FILLER_39_140 ();
 sg13g2_fill_1 FILLER_39_144 ();
 sg13g2_decap_4 FILLER_39_178 ();
 sg13g2_fill_2 FILLER_39_182 ();
 sg13g2_fill_1 FILLER_39_213 ();
 sg13g2_fill_1 FILLER_39_227 ();
 sg13g2_fill_1 FILLER_39_235 ();
 sg13g2_fill_1 FILLER_39_239 ();
 sg13g2_fill_1 FILLER_39_248 ();
 sg13g2_fill_1 FILLER_39_254 ();
 sg13g2_fill_2 FILLER_39_272 ();
 sg13g2_fill_2 FILLER_39_279 ();
 sg13g2_fill_1 FILLER_39_281 ();
 sg13g2_fill_2 FILLER_39_287 ();
 sg13g2_fill_1 FILLER_39_289 ();
 sg13g2_fill_2 FILLER_39_307 ();
 sg13g2_decap_4 FILLER_39_314 ();
 sg13g2_fill_2 FILLER_39_328 ();
 sg13g2_decap_4 FILLER_39_334 ();
 sg13g2_fill_2 FILLER_39_363 ();
 sg13g2_fill_2 FILLER_39_375 ();
 sg13g2_decap_4 FILLER_39_381 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_4 FILLER_40_84 ();
 sg13g2_fill_2 FILLER_40_88 ();
 sg13g2_decap_8 FILLER_40_136 ();
 sg13g2_fill_2 FILLER_40_143 ();
 sg13g2_fill_1 FILLER_40_145 ();
 sg13g2_decap_8 FILLER_40_180 ();
 sg13g2_fill_1 FILLER_40_187 ();
 sg13g2_decap_8 FILLER_40_192 ();
 sg13g2_decap_4 FILLER_40_199 ();
 sg13g2_fill_2 FILLER_40_203 ();
 sg13g2_decap_4 FILLER_40_216 ();
 sg13g2_fill_1 FILLER_40_220 ();
 sg13g2_fill_1 FILLER_40_224 ();
 sg13g2_fill_1 FILLER_40_229 ();
 sg13g2_fill_1 FILLER_40_234 ();
 sg13g2_fill_1 FILLER_40_239 ();
 sg13g2_fill_1 FILLER_40_251 ();
 sg13g2_decap_4 FILLER_40_257 ();
 sg13g2_fill_1 FILLER_40_261 ();
 sg13g2_fill_1 FILLER_40_279 ();
 sg13g2_decap_4 FILLER_40_306 ();
 sg13g2_fill_1 FILLER_40_310 ();
 sg13g2_fill_2 FILLER_40_321 ();
 sg13g2_decap_4 FILLER_40_349 ();
 sg13g2_decap_8 FILLER_40_358 ();
 sg13g2_fill_2 FILLER_40_365 ();
 sg13g2_decap_4 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_381 ();
 sg13g2_decap_4 FILLER_40_388 ();
 sg13g2_fill_2 FILLER_40_392 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_4 FILLER_41_77 ();
 sg13g2_fill_2 FILLER_41_81 ();
 sg13g2_decap_4 FILLER_41_122 ();
 sg13g2_fill_2 FILLER_41_141 ();
 sg13g2_fill_1 FILLER_41_143 ();
 sg13g2_decap_4 FILLER_41_148 ();
 sg13g2_fill_1 FILLER_41_152 ();
 sg13g2_fill_2 FILLER_41_168 ();
 sg13g2_fill_2 FILLER_41_175 ();
 sg13g2_fill_1 FILLER_41_177 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_fill_2 FILLER_41_188 ();
 sg13g2_fill_1 FILLER_41_190 ();
 sg13g2_fill_2 FILLER_41_219 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_decap_8 FILLER_41_226 ();
 sg13g2_decap_8 FILLER_41_233 ();
 sg13g2_decap_4 FILLER_41_240 ();
 sg13g2_fill_1 FILLER_41_244 ();
 sg13g2_fill_1 FILLER_41_249 ();
 sg13g2_fill_1 FILLER_41_253 ();
 sg13g2_decap_8 FILLER_41_258 ();
 sg13g2_fill_2 FILLER_41_265 ();
 sg13g2_fill_2 FILLER_41_272 ();
 sg13g2_fill_1 FILLER_41_274 ();
 sg13g2_decap_4 FILLER_41_280 ();
 sg13g2_fill_2 FILLER_41_284 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_4 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_fill_2 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_345 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_decap_4 FILLER_41_356 ();
 sg13g2_fill_2 FILLER_41_360 ();
 sg13g2_fill_2 FILLER_41_422 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_4 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_92 ();
 sg13g2_decap_8 FILLER_42_99 ();
 sg13g2_fill_2 FILLER_42_106 ();
 sg13g2_fill_1 FILLER_42_108 ();
 sg13g2_fill_2 FILLER_42_131 ();
 sg13g2_fill_1 FILLER_42_147 ();
 sg13g2_fill_1 FILLER_42_155 ();
 sg13g2_fill_1 FILLER_42_161 ();
 sg13g2_fill_1 FILLER_42_172 ();
 sg13g2_fill_1 FILLER_42_178 ();
 sg13g2_fill_1 FILLER_42_186 ();
 sg13g2_fill_1 FILLER_42_220 ();
 sg13g2_decap_4 FILLER_42_229 ();
 sg13g2_decap_8 FILLER_42_289 ();
 sg13g2_fill_2 FILLER_42_296 ();
 sg13g2_fill_1 FILLER_42_298 ();
 sg13g2_decap_4 FILLER_42_311 ();
 sg13g2_fill_2 FILLER_42_325 ();
 sg13g2_decap_4 FILLER_42_332 ();
 sg13g2_fill_2 FILLER_42_360 ();
 sg13g2_fill_2 FILLER_42_368 ();
 sg13g2_decap_4 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_4 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_88 ();
 sg13g2_fill_1 FILLER_43_112 ();
 sg13g2_fill_2 FILLER_43_149 ();
 sg13g2_fill_1 FILLER_43_151 ();
 sg13g2_fill_2 FILLER_43_156 ();
 sg13g2_fill_1 FILLER_43_162 ();
 sg13g2_fill_1 FILLER_43_170 ();
 sg13g2_fill_2 FILLER_43_181 ();
 sg13g2_fill_1 FILLER_43_193 ();
 sg13g2_fill_2 FILLER_43_202 ();
 sg13g2_fill_1 FILLER_43_208 ();
 sg13g2_fill_2 FILLER_43_238 ();
 sg13g2_decap_4 FILLER_43_282 ();
 sg13g2_fill_2 FILLER_43_286 ();
 sg13g2_fill_2 FILLER_43_309 ();
 sg13g2_fill_2 FILLER_43_341 ();
 sg13g2_fill_1 FILLER_43_357 ();
 sg13g2_fill_1 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_374 ();
 sg13g2_fill_1 FILLER_43_380 ();
 sg13g2_fill_1 FILLER_43_391 ();
 sg13g2_fill_1 FILLER_43_402 ();
 sg13g2_fill_1 FILLER_43_411 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_fill_1 FILLER_44_115 ();
 sg13g2_fill_2 FILLER_44_143 ();
 sg13g2_fill_2 FILLER_44_163 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_decap_4 FILLER_44_238 ();
 sg13g2_fill_2 FILLER_44_242 ();
 sg13g2_fill_1 FILLER_44_357 ();
 sg13g2_fill_1 FILLER_44_362 ();
 sg13g2_fill_1 FILLER_44_413 ();
 sg13g2_fill_2 FILLER_44_427 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_4 FILLER_45_91 ();
 sg13g2_fill_2 FILLER_45_95 ();
 sg13g2_fill_1 FILLER_45_102 ();
 sg13g2_fill_1 FILLER_45_116 ();
 sg13g2_decap_4 FILLER_45_136 ();
 sg13g2_fill_2 FILLER_45_140 ();
 sg13g2_fill_2 FILLER_45_152 ();
 sg13g2_fill_1 FILLER_45_160 ();
 sg13g2_fill_2 FILLER_45_164 ();
 sg13g2_fill_2 FILLER_45_186 ();
 sg13g2_fill_1 FILLER_45_188 ();
 sg13g2_fill_1 FILLER_45_197 ();
 sg13g2_fill_1 FILLER_45_220 ();
 sg13g2_decap_4 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_259 ();
 sg13g2_fill_2 FILLER_45_265 ();
 sg13g2_fill_1 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_320 ();
 sg13g2_fill_1 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_358 ();
 sg13g2_fill_2 FILLER_45_365 ();
 sg13g2_fill_1 FILLER_45_367 ();
 sg13g2_fill_1 FILLER_45_396 ();
 sg13g2_decap_4 FILLER_45_406 ();
 sg13g2_fill_2 FILLER_45_410 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_fill_2 FILLER_46_84 ();
 sg13g2_decap_4 FILLER_46_103 ();
 sg13g2_fill_1 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_206 ();
 sg13g2_fill_2 FILLER_46_222 ();
 sg13g2_decap_8 FILLER_46_241 ();
 sg13g2_decap_8 FILLER_46_248 ();
 sg13g2_decap_4 FILLER_46_296 ();
 sg13g2_fill_1 FILLER_46_304 ();
 sg13g2_fill_1 FILLER_46_325 ();
 sg13g2_fill_1 FILLER_46_336 ();
 sg13g2_decap_4 FILLER_46_342 ();
 sg13g2_fill_2 FILLER_46_346 ();
 sg13g2_decap_4 FILLER_46_358 ();
 sg13g2_fill_1 FILLER_46_362 ();
 sg13g2_decap_8 FILLER_46_368 ();
 sg13g2_decap_4 FILLER_46_375 ();
 sg13g2_fill_1 FILLER_46_379 ();
 sg13g2_fill_1 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_fill_1 FILLER_46_406 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_fill_1 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_136 ();
 sg13g2_fill_1 FILLER_47_148 ();
 sg13g2_fill_1 FILLER_47_153 ();
 sg13g2_fill_1 FILLER_47_159 ();
 sg13g2_fill_1 FILLER_47_165 ();
 sg13g2_fill_1 FILLER_47_176 ();
 sg13g2_fill_1 FILLER_47_181 ();
 sg13g2_fill_1 FILLER_47_199 ();
 sg13g2_fill_2 FILLER_47_222 ();
 sg13g2_fill_1 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_242 ();
 sg13g2_decap_8 FILLER_47_249 ();
 sg13g2_decap_8 FILLER_47_256 ();
 sg13g2_decap_4 FILLER_47_263 ();
 sg13g2_fill_1 FILLER_47_267 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_fill_1 FILLER_47_284 ();
 sg13g2_fill_2 FILLER_47_347 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_4 FILLER_47_378 ();
 sg13g2_decap_4 FILLER_47_396 ();
 sg13g2_decap_4 FILLER_47_424 ();
 sg13g2_fill_2 FILLER_47_428 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_129 ();
 sg13g2_fill_2 FILLER_48_136 ();
 sg13g2_fill_1 FILLER_48_138 ();
 sg13g2_decap_4 FILLER_48_193 ();
 sg13g2_fill_2 FILLER_48_201 ();
 sg13g2_fill_2 FILLER_48_207 ();
 sg13g2_fill_1 FILLER_48_209 ();
 sg13g2_decap_8 FILLER_48_227 ();
 sg13g2_decap_4 FILLER_48_234 ();
 sg13g2_fill_1 FILLER_48_238 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_2 FILLER_48_271 ();
 sg13g2_fill_2 FILLER_48_306 ();
 sg13g2_fill_2 FILLER_48_319 ();
 sg13g2_fill_1 FILLER_48_321 ();
 sg13g2_fill_1 FILLER_48_331 ();
 sg13g2_decap_4 FILLER_48_376 ();
 sg13g2_fill_2 FILLER_48_380 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_84 ();
 sg13g2_fill_1 FILLER_49_115 ();
 sg13g2_fill_2 FILLER_49_132 ();
 sg13g2_fill_1 FILLER_49_134 ();
 sg13g2_fill_2 FILLER_49_152 ();
 sg13g2_decap_4 FILLER_49_159 ();
 sg13g2_decap_8 FILLER_49_173 ();
 sg13g2_fill_1 FILLER_49_206 ();
 sg13g2_fill_2 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_230 ();
 sg13g2_decap_8 FILLER_49_237 ();
 sg13g2_fill_1 FILLER_49_244 ();
 sg13g2_decap_4 FILLER_49_250 ();
 sg13g2_fill_2 FILLER_49_254 ();
 sg13g2_fill_1 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_265 ();
 sg13g2_fill_1 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_303 ();
 sg13g2_fill_2 FILLER_49_310 ();
 sg13g2_fill_1 FILLER_49_312 ();
 sg13g2_fill_2 FILLER_49_336 ();
 sg13g2_fill_1 FILLER_49_338 ();
 sg13g2_fill_2 FILLER_49_361 ();
 sg13g2_fill_1 FILLER_49_363 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_4 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_77 ();
 sg13g2_fill_1 FILLER_50_79 ();
 sg13g2_fill_2 FILLER_50_106 ();
 sg13g2_fill_1 FILLER_50_108 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_fill_2 FILLER_50_147 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_decap_8 FILLER_50_158 ();
 sg13g2_decap_8 FILLER_50_165 ();
 sg13g2_decap_8 FILLER_50_172 ();
 sg13g2_decap_8 FILLER_50_179 ();
 sg13g2_fill_2 FILLER_50_186 ();
 sg13g2_fill_1 FILLER_50_188 ();
 sg13g2_decap_8 FILLER_50_193 ();
 sg13g2_fill_2 FILLER_50_200 ();
 sg13g2_fill_1 FILLER_50_202 ();
 sg13g2_fill_1 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_238 ();
 sg13g2_fill_1 FILLER_50_244 ();
 sg13g2_fill_1 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_286 ();
 sg13g2_fill_1 FILLER_50_288 ();
 sg13g2_fill_1 FILLER_50_295 ();
 sg13g2_fill_2 FILLER_50_317 ();
 sg13g2_fill_2 FILLER_50_323 ();
 sg13g2_fill_1 FILLER_50_325 ();
 sg13g2_fill_1 FILLER_50_338 ();
 sg13g2_fill_2 FILLER_50_356 ();
 sg13g2_fill_1 FILLER_50_400 ();
 sg13g2_fill_2 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_fill_2 FILLER_51_84 ();
 sg13g2_fill_1 FILLER_51_86 ();
 sg13g2_fill_1 FILLER_51_98 ();
 sg13g2_fill_1 FILLER_51_103 ();
 sg13g2_fill_1 FILLER_51_117 ();
 sg13g2_decap_8 FILLER_51_128 ();
 sg13g2_decap_4 FILLER_51_139 ();
 sg13g2_fill_1 FILLER_51_177 ();
 sg13g2_decap_8 FILLER_51_183 ();
 sg13g2_fill_2 FILLER_51_190 ();
 sg13g2_fill_1 FILLER_51_192 ();
 sg13g2_fill_1 FILLER_51_217 ();
 sg13g2_fill_1 FILLER_51_269 ();
 sg13g2_fill_2 FILLER_51_312 ();
 sg13g2_decap_4 FILLER_51_358 ();
 sg13g2_fill_2 FILLER_51_362 ();
 sg13g2_fill_1 FILLER_51_370 ();
 sg13g2_fill_1 FILLER_51_402 ();
 sg13g2_fill_1 FILLER_51_407 ();
 sg13g2_fill_1 FILLER_51_429 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_98 ();
 sg13g2_fill_1 FILLER_52_100 ();
 sg13g2_fill_2 FILLER_52_106 ();
 sg13g2_fill_1 FILLER_52_113 ();
 sg13g2_decap_8 FILLER_52_121 ();
 sg13g2_fill_2 FILLER_52_128 ();
 sg13g2_fill_1 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_151 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_1 FILLER_52_187 ();
 sg13g2_fill_2 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_200 ();
 sg13g2_fill_1 FILLER_52_223 ();
 sg13g2_fill_2 FILLER_52_229 ();
 sg13g2_fill_2 FILLER_52_297 ();
 sg13g2_fill_2 FILLER_52_309 ();
 sg13g2_fill_1 FILLER_52_311 ();
 sg13g2_fill_2 FILLER_52_340 ();
 sg13g2_fill_1 FILLER_52_370 ();
 sg13g2_decap_4 FILLER_52_387 ();
 sg13g2_decap_4 FILLER_52_426 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_fill_1 FILLER_53_120 ();
 sg13g2_fill_2 FILLER_53_162 ();
 sg13g2_fill_1 FILLER_53_164 ();
 sg13g2_fill_2 FILLER_53_239 ();
 sg13g2_fill_2 FILLER_53_246 ();
 sg13g2_fill_2 FILLER_53_253 ();
 sg13g2_decap_8 FILLER_53_260 ();
 sg13g2_fill_1 FILLER_53_267 ();
 sg13g2_decap_4 FILLER_53_278 ();
 sg13g2_fill_2 FILLER_53_282 ();
 sg13g2_decap_4 FILLER_53_288 ();
 sg13g2_fill_1 FILLER_53_324 ();
 sg13g2_fill_2 FILLER_53_351 ();
 sg13g2_fill_1 FILLER_53_353 ();
 sg13g2_decap_4 FILLER_53_358 ();
 sg13g2_decap_4 FILLER_53_389 ();
 sg13g2_fill_1 FILLER_53_393 ();
 sg13g2_decap_8 FILLER_53_402 ();
 sg13g2_fill_2 FILLER_53_409 ();
 sg13g2_fill_1 FILLER_53_411 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_84 ();
 sg13g2_fill_1 FILLER_54_86 ();
 sg13g2_fill_2 FILLER_54_133 ();
 sg13g2_fill_1 FILLER_54_135 ();
 sg13g2_fill_1 FILLER_54_147 ();
 sg13g2_fill_2 FILLER_54_179 ();
 sg13g2_fill_1 FILLER_54_181 ();
 sg13g2_fill_2 FILLER_54_218 ();
 sg13g2_fill_1 FILLER_54_225 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_decap_8 FILLER_54_239 ();
 sg13g2_decap_8 FILLER_54_246 ();
 sg13g2_decap_4 FILLER_54_253 ();
 sg13g2_fill_1 FILLER_54_257 ();
 sg13g2_decap_8 FILLER_54_267 ();
 sg13g2_fill_2 FILLER_54_274 ();
 sg13g2_decap_4 FILLER_54_287 ();
 sg13g2_fill_1 FILLER_54_314 ();
 sg13g2_fill_1 FILLER_54_331 ();
 sg13g2_decap_8 FILLER_54_357 ();
 sg13g2_fill_2 FILLER_54_364 ();
 sg13g2_fill_1 FILLER_54_366 ();
 sg13g2_fill_2 FILLER_54_386 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_4 FILLER_55_84 ();
 sg13g2_fill_2 FILLER_55_88 ();
 sg13g2_fill_2 FILLER_55_131 ();
 sg13g2_fill_1 FILLER_55_133 ();
 sg13g2_decap_4 FILLER_55_143 ();
 sg13g2_fill_1 FILLER_55_147 ();
 sg13g2_fill_2 FILLER_55_179 ();
 sg13g2_fill_1 FILLER_55_202 ();
 sg13g2_decap_4 FILLER_55_239 ();
 sg13g2_decap_8 FILLER_55_247 ();
 sg13g2_fill_2 FILLER_55_271 ();
 sg13g2_fill_1 FILLER_55_273 ();
 sg13g2_fill_2 FILLER_55_287 ();
 sg13g2_fill_1 FILLER_55_310 ();
 sg13g2_fill_1 FILLER_55_338 ();
 sg13g2_fill_1 FILLER_55_355 ();
 sg13g2_fill_1 FILLER_55_366 ();
 sg13g2_fill_1 FILLER_55_371 ();
 sg13g2_fill_1 FILLER_55_382 ();
 sg13g2_fill_1 FILLER_55_387 ();
 sg13g2_fill_2 FILLER_55_393 ();
 sg13g2_fill_1 FILLER_55_412 ();
 sg13g2_decap_4 FILLER_55_418 ();
 sg13g2_fill_1 FILLER_55_422 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_4 FILLER_56_105 ();
 sg13g2_fill_2 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_127 ();
 sg13g2_fill_1 FILLER_56_134 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_4 FILLER_56_152 ();
 sg13g2_decap_4 FILLER_56_160 ();
 sg13g2_fill_2 FILLER_56_174 ();
 sg13g2_fill_1 FILLER_56_176 ();
 sg13g2_decap_8 FILLER_56_200 ();
 sg13g2_fill_1 FILLER_56_207 ();
 sg13g2_decap_8 FILLER_56_212 ();
 sg13g2_fill_2 FILLER_56_293 ();
 sg13g2_fill_1 FILLER_56_295 ();
 sg13g2_decap_4 FILLER_56_305 ();
 sg13g2_fill_2 FILLER_56_309 ();
 sg13g2_fill_1 FILLER_56_323 ();
 sg13g2_decap_4 FILLER_56_329 ();
 sg13g2_fill_1 FILLER_56_333 ();
 sg13g2_fill_1 FILLER_56_337 ();
 sg13g2_fill_1 FILLER_56_348 ();
 sg13g2_fill_1 FILLER_56_359 ();
 sg13g2_fill_2 FILLER_56_365 ();
 sg13g2_fill_1 FILLER_56_388 ();
 sg13g2_fill_1 FILLER_56_424 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_4 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_112 ();
 sg13g2_fill_1 FILLER_57_123 ();
 sg13g2_fill_2 FILLER_57_128 ();
 sg13g2_decap_4 FILLER_57_165 ();
 sg13g2_decap_8 FILLER_57_186 ();
 sg13g2_fill_1 FILLER_57_193 ();
 sg13g2_decap_4 FILLER_57_215 ();
 sg13g2_fill_1 FILLER_57_255 ();
 sg13g2_fill_1 FILLER_57_266 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_fill_1 FILLER_57_289 ();
 sg13g2_fill_1 FILLER_57_295 ();
 sg13g2_fill_1 FILLER_57_352 ();
 sg13g2_fill_2 FILLER_57_370 ();
 sg13g2_fill_1 FILLER_57_372 ();
 sg13g2_fill_1 FILLER_57_399 ();
 sg13g2_fill_1 FILLER_57_405 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_4 FILLER_58_77 ();
 sg13g2_fill_1 FILLER_58_81 ();
 sg13g2_fill_1 FILLER_58_113 ();
 sg13g2_fill_2 FILLER_58_170 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_fill_1 FILLER_58_201 ();
 sg13g2_fill_2 FILLER_58_207 ();
 sg13g2_fill_1 FILLER_58_209 ();
 sg13g2_fill_1 FILLER_58_214 ();
 sg13g2_fill_1 FILLER_58_220 ();
 sg13g2_fill_1 FILLER_58_226 ();
 sg13g2_fill_1 FILLER_58_237 ();
 sg13g2_fill_1 FILLER_58_246 ();
 sg13g2_fill_2 FILLER_58_256 ();
 sg13g2_fill_1 FILLER_58_268 ();
 sg13g2_fill_1 FILLER_58_273 ();
 sg13g2_fill_1 FILLER_58_278 ();
 sg13g2_fill_2 FILLER_58_292 ();
 sg13g2_fill_1 FILLER_58_342 ();
 sg13g2_fill_1 FILLER_58_369 ();
 sg13g2_decap_8 FILLER_58_395 ();
 sg13g2_decap_8 FILLER_58_402 ();
 sg13g2_fill_2 FILLER_58_409 ();
 sg13g2_fill_1 FILLER_58_411 ();
 sg13g2_fill_2 FILLER_58_421 ();
 sg13g2_fill_2 FILLER_58_427 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_4 FILLER_59_84 ();
 sg13g2_fill_1 FILLER_59_88 ();
 sg13g2_decap_8 FILLER_59_93 ();
 sg13g2_decap_4 FILLER_59_100 ();
 sg13g2_fill_2 FILLER_59_104 ();
 sg13g2_decap_4 FILLER_59_110 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_142 ();
 sg13g2_fill_1 FILLER_59_148 ();
 sg13g2_fill_1 FILLER_59_162 ();
 sg13g2_fill_2 FILLER_59_167 ();
 sg13g2_fill_1 FILLER_59_169 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_fill_2 FILLER_59_182 ();
 sg13g2_decap_4 FILLER_59_228 ();
 sg13g2_fill_1 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_306 ();
 sg13g2_fill_1 FILLER_59_311 ();
 sg13g2_fill_1 FILLER_59_316 ();
 sg13g2_fill_1 FILLER_59_330 ();
 sg13g2_decap_4 FILLER_59_336 ();
 sg13g2_fill_2 FILLER_59_345 ();
 sg13g2_decap_4 FILLER_59_352 ();
 sg13g2_decap_4 FILLER_59_360 ();
 sg13g2_fill_2 FILLER_59_364 ();
 sg13g2_decap_8 FILLER_59_370 ();
 sg13g2_fill_1 FILLER_59_377 ();
 sg13g2_fill_2 FILLER_59_395 ();
 sg13g2_fill_2 FILLER_59_401 ();
 sg13g2_fill_1 FILLER_59_403 ();
 sg13g2_decap_4 FILLER_59_425 ();
 sg13g2_fill_1 FILLER_59_429 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_4 FILLER_60_91 ();
 sg13g2_fill_1 FILLER_60_124 ();
 sg13g2_fill_1 FILLER_60_137 ();
 sg13g2_fill_1 FILLER_60_142 ();
 sg13g2_fill_2 FILLER_60_151 ();
 sg13g2_fill_2 FILLER_60_162 ();
 sg13g2_fill_2 FILLER_60_178 ();
 sg13g2_decap_8 FILLER_60_183 ();
 sg13g2_fill_2 FILLER_60_190 ();
 sg13g2_fill_2 FILLER_60_251 ();
 sg13g2_fill_1 FILLER_60_258 ();
 sg13g2_fill_1 FILLER_60_276 ();
 sg13g2_fill_1 FILLER_60_307 ();
 sg13g2_decap_4 FILLER_60_325 ();
 sg13g2_fill_1 FILLER_60_329 ();
 sg13g2_fill_1 FILLER_60_350 ();
 sg13g2_fill_2 FILLER_60_355 ();
 sg13g2_decap_4 FILLER_60_369 ();
 sg13g2_decap_4 FILLER_60_379 ();
 sg13g2_decap_8 FILLER_60_392 ();
 sg13g2_decap_4 FILLER_60_399 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_4 FILLER_61_91 ();
 sg13g2_fill_1 FILLER_61_116 ();
 sg13g2_fill_2 FILLER_61_127 ();
 sg13g2_decap_8 FILLER_61_159 ();
 sg13g2_decap_8 FILLER_61_166 ();
 sg13g2_fill_1 FILLER_61_173 ();
 sg13g2_fill_2 FILLER_61_189 ();
 sg13g2_fill_1 FILLER_61_191 ();
 sg13g2_decap_8 FILLER_61_200 ();
 sg13g2_fill_2 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_223 ();
 sg13g2_fill_2 FILLER_61_229 ();
 sg13g2_fill_1 FILLER_61_231 ();
 sg13g2_fill_2 FILLER_61_241 ();
 sg13g2_fill_1 FILLER_61_243 ();
 sg13g2_fill_1 FILLER_61_336 ();
 sg13g2_decap_4 FILLER_61_352 ();
 sg13g2_fill_1 FILLER_61_356 ();
 sg13g2_fill_2 FILLER_61_374 ();
 sg13g2_fill_1 FILLER_61_376 ();
 sg13g2_fill_1 FILLER_61_394 ();
 sg13g2_fill_1 FILLER_61_405 ();
 sg13g2_fill_1 FILLER_61_413 ();
 sg13g2_fill_2 FILLER_61_423 ();
 sg13g2_fill_1 FILLER_61_429 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_4 FILLER_62_91 ();
 sg13g2_fill_2 FILLER_62_95 ();
 sg13g2_fill_1 FILLER_62_114 ();
 sg13g2_fill_1 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_134 ();
 sg13g2_fill_2 FILLER_62_139 ();
 sg13g2_fill_2 FILLER_62_184 ();
 sg13g2_fill_2 FILLER_62_212 ();
 sg13g2_fill_1 FILLER_62_214 ();
 sg13g2_decap_8 FILLER_62_235 ();
 sg13g2_decap_8 FILLER_62_242 ();
 sg13g2_fill_1 FILLER_62_249 ();
 sg13g2_decap_8 FILLER_62_254 ();
 sg13g2_fill_2 FILLER_62_266 ();
 sg13g2_fill_1 FILLER_62_268 ();
 sg13g2_fill_1 FILLER_62_273 ();
 sg13g2_decap_4 FILLER_62_291 ();
 sg13g2_fill_1 FILLER_62_295 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_decap_4 FILLER_62_308 ();
 sg13g2_fill_2 FILLER_62_312 ();
 sg13g2_fill_2 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_328 ();
 sg13g2_fill_2 FILLER_62_335 ();
 sg13g2_fill_2 FILLER_62_340 ();
 sg13g2_fill_2 FILLER_62_347 ();
 sg13g2_fill_2 FILLER_62_354 ();
 sg13g2_fill_1 FILLER_62_356 ();
 sg13g2_fill_1 FILLER_62_367 ();
 sg13g2_fill_2 FILLER_62_399 ();
 sg13g2_fill_1 FILLER_62_401 ();
 sg13g2_fill_2 FILLER_62_427 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_fill_2 FILLER_63_84 ();
 sg13g2_decap_4 FILLER_63_133 ();
 sg13g2_fill_1 FILLER_63_137 ();
 sg13g2_fill_2 FILLER_63_167 ();
 sg13g2_fill_1 FILLER_63_169 ();
 sg13g2_fill_1 FILLER_63_188 ();
 sg13g2_fill_2 FILLER_63_206 ();
 sg13g2_fill_2 FILLER_63_225 ();
 sg13g2_decap_4 FILLER_63_237 ();
 sg13g2_fill_2 FILLER_63_241 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_fill_1 FILLER_63_269 ();
 sg13g2_decap_4 FILLER_63_292 ();
 sg13g2_fill_2 FILLER_63_296 ();
 sg13g2_decap_4 FILLER_63_302 ();
 sg13g2_fill_1 FILLER_63_327 ();
 sg13g2_fill_2 FILLER_63_333 ();
 sg13g2_fill_1 FILLER_63_365 ();
 sg13g2_fill_2 FILLER_63_376 ();
 sg13g2_decap_8 FILLER_63_423 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_95 ();
 sg13g2_fill_1 FILLER_64_106 ();
 sg13g2_decap_4 FILLER_64_127 ();
 sg13g2_fill_1 FILLER_64_137 ();
 sg13g2_fill_1 FILLER_64_145 ();
 sg13g2_fill_2 FILLER_64_154 ();
 sg13g2_fill_1 FILLER_64_160 ();
 sg13g2_decap_4 FILLER_64_191 ();
 sg13g2_fill_1 FILLER_64_199 ();
 sg13g2_fill_2 FILLER_64_252 ();
 sg13g2_fill_1 FILLER_64_254 ();
 sg13g2_fill_1 FILLER_64_275 ();
 sg13g2_fill_2 FILLER_64_326 ();
 sg13g2_fill_1 FILLER_64_328 ();
 sg13g2_fill_1 FILLER_64_334 ();
 sg13g2_fill_2 FILLER_64_340 ();
 sg13g2_fill_1 FILLER_64_342 ();
 sg13g2_fill_1 FILLER_64_400 ();
 sg13g2_fill_1 FILLER_64_411 ();
 sg13g2_fill_1 FILLER_64_429 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_4 FILLER_65_98 ();
 sg13g2_fill_1 FILLER_65_131 ();
 sg13g2_decap_8 FILLER_65_137 ();
 sg13g2_fill_2 FILLER_65_144 ();
 sg13g2_fill_2 FILLER_65_184 ();
 sg13g2_fill_1 FILLER_65_186 ();
 sg13g2_fill_1 FILLER_65_192 ();
 sg13g2_decap_8 FILLER_65_198 ();
 sg13g2_fill_2 FILLER_65_205 ();
 sg13g2_fill_1 FILLER_65_207 ();
 sg13g2_decap_4 FILLER_65_212 ();
 sg13g2_fill_1 FILLER_65_216 ();
 sg13g2_fill_2 FILLER_65_221 ();
 sg13g2_decap_4 FILLER_65_233 ();
 sg13g2_fill_1 FILLER_65_237 ();
 sg13g2_fill_1 FILLER_65_262 ();
 sg13g2_fill_2 FILLER_65_266 ();
 sg13g2_fill_2 FILLER_65_292 ();
 sg13g2_fill_1 FILLER_65_298 ();
 sg13g2_fill_1 FILLER_65_321 ();
 sg13g2_decap_8 FILLER_65_391 ();
 sg13g2_fill_2 FILLER_65_422 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_4 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_fill_2 FILLER_66_119 ();
 sg13g2_fill_2 FILLER_66_140 ();
 sg13g2_fill_1 FILLER_66_142 ();
 sg13g2_decap_4 FILLER_66_147 ();
 sg13g2_fill_2 FILLER_66_151 ();
 sg13g2_fill_1 FILLER_66_170 ();
 sg13g2_fill_2 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_195 ();
 sg13g2_fill_2 FILLER_66_202 ();
 sg13g2_decap_4 FILLER_66_209 ();
 sg13g2_fill_1 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_235 ();
 sg13g2_decap_4 FILLER_66_242 ();
 sg13g2_fill_1 FILLER_66_246 ();
 sg13g2_decap_4 FILLER_66_262 ();
 sg13g2_fill_2 FILLER_66_266 ();
 sg13g2_fill_2 FILLER_66_272 ();
 sg13g2_fill_1 FILLER_66_274 ();
 sg13g2_fill_1 FILLER_66_295 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_318 ();
 sg13g2_fill_1 FILLER_66_341 ();
 sg13g2_fill_2 FILLER_66_405 ();
 sg13g2_fill_1 FILLER_66_429 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_4 FILLER_67_91 ();
 sg13g2_fill_1 FILLER_67_95 ();
 sg13g2_fill_1 FILLER_67_150 ();
 sg13g2_decap_4 FILLER_67_164 ();
 sg13g2_fill_2 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_237 ();
 sg13g2_fill_2 FILLER_67_244 ();
 sg13g2_fill_1 FILLER_67_246 ();
 sg13g2_fill_1 FILLER_67_262 ();
 sg13g2_fill_1 FILLER_67_268 ();
 sg13g2_fill_1 FILLER_67_279 ();
 sg13g2_decap_4 FILLER_67_297 ();
 sg13g2_fill_2 FILLER_67_301 ();
 sg13g2_fill_1 FILLER_67_310 ();
 sg13g2_fill_1 FILLER_67_321 ();
 sg13g2_fill_1 FILLER_67_341 ();
 sg13g2_fill_1 FILLER_67_347 ();
 sg13g2_fill_2 FILLER_67_379 ();
 sg13g2_fill_1 FILLER_67_429 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_fill_2 FILLER_68_125 ();
 sg13g2_fill_1 FILLER_68_127 ();
 sg13g2_fill_1 FILLER_68_146 ();
 sg13g2_fill_1 FILLER_68_151 ();
 sg13g2_fill_1 FILLER_68_156 ();
 sg13g2_fill_2 FILLER_68_161 ();
 sg13g2_fill_1 FILLER_68_168 ();
 sg13g2_fill_1 FILLER_68_173 ();
 sg13g2_fill_1 FILLER_68_192 ();
 sg13g2_decap_4 FILLER_68_196 ();
 sg13g2_fill_1 FILLER_68_200 ();
 sg13g2_fill_2 FILLER_68_209 ();
 sg13g2_fill_1 FILLER_68_211 ();
 sg13g2_fill_1 FILLER_68_219 ();
 sg13g2_fill_1 FILLER_68_227 ();
 sg13g2_fill_1 FILLER_68_239 ();
 sg13g2_fill_1 FILLER_68_249 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_2 FILLER_68_298 ();
 sg13g2_fill_1 FILLER_68_300 ();
 sg13g2_decap_8 FILLER_68_311 ();
 sg13g2_fill_2 FILLER_68_318 ();
 sg13g2_decap_4 FILLER_68_323 ();
 sg13g2_fill_2 FILLER_68_346 ();
 sg13g2_fill_1 FILLER_68_379 ();
 sg13g2_fill_1 FILLER_68_385 ();
 sg13g2_fill_1 FILLER_68_399 ();
 sg13g2_fill_1 FILLER_68_404 ();
 sg13g2_fill_2 FILLER_68_415 ();
 sg13g2_fill_2 FILLER_68_427 ();
 sg13g2_fill_1 FILLER_68_429 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_fill_2 FILLER_69_105 ();
 sg13g2_fill_1 FILLER_69_107 ();
 sg13g2_fill_1 FILLER_69_113 ();
 sg13g2_fill_2 FILLER_69_140 ();
 sg13g2_fill_1 FILLER_69_172 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_fill_1 FILLER_69_186 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_208 ();
 sg13g2_fill_1 FILLER_69_222 ();
 sg13g2_fill_2 FILLER_69_300 ();
 sg13g2_decap_8 FILLER_69_317 ();
 sg13g2_decap_8 FILLER_69_324 ();
 sg13g2_decap_4 FILLER_69_331 ();
 sg13g2_fill_1 FILLER_69_365 ();
 sg13g2_fill_2 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_fill_2 FILLER_69_410 ();
 sg13g2_decap_8 FILLER_69_419 ();
 sg13g2_decap_4 FILLER_69_426 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_fill_2 FILLER_70_131 ();
 sg13g2_fill_1 FILLER_70_150 ();
 sg13g2_fill_1 FILLER_70_156 ();
 sg13g2_fill_1 FILLER_70_175 ();
 sg13g2_fill_2 FILLER_70_197 ();
 sg13g2_fill_1 FILLER_70_210 ();
 sg13g2_fill_2 FILLER_70_255 ();
 sg13g2_fill_2 FILLER_70_267 ();
 sg13g2_fill_2 FILLER_70_274 ();
 sg13g2_fill_1 FILLER_70_323 ();
 sg13g2_fill_1 FILLER_70_329 ();
 sg13g2_fill_1 FILLER_70_340 ();
 sg13g2_decap_8 FILLER_70_344 ();
 sg13g2_fill_2 FILLER_70_351 ();
 sg13g2_fill_1 FILLER_70_353 ();
 sg13g2_decap_8 FILLER_70_367 ();
 sg13g2_fill_1 FILLER_70_374 ();
 sg13g2_decap_8 FILLER_70_379 ();
 sg13g2_decap_4 FILLER_70_386 ();
 sg13g2_fill_1 FILLER_70_394 ();
 sg13g2_fill_1 FILLER_70_413 ();
 sg13g2_fill_1 FILLER_70_429 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_4 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_106 ();
 sg13g2_fill_2 FILLER_71_113 ();
 sg13g2_fill_1 FILLER_71_115 ();
 sg13g2_fill_1 FILLER_71_141 ();
 sg13g2_fill_2 FILLER_71_145 ();
 sg13g2_fill_1 FILLER_71_153 ();
 sg13g2_fill_1 FILLER_71_161 ();
 sg13g2_fill_1 FILLER_71_167 ();
 sg13g2_fill_1 FILLER_71_174 ();
 sg13g2_fill_2 FILLER_71_185 ();
 sg13g2_decap_8 FILLER_71_191 ();
 sg13g2_decap_8 FILLER_71_198 ();
 sg13g2_fill_1 FILLER_71_205 ();
 sg13g2_fill_1 FILLER_71_211 ();
 sg13g2_fill_1 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_228 ();
 sg13g2_fill_1 FILLER_71_235 ();
 sg13g2_decap_8 FILLER_71_243 ();
 sg13g2_decap_4 FILLER_71_250 ();
 sg13g2_fill_2 FILLER_71_254 ();
 sg13g2_fill_1 FILLER_71_356 ();
 sg13g2_fill_1 FILLER_71_405 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_fill_2 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_190 ();
 sg13g2_decap_8 FILLER_72_197 ();
 sg13g2_fill_2 FILLER_72_221 ();
 sg13g2_decap_8 FILLER_72_241 ();
 sg13g2_decap_8 FILLER_72_248 ();
 sg13g2_decap_8 FILLER_72_255 ();
 sg13g2_fill_1 FILLER_72_262 ();
 sg13g2_decap_8 FILLER_72_276 ();
 sg13g2_decap_8 FILLER_72_283 ();
 sg13g2_fill_2 FILLER_72_299 ();
 sg13g2_fill_1 FILLER_72_312 ();
 sg13g2_fill_1 FILLER_72_318 ();
 sg13g2_fill_2 FILLER_72_324 ();
 sg13g2_fill_1 FILLER_72_402 ();
 sg13g2_fill_2 FILLER_72_428 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_4 FILLER_73_105 ();
 sg13g2_fill_2 FILLER_73_109 ();
 sg13g2_fill_1 FILLER_73_128 ();
 sg13g2_fill_1 FILLER_73_133 ();
 sg13g2_fill_2 FILLER_73_139 ();
 sg13g2_fill_2 FILLER_73_151 ();
 sg13g2_decap_8 FILLER_73_156 ();
 sg13g2_fill_1 FILLER_73_179 ();
 sg13g2_fill_2 FILLER_73_190 ();
 sg13g2_fill_1 FILLER_73_202 ();
 sg13g2_fill_2 FILLER_73_208 ();
 sg13g2_fill_2 FILLER_73_256 ();
 sg13g2_fill_2 FILLER_73_284 ();
 sg13g2_fill_1 FILLER_73_286 ();
 sg13g2_fill_1 FILLER_73_292 ();
 sg13g2_decap_8 FILLER_73_297 ();
 sg13g2_fill_1 FILLER_73_304 ();
 sg13g2_fill_1 FILLER_73_314 ();
 sg13g2_fill_2 FILLER_73_331 ();
 sg13g2_fill_1 FILLER_73_333 ();
 sg13g2_decap_4 FILLER_73_384 ();
 sg13g2_fill_1 FILLER_73_395 ();
 sg13g2_fill_1 FILLER_73_404 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_fill_2 FILLER_74_105 ();
 sg13g2_fill_1 FILLER_74_107 ();
 sg13g2_decap_8 FILLER_74_125 ();
 sg13g2_decap_8 FILLER_74_132 ();
 sg13g2_decap_4 FILLER_74_139 ();
 sg13g2_fill_1 FILLER_74_143 ();
 sg13g2_fill_1 FILLER_74_148 ();
 sg13g2_fill_2 FILLER_74_154 ();
 sg13g2_fill_2 FILLER_74_161 ();
 sg13g2_fill_1 FILLER_74_168 ();
 sg13g2_fill_1 FILLER_74_272 ();
 sg13g2_fill_2 FILLER_74_279 ();
 sg13g2_fill_1 FILLER_74_281 ();
 sg13g2_fill_1 FILLER_74_308 ();
 sg13g2_fill_2 FILLER_74_338 ();
 sg13g2_fill_2 FILLER_74_364 ();
 sg13g2_fill_2 FILLER_74_384 ();
 sg13g2_decap_4 FILLER_74_390 ();
 sg13g2_fill_2 FILLER_74_394 ();
 sg13g2_fill_1 FILLER_74_409 ();
 sg13g2_fill_2 FILLER_74_422 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_4 FILLER_75_126 ();
 sg13g2_fill_1 FILLER_75_130 ();
 sg13g2_decap_4 FILLER_75_175 ();
 sg13g2_fill_1 FILLER_75_179 ();
 sg13g2_decap_4 FILLER_75_217 ();
 sg13g2_fill_2 FILLER_75_221 ();
 sg13g2_fill_1 FILLER_75_228 ();
 sg13g2_fill_2 FILLER_75_239 ();
 sg13g2_fill_1 FILLER_75_261 ();
 sg13g2_decap_8 FILLER_75_307 ();
 sg13g2_fill_2 FILLER_75_319 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_fill_2 FILLER_75_349 ();
 sg13g2_fill_1 FILLER_75_351 ();
 sg13g2_fill_1 FILLER_75_356 ();
 sg13g2_fill_2 FILLER_75_361 ();
 sg13g2_fill_1 FILLER_75_373 ();
 sg13g2_fill_1 FILLER_75_405 ();
 sg13g2_fill_2 FILLER_75_428 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_4 FILLER_76_105 ();
 sg13g2_fill_2 FILLER_76_109 ();
 sg13g2_fill_1 FILLER_76_141 ();
 sg13g2_decap_4 FILLER_76_181 ();
 sg13g2_fill_2 FILLER_76_212 ();
 sg13g2_fill_2 FILLER_76_231 ();
 sg13g2_fill_2 FILLER_76_261 ();
 sg13g2_fill_1 FILLER_76_263 ();
 sg13g2_fill_1 FILLER_76_286 ();
 sg13g2_fill_1 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_301 ();
 sg13g2_fill_2 FILLER_76_407 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_fill_2 FILLER_77_173 ();
 sg13g2_decap_8 FILLER_77_191 ();
 sg13g2_fill_1 FILLER_77_198 ();
 sg13g2_decap_8 FILLER_77_234 ();
 sg13g2_fill_1 FILLER_77_241 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_fill_1 FILLER_77_290 ();
 sg13g2_fill_1 FILLER_77_393 ();
 sg13g2_fill_1 FILLER_77_399 ();
 sg13g2_fill_1 FILLER_77_410 ();
 sg13g2_fill_2 FILLER_77_428 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_4 FILLER_78_119 ();
 sg13g2_fill_2 FILLER_78_199 ();
 sg13g2_fill_2 FILLER_78_252 ();
 sg13g2_fill_2 FILLER_78_258 ();
 sg13g2_fill_1 FILLER_78_260 ();
 sg13g2_fill_1 FILLER_78_305 ();
 sg13g2_fill_1 FILLER_78_310 ();
 sg13g2_fill_1 FILLER_78_314 ();
 sg13g2_fill_1 FILLER_78_336 ();
 sg13g2_fill_1 FILLER_78_342 ();
 sg13g2_fill_1 FILLER_78_368 ();
 sg13g2_fill_1 FILLER_78_390 ();
 sg13g2_fill_2 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_419 ();
 sg13g2_decap_4 FILLER_78_426 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_4 FILLER_79_70 ();
 sg13g2_fill_2 FILLER_79_74 ();
 sg13g2_decap_4 FILLER_79_80 ();
 sg13g2_decap_8 FILLER_79_88 ();
 sg13g2_decap_8 FILLER_79_95 ();
 sg13g2_fill_2 FILLER_79_102 ();
 sg13g2_fill_2 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_114 ();
 sg13g2_fill_1 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_124 ();
 sg13g2_fill_1 FILLER_79_184 ();
 sg13g2_fill_2 FILLER_79_232 ();
 sg13g2_fill_1 FILLER_79_234 ();
 sg13g2_fill_1 FILLER_79_338 ();
 sg13g2_fill_1 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_fill_2 FILLER_79_427 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_89 ();
 sg13g2_fill_1 FILLER_80_94 ();
 sg13g2_fill_1 FILLER_80_103 ();
 sg13g2_fill_1 FILLER_80_124 ();
 sg13g2_fill_1 FILLER_80_167 ();
 sg13g2_fill_1 FILLER_80_176 ();
 sg13g2_fill_2 FILLER_80_201 ();
 sg13g2_fill_2 FILLER_80_219 ();
 sg13g2_decap_4 FILLER_80_241 ();
 sg13g2_fill_2 FILLER_80_245 ();
 sg13g2_fill_1 FILLER_80_251 ();
 sg13g2_fill_2 FILLER_80_264 ();
 sg13g2_fill_1 FILLER_80_266 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_fill_1 FILLER_80_277 ();
 sg13g2_fill_1 FILLER_80_282 ();
 sg13g2_fill_2 FILLER_80_287 ();
 sg13g2_fill_1 FILLER_80_303 ();
 sg13g2_decap_8 FILLER_80_410 ();
 sg13g2_decap_8 FILLER_80_417 ();
 sg13g2_decap_4 FILLER_80_424 ();
 sg13g2_fill_2 FILLER_80_428 ();
endmodule
