module tt_um_rajum_iterativeMAC (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire clknet_0_clk;
 wire \ad.a[0] ;
 wire \ad.a[10] ;
 wire \ad.a[11] ;
 wire \ad.a[12] ;
 wire \ad.a[13] ;
 wire \ad.a[14] ;
 wire \ad.a[15] ;
 wire \ad.a[16] ;
 wire \ad.a[17] ;
 wire \ad.a[18] ;
 wire \ad.a[19] ;
 wire \ad.a[1] ;
 wire \ad.a[20] ;
 wire \ad.a[21] ;
 wire \ad.a[22] ;
 wire \ad.a[23] ;
 wire \ad.a[24] ;
 wire \ad.a[25] ;
 wire \ad.a[26] ;
 wire \ad.a[27] ;
 wire \ad.a[28] ;
 wire \ad.a[29] ;
 wire \ad.a[2] ;
 wire \ad.a[30] ;
 wire \ad.a[31] ;
 wire \ad.a[3] ;
 wire \ad.a[4] ;
 wire \ad.a[5] ;
 wire \ad.a[6] ;
 wire \ad.a[7] ;
 wire \ad.a[8] ;
 wire \ad.a[9] ;
 wire \inp_a[0] ;
 wire \inp_a[1] ;
 wire \inp_a[2] ;
 wire \inp_a[3] ;
 wire \inp_a[4] ;
 wire \inp_a[5] ;
 wire \inp_a[6] ;
 wire mode;
 wire \result[0] ;
 wire \result[10] ;
 wire \result[11] ;
 wire \result[12] ;
 wire \result[13] ;
 wire \result[14] ;
 wire \result[15] ;
 wire \result[16] ;
 wire \result[17] ;
 wire \result[18] ;
 wire \result[19] ;
 wire \result[1] ;
 wire \result[20] ;
 wire \result[21] ;
 wire \result[22] ;
 wire \result[23] ;
 wire \result[24] ;
 wire \result[25] ;
 wire \result[26] ;
 wire \result[27] ;
 wire \result[28] ;
 wire \result[29] ;
 wire \result[2] ;
 wire \result[30] ;
 wire \result[31] ;
 wire \result[3] ;
 wire \result[4] ;
 wire \result[5] ;
 wire \result[6] ;
 wire \result[7] ;
 wire \result[8] ;
 wire \result[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _1434_ (.A(ui_in[0]),
    .X(_0552_));
 sg13g2_buf_1 _1435_ (.A(_0552_),
    .X(_0553_));
 sg13g2_buf_8 _1436_ (.A(\inp_a[0] ),
    .X(_0554_));
 sg13g2_buf_1 _1437_ (.A(net100),
    .X(_0555_));
 sg13g2_buf_1 _1438_ (.A(rst_n),
    .X(_0556_));
 sg13g2_mux2_1 _1439_ (.A0(net101),
    .A1(net92),
    .S(_0556_),
    .X(_0010_));
 sg13g2_buf_1 _1440_ (.A(net1),
    .X(_0557_));
 sg13g2_buf_1 _1441_ (.A(\inp_a[1] ),
    .X(_0558_));
 sg13g2_mux2_1 _1442_ (.A0(net107),
    .A1(_0558_),
    .S(net108),
    .X(_0011_));
 sg13g2_buf_1 _1443_ (.A(net2),
    .X(_0559_));
 sg13g2_buf_8 _1444_ (.A(\inp_a[2] ),
    .X(_0560_));
 sg13g2_buf_1 _1445_ (.A(net98),
    .X(_0561_));
 sg13g2_mux2_1 _1446_ (.A0(net106),
    .A1(_0561_),
    .S(_0556_),
    .X(_0012_));
 sg13g2_buf_1 _1447_ (.A(net3),
    .X(_0562_));
 sg13g2_buf_2 _1448_ (.A(\inp_a[3] ),
    .X(_0563_));
 sg13g2_buf_1 _1449_ (.A(_0563_),
    .X(_0564_));
 sg13g2_mux2_1 _1450_ (.A0(net105),
    .A1(net90),
    .S(net108),
    .X(_0013_));
 sg13g2_buf_2 _1451_ (.A(ui_in[4]),
    .X(_0565_));
 sg13g2_buf_8 _1452_ (.A(\inp_a[4] ),
    .X(_0566_));
 sg13g2_buf_1 _1453_ (.A(_0566_),
    .X(_0567_));
 sg13g2_mux2_1 _1454_ (.A0(net104),
    .A1(_0567_),
    .S(net108),
    .X(_0014_));
 sg13g2_buf_2 _1455_ (.A(ui_in[5]),
    .X(_0568_));
 sg13g2_buf_1 _1456_ (.A(_0568_),
    .X(_0569_));
 sg13g2_inv_1 _1457_ (.Y(_0570_),
    .A(net97));
 sg13g2_buf_1 _1458_ (.A(net108),
    .X(_0571_));
 sg13g2_buf_2 _1459_ (.A(\inp_a[5] ),
    .X(_0572_));
 sg13g2_buf_1 _1460_ (.A(_0572_),
    .X(_0573_));
 sg13g2_nand2_1 _1461_ (.Y(_0574_),
    .A(net88),
    .B(net96));
 sg13g2_o21ai_1 _1462_ (.B1(_0574_),
    .Y(_0015_),
    .A1(_0570_),
    .A2(net96));
 sg13g2_buf_2 _1463_ (.A(ui_in[6]),
    .X(_0575_));
 sg13g2_buf_1 _1464_ (.A(_0575_),
    .X(_0576_));
 sg13g2_inv_1 _1465_ (.Y(_0577_),
    .A(net95));
 sg13g2_buf_1 _1466_ (.A(\inp_a[6] ),
    .X(_0578_));
 sg13g2_buf_1 _1467_ (.A(_0578_),
    .X(_0579_));
 sg13g2_nand2_1 _1468_ (.Y(_0580_),
    .A(net87),
    .B(net96));
 sg13g2_o21ai_1 _1469_ (.B1(_0580_),
    .Y(_0016_),
    .A1(_0577_),
    .A2(net96));
 sg13g2_buf_1 _1470_ (.A(ui_in[7]),
    .X(_0581_));
 sg13g2_buf_1 _1471_ (.A(net103),
    .X(_0582_));
 sg13g2_mux2_1 _1472_ (.A0(_0582_),
    .A1(mode),
    .S(net108),
    .X(_0017_));
 sg13g2_inv_1 _1473_ (.Y(_0583_),
    .A(net108));
 sg13g2_buf_1 _1474_ (.A(_0583_),
    .X(_0584_));
 sg13g2_buf_1 _1475_ (.A(net86),
    .X(_0585_));
 sg13g2_buf_1 _1476_ (.A(\state[0] ),
    .X(_0586_));
 sg13g2_buf_1 _1477_ (.A(_0586_),
    .X(_0587_));
 sg13g2_buf_1 _1478_ (.A(net85),
    .X(_0588_));
 sg13g2_buf_1 _1479_ (.A(net75),
    .X(_0589_));
 sg13g2_buf_2 _1480_ (.A(\state[1] ),
    .X(_0590_));
 sg13g2_buf_1 _1481_ (.A(_0590_),
    .X(_0591_));
 sg13g2_buf_1 _1482_ (.A(net84),
    .X(_0592_));
 sg13g2_buf_1 _1483_ (.A(net74),
    .X(_0593_));
 sg13g2_nor2_1 _1484_ (.A(net68),
    .B(net67),
    .Y(_0594_));
 sg13g2_and2_1 _1485_ (.A(_0004_),
    .B(_0594_),
    .X(_0595_));
 sg13g2_buf_1 _1486_ (.A(_0595_),
    .X(_0596_));
 sg13g2_buf_1 _1487_ (.A(net53),
    .X(_0597_));
 sg13g2_buf_1 _1488_ (.A(\ad.a[0] ),
    .X(_0598_));
 sg13g2_buf_1 _1489_ (.A(\state[2] ),
    .X(_0599_));
 sg13g2_and2_1 _1490_ (.A(_0555_),
    .B(net101),
    .X(_0600_));
 sg13g2_nor2b_1 _1491_ (.A(net93),
    .B_N(net4),
    .Y(_0601_));
 sg13g2_a21oi_1 _1492_ (.A1(net93),
    .A2(_0600_),
    .Y(_0602_),
    .B1(_0601_));
 sg13g2_inv_2 _1493_ (.Y(_0603_),
    .A(_0586_));
 sg13g2_nand2_1 _1494_ (.Y(_0604_),
    .A(_0603_),
    .B(_0590_));
 sg13g2_nand2_1 _1495_ (.Y(_0605_),
    .A(\state[2] ),
    .B(net4));
 sg13g2_nor2_1 _1496_ (.A(_0590_),
    .B(_0605_),
    .Y(_0606_));
 sg13g2_nand2_1 _1497_ (.Y(_0607_),
    .A(_0555_),
    .B(_0553_));
 sg13g2_inv_1 _1498_ (.Y(_0608_),
    .A(\state[2] ));
 sg13g2_nand2_2 _1499_ (.Y(_0609_),
    .A(_0590_),
    .B(_0608_));
 sg13g2_nor2_1 _1500_ (.A(_0607_),
    .B(_0609_),
    .Y(_0610_));
 sg13g2_o21ai_1 _1501_ (.B1(_0586_),
    .Y(_0611_),
    .A1(_0606_),
    .A2(_0610_));
 sg13g2_o21ai_1 _1502_ (.B1(_0611_),
    .Y(_0612_),
    .A1(_0602_),
    .A2(_0604_));
 sg13g2_nand2_1 _1503_ (.Y(_0613_),
    .A(_0566_),
    .B(net1));
 sg13g2_nand2_1 _1504_ (.Y(_0614_),
    .A(_0572_),
    .B(_0552_));
 sg13g2_nand2_1 _1505_ (.Y(_0615_),
    .A(_0613_),
    .B(_0614_));
 sg13g2_nand2_2 _1506_ (.Y(_0616_),
    .A(_0563_),
    .B(net106));
 sg13g2_o21ai_1 _1507_ (.B1(_0616_),
    .Y(_0617_),
    .A1(_0613_),
    .A2(_0614_));
 sg13g2_nand2_2 _1508_ (.Y(_0618_),
    .A(_0615_),
    .B(_0617_));
 sg13g2_nand2_2 _1509_ (.Y(_0619_),
    .A(net98),
    .B(net104));
 sg13g2_nand2_1 _1510_ (.Y(_0620_),
    .A(_0575_),
    .B(net100));
 sg13g2_nand2_1 _1511_ (.Y(_0621_),
    .A(\inp_a[1] ),
    .B(_0568_));
 sg13g2_xor2_1 _1512_ (.B(_0621_),
    .A(_0620_),
    .X(_0622_));
 sg13g2_xor2_1 _1513_ (.B(_0622_),
    .A(_0619_),
    .X(_0623_));
 sg13g2_nand2_1 _1514_ (.Y(_0624_),
    .A(_0618_),
    .B(_0623_));
 sg13g2_xnor2_1 _1515_ (.Y(_0625_),
    .A(_0619_),
    .B(_0622_));
 sg13g2_nand2_1 _1516_ (.Y(_0626_),
    .A(_0618_),
    .B(_0625_));
 sg13g2_nand2_2 _1517_ (.Y(_0627_),
    .A(net98),
    .B(net105));
 sg13g2_nand2_1 _1518_ (.Y(_0628_),
    .A(net100),
    .B(_0568_));
 sg13g2_nand2_1 _1519_ (.Y(_0629_),
    .A(net99),
    .B(_0565_));
 sg13g2_a21o_1 _1520_ (.A2(_0628_),
    .A1(_0627_),
    .B1(_0629_),
    .X(_0630_));
 sg13g2_o21ai_1 _1521_ (.B1(_0630_),
    .Y(_0631_),
    .A1(_0627_),
    .A2(_0628_));
 sg13g2_nand2_2 _1522_ (.Y(_0632_),
    .A(_0572_),
    .B(net107));
 sg13g2_nand2_1 _1523_ (.Y(_0633_),
    .A(_0563_),
    .B(net105));
 sg13g2_nand2_1 _1524_ (.Y(_0634_),
    .A(_0566_),
    .B(net2));
 sg13g2_xor2_1 _1525_ (.B(_0634_),
    .A(_0633_),
    .X(_0635_));
 sg13g2_xor2_1 _1526_ (.B(_0635_),
    .A(_0632_),
    .X(_0636_));
 sg13g2_xnor2_1 _1527_ (.Y(_0637_),
    .A(_0631_),
    .B(_0636_));
 sg13g2_mux2_1 _1528_ (.A0(_0624_),
    .A1(_0626_),
    .S(_0637_),
    .X(_0638_));
 sg13g2_and2_1 _1529_ (.A(net100),
    .B(_0568_),
    .X(_0639_));
 sg13g2_xnor2_1 _1530_ (.Y(_0640_),
    .A(_0639_),
    .B(_0629_));
 sg13g2_xnor2_1 _1531_ (.Y(_0641_),
    .A(_0627_),
    .B(_0640_));
 sg13g2_nand2_2 _1532_ (.Y(_0642_),
    .A(_0566_),
    .B(_0552_));
 sg13g2_nand2_1 _1533_ (.Y(_0643_),
    .A(_0563_),
    .B(net107));
 sg13g2_nand2_2 _1534_ (.Y(_0644_),
    .A(_0572_),
    .B(net106));
 sg13g2_nor3_1 _1535_ (.A(_0642_),
    .B(_0643_),
    .C(_0644_),
    .Y(_0645_));
 sg13g2_nor2_1 _1536_ (.A(_0641_),
    .B(_0645_),
    .Y(_0646_));
 sg13g2_xor2_1 _1537_ (.B(_0614_),
    .A(_0613_),
    .X(_0647_));
 sg13g2_xnor2_1 _1538_ (.Y(_0648_),
    .A(_0616_),
    .B(_0647_));
 sg13g2_nand2_1 _1539_ (.Y(_0649_),
    .A(net98),
    .B(net2));
 sg13g2_nand2_1 _1540_ (.Y(_0650_),
    .A(net100),
    .B(net104));
 sg13g2_nand2_2 _1541_ (.Y(_0651_),
    .A(net99),
    .B(net105));
 sg13g2_a21o_1 _1542_ (.A2(_0650_),
    .A1(_0649_),
    .B1(_0651_),
    .X(_0652_));
 sg13g2_o21ai_1 _1543_ (.B1(_0652_),
    .Y(_0653_),
    .A1(_0649_),
    .A2(_0650_));
 sg13g2_a21o_1 _1544_ (.A2(_0648_),
    .A1(_0641_),
    .B1(_0653_),
    .X(_0654_));
 sg13g2_nor2b_1 _1545_ (.A(_0646_),
    .B_N(_0654_),
    .Y(_0655_));
 sg13g2_nand2_1 _1546_ (.Y(_0656_),
    .A(_0653_),
    .B(_0648_));
 sg13g2_nand2_1 _1547_ (.Y(_0657_),
    .A(_0656_),
    .B(_0618_));
 sg13g2_xnor2_1 _1548_ (.Y(_0658_),
    .A(_0623_),
    .B(_0637_));
 sg13g2_a22oi_1 _1549_ (.Y(_0659_),
    .B1(_0657_),
    .B2(_0658_),
    .A2(_0655_),
    .A1(_0638_));
 sg13g2_buf_2 _1550_ (.A(_0659_),
    .X(_0660_));
 sg13g2_nand2_1 _1551_ (.Y(_0661_),
    .A(net107),
    .B(_0578_));
 sg13g2_and2_1 _1552_ (.A(\inp_a[1] ),
    .B(_0575_),
    .X(_0662_));
 sg13g2_buf_1 _1553_ (.A(_0662_),
    .X(_0663_));
 sg13g2_nand2_1 _1554_ (.Y(_0664_),
    .A(net91),
    .B(_0569_));
 sg13g2_and2_1 _1555_ (.A(net103),
    .B(net100),
    .X(_0665_));
 sg13g2_xnor2_1 _1556_ (.Y(_0666_),
    .A(_0664_),
    .B(_0665_));
 sg13g2_xnor2_1 _1557_ (.Y(_0667_),
    .A(_0663_),
    .B(_0666_));
 sg13g2_a21o_1 _1558_ (.A2(_0620_),
    .A1(_0619_),
    .B1(_0621_),
    .X(_0668_));
 sg13g2_o21ai_1 _1559_ (.B1(_0668_),
    .Y(_0669_),
    .A1(_0619_),
    .A2(_0620_));
 sg13g2_buf_2 _1560_ (.A(_0669_),
    .X(_0670_));
 sg13g2_nand2_1 _1561_ (.Y(_0671_),
    .A(_0566_),
    .B(net3));
 sg13g2_nand2_1 _1562_ (.Y(_0672_),
    .A(_0563_),
    .B(net104));
 sg13g2_xor2_1 _1563_ (.B(_0672_),
    .A(_0671_),
    .X(_0673_));
 sg13g2_xor2_1 _1564_ (.B(_0673_),
    .A(_0644_),
    .X(_0674_));
 sg13g2_xnor2_1 _1565_ (.Y(_0675_),
    .A(_0670_),
    .B(_0674_));
 sg13g2_xnor2_1 _1566_ (.Y(_0676_),
    .A(_0667_),
    .B(_0675_));
 sg13g2_xnor2_1 _1567_ (.Y(_0677_),
    .A(_0632_),
    .B(_0635_));
 sg13g2_a21o_1 _1568_ (.A2(_0625_),
    .A1(_0677_),
    .B1(_0631_),
    .X(_0678_));
 sg13g2_nand2_1 _1569_ (.Y(_0679_),
    .A(_0632_),
    .B(_0634_));
 sg13g2_o21ai_1 _1570_ (.B1(_0633_),
    .Y(_0680_),
    .A1(_0632_),
    .A2(_0634_));
 sg13g2_nand2_1 _1571_ (.Y(_0681_),
    .A(_0679_),
    .B(_0680_));
 sg13g2_a21oi_1 _1572_ (.A1(_0636_),
    .A2(_0623_),
    .Y(_0682_),
    .B1(_0681_));
 sg13g2_and2_1 _1573_ (.A(_0679_),
    .B(_0680_),
    .X(_0683_));
 sg13g2_a21oi_1 _1574_ (.A1(_0677_),
    .A2(_0625_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_o21ai_1 _1575_ (.B1(_0631_),
    .Y(_0685_),
    .A1(_0677_),
    .A2(_0625_));
 sg13g2_a22oi_1 _1576_ (.Y(_0686_),
    .B1(_0684_),
    .B2(_0685_),
    .A2(_0682_),
    .A1(_0678_));
 sg13g2_xnor2_1 _1577_ (.Y(_0687_),
    .A(_0676_),
    .B(_0686_));
 sg13g2_xor2_1 _1578_ (.B(_0687_),
    .A(_0661_),
    .X(_0688_));
 sg13g2_xnor2_1 _1579_ (.Y(_0689_),
    .A(_0660_),
    .B(_0688_));
 sg13g2_xor2_1 _1580_ (.B(_0647_),
    .A(_0616_),
    .X(_0690_));
 sg13g2_xnor2_1 _1581_ (.Y(_0691_),
    .A(_0653_),
    .B(_0690_));
 sg13g2_xnor2_1 _1582_ (.Y(_0692_),
    .A(_0641_),
    .B(_0691_));
 sg13g2_nand2b_1 _1583_ (.Y(_0693_),
    .B(_0642_),
    .A_N(_0651_));
 sg13g2_nand2_1 _1584_ (.Y(_0694_),
    .A(_0651_),
    .B(_0642_));
 sg13g2_xnor2_1 _1585_ (.Y(_0695_),
    .A(_0649_),
    .B(_0650_));
 sg13g2_mux2_1 _1586_ (.A0(_0693_),
    .A1(_0694_),
    .S(_0695_),
    .X(_0696_));
 sg13g2_and2_1 _1587_ (.A(_0564_),
    .B(net107),
    .X(_0697_));
 sg13g2_a22oi_1 _1588_ (.Y(_0698_),
    .B1(net107),
    .B2(_0560_),
    .A2(net105),
    .A1(net100));
 sg13g2_nand2_1 _1589_ (.Y(_0699_),
    .A(net99),
    .B(net106));
 sg13g2_nand4_1 _1590_ (.B(net100),
    .C(_0562_),
    .A(_0560_),
    .Y(_0700_),
    .D(net107));
 sg13g2_o21ai_1 _1591_ (.B1(_0700_),
    .Y(_0701_),
    .A1(_0698_),
    .A2(_0699_));
 sg13g2_buf_1 _1592_ (.A(_0701_),
    .X(_0702_));
 sg13g2_or2_1 _1593_ (.X(_0703_),
    .B(_0702_),
    .A(_0697_));
 sg13g2_nor2b_1 _1594_ (.A(_0642_),
    .B_N(_0651_),
    .Y(_0704_));
 sg13g2_nor2_1 _1595_ (.A(_0651_),
    .B(_0642_),
    .Y(_0705_));
 sg13g2_mux2_1 _1596_ (.A0(_0704_),
    .A1(_0705_),
    .S(_0695_),
    .X(_0706_));
 sg13g2_buf_2 _1597_ (.A(_0706_),
    .X(_0707_));
 sg13g2_and2_1 _1598_ (.A(_0697_),
    .B(_0702_),
    .X(_0708_));
 sg13g2_buf_1 _1599_ (.A(_0708_),
    .X(_0709_));
 sg13g2_or2_1 _1600_ (.X(_0710_),
    .B(_0709_),
    .A(_0707_));
 sg13g2_a21oi_1 _1601_ (.A1(_0696_),
    .A2(_0703_),
    .Y(_0711_),
    .B1(_0710_));
 sg13g2_nand2_1 _1602_ (.Y(_0712_),
    .A(_0707_),
    .B(_0709_));
 sg13g2_o21ai_1 _1603_ (.B1(_0712_),
    .Y(_0713_),
    .A1(_0692_),
    .A2(_0711_));
 sg13g2_buf_1 _1604_ (.A(_0713_),
    .X(_0714_));
 sg13g2_o21ai_1 _1605_ (.B1(_0696_),
    .Y(_0715_),
    .A1(_0702_),
    .A2(_0707_));
 sg13g2_nor2_1 _1606_ (.A(_0696_),
    .B(_0702_),
    .Y(_0716_));
 sg13g2_a221oi_1 _1607_ (.B2(_0643_),
    .C1(_0716_),
    .B1(_0715_),
    .A1(_0707_),
    .Y(_0717_),
    .A2(_0709_));
 sg13g2_xnor2_1 _1608_ (.Y(_0718_),
    .A(_0692_),
    .B(_0717_));
 sg13g2_xnor2_1 _1609_ (.Y(_0719_),
    .A(_0651_),
    .B(_0695_));
 sg13g2_xnor2_1 _1610_ (.Y(_0720_),
    .A(_0642_),
    .B(_0643_));
 sg13g2_xnor2_1 _1611_ (.Y(_0721_),
    .A(_0702_),
    .B(_0720_));
 sg13g2_xnor2_1 _1612_ (.Y(_0722_),
    .A(_0719_),
    .B(_0721_));
 sg13g2_nand2_1 _1613_ (.Y(_0723_),
    .A(net98),
    .B(_0557_));
 sg13g2_nand2_1 _1614_ (.Y(_0724_),
    .A(net92),
    .B(_0562_));
 sg13g2_xnor2_1 _1615_ (.Y(_0725_),
    .A(_0723_),
    .B(_0724_));
 sg13g2_xnor2_1 _1616_ (.Y(_0726_),
    .A(_0699_),
    .B(_0725_));
 sg13g2_nand2_1 _1617_ (.Y(_0727_),
    .A(\inp_a[1] ),
    .B(_0557_));
 sg13g2_a22oi_1 _1618_ (.Y(_0728_),
    .B1(_0552_),
    .B2(net98),
    .A2(net106),
    .A1(_0554_));
 sg13g2_nand4_1 _1619_ (.B(_0554_),
    .C(net106),
    .A(net98),
    .Y(_0729_),
    .D(_0552_));
 sg13g2_o21ai_1 _1620_ (.B1(_0729_),
    .Y(_0730_),
    .A1(_0727_),
    .A2(_0728_));
 sg13g2_nand2_1 _1621_ (.Y(_0731_),
    .A(_0564_),
    .B(net101));
 sg13g2_nor2b_1 _1622_ (.A(_0730_),
    .B_N(_0731_),
    .Y(_0732_));
 sg13g2_nand2b_1 _1623_ (.Y(_0733_),
    .B(_0730_),
    .A_N(_0731_));
 sg13g2_o21ai_1 _1624_ (.B1(_0733_),
    .Y(_0734_),
    .A1(_0726_),
    .A2(_0732_));
 sg13g2_nand2_1 _1625_ (.Y(_0735_),
    .A(_0722_),
    .B(_0734_));
 sg13g2_xor2_1 _1626_ (.B(_0559_),
    .A(_0561_),
    .X(_0736_));
 sg13g2_nor3_1 _1627_ (.A(_0607_),
    .B(_0727_),
    .C(_0736_),
    .Y(_0737_));
 sg13g2_xnor2_1 _1628_ (.Y(_0738_),
    .A(_0731_),
    .B(_0730_));
 sg13g2_xnor2_1 _1629_ (.Y(_0739_),
    .A(_0726_),
    .B(_0738_));
 sg13g2_nand2_1 _1630_ (.Y(_0740_),
    .A(_0737_),
    .B(_0739_));
 sg13g2_nor2_1 _1631_ (.A(_0722_),
    .B(_0734_),
    .Y(_0741_));
 sg13g2_a21oi_2 _1632_ (.B1(_0741_),
    .Y(_0742_),
    .A2(_0740_),
    .A1(_0735_));
 sg13g2_nand3_1 _1633_ (.B(_0718_),
    .C(_0742_),
    .A(net37),
    .Y(_0743_));
 sg13g2_nand2_1 _1634_ (.Y(_0744_),
    .A(net87),
    .B(net101));
 sg13g2_a21oi_1 _1635_ (.A1(_0718_),
    .A2(_0742_),
    .Y(_0745_),
    .B1(net37));
 sg13g2_a21oi_1 _1636_ (.A1(_0743_),
    .A2(_0744_),
    .Y(_0746_),
    .B1(_0745_));
 sg13g2_nand2_1 _1637_ (.Y(_0747_),
    .A(_0689_),
    .B(_0746_));
 sg13g2_and2_1 _1638_ (.A(_0578_),
    .B(net101),
    .X(_0748_));
 sg13g2_buf_1 _1639_ (.A(_0748_),
    .X(_0749_));
 sg13g2_a21o_1 _1640_ (.A2(_0703_),
    .A1(_0696_),
    .B1(_0710_),
    .X(_0750_));
 sg13g2_xor2_1 _1641_ (.B(_0640_),
    .A(_0627_),
    .X(_0751_));
 sg13g2_xnor2_1 _1642_ (.Y(_0752_),
    .A(_0751_),
    .B(_0691_));
 sg13g2_a22oi_1 _1643_ (.Y(_0753_),
    .B1(_0750_),
    .B2(_0752_),
    .A2(_0709_),
    .A1(_0707_));
 sg13g2_xnor2_1 _1644_ (.Y(_0754_),
    .A(_0752_),
    .B(_0717_));
 sg13g2_a21o_1 _1645_ (.A2(_0740_),
    .A1(_0735_),
    .B1(_0741_),
    .X(_0755_));
 sg13g2_buf_1 _1646_ (.A(_0755_),
    .X(_0756_));
 sg13g2_nand2_1 _1647_ (.Y(_0757_),
    .A(_0641_),
    .B(_0648_));
 sg13g2_nor2b_1 _1648_ (.A(_0653_),
    .B_N(_0618_),
    .Y(_0758_));
 sg13g2_a21oi_1 _1649_ (.A1(_0751_),
    .A2(_0690_),
    .Y(_0759_),
    .B1(_0618_));
 sg13g2_and3_1 _1650_ (.X(_0760_),
    .A(_0751_),
    .B(_0690_),
    .C(_0618_));
 sg13g2_a221oi_1 _1651_ (.B2(_0654_),
    .C1(_0760_),
    .B1(_0759_),
    .A1(_0757_),
    .Y(_0761_),
    .A2(_0758_));
 sg13g2_xnor2_1 _1652_ (.Y(_0762_),
    .A(_0658_),
    .B(_0761_));
 sg13g2_nor4_1 _1653_ (.A(_0753_),
    .B(_0754_),
    .C(_0756_),
    .D(_0762_),
    .Y(_0763_));
 sg13g2_xor2_1 _1654_ (.B(_0761_),
    .A(_0658_),
    .X(_0764_));
 sg13g2_and4_1 _1655_ (.A(_0718_),
    .B(_0742_),
    .C(_0660_),
    .D(_0764_),
    .X(_0765_));
 sg13g2_a22oi_1 _1656_ (.Y(_0766_),
    .B1(_0765_),
    .B2(_0688_),
    .A2(_0763_),
    .A1(_0749_));
 sg13g2_or4_1 _1657_ (.A(_0754_),
    .B(_0756_),
    .C(_0660_),
    .D(_0762_),
    .X(_0767_));
 sg13g2_nand3_1 _1658_ (.B(_0660_),
    .C(_0764_),
    .A(net37),
    .Y(_0768_));
 sg13g2_mux2_1 _1659_ (.A0(_0767_),
    .A1(_0768_),
    .S(_0688_),
    .X(_0769_));
 sg13g2_nand3b_1 _1660_ (.B(_0764_),
    .C(_0714_),
    .Y(_0770_),
    .A_N(_0660_));
 sg13g2_nand3_1 _1661_ (.B(_0764_),
    .C(_0749_),
    .A(_0660_),
    .Y(_0771_));
 sg13g2_mux2_1 _1662_ (.A0(_0770_),
    .A1(_0771_),
    .S(_0688_),
    .X(_0772_));
 sg13g2_or4_1 _1663_ (.A(_0660_),
    .B(_0688_),
    .C(_0762_),
    .D(_0744_),
    .X(_0773_));
 sg13g2_and4_1 _1664_ (.A(_0766_),
    .B(_0769_),
    .C(_0772_),
    .D(_0773_),
    .X(_0774_));
 sg13g2_buf_1 _1665_ (.A(_0774_),
    .X(_0775_));
 sg13g2_nand2_1 _1666_ (.Y(_0776_),
    .A(_0747_),
    .B(_0775_));
 sg13g2_nor2b_1 _1667_ (.A(net92),
    .B_N(net91),
    .Y(_0777_));
 sg13g2_nand4_1 _1668_ (.B(net99),
    .C(_0570_),
    .A(_0581_),
    .Y(_0778_),
    .D(_0777_));
 sg13g2_inv_1 _1669_ (.Y(_0779_),
    .A(net91));
 sg13g2_nor2b_1 _1670_ (.A(net99),
    .B_N(net103),
    .Y(_0780_));
 sg13g2_a22oi_1 _1671_ (.Y(_0781_),
    .B1(_0639_),
    .B2(_0780_),
    .A2(net92),
    .A1(_0779_));
 sg13g2_a21o_1 _1672_ (.A2(_0781_),
    .A1(_0778_),
    .B1(_0577_),
    .X(_0782_));
 sg13g2_nand3b_1 _1673_ (.B(net92),
    .C(net91),
    .Y(_0783_),
    .A_N(_0575_));
 sg13g2_a21oi_1 _1674_ (.A1(net103),
    .A2(_0783_),
    .Y(_0784_),
    .B1(_0621_));
 sg13g2_nand2_2 _1675_ (.Y(_0785_),
    .A(net103),
    .B(net91));
 sg13g2_a22oi_1 _1676_ (.Y(_0786_),
    .B1(net91),
    .B2(net95),
    .A2(net99),
    .A1(net103));
 sg13g2_o21ai_1 _1677_ (.B1(_0786_),
    .Y(_0787_),
    .A1(_0628_),
    .A2(_0785_));
 sg13g2_nor2b_1 _1678_ (.A(_0784_),
    .B_N(_0787_),
    .Y(_0788_));
 sg13g2_nand2_2 _1679_ (.Y(_0789_),
    .A(_0572_),
    .B(net105));
 sg13g2_nand2_1 _1680_ (.Y(_0790_),
    .A(_0566_),
    .B(net104));
 sg13g2_nand2_1 _1681_ (.Y(_0791_),
    .A(net97),
    .B(net90));
 sg13g2_xor2_1 _1682_ (.B(_0791_),
    .A(_0790_),
    .X(_0792_));
 sg13g2_xor2_1 _1683_ (.B(_0792_),
    .A(_0789_),
    .X(_0793_));
 sg13g2_a21o_1 _1684_ (.A2(_0788_),
    .A1(_0782_),
    .B1(_0793_),
    .X(_0794_));
 sg13g2_nand3_1 _1685_ (.B(_0782_),
    .C(_0788_),
    .A(_0793_),
    .Y(_0795_));
 sg13g2_nand2_1 _1686_ (.Y(_0796_),
    .A(_0794_),
    .B(_0795_));
 sg13g2_nand2_2 _1687_ (.Y(_0797_),
    .A(net99),
    .B(_0575_));
 sg13g2_xnor2_1 _1688_ (.Y(_0798_),
    .A(_0797_),
    .B(_0666_));
 sg13g2_xnor2_1 _1689_ (.Y(_0799_),
    .A(_0644_),
    .B(_0673_));
 sg13g2_a21o_1 _1690_ (.A2(_0799_),
    .A1(_0798_),
    .B1(_0670_),
    .X(_0800_));
 sg13g2_nand2_1 _1691_ (.Y(_0801_),
    .A(_0644_),
    .B(_0671_));
 sg13g2_o21ai_1 _1692_ (.B1(_0672_),
    .Y(_0802_),
    .A1(_0644_),
    .A2(_0671_));
 sg13g2_nand2_1 _1693_ (.Y(_0803_),
    .A(_0801_),
    .B(_0802_));
 sg13g2_a21oi_1 _1694_ (.A1(_0667_),
    .A2(_0674_),
    .Y(_0804_),
    .B1(_0803_));
 sg13g2_and2_1 _1695_ (.A(_0801_),
    .B(_0802_),
    .X(_0805_));
 sg13g2_nor2_1 _1696_ (.A(_0670_),
    .B(_0805_),
    .Y(_0806_));
 sg13g2_nand2_1 _1697_ (.Y(_0807_),
    .A(_0798_),
    .B(_0799_));
 sg13g2_nor3_1 _1698_ (.A(_0798_),
    .B(_0799_),
    .C(_0805_),
    .Y(_0808_));
 sg13g2_a221oi_1 _1699_ (.B2(_0807_),
    .C1(_0808_),
    .B1(_0806_),
    .A1(_0800_),
    .Y(_0809_),
    .A2(_0804_));
 sg13g2_xnor2_1 _1700_ (.Y(_0810_),
    .A(_0796_),
    .B(_0809_));
 sg13g2_xnor2_1 _1701_ (.Y(_0811_),
    .A(_0798_),
    .B(_0675_));
 sg13g2_nand2_1 _1702_ (.Y(_0812_),
    .A(_0678_),
    .B(_0682_));
 sg13g2_and2_1 _1703_ (.A(_0685_),
    .B(_0684_),
    .X(_0813_));
 sg13g2_a221oi_1 _1704_ (.B2(_0812_),
    .C1(_0813_),
    .B1(_0811_),
    .A1(net106),
    .Y(_0814_),
    .A2(_0579_));
 sg13g2_nand2_1 _1705_ (.Y(_0815_),
    .A(_0677_),
    .B(_0625_));
 sg13g2_xnor2_1 _1706_ (.Y(_0816_),
    .A(_0670_),
    .B(_0799_));
 sg13g2_nor2_1 _1707_ (.A(_0798_),
    .B(_0683_),
    .Y(_0817_));
 sg13g2_a22oi_1 _1708_ (.Y(_0818_),
    .B1(_0816_),
    .B2(_0817_),
    .A2(_0685_),
    .A1(_0815_));
 sg13g2_nand3_1 _1709_ (.B(_0675_),
    .C(_0681_),
    .A(_0798_),
    .Y(_0819_));
 sg13g2_nand2_1 _1710_ (.Y(_0820_),
    .A(net106),
    .B(_0579_));
 sg13g2_a221oi_1 _1711_ (.B2(_0819_),
    .C1(_0820_),
    .B1(_0818_),
    .A1(_0676_),
    .Y(_0821_),
    .A2(_0683_));
 sg13g2_or3_1 _1712_ (.A(_0810_),
    .B(_0814_),
    .C(_0821_),
    .X(_0822_));
 sg13g2_o21ai_1 _1713_ (.B1(_0810_),
    .Y(_0823_),
    .A1(_0814_),
    .A2(_0821_));
 sg13g2_a21o_1 _1714_ (.A2(_0687_),
    .A1(_0661_),
    .B1(_0660_),
    .X(_0824_));
 sg13g2_or2_1 _1715_ (.X(_0825_),
    .B(_0687_),
    .A(_0661_));
 sg13g2_a22oi_1 _1716_ (.Y(_0826_),
    .B1(_0824_),
    .B2(_0825_),
    .A2(_0823_),
    .A1(_0822_));
 sg13g2_nand4_1 _1717_ (.B(_0822_),
    .C(_0823_),
    .A(_0825_),
    .Y(_0827_),
    .D(_0824_));
 sg13g2_buf_1 _1718_ (.A(_0827_),
    .X(_0828_));
 sg13g2_nand2b_1 _1719_ (.Y(_0829_),
    .B(_0828_),
    .A_N(_0826_));
 sg13g2_xnor2_1 _1720_ (.Y(_0830_),
    .A(_0776_),
    .B(_0829_));
 sg13g2_nor2_1 _1721_ (.A(_0612_),
    .B(_0830_),
    .Y(_0831_));
 sg13g2_xnor2_1 _1722_ (.Y(_0832_),
    .A(_0598_),
    .B(_0831_));
 sg13g2_buf_1 _1723_ (.A(net93),
    .X(_0833_));
 sg13g2_buf_1 _1724_ (.A(_0604_),
    .X(_0834_));
 sg13g2_inv_1 _1725_ (.Y(_0835_),
    .A(_0590_));
 sg13g2_nand2_1 _1726_ (.Y(_0836_),
    .A(_0586_),
    .B(net82));
 sg13g2_nand3_1 _1727_ (.B(net66),
    .C(_0836_),
    .A(net83),
    .Y(_0837_));
 sg13g2_buf_1 _1728_ (.A(_0837_),
    .X(_0838_));
 sg13g2_buf_1 _1729_ (.A(net57),
    .X(_0839_));
 sg13g2_nor2_2 _1730_ (.A(net53),
    .B(net52),
    .Y(_0840_));
 sg13g2_a22oi_1 _1731_ (.Y(_0841_),
    .B1(_0832_),
    .B2(_0840_),
    .A2(net46),
    .A1(\result[0] ));
 sg13g2_nor2_1 _1732_ (.A(net76),
    .B(_0841_),
    .Y(_0018_));
 sg13g2_buf_1 _1733_ (.A(net53),
    .X(_0842_));
 sg13g2_buf_1 _1734_ (.A(net45),
    .X(_0843_));
 sg13g2_nand2_1 _1735_ (.Y(_0844_),
    .A(\result[10] ),
    .B(net41));
 sg13g2_nand2_1 _1736_ (.Y(_0845_),
    .A(_0004_),
    .B(_0594_));
 sg13g2_buf_1 _1737_ (.A(_0845_),
    .X(_0846_));
 sg13g2_buf_1 _1738_ (.A(net51),
    .X(_0847_));
 sg13g2_buf_1 _1739_ (.A(net57),
    .X(_0848_));
 sg13g2_nor2_2 _1740_ (.A(_0603_),
    .B(_0590_),
    .Y(_0849_));
 sg13g2_buf_1 _1741_ (.A(_0849_),
    .X(_0850_));
 sg13g2_nand2_1 _1742_ (.Y(_0851_),
    .A(net92),
    .B(net107));
 sg13g2_nand2_1 _1743_ (.Y(_0852_),
    .A(_0558_),
    .B(net101));
 sg13g2_xnor2_1 _1744_ (.Y(_0853_),
    .A(_0851_),
    .B(_0852_));
 sg13g2_nor2_1 _1745_ (.A(net93),
    .B(net5),
    .Y(_0854_));
 sg13g2_a21oi_1 _1746_ (.A1(net93),
    .A2(_0853_),
    .Y(_0855_),
    .B1(_0854_));
 sg13g2_nand3b_1 _1747_ (.B(_0747_),
    .C(_0775_),
    .Y(_0856_),
    .A_N(_0826_));
 sg13g2_buf_2 _1748_ (.A(_0856_),
    .X(_0857_));
 sg13g2_a22oi_1 _1749_ (.Y(_0858_),
    .B1(_0818_),
    .B2(_0819_),
    .A2(_0683_),
    .A1(_0676_));
 sg13g2_nand2_1 _1750_ (.Y(_0859_),
    .A(_0810_),
    .B(_0858_));
 sg13g2_o21ai_1 _1751_ (.B1(_0820_),
    .Y(_0860_),
    .A1(_0810_),
    .A2(_0858_));
 sg13g2_nand2_1 _1752_ (.Y(_0861_),
    .A(net105),
    .B(_0578_));
 sg13g2_xnor2_1 _1753_ (.Y(_0862_),
    .A(_0789_),
    .B(_0792_));
 sg13g2_nand3_1 _1754_ (.B(_0782_),
    .C(_0788_),
    .A(_0862_),
    .Y(_0863_));
 sg13g2_buf_1 _1755_ (.A(_0863_),
    .X(_0864_));
 sg13g2_inv_1 _1756_ (.Y(_0865_),
    .A(net99));
 sg13g2_nand2b_1 _1757_ (.Y(_0866_),
    .B(net97),
    .A_N(_0576_));
 sg13g2_mux2_1 _1758_ (.A0(_0577_),
    .A1(_0866_),
    .S(net91),
    .X(_0867_));
 sg13g2_nand4_1 _1759_ (.B(net91),
    .C(net95),
    .A(_0865_),
    .Y(_0868_),
    .D(_0569_));
 sg13g2_o21ai_1 _1760_ (.B1(_0868_),
    .Y(_0869_),
    .A1(_0865_),
    .A2(_0867_));
 sg13g2_nor3_1 _1761_ (.A(_0582_),
    .B(_0797_),
    .C(_0664_),
    .Y(_0870_));
 sg13g2_a21oi_1 _1762_ (.A1(_0665_),
    .A2(_0869_),
    .Y(_0871_),
    .B1(_0870_));
 sg13g2_and2_1 _1763_ (.A(_0575_),
    .B(_0563_),
    .X(_0872_));
 sg13g2_buf_1 _1764_ (.A(_0872_),
    .X(_0873_));
 sg13g2_o21ai_1 _1765_ (.B1(_0873_),
    .Y(_0874_),
    .A1(_0663_),
    .A2(_0785_));
 sg13g2_nand2_2 _1766_ (.Y(_0875_),
    .A(_0575_),
    .B(net90));
 sg13g2_o21ai_1 _1767_ (.B1(_0875_),
    .Y(_0876_),
    .A1(_0663_),
    .A2(_0785_));
 sg13g2_nand2_1 _1768_ (.Y(_0877_),
    .A(net104),
    .B(_0572_));
 sg13g2_nand2_2 _1769_ (.Y(_0878_),
    .A(_0568_),
    .B(_0566_));
 sg13g2_xnor2_1 _1770_ (.Y(_0879_),
    .A(_0877_),
    .B(_0878_));
 sg13g2_mux2_1 _1771_ (.A0(_0874_),
    .A1(_0876_),
    .S(_0879_),
    .X(_0880_));
 sg13g2_buf_1 _1772_ (.A(_0880_),
    .X(_0881_));
 sg13g2_and2_1 _1773_ (.A(net103),
    .B(net98),
    .X(_0882_));
 sg13g2_buf_2 _1774_ (.A(_0882_),
    .X(_0883_));
 sg13g2_nand3_1 _1775_ (.B(_0883_),
    .C(_0875_),
    .A(_0797_),
    .Y(_0884_));
 sg13g2_nand3_1 _1776_ (.B(_0883_),
    .C(_0873_),
    .A(_0797_),
    .Y(_0885_));
 sg13g2_mux2_1 _1777_ (.A0(_0884_),
    .A1(_0885_),
    .S(_0879_),
    .X(_0886_));
 sg13g2_buf_1 _1778_ (.A(_0886_),
    .X(_0887_));
 sg13g2_nand2_1 _1779_ (.Y(_0888_),
    .A(_0789_),
    .B(_0790_));
 sg13g2_o21ai_1 _1780_ (.B1(_0791_),
    .Y(_0889_),
    .A1(_0789_),
    .A2(_0790_));
 sg13g2_nand2_1 _1781_ (.Y(_0890_),
    .A(_0888_),
    .B(_0889_));
 sg13g2_nand3_1 _1782_ (.B(_0887_),
    .C(_0890_),
    .A(_0881_),
    .Y(_0891_));
 sg13g2_a21o_1 _1783_ (.A2(_0887_),
    .A1(_0881_),
    .B1(_0890_),
    .X(_0892_));
 sg13g2_a22oi_1 _1784_ (.Y(_0893_),
    .B1(_0891_),
    .B2(_0892_),
    .A2(net61),
    .A1(net49));
 sg13g2_and4_1 _1785_ (.A(net49),
    .B(net61),
    .C(_0891_),
    .D(_0892_),
    .X(_0894_));
 sg13g2_nor3_1 _1786_ (.A(_0861_),
    .B(_0893_),
    .C(_0894_),
    .Y(_0895_));
 sg13g2_and2_1 _1787_ (.A(net105),
    .B(_0578_),
    .X(_0896_));
 sg13g2_buf_1 _1788_ (.A(_0896_),
    .X(_0897_));
 sg13g2_and2_1 _1789_ (.A(_0888_),
    .B(_0889_),
    .X(_0898_));
 sg13g2_nand3_1 _1790_ (.B(_0887_),
    .C(_0898_),
    .A(_0881_),
    .Y(_0899_));
 sg13g2_buf_2 _1791_ (.A(_0899_),
    .X(_0900_));
 sg13g2_a21o_1 _1792_ (.A2(_0887_),
    .A1(_0881_),
    .B1(_0898_),
    .X(_0901_));
 sg13g2_buf_2 _1793_ (.A(_0901_),
    .X(_0902_));
 sg13g2_and4_1 _1794_ (.A(net49),
    .B(net61),
    .C(_0900_),
    .D(_0902_),
    .X(_0903_));
 sg13g2_a22oi_1 _1795_ (.Y(_0904_),
    .B1(_0900_),
    .B2(_0902_),
    .A2(_0871_),
    .A1(_0864_));
 sg13g2_nor3_1 _1796_ (.A(_0897_),
    .B(_0903_),
    .C(_0904_),
    .Y(_0905_));
 sg13g2_o21ai_1 _1797_ (.B1(_0670_),
    .Y(_0906_),
    .A1(_0798_),
    .A2(_0799_));
 sg13g2_nand2_1 _1798_ (.Y(_0907_),
    .A(_0807_),
    .B(_0906_));
 sg13g2_nand3_1 _1799_ (.B(_0794_),
    .C(_0795_),
    .A(_0803_),
    .Y(_0908_));
 sg13g2_a21oi_1 _1800_ (.A1(_0794_),
    .A2(_0795_),
    .Y(_0909_),
    .B1(_0803_));
 sg13g2_a21oi_1 _1801_ (.A1(_0907_),
    .A2(_0908_),
    .Y(_0910_),
    .B1(_0909_));
 sg13g2_o21ai_1 _1802_ (.B1(_0910_),
    .Y(_0911_),
    .A1(_0895_),
    .A2(_0905_));
 sg13g2_a21o_1 _1803_ (.A2(_0908_),
    .A1(_0907_),
    .B1(_0909_),
    .X(_0912_));
 sg13g2_o21ai_1 _1804_ (.B1(_0897_),
    .Y(_0913_),
    .A1(_0903_),
    .A2(_0904_));
 sg13g2_o21ai_1 _1805_ (.B1(_0861_),
    .Y(_0914_),
    .A1(_0893_),
    .A2(_0894_));
 sg13g2_nand3_1 _1806_ (.B(_0913_),
    .C(_0914_),
    .A(_0912_),
    .Y(_0915_));
 sg13g2_a22oi_1 _1807_ (.Y(_0916_),
    .B1(_0911_),
    .B2(_0915_),
    .A2(_0860_),
    .A1(_0859_));
 sg13g2_nand4_1 _1808_ (.B(_0860_),
    .C(_0911_),
    .A(_0859_),
    .Y(_0917_),
    .D(_0915_));
 sg13g2_nand2b_1 _1809_ (.Y(_0918_),
    .B(_0917_),
    .A_N(_0916_));
 sg13g2_a21oi_1 _1810_ (.A1(_0828_),
    .A2(_0857_),
    .Y(_0919_),
    .B1(_0918_));
 sg13g2_and3_1 _1811_ (.X(_0920_),
    .A(_0828_),
    .B(_0857_),
    .C(_0918_));
 sg13g2_buf_1 _1812_ (.A(_0608_),
    .X(_0921_));
 sg13g2_o21ai_1 _1813_ (.B1(net81),
    .Y(_0922_),
    .A1(_0919_),
    .A2(_0920_));
 sg13g2_buf_1 _1814_ (.A(_0833_),
    .X(_0923_));
 sg13g2_nor2_1 _1815_ (.A(net73),
    .B(_0853_),
    .Y(_0924_));
 sg13g2_nor2_1 _1816_ (.A(net85),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_o21ai_1 _1817_ (.B1(net73),
    .Y(_0926_),
    .A1(_0919_),
    .A2(_0920_));
 sg13g2_a221oi_1 _1818_ (.B2(_0926_),
    .C1(net82),
    .B1(_0925_),
    .A1(net75),
    .Y(_0927_),
    .A2(_0922_));
 sg13g2_a21o_1 _1819_ (.A2(_0855_),
    .A1(net65),
    .B1(_0927_),
    .X(_0928_));
 sg13g2_nor2_1 _1820_ (.A(\ad.a[9] ),
    .B(_0928_),
    .Y(_0929_));
 sg13g2_inv_1 _1821_ (.Y(_0930_),
    .A(_0602_));
 sg13g2_buf_1 _1822_ (.A(_0923_),
    .X(_0931_));
 sg13g2_nor2_1 _1823_ (.A(net64),
    .B(_0607_),
    .Y(_0932_));
 sg13g2_a21oi_1 _1824_ (.A1(net64),
    .A2(_0830_),
    .Y(_0933_),
    .B1(_0932_));
 sg13g2_nor2_1 _1825_ (.A(_0603_),
    .B(net73),
    .Y(_0934_));
 sg13g2_nand2_1 _1826_ (.Y(_0935_),
    .A(_0830_),
    .B(net63));
 sg13g2_o21ai_1 _1827_ (.B1(_0935_),
    .Y(_0936_),
    .A1(net75),
    .A2(_0933_));
 sg13g2_a22oi_1 _1828_ (.Y(_0937_),
    .B1(_0936_),
    .B2(_0592_),
    .A2(net65),
    .A1(_0930_));
 sg13g2_inv_1 _1829_ (.Y(_0938_),
    .A(\ad.a[5] ));
 sg13g2_inv_1 _1830_ (.Y(_0939_),
    .A(\ad.a[6] ));
 sg13g2_nor2_1 _1831_ (.A(_0586_),
    .B(_0835_),
    .Y(_0940_));
 sg13g2_buf_1 _1832_ (.A(_0940_),
    .X(_0941_));
 sg13g2_a221oi_1 _1833_ (.B2(_0752_),
    .C1(_0608_),
    .B1(_0750_),
    .A1(_0707_),
    .Y(_0942_),
    .A2(_0709_));
 sg13g2_o21ai_1 _1834_ (.B1(_0942_),
    .Y(_0943_),
    .A1(_0754_),
    .A2(_0756_));
 sg13g2_nand4_1 _1835_ (.B(net37),
    .C(_0718_),
    .A(net93),
    .Y(_0944_),
    .D(_0742_));
 sg13g2_xnor2_1 _1836_ (.Y(_0945_),
    .A(_0764_),
    .B(_0749_));
 sg13g2_a21o_1 _1837_ (.A2(_0944_),
    .A1(_0943_),
    .B1(_0945_),
    .X(_0946_));
 sg13g2_nand2_1 _1838_ (.Y(_0947_),
    .A(_0718_),
    .B(_0742_));
 sg13g2_nand4_1 _1839_ (.B(net37),
    .C(_0947_),
    .A(net83),
    .Y(_0948_),
    .D(_0945_));
 sg13g2_nor2_1 _1840_ (.A(_0754_),
    .B(_0756_),
    .Y(_0949_));
 sg13g2_nand3_1 _1841_ (.B(_0945_),
    .C(_0942_),
    .A(_0949_),
    .Y(_0950_));
 sg13g2_nand2_1 _1842_ (.Y(_0951_),
    .A(net81),
    .B(net10));
 sg13g2_nand4_1 _1843_ (.B(_0948_),
    .C(_0950_),
    .A(_0946_),
    .Y(_0952_),
    .D(_0951_));
 sg13g2_nand2_1 _1844_ (.Y(_0953_),
    .A(net93),
    .B(net10));
 sg13g2_nor2_1 _1845_ (.A(net84),
    .B(_0953_),
    .Y(_0954_));
 sg13g2_inv_1 _1846_ (.Y(_0955_),
    .A(_0954_));
 sg13g2_a221oi_1 _1847_ (.B2(_0752_),
    .C1(_0609_),
    .B1(_0750_),
    .A1(_0707_),
    .Y(_0956_),
    .A2(_0709_));
 sg13g2_o21ai_1 _1848_ (.B1(_0956_),
    .Y(_0957_),
    .A1(_0754_),
    .A2(_0756_));
 sg13g2_nor2_1 _1849_ (.A(net82),
    .B(net93),
    .Y(_0958_));
 sg13g2_nand4_1 _1850_ (.B(_0714_),
    .C(_0718_),
    .A(net72),
    .Y(_0959_),
    .D(_0742_));
 sg13g2_a21o_1 _1851_ (.A2(_0959_),
    .A1(_0957_),
    .B1(_0945_),
    .X(_0960_));
 sg13g2_nand4_1 _1852_ (.B(net37),
    .C(_0947_),
    .A(net72),
    .Y(_0961_),
    .D(_0945_));
 sg13g2_nand3_1 _1853_ (.B(_0945_),
    .C(_0956_),
    .A(_0949_),
    .Y(_0962_));
 sg13g2_nand4_1 _1854_ (.B(_0960_),
    .C(_0961_),
    .A(_0955_),
    .Y(_0963_),
    .D(_0962_));
 sg13g2_a22oi_1 _1855_ (.Y(_0964_),
    .B1(_0963_),
    .B2(net85),
    .A2(_0952_),
    .A1(net62));
 sg13g2_and2_1 _1856_ (.A(_0939_),
    .B(_0964_),
    .X(_0965_));
 sg13g2_nor2_1 _1857_ (.A(_0939_),
    .B(_0838_),
    .Y(_0966_));
 sg13g2_and2_1 _1858_ (.A(_0859_),
    .B(_0860_),
    .X(_0967_));
 sg13g2_and2_1 _1859_ (.A(_0911_),
    .B(_0915_),
    .X(_0968_));
 sg13g2_a221oi_1 _1860_ (.B2(_0968_),
    .C1(_0826_),
    .B1(_0967_),
    .A1(_0689_),
    .Y(_0969_),
    .A2(_0746_));
 sg13g2_and2_1 _1861_ (.A(_0775_),
    .B(_0969_),
    .X(_0970_));
 sg13g2_nand2_1 _1862_ (.Y(_0971_),
    .A(_0797_),
    .B(_0873_));
 sg13g2_nand2_1 _1863_ (.Y(_0972_),
    .A(_0797_),
    .B(_0875_));
 sg13g2_mux2_1 _1864_ (.A0(_0971_),
    .A1(_0972_),
    .S(_0879_),
    .X(_0973_));
 sg13g2_buf_1 _1865_ (.A(_0973_),
    .X(_0974_));
 sg13g2_nand2_1 _1866_ (.Y(_0975_),
    .A(_0883_),
    .B(_0974_));
 sg13g2_nand2_1 _1867_ (.Y(_0976_),
    .A(_0877_),
    .B(_0878_));
 sg13g2_o21ai_1 _1868_ (.B1(_0875_),
    .Y(_0977_),
    .A1(_0877_),
    .A2(_0878_));
 sg13g2_nand2_2 _1869_ (.Y(_0978_),
    .A(_0976_),
    .B(_0977_));
 sg13g2_nand2_1 _1870_ (.Y(_0979_),
    .A(net97),
    .B(_0572_));
 sg13g2_and2_1 _1871_ (.A(net103),
    .B(net90),
    .X(_0980_));
 sg13g2_nand2_1 _1872_ (.Y(_0981_),
    .A(_0575_),
    .B(_0566_));
 sg13g2_xnor2_1 _1873_ (.Y(_0982_),
    .A(_0980_),
    .B(_0981_));
 sg13g2_xnor2_1 _1874_ (.Y(_0983_),
    .A(_0979_),
    .B(_0982_));
 sg13g2_nand2b_1 _1875_ (.Y(_0984_),
    .B(_0983_),
    .A_N(_0978_));
 sg13g2_nor2b_1 _1876_ (.A(_0983_),
    .B_N(_0978_),
    .Y(_0985_));
 sg13g2_a21oi_2 _1877_ (.B1(_0985_),
    .Y(_0986_),
    .A2(_0984_),
    .A1(_0975_));
 sg13g2_nand2_1 _1878_ (.Y(_0987_),
    .A(net97),
    .B(net87));
 sg13g2_inv_1 _1879_ (.Y(_0988_),
    .A(net88));
 sg13g2_nand2_1 _1880_ (.Y(_0989_),
    .A(_0567_),
    .B(net88));
 sg13g2_or2_1 _1881_ (.X(_0990_),
    .B(net90),
    .A(net97));
 sg13g2_nand3b_1 _1882_ (.B(net90),
    .C(net97),
    .Y(_0991_),
    .A_N(net89));
 sg13g2_o21ai_1 _1883_ (.B1(_0991_),
    .Y(_0992_),
    .A1(_0989_),
    .A2(_0990_));
 sg13g2_a22oi_1 _1884_ (.Y(_0993_),
    .B1(_0992_),
    .B2(net94),
    .A2(_0988_),
    .A1(net90));
 sg13g2_nand2_1 _1885_ (.Y(_0994_),
    .A(net94),
    .B(net88));
 sg13g2_or2_1 _1886_ (.X(_0995_),
    .B(_0994_),
    .A(_0791_));
 sg13g2_a22oi_1 _1887_ (.Y(_0996_),
    .B1(net88),
    .B2(net95),
    .A2(net89),
    .A1(net94));
 sg13g2_nand3b_1 _1888_ (.B(net90),
    .C(net88),
    .Y(_0997_),
    .A_N(net95));
 sg13g2_a21oi_1 _1889_ (.A1(net94),
    .A2(_0997_),
    .Y(_0998_),
    .B1(_0878_));
 sg13g2_a21oi_1 _1890_ (.A1(_0995_),
    .A2(_0996_),
    .Y(_0999_),
    .B1(_0998_));
 sg13g2_o21ai_1 _1891_ (.B1(_0999_),
    .Y(_1000_),
    .A1(_0577_),
    .A2(_0993_));
 sg13g2_nor2_1 _1892_ (.A(_0987_),
    .B(_1000_),
    .Y(_1001_));
 sg13g2_nand2_1 _1893_ (.Y(_1002_),
    .A(_0987_),
    .B(_1000_));
 sg13g2_o21ai_1 _1894_ (.B1(_1002_),
    .Y(_1003_),
    .A1(_0986_),
    .A2(_1001_));
 sg13g2_buf_2 _1895_ (.A(_1003_),
    .X(_1004_));
 sg13g2_nand2b_1 _1896_ (.Y(_1005_),
    .B(net89),
    .A_N(net88));
 sg13g2_nand3b_1 _1897_ (.B(net88),
    .C(net97),
    .Y(_1006_),
    .A_N(net89));
 sg13g2_a21oi_1 _1898_ (.A1(_1005_),
    .A2(_1006_),
    .Y(_1007_),
    .B1(_0577_));
 sg13g2_nor3_1 _1899_ (.A(_0576_),
    .B(_0570_),
    .C(_0989_),
    .Y(_1008_));
 sg13g2_o21ai_1 _1900_ (.B1(_0980_),
    .Y(_1009_),
    .A1(_1007_),
    .A2(_1008_));
 sg13g2_or3_1 _1901_ (.A(net94),
    .B(_0979_),
    .C(_0981_),
    .X(_1010_));
 sg13g2_nand2_1 _1902_ (.Y(_1011_),
    .A(_1009_),
    .B(_1010_));
 sg13g2_nand2_1 _1903_ (.Y(_1012_),
    .A(net95),
    .B(net87));
 sg13g2_nor2_1 _1904_ (.A(net89),
    .B(_0994_),
    .Y(_1013_));
 sg13g2_mux2_1 _1905_ (.A0(net89),
    .A1(_1013_),
    .S(net87),
    .X(_1014_));
 sg13g2_a22oi_1 _1906_ (.Y(_1015_),
    .B1(_1014_),
    .B2(net95),
    .A2(_1012_),
    .A1(_0994_));
 sg13g2_xnor2_1 _1907_ (.Y(_1016_),
    .A(_1011_),
    .B(_1015_));
 sg13g2_xnor2_1 _1908_ (.Y(_1017_),
    .A(_1004_),
    .B(_1016_));
 sg13g2_inv_1 _1909_ (.Y(_1018_),
    .A(net87));
 sg13g2_and2_1 _1910_ (.A(_1009_),
    .B(_1010_),
    .X(_1019_));
 sg13g2_buf_1 _1911_ (.A(_1019_),
    .X(_1020_));
 sg13g2_a21oi_1 _1912_ (.A1(net87),
    .A2(_1020_),
    .Y(_1021_),
    .B1(_0981_));
 sg13g2_a21oi_1 _1913_ (.A1(_1018_),
    .A2(_1011_),
    .Y(_1022_),
    .B1(_1021_));
 sg13g2_o21ai_1 _1914_ (.B1(_0577_),
    .Y(_1023_),
    .A1(_0988_),
    .A2(_1009_));
 sg13g2_o21ai_1 _1915_ (.B1(_1023_),
    .Y(_1024_),
    .A1(_0573_),
    .A2(_1011_));
 sg13g2_nand2_1 _1916_ (.Y(_1025_),
    .A(net87),
    .B(_1024_));
 sg13g2_o21ai_1 _1917_ (.B1(_1025_),
    .Y(_1026_),
    .A1(_0988_),
    .A2(_1022_));
 sg13g2_nor3_1 _1918_ (.A(net94),
    .B(_1020_),
    .C(_1012_),
    .Y(_1027_));
 sg13g2_a21o_1 _1919_ (.A2(_1026_),
    .A1(net94),
    .B1(_1027_),
    .X(_1028_));
 sg13g2_buf_1 _1920_ (.A(_1028_),
    .X(_1029_));
 sg13g2_nand2b_1 _1921_ (.Y(_1030_),
    .B(_1029_),
    .A_N(_1017_));
 sg13g2_and4_1 _1922_ (.A(_0825_),
    .B(_0822_),
    .C(_0823_),
    .D(_0824_),
    .X(_1031_));
 sg13g2_a21o_1 _1923_ (.A2(_0917_),
    .A1(_1031_),
    .B1(_0916_),
    .X(_1032_));
 sg13g2_buf_2 _1924_ (.A(_1032_),
    .X(_1033_));
 sg13g2_and2_1 _1925_ (.A(net49),
    .B(net61),
    .X(_1034_));
 sg13g2_nor2_1 _1926_ (.A(_1034_),
    .B(_0900_),
    .Y(_1035_));
 sg13g2_nand3_1 _1927_ (.B(net61),
    .C(_0900_),
    .A(net49),
    .Y(_1036_));
 sg13g2_buf_1 _1928_ (.A(_1036_),
    .X(_1037_));
 sg13g2_and3_1 _1929_ (.X(_1038_),
    .A(_0897_),
    .B(_0902_),
    .C(_1037_));
 sg13g2_o21ai_1 _1930_ (.B1(_0912_),
    .Y(_1039_),
    .A1(_1035_),
    .A2(_1038_));
 sg13g2_a21oi_2 _1931_ (.B1(_0898_),
    .Y(_1040_),
    .A2(_0887_),
    .A1(_0881_));
 sg13g2_nand2_1 _1932_ (.Y(_1041_),
    .A(_0861_),
    .B(_1040_));
 sg13g2_nand3_1 _1933_ (.B(net61),
    .C(_1040_),
    .A(net49),
    .Y(_1042_));
 sg13g2_nand4_1 _1934_ (.B(net49),
    .C(net61),
    .A(_0861_),
    .Y(_1043_),
    .D(_0900_));
 sg13g2_nand3_1 _1935_ (.B(_1042_),
    .C(_1043_),
    .A(_1041_),
    .Y(_1044_));
 sg13g2_nor2_1 _1936_ (.A(_0897_),
    .B(_1042_),
    .Y(_1045_));
 sg13g2_a221oi_1 _1937_ (.B2(_0910_),
    .C1(_1045_),
    .B1(_1044_),
    .A1(_0897_),
    .Y(_1046_),
    .A2(_1035_));
 sg13g2_nor2_1 _1938_ (.A(_0663_),
    .B(_0875_),
    .Y(_1047_));
 sg13g2_nor2_1 _1939_ (.A(_0663_),
    .B(_0873_),
    .Y(_1048_));
 sg13g2_mux2_1 _1940_ (.A0(_1047_),
    .A1(_1048_),
    .S(_0879_),
    .X(_1049_));
 sg13g2_and2_1 _1941_ (.A(net104),
    .B(_0578_),
    .X(_1050_));
 sg13g2_buf_1 _1942_ (.A(_1050_),
    .X(_1051_));
 sg13g2_o21ai_1 _1943_ (.B1(_1051_),
    .Y(_1052_),
    .A1(_0785_),
    .A2(_1049_));
 sg13g2_nand3_1 _1944_ (.B(_0974_),
    .C(_1051_),
    .A(_0883_),
    .Y(_1053_));
 sg13g2_xnor2_1 _1945_ (.Y(_1054_),
    .A(_0978_),
    .B(_0983_));
 sg13g2_mux2_1 _1946_ (.A0(_1052_),
    .A1(_1053_),
    .S(_1054_),
    .X(_1055_));
 sg13g2_nand2_1 _1947_ (.Y(_1056_),
    .A(net104),
    .B(_0578_));
 sg13g2_nand3_1 _1948_ (.B(_0974_),
    .C(_1056_),
    .A(_0883_),
    .Y(_1057_));
 sg13g2_o21ai_1 _1949_ (.B1(_1056_),
    .Y(_1058_),
    .A1(_0785_),
    .A2(_1049_));
 sg13g2_mux2_1 _1950_ (.A0(_1057_),
    .A1(_1058_),
    .S(_1054_),
    .X(_1059_));
 sg13g2_and2_1 _1951_ (.A(_1055_),
    .B(_1059_),
    .X(_1060_));
 sg13g2_a21oi_1 _1952_ (.A1(_1039_),
    .A2(_1046_),
    .Y(_1061_),
    .B1(_1060_));
 sg13g2_and3_1 _1953_ (.X(_1062_),
    .A(_1060_),
    .B(_1039_),
    .C(_1046_));
 sg13g2_a221oi_1 _1954_ (.B2(_0883_),
    .C1(_0983_),
    .B1(_0974_),
    .A1(_0976_),
    .Y(_1063_),
    .A2(_0977_));
 sg13g2_a21oi_1 _1955_ (.A1(_0902_),
    .A2(_1037_),
    .Y(_1064_),
    .B1(_0986_));
 sg13g2_or2_1 _1956_ (.X(_1065_),
    .B(_1064_),
    .A(_1063_));
 sg13g2_xor2_1 _1957_ (.B(_1000_),
    .A(_0987_),
    .X(_1066_));
 sg13g2_nor2_1 _1958_ (.A(_1051_),
    .B(_1066_),
    .Y(_1067_));
 sg13g2_a21oi_1 _1959_ (.A1(_0883_),
    .A2(_0974_),
    .Y(_1068_),
    .B1(_1051_));
 sg13g2_nor3_1 _1960_ (.A(_1040_),
    .B(_0984_),
    .C(_1068_),
    .Y(_1069_));
 sg13g2_and2_1 _1961_ (.A(_0900_),
    .B(_1063_),
    .X(_1070_));
 sg13g2_and2_1 _1962_ (.A(_1040_),
    .B(_1063_),
    .X(_1071_));
 sg13g2_a221oi_1 _1963_ (.B2(_1034_),
    .C1(_1071_),
    .B1(_1070_),
    .A1(_1037_),
    .Y(_1072_),
    .A2(_1069_));
 sg13g2_nand4_1 _1964_ (.B(net61),
    .C(_0900_),
    .A(net49),
    .Y(_1073_),
    .D(_0978_));
 sg13g2_a21oi_1 _1965_ (.A1(_1040_),
    .A2(_0978_),
    .Y(_1074_),
    .B1(_1053_));
 sg13g2_nand3_1 _1966_ (.B(_1073_),
    .C(_1074_),
    .A(_0983_),
    .Y(_1075_));
 sg13g2_and3_1 _1967_ (.X(_1076_),
    .A(_1066_),
    .B(_1072_),
    .C(_1075_));
 sg13g2_o21ai_1 _1968_ (.B1(_1056_),
    .Y(_1077_),
    .A1(_1063_),
    .A2(_1064_));
 sg13g2_a21oi_1 _1969_ (.A1(_1072_),
    .A2(_1075_),
    .Y(_1078_),
    .B1(_1066_));
 sg13g2_a221oi_1 _1970_ (.B2(_1077_),
    .C1(_1078_),
    .B1(_1076_),
    .A1(_1065_),
    .Y(_1079_),
    .A2(_1067_));
 sg13g2_o21ai_1 _1971_ (.B1(_1079_),
    .Y(_1080_),
    .A1(_1061_),
    .A2(_1062_));
 sg13g2_or3_1 _1972_ (.A(_1030_),
    .B(_1033_),
    .C(_1080_),
    .X(_1081_));
 sg13g2_nand2b_1 _1973_ (.Y(_1082_),
    .B(_0981_),
    .A_N(_0994_));
 sg13g2_a22oi_1 _1974_ (.Y(_1083_),
    .B1(_1012_),
    .B2(_1082_),
    .A2(_1020_),
    .A1(_1004_));
 sg13g2_nor2_1 _1975_ (.A(_1004_),
    .B(_1020_),
    .Y(_1084_));
 sg13g2_nor3_1 _1976_ (.A(net89),
    .B(_0994_),
    .C(_1012_),
    .Y(_1085_));
 sg13g2_nor3_1 _1977_ (.A(_1083_),
    .B(_1084_),
    .C(_1085_),
    .Y(_1086_));
 sg13g2_nand3_1 _1978_ (.B(net89),
    .C(_0573_),
    .A(net95),
    .Y(_1087_));
 sg13g2_a21oi_1 _1979_ (.A1(_1086_),
    .A2(_1087_),
    .Y(_1088_),
    .B1(_1018_));
 sg13g2_nor2b_1 _1980_ (.A(_1017_),
    .B_N(_1029_),
    .Y(_1089_));
 sg13g2_xnor2_1 _1981_ (.Y(_1090_),
    .A(_0975_),
    .B(_1054_));
 sg13g2_and2_1 _1982_ (.A(_0902_),
    .B(_1037_),
    .X(_1091_));
 sg13g2_nor2_1 _1983_ (.A(_1090_),
    .B(_1091_),
    .Y(_1092_));
 sg13g2_a21oi_1 _1984_ (.A1(_1090_),
    .A2(_1091_),
    .Y(_1093_),
    .B1(_1051_));
 sg13g2_nor2_2 _1985_ (.A(_1092_),
    .B(_1093_),
    .Y(_1094_));
 sg13g2_and4_1 _1986_ (.A(_0902_),
    .B(_1037_),
    .C(_1055_),
    .D(_1059_),
    .X(_1095_));
 sg13g2_a22oi_1 _1987_ (.Y(_1096_),
    .B1(_1055_),
    .B2(_1059_),
    .A2(_1037_),
    .A1(_0902_));
 sg13g2_or2_1 _1988_ (.X(_1097_),
    .B(_1096_),
    .A(_1095_));
 sg13g2_buf_1 _1989_ (.A(_1097_),
    .X(_1098_));
 sg13g2_o21ai_1 _1990_ (.B1(_0913_),
    .Y(_1099_),
    .A1(_0910_),
    .A2(_0905_));
 sg13g2_xor2_1 _1991_ (.B(_1066_),
    .A(_0986_),
    .X(_1100_));
 sg13g2_a21o_1 _1992_ (.A2(_1099_),
    .A1(_1098_),
    .B1(_1100_),
    .X(_1101_));
 sg13g2_and3_1 _1993_ (.X(_1102_),
    .A(_1098_),
    .B(_1100_),
    .C(_1099_));
 sg13g2_a21o_1 _1994_ (.A2(_1101_),
    .A1(_1094_),
    .B1(_1102_),
    .X(_1103_));
 sg13g2_a22oi_1 _1995_ (.Y(_1104_),
    .B1(_1089_),
    .B2(_1103_),
    .A2(_1088_),
    .A1(net94));
 sg13g2_o21ai_1 _1996_ (.B1(_1104_),
    .Y(_1105_),
    .A1(_0970_),
    .A2(_1081_));
 sg13g2_buf_1 _1997_ (.A(_1105_),
    .X(_1106_));
 sg13g2_mux2_1 _1998_ (.A0(_0965_),
    .A1(_0966_),
    .S(net36),
    .X(_1107_));
 sg13g2_nand3_1 _1999_ (.B(_0838_),
    .C(_0964_),
    .A(_0939_),
    .Y(_1108_));
 sg13g2_o21ai_1 _2000_ (.B1(_1108_),
    .Y(_1109_),
    .A1(_0939_),
    .A2(_0964_));
 sg13g2_inv_1 _2001_ (.Y(_1110_),
    .A(\ad.a[7] ));
 sg13g2_nor2_1 _2002_ (.A(_0603_),
    .B(net82),
    .Y(_1111_));
 sg13g2_nand3_1 _2003_ (.B(_0689_),
    .C(_1111_),
    .A(_0921_),
    .Y(_1112_));
 sg13g2_nand3_1 _2004_ (.B(net62),
    .C(_0689_),
    .A(net83),
    .Y(_1113_));
 sg13g2_nor2_1 _2005_ (.A(net37),
    .B(_0749_),
    .Y(_1114_));
 sg13g2_o21ai_1 _2006_ (.B1(_0762_),
    .Y(_1115_),
    .A1(_0753_),
    .A2(_0744_));
 sg13g2_nand2b_1 _2007_ (.Y(_1116_),
    .B(_1115_),
    .A_N(_1114_));
 sg13g2_nor4_1 _2008_ (.A(_0753_),
    .B(_0947_),
    .C(_0762_),
    .D(_0744_),
    .Y(_1117_));
 sg13g2_a221oi_1 _2009_ (.B2(_0947_),
    .C1(_1117_),
    .B1(_1116_),
    .A1(_0762_),
    .Y(_1118_),
    .A2(_1114_));
 sg13g2_a21o_1 _2010_ (.A2(_1113_),
    .A1(_1112_),
    .B1(_1118_),
    .X(_1119_));
 sg13g2_nand2_2 _2011_ (.Y(_1120_),
    .A(net85),
    .B(_0590_));
 sg13g2_nor3_1 _2012_ (.A(net83),
    .B(_0689_),
    .C(_1120_),
    .Y(_1121_));
 sg13g2_nor3_1 _2013_ (.A(net81),
    .B(net66),
    .C(_0689_),
    .Y(_1122_));
 sg13g2_o21ai_1 _2014_ (.B1(_1118_),
    .Y(_1123_),
    .A1(_1121_),
    .A2(_1122_));
 sg13g2_and2_1 _2015_ (.A(net83),
    .B(net11),
    .X(_1124_));
 sg13g2_nor2b_1 _2016_ (.A(net83),
    .B_N(net11),
    .Y(_1125_));
 sg13g2_a22oi_1 _2017_ (.Y(_1126_),
    .B1(_1125_),
    .B2(_0941_),
    .A2(_1124_),
    .A1(_0849_));
 sg13g2_and3_1 _2018_ (.X(_1127_),
    .A(_1119_),
    .B(_1123_),
    .C(_1126_));
 sg13g2_xnor2_1 _2019_ (.Y(_1128_),
    .A(_1110_),
    .B(_1127_));
 sg13g2_nor4_1 _2020_ (.A(_0938_),
    .B(_1107_),
    .C(_1109_),
    .D(_1128_),
    .Y(_1129_));
 sg13g2_inv_1 _2021_ (.Y(_1130_),
    .A(\ad.a[4] ));
 sg13g2_nor3_2 _2022_ (.A(_0608_),
    .B(_0940_),
    .C(_0849_),
    .Y(_1131_));
 sg13g2_nor2_2 _2023_ (.A(_1061_),
    .B(_1062_),
    .Y(_1132_));
 sg13g2_nand3_1 _2024_ (.B(_1131_),
    .C(_1132_),
    .A(\ad.a[2] ),
    .Y(_1133_));
 sg13g2_or3_1 _2025_ (.A(_0970_),
    .B(_1033_),
    .C(_1133_),
    .X(_1134_));
 sg13g2_inv_1 _2026_ (.Y(_1135_),
    .A(\ad.a[2] ));
 sg13g2_nor3_1 _2027_ (.A(_1135_),
    .B(_0837_),
    .C(_1132_),
    .Y(_1136_));
 sg13g2_nand2_1 _2028_ (.Y(_1137_),
    .A(_0970_),
    .B(_1136_));
 sg13g2_nand2_1 _2029_ (.Y(_1138_),
    .A(net101),
    .B(_0777_));
 sg13g2_nand3b_1 _2030_ (.B(_0559_),
    .C(net92),
    .Y(_1139_),
    .A_N(_0553_));
 sg13g2_a21oi_1 _2031_ (.A1(_1138_),
    .A2(_1139_),
    .Y(_1140_),
    .B1(_0727_));
 sg13g2_inv_1 _2032_ (.Y(_1141_),
    .A(_0728_));
 sg13g2_a21oi_1 _2033_ (.A1(net92),
    .A2(net101),
    .Y(_1142_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2034_ (.B1(_0729_),
    .Y(_1143_),
    .A1(_1141_),
    .A2(_1142_));
 sg13g2_nor2_1 _2035_ (.A(_1140_),
    .B(_1143_),
    .Y(_1144_));
 sg13g2_nand2_1 _2036_ (.Y(_1145_),
    .A(_0599_),
    .B(net6));
 sg13g2_nor2_1 _2037_ (.A(net84),
    .B(_1145_),
    .Y(_1146_));
 sg13g2_a21oi_1 _2038_ (.A1(net72),
    .A2(_1144_),
    .Y(_1147_),
    .B1(_1146_));
 sg13g2_mux2_1 _2039_ (.A0(net6),
    .A1(_1144_),
    .S(net83),
    .X(_1148_));
 sg13g2_nand2_1 _2040_ (.Y(_1149_),
    .A(_0941_),
    .B(_1148_));
 sg13g2_o21ai_1 _2041_ (.B1(_1149_),
    .Y(_1150_),
    .A1(_0603_),
    .A2(_1147_));
 sg13g2_a22oi_1 _2042_ (.Y(_1151_),
    .B1(_1136_),
    .B2(_1033_),
    .A2(_1150_),
    .A1(\ad.a[2] ));
 sg13g2_nand3_1 _2043_ (.B(_1137_),
    .C(_1151_),
    .A(_1134_),
    .Y(_1152_));
 sg13g2_inv_1 _2044_ (.Y(_1153_),
    .A(\ad.a[1] ));
 sg13g2_and2_1 _2045_ (.A(_0598_),
    .B(_1131_),
    .X(_1154_));
 sg13g2_o21ai_1 _2046_ (.B1(_1154_),
    .Y(_1155_),
    .A1(_0826_),
    .A2(_1031_));
 sg13g2_a21oi_1 _2047_ (.A1(_0747_),
    .A2(_0775_),
    .Y(_1156_),
    .B1(_1155_));
 sg13g2_and2_1 _2048_ (.A(_0689_),
    .B(_0746_),
    .X(_1157_));
 sg13g2_nand4_1 _2049_ (.B(_0769_),
    .C(_0772_),
    .A(_0766_),
    .Y(_1158_),
    .D(_0773_));
 sg13g2_nand2_1 _2050_ (.Y(_1159_),
    .A(_0598_),
    .B(_1131_));
 sg13g2_nor4_2 _2051_ (.A(_1157_),
    .B(_1158_),
    .C(_0829_),
    .Y(_1160_),
    .D(_1159_));
 sg13g2_and2_1 _2052_ (.A(_0598_),
    .B(_0612_),
    .X(_1161_));
 sg13g2_nor3_2 _2053_ (.A(_1156_),
    .B(_1160_),
    .C(_1161_),
    .Y(_1162_));
 sg13g2_nand2_1 _2054_ (.Y(_1163_),
    .A(_0599_),
    .B(net5));
 sg13g2_nand2b_1 _2055_ (.Y(_1164_),
    .B(net82),
    .A_N(_1163_));
 sg13g2_o21ai_1 _2056_ (.B1(_1164_),
    .Y(_1165_),
    .A1(_0609_),
    .A2(_0853_));
 sg13g2_a22oi_1 _2057_ (.Y(_1166_),
    .B1(_1165_),
    .B2(net85),
    .A2(_0855_),
    .A1(net62));
 sg13g2_inv_1 _2058_ (.Y(_1167_),
    .A(_1166_));
 sg13g2_nor4_1 _2059_ (.A(_1156_),
    .B(_1160_),
    .C(_1161_),
    .D(_1167_),
    .Y(_1168_));
 sg13g2_o21ai_1 _2060_ (.B1(_0828_),
    .Y(_1169_),
    .A1(_1157_),
    .A2(_1158_));
 sg13g2_nor3_1 _2061_ (.A(_0826_),
    .B(_0837_),
    .C(_0918_),
    .Y(_1170_));
 sg13g2_and3_1 _2062_ (.X(_1171_),
    .A(_0828_),
    .B(_1131_),
    .C(_0918_));
 sg13g2_a22oi_1 _2063_ (.Y(_1172_),
    .B1(_1171_),
    .B2(_0857_),
    .A2(_1170_),
    .A1(_1169_));
 sg13g2_nand2_1 _2064_ (.Y(_1173_),
    .A(_1153_),
    .B(_1166_));
 sg13g2_a221oi_1 _2065_ (.B2(_0857_),
    .C1(_1173_),
    .B1(_1171_),
    .A1(_1169_),
    .Y(_1174_),
    .A2(_1170_));
 sg13g2_a221oi_1 _2066_ (.B2(_1172_),
    .C1(_1174_),
    .B1(_1168_),
    .A1(_1153_),
    .Y(_1175_),
    .A2(_1162_));
 sg13g2_or2_1 _2067_ (.X(_1176_),
    .B(_1175_),
    .A(_1152_));
 sg13g2_nor3_1 _2068_ (.A(_1031_),
    .B(_0918_),
    .C(_1132_),
    .Y(_1177_));
 sg13g2_nand2_1 _2069_ (.Y(_1178_),
    .A(_0859_),
    .B(_0860_));
 sg13g2_or3_1 _2070_ (.A(_0895_),
    .B(_1095_),
    .C(_1096_),
    .X(_1179_));
 sg13g2_a22oi_1 _2071_ (.Y(_1180_),
    .B1(_1179_),
    .B2(_0912_),
    .A2(_1098_),
    .A1(_0914_));
 sg13g2_nand2_1 _2072_ (.Y(_1181_),
    .A(_1098_),
    .B(_1099_));
 sg13g2_o21ai_1 _2073_ (.B1(_1181_),
    .Y(_1182_),
    .A1(_1178_),
    .A2(_1180_));
 sg13g2_xor2_1 _2074_ (.B(_0739_),
    .A(_0737_),
    .X(_1183_));
 sg13g2_and2_1 _2075_ (.A(_0608_),
    .B(_1183_),
    .X(_1184_));
 sg13g2_nand2_1 _2076_ (.Y(_1185_),
    .A(_0603_),
    .B(net82));
 sg13g2_o21ai_1 _2077_ (.B1(_1185_),
    .Y(_1186_),
    .A1(_1120_),
    .A2(_1184_));
 sg13g2_a21o_1 _2078_ (.A2(_1067_),
    .A1(_1065_),
    .B1(_1078_),
    .X(_1187_));
 sg13g2_a21o_1 _2079_ (.A2(_1076_),
    .A1(_1077_),
    .B1(_1187_),
    .X(_1188_));
 sg13g2_nand3b_1 _2080_ (.B(_1186_),
    .C(_1188_),
    .Y(_1189_),
    .A_N(_1182_));
 sg13g2_a21o_1 _2081_ (.A2(_1177_),
    .A1(_0857_),
    .B1(_1189_),
    .X(_1190_));
 sg13g2_and2_1 _2082_ (.A(_1079_),
    .B(_1186_),
    .X(_1191_));
 sg13g2_nand3_1 _2083_ (.B(_1177_),
    .C(_1191_),
    .A(_0857_),
    .Y(_1192_));
 sg13g2_inv_1 _2084_ (.Y(_1193_),
    .A(net7));
 sg13g2_nand2_1 _2085_ (.Y(_1194_),
    .A(_0587_),
    .B(_1183_));
 sg13g2_o21ai_1 _2086_ (.B1(_1194_),
    .Y(_1195_),
    .A1(_0587_),
    .A2(_1193_));
 sg13g2_nand2_1 _2087_ (.Y(_1196_),
    .A(net72),
    .B(_1195_));
 sg13g2_a21oi_1 _2088_ (.A1(_1193_),
    .A2(_0849_),
    .Y(_1197_),
    .B1(net81));
 sg13g2_o21ai_1 _2089_ (.B1(_1197_),
    .Y(_1198_),
    .A1(net66),
    .A2(_1183_));
 sg13g2_a22oi_1 _2090_ (.Y(_1199_),
    .B1(_1182_),
    .B2(_1191_),
    .A2(_1198_),
    .A1(_1196_));
 sg13g2_nand3_1 _2091_ (.B(_1192_),
    .C(_1199_),
    .A(_1190_),
    .Y(_1200_));
 sg13g2_a21oi_1 _2092_ (.A1(_0775_),
    .A2(_0969_),
    .Y(_1201_),
    .B1(_1033_));
 sg13g2_xnor2_1 _2093_ (.Y(_1202_),
    .A(_1132_),
    .B(_1201_));
 sg13g2_or2_1 _2094_ (.X(_1203_),
    .B(_1150_),
    .A(\ad.a[2] ));
 sg13g2_a21oi_2 _2095_ (.B1(_1203_),
    .Y(_1204_),
    .A2(_1202_),
    .A1(_1131_));
 sg13g2_nor2_1 _2096_ (.A(_1200_),
    .B(_1204_),
    .Y(_1205_));
 sg13g2_inv_1 _2097_ (.Y(_1206_),
    .A(net8));
 sg13g2_xor2_1 _2098_ (.B(_0734_),
    .A(_0722_),
    .X(_1207_));
 sg13g2_xnor2_1 _2099_ (.Y(_1208_),
    .A(_0740_),
    .B(_1207_));
 sg13g2_nand2_1 _2100_ (.Y(_1209_),
    .A(net85),
    .B(_1208_));
 sg13g2_o21ai_1 _2101_ (.B1(_1209_),
    .Y(_1210_),
    .A1(net85),
    .A2(_1206_));
 sg13g2_nand2_1 _2102_ (.Y(_1211_),
    .A(net72),
    .B(_1210_));
 sg13g2_a21o_1 _2103_ (.A2(_0969_),
    .A1(_0775_),
    .B1(_1033_),
    .X(_1212_));
 sg13g2_a21oi_2 _2104_ (.B1(_1102_),
    .Y(_1213_),
    .A2(_1101_),
    .A1(_1094_));
 sg13g2_and3_1 _2105_ (.X(_1214_),
    .A(_1111_),
    .B(_1017_),
    .C(_1213_));
 sg13g2_o21ai_1 _2106_ (.B1(_1214_),
    .Y(_1215_),
    .A1(_1080_),
    .A2(_1212_));
 sg13g2_nor2_1 _2107_ (.A(_1132_),
    .B(_1188_),
    .Y(_1216_));
 sg13g2_nor2_1 _2108_ (.A(_1120_),
    .B(_1017_),
    .Y(_1217_));
 sg13g2_nand3_1 _2109_ (.B(_1201_),
    .C(_1217_),
    .A(_1216_),
    .Y(_1218_));
 sg13g2_a22oi_1 _2110_ (.Y(_1219_),
    .B1(_1103_),
    .B2(_1217_),
    .A2(net65),
    .A1(_1206_));
 sg13g2_nand3_1 _2111_ (.B(_1218_),
    .C(_1219_),
    .A(_1215_),
    .Y(_1220_));
 sg13g2_nor2_1 _2112_ (.A(net84),
    .B(_1017_),
    .Y(_1221_));
 sg13g2_nand3_1 _2113_ (.B(_1080_),
    .C(_1221_),
    .A(_1213_),
    .Y(_1222_));
 sg13g2_nand3_1 _2114_ (.B(_1033_),
    .C(_1221_),
    .A(_1213_),
    .Y(_1223_));
 sg13g2_nand4_1 _2115_ (.B(_1213_),
    .C(_0969_),
    .A(_0775_),
    .Y(_1224_),
    .D(_1221_));
 sg13g2_nand3_1 _2116_ (.B(_1223_),
    .C(_1224_),
    .A(_1222_),
    .Y(_1225_));
 sg13g2_nand2_1 _2117_ (.Y(_1226_),
    .A(_0835_),
    .B(_1017_));
 sg13g2_nor2_1 _2118_ (.A(_1213_),
    .B(_1226_),
    .Y(_1227_));
 sg13g2_nor4_1 _2119_ (.A(_0970_),
    .B(_1033_),
    .C(_1080_),
    .D(_1226_),
    .Y(_1228_));
 sg13g2_nor3_1 _2120_ (.A(_1225_),
    .B(_1227_),
    .C(_1228_),
    .Y(_1229_));
 sg13g2_a221oi_1 _2121_ (.B2(_0591_),
    .C1(net85),
    .B1(_1208_),
    .A1(net8),
    .Y(_1230_),
    .A2(net72));
 sg13g2_a21oi_1 _2122_ (.A1(_0591_),
    .A2(_1210_),
    .Y(_1231_),
    .B1(_0833_));
 sg13g2_a221oi_1 _2123_ (.B2(_1230_),
    .C1(_1231_),
    .B1(_1229_),
    .A1(_1211_),
    .Y(_1232_),
    .A2(_1220_));
 sg13g2_buf_1 _2124_ (.A(_1232_),
    .X(_1233_));
 sg13g2_a21oi_1 _2125_ (.A1(_1176_),
    .A2(_1205_),
    .Y(_1234_),
    .B1(_1233_));
 sg13g2_nand3_1 _2126_ (.B(_1176_),
    .C(_1205_),
    .A(_1233_),
    .Y(_1235_));
 sg13g2_o21ai_1 _2127_ (.B1(_1235_),
    .Y(_1236_),
    .A1(_1130_),
    .A2(_1234_));
 sg13g2_a21o_1 _2128_ (.A2(_1177_),
    .A1(_0857_),
    .B1(_1182_),
    .X(_1237_));
 sg13g2_o21ai_1 _2129_ (.B1(_1100_),
    .Y(_1238_),
    .A1(_1094_),
    .A2(_1237_));
 sg13g2_nand2_1 _2130_ (.Y(_1239_),
    .A(_1094_),
    .B(_1237_));
 sg13g2_a221oi_1 _2131_ (.B2(_1239_),
    .C1(_1029_),
    .B1(_1238_),
    .A1(_1004_),
    .Y(_1240_),
    .A2(_1016_));
 sg13g2_a21oi_1 _2132_ (.A1(_1216_),
    .A2(_1201_),
    .Y(_1241_),
    .B1(_1103_));
 sg13g2_nand3_1 _2133_ (.B(_1029_),
    .C(_1241_),
    .A(_1016_),
    .Y(_1242_));
 sg13g2_nand3_1 _2134_ (.B(_1029_),
    .C(_1241_),
    .A(_1004_),
    .Y(_1243_));
 sg13g2_and2_1 _2135_ (.A(_1004_),
    .B(_1016_),
    .X(_1244_));
 sg13g2_nor3_1 _2136_ (.A(_1004_),
    .B(_1016_),
    .C(_1029_),
    .Y(_1245_));
 sg13g2_a21oi_1 _2137_ (.A1(_1029_),
    .A2(_1244_),
    .Y(_1246_),
    .B1(_1245_));
 sg13g2_nand3_1 _2138_ (.B(_1243_),
    .C(_1246_),
    .A(_1242_),
    .Y(_1247_));
 sg13g2_nor2_1 _2139_ (.A(net81),
    .B(_1120_),
    .Y(_1248_));
 sg13g2_o21ai_1 _2140_ (.B1(_1248_),
    .Y(_1249_),
    .A1(_1240_),
    .A2(_1247_));
 sg13g2_nor2_1 _2141_ (.A(net81),
    .B(_1185_),
    .Y(_1250_));
 sg13g2_o21ai_1 _2142_ (.B1(_1250_),
    .Y(_1251_),
    .A1(_1240_),
    .A2(_1247_));
 sg13g2_nor2b_1 _2143_ (.A(net73),
    .B_N(net9),
    .Y(_1252_));
 sg13g2_xnor2_1 _2144_ (.Y(_1253_),
    .A(_0718_),
    .B(_0756_));
 sg13g2_inv_1 _2145_ (.Y(_1254_),
    .A(_1253_));
 sg13g2_nor2_1 _2146_ (.A(net81),
    .B(_1254_),
    .Y(_1255_));
 sg13g2_o21ai_1 _2147_ (.B1(net62),
    .Y(_1256_),
    .A1(_1252_),
    .A2(_1255_));
 sg13g2_nand2_1 _2148_ (.Y(_1257_),
    .A(net83),
    .B(net9));
 sg13g2_nor2_1 _2149_ (.A(net84),
    .B(_1257_),
    .Y(_1258_));
 sg13g2_nor2_1 _2150_ (.A(_0609_),
    .B(_1254_),
    .Y(_1259_));
 sg13g2_o21ai_1 _2151_ (.B1(net75),
    .Y(_1260_),
    .A1(_1258_),
    .A2(_1259_));
 sg13g2_nand4_1 _2152_ (.B(_1251_),
    .C(_1256_),
    .A(_1249_),
    .Y(_1261_),
    .D(_1260_));
 sg13g2_buf_2 _2153_ (.A(_1261_),
    .X(_1262_));
 sg13g2_nor3_1 _2154_ (.A(_1107_),
    .B(_1109_),
    .C(_1128_),
    .Y(_1263_));
 sg13g2_nor2_1 _2155_ (.A(\ad.a[4] ),
    .B(_1233_),
    .Y(_1264_));
 sg13g2_and3_1 _2156_ (.X(_1265_),
    .A(_1190_),
    .B(_1192_),
    .C(_1199_));
 sg13g2_or3_1 _2157_ (.A(_1152_),
    .B(_1175_),
    .C(_1265_),
    .X(_1266_));
 sg13g2_buf_1 _2158_ (.A(_1266_),
    .X(_1267_));
 sg13g2_inv_1 _2159_ (.Y(_1268_),
    .A(\ad.a[3] ));
 sg13g2_a21oi_2 _2160_ (.B1(_1268_),
    .Y(_1269_),
    .A2(_1204_),
    .A1(_1200_));
 sg13g2_nand3_1 _2161_ (.B(_1267_),
    .C(_1269_),
    .A(_1129_),
    .Y(_1270_));
 sg13g2_nand3_1 _2162_ (.B(_1123_),
    .C(_1126_),
    .A(_1119_),
    .Y(_1271_));
 sg13g2_buf_1 _2163_ (.A(_1131_),
    .X(_1272_));
 sg13g2_nand2_1 _2164_ (.Y(_1273_),
    .A(net60),
    .B(net36));
 sg13g2_a221oi_1 _2165_ (.B2(_1110_),
    .C1(_0939_),
    .B1(_1127_),
    .A1(_0964_),
    .Y(_1274_),
    .A2(_1273_));
 sg13g2_a21oi_1 _2166_ (.A1(\ad.a[7] ),
    .A2(_1271_),
    .Y(_1275_),
    .B1(_1274_));
 sg13g2_o21ai_1 _2167_ (.B1(_1275_),
    .Y(_1276_),
    .A1(_1264_),
    .A2(_1270_));
 sg13g2_a221oi_1 _2168_ (.B2(_1263_),
    .C1(_1276_),
    .B1(_1262_),
    .A1(_1129_),
    .Y(_1277_),
    .A2(_1236_));
 sg13g2_and3_1 _2169_ (.X(_1278_),
    .A(_1233_),
    .B(_1267_),
    .C(_1269_));
 sg13g2_and3_1 _2170_ (.X(_1279_),
    .A(\ad.a[4] ),
    .B(_1267_),
    .C(_1269_));
 sg13g2_nand2_1 _2171_ (.Y(_1280_),
    .A(_0938_),
    .B(_1275_));
 sg13g2_nor4_2 _2172_ (.A(_1236_),
    .B(_1278_),
    .C(_1279_),
    .Y(_1281_),
    .D(_1280_));
 sg13g2_or2_1 _2173_ (.X(_1282_),
    .B(_1281_),
    .A(_1277_));
 sg13g2_nor3_1 _2174_ (.A(_0937_),
    .B(_1277_),
    .C(_1281_),
    .Y(_1283_));
 sg13g2_nor2_1 _2175_ (.A(\ad.a[8] ),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_a21oi_2 _2176_ (.B1(_1284_),
    .Y(_1285_),
    .A2(_1282_),
    .A1(_0937_));
 sg13g2_and2_1 _2177_ (.A(\ad.a[9] ),
    .B(_0928_),
    .X(_1286_));
 sg13g2_buf_1 _2178_ (.A(_1286_),
    .X(_1287_));
 sg13g2_nor2_1 _2179_ (.A(_1285_),
    .B(_1287_),
    .Y(_1288_));
 sg13g2_nor2_1 _2180_ (.A(_0929_),
    .B(_1288_),
    .Y(_1289_));
 sg13g2_nor3_1 _2181_ (.A(_0923_),
    .B(_1140_),
    .C(_1143_),
    .Y(_1290_));
 sg13g2_a21oi_1 _2182_ (.A1(net64),
    .A2(_1202_),
    .Y(_1291_),
    .B1(_1290_));
 sg13g2_nand2_1 _2183_ (.Y(_1292_),
    .A(net63),
    .B(_1202_));
 sg13g2_o21ai_1 _2184_ (.B1(_1292_),
    .Y(_1293_),
    .A1(_0588_),
    .A2(_1291_));
 sg13g2_a22oi_1 _2185_ (.Y(_1294_),
    .B1(_1293_),
    .B2(net74),
    .A2(_1148_),
    .A1(net65));
 sg13g2_inv_1 _2186_ (.Y(_1295_),
    .A(_1294_));
 sg13g2_nor2_1 _2187_ (.A(_1289_),
    .B(_1295_),
    .Y(_1296_));
 sg13g2_nand2_1 _2188_ (.Y(_1297_),
    .A(_1289_),
    .B(_1295_));
 sg13g2_nor2b_1 _2189_ (.A(_1296_),
    .B_N(_1297_),
    .Y(_1298_));
 sg13g2_xnor2_1 _2190_ (.Y(_1299_),
    .A(\ad.a[10] ),
    .B(_1298_));
 sg13g2_nand2_1 _2191_ (.Y(_1300_),
    .A(\result[2] ),
    .B(net52));
 sg13g2_o21ai_1 _2192_ (.B1(_1300_),
    .Y(_1301_),
    .A1(net50),
    .A2(_1299_));
 sg13g2_nand2_1 _2193_ (.Y(_1302_),
    .A(net44),
    .B(_1301_));
 sg13g2_buf_1 _2194_ (.A(_0583_),
    .X(_1303_));
 sg13g2_a21oi_1 _2195_ (.A1(_0844_),
    .A2(_1302_),
    .Y(_0019_),
    .B1(net80));
 sg13g2_buf_1 _2196_ (.A(net45),
    .X(_1304_));
 sg13g2_inv_1 _2197_ (.Y(_1305_),
    .A(\ad.a[11] ));
 sg13g2_nand2_1 _2198_ (.Y(_1306_),
    .A(net73),
    .B(_1183_));
 sg13g2_o21ai_1 _2199_ (.B1(_1306_),
    .Y(_1307_),
    .A1(net73),
    .A2(_1193_));
 sg13g2_xnor2_1 _2200_ (.Y(_1308_),
    .A(_1079_),
    .B(_1237_));
 sg13g2_inv_1 _2201_ (.Y(_1309_),
    .A(_1184_));
 sg13g2_o21ai_1 _2202_ (.B1(_1309_),
    .Y(_1310_),
    .A1(net81),
    .A2(_1308_));
 sg13g2_nor3_1 _2203_ (.A(net73),
    .B(_1120_),
    .C(_1308_),
    .Y(_1311_));
 sg13g2_a221oi_1 _2204_ (.B2(net62),
    .C1(_1311_),
    .B1(_1310_),
    .A1(net65),
    .Y(_1312_),
    .A2(_1307_));
 sg13g2_buf_1 _2205_ (.A(_1312_),
    .X(_1313_));
 sg13g2_xnor2_1 _2206_ (.Y(_1314_),
    .A(_1305_),
    .B(_1313_));
 sg13g2_inv_1 _2207_ (.Y(_1315_),
    .A(\ad.a[10] ));
 sg13g2_a21oi_1 _2208_ (.A1(_1315_),
    .A2(_1297_),
    .Y(_1316_),
    .B1(_1296_));
 sg13g2_xnor2_1 _2209_ (.Y(_1317_),
    .A(_1314_),
    .B(_1316_));
 sg13g2_nand2_1 _2210_ (.Y(_1318_),
    .A(net60),
    .B(_1317_));
 sg13g2_nand2_1 _2211_ (.Y(_1319_),
    .A(\result[3] ),
    .B(net52));
 sg13g2_buf_1 _2212_ (.A(net53),
    .X(_1320_));
 sg13g2_a21oi_1 _2213_ (.A1(_1318_),
    .A2(_1319_),
    .Y(_1321_),
    .B1(net43));
 sg13g2_a21oi_1 _2214_ (.A1(\result[11] ),
    .A2(net40),
    .Y(_1322_),
    .B1(_1321_));
 sg13g2_nor2_1 _2215_ (.A(net76),
    .B(_1322_),
    .Y(_0020_));
 sg13g2_nand2_1 _2216_ (.Y(_1323_),
    .A(\result[12] ),
    .B(net41));
 sg13g2_xnor2_1 _2217_ (.Y(_1324_),
    .A(_1017_),
    .B(_1241_));
 sg13g2_nor2_1 _2218_ (.A(net64),
    .B(_1324_),
    .Y(_1325_));
 sg13g2_buf_1 _2219_ (.A(_0921_),
    .X(_1326_));
 sg13g2_nand2_1 _2220_ (.Y(_1327_),
    .A(net71),
    .B(_1208_));
 sg13g2_o21ai_1 _2221_ (.B1(_1327_),
    .Y(_1328_),
    .A1(net71),
    .A2(_1324_));
 sg13g2_nor2_1 _2222_ (.A(net73),
    .B(_1206_),
    .Y(_1329_));
 sg13g2_a21oi_1 _2223_ (.A1(net64),
    .A2(_1208_),
    .Y(_1330_),
    .B1(_1329_));
 sg13g2_nor2_1 _2224_ (.A(_0836_),
    .B(_1330_),
    .Y(_1331_));
 sg13g2_a221oi_1 _2225_ (.B2(net62),
    .C1(_1331_),
    .B1(_1328_),
    .A1(_1111_),
    .Y(_1332_),
    .A2(_1325_));
 sg13g2_xnor2_1 _2226_ (.Y(_1333_),
    .A(\ad.a[12] ),
    .B(_1332_));
 sg13g2_nand2_1 _2227_ (.Y(_1334_),
    .A(_1305_),
    .B(_1313_));
 sg13g2_nand2_1 _2228_ (.Y(_1335_),
    .A(_1315_),
    .B(_1294_));
 sg13g2_a21o_1 _2229_ (.A2(_1285_),
    .A1(_0928_),
    .B1(\ad.a[9] ),
    .X(_1336_));
 sg13g2_o21ai_1 _2230_ (.B1(_1336_),
    .Y(_1337_),
    .A1(_0928_),
    .A2(_1285_));
 sg13g2_o21ai_1 _2231_ (.B1(_1337_),
    .Y(_1338_),
    .A1(_1315_),
    .A2(_1294_));
 sg13g2_nand2_1 _2232_ (.Y(_1339_),
    .A(_1335_),
    .B(_1338_));
 sg13g2_o21ai_1 _2233_ (.B1(_1339_),
    .Y(_1340_),
    .A1(_1305_),
    .A2(_1313_));
 sg13g2_nand2_1 _2234_ (.Y(_1341_),
    .A(_1334_),
    .B(_1340_));
 sg13g2_xor2_1 _2235_ (.B(_1341_),
    .A(_1333_),
    .X(_1342_));
 sg13g2_nand2_1 _2236_ (.Y(_1343_),
    .A(\result[4] ),
    .B(net57));
 sg13g2_o21ai_1 _2237_ (.B1(_1343_),
    .Y(_1344_),
    .A1(net50),
    .A2(_1342_));
 sg13g2_nand2_1 _2238_ (.Y(_1345_),
    .A(net44),
    .B(_1344_));
 sg13g2_buf_1 _2239_ (.A(_0583_),
    .X(_1346_));
 sg13g2_a21oi_1 _2240_ (.A1(_1323_),
    .A2(_1345_),
    .Y(_0021_),
    .B1(net79));
 sg13g2_nor3_1 _2241_ (.A(_1305_),
    .B(_1313_),
    .C(_1332_),
    .Y(_1347_));
 sg13g2_o21ai_1 _2242_ (.B1(_1332_),
    .Y(_1348_),
    .A1(_1305_),
    .A2(_1313_));
 sg13g2_o21ai_1 _2243_ (.B1(_1348_),
    .Y(_1349_),
    .A1(\ad.a[12] ),
    .A2(_1347_));
 sg13g2_nor2b_1 _2244_ (.A(_1314_),
    .B_N(_1333_),
    .Y(_1350_));
 sg13g2_o21ai_1 _2245_ (.B1(_1297_),
    .Y(_1351_),
    .A1(_1315_),
    .A2(_1296_));
 sg13g2_nand2_1 _2246_ (.Y(_1352_),
    .A(_1350_),
    .B(_1351_));
 sg13g2_and2_1 _2247_ (.A(_1349_),
    .B(_1352_),
    .X(_1353_));
 sg13g2_o21ai_1 _2248_ (.B1(net65),
    .Y(_1354_),
    .A1(_1252_),
    .A2(_1255_));
 sg13g2_buf_1 _2249_ (.A(_0603_),
    .X(_1355_));
 sg13g2_nor2_1 _2250_ (.A(_1240_),
    .B(_1247_),
    .Y(_1356_));
 sg13g2_nor3_1 _2251_ (.A(net70),
    .B(net64),
    .C(_1356_),
    .Y(_1357_));
 sg13g2_o21ai_1 _2252_ (.B1(net64),
    .Y(_1358_),
    .A1(_1240_),
    .A2(_1247_));
 sg13g2_nand2_1 _2253_ (.Y(_1359_),
    .A(net71),
    .B(_1253_));
 sg13g2_a21oi_1 _2254_ (.A1(_1358_),
    .A2(_1359_),
    .Y(_1360_),
    .B1(net75));
 sg13g2_o21ai_1 _2255_ (.B1(net74),
    .Y(_1361_),
    .A1(_1357_),
    .A2(_1360_));
 sg13g2_nand2_1 _2256_ (.Y(_1362_),
    .A(_1354_),
    .B(_1361_));
 sg13g2_xor2_1 _2257_ (.B(_1362_),
    .A(\ad.a[13] ),
    .X(_1363_));
 sg13g2_xnor2_1 _2258_ (.Y(_1364_),
    .A(_1353_),
    .B(_1363_));
 sg13g2_nand2_1 _2259_ (.Y(_1365_),
    .A(net60),
    .B(_1364_));
 sg13g2_nand2_1 _2260_ (.Y(_1366_),
    .A(\result[5] ),
    .B(net52));
 sg13g2_a21oi_1 _2261_ (.A1(_1365_),
    .A2(_1366_),
    .Y(_1367_),
    .B1(net43));
 sg13g2_a21oi_1 _2262_ (.A1(\result[13] ),
    .A2(net40),
    .Y(_1368_),
    .B1(_1367_));
 sg13g2_nor2_1 _2263_ (.A(net76),
    .B(_1368_),
    .Y(_0022_));
 sg13g2_nand2_1 _2264_ (.Y(_0085_),
    .A(\result[14] ),
    .B(net41));
 sg13g2_xnor2_1 _2265_ (.Y(_0086_),
    .A(net37),
    .B(_0945_));
 sg13g2_xnor2_1 _2266_ (.Y(_0087_),
    .A(_0949_),
    .B(_0086_));
 sg13g2_nor2_1 _2267_ (.A(_0931_),
    .B(_0087_),
    .Y(_0088_));
 sg13g2_a21oi_1 _2268_ (.A1(_0931_),
    .A2(net36),
    .Y(_0089_),
    .B1(_0088_));
 sg13g2_nand2_1 _2269_ (.Y(_0090_),
    .A(net63),
    .B(_1106_));
 sg13g2_o21ai_1 _2270_ (.B1(_0090_),
    .Y(_0091_),
    .A1(_0588_),
    .A2(_0089_));
 sg13g2_a22oi_1 _2271_ (.Y(_0092_),
    .B1(_0091_),
    .B2(net74),
    .A2(_0952_),
    .A1(net65));
 sg13g2_o21ai_1 _2272_ (.B1(_0937_),
    .Y(_0093_),
    .A1(_1277_),
    .A2(_1281_));
 sg13g2_a21oi_1 _2273_ (.A1(\ad.a[8] ),
    .A2(_0093_),
    .Y(_0094_),
    .B1(_1283_));
 sg13g2_nand3b_1 _2274_ (.B(_1335_),
    .C(_1350_),
    .Y(_0095_),
    .A_N(_0929_));
 sg13g2_inv_1 _2275_ (.Y(_0096_),
    .A(_1287_));
 sg13g2_o21ai_1 _2276_ (.B1(\ad.a[10] ),
    .Y(_0097_),
    .A1(_1287_),
    .A2(_1295_));
 sg13g2_o21ai_1 _2277_ (.B1(_0097_),
    .Y(_0098_),
    .A1(_0096_),
    .A2(_1294_));
 sg13g2_nand2_1 _2278_ (.Y(_0099_),
    .A(_1350_),
    .B(_0098_));
 sg13g2_o21ai_1 _2279_ (.B1(_0099_),
    .Y(_0100_),
    .A1(_0094_),
    .A2(_0095_));
 sg13g2_nand2b_1 _2280_ (.Y(_0101_),
    .B(_1349_),
    .A_N(_0100_));
 sg13g2_a21oi_1 _2281_ (.A1(\ad.a[13] ),
    .A2(_1362_),
    .Y(_0102_),
    .B1(_0101_));
 sg13g2_or2_1 _2282_ (.X(_0103_),
    .B(_1362_),
    .A(\ad.a[13] ));
 sg13g2_nand2b_1 _2283_ (.Y(_0104_),
    .B(_0103_),
    .A_N(_0102_));
 sg13g2_xor2_1 _2284_ (.B(_0104_),
    .A(_0092_),
    .X(_0105_));
 sg13g2_xnor2_1 _2285_ (.Y(_0106_),
    .A(\ad.a[14] ),
    .B(_0105_));
 sg13g2_nand2_1 _2286_ (.Y(_0107_),
    .A(\result[6] ),
    .B(net57));
 sg13g2_o21ai_1 _2287_ (.B1(_0107_),
    .Y(_0108_),
    .A1(net50),
    .A2(_0106_));
 sg13g2_nand2_1 _2288_ (.Y(_0109_),
    .A(_0847_),
    .B(_0108_));
 sg13g2_a21oi_1 _2289_ (.A1(_0085_),
    .A2(_0109_),
    .Y(_0023_),
    .B1(net79));
 sg13g2_nand2_1 _2290_ (.Y(_0110_),
    .A(\result[15] ),
    .B(net41));
 sg13g2_buf_1 _2291_ (.A(\ad.a[15] ),
    .X(_0111_));
 sg13g2_buf_1 _2292_ (.A(net64),
    .X(_0112_));
 sg13g2_xnor2_1 _2293_ (.Y(_0113_),
    .A(_0689_),
    .B(_1118_));
 sg13g2_nor2_1 _2294_ (.A(net59),
    .B(_0113_),
    .Y(_0114_));
 sg13g2_nor2_1 _2295_ (.A(net71),
    .B(_0113_),
    .Y(_0115_));
 sg13g2_or2_1 _2296_ (.X(_0116_),
    .B(_0115_),
    .A(_1125_));
 sg13g2_a22oi_1 _2297_ (.Y(_0117_),
    .B1(_0116_),
    .B2(net65),
    .A2(_0114_),
    .A1(net62));
 sg13g2_buf_1 _2298_ (.A(_0117_),
    .X(_0118_));
 sg13g2_nand2b_1 _2299_ (.Y(_0119_),
    .B(_0092_),
    .A_N(\ad.a[14] ));
 sg13g2_and2_1 _2300_ (.A(_0103_),
    .B(_0119_),
    .X(_0120_));
 sg13g2_nand2b_1 _2301_ (.Y(_0121_),
    .B(\ad.a[14] ),
    .A_N(_0092_));
 sg13g2_a21oi_1 _2302_ (.A1(_1354_),
    .A2(_1361_),
    .Y(_0122_),
    .B1(_1349_));
 sg13g2_nand3_1 _2303_ (.B(_1354_),
    .C(_1361_),
    .A(_1349_),
    .Y(_0123_));
 sg13g2_o21ai_1 _2304_ (.B1(_0123_),
    .Y(_0124_),
    .A1(\ad.a[13] ),
    .A2(_0122_));
 sg13g2_inv_1 _2305_ (.Y(_0125_),
    .A(_0119_));
 sg13g2_a21oi_1 _2306_ (.A1(_0121_),
    .A2(_0124_),
    .Y(_0126_),
    .B1(_0125_));
 sg13g2_a21oi_2 _2307_ (.B1(_0126_),
    .Y(_0127_),
    .A2(_0120_),
    .A1(_0100_));
 sg13g2_xnor2_1 _2308_ (.Y(_0128_),
    .A(_0118_),
    .B(_0127_));
 sg13g2_xor2_1 _2309_ (.B(_0128_),
    .A(_0111_),
    .X(_0129_));
 sg13g2_nand2_1 _2310_ (.Y(_0130_),
    .A(\result[7] ),
    .B(net57));
 sg13g2_o21ai_1 _2311_ (.B1(_0130_),
    .Y(_0131_),
    .A1(net50),
    .A2(_0129_));
 sg13g2_nand2_1 _2312_ (.Y(_0132_),
    .A(_0847_),
    .B(_0131_));
 sg13g2_a21oi_1 _2313_ (.A1(_0110_),
    .A2(_0132_),
    .Y(_0024_),
    .B1(net79));
 sg13g2_buf_1 _2314_ (.A(net57),
    .X(_0133_));
 sg13g2_and2_1 _2315_ (.A(net84),
    .B(_0605_),
    .X(_0134_));
 sg13g2_a21oi_1 _2316_ (.A1(net82),
    .A2(_0933_),
    .Y(_0135_),
    .B1(_0134_));
 sg13g2_a21oi_1 _2317_ (.A1(net72),
    .A2(_0830_),
    .Y(_0136_),
    .B1(_0606_));
 sg13g2_nor2_1 _2318_ (.A(net75),
    .B(_0136_),
    .Y(_0137_));
 sg13g2_a21oi_1 _2319_ (.A1(net75),
    .A2(_0135_),
    .Y(_0138_),
    .B1(_0137_));
 sg13g2_xnor2_1 _2320_ (.Y(_0139_),
    .A(_0005_),
    .B(_0138_));
 sg13g2_and2_1 _2321_ (.A(_0100_),
    .B(_0120_),
    .X(_0140_));
 sg13g2_nand2b_1 _2322_ (.Y(_0141_),
    .B(_0118_),
    .A_N(_0126_));
 sg13g2_o21ai_1 _2323_ (.B1(_0111_),
    .Y(_0142_),
    .A1(_0140_),
    .A2(_0141_));
 sg13g2_or2_1 _2324_ (.X(_0143_),
    .B(_0127_),
    .A(_0118_));
 sg13g2_and2_1 _2325_ (.A(_0142_),
    .B(_0143_),
    .X(_0144_));
 sg13g2_xnor2_1 _2326_ (.Y(_0145_),
    .A(_0139_),
    .B(_0144_));
 sg13g2_nor2_2 _2327_ (.A(net53),
    .B(_1272_),
    .Y(_0146_));
 sg13g2_buf_1 _2328_ (.A(_0146_),
    .X(_0147_));
 sg13g2_a22oi_1 _2329_ (.Y(_0148_),
    .B1(net39),
    .B2(\result[8] ),
    .A2(_0600_),
    .A1(net53));
 sg13g2_o21ai_1 _2330_ (.B1(_0148_),
    .Y(_0149_),
    .A1(net48),
    .A2(_0145_));
 sg13g2_and2_1 _2331_ (.A(_0571_),
    .B(_0149_),
    .X(_0025_));
 sg13g2_nor2_1 _2332_ (.A(_0919_),
    .B(_0920_),
    .Y(_0150_));
 sg13g2_o21ai_1 _2333_ (.B1(_1164_),
    .Y(_0151_),
    .A1(_0609_),
    .A2(_0150_));
 sg13g2_nor2_1 _2334_ (.A(net84),
    .B(_0924_),
    .Y(_0152_));
 sg13g2_a221oi_1 _2335_ (.B2(_0926_),
    .C1(net70),
    .B1(_0152_),
    .A1(net84),
    .Y(_0153_),
    .A2(_1163_));
 sg13g2_a21oi_1 _2336_ (.A1(net70),
    .A2(_0151_),
    .Y(_0154_),
    .B1(_0153_));
 sg13g2_xnor2_1 _2337_ (.Y(_0155_),
    .A(_0006_),
    .B(_0154_));
 sg13g2_inv_1 _2338_ (.Y(_0156_),
    .A(_0155_));
 sg13g2_nor2b_1 _2339_ (.A(_0138_),
    .B_N(\ad.a[16] ),
    .Y(_0157_));
 sg13g2_a21oi_1 _2340_ (.A1(_0142_),
    .A2(_0143_),
    .Y(_0158_),
    .B1(_0139_));
 sg13g2_nor2_1 _2341_ (.A(_0157_),
    .B(_0158_),
    .Y(_0159_));
 sg13g2_xnor2_1 _2342_ (.Y(_0160_),
    .A(_0156_),
    .B(_0159_));
 sg13g2_buf_1 _2343_ (.A(net60),
    .X(_0161_));
 sg13g2_buf_1 _2344_ (.A(_0845_),
    .X(_0162_));
 sg13g2_nor2_1 _2345_ (.A(net47),
    .B(_0853_),
    .Y(_0163_));
 sg13g2_a221oi_1 _2346_ (.B2(net56),
    .C1(_0163_),
    .B1(_0160_),
    .A1(\result[9] ),
    .Y(_0164_),
    .A2(net39));
 sg13g2_nor2_1 _2347_ (.A(net76),
    .B(_0164_),
    .Y(_0026_));
 sg13g2_buf_1 _2348_ (.A(net53),
    .X(_0165_));
 sg13g2_buf_1 _2349_ (.A(_0146_),
    .X(_0166_));
 sg13g2_a22oi_1 _2350_ (.Y(_0167_),
    .B1(net38),
    .B2(\result[10] ),
    .A2(_1144_),
    .A1(net42));
 sg13g2_buf_1 _2351_ (.A(net82),
    .X(_0168_));
 sg13g2_and2_1 _2352_ (.A(net74),
    .B(_1145_),
    .X(_0169_));
 sg13g2_a21oi_1 _2353_ (.A1(net69),
    .A2(_1291_),
    .Y(_0170_),
    .B1(_0169_));
 sg13g2_a21oi_1 _2354_ (.A1(net72),
    .A2(_1202_),
    .Y(_0171_),
    .B1(_1146_));
 sg13g2_nor2_1 _2355_ (.A(net75),
    .B(_0171_),
    .Y(_0172_));
 sg13g2_a21oi_2 _2356_ (.B1(_0172_),
    .Y(_0173_),
    .A2(_0170_),
    .A1(net68));
 sg13g2_or2_1 _2357_ (.X(_0174_),
    .B(_0155_),
    .A(_0139_));
 sg13g2_buf_1 _2358_ (.A(_0174_),
    .X(_0175_));
 sg13g2_nor2b_1 _2359_ (.A(_0154_),
    .B_N(\ad.a[17] ),
    .Y(_0176_));
 sg13g2_a21oi_1 _2360_ (.A1(_0156_),
    .A2(_0157_),
    .Y(_0177_),
    .B1(_0176_));
 sg13g2_o21ai_1 _2361_ (.B1(_0177_),
    .Y(_0178_),
    .A1(_0144_),
    .A2(_0175_));
 sg13g2_xor2_1 _2362_ (.B(_0178_),
    .A(_0173_),
    .X(_0179_));
 sg13g2_xnor2_1 _2363_ (.Y(_0180_),
    .A(\ad.a[18] ),
    .B(_0179_));
 sg13g2_nand2_1 _2364_ (.Y(_0181_),
    .A(net56),
    .B(_0180_));
 sg13g2_a21oi_1 _2365_ (.A1(_0167_),
    .A2(_0181_),
    .Y(_0027_),
    .B1(net79));
 sg13g2_inv_1 _2366_ (.Y(_0182_),
    .A(\ad.a[19] ));
 sg13g2_nand2_1 _2367_ (.Y(_0183_),
    .A(net59),
    .B(net7));
 sg13g2_nand2_1 _2368_ (.Y(_0184_),
    .A(net74),
    .B(_0183_));
 sg13g2_o21ai_1 _2369_ (.B1(_0184_),
    .Y(_0185_),
    .A1(net74),
    .A2(_1310_));
 sg13g2_nor3_1 _2370_ (.A(net69),
    .B(net59),
    .C(_1308_),
    .Y(_0186_));
 sg13g2_nor2_1 _2371_ (.A(net74),
    .B(_0183_),
    .Y(_0187_));
 sg13g2_o21ai_1 _2372_ (.B1(net70),
    .Y(_0188_),
    .A1(_0186_),
    .A2(_0187_));
 sg13g2_o21ai_1 _2373_ (.B1(_0188_),
    .Y(_0189_),
    .A1(net70),
    .A2(_0185_));
 sg13g2_nor2b_1 _2374_ (.A(_0176_),
    .B_N(_0173_),
    .Y(_0190_));
 sg13g2_o21ai_1 _2375_ (.B1(_0156_),
    .Y(_0191_),
    .A1(_0157_),
    .A2(_0158_));
 sg13g2_inv_1 _2376_ (.Y(_0192_),
    .A(\ad.a[18] ));
 sg13g2_a21oi_1 _2377_ (.A1(_0190_),
    .A2(_0191_),
    .Y(_0193_),
    .B1(_0192_));
 sg13g2_nor2b_1 _2378_ (.A(_0118_),
    .B_N(_0111_),
    .Y(_0194_));
 sg13g2_nand2b_1 _2379_ (.Y(_0195_),
    .B(_0194_),
    .A_N(_0175_));
 sg13g2_a21oi_1 _2380_ (.A1(_0177_),
    .A2(_0195_),
    .Y(_0196_),
    .B1(_0173_));
 sg13g2_nor2b_1 _2381_ (.A(_0111_),
    .B_N(_0118_),
    .Y(_0197_));
 sg13g2_nor4_1 _2382_ (.A(_0127_),
    .B(_0173_),
    .C(_0175_),
    .D(_0197_),
    .Y(_0198_));
 sg13g2_or2_1 _2383_ (.X(_0199_),
    .B(_0198_),
    .A(_0196_));
 sg13g2_nor3_1 _2384_ (.A(_0189_),
    .B(_0193_),
    .C(_0199_),
    .Y(_0200_));
 sg13g2_o21ai_1 _2385_ (.B1(_0189_),
    .Y(_0201_),
    .A1(_0193_),
    .A2(_0199_));
 sg13g2_nor2b_1 _2386_ (.A(_0200_),
    .B_N(_0201_),
    .Y(_0202_));
 sg13g2_xnor2_1 _2387_ (.Y(_0203_),
    .A(_0182_),
    .B(_0202_));
 sg13g2_nand2_1 _2388_ (.Y(_0204_),
    .A(net56),
    .B(_0203_));
 sg13g2_a22oi_1 _2389_ (.Y(_0205_),
    .B1(net38),
    .B2(\result[11] ),
    .A2(_1183_),
    .A1(net43));
 sg13g2_a21oi_1 _2390_ (.A1(_0204_),
    .A2(_0205_),
    .Y(_0028_),
    .B1(net79));
 sg13g2_nand2_1 _2391_ (.Y(_0206_),
    .A(_1172_),
    .B(_1166_));
 sg13g2_xnor2_1 _2392_ (.Y(_0207_),
    .A(_1153_),
    .B(_1162_));
 sg13g2_xnor2_1 _2393_ (.Y(_0208_),
    .A(_0206_),
    .B(_0207_));
 sg13g2_a22oi_1 _2394_ (.Y(_0209_),
    .B1(_0840_),
    .B2(_0208_),
    .A2(net46),
    .A1(\result[1] ));
 sg13g2_nor2_1 _2395_ (.A(net76),
    .B(_0209_),
    .Y(_0029_));
 sg13g2_a22oi_1 _2396_ (.Y(_0210_),
    .B1(net38),
    .B2(\result[12] ),
    .A2(_1208_),
    .A1(net42));
 sg13g2_xnor2_1 _2397_ (.Y(_0211_),
    .A(_0192_),
    .B(_0173_));
 sg13g2_nor4_1 _2398_ (.A(_0127_),
    .B(_0175_),
    .C(_0197_),
    .D(_0211_),
    .Y(_0212_));
 sg13g2_inv_1 _2399_ (.Y(_0213_),
    .A(_0139_));
 sg13g2_a21oi_1 _2400_ (.A1(_0213_),
    .A2(_0194_),
    .Y(_0214_),
    .B1(_0157_));
 sg13g2_o21ai_1 _2401_ (.B1(_0190_),
    .Y(_0215_),
    .A1(_0155_),
    .A2(_0214_));
 sg13g2_a21o_1 _2402_ (.A2(_0215_),
    .A1(\ad.a[18] ),
    .B1(_0196_),
    .X(_0216_));
 sg13g2_o21ai_1 _2403_ (.B1(_0189_),
    .Y(_0217_),
    .A1(_0212_),
    .A2(_0216_));
 sg13g2_nor3_1 _2404_ (.A(_0189_),
    .B(_0212_),
    .C(_0216_),
    .Y(_0218_));
 sg13g2_a21oi_1 _2405_ (.A1(_0182_),
    .A2(_0217_),
    .Y(_0219_),
    .B1(_0218_));
 sg13g2_nand2_1 _2406_ (.Y(_0220_),
    .A(_0112_),
    .B(net8));
 sg13g2_nor2_1 _2407_ (.A(net67),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_a21oi_1 _2408_ (.A1(net67),
    .A2(_1325_),
    .Y(_0222_),
    .B1(_0221_));
 sg13g2_nor2_1 _2409_ (.A(net69),
    .B(net71),
    .Y(_0223_));
 sg13g2_a221oi_1 _2410_ (.B2(net69),
    .C1(net70),
    .B1(_1328_),
    .A1(net8),
    .Y(_0224_),
    .A2(_0223_));
 sg13g2_a21oi_2 _2411_ (.B1(_0224_),
    .Y(_0225_),
    .A2(_0222_),
    .A1(net70));
 sg13g2_xnor2_1 _2412_ (.Y(_0226_),
    .A(\ad.a[20] ),
    .B(_0225_));
 sg13g2_xnor2_1 _2413_ (.Y(_0227_),
    .A(_0219_),
    .B(_0226_));
 sg13g2_nand2_1 _2414_ (.Y(_0228_),
    .A(net56),
    .B(_0227_));
 sg13g2_a21oi_1 _2415_ (.A1(_0210_),
    .A2(_0228_),
    .Y(_0030_),
    .B1(_1346_));
 sg13g2_a22oi_1 _2416_ (.Y(_0229_),
    .B1(net38),
    .B2(\result[13] ),
    .A2(_1253_),
    .A1(net42));
 sg13g2_buf_2 _2417_ (.A(\ad.a[21] ),
    .X(_0230_));
 sg13g2_nor3_1 _2418_ (.A(net69),
    .B(net59),
    .C(_1356_),
    .Y(_0231_));
 sg13g2_nor2_1 _2419_ (.A(_1258_),
    .B(_0231_),
    .Y(_0232_));
 sg13g2_nand2_1 _2420_ (.Y(_0233_),
    .A(net67),
    .B(_1257_));
 sg13g2_nand3_1 _2421_ (.B(_1358_),
    .C(_1359_),
    .A(net69),
    .Y(_0234_));
 sg13g2_nand3_1 _2422_ (.B(_0233_),
    .C(_0234_),
    .A(net68),
    .Y(_0235_));
 sg13g2_o21ai_1 _2423_ (.B1(_0235_),
    .Y(_0236_),
    .A1(net68),
    .A2(_0232_));
 sg13g2_inv_1 _2424_ (.Y(_0237_),
    .A(_0236_));
 sg13g2_and2_1 _2425_ (.A(\ad.a[20] ),
    .B(_0225_),
    .X(_0238_));
 sg13g2_a21oi_1 _2426_ (.A1(_0182_),
    .A2(_0201_),
    .Y(_0239_),
    .B1(_0200_));
 sg13g2_or2_1 _2427_ (.X(_0240_),
    .B(_0225_),
    .A(\ad.a[20] ));
 sg13g2_o21ai_1 _2428_ (.B1(_0240_),
    .Y(_0241_),
    .A1(_0238_),
    .A2(_0239_));
 sg13g2_xnor2_1 _2429_ (.Y(_0242_),
    .A(_0237_),
    .B(_0241_));
 sg13g2_xnor2_1 _2430_ (.Y(_0243_),
    .A(_0230_),
    .B(_0242_));
 sg13g2_nand2_1 _2431_ (.Y(_0244_),
    .A(net56),
    .B(_0243_));
 sg13g2_a21oi_1 _2432_ (.A1(_0229_),
    .A2(_0244_),
    .Y(_0031_),
    .B1(net79));
 sg13g2_a21o_1 _2433_ (.A2(_0225_),
    .A1(_0219_),
    .B1(\ad.a[20] ),
    .X(_0245_));
 sg13g2_or2_1 _2434_ (.X(_0246_),
    .B(_0225_),
    .A(_0219_));
 sg13g2_a22oi_1 _2435_ (.Y(_0247_),
    .B1(_0245_),
    .B2(_0246_),
    .A2(_0236_),
    .A1(_0230_));
 sg13g2_nor2_1 _2436_ (.A(_0230_),
    .B(_0236_),
    .Y(_0248_));
 sg13g2_or2_1 _2437_ (.X(_0249_),
    .B(_0248_),
    .A(_0247_));
 sg13g2_buf_1 _2438_ (.A(_0249_),
    .X(_0250_));
 sg13g2_buf_2 _2439_ (.A(\ad.a[22] ),
    .X(_0251_));
 sg13g2_and2_1 _2440_ (.A(_0592_),
    .B(_0953_),
    .X(_0252_));
 sg13g2_a21oi_1 _2441_ (.A1(net69),
    .A2(_0089_),
    .Y(_0253_),
    .B1(_0252_));
 sg13g2_a21oi_1 _2442_ (.A1(_0958_),
    .A2(net36),
    .Y(_0254_),
    .B1(_0954_));
 sg13g2_nor2_1 _2443_ (.A(net68),
    .B(_0254_),
    .Y(_0255_));
 sg13g2_a21oi_2 _2444_ (.B1(_0255_),
    .Y(_0256_),
    .A2(_0253_),
    .A1(_0589_));
 sg13g2_xnor2_1 _2445_ (.Y(_0257_),
    .A(_0251_),
    .B(_0256_));
 sg13g2_xnor2_1 _2446_ (.Y(_0258_),
    .A(_0250_),
    .B(_0257_));
 sg13g2_buf_1 _2447_ (.A(net60),
    .X(_0259_));
 sg13g2_nor2_1 _2448_ (.A(net47),
    .B(_0087_),
    .Y(_0260_));
 sg13g2_a221oi_1 _2449_ (.B2(net55),
    .C1(_0260_),
    .B1(_0258_),
    .A1(\result[14] ),
    .Y(_0261_),
    .A2(net39));
 sg13g2_nor2_1 _2450_ (.A(_0585_),
    .B(_0261_),
    .Y(_0032_));
 sg13g2_nor3_1 _2451_ (.A(net67),
    .B(net59),
    .C(_0113_),
    .Y(_0262_));
 sg13g2_a21oi_1 _2452_ (.A1(net67),
    .A2(_1124_),
    .Y(_0263_),
    .B1(_0262_));
 sg13g2_nand2_1 _2453_ (.Y(_0264_),
    .A(_0594_),
    .B(_1124_));
 sg13g2_o21ai_1 _2454_ (.B1(_0264_),
    .Y(_0265_),
    .A1(net70),
    .A2(_0263_));
 sg13g2_xor2_1 _2455_ (.B(_0265_),
    .A(_0007_),
    .X(_0266_));
 sg13g2_inv_1 _2456_ (.Y(_0267_),
    .A(_0266_));
 sg13g2_inv_1 _2457_ (.Y(_0268_),
    .A(_0230_));
 sg13g2_inv_1 _2458_ (.Y(_0269_),
    .A(_0251_));
 sg13g2_a221oi_1 _2459_ (.B2(_0269_),
    .C1(_0241_),
    .B1(_0256_),
    .A1(_0268_),
    .Y(_0270_),
    .A2(_0237_));
 sg13g2_nand2b_1 _2460_ (.Y(_0271_),
    .B(_0251_),
    .A_N(_0256_));
 sg13g2_nand3b_1 _2461_ (.B(_0230_),
    .C(_0236_),
    .Y(_0272_),
    .A_N(_0256_));
 sg13g2_nand3_1 _2462_ (.B(_0251_),
    .C(_0236_),
    .A(_0230_),
    .Y(_0273_));
 sg13g2_nand3_1 _2463_ (.B(_0272_),
    .C(_0273_),
    .A(_0271_),
    .Y(_0274_));
 sg13g2_nor2_1 _2464_ (.A(_0270_),
    .B(_0274_),
    .Y(_0275_));
 sg13g2_xnor2_1 _2465_ (.Y(_0276_),
    .A(_0267_),
    .B(_0275_));
 sg13g2_nor2_1 _2466_ (.A(net47),
    .B(_0113_),
    .Y(_0277_));
 sg13g2_a221oi_1 _2467_ (.B2(net55),
    .C1(_0277_),
    .B1(_0276_),
    .A1(\result[15] ),
    .Y(_0278_),
    .A2(net39));
 sg13g2_nor2_1 _2468_ (.A(_0585_),
    .B(_0278_),
    .Y(_0033_));
 sg13g2_mux2_1 _2469_ (.A0(net4),
    .A1(_0830_),
    .S(_0168_),
    .X(_0279_));
 sg13g2_nor2_1 _2470_ (.A(net66),
    .B(_0605_),
    .Y(_0280_));
 sg13g2_a21oi_1 _2471_ (.A1(net63),
    .A2(_0279_),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_xnor2_1 _2472_ (.Y(_0282_),
    .A(_0008_),
    .B(_0281_));
 sg13g2_inv_1 _2473_ (.Y(_0283_),
    .A(_0282_));
 sg13g2_nand2_1 _2474_ (.Y(_0284_),
    .A(_0257_),
    .B(_0267_));
 sg13g2_nand2_1 _2475_ (.Y(_0285_),
    .A(\ad.a[23] ),
    .B(_0265_));
 sg13g2_o21ai_1 _2476_ (.B1(_0285_),
    .Y(_0286_),
    .A1(_0271_),
    .A2(_0266_));
 sg13g2_inv_1 _2477_ (.Y(_0287_),
    .A(_0286_));
 sg13g2_o21ai_1 _2478_ (.B1(_0287_),
    .Y(_0288_),
    .A1(_0250_),
    .A2(_0284_));
 sg13g2_xnor2_1 _2479_ (.Y(_0289_),
    .A(_0283_),
    .B(_0288_));
 sg13g2_a22oi_1 _2480_ (.Y(_0290_),
    .B1(_0147_),
    .B2(\result[16] ),
    .A2(_0830_),
    .A1(net53));
 sg13g2_o21ai_1 _2481_ (.B1(_0290_),
    .Y(_0291_),
    .A1(_0133_),
    .A2(_0289_));
 sg13g2_and2_1 _2482_ (.A(net96),
    .B(_0291_),
    .X(_0034_));
 sg13g2_nand2_1 _2483_ (.Y(_0292_),
    .A(_0593_),
    .B(net5));
 sg13g2_o21ai_1 _2484_ (.B1(_0292_),
    .Y(_0293_),
    .A1(net67),
    .A2(_0150_));
 sg13g2_nand2_1 _2485_ (.Y(_0294_),
    .A(net63),
    .B(_0293_));
 sg13g2_o21ai_1 _2486_ (.B1(_0294_),
    .Y(_0295_),
    .A1(net66),
    .A2(_1163_));
 sg13g2_xor2_1 _2487_ (.B(_0295_),
    .A(_0009_),
    .X(_0296_));
 sg13g2_nor2b_1 _2488_ (.A(_0281_),
    .B_N(\ad.a[24] ),
    .Y(_0297_));
 sg13g2_o21ai_1 _2489_ (.B1(_0267_),
    .Y(_0298_),
    .A1(_0270_),
    .A2(_0274_));
 sg13g2_a21oi_1 _2490_ (.A1(_0285_),
    .A2(_0298_),
    .Y(_0299_),
    .B1(_0282_));
 sg13g2_nor2_1 _2491_ (.A(_0297_),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_xnor2_1 _2492_ (.Y(_0301_),
    .A(_0296_),
    .B(_0300_));
 sg13g2_nor2_1 _2493_ (.A(_0846_),
    .B(_0150_),
    .Y(_0302_));
 sg13g2_a21oi_1 _2494_ (.A1(\result[17] ),
    .A2(_0146_),
    .Y(_0303_),
    .B1(_0302_));
 sg13g2_o21ai_1 _2495_ (.B1(_0303_),
    .Y(_0304_),
    .A1(net50),
    .A2(_0301_));
 sg13g2_and2_1 _2496_ (.A(net96),
    .B(_0304_),
    .X(_0035_));
 sg13g2_a21oi_1 _2497_ (.A1(_0283_),
    .A2(_0286_),
    .Y(_0305_),
    .B1(_0297_));
 sg13g2_nand2_1 _2498_ (.Y(_0306_),
    .A(\ad.a[25] ),
    .B(_0295_));
 sg13g2_o21ai_1 _2499_ (.B1(_0306_),
    .Y(_0307_),
    .A1(_0296_),
    .A2(_0305_));
 sg13g2_or2_1 _2500_ (.X(_0308_),
    .B(_0296_),
    .A(_0282_));
 sg13g2_nor4_1 _2501_ (.A(_0247_),
    .B(_0248_),
    .C(_0284_),
    .D(_0308_),
    .Y(_0309_));
 sg13g2_nor2_1 _2502_ (.A(_0307_),
    .B(_0309_),
    .Y(_0310_));
 sg13g2_buf_1 _2503_ (.A(_0593_),
    .X(_0311_));
 sg13g2_xnor2_1 _2504_ (.Y(_0312_),
    .A(_1132_),
    .B(_1212_));
 sg13g2_nand2_1 _2505_ (.Y(_0313_),
    .A(net67),
    .B(net6));
 sg13g2_o21ai_1 _2506_ (.B1(_0313_),
    .Y(_0314_),
    .A1(net58),
    .A2(_0312_));
 sg13g2_nor2_1 _2507_ (.A(net66),
    .B(_1145_),
    .Y(_0315_));
 sg13g2_a21oi_1 _2508_ (.A1(net63),
    .A2(_0314_),
    .Y(_0316_),
    .B1(_0315_));
 sg13g2_xnor2_1 _2509_ (.Y(_0317_),
    .A(_0000_),
    .B(_0316_));
 sg13g2_xnor2_1 _2510_ (.Y(_0318_),
    .A(_0310_),
    .B(_0317_));
 sg13g2_a22oi_1 _2511_ (.Y(_0319_),
    .B1(net39),
    .B2(\result[18] ),
    .A2(_1202_),
    .A1(_0596_));
 sg13g2_o21ai_1 _2512_ (.B1(_0319_),
    .Y(_0320_),
    .A1(net50),
    .A2(_0318_));
 sg13g2_and2_1 _2513_ (.A(net96),
    .B(_0320_),
    .X(_0036_));
 sg13g2_inv_1 _2514_ (.Y(_0321_),
    .A(_1308_));
 sg13g2_a22oi_1 _2515_ (.Y(_0322_),
    .B1(net38),
    .B2(\result[19] ),
    .A2(_0321_),
    .A1(_0165_));
 sg13g2_a21oi_1 _2516_ (.A1(_0285_),
    .A2(_0298_),
    .Y(_0323_),
    .B1(_0308_));
 sg13g2_nand2b_1 _2517_ (.Y(_0324_),
    .B(_0297_),
    .A_N(_0009_));
 sg13g2_and2_1 _2518_ (.A(_0009_),
    .B(_0297_),
    .X(_0325_));
 sg13g2_o21ai_1 _2519_ (.B1(_0295_),
    .Y(_0326_),
    .A1(\ad.a[25] ),
    .A2(_0325_));
 sg13g2_o21ai_1 _2520_ (.B1(_0326_),
    .Y(_0327_),
    .A1(_0295_),
    .A2(_0324_));
 sg13g2_inv_1 _2521_ (.Y(_0328_),
    .A(_0317_));
 sg13g2_o21ai_1 _2522_ (.B1(_0328_),
    .Y(_0329_),
    .A1(_0323_),
    .A2(_0327_));
 sg13g2_inv_1 _2523_ (.Y(_0330_),
    .A(_0316_));
 sg13g2_nand2_1 _2524_ (.Y(_0331_),
    .A(\ad.a[26] ),
    .B(_0330_));
 sg13g2_nand2_1 _2525_ (.Y(_0332_),
    .A(_0329_),
    .B(_0331_));
 sg13g2_nand2_1 _2526_ (.Y(_0333_),
    .A(net58),
    .B(net7));
 sg13g2_o21ai_1 _2527_ (.B1(_0333_),
    .Y(_0334_),
    .A1(net58),
    .A2(_1308_));
 sg13g2_nand2_1 _2528_ (.Y(_0335_),
    .A(net63),
    .B(_0334_));
 sg13g2_o21ai_1 _2529_ (.B1(_0335_),
    .Y(_0336_),
    .A1(net66),
    .A2(_0183_));
 sg13g2_xnor2_1 _2530_ (.Y(_0337_),
    .A(_0001_),
    .B(_0336_));
 sg13g2_inv_1 _2531_ (.Y(_0338_),
    .A(_0337_));
 sg13g2_xnor2_1 _2532_ (.Y(_0339_),
    .A(_0332_),
    .B(_0338_));
 sg13g2_nand2_1 _2533_ (.Y(_0340_),
    .A(net56),
    .B(_0339_));
 sg13g2_a21oi_1 _2534_ (.A1(_0322_),
    .A2(_0340_),
    .Y(_0037_),
    .B1(net79));
 sg13g2_nand2_1 _2535_ (.Y(_0341_),
    .A(net58),
    .B(net8));
 sg13g2_nand2_1 _2536_ (.Y(_0342_),
    .A(net68),
    .B(_1326_));
 sg13g2_a21oi_1 _2537_ (.A1(_1229_),
    .A2(_0341_),
    .Y(_0343_),
    .B1(_0342_));
 sg13g2_or2_1 _2538_ (.X(_0344_),
    .B(_0220_),
    .A(_0834_));
 sg13g2_nand2b_1 _2539_ (.Y(_0345_),
    .B(_0344_),
    .A_N(_0343_));
 sg13g2_xor2_1 _2540_ (.B(_0345_),
    .A(_0002_),
    .X(_0346_));
 sg13g2_and2_1 _2541_ (.A(\ad.a[27] ),
    .B(_0336_),
    .X(_0347_));
 sg13g2_inv_1 _2542_ (.Y(_0348_),
    .A(_0347_));
 sg13g2_inv_1 _2543_ (.Y(_0349_),
    .A(\ad.a[26] ));
 sg13g2_o21ai_1 _2544_ (.B1(_0000_),
    .Y(_0350_),
    .A1(_0307_),
    .A2(_0309_));
 sg13g2_a21oi_1 _2545_ (.A1(_0349_),
    .A2(_0350_),
    .Y(_0351_),
    .B1(_0316_));
 sg13g2_nor3_1 _2546_ (.A(_0000_),
    .B(_0310_),
    .C(_0330_),
    .Y(_0352_));
 sg13g2_o21ai_1 _2547_ (.B1(_0337_),
    .Y(_0353_),
    .A1(_0351_),
    .A2(_0352_));
 sg13g2_nand2_1 _2548_ (.Y(_0354_),
    .A(_0348_),
    .B(_0353_));
 sg13g2_xor2_1 _2549_ (.B(_0354_),
    .A(_0346_),
    .X(_0355_));
 sg13g2_inv_1 _2550_ (.Y(_0356_),
    .A(_1324_));
 sg13g2_a22oi_1 _2551_ (.Y(_0357_),
    .B1(_0146_),
    .B2(\result[20] ),
    .A2(_0356_),
    .A1(_0596_));
 sg13g2_o21ai_1 _2552_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_0848_),
    .A2(_0355_));
 sg13g2_and2_1 _2553_ (.A(_0571_),
    .B(_0358_),
    .X(_0038_));
 sg13g2_inv_1 _2554_ (.Y(_0359_),
    .A(\ad.a[29] ));
 sg13g2_nand2_2 _2555_ (.Y(_0360_),
    .A(\ad.a[28] ),
    .B(_0345_));
 sg13g2_a21o_1 _2556_ (.A2(_0331_),
    .A1(_0329_),
    .B1(_0338_),
    .X(_0361_));
 sg13g2_a21o_1 _2557_ (.A2(_0361_),
    .A1(_0348_),
    .B1(_0346_),
    .X(_0362_));
 sg13g2_nand2_1 _2558_ (.Y(_0363_),
    .A(net58),
    .B(net9));
 sg13g2_o21ai_1 _2559_ (.B1(_0363_),
    .Y(_0364_),
    .A1(net58),
    .A2(_1356_));
 sg13g2_nand2_1 _2560_ (.Y(_0365_),
    .A(net63),
    .B(_0364_));
 sg13g2_o21ai_1 _2561_ (.B1(_0365_),
    .Y(_0366_),
    .A1(net66),
    .A2(_1257_));
 sg13g2_a21oi_1 _2562_ (.A1(_0360_),
    .A2(_0362_),
    .Y(_0367_),
    .B1(_0366_));
 sg13g2_and3_1 _2563_ (.X(_0368_),
    .A(_0366_),
    .B(_0360_),
    .C(_0362_));
 sg13g2_nor3_1 _2564_ (.A(_0359_),
    .B(_0367_),
    .C(_0368_),
    .Y(_0369_));
 sg13g2_a21o_1 _2565_ (.A2(_0362_),
    .A1(_0360_),
    .B1(_0366_),
    .X(_0370_));
 sg13g2_nand3_1 _2566_ (.B(_0360_),
    .C(_0362_),
    .A(_0366_),
    .Y(_0371_));
 sg13g2_a21oi_1 _2567_ (.A1(_0370_),
    .A2(_0371_),
    .Y(_0372_),
    .B1(\ad.a[29] ));
 sg13g2_o21ai_1 _2568_ (.B1(_0161_),
    .Y(_0373_),
    .A1(_0369_),
    .A2(_0372_));
 sg13g2_inv_1 _2569_ (.Y(_0374_),
    .A(_1356_));
 sg13g2_a22oi_1 _2570_ (.Y(_0375_),
    .B1(net38),
    .B2(\result[21] ),
    .A2(_0374_),
    .A1(_1320_));
 sg13g2_a21oi_1 _2571_ (.A1(_0373_),
    .A2(_0375_),
    .Y(_0039_),
    .B1(net79));
 sg13g2_nor2_1 _2572_ (.A(_1152_),
    .B(_1204_),
    .Y(_0376_));
 sg13g2_xor2_1 _2573_ (.B(_0376_),
    .A(_1175_),
    .X(_0377_));
 sg13g2_a22oi_1 _2574_ (.Y(_0378_),
    .B1(_0840_),
    .B2(_0377_),
    .A2(net42),
    .A1(\result[2] ));
 sg13g2_nor2_1 _2575_ (.A(net76),
    .B(_0378_),
    .Y(_0040_));
 sg13g2_a22oi_1 _2576_ (.Y(_0379_),
    .B1(_0166_),
    .B2(\result[22] ),
    .A2(net36),
    .A1(_0165_));
 sg13g2_inv_1 _2577_ (.Y(_0380_),
    .A(\ad.a[30] ));
 sg13g2_mux2_1 _2578_ (.A0(net10),
    .A1(net36),
    .S(net69),
    .X(_0381_));
 sg13g2_nor2_1 _2579_ (.A(_0834_),
    .B(_0953_),
    .Y(_0382_));
 sg13g2_a21oi_2 _2580_ (.B1(_0382_),
    .Y(_0383_),
    .A2(_0381_),
    .A1(_0934_));
 sg13g2_a21o_1 _2581_ (.A2(_0353_),
    .A1(_0348_),
    .B1(_0346_),
    .X(_0384_));
 sg13g2_inv_1 _2582_ (.Y(_0385_),
    .A(_0366_));
 sg13g2_a21o_1 _2583_ (.A2(_0384_),
    .A1(_0360_),
    .B1(_0385_),
    .X(_0386_));
 sg13g2_and3_1 _2584_ (.X(_0387_),
    .A(_0385_),
    .B(_0360_),
    .C(_0384_));
 sg13g2_buf_1 _2585_ (.A(_0387_),
    .X(_0388_));
 sg13g2_a21oi_1 _2586_ (.A1(_0359_),
    .A2(_0386_),
    .Y(_0389_),
    .B1(_0388_));
 sg13g2_xnor2_1 _2587_ (.Y(_0390_),
    .A(_0383_),
    .B(_0389_));
 sg13g2_xnor2_1 _2588_ (.Y(_0391_),
    .A(_0380_),
    .B(_0390_));
 sg13g2_nand2_1 _2589_ (.Y(_0392_),
    .A(_0161_),
    .B(_0391_));
 sg13g2_a21oi_1 _2590_ (.A1(_0379_),
    .A2(_0392_),
    .Y(_0041_),
    .B1(_1346_));
 sg13g2_nor3_1 _2591_ (.A(_0359_),
    .B(_0383_),
    .C(_0388_),
    .Y(_0393_));
 sg13g2_nor2_1 _2592_ (.A(_0383_),
    .B(_0386_),
    .Y(_0394_));
 sg13g2_nor3_1 _2593_ (.A(_0380_),
    .B(_0388_),
    .C(_0386_),
    .Y(_0395_));
 sg13g2_nand2_1 _2594_ (.Y(_0396_),
    .A(\ad.a[29] ),
    .B(\ad.a[30] ));
 sg13g2_nand2b_1 _2595_ (.Y(_0397_),
    .B(\ad.a[30] ),
    .A_N(_0383_));
 sg13g2_o21ai_1 _2596_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_0388_),
    .A2(_0396_));
 sg13g2_nor4_1 _2597_ (.A(_0393_),
    .B(_0394_),
    .C(_0395_),
    .D(_0398_),
    .Y(_0399_));
 sg13g2_xor2_1 _2598_ (.B(net59),
    .A(_0589_),
    .X(_0400_));
 sg13g2_nand3_1 _2599_ (.B(net11),
    .C(_0400_),
    .A(_0311_),
    .Y(_0401_));
 sg13g2_xor2_1 _2600_ (.B(_0401_),
    .A(\ad.a[31] ),
    .X(_0402_));
 sg13g2_xnor2_1 _2601_ (.Y(_0403_),
    .A(_0399_),
    .B(_0402_));
 sg13g2_nand3_1 _2602_ (.B(net51),
    .C(_0839_),
    .A(\result[23] ),
    .Y(_0404_));
 sg13g2_o21ai_1 _2603_ (.B1(_0404_),
    .Y(_0405_),
    .A1(_0848_),
    .A2(_0403_));
 sg13g2_and2_1 _2604_ (.A(net96),
    .B(_0405_),
    .X(_0042_));
 sg13g2_nor2_1 _2605_ (.A(_1152_),
    .B(_1175_),
    .Y(_0406_));
 sg13g2_or2_1 _2606_ (.X(_0407_),
    .B(_1204_),
    .A(_0406_));
 sg13g2_xnor2_1 _2607_ (.Y(_0408_),
    .A(_1265_),
    .B(_0407_));
 sg13g2_xnor2_1 _2608_ (.Y(_0409_),
    .A(_1268_),
    .B(_0408_));
 sg13g2_a22oi_1 _2609_ (.Y(_0410_),
    .B1(_0840_),
    .B2(_0409_),
    .A2(net42),
    .A1(\result[3] ));
 sg13g2_nor2_1 _2610_ (.A(net76),
    .B(_0410_),
    .Y(_0043_));
 sg13g2_a22oi_1 _2611_ (.Y(_0411_),
    .B1(_1267_),
    .B2(_1269_),
    .A2(_1205_),
    .A1(_1176_));
 sg13g2_xnor2_1 _2612_ (.Y(_0412_),
    .A(_1233_),
    .B(_0411_));
 sg13g2_xnor2_1 _2613_ (.Y(_0413_),
    .A(_1130_),
    .B(_0412_));
 sg13g2_a22oi_1 _2614_ (.Y(_0414_),
    .B1(_0840_),
    .B2(_0413_),
    .A2(net42),
    .A1(\result[4] ));
 sg13g2_nor2_1 _2615_ (.A(net76),
    .B(_0414_),
    .Y(_0044_));
 sg13g2_nand2_1 _2616_ (.Y(_0415_),
    .A(\result[5] ),
    .B(_0843_));
 sg13g2_or3_1 _2617_ (.A(_1236_),
    .B(_1278_),
    .C(_1279_),
    .X(_0416_));
 sg13g2_buf_1 _2618_ (.A(_0416_),
    .X(_0417_));
 sg13g2_xor2_1 _2619_ (.B(_0417_),
    .A(_1262_),
    .X(_0418_));
 sg13g2_xnor2_1 _2620_ (.Y(_0419_),
    .A(_0938_),
    .B(_0418_));
 sg13g2_nand3_1 _2621_ (.B(net56),
    .C(_0419_),
    .A(net44),
    .Y(_0420_));
 sg13g2_buf_1 _2622_ (.A(_0583_),
    .X(_0421_));
 sg13g2_a21oi_1 _2623_ (.A1(_0415_),
    .A2(_0420_),
    .Y(_0045_),
    .B1(net78));
 sg13g2_buf_1 _2624_ (.A(_0583_),
    .X(_0422_));
 sg13g2_nor2_1 _2625_ (.A(_1107_),
    .B(_1109_),
    .Y(_0423_));
 sg13g2_o21ai_1 _2626_ (.B1(\ad.a[5] ),
    .Y(_0424_),
    .A1(_1262_),
    .A2(_0417_));
 sg13g2_inv_1 _2627_ (.Y(_0425_),
    .A(_0424_));
 sg13g2_a21oi_2 _2628_ (.B1(_0425_),
    .Y(_0426_),
    .A2(_0417_),
    .A1(_1262_));
 sg13g2_xor2_1 _2629_ (.B(_0426_),
    .A(_0423_),
    .X(_0427_));
 sg13g2_nor3_1 _2630_ (.A(net43),
    .B(net50),
    .C(_0427_),
    .Y(_0428_));
 sg13g2_a21oi_1 _2631_ (.A1(\result[6] ),
    .A2(net40),
    .Y(_0429_),
    .B1(_0428_));
 sg13g2_nor2_1 _2632_ (.A(net77),
    .B(_0429_),
    .Y(_0046_));
 sg13g2_nand2_1 _2633_ (.Y(_0430_),
    .A(\result[7] ),
    .B(net41));
 sg13g2_and2_1 _2634_ (.A(net62),
    .B(_0952_),
    .X(_0431_));
 sg13g2_a21o_1 _2635_ (.A2(_0963_),
    .A1(net68),
    .B1(_0431_),
    .X(_0432_));
 sg13g2_a21oi_1 _2636_ (.A1(net60),
    .A2(net36),
    .Y(_0433_),
    .B1(_0432_));
 sg13g2_nand2_1 _2637_ (.Y(_0434_),
    .A(_0433_),
    .B(_0426_));
 sg13g2_nor2_1 _2638_ (.A(_0433_),
    .B(_0426_),
    .Y(_0435_));
 sg13g2_a21oi_1 _2639_ (.A1(\ad.a[6] ),
    .A2(_0434_),
    .Y(_0436_),
    .B1(_0435_));
 sg13g2_xor2_1 _2640_ (.B(_0436_),
    .A(_1128_),
    .X(_0437_));
 sg13g2_nand3_1 _2641_ (.B(net56),
    .C(_0437_),
    .A(net44),
    .Y(_0438_));
 sg13g2_a21oi_1 _2642_ (.A1(_0430_),
    .A2(_0438_),
    .Y(_0047_),
    .B1(net78));
 sg13g2_xnor2_1 _2643_ (.Y(_0439_),
    .A(\ad.a[8] ),
    .B(_0937_));
 sg13g2_xnor2_1 _2644_ (.Y(_0440_),
    .A(_1282_),
    .B(_0439_));
 sg13g2_nand2_1 _2645_ (.Y(_0441_),
    .A(net60),
    .B(_0440_));
 sg13g2_nand2_1 _2646_ (.Y(_0442_),
    .A(\result[0] ),
    .B(net52));
 sg13g2_a21oi_1 _2647_ (.A1(_0441_),
    .A2(_0442_),
    .Y(_0443_),
    .B1(net43));
 sg13g2_a21oi_1 _2648_ (.A1(\result[8] ),
    .A2(net40),
    .Y(_0444_),
    .B1(_0443_));
 sg13g2_nor2_1 _2649_ (.A(net77),
    .B(_0444_),
    .Y(_0048_));
 sg13g2_nand2_1 _2650_ (.Y(_0445_),
    .A(\result[9] ),
    .B(_0843_));
 sg13g2_nor2_1 _2651_ (.A(_0929_),
    .B(_1287_),
    .Y(_0446_));
 sg13g2_xnor2_1 _2652_ (.Y(_0447_),
    .A(_1285_),
    .B(_0446_));
 sg13g2_nand2_1 _2653_ (.Y(_0448_),
    .A(\result[1] ),
    .B(net57));
 sg13g2_o21ai_1 _2654_ (.B1(_0448_),
    .Y(_0449_),
    .A1(net50),
    .A2(_0447_));
 sg13g2_nand2_1 _2655_ (.Y(_0450_),
    .A(net44),
    .B(_0449_));
 sg13g2_a21oi_1 _2656_ (.A1(_0445_),
    .A2(_0450_),
    .Y(_0049_),
    .B1(net78));
 sg13g2_or4_1 _2657_ (.A(net36),
    .B(_0356_),
    .C(_0321_),
    .D(_0374_),
    .X(_0451_));
 sg13g2_buf_1 _2658_ (.A(_0451_),
    .X(_0452_));
 sg13g2_nand2_1 _2659_ (.Y(_0453_),
    .A(net71),
    .B(_0452_));
 sg13g2_a21o_1 _2660_ (.A2(_0453_),
    .A1(_0003_),
    .B1(_0168_),
    .X(_0454_));
 sg13g2_o21ai_1 _2661_ (.B1(_0454_),
    .Y(_0455_),
    .A1(net59),
    .A2(_0003_));
 sg13g2_a21oi_1 _2662_ (.A1(net19),
    .A2(_0850_),
    .Y(_0456_),
    .B1(_0452_));
 sg13g2_nor2_1 _2663_ (.A(_1326_),
    .B(_0836_),
    .Y(_0457_));
 sg13g2_a21oi_1 _2664_ (.A1(net71),
    .A2(_0456_),
    .Y(_0458_),
    .B1(_0457_));
 sg13g2_o21ai_1 _2665_ (.B1(net108),
    .Y(_0459_),
    .A1(_0003_),
    .A2(_0458_));
 sg13g2_a21oi_1 _2666_ (.A1(_1355_),
    .A2(_0455_),
    .Y(_0050_),
    .B1(_0459_));
 sg13g2_o21ai_1 _2667_ (.B1(net71),
    .Y(_0460_),
    .A1(net19),
    .A2(_0452_));
 sg13g2_nand2_1 _2668_ (.Y(_0461_),
    .A(net68),
    .B(_0453_));
 sg13g2_a22oi_1 _2669_ (.Y(_0462_),
    .B1(_0461_),
    .B2(net58),
    .A2(_0460_),
    .A1(_0850_));
 sg13g2_nor2_1 _2670_ (.A(_0422_),
    .B(_0462_),
    .Y(_0051_));
 sg13g2_nor2b_1 _2671_ (.A(net19),
    .B_N(_0452_),
    .Y(_0463_));
 sg13g2_nor3_1 _2672_ (.A(net58),
    .B(_0112_),
    .C(_0463_),
    .Y(_0464_));
 sg13g2_o21ai_1 _2673_ (.B1(_0311_),
    .Y(_0465_),
    .A1(net59),
    .A2(_0452_));
 sg13g2_and2_1 _2674_ (.A(_1355_),
    .B(_0465_),
    .X(_0466_));
 sg13g2_nor4_1 _2675_ (.A(net86),
    .B(_1248_),
    .C(_0464_),
    .D(_0466_),
    .Y(_0052_));
 sg13g2_nor2_1 _2676_ (.A(_0612_),
    .B(net55),
    .Y(_0467_));
 sg13g2_nor2_1 _2677_ (.A(net42),
    .B(_0467_),
    .Y(_0468_));
 sg13g2_o21ai_1 _2678_ (.B1(net108),
    .Y(_0469_),
    .A1(_0598_),
    .A2(_0612_));
 sg13g2_a21oi_1 _2679_ (.A1(_0598_),
    .A2(_0468_),
    .Y(_0053_),
    .B1(_0469_));
 sg13g2_buf_1 _2680_ (.A(net60),
    .X(_0470_));
 sg13g2_o21ai_1 _2681_ (.B1(net47),
    .Y(_0471_),
    .A1(net54),
    .A2(_1298_));
 sg13g2_nand2_1 _2682_ (.Y(_0472_),
    .A(\ad.a[10] ),
    .B(_0471_));
 sg13g2_nand3_1 _2683_ (.B(_1298_),
    .C(net39),
    .A(_1315_),
    .Y(_0473_));
 sg13g2_a21oi_1 _2684_ (.A1(_0472_),
    .A2(_0473_),
    .Y(_0054_),
    .B1(net78));
 sg13g2_nand2_1 _2685_ (.Y(_0474_),
    .A(\ad.a[11] ),
    .B(net41));
 sg13g2_nand3_1 _2686_ (.B(net48),
    .C(_1317_),
    .A(net44),
    .Y(_0475_));
 sg13g2_a21oi_1 _2687_ (.A1(_0474_),
    .A2(_0475_),
    .Y(_0055_),
    .B1(net78));
 sg13g2_nor3_1 _2688_ (.A(net43),
    .B(net55),
    .C(_1342_),
    .Y(_0476_));
 sg13g2_a21oi_1 _2689_ (.A1(\ad.a[12] ),
    .A2(net46),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_nor2_1 _2690_ (.A(net77),
    .B(_0477_),
    .Y(_0056_));
 sg13g2_nand2_1 _2691_ (.Y(_0478_),
    .A(\ad.a[13] ),
    .B(net41));
 sg13g2_nand3_1 _2692_ (.B(net48),
    .C(_1364_),
    .A(net44),
    .Y(_0479_));
 sg13g2_a21oi_1 _2693_ (.A1(_0478_),
    .A2(_0479_),
    .Y(_0057_),
    .B1(net78));
 sg13g2_o21ai_1 _2694_ (.B1(net47),
    .Y(_0480_),
    .A1(net54),
    .A2(_0105_));
 sg13g2_nand2_1 _2695_ (.Y(_0481_),
    .A(\ad.a[14] ),
    .B(_0480_));
 sg13g2_nand3b_1 _2696_ (.B(_0105_),
    .C(net39),
    .Y(_0482_),
    .A_N(\ad.a[14] ));
 sg13g2_a21oi_1 _2697_ (.A1(_0481_),
    .A2(_0482_),
    .Y(_0058_),
    .B1(net78));
 sg13g2_a21o_1 _2698_ (.A2(_0128_),
    .A1(_0839_),
    .B1(net45),
    .X(_0483_));
 sg13g2_nand2_2 _2699_ (.Y(_0484_),
    .A(_0845_),
    .B(net57));
 sg13g2_nor3_1 _2700_ (.A(_0111_),
    .B(_0128_),
    .C(_0484_),
    .Y(_0485_));
 sg13g2_a21oi_1 _2701_ (.A1(_0111_),
    .A2(_0483_),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_nor2_1 _2702_ (.A(net77),
    .B(_0486_),
    .Y(_0059_));
 sg13g2_nor3_1 _2703_ (.A(net43),
    .B(net55),
    .C(_0145_),
    .Y(_0487_));
 sg13g2_a21oi_1 _2704_ (.A1(\ad.a[16] ),
    .A2(net46),
    .Y(_0488_),
    .B1(_0487_));
 sg13g2_nor2_1 _2705_ (.A(net77),
    .B(_0488_),
    .Y(_0060_));
 sg13g2_nand2_1 _2706_ (.Y(_0489_),
    .A(\ad.a[17] ),
    .B(net41));
 sg13g2_nand3_1 _2707_ (.B(net48),
    .C(_0160_),
    .A(net44),
    .Y(_0490_));
 sg13g2_a21oi_1 _2708_ (.A1(_0489_),
    .A2(_0490_),
    .Y(_0061_),
    .B1(net78));
 sg13g2_a21o_1 _2709_ (.A2(_0179_),
    .A1(net52),
    .B1(net45),
    .X(_0491_));
 sg13g2_nor3_1 _2710_ (.A(\ad.a[18] ),
    .B(_0484_),
    .C(_0179_),
    .Y(_0492_));
 sg13g2_a21oi_1 _2711_ (.A1(\ad.a[18] ),
    .A2(_0491_),
    .Y(_0493_),
    .B1(_0492_));
 sg13g2_nor2_1 _2712_ (.A(net77),
    .B(_0493_),
    .Y(_0062_));
 sg13g2_o21ai_1 _2713_ (.B1(net51),
    .Y(_0494_),
    .A1(_0470_),
    .A2(_0202_));
 sg13g2_nand2_1 _2714_ (.Y(_0495_),
    .A(\ad.a[19] ),
    .B(_0494_));
 sg13g2_nand3_1 _2715_ (.B(net38),
    .C(_0202_),
    .A(_0182_),
    .Y(_0496_));
 sg13g2_a21oi_1 _2716_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0063_),
    .B1(_0421_));
 sg13g2_xnor2_1 _2717_ (.Y(_0497_),
    .A(_1162_),
    .B(_1167_));
 sg13g2_o21ai_1 _2718_ (.B1(net51),
    .Y(_0498_),
    .A1(net54),
    .A2(_0497_));
 sg13g2_nor2_1 _2719_ (.A(\ad.a[1] ),
    .B(_0484_),
    .Y(_0499_));
 sg13g2_a22oi_1 _2720_ (.Y(_0500_),
    .B1(_0499_),
    .B2(_0497_),
    .A2(_0498_),
    .A1(\ad.a[1] ));
 sg13g2_nor2_1 _2721_ (.A(net77),
    .B(_0500_),
    .Y(_0064_));
 sg13g2_nand2_1 _2722_ (.Y(_0501_),
    .A(\ad.a[20] ),
    .B(net40));
 sg13g2_nand3_1 _2723_ (.B(net48),
    .C(_0227_),
    .A(net47),
    .Y(_0502_));
 sg13g2_a21oi_1 _2724_ (.A1(_0501_),
    .A2(_0502_),
    .Y(_0065_),
    .B1(_0421_));
 sg13g2_a21o_1 _2725_ (.A2(_0242_),
    .A1(net52),
    .B1(net45),
    .X(_0503_));
 sg13g2_nor3_1 _2726_ (.A(_0230_),
    .B(_0484_),
    .C(_0242_),
    .Y(_0504_));
 sg13g2_a21oi_1 _2727_ (.A1(_0230_),
    .A2(_0503_),
    .Y(_0505_),
    .B1(_0504_));
 sg13g2_nor2_1 _2728_ (.A(net77),
    .B(_0505_),
    .Y(_0066_));
 sg13g2_xnor2_1 _2729_ (.Y(_0506_),
    .A(_0250_),
    .B(_0256_));
 sg13g2_a21o_1 _2730_ (.A2(_0506_),
    .A1(net52),
    .B1(net45),
    .X(_0507_));
 sg13g2_nor3_1 _2731_ (.A(_0251_),
    .B(_0484_),
    .C(_0506_),
    .Y(_0508_));
 sg13g2_a21oi_1 _2732_ (.A1(_0251_),
    .A2(_0507_),
    .Y(_0509_),
    .B1(_0508_));
 sg13g2_nor2_1 _2733_ (.A(_0422_),
    .B(_0509_),
    .Y(_0067_));
 sg13g2_nand2_1 _2734_ (.Y(_0510_),
    .A(\ad.a[23] ),
    .B(net40));
 sg13g2_nand3_1 _2735_ (.B(net48),
    .C(_0276_),
    .A(_0162_),
    .Y(_0511_));
 sg13g2_a21oi_1 _2736_ (.A1(_0510_),
    .A2(_0511_),
    .Y(_0068_),
    .B1(net86));
 sg13g2_nor3_1 _2737_ (.A(net43),
    .B(net55),
    .C(_0289_),
    .Y(_0512_));
 sg13g2_a21oi_1 _2738_ (.A1(\ad.a[24] ),
    .A2(net46),
    .Y(_0513_),
    .B1(_0512_));
 sg13g2_nor2_1 _2739_ (.A(net80),
    .B(_0513_),
    .Y(_0069_));
 sg13g2_nor3_1 _2740_ (.A(_1320_),
    .B(net55),
    .C(_0301_),
    .Y(_0514_));
 sg13g2_a21oi_1 _2741_ (.A1(\ad.a[25] ),
    .A2(net46),
    .Y(_0515_),
    .B1(_0514_));
 sg13g2_nor2_1 _2742_ (.A(net80),
    .B(_0515_),
    .Y(_0070_));
 sg13g2_nor3_1 _2743_ (.A(_0842_),
    .B(net55),
    .C(_0318_),
    .Y(_0516_));
 sg13g2_a21oi_1 _2744_ (.A1(\ad.a[26] ),
    .A2(net46),
    .Y(_0517_),
    .B1(_0516_));
 sg13g2_nor2_1 _2745_ (.A(net80),
    .B(_0517_),
    .Y(_0071_));
 sg13g2_nand2_1 _2746_ (.Y(_0518_),
    .A(\ad.a[27] ),
    .B(_1304_));
 sg13g2_nand3_1 _2747_ (.B(_0133_),
    .C(_0339_),
    .A(_0162_),
    .Y(_0519_));
 sg13g2_a21oi_1 _2748_ (.A1(_0518_),
    .A2(_0519_),
    .Y(_0072_),
    .B1(net86));
 sg13g2_nor3_1 _2749_ (.A(_0842_),
    .B(_0259_),
    .C(_0355_),
    .Y(_0520_));
 sg13g2_a21oi_1 _2750_ (.A1(\ad.a[28] ),
    .A2(_0597_),
    .Y(_0521_),
    .B1(_0520_));
 sg13g2_nor2_1 _2751_ (.A(_1303_),
    .B(_0521_),
    .Y(_0073_));
 sg13g2_nand2_1 _2752_ (.Y(_0522_),
    .A(\ad.a[29] ),
    .B(_1304_));
 sg13g2_nor4_1 _2753_ (.A(_0359_),
    .B(_1272_),
    .C(_0367_),
    .D(_0368_),
    .Y(_0523_));
 sg13g2_nand2_1 _2754_ (.Y(_0524_),
    .A(_0359_),
    .B(_0146_));
 sg13g2_a21oi_1 _2755_ (.A1(_0370_),
    .A2(_0371_),
    .Y(_0525_),
    .B1(_0524_));
 sg13g2_nor2_1 _2756_ (.A(_0523_),
    .B(_0525_),
    .Y(_0526_));
 sg13g2_a21oi_1 _2757_ (.A1(_0522_),
    .A2(_0526_),
    .Y(_0074_),
    .B1(_0584_));
 sg13g2_a22oi_1 _2758_ (.Y(_0527_),
    .B1(net38),
    .B2(_0377_),
    .A2(net42),
    .A1(\ad.a[2] ));
 sg13g2_nor2_1 _2759_ (.A(net80),
    .B(_0527_),
    .Y(_0075_));
 sg13g2_o21ai_1 _2760_ (.B1(_0846_),
    .Y(_0528_),
    .A1(_0470_),
    .A2(_0390_));
 sg13g2_nand2_1 _2761_ (.Y(_0529_),
    .A(\ad.a[30] ),
    .B(_0528_));
 sg13g2_nand3_1 _2762_ (.B(_0166_),
    .C(_0390_),
    .A(_0380_),
    .Y(_0530_));
 sg13g2_a21oi_1 _2763_ (.A1(_0529_),
    .A2(_0530_),
    .Y(_0076_),
    .B1(_0584_));
 sg13g2_nor3_1 _2764_ (.A(net45),
    .B(_0259_),
    .C(_0403_),
    .Y(_0531_));
 sg13g2_a21oi_1 _2765_ (.A1(\ad.a[31] ),
    .A2(_0597_),
    .Y(_0532_),
    .B1(_0531_));
 sg13g2_nor2_1 _2766_ (.A(_1303_),
    .B(_0532_),
    .Y(_0077_));
 sg13g2_o21ai_1 _2767_ (.B1(net51),
    .Y(_0533_),
    .A1(net54),
    .A2(_0408_));
 sg13g2_nor2_1 _2768_ (.A(\ad.a[3] ),
    .B(_0484_),
    .Y(_0534_));
 sg13g2_a22oi_1 _2769_ (.Y(_0535_),
    .B1(_0534_),
    .B2(_0408_),
    .A2(_0533_),
    .A1(\ad.a[3] ));
 sg13g2_nor2_1 _2770_ (.A(net80),
    .B(_0535_),
    .Y(_0078_));
 sg13g2_o21ai_1 _2771_ (.B1(net51),
    .Y(_0536_),
    .A1(net54),
    .A2(_0412_));
 sg13g2_nor2_1 _2772_ (.A(\ad.a[4] ),
    .B(_0484_),
    .Y(_0537_));
 sg13g2_a22oi_1 _2773_ (.Y(_0538_),
    .B1(_0537_),
    .B2(_0412_),
    .A2(_0536_),
    .A1(\ad.a[4] ));
 sg13g2_nor2_1 _2774_ (.A(net80),
    .B(_0538_),
    .Y(_0079_));
 sg13g2_o21ai_1 _2775_ (.B1(net51),
    .Y(_0539_),
    .A1(net54),
    .A2(_0418_));
 sg13g2_nand2_1 _2776_ (.Y(_0540_),
    .A(\ad.a[5] ),
    .B(_0539_));
 sg13g2_nand3_1 _2777_ (.B(net39),
    .C(_0418_),
    .A(_0938_),
    .Y(_0541_));
 sg13g2_a21oi_1 _2778_ (.A1(_0540_),
    .A2(_0541_),
    .Y(_0080_),
    .B1(net86));
 sg13g2_xnor2_1 _2779_ (.Y(_0542_),
    .A(_0432_),
    .B(_0426_));
 sg13g2_o21ai_1 _2780_ (.B1(net51),
    .Y(_0543_),
    .A1(net54),
    .A2(_0542_));
 sg13g2_nand2_1 _2781_ (.Y(_0544_),
    .A(\ad.a[6] ),
    .B(_0543_));
 sg13g2_nand3_1 _2782_ (.B(_0147_),
    .C(_0542_),
    .A(_0939_),
    .Y(_0545_));
 sg13g2_a21oi_1 _2783_ (.A1(_0544_),
    .A2(_0545_),
    .Y(_0081_),
    .B1(net86));
 sg13g2_nand2_1 _2784_ (.Y(_0546_),
    .A(\ad.a[7] ),
    .B(net40));
 sg13g2_nand3_1 _2785_ (.B(net48),
    .C(_0437_),
    .A(net47),
    .Y(_0547_));
 sg13g2_a21oi_1 _2786_ (.A1(_0546_),
    .A2(_0547_),
    .Y(_0082_),
    .B1(net86));
 sg13g2_nand2_1 _2787_ (.Y(_0548_),
    .A(\ad.a[8] ),
    .B(net40));
 sg13g2_nand3_1 _2788_ (.B(net48),
    .C(_0440_),
    .A(net47),
    .Y(_0549_));
 sg13g2_a21oi_1 _2789_ (.A1(_0548_),
    .A2(_0549_),
    .Y(_0083_),
    .B1(net86));
 sg13g2_nor3_1 _2790_ (.A(net45),
    .B(net54),
    .C(_0447_),
    .Y(_0550_));
 sg13g2_a21oi_1 _2791_ (.A1(\ad.a[9] ),
    .A2(net46),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_nor2_1 _2792_ (.A(net80),
    .B(_0551_),
    .Y(_0084_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _2794_ (.A(net102),
    .X(net12));
 sg13g2_buf_1 _2795_ (.A(net102),
    .X(net13));
 sg13g2_buf_1 _2796_ (.A(net102),
    .X(net14));
 sg13g2_buf_1 _2797_ (.A(net102),
    .X(net15));
 sg13g2_buf_1 _2798_ (.A(net102),
    .X(net16));
 sg13g2_buf_1 _2799_ (.A(net102),
    .X(net17));
 sg13g2_buf_1 _2800_ (.A(net102),
    .X(net18));
 sg13g2_buf_1 _2801_ (.A(\result[16] ),
    .X(net20));
 sg13g2_buf_1 _2802_ (.A(\result[17] ),
    .X(net21));
 sg13g2_buf_1 _2803_ (.A(\result[18] ),
    .X(net22));
 sg13g2_buf_1 _2804_ (.A(\result[19] ),
    .X(net23));
 sg13g2_buf_1 _2805_ (.A(\result[20] ),
    .X(net24));
 sg13g2_buf_1 _2806_ (.A(\result[21] ),
    .X(net25));
 sg13g2_buf_1 _2807_ (.A(\result[22] ),
    .X(net26));
 sg13g2_buf_1 _2808_ (.A(\result[23] ),
    .X(net27));
 sg13g2_buf_1 _2809_ (.A(\result[24] ),
    .X(net28));
 sg13g2_buf_1 _2810_ (.A(\result[25] ),
    .X(net29));
 sg13g2_buf_1 _2811_ (.A(\result[26] ),
    .X(net30));
 sg13g2_buf_1 _2812_ (.A(\result[27] ),
    .X(net31));
 sg13g2_buf_1 _2813_ (.A(\result[28] ),
    .X(net32));
 sg13g2_buf_1 _2814_ (.A(\result[29] ),
    .X(net33));
 sg13g2_buf_1 _2815_ (.A(\result[30] ),
    .X(net34));
 sg13g2_buf_1 _2816_ (.A(\result[31] ),
    .X(net35));
 sg13g2_dfrbp_1 \inp_a[0]$_DFFE_PN_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net109),
    .D(_0010_),
    .Q_N(_1432_),
    .Q(\inp_a[0] ));
 sg13g2_dfrbp_1 \inp_a[1]$_DFFE_PN_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net110),
    .D(_0011_),
    .Q_N(_1431_),
    .Q(\inp_a[1] ));
 sg13g2_dfrbp_1 \inp_a[2]$_DFFE_PN_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net111),
    .D(_0012_),
    .Q_N(_1430_),
    .Q(\inp_a[2] ));
 sg13g2_dfrbp_1 \inp_a[3]$_DFFE_PN_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net112),
    .D(_0013_),
    .Q_N(_1429_),
    .Q(\inp_a[3] ));
 sg13g2_dfrbp_1 \inp_a[4]$_DFFE_PN_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net113),
    .D(_0014_),
    .Q_N(_1428_),
    .Q(\inp_a[4] ));
 sg13g2_dfrbp_1 \inp_a[5]$_DFFE_PN_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net114),
    .D(_0015_),
    .Q_N(_1427_),
    .Q(\inp_a[5] ));
 sg13g2_dfrbp_1 \inp_a[6]$_DFFE_PN_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net115),
    .D(_0016_),
    .Q_N(_1426_),
    .Q(\inp_a[6] ));
 sg13g2_dfrbp_1 \mode$_DFFE_PN_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net116),
    .D(_0017_),
    .Q_N(net19),
    .Q(mode));
 sg13g2_dfrbp_1 \result[0]$_SDFFE_PN0N_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net117),
    .D(_0018_),
    .Q_N(_1425_),
    .Q(\result[0] ));
 sg13g2_dfrbp_1 \result[10]$_SDFFE_PN0N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net118),
    .D(_0019_),
    .Q_N(_1424_),
    .Q(\result[10] ));
 sg13g2_dfrbp_1 \result[11]$_SDFFE_PN0N_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net119),
    .D(_0020_),
    .Q_N(_1423_),
    .Q(\result[11] ));
 sg13g2_dfrbp_1 \result[12]$_SDFFE_PN0N_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net120),
    .D(_0021_),
    .Q_N(_1422_),
    .Q(\result[12] ));
 sg13g2_dfrbp_1 \result[13]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net121),
    .D(_0022_),
    .Q_N(_1421_),
    .Q(\result[13] ));
 sg13g2_dfrbp_1 \result[14]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net122),
    .D(_0023_),
    .Q_N(_1420_),
    .Q(\result[14] ));
 sg13g2_dfrbp_1 \result[15]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net123),
    .D(_0024_),
    .Q_N(_1419_),
    .Q(\result[15] ));
 sg13g2_dfrbp_1 \result[16]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net124),
    .D(_0025_),
    .Q_N(_1418_),
    .Q(\result[16] ));
 sg13g2_dfrbp_1 \result[17]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net125),
    .D(_0026_),
    .Q_N(_1417_),
    .Q(\result[17] ));
 sg13g2_dfrbp_1 \result[18]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net126),
    .D(_0027_),
    .Q_N(_1416_),
    .Q(\result[18] ));
 sg13g2_dfrbp_1 \result[19]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net127),
    .D(_0028_),
    .Q_N(_1415_),
    .Q(\result[19] ));
 sg13g2_dfrbp_1 \result[1]$_SDFFE_PN0N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net128),
    .D(_0029_),
    .Q_N(_1414_),
    .Q(\result[1] ));
 sg13g2_dfrbp_1 \result[20]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net129),
    .D(_0030_),
    .Q_N(_1413_),
    .Q(\result[20] ));
 sg13g2_dfrbp_1 \result[21]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net130),
    .D(_0031_),
    .Q_N(_1412_),
    .Q(\result[21] ));
 sg13g2_dfrbp_1 \result[22]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net131),
    .D(_0032_),
    .Q_N(_1411_),
    .Q(\result[22] ));
 sg13g2_dfrbp_1 \result[23]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net132),
    .D(_0033_),
    .Q_N(_1410_),
    .Q(\result[23] ));
 sg13g2_dfrbp_1 \result[24]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net133),
    .D(_0034_),
    .Q_N(_1409_),
    .Q(\result[24] ));
 sg13g2_dfrbp_1 \result[25]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net134),
    .D(_0035_),
    .Q_N(_1408_),
    .Q(\result[25] ));
 sg13g2_dfrbp_1 \result[26]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net135),
    .D(_0036_),
    .Q_N(_1407_),
    .Q(\result[26] ));
 sg13g2_dfrbp_1 \result[27]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net136),
    .D(_0037_),
    .Q_N(_1406_),
    .Q(\result[27] ));
 sg13g2_dfrbp_1 \result[28]$_SDFF_PN0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net137),
    .D(_0038_),
    .Q_N(_1405_),
    .Q(\result[28] ));
 sg13g2_dfrbp_1 \result[29]$_SDFF_PN0_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net138),
    .D(_0039_),
    .Q_N(_1404_),
    .Q(\result[29] ));
 sg13g2_dfrbp_1 \result[2]$_SDFFE_PN0N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net139),
    .D(_0040_),
    .Q_N(_1403_),
    .Q(\result[2] ));
 sg13g2_dfrbp_1 \result[30]$_SDFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net140),
    .D(_0041_),
    .Q_N(_1402_),
    .Q(\result[30] ));
 sg13g2_dfrbp_1 \result[31]$_SDFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net141),
    .D(_0042_),
    .Q_N(_1401_),
    .Q(\result[31] ));
 sg13g2_dfrbp_1 \result[3]$_SDFFE_PN0N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net142),
    .D(_0043_),
    .Q_N(_1400_),
    .Q(\result[3] ));
 sg13g2_dfrbp_1 \result[4]$_SDFFE_PN0N_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net143),
    .D(_0044_),
    .Q_N(_1399_),
    .Q(\result[4] ));
 sg13g2_dfrbp_1 \result[5]$_SDFFE_PN0N_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net144),
    .D(_0045_),
    .Q_N(_1398_),
    .Q(\result[5] ));
 sg13g2_dfrbp_1 \result[6]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net145),
    .D(_0046_),
    .Q_N(_1397_),
    .Q(\result[6] ));
 sg13g2_dfrbp_1 \result[7]$_SDFFE_PN0N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net146),
    .D(_0047_),
    .Q_N(_1396_),
    .Q(\result[7] ));
 sg13g2_dfrbp_1 \result[8]$_SDFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net147),
    .D(_0048_),
    .Q_N(_1395_),
    .Q(\result[8] ));
 sg13g2_dfrbp_1 \result[9]$_SDFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net148),
    .D(_0049_),
    .Q_N(_1394_),
    .Q(\result[9] ));
 sg13g2_dfrbp_1 \state[0]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net149),
    .D(_0050_),
    .Q_N(_0003_),
    .Q(\state[0] ));
 sg13g2_dfrbp_1 \state[1]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net150),
    .D(_0051_),
    .Q_N(_1393_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 \state[2]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net151),
    .D(_0052_),
    .Q_N(_0004_),
    .Q(\state[2] ));
 sg13g2_dfrbp_1 \sum[0]$_SDFFE_PN0N_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net152),
    .D(_0053_),
    .Q_N(_1392_),
    .Q(\ad.a[0] ));
 sg13g2_dfrbp_1 \sum[10]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net153),
    .D(_0054_),
    .Q_N(_1391_),
    .Q(\ad.a[10] ));
 sg13g2_dfrbp_1 \sum[11]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net154),
    .D(_0055_),
    .Q_N(_1390_),
    .Q(\ad.a[11] ));
 sg13g2_dfrbp_1 \sum[12]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net155),
    .D(_0056_),
    .Q_N(_1389_),
    .Q(\ad.a[12] ));
 sg13g2_dfrbp_1 \sum[13]$_SDFFE_PN0N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net156),
    .D(_0057_),
    .Q_N(_1388_),
    .Q(\ad.a[13] ));
 sg13g2_dfrbp_1 \sum[14]$_SDFFE_PN0N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net157),
    .D(_0058_),
    .Q_N(_1387_),
    .Q(\ad.a[14] ));
 sg13g2_dfrbp_1 \sum[15]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net158),
    .D(_0059_),
    .Q_N(_1386_),
    .Q(\ad.a[15] ));
 sg13g2_dfrbp_1 \sum[16]$_SDFFE_PN0N_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net159),
    .D(_0060_),
    .Q_N(_0005_),
    .Q(\ad.a[16] ));
 sg13g2_dfrbp_1 \sum[17]$_SDFFE_PN0N_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net160),
    .D(_0061_),
    .Q_N(_0006_),
    .Q(\ad.a[17] ));
 sg13g2_dfrbp_1 \sum[18]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net161),
    .D(_0062_),
    .Q_N(_1385_),
    .Q(\ad.a[18] ));
 sg13g2_dfrbp_1 \sum[19]$_SDFFE_PN0N_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net162),
    .D(_0063_),
    .Q_N(_1384_),
    .Q(\ad.a[19] ));
 sg13g2_dfrbp_1 \sum[1]$_SDFFE_PN0N_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net163),
    .D(_0064_),
    .Q_N(_1383_),
    .Q(\ad.a[1] ));
 sg13g2_dfrbp_1 \sum[20]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net164),
    .D(_0065_),
    .Q_N(_1382_),
    .Q(\ad.a[20] ));
 sg13g2_dfrbp_1 \sum[21]$_SDFFE_PN0N_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net165),
    .D(_0066_),
    .Q_N(_1381_),
    .Q(\ad.a[21] ));
 sg13g2_dfrbp_1 \sum[22]$_SDFFE_PN0N_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net166),
    .D(_0067_),
    .Q_N(_1380_),
    .Q(\ad.a[22] ));
 sg13g2_dfrbp_1 \sum[23]$_SDFFE_PN0N_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net167),
    .D(_0068_),
    .Q_N(_0007_),
    .Q(\ad.a[23] ));
 sg13g2_dfrbp_1 \sum[24]$_SDFFE_PN0N_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net168),
    .D(_0069_),
    .Q_N(_0008_),
    .Q(\ad.a[24] ));
 sg13g2_dfrbp_1 \sum[25]$_SDFFE_PN0N_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net169),
    .D(_0070_),
    .Q_N(_0009_),
    .Q(\ad.a[25] ));
 sg13g2_dfrbp_1 \sum[26]$_SDFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net170),
    .D(_0071_),
    .Q_N(_0000_),
    .Q(\ad.a[26] ));
 sg13g2_dfrbp_1 \sum[27]$_SDFFE_PN0N_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net171),
    .D(_0072_),
    .Q_N(_0001_),
    .Q(\ad.a[27] ));
 sg13g2_dfrbp_1 \sum[28]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net172),
    .D(_0073_),
    .Q_N(_0002_),
    .Q(\ad.a[28] ));
 sg13g2_dfrbp_1 \sum[29]$_SDFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net173),
    .D(_0074_),
    .Q_N(_1379_),
    .Q(\ad.a[29] ));
 sg13g2_dfrbp_1 \sum[2]$_SDFFE_PN0N_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net174),
    .D(_0075_),
    .Q_N(_1378_),
    .Q(\ad.a[2] ));
 sg13g2_dfrbp_1 \sum[30]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net175),
    .D(_0076_),
    .Q_N(_1377_),
    .Q(\ad.a[30] ));
 sg13g2_dfrbp_1 \sum[31]$_SDFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net176),
    .D(_0077_),
    .Q_N(_1376_),
    .Q(\ad.a[31] ));
 sg13g2_dfrbp_1 \sum[3]$_SDFFE_PN0N_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net177),
    .D(_0078_),
    .Q_N(_1375_),
    .Q(\ad.a[3] ));
 sg13g2_dfrbp_1 \sum[4]$_SDFFE_PN0N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net178),
    .D(_0079_),
    .Q_N(_1374_),
    .Q(\ad.a[4] ));
 sg13g2_dfrbp_1 \sum[5]$_SDFFE_PN0N_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net179),
    .D(_0080_),
    .Q_N(_1373_),
    .Q(\ad.a[5] ));
 sg13g2_dfrbp_1 \sum[6]$_SDFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net180),
    .D(_0081_),
    .Q_N(_1372_),
    .Q(\ad.a[6] ));
 sg13g2_dfrbp_1 \sum[7]$_SDFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net181),
    .D(_0082_),
    .Q_N(_1371_),
    .Q(\ad.a[7] ));
 sg13g2_dfrbp_1 \sum[8]$_SDFFE_PN0N_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net182),
    .D(_0083_),
    .Q_N(_1370_),
    .Q(\ad.a[8] ));
 sg13g2_dfrbp_1 \sum[9]$_SDFFE_PN0N_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net183),
    .D(_0084_),
    .Q_N(_1369_),
    .Q(\ad.a[9] ));
 sg13g2_buf_1 input1 (.A(ui_in[1]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[0]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[1]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[2]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[3]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[4]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[5]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[6]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[7]),
    .X(net11));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[0]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[1]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[2]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[4]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[5]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[6]));
 sg13g2_buf_1 output19 (.A(net102),
    .X(uio_oe[7]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[0]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[1]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[2]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[3]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[4]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_out[5]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[6]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[7]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[0]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[1]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[2]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[3]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[4]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uo_out[5]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[6]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout36 (.A(_1106_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0714_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0166_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0147_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1304_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0843_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0165_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1320_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0847_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0842_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0597_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0162_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0133_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0864_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0848_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0846_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0839_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0596_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0470_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0259_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0161_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0838_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0311_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0112_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1272_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0871_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0941_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0934_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0931_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0850_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0834_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0593_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0589_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0168_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1355_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1326_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0958_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0923_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0592_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0588_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0585_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0422_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0421_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1346_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1303_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0921_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0835_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0833_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0591_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0587_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0584_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0579_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0573_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0567_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0564_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0561_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0555_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0599_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0582_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0576_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0571_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0569_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0560_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0558_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0554_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0553_),
    .X(net101));
 sg13g2_buf_1 fanout102 (.A(net19),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0581_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0565_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0562_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0559_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0557_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0556_),
    .X(net108));
 sg13g2_tiehi \inp_a[0]$_DFFE_PN__109  (.L_HI(net109));
 sg13g2_tiehi \inp_a[1]$_DFFE_PN__110  (.L_HI(net110));
 sg13g2_tiehi \inp_a[2]$_DFFE_PN__111  (.L_HI(net111));
 sg13g2_tiehi \inp_a[3]$_DFFE_PN__112  (.L_HI(net112));
 sg13g2_tiehi \inp_a[4]$_DFFE_PN__113  (.L_HI(net113));
 sg13g2_tiehi \inp_a[5]$_DFFE_PN__114  (.L_HI(net114));
 sg13g2_tiehi \inp_a[6]$_DFFE_PN__115  (.L_HI(net115));
 sg13g2_tiehi \mode$_DFFE_PN__116  (.L_HI(net116));
 sg13g2_tiehi \result[0]$_SDFFE_PN0N__117  (.L_HI(net117));
 sg13g2_tiehi \result[10]$_SDFFE_PN0N__118  (.L_HI(net118));
 sg13g2_tiehi \result[11]$_SDFFE_PN0N__119  (.L_HI(net119));
 sg13g2_tiehi \result[12]$_SDFFE_PN0N__120  (.L_HI(net120));
 sg13g2_tiehi \result[13]$_SDFFE_PN0N__121  (.L_HI(net121));
 sg13g2_tiehi \result[14]$_SDFFE_PN0N__122  (.L_HI(net122));
 sg13g2_tiehi \result[15]$_SDFFE_PN0N__123  (.L_HI(net123));
 sg13g2_tiehi \result[16]$_SDFF_PN0__124  (.L_HI(net124));
 sg13g2_tiehi \result[17]$_SDFF_PN0__125  (.L_HI(net125));
 sg13g2_tiehi \result[18]$_SDFF_PN0__126  (.L_HI(net126));
 sg13g2_tiehi \result[19]$_SDFF_PN0__127  (.L_HI(net127));
 sg13g2_tiehi \result[1]$_SDFFE_PN0N__128  (.L_HI(net128));
 sg13g2_tiehi \result[20]$_SDFF_PN0__129  (.L_HI(net129));
 sg13g2_tiehi \result[21]$_SDFF_PN0__130  (.L_HI(net130));
 sg13g2_tiehi \result[22]$_SDFF_PN0__131  (.L_HI(net131));
 sg13g2_tiehi \result[23]$_SDFF_PN0__132  (.L_HI(net132));
 sg13g2_tiehi \result[24]$_SDFF_PN0__133  (.L_HI(net133));
 sg13g2_tiehi \result[25]$_SDFF_PN0__134  (.L_HI(net134));
 sg13g2_tiehi \result[26]$_SDFF_PN0__135  (.L_HI(net135));
 sg13g2_tiehi \result[27]$_SDFF_PN0__136  (.L_HI(net136));
 sg13g2_tiehi \result[28]$_SDFF_PN0__137  (.L_HI(net137));
 sg13g2_tiehi \result[29]$_SDFF_PN0__138  (.L_HI(net138));
 sg13g2_tiehi \result[2]$_SDFFE_PN0N__139  (.L_HI(net139));
 sg13g2_tiehi \result[30]$_SDFF_PN0__140  (.L_HI(net140));
 sg13g2_tiehi \result[31]$_SDFF_PN0__141  (.L_HI(net141));
 sg13g2_tiehi \result[3]$_SDFFE_PN0N__142  (.L_HI(net142));
 sg13g2_tiehi \result[4]$_SDFFE_PN0N__143  (.L_HI(net143));
 sg13g2_tiehi \result[5]$_SDFFE_PN0N__144  (.L_HI(net144));
 sg13g2_tiehi \result[6]$_SDFFE_PN0N__145  (.L_HI(net145));
 sg13g2_tiehi \result[7]$_SDFFE_PN0N__146  (.L_HI(net146));
 sg13g2_tiehi \result[8]$_SDFFE_PN0N__147  (.L_HI(net147));
 sg13g2_tiehi \result[9]$_SDFFE_PN0N__148  (.L_HI(net148));
 sg13g2_tiehi \state[0]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \state[1]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \state[2]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \sum[0]$_SDFFE_PN0N__152  (.L_HI(net152));
 sg13g2_tiehi \sum[10]$_SDFFE_PN0N__153  (.L_HI(net153));
 sg13g2_tiehi \sum[11]$_SDFFE_PN0N__154  (.L_HI(net154));
 sg13g2_tiehi \sum[12]$_SDFFE_PN0N__155  (.L_HI(net155));
 sg13g2_tiehi \sum[13]$_SDFFE_PN0N__156  (.L_HI(net156));
 sg13g2_tiehi \sum[14]$_SDFFE_PN0N__157  (.L_HI(net157));
 sg13g2_tiehi \sum[15]$_SDFFE_PN0N__158  (.L_HI(net158));
 sg13g2_tiehi \sum[16]$_SDFFE_PN0N__159  (.L_HI(net159));
 sg13g2_tiehi \sum[17]$_SDFFE_PN0N__160  (.L_HI(net160));
 sg13g2_tiehi \sum[18]$_SDFFE_PN0N__161  (.L_HI(net161));
 sg13g2_tiehi \sum[19]$_SDFFE_PN0N__162  (.L_HI(net162));
 sg13g2_tiehi \sum[1]$_SDFFE_PN0N__163  (.L_HI(net163));
 sg13g2_tiehi \sum[20]$_SDFFE_PN0N__164  (.L_HI(net164));
 sg13g2_tiehi \sum[21]$_SDFFE_PN0N__165  (.L_HI(net165));
 sg13g2_tiehi \sum[22]$_SDFFE_PN0N__166  (.L_HI(net166));
 sg13g2_tiehi \sum[23]$_SDFFE_PN0N__167  (.L_HI(net167));
 sg13g2_tiehi \sum[24]$_SDFFE_PN0N__168  (.L_HI(net168));
 sg13g2_tiehi \sum[25]$_SDFFE_PN0N__169  (.L_HI(net169));
 sg13g2_tiehi \sum[26]$_SDFFE_PN0N__170  (.L_HI(net170));
 sg13g2_tiehi \sum[27]$_SDFFE_PN0N__171  (.L_HI(net171));
 sg13g2_tiehi \sum[28]$_SDFFE_PN0N__172  (.L_HI(net172));
 sg13g2_tiehi \sum[29]$_SDFFE_PN0N__173  (.L_HI(net173));
 sg13g2_tiehi \sum[2]$_SDFFE_PN0N__174  (.L_HI(net174));
 sg13g2_tiehi \sum[30]$_SDFFE_PN0N__175  (.L_HI(net175));
 sg13g2_tiehi \sum[31]$_SDFFE_PN0N__176  (.L_HI(net176));
 sg13g2_tiehi \sum[3]$_SDFFE_PN0N__177  (.L_HI(net177));
 sg13g2_tiehi \sum[4]$_SDFFE_PN0N__178  (.L_HI(net178));
 sg13g2_tiehi \sum[5]$_SDFFE_PN0N__179  (.L_HI(net179));
 sg13g2_tiehi \sum[6]$_SDFFE_PN0N__180  (.L_HI(net180));
 sg13g2_tiehi \sum[7]$_SDFFE_PN0N__181  (.L_HI(net181));
 sg13g2_tiehi \sum[8]$_SDFFE_PN0N__182  (.L_HI(net182));
 sg13g2_tiehi \sum[9]$_SDFFE_PN0N__183  (.L_HI(net183));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_4 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_170 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_184 ();
 sg13g2_decap_4 FILLER_0_191 ();
 sg13g2_fill_2 FILLER_0_195 ();
 sg13g2_decap_8 FILLER_0_202 ();
 sg13g2_decap_4 FILLER_0_209 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_fill_1 FILLER_0_229 ();
 sg13g2_decap_4 FILLER_0_240 ();
 sg13g2_fill_2 FILLER_0_244 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_340 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_354 ();
 sg13g2_decap_8 FILLER_0_361 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_4 FILLER_0_424 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_4 FILLER_1_119 ();
 sg13g2_fill_1 FILLER_1_123 ();
 sg13g2_decap_4 FILLER_1_132 ();
 sg13g2_fill_2 FILLER_1_136 ();
 sg13g2_decap_4 FILLER_1_143 ();
 sg13g2_fill_1 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_152 ();
 sg13g2_fill_1 FILLER_1_159 ();
 sg13g2_fill_1 FILLER_1_175 ();
 sg13g2_decap_4 FILLER_1_186 ();
 sg13g2_fill_2 FILLER_1_222 ();
 sg13g2_fill_1 FILLER_1_244 ();
 sg13g2_decap_8 FILLER_1_269 ();
 sg13g2_decap_8 FILLER_1_293 ();
 sg13g2_decap_8 FILLER_1_300 ();
 sg13g2_decap_8 FILLER_1_307 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_349 ();
 sg13g2_decap_4 FILLER_1_356 ();
 sg13g2_fill_2 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_decap_8 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_1_415 ();
 sg13g2_decap_8 FILLER_1_422 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_fill_2 FILLER_2_134 ();
 sg13g2_fill_1 FILLER_2_144 ();
 sg13g2_fill_2 FILLER_2_150 ();
 sg13g2_fill_2 FILLER_2_157 ();
 sg13g2_fill_2 FILLER_2_169 ();
 sg13g2_fill_1 FILLER_2_171 ();
 sg13g2_decap_4 FILLER_2_186 ();
 sg13g2_fill_1 FILLER_2_190 ();
 sg13g2_fill_2 FILLER_2_201 ();
 sg13g2_decap_8 FILLER_2_218 ();
 sg13g2_decap_4 FILLER_2_225 ();
 sg13g2_fill_1 FILLER_2_229 ();
 sg13g2_fill_1 FILLER_2_253 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_4 FILLER_2_273 ();
 sg13g2_fill_1 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_292 ();
 sg13g2_fill_2 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_325 ();
 sg13g2_fill_2 FILLER_2_332 ();
 sg13g2_fill_2 FILLER_2_339 ();
 sg13g2_fill_1 FILLER_2_354 ();
 sg13g2_fill_2 FILLER_2_375 ();
 sg13g2_fill_1 FILLER_2_377 ();
 sg13g2_fill_2 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_428 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_4 FILLER_3_126 ();
 sg13g2_fill_2 FILLER_3_135 ();
 sg13g2_fill_1 FILLER_3_137 ();
 sg13g2_decap_4 FILLER_3_148 ();
 sg13g2_decap_8 FILLER_3_163 ();
 sg13g2_decap_8 FILLER_3_170 ();
 sg13g2_fill_1 FILLER_3_177 ();
 sg13g2_decap_4 FILLER_3_193 ();
 sg13g2_fill_1 FILLER_3_197 ();
 sg13g2_fill_2 FILLER_3_214 ();
 sg13g2_fill_1 FILLER_3_221 ();
 sg13g2_fill_1 FILLER_3_226 ();
 sg13g2_fill_1 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_237 ();
 sg13g2_decap_8 FILLER_3_244 ();
 sg13g2_decap_4 FILLER_3_259 ();
 sg13g2_fill_1 FILLER_3_267 ();
 sg13g2_fill_1 FILLER_3_277 ();
 sg13g2_fill_1 FILLER_3_288 ();
 sg13g2_decap_4 FILLER_3_296 ();
 sg13g2_decap_4 FILLER_3_304 ();
 sg13g2_decap_4 FILLER_3_312 ();
 sg13g2_fill_2 FILLER_3_316 ();
 sg13g2_fill_2 FILLER_3_328 ();
 sg13g2_fill_1 FILLER_3_330 ();
 sg13g2_fill_1 FILLER_3_346 ();
 sg13g2_fill_2 FILLER_3_352 ();
 sg13g2_decap_8 FILLER_3_365 ();
 sg13g2_fill_1 FILLER_3_372 ();
 sg13g2_fill_2 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_decap_4 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_421 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_decap_4 FILLER_4_137 ();
 sg13g2_fill_1 FILLER_4_141 ();
 sg13g2_fill_1 FILLER_4_165 ();
 sg13g2_fill_1 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_185 ();
 sg13g2_fill_1 FILLER_4_206 ();
 sg13g2_fill_2 FILLER_4_212 ();
 sg13g2_fill_1 FILLER_4_214 ();
 sg13g2_fill_2 FILLER_4_224 ();
 sg13g2_fill_1 FILLER_4_226 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_fill_2 FILLER_4_238 ();
 sg13g2_fill_1 FILLER_4_240 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_fill_2 FILLER_4_260 ();
 sg13g2_fill_2 FILLER_4_266 ();
 sg13g2_decap_4 FILLER_4_288 ();
 sg13g2_fill_1 FILLER_4_292 ();
 sg13g2_fill_2 FILLER_4_309 ();
 sg13g2_fill_1 FILLER_4_311 ();
 sg13g2_fill_2 FILLER_4_324 ();
 sg13g2_fill_1 FILLER_4_326 ();
 sg13g2_decap_4 FILLER_4_340 ();
 sg13g2_fill_2 FILLER_4_344 ();
 sg13g2_decap_4 FILLER_4_365 ();
 sg13g2_fill_2 FILLER_4_369 ();
 sg13g2_fill_2 FILLER_4_389 ();
 sg13g2_fill_1 FILLER_4_395 ();
 sg13g2_fill_2 FILLER_4_400 ();
 sg13g2_fill_1 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_fill_2 FILLER_5_126 ();
 sg13g2_decap_4 FILLER_5_134 ();
 sg13g2_decap_8 FILLER_5_153 ();
 sg13g2_fill_1 FILLER_5_160 ();
 sg13g2_decap_4 FILLER_5_165 ();
 sg13g2_fill_1 FILLER_5_169 ();
 sg13g2_decap_8 FILLER_5_185 ();
 sg13g2_fill_2 FILLER_5_192 ();
 sg13g2_decap_4 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_218 ();
 sg13g2_fill_1 FILLER_5_227 ();
 sg13g2_fill_2 FILLER_5_232 ();
 sg13g2_fill_2 FILLER_5_239 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_4 FILLER_5_266 ();
 sg13g2_fill_1 FILLER_5_270 ();
 sg13g2_decap_4 FILLER_5_320 ();
 sg13g2_fill_2 FILLER_5_324 ();
 sg13g2_fill_2 FILLER_5_337 ();
 sg13g2_decap_4 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_fill_2 FILLER_5_376 ();
 sg13g2_fill_1 FILLER_5_378 ();
 sg13g2_fill_2 FILLER_5_391 ();
 sg13g2_fill_1 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_4 FILLER_5_424 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_fill_2 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_135 ();
 sg13g2_fill_2 FILLER_6_152 ();
 sg13g2_decap_4 FILLER_6_161 ();
 sg13g2_fill_1 FILLER_6_165 ();
 sg13g2_fill_2 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_187 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_220 ();
 sg13g2_decap_4 FILLER_6_227 ();
 sg13g2_fill_2 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_4 FILLER_6_272 ();
 sg13g2_fill_1 FILLER_6_285 ();
 sg13g2_fill_2 FILLER_6_294 ();
 sg13g2_fill_2 FILLER_6_301 ();
 sg13g2_decap_4 FILLER_6_308 ();
 sg13g2_fill_1 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_316 ();
 sg13g2_fill_2 FILLER_6_323 ();
 sg13g2_decap_4 FILLER_6_331 ();
 sg13g2_fill_1 FILLER_6_335 ();
 sg13g2_decap_4 FILLER_6_341 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_4 FILLER_6_394 ();
 sg13g2_fill_1 FILLER_6_398 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_4 FILLER_6_424 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_fill_2 FILLER_7_133 ();
 sg13g2_fill_1 FILLER_7_135 ();
 sg13g2_decap_8 FILLER_7_151 ();
 sg13g2_decap_8 FILLER_7_158 ();
 sg13g2_decap_4 FILLER_7_165 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_decap_4 FILLER_7_187 ();
 sg13g2_fill_2 FILLER_7_191 ();
 sg13g2_decap_8 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_204 ();
 sg13g2_decap_4 FILLER_7_209 ();
 sg13g2_fill_1 FILLER_7_213 ();
 sg13g2_decap_8 FILLER_7_228 ();
 sg13g2_decap_8 FILLER_7_235 ();
 sg13g2_decap_4 FILLER_7_242 ();
 sg13g2_fill_2 FILLER_7_246 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_fill_1 FILLER_7_274 ();
 sg13g2_fill_2 FILLER_7_280 ();
 sg13g2_fill_2 FILLER_7_286 ();
 sg13g2_decap_8 FILLER_7_293 ();
 sg13g2_decap_8 FILLER_7_300 ();
 sg13g2_fill_2 FILLER_7_307 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_fill_2 FILLER_7_319 ();
 sg13g2_decap_4 FILLER_7_342 ();
 sg13g2_fill_2 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_356 ();
 sg13g2_decap_4 FILLER_7_363 ();
 sg13g2_fill_1 FILLER_7_367 ();
 sg13g2_fill_1 FILLER_7_384 ();
 sg13g2_fill_1 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_71 ();
 sg13g2_decap_8 FILLER_8_78 ();
 sg13g2_decap_8 FILLER_8_85 ();
 sg13g2_fill_2 FILLER_8_92 ();
 sg13g2_fill_1 FILLER_8_94 ();
 sg13g2_fill_1 FILLER_8_121 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_140 ();
 sg13g2_fill_1 FILLER_8_142 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_4 FILLER_8_175 ();
 sg13g2_fill_1 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_191 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_fill_1 FILLER_8_200 ();
 sg13g2_decap_4 FILLER_8_206 ();
 sg13g2_fill_2 FILLER_8_214 ();
 sg13g2_fill_1 FILLER_8_216 ();
 sg13g2_decap_8 FILLER_8_237 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_fill_2 FILLER_8_251 ();
 sg13g2_fill_1 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_292 ();
 sg13g2_decap_8 FILLER_8_299 ();
 sg13g2_fill_1 FILLER_8_306 ();
 sg13g2_decap_8 FILLER_8_311 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_decap_8 FILLER_8_325 ();
 sg13g2_decap_4 FILLER_8_332 ();
 sg13g2_fill_2 FILLER_8_336 ();
 sg13g2_decap_4 FILLER_8_345 ();
 sg13g2_fill_2 FILLER_8_349 ();
 sg13g2_fill_2 FILLER_8_355 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_414 ();
 sg13g2_decap_8 FILLER_8_421 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_4 FILLER_9_42 ();
 sg13g2_fill_1 FILLER_9_46 ();
 sg13g2_decap_8 FILLER_9_51 ();
 sg13g2_decap_4 FILLER_9_58 ();
 sg13g2_fill_1 FILLER_9_62 ();
 sg13g2_fill_2 FILLER_9_93 ();
 sg13g2_fill_1 FILLER_9_95 ();
 sg13g2_fill_2 FILLER_9_108 ();
 sg13g2_decap_8 FILLER_9_166 ();
 sg13g2_fill_1 FILLER_9_173 ();
 sg13g2_fill_1 FILLER_9_188 ();
 sg13g2_fill_2 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_fill_2 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_4 FILLER_9_265 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_decap_4 FILLER_9_279 ();
 sg13g2_decap_4 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_346 ();
 sg13g2_fill_1 FILLER_9_360 ();
 sg13g2_fill_1 FILLER_9_365 ();
 sg13g2_fill_1 FILLER_9_388 ();
 sg13g2_decap_4 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_fill_1 FILLER_9_409 ();
 sg13g2_decap_8 FILLER_9_418 ();
 sg13g2_decap_4 FILLER_9_425 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_4 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_fill_2 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_72 ();
 sg13g2_fill_1 FILLER_10_102 ();
 sg13g2_fill_2 FILLER_10_111 ();
 sg13g2_fill_2 FILLER_10_118 ();
 sg13g2_fill_2 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_142 ();
 sg13g2_decap_8 FILLER_10_149 ();
 sg13g2_fill_1 FILLER_10_156 ();
 sg13g2_decap_4 FILLER_10_169 ();
 sg13g2_fill_2 FILLER_10_173 ();
 sg13g2_fill_2 FILLER_10_182 ();
 sg13g2_fill_1 FILLER_10_184 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_decap_8 FILLER_10_218 ();
 sg13g2_decap_8 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_232 ();
 sg13g2_fill_1 FILLER_10_244 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_fill_2 FILLER_10_265 ();
 sg13g2_fill_1 FILLER_10_267 ();
 sg13g2_fill_1 FILLER_10_298 ();
 sg13g2_decap_4 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_4 FILLER_10_369 ();
 sg13g2_decap_4 FILLER_10_386 ();
 sg13g2_fill_2 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_48 ();
 sg13g2_decap_8 FILLER_11_58 ();
 sg13g2_decap_4 FILLER_11_65 ();
 sg13g2_fill_2 FILLER_11_69 ();
 sg13g2_decap_8 FILLER_11_75 ();
 sg13g2_decap_4 FILLER_11_82 ();
 sg13g2_fill_2 FILLER_11_86 ();
 sg13g2_fill_2 FILLER_11_109 ();
 sg13g2_fill_2 FILLER_11_119 ();
 sg13g2_fill_1 FILLER_11_121 ();
 sg13g2_decap_4 FILLER_11_129 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_fill_2 FILLER_11_145 ();
 sg13g2_decap_8 FILLER_11_156 ();
 sg13g2_decap_4 FILLER_11_163 ();
 sg13g2_fill_2 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_176 ();
 sg13g2_fill_2 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_4 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_fill_1 FILLER_11_238 ();
 sg13g2_fill_2 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_decap_8 FILLER_11_278 ();
 sg13g2_decap_4 FILLER_11_285 ();
 sg13g2_decap_4 FILLER_11_302 ();
 sg13g2_decap_8 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_325 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_decap_4 FILLER_11_343 ();
 sg13g2_fill_2 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_362 ();
 sg13g2_fill_2 FILLER_11_369 ();
 sg13g2_fill_2 FILLER_11_388 ();
 sg13g2_fill_1 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_4 FILLER_12_32 ();
 sg13g2_fill_1 FILLER_12_40 ();
 sg13g2_fill_1 FILLER_12_47 ();
 sg13g2_fill_2 FILLER_12_74 ();
 sg13g2_fill_1 FILLER_12_76 ();
 sg13g2_decap_4 FILLER_12_83 ();
 sg13g2_fill_1 FILLER_12_87 ();
 sg13g2_fill_2 FILLER_12_96 ();
 sg13g2_fill_2 FILLER_12_104 ();
 sg13g2_fill_1 FILLER_12_106 ();
 sg13g2_fill_1 FILLER_12_112 ();
 sg13g2_decap_4 FILLER_12_121 ();
 sg13g2_fill_2 FILLER_12_129 ();
 sg13g2_fill_1 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_140 ();
 sg13g2_fill_1 FILLER_12_150 ();
 sg13g2_fill_1 FILLER_12_159 ();
 sg13g2_fill_1 FILLER_12_164 ();
 sg13g2_fill_1 FILLER_12_179 ();
 sg13g2_fill_2 FILLER_12_185 ();
 sg13g2_fill_2 FILLER_12_205 ();
 sg13g2_fill_1 FILLER_12_207 ();
 sg13g2_fill_1 FILLER_12_211 ();
 sg13g2_fill_2 FILLER_12_223 ();
 sg13g2_decap_8 FILLER_12_229 ();
 sg13g2_decap_4 FILLER_12_236 ();
 sg13g2_fill_2 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_4 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_318 ();
 sg13g2_decap_4 FILLER_12_325 ();
 sg13g2_fill_1 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_339 ();
 sg13g2_fill_2 FILLER_12_346 ();
 sg13g2_fill_1 FILLER_12_348 ();
 sg13g2_fill_2 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_fill_1 FILLER_12_383 ();
 sg13g2_fill_2 FILLER_12_390 ();
 sg13g2_fill_1 FILLER_12_392 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_1 FILLER_12_418 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_15 ();
 sg13g2_fill_1 FILLER_13_43 ();
 sg13g2_decap_8 FILLER_13_50 ();
 sg13g2_decap_8 FILLER_13_57 ();
 sg13g2_decap_8 FILLER_13_64 ();
 sg13g2_decap_8 FILLER_13_71 ();
 sg13g2_fill_2 FILLER_13_78 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_fill_2 FILLER_13_109 ();
 sg13g2_decap_8 FILLER_13_117 ();
 sg13g2_decap_8 FILLER_13_124 ();
 sg13g2_decap_8 FILLER_13_131 ();
 sg13g2_fill_2 FILLER_13_163 ();
 sg13g2_fill_1 FILLER_13_165 ();
 sg13g2_fill_1 FILLER_13_170 ();
 sg13g2_fill_2 FILLER_13_176 ();
 sg13g2_fill_1 FILLER_13_190 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_233 ();
 sg13g2_decap_4 FILLER_13_240 ();
 sg13g2_fill_1 FILLER_13_244 ();
 sg13g2_fill_1 FILLER_13_251 ();
 sg13g2_decap_8 FILLER_13_260 ();
 sg13g2_decap_8 FILLER_13_267 ();
 sg13g2_decap_8 FILLER_13_274 ();
 sg13g2_decap_4 FILLER_13_281 ();
 sg13g2_fill_1 FILLER_13_285 ();
 sg13g2_decap_4 FILLER_13_298 ();
 sg13g2_decap_4 FILLER_13_314 ();
 sg13g2_fill_1 FILLER_13_318 ();
 sg13g2_fill_2 FILLER_13_327 ();
 sg13g2_decap_4 FILLER_13_341 ();
 sg13g2_decap_8 FILLER_13_349 ();
 sg13g2_decap_8 FILLER_13_356 ();
 sg13g2_decap_8 FILLER_13_363 ();
 sg13g2_fill_1 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_4 FILLER_13_391 ();
 sg13g2_fill_1 FILLER_13_395 ();
 sg13g2_fill_2 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_fill_1 FILLER_14_40 ();
 sg13g2_decap_8 FILLER_14_47 ();
 sg13g2_fill_2 FILLER_14_54 ();
 sg13g2_fill_1 FILLER_14_56 ();
 sg13g2_decap_4 FILLER_14_93 ();
 sg13g2_fill_2 FILLER_14_97 ();
 sg13g2_fill_2 FILLER_14_106 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_decap_4 FILLER_14_131 ();
 sg13g2_fill_1 FILLER_14_135 ();
 sg13g2_fill_2 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_152 ();
 sg13g2_decap_8 FILLER_14_157 ();
 sg13g2_decap_4 FILLER_14_164 ();
 sg13g2_fill_2 FILLER_14_173 ();
 sg13g2_fill_2 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_181 ();
 sg13g2_fill_2 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_4 FILLER_14_207 ();
 sg13g2_fill_2 FILLER_14_211 ();
 sg13g2_decap_4 FILLER_14_225 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_4 FILLER_14_266 ();
 sg13g2_decap_4 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_300 ();
 sg13g2_decap_8 FILLER_14_321 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_4 FILLER_14_371 ();
 sg13g2_fill_2 FILLER_14_375 ();
 sg13g2_decap_4 FILLER_14_381 ();
 sg13g2_decap_4 FILLER_14_389 ();
 sg13g2_fill_1 FILLER_14_399 ();
 sg13g2_fill_1 FILLER_14_406 ();
 sg13g2_fill_2 FILLER_14_419 ();
 sg13g2_fill_1 FILLER_14_421 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_22 ();
 sg13g2_decap_8 FILLER_15_29 ();
 sg13g2_fill_1 FILLER_15_40 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_4 FILLER_15_56 ();
 sg13g2_fill_2 FILLER_15_60 ();
 sg13g2_fill_1 FILLER_15_70 ();
 sg13g2_decap_4 FILLER_15_76 ();
 sg13g2_decap_4 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_fill_1 FILLER_15_92 ();
 sg13g2_decap_4 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_4 FILLER_15_141 ();
 sg13g2_decap_8 FILLER_15_149 ();
 sg13g2_decap_8 FILLER_15_156 ();
 sg13g2_fill_2 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_165 ();
 sg13g2_decap_4 FILLER_15_171 ();
 sg13g2_decap_4 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_191 ();
 sg13g2_decap_8 FILLER_15_198 ();
 sg13g2_decap_4 FILLER_15_205 ();
 sg13g2_fill_1 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_226 ();
 sg13g2_fill_2 FILLER_15_233 ();
 sg13g2_fill_1 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_4 FILLER_15_268 ();
 sg13g2_fill_2 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_fill_2 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_4 FILLER_15_348 ();
 sg13g2_fill_2 FILLER_15_372 ();
 sg13g2_fill_1 FILLER_15_374 ();
 sg13g2_decap_4 FILLER_15_379 ();
 sg13g2_fill_1 FILLER_15_383 ();
 sg13g2_fill_2 FILLER_15_390 ();
 sg13g2_fill_1 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_418 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_9 ();
 sg13g2_fill_2 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_48 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_fill_1 FILLER_16_89 ();
 sg13g2_fill_1 FILLER_16_114 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_decap_4 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_fill_2 FILLER_16_149 ();
 sg13g2_fill_1 FILLER_16_160 ();
 sg13g2_fill_2 FILLER_16_165 ();
 sg13g2_fill_2 FILLER_16_176 ();
 sg13g2_fill_1 FILLER_16_178 ();
 sg13g2_decap_8 FILLER_16_208 ();
 sg13g2_decap_8 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_222 ();
 sg13g2_decap_4 FILLER_16_229 ();
 sg13g2_fill_1 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_249 ();
 sg13g2_decap_4 FILLER_16_260 ();
 sg13g2_fill_1 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_291 ();
 sg13g2_decap_4 FILLER_16_296 ();
 sg13g2_decap_4 FILLER_16_323 ();
 sg13g2_fill_2 FILLER_16_327 ();
 sg13g2_fill_2 FILLER_16_350 ();
 sg13g2_decap_4 FILLER_16_356 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_decap_4 FILLER_16_381 ();
 sg13g2_fill_1 FILLER_16_385 ();
 sg13g2_fill_2 FILLER_16_398 ();
 sg13g2_fill_1 FILLER_16_404 ();
 sg13g2_decap_4 FILLER_16_409 ();
 sg13g2_fill_2 FILLER_16_417 ();
 sg13g2_fill_1 FILLER_16_419 ();
 sg13g2_decap_4 FILLER_16_425 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_38 ();
 sg13g2_decap_4 FILLER_17_54 ();
 sg13g2_fill_1 FILLER_17_58 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_103 ();
 sg13g2_decap_8 FILLER_17_121 ();
 sg13g2_fill_2 FILLER_17_128 ();
 sg13g2_decap_8 FILLER_17_134 ();
 sg13g2_fill_2 FILLER_17_141 ();
 sg13g2_fill_2 FILLER_17_176 ();
 sg13g2_decap_4 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_187 ();
 sg13g2_decap_8 FILLER_17_193 ();
 sg13g2_fill_2 FILLER_17_200 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_218 ();
 sg13g2_decap_4 FILLER_17_225 ();
 sg13g2_fill_1 FILLER_17_229 ();
 sg13g2_decap_8 FILLER_17_234 ();
 sg13g2_decap_8 FILLER_17_241 ();
 sg13g2_fill_2 FILLER_17_248 ();
 sg13g2_fill_1 FILLER_17_250 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_decap_4 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_fill_1 FILLER_17_326 ();
 sg13g2_decap_4 FILLER_17_333 ();
 sg13g2_decap_4 FILLER_17_342 ();
 sg13g2_decap_4 FILLER_17_351 ();
 sg13g2_decap_4 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_373 ();
 sg13g2_fill_2 FILLER_17_384 ();
 sg13g2_fill_1 FILLER_17_386 ();
 sg13g2_decap_4 FILLER_17_400 ();
 sg13g2_fill_1 FILLER_17_404 ();
 sg13g2_fill_2 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_422 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_4 FILLER_18_7 ();
 sg13g2_fill_1 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_16 ();
 sg13g2_fill_1 FILLER_18_31 ();
 sg13g2_fill_1 FILLER_18_44 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_55 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_fill_2 FILLER_18_75 ();
 sg13g2_decap_8 FILLER_18_82 ();
 sg13g2_decap_4 FILLER_18_89 ();
 sg13g2_fill_2 FILLER_18_93 ();
 sg13g2_fill_2 FILLER_18_100 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_fill_1 FILLER_18_158 ();
 sg13g2_fill_2 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_184 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_decap_4 FILLER_18_269 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_283 ();
 sg13g2_fill_1 FILLER_18_285 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_1 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_318 ();
 sg13g2_fill_1 FILLER_18_325 ();
 sg13g2_decap_4 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_fill_2 FILLER_18_373 ();
 sg13g2_fill_1 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_412 ();
 sg13g2_decap_8 FILLER_18_419 ();
 sg13g2_decap_4 FILLER_18_426 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_decap_4 FILLER_19_60 ();
 sg13g2_fill_1 FILLER_19_64 ();
 sg13g2_decap_8 FILLER_19_75 ();
 sg13g2_decap_4 FILLER_19_91 ();
 sg13g2_fill_2 FILLER_19_104 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_fill_1 FILLER_19_130 ();
 sg13g2_decap_4 FILLER_19_135 ();
 sg13g2_decap_4 FILLER_19_143 ();
 sg13g2_fill_2 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_decap_8 FILLER_19_157 ();
 sg13g2_decap_4 FILLER_19_164 ();
 sg13g2_decap_8 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_180 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_decap_4 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_206 ();
 sg13g2_decap_4 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_237 ();
 sg13g2_decap_4 FILLER_19_244 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_4 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_decap_4 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_317 ();
 sg13g2_fill_2 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_decap_8 FILLER_19_341 ();
 sg13g2_decap_4 FILLER_19_348 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_fill_1 FILLER_19_369 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_15 ();
 sg13g2_decap_4 FILLER_20_22 ();
 sg13g2_fill_1 FILLER_20_37 ();
 sg13g2_decap_4 FILLER_20_46 ();
 sg13g2_fill_1 FILLER_20_66 ();
 sg13g2_decap_4 FILLER_20_75 ();
 sg13g2_fill_2 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_fill_1 FILLER_20_126 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_decap_8 FILLER_20_169 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_201 ();
 sg13g2_decap_4 FILLER_20_208 ();
 sg13g2_decap_8 FILLER_20_230 ();
 sg13g2_decap_8 FILLER_20_237 ();
 sg13g2_fill_2 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_259 ();
 sg13g2_fill_2 FILLER_20_270 ();
 sg13g2_fill_1 FILLER_20_272 ();
 sg13g2_decap_8 FILLER_20_289 ();
 sg13g2_decap_4 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_313 ();
 sg13g2_fill_2 FILLER_20_320 ();
 sg13g2_fill_1 FILLER_20_334 ();
 sg13g2_fill_2 FILLER_20_367 ();
 sg13g2_decap_4 FILLER_20_373 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_fill_1 FILLER_20_401 ();
 sg13g2_decap_8 FILLER_20_414 ();
 sg13g2_decap_8 FILLER_20_421 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_32 ();
 sg13g2_fill_1 FILLER_21_38 ();
 sg13g2_fill_1 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_55 ();
 sg13g2_decap_8 FILLER_21_62 ();
 sg13g2_decap_8 FILLER_21_69 ();
 sg13g2_fill_2 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_78 ();
 sg13g2_decap_4 FILLER_21_87 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_decap_4 FILLER_21_97 ();
 sg13g2_fill_2 FILLER_21_101 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_129 ();
 sg13g2_fill_2 FILLER_21_136 ();
 sg13g2_decap_4 FILLER_21_143 ();
 sg13g2_fill_2 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_fill_2 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_fill_1 FILLER_21_182 ();
 sg13g2_fill_1 FILLER_21_191 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_207 ();
 sg13g2_fill_2 FILLER_21_222 ();
 sg13g2_fill_2 FILLER_21_228 ();
 sg13g2_fill_1 FILLER_21_230 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_fill_2 FILLER_21_282 ();
 sg13g2_fill_2 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_297 ();
 sg13g2_fill_2 FILLER_21_304 ();
 sg13g2_fill_1 FILLER_21_306 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_fill_1 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_4 FILLER_21_364 ();
 sg13g2_fill_1 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_fill_2 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_414 ();
 sg13g2_decap_8 FILLER_21_421 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_fill_2 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_36 ();
 sg13g2_fill_2 FILLER_22_43 ();
 sg13g2_fill_2 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_103 ();
 sg13g2_decap_4 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_149 ();
 sg13g2_decap_4 FILLER_22_156 ();
 sg13g2_fill_2 FILLER_22_160 ();
 sg13g2_decap_8 FILLER_22_167 ();
 sg13g2_decap_4 FILLER_22_174 ();
 sg13g2_decap_4 FILLER_22_195 ();
 sg13g2_fill_2 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_233 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_decap_4 FILLER_22_252 ();
 sg13g2_fill_2 FILLER_22_264 ();
 sg13g2_fill_2 FILLER_22_271 ();
 sg13g2_fill_2 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_fill_2 FILLER_22_362 ();
 sg13g2_fill_1 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_27 ();
 sg13g2_decap_8 FILLER_23_33 ();
 sg13g2_decap_4 FILLER_23_43 ();
 sg13g2_fill_2 FILLER_23_47 ();
 sg13g2_decap_8 FILLER_23_59 ();
 sg13g2_fill_2 FILLER_23_66 ();
 sg13g2_decap_4 FILLER_23_87 ();
 sg13g2_decap_8 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_108 ();
 sg13g2_decap_8 FILLER_23_117 ();
 sg13g2_fill_2 FILLER_23_124 ();
 sg13g2_fill_2 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_205 ();
 sg13g2_decap_8 FILLER_23_212 ();
 sg13g2_fill_2 FILLER_23_219 ();
 sg13g2_fill_2 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_fill_2 FILLER_23_299 ();
 sg13g2_fill_2 FILLER_23_311 ();
 sg13g2_fill_1 FILLER_23_318 ();
 sg13g2_decap_4 FILLER_23_327 ();
 sg13g2_fill_2 FILLER_23_331 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_fill_2 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_4 FILLER_23_400 ();
 sg13g2_decap_4 FILLER_23_408 ();
 sg13g2_fill_2 FILLER_23_412 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_fill_2 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_31 ();
 sg13g2_decap_8 FILLER_24_38 ();
 sg13g2_fill_1 FILLER_24_45 ();
 sg13g2_decap_8 FILLER_24_59 ();
 sg13g2_fill_1 FILLER_24_66 ();
 sg13g2_decap_4 FILLER_24_71 ();
 sg13g2_fill_2 FILLER_24_79 ();
 sg13g2_decap_8 FILLER_24_85 ();
 sg13g2_decap_4 FILLER_24_92 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_136 ();
 sg13g2_decap_4 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_decap_4 FILLER_24_184 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_194 ();
 sg13g2_decap_4 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_243 ();
 sg13g2_decap_4 FILLER_24_274 ();
 sg13g2_fill_1 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_303 ();
 sg13g2_fill_1 FILLER_24_313 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_2 FILLER_24_389 ();
 sg13g2_fill_1 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_4 FILLER_24_425 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_27 ();
 sg13g2_fill_1 FILLER_25_31 ();
 sg13g2_fill_2 FILLER_25_41 ();
 sg13g2_decap_4 FILLER_25_94 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_fill_1 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_114 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_fill_1 FILLER_25_166 ();
 sg13g2_decap_8 FILLER_25_173 ();
 sg13g2_decap_8 FILLER_25_180 ();
 sg13g2_decap_8 FILLER_25_187 ();
 sg13g2_fill_2 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_219 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_263 ();
 sg13g2_fill_2 FILLER_25_268 ();
 sg13g2_fill_1 FILLER_25_318 ();
 sg13g2_decap_4 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_327 ();
 sg13g2_decap_8 FILLER_25_339 ();
 sg13g2_fill_2 FILLER_25_346 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_4 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_fill_2 FILLER_26_25 ();
 sg13g2_fill_2 FILLER_26_39 ();
 sg13g2_fill_2 FILLER_26_54 ();
 sg13g2_fill_2 FILLER_26_61 ();
 sg13g2_fill_1 FILLER_26_68 ();
 sg13g2_fill_2 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_103 ();
 sg13g2_fill_1 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_112 ();
 sg13g2_decap_4 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_148 ();
 sg13g2_decap_8 FILLER_26_155 ();
 sg13g2_decap_8 FILLER_26_162 ();
 sg13g2_decap_4 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_fill_2 FILLER_26_238 ();
 sg13g2_fill_1 FILLER_26_240 ();
 sg13g2_decap_4 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_fill_2 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_4 FILLER_26_294 ();
 sg13g2_fill_2 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_decap_4 FILLER_26_320 ();
 sg13g2_fill_1 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_350 ();
 sg13g2_decap_4 FILLER_26_356 ();
 sg13g2_fill_1 FILLER_26_360 ();
 sg13g2_decap_4 FILLER_26_365 ();
 sg13g2_fill_1 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_12 ();
 sg13g2_fill_2 FILLER_27_19 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_60 ();
 sg13g2_decap_4 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_74 ();
 sg13g2_decap_4 FILLER_27_80 ();
 sg13g2_decap_4 FILLER_27_88 ();
 sg13g2_fill_2 FILLER_27_97 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_fill_2 FILLER_27_104 ();
 sg13g2_decap_8 FILLER_27_115 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_127 ();
 sg13g2_fill_1 FILLER_27_134 ();
 sg13g2_decap_4 FILLER_27_143 ();
 sg13g2_fill_2 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_155 ();
 sg13g2_decap_4 FILLER_27_162 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_fill_2 FILLER_27_192 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_296 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_303 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_fill_2 FILLER_27_317 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_decap_4 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_8 FILLER_27_403 ();
 sg13g2_decap_8 FILLER_27_410 ();
 sg13g2_decap_8 FILLER_27_417 ();
 sg13g2_decap_4 FILLER_27_424 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_28 ();
 sg13g2_fill_1 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_38 ();
 sg13g2_decap_8 FILLER_28_45 ();
 sg13g2_fill_1 FILLER_28_52 ();
 sg13g2_fill_2 FILLER_28_71 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_decap_4 FILLER_28_86 ();
 sg13g2_fill_1 FILLER_28_90 ();
 sg13g2_decap_8 FILLER_28_96 ();
 sg13g2_decap_8 FILLER_28_108 ();
 sg13g2_decap_8 FILLER_28_115 ();
 sg13g2_decap_8 FILLER_28_122 ();
 sg13g2_decap_4 FILLER_28_129 ();
 sg13g2_fill_2 FILLER_28_133 ();
 sg13g2_decap_4 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_decap_4 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_195 ();
 sg13g2_fill_1 FILLER_28_199 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_226 ();
 sg13g2_decap_4 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_decap_8 FILLER_28_277 ();
 sg13g2_fill_2 FILLER_28_284 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_2 FILLER_28_310 ();
 sg13g2_fill_2 FILLER_28_328 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_fill_1 FILLER_28_361 ();
 sg13g2_fill_2 FILLER_28_395 ();
 sg13g2_fill_2 FILLER_28_402 ();
 sg13g2_decap_4 FILLER_29_31 ();
 sg13g2_decap_8 FILLER_29_39 ();
 sg13g2_fill_2 FILLER_29_46 ();
 sg13g2_fill_2 FILLER_29_68 ();
 sg13g2_fill_1 FILLER_29_101 ();
 sg13g2_decap_8 FILLER_29_138 ();
 sg13g2_fill_2 FILLER_29_145 ();
 sg13g2_fill_2 FILLER_29_155 ();
 sg13g2_fill_2 FILLER_29_163 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_179 ();
 sg13g2_decap_8 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_fill_2 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_205 ();
 sg13g2_fill_2 FILLER_29_229 ();
 sg13g2_decap_4 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_fill_1 FILLER_29_266 ();
 sg13g2_decap_4 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_280 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_fill_2 FILLER_29_305 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_decap_8 FILLER_29_328 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_354 ();
 sg13g2_decap_4 FILLER_29_397 ();
 sg13g2_decap_8 FILLER_29_404 ();
 sg13g2_fill_2 FILLER_29_415 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_11 ();
 sg13g2_decap_4 FILLER_30_18 ();
 sg13g2_fill_2 FILLER_30_31 ();
 sg13g2_decap_8 FILLER_30_37 ();
 sg13g2_fill_2 FILLER_30_44 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_decap_4 FILLER_30_111 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_decap_4 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_decap_8 FILLER_30_209 ();
 sg13g2_fill_2 FILLER_30_216 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_236 ();
 sg13g2_fill_2 FILLER_30_241 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_decap_4 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_decap_4 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_285 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_decap_4 FILLER_30_308 ();
 sg13g2_fill_1 FILLER_30_316 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_359 ();
 sg13g2_decap_4 FILLER_30_367 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_decap_4 FILLER_30_383 ();
 sg13g2_fill_1 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_422 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_30 ();
 sg13g2_fill_2 FILLER_31_39 ();
 sg13g2_fill_1 FILLER_31_41 ();
 sg13g2_fill_2 FILLER_31_47 ();
 sg13g2_fill_2 FILLER_31_54 ();
 sg13g2_fill_1 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_4 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_fill_2 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_142 ();
 sg13g2_decap_8 FILLER_31_148 ();
 sg13g2_fill_1 FILLER_31_155 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_178 ();
 sg13g2_fill_2 FILLER_31_185 ();
 sg13g2_fill_1 FILLER_31_187 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_204 ();
 sg13g2_decap_4 FILLER_31_211 ();
 sg13g2_fill_2 FILLER_31_221 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_decap_4 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_255 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_2 FILLER_31_292 ();
 sg13g2_fill_1 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_decap_4 FILLER_31_314 ();
 sg13g2_fill_2 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_325 ();
 sg13g2_decap_4 FILLER_31_330 ();
 sg13g2_fill_2 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_fill_1 FILLER_31_354 ();
 sg13g2_fill_1 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_4 FILLER_31_381 ();
 sg13g2_fill_1 FILLER_31_385 ();
 sg13g2_fill_1 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_415 ();
 sg13g2_decap_8 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_15 ();
 sg13g2_fill_1 FILLER_32_22 ();
 sg13g2_decap_4 FILLER_32_27 ();
 sg13g2_fill_1 FILLER_32_31 ();
 sg13g2_decap_8 FILLER_32_37 ();
 sg13g2_fill_1 FILLER_32_44 ();
 sg13g2_fill_1 FILLER_32_64 ();
 sg13g2_decap_8 FILLER_32_80 ();
 sg13g2_decap_8 FILLER_32_87 ();
 sg13g2_decap_8 FILLER_32_94 ();
 sg13g2_decap_4 FILLER_32_101 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_111 ();
 sg13g2_fill_2 FILLER_32_117 ();
 sg13g2_fill_1 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_136 ();
 sg13g2_decap_4 FILLER_32_143 ();
 sg13g2_fill_2 FILLER_32_156 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_233 ();
 sg13g2_fill_2 FILLER_32_239 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_fill_2 FILLER_32_279 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_fill_2 FILLER_32_312 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_fill_2 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_346 ();
 sg13g2_decap_8 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_384 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_fill_2 FILLER_32_397 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_fill_2 FILLER_32_409 ();
 sg13g2_decap_8 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_decap_4 FILLER_33_18 ();
 sg13g2_fill_1 FILLER_33_22 ();
 sg13g2_fill_1 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_57 ();
 sg13g2_fill_1 FILLER_33_59 ();
 sg13g2_decap_4 FILLER_33_65 ();
 sg13g2_fill_2 FILLER_33_69 ();
 sg13g2_decap_8 FILLER_33_76 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_fill_2 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_153 ();
 sg13g2_decap_4 FILLER_33_170 ();
 sg13g2_fill_1 FILLER_33_174 ();
 sg13g2_fill_2 FILLER_33_188 ();
 sg13g2_fill_1 FILLER_33_190 ();
 sg13g2_decap_8 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_226 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_decap_4 FILLER_33_239 ();
 sg13g2_fill_1 FILLER_33_243 ();
 sg13g2_decap_8 FILLER_33_248 ();
 sg13g2_decap_4 FILLER_33_255 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_decap_4 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_292 ();
 sg13g2_decap_8 FILLER_33_299 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_fill_2 FILLER_33_319 ();
 sg13g2_fill_1 FILLER_33_321 ();
 sg13g2_decap_8 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_349 ();
 sg13g2_fill_2 FILLER_33_356 ();
 sg13g2_decap_4 FILLER_33_363 ();
 sg13g2_decap_4 FILLER_33_376 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_decap_4 FILLER_33_398 ();
 sg13g2_fill_2 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_31 ();
 sg13g2_decap_8 FILLER_34_38 ();
 sg13g2_decap_4 FILLER_34_45 ();
 sg13g2_fill_2 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_68 ();
 sg13g2_fill_2 FILLER_34_77 ();
 sg13g2_decap_4 FILLER_34_89 ();
 sg13g2_decap_8 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_decap_8 FILLER_34_122 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_fill_1 FILLER_34_142 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_fill_2 FILLER_34_161 ();
 sg13g2_fill_1 FILLER_34_163 ();
 sg13g2_fill_2 FILLER_34_177 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_203 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_decap_4 FILLER_34_292 ();
 sg13g2_fill_2 FILLER_34_296 ();
 sg13g2_fill_1 FILLER_34_307 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_fill_1 FILLER_34_352 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_decap_4 FILLER_34_375 ();
 sg13g2_fill_2 FILLER_34_379 ();
 sg13g2_fill_2 FILLER_34_385 ();
 sg13g2_fill_1 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_418 ();
 sg13g2_decap_4 FILLER_34_425 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_11 ();
 sg13g2_decap_4 FILLER_35_18 ();
 sg13g2_fill_1 FILLER_35_22 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_4 FILLER_35_35 ();
 sg13g2_decap_4 FILLER_35_51 ();
 sg13g2_fill_2 FILLER_35_55 ();
 sg13g2_decap_8 FILLER_35_76 ();
 sg13g2_decap_4 FILLER_35_83 ();
 sg13g2_fill_1 FILLER_35_87 ();
 sg13g2_decap_4 FILLER_35_93 ();
 sg13g2_fill_1 FILLER_35_97 ();
 sg13g2_fill_1 FILLER_35_124 ();
 sg13g2_decap_8 FILLER_35_151 ();
 sg13g2_fill_1 FILLER_35_166 ();
 sg13g2_fill_1 FILLER_35_171 ();
 sg13g2_fill_1 FILLER_35_177 ();
 sg13g2_fill_1 FILLER_35_189 ();
 sg13g2_decap_4 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_35_202 ();
 sg13g2_fill_2 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_223 ();
 sg13g2_decap_8 FILLER_35_230 ();
 sg13g2_decap_8 FILLER_35_237 ();
 sg13g2_decap_8 FILLER_35_244 ();
 sg13g2_decap_8 FILLER_35_251 ();
 sg13g2_decap_4 FILLER_35_258 ();
 sg13g2_fill_1 FILLER_35_262 ();
 sg13g2_fill_1 FILLER_35_272 ();
 sg13g2_decap_4 FILLER_35_277 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_303 ();
 sg13g2_decap_8 FILLER_35_318 ();
 sg13g2_decap_8 FILLER_35_325 ();
 sg13g2_fill_2 FILLER_35_332 ();
 sg13g2_fill_2 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_345 ();
 sg13g2_decap_4 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_fill_1 FILLER_35_380 ();
 sg13g2_decap_4 FILLER_35_402 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_412 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_decap_8 FILLER_36_26 ();
 sg13g2_decap_8 FILLER_36_33 ();
 sg13g2_decap_4 FILLER_36_45 ();
 sg13g2_fill_1 FILLER_36_49 ();
 sg13g2_fill_2 FILLER_36_62 ();
 sg13g2_fill_1 FILLER_36_64 ();
 sg13g2_decap_8 FILLER_36_73 ();
 sg13g2_decap_4 FILLER_36_80 ();
 sg13g2_decap_8 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_103 ();
 sg13g2_fill_1 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_117 ();
 sg13g2_decap_8 FILLER_36_124 ();
 sg13g2_decap_4 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_156 ();
 sg13g2_decap_8 FILLER_36_163 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_229 ();
 sg13g2_fill_1 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_decap_4 FILLER_36_298 ();
 sg13g2_fill_2 FILLER_36_302 ();
 sg13g2_decap_4 FILLER_36_330 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_362 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_fill_2 FILLER_36_370 ();
 sg13g2_fill_1 FILLER_36_372 ();
 sg13g2_fill_2 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_fill_2 FILLER_36_398 ();
 sg13g2_fill_1 FILLER_36_400 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_fill_2 FILLER_37_41 ();
 sg13g2_fill_2 FILLER_37_47 ();
 sg13g2_fill_1 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_54 ();
 sg13g2_decap_4 FILLER_37_60 ();
 sg13g2_fill_1 FILLER_37_72 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_decap_4 FILLER_37_103 ();
 sg13g2_fill_2 FILLER_37_107 ();
 sg13g2_fill_1 FILLER_37_140 ();
 sg13g2_fill_1 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_184 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_276 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_decap_4 FILLER_37_340 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_decap_4 FILLER_37_354 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_fill_2 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_19 ();
 sg13g2_fill_2 FILLER_38_26 ();
 sg13g2_decap_4 FILLER_38_58 ();
 sg13g2_fill_2 FILLER_38_62 ();
 sg13g2_fill_2 FILLER_38_90 ();
 sg13g2_fill_2 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_122 ();
 sg13g2_fill_1 FILLER_38_131 ();
 sg13g2_decap_4 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_155 ();
 sg13g2_decap_4 FILLER_38_192 ();
 sg13g2_fill_2 FILLER_38_196 ();
 sg13g2_decap_4 FILLER_38_202 ();
 sg13g2_fill_1 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_211 ();
 sg13g2_fill_2 FILLER_38_216 ();
 sg13g2_fill_1 FILLER_38_218 ();
 sg13g2_decap_4 FILLER_38_231 ();
 sg13g2_fill_1 FILLER_38_251 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_347 ();
 sg13g2_decap_4 FILLER_38_353 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_fill_1 FILLER_38_369 ();
 sg13g2_fill_1 FILLER_38_374 ();
 sg13g2_fill_2 FILLER_38_383 ();
 sg13g2_fill_1 FILLER_38_385 ();
 sg13g2_fill_2 FILLER_38_390 ();
 sg13g2_fill_2 FILLER_38_396 ();
 sg13g2_fill_1 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_decap_4 FILLER_38_411 ();
 sg13g2_decap_8 FILLER_38_419 ();
 sg13g2_decap_4 FILLER_38_426 ();
endmodule
