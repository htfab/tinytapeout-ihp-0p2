module tt_um_jayjaywong12 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire clknet_leaf_0_clk;
 wire net182;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[16][0] ;
 wire \mem[16][1] ;
 wire \mem[16][2] ;
 wire \mem[16][3] ;
 wire \mem[17][0] ;
 wire \mem[17][1] ;
 wire \mem[17][2] ;
 wire \mem[17][3] ;
 wire \mem[18][0] ;
 wire \mem[18][1] ;
 wire \mem[18][2] ;
 wire \mem[18][3] ;
 wire \mem[19][0] ;
 wire \mem[19][1] ;
 wire \mem[19][2] ;
 wire \mem[19][3] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[20][0] ;
 wire \mem[20][1] ;
 wire \mem[20][2] ;
 wire \mem[20][3] ;
 wire \mem[21][0] ;
 wire \mem[21][1] ;
 wire \mem[21][2] ;
 wire \mem[21][3] ;
 wire \mem[22][0] ;
 wire \mem[22][1] ;
 wire \mem[22][2] ;
 wire \mem[22][3] ;
 wire \mem[23][0] ;
 wire \mem[23][1] ;
 wire \mem[23][2] ;
 wire \mem[23][3] ;
 wire \mem[24][0] ;
 wire \mem[24][1] ;
 wire \mem[24][2] ;
 wire \mem[24][3] ;
 wire \mem[25][0] ;
 wire \mem[25][1] ;
 wire \mem[25][2] ;
 wire \mem[25][3] ;
 wire \mem[26][0] ;
 wire \mem[26][1] ;
 wire \mem[26][2] ;
 wire \mem[26][3] ;
 wire \mem[27][0] ;
 wire \mem[27][1] ;
 wire \mem[27][2] ;
 wire \mem[27][3] ;
 wire \mem[28][0] ;
 wire \mem[28][1] ;
 wire \mem[28][2] ;
 wire \mem[28][3] ;
 wire \mem[29][0] ;
 wire \mem[29][1] ;
 wire \mem[29][2] ;
 wire \mem[29][3] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[30][0] ;
 wire \mem[30][1] ;
 wire \mem[30][2] ;
 wire \mem[30][3] ;
 wire \mem[31][0] ;
 wire \mem[31][1] ;
 wire \mem[31][2] ;
 wire \mem[31][3] ;
 wire \mem[32][0] ;
 wire \mem[32][1] ;
 wire \mem[32][2] ;
 wire \mem[32][3] ;
 wire \mem[35][0] ;
 wire \mem[35][1] ;
 wire \mem[35][2] ;
 wire \mem[35][3] ;
 wire \mem[36][0] ;
 wire \mem[36][1] ;
 wire \mem[36][2] ;
 wire \mem[36][3] ;
 wire \mem[37][0] ;
 wire \mem[37][1] ;
 wire \mem[37][2] ;
 wire \mem[37][3] ;
 wire \mem[38][0] ;
 wire \mem[38][1] ;
 wire \mem[38][2] ;
 wire \mem[38][3] ;
 wire \mem[39][0] ;
 wire \mem[39][1] ;
 wire \mem[39][2] ;
 wire \mem[39][3] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[40][0] ;
 wire \mem[40][1] ;
 wire \mem[40][2] ;
 wire \mem[40][3] ;
 wire \mem[41][0] ;
 wire \mem[41][1] ;
 wire \mem[41][2] ;
 wire \mem[41][3] ;
 wire \mem[42][0] ;
 wire \mem[42][1] ;
 wire \mem[42][2] ;
 wire \mem[42][3] ;
 wire \mem[43][0] ;
 wire \mem[43][1] ;
 wire \mem[43][2] ;
 wire \mem[43][3] ;
 wire \mem[44][0] ;
 wire \mem[44][1] ;
 wire \mem[44][2] ;
 wire \mem[44][3] ;
 wire \mem[45][0] ;
 wire \mem[45][1] ;
 wire \mem[45][2] ;
 wire \mem[45][3] ;
 wire \mem[46][0] ;
 wire \mem[46][1] ;
 wire \mem[46][2] ;
 wire \mem[46][3] ;
 wire \mem[47][0] ;
 wire \mem[47][1] ;
 wire \mem[47][2] ;
 wire \mem[47][3] ;
 wire \mem[48][0] ;
 wire \mem[48][1] ;
 wire \mem[48][2] ;
 wire \mem[48][3] ;
 wire \mem[49][0] ;
 wire \mem[49][1] ;
 wire \mem[49][2] ;
 wire \mem[49][3] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[50][0] ;
 wire \mem[50][1] ;
 wire \mem[50][2] ;
 wire \mem[50][3] ;
 wire \mem[51][0] ;
 wire \mem[51][1] ;
 wire \mem[51][2] ;
 wire \mem[51][3] ;
 wire \mem[52][0] ;
 wire \mem[52][1] ;
 wire \mem[52][2] ;
 wire \mem[52][3] ;
 wire \mem[53][0] ;
 wire \mem[53][1] ;
 wire \mem[53][2] ;
 wire \mem[53][3] ;
 wire \mem[54][0] ;
 wire \mem[54][1] ;
 wire \mem[54][2] ;
 wire \mem[54][3] ;
 wire \mem[55][0] ;
 wire \mem[55][1] ;
 wire \mem[55][2] ;
 wire \mem[55][3] ;
 wire \mem[56][0] ;
 wire \mem[56][1] ;
 wire \mem[56][2] ;
 wire \mem[56][3] ;
 wire \mem[57][0] ;
 wire \mem[57][1] ;
 wire \mem[57][2] ;
 wire \mem[57][3] ;
 wire \mem[58][0] ;
 wire \mem[58][1] ;
 wire \mem[58][2] ;
 wire \mem[58][3] ;
 wire \mem[59][0] ;
 wire \mem[59][1] ;
 wire \mem[59][2] ;
 wire \mem[59][3] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[60][0] ;
 wire \mem[60][1] ;
 wire \mem[60][2] ;
 wire \mem[60][3] ;
 wire \mem[61][0] ;
 wire \mem[61][1] ;
 wire \mem[61][2] ;
 wire \mem[61][3] ;
 wire \mem[62][0] ;
 wire \mem[62][1] ;
 wire \mem[62][2] ;
 wire \mem[62][3] ;
 wire \mem[63][0] ;
 wire \mem[63][1] ;
 wire \mem[63][2] ;
 wire \mem[63][3] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \prev_acc[0] ;
 wire \prev_acc[1] ;
 wire \prev_acc[2] ;
 wire \prev_acc[3] ;
 wire \prev_acc[4] ;
 wire \prev_acc[5] ;
 wire \prev_acc[6] ;
 wire \prev_acc[7] ;
 wire \products[0][0] ;
 wire \products[0][1] ;
 wire \products[0][2] ;
 wire \products[0][3] ;
 wire \products[0][4] ;
 wire \products[0][5] ;
 wire \products[0][6] ;
 wire \products[0][7] ;
 wire \products[10][0] ;
 wire \products[10][1] ;
 wire \products[10][2] ;
 wire \products[10][3] ;
 wire \products[10][4] ;
 wire \products[10][5] ;
 wire \products[10][6] ;
 wire \products[10][7] ;
 wire \products[11][0] ;
 wire \products[11][1] ;
 wire \products[11][2] ;
 wire \products[11][3] ;
 wire \products[11][4] ;
 wire \products[11][5] ;
 wire \products[11][6] ;
 wire \products[11][7] ;
 wire \products[12][0] ;
 wire \products[12][1] ;
 wire \products[12][2] ;
 wire \products[12][3] ;
 wire \products[12][4] ;
 wire \products[12][5] ;
 wire \products[12][6] ;
 wire \products[12][7] ;
 wire \products[13][0] ;
 wire \products[13][1] ;
 wire \products[13][2] ;
 wire \products[13][3] ;
 wire \products[13][4] ;
 wire \products[13][5] ;
 wire \products[13][6] ;
 wire \products[13][7] ;
 wire \products[14][0] ;
 wire \products[14][1] ;
 wire \products[14][2] ;
 wire \products[14][3] ;
 wire \products[14][4] ;
 wire \products[14][5] ;
 wire \products[14][6] ;
 wire \products[14][7] ;
 wire \products[15][0] ;
 wire \products[15][1] ;
 wire \products[15][2] ;
 wire \products[15][3] ;
 wire \products[15][4] ;
 wire \products[15][5] ;
 wire \products[15][6] ;
 wire \products[15][7] ;
 wire \products[1][0] ;
 wire \products[1][1] ;
 wire \products[1][2] ;
 wire \products[1][3] ;
 wire \products[1][4] ;
 wire \products[1][5] ;
 wire \products[1][6] ;
 wire \products[1][7] ;
 wire \products[2][0] ;
 wire \products[2][1] ;
 wire \products[2][2] ;
 wire \products[2][3] ;
 wire \products[2][4] ;
 wire \products[2][5] ;
 wire \products[2][6] ;
 wire \products[2][7] ;
 wire \products[3][0] ;
 wire \products[3][1] ;
 wire \products[3][2] ;
 wire \products[3][3] ;
 wire \products[3][4] ;
 wire \products[3][5] ;
 wire \products[3][6] ;
 wire \products[3][7] ;
 wire \products[4][0] ;
 wire \products[4][1] ;
 wire \products[4][2] ;
 wire \products[4][3] ;
 wire \products[4][4] ;
 wire \products[4][5] ;
 wire \products[4][6] ;
 wire \products[4][7] ;
 wire \products[5][0] ;
 wire \products[5][1] ;
 wire \products[5][2] ;
 wire \products[5][3] ;
 wire \products[5][4] ;
 wire \products[5][5] ;
 wire \products[5][6] ;
 wire \products[5][7] ;
 wire \products[6][0] ;
 wire \products[6][1] ;
 wire \products[6][2] ;
 wire \products[6][3] ;
 wire \products[6][4] ;
 wire \products[6][5] ;
 wire \products[6][6] ;
 wire \products[6][7] ;
 wire \products[7][0] ;
 wire \products[7][1] ;
 wire \products[7][2] ;
 wire \products[7][3] ;
 wire \products[7][4] ;
 wire \products[7][5] ;
 wire \products[7][6] ;
 wire \products[7][7] ;
 wire \products[8][0] ;
 wire \products[8][1] ;
 wire \products[8][2] ;
 wire \products[8][3] ;
 wire \products[8][4] ;
 wire \products[8][5] ;
 wire \products[8][6] ;
 wire \products[8][7] ;
 wire \products[9][0] ;
 wire \products[9][1] ;
 wire \products[9][2] ;
 wire \products[9][3] ;
 wire \products[9][4] ;
 wire \products[9][5] ;
 wire \products[9][6] ;
 wire \products[9][7] ;
 wire read_operation;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_inv_1 _3190_ (.Y(_2605_),
    .A(net2));
 sg13g2_buf_1 _3191_ (.A(rst_n),
    .X(_2606_));
 sg13g2_buf_1 _3192_ (.A(net15),
    .X(_2607_));
 sg13g2_buf_1 _3193_ (.A(net16),
    .X(_2608_));
 sg13g2_nand2_1 _3194_ (.Y(_2609_),
    .A(_2607_),
    .B(_2608_));
 sg13g2_nand4_1 _3195_ (.B(_2605_),
    .C(_2606_),
    .A(net1),
    .Y(_2610_),
    .D(_2609_));
 sg13g2_buf_1 _3196_ (.A(_2610_),
    .X(_2611_));
 sg13g2_buf_1 _3197_ (.A(_2611_),
    .X(_2612_));
 sg13g2_xor2_1 _3198_ (.B(\products[9][0] ),
    .A(\products[8][0] ),
    .X(_2613_));
 sg13g2_xnor2_1 _3199_ (.Y(_2614_),
    .A(\products[14][0] ),
    .B(\products[1][0] ));
 sg13g2_xnor2_1 _3200_ (.Y(_2615_),
    .A(\products[15][0] ),
    .B(_2614_));
 sg13g2_xnor2_1 _3201_ (.Y(_2616_),
    .A(\products[11][0] ),
    .B(\products[13][0] ));
 sg13g2_xnor2_1 _3202_ (.Y(_2617_),
    .A(\products[12][0] ),
    .B(_2616_));
 sg13g2_buf_1 _3203_ (.A(\prev_acc[0] ),
    .X(_2618_));
 sg13g2_xnor2_1 _3204_ (.Y(_2619_),
    .A(_2618_),
    .B(\products[10][0] ));
 sg13g2_xnor2_1 _3205_ (.Y(_2620_),
    .A(\products[0][0] ),
    .B(_2619_));
 sg13g2_xor2_1 _3206_ (.B(_2620_),
    .A(_2617_),
    .X(_2621_));
 sg13g2_xor2_1 _3207_ (.B(_2621_),
    .A(_2615_),
    .X(_2622_));
 sg13g2_xnor2_1 _3208_ (.Y(_2623_),
    .A(\products[5][0] ),
    .B(\products[7][0] ));
 sg13g2_xnor2_1 _3209_ (.Y(_2624_),
    .A(\products[6][0] ),
    .B(_2623_));
 sg13g2_xnor2_1 _3210_ (.Y(_2625_),
    .A(\products[2][0] ),
    .B(\products[4][0] ));
 sg13g2_xnor2_1 _3211_ (.Y(_2626_),
    .A(\products[3][0] ),
    .B(_2625_));
 sg13g2_xor2_1 _3212_ (.B(_2626_),
    .A(_2624_),
    .X(_2627_));
 sg13g2_xor2_1 _3213_ (.B(_2627_),
    .A(_2622_),
    .X(_2628_));
 sg13g2_xnor2_1 _3214_ (.Y(_2629_),
    .A(_2613_),
    .B(_2628_));
 sg13g2_nor2_1 _3215_ (.A(net3),
    .B(_2612_),
    .Y(_2630_));
 sg13g2_a21oi_1 _3216_ (.A1(_2612_),
    .A2(_2629_),
    .Y(_2631_),
    .B1(_2630_));
 sg13g2_buf_1 _3217_ (.A(_2631_),
    .X(_2632_));
 sg13g2_buf_1 _3218_ (.A(net52),
    .X(_2633_));
 sg13g2_buf_1 _3219_ (.A(\mem[0][0] ),
    .X(_2634_));
 sg13g2_buf_2 _3220_ (.A(ui_in[0]),
    .X(_2635_));
 sg13g2_buf_1 _3221_ (.A(ui_in[1]),
    .X(_2636_));
 sg13g2_buf_1 _3222_ (.A(ui_in[2]),
    .X(_2637_));
 sg13g2_nor4_1 _3223_ (.A(_2635_),
    .B(_2636_),
    .C(_2637_),
    .D(net58),
    .Y(_2638_));
 sg13g2_buf_4 _3224_ (.X(_2639_),
    .A(_2638_));
 sg13g2_buf_1 _3225_ (.A(ui_in[3]),
    .X(_2640_));
 sg13g2_buf_1 _3226_ (.A(ui_in[4]),
    .X(_2641_));
 sg13g2_buf_1 _3227_ (.A(ui_in[5]),
    .X(_2642_));
 sg13g2_nor4_1 _3228_ (.A(_2640_),
    .B(net177),
    .C(net176),
    .D(net58),
    .Y(_2643_));
 sg13g2_buf_4 _3229_ (.X(_2644_),
    .A(_2643_));
 sg13g2_nand2_2 _3230_ (.Y(_2645_),
    .A(_2639_),
    .B(_2644_));
 sg13g2_mux2_1 _3231_ (.A0(net51),
    .A1(net175),
    .S(_2645_),
    .X(_0001_));
 sg13g2_and4_1 _3232_ (.A(net1),
    .B(_2605_),
    .C(_2606_),
    .D(_2609_),
    .X(_2646_));
 sg13g2_buf_2 _3233_ (.A(_2646_),
    .X(_2647_));
 sg13g2_nand2_1 _3234_ (.Y(_2648_),
    .A(_2617_),
    .B(_2620_));
 sg13g2_nand2_1 _3235_ (.Y(_2649_),
    .A(\products[11][0] ),
    .B(\products[13][0] ));
 sg13g2_o21ai_1 _3236_ (.B1(\products[12][0] ),
    .Y(_2650_),
    .A1(\products[11][0] ),
    .A2(\products[13][0] ));
 sg13g2_nand2_1 _3237_ (.Y(_2651_),
    .A(\products[14][0] ),
    .B(\products[1][0] ));
 sg13g2_o21ai_1 _3238_ (.B1(\products[15][0] ),
    .Y(_2652_),
    .A1(\products[14][0] ),
    .A2(\products[1][0] ));
 sg13g2_a22oi_1 _3239_ (.Y(_2653_),
    .B1(_2651_),
    .B2(_2652_),
    .A2(_2650_),
    .A1(_2649_));
 sg13g2_and4_1 _3240_ (.A(_2649_),
    .B(_2650_),
    .C(_2651_),
    .D(_2652_),
    .X(_2654_));
 sg13g2_buf_8 _3241_ (.A(\products[14][1] ),
    .X(_2655_));
 sg13g2_buf_8 _3242_ (.A(\products[1][1] ),
    .X(_2656_));
 sg13g2_xnor2_1 _3243_ (.Y(_2657_),
    .A(_2655_),
    .B(_2656_));
 sg13g2_xnor2_1 _3244_ (.Y(_2658_),
    .A(\products[15][1] ),
    .B(_2657_));
 sg13g2_o21ai_1 _3245_ (.B1(_2658_),
    .Y(_2659_),
    .A1(_2653_),
    .A2(_2654_));
 sg13g2_buf_1 _3246_ (.A(_2659_),
    .X(_2660_));
 sg13g2_or3_1 _3247_ (.A(_2653_),
    .B(_2654_),
    .C(_2658_),
    .X(_2661_));
 sg13g2_buf_1 _3248_ (.A(_2661_),
    .X(_2662_));
 sg13g2_nand3_1 _3249_ (.B(_2660_),
    .C(_2662_),
    .A(_2648_),
    .Y(_2663_));
 sg13g2_a21o_1 _3250_ (.A2(_2662_),
    .A1(_2660_),
    .B1(_2648_),
    .X(_2664_));
 sg13g2_buf_2 _3251_ (.A(\prev_acc[1] ),
    .X(_2665_));
 sg13g2_xnor2_1 _3252_ (.Y(_2666_),
    .A(_2665_),
    .B(\products[10][1] ));
 sg13g2_xnor2_1 _3253_ (.Y(_2667_),
    .A(\products[0][1] ),
    .B(_2666_));
 sg13g2_nor2_1 _3254_ (.A(_2618_),
    .B(\products[10][0] ),
    .Y(_2668_));
 sg13g2_a21oi_1 _3255_ (.A1(_2618_),
    .A2(\products[10][0] ),
    .Y(_2669_),
    .B1(\products[0][0] ));
 sg13g2_nor2_1 _3256_ (.A(_2668_),
    .B(_2669_),
    .Y(_2670_));
 sg13g2_buf_1 _3257_ (.A(\products[11][1] ),
    .X(_2671_));
 sg13g2_buf_1 _3258_ (.A(\products[13][1] ),
    .X(_2672_));
 sg13g2_xnor2_1 _3259_ (.Y(_2673_),
    .A(_2671_),
    .B(_2672_));
 sg13g2_xnor2_1 _3260_ (.Y(_2674_),
    .A(\products[12][1] ),
    .B(_2673_));
 sg13g2_xor2_1 _3261_ (.B(_2674_),
    .A(_2670_),
    .X(_2675_));
 sg13g2_xnor2_1 _3262_ (.Y(_2676_),
    .A(_2667_),
    .B(_2675_));
 sg13g2_a21oi_1 _3263_ (.A1(_2663_),
    .A2(_2664_),
    .Y(_2677_),
    .B1(_2676_));
 sg13g2_xor2_1 _3264_ (.B(_2675_),
    .A(_2667_),
    .X(_2678_));
 sg13g2_and3_1 _3265_ (.X(_2679_),
    .A(_2648_),
    .B(_2660_),
    .C(_2662_));
 sg13g2_a21oi_1 _3266_ (.A1(_2660_),
    .A2(_2662_),
    .Y(_2680_),
    .B1(_2648_));
 sg13g2_nor3_1 _3267_ (.A(_2678_),
    .B(_2679_),
    .C(_2680_),
    .Y(_2681_));
 sg13g2_or2_1 _3268_ (.X(_2682_),
    .B(_2681_),
    .A(_2677_));
 sg13g2_nand2_1 _3269_ (.Y(_2683_),
    .A(_2615_),
    .B(_2621_));
 sg13g2_inv_1 _3270_ (.Y(_2684_),
    .A(_2683_));
 sg13g2_nand2_1 _3271_ (.Y(_2685_),
    .A(_2624_),
    .B(_2626_));
 sg13g2_xnor2_1 _3272_ (.Y(_2686_),
    .A(\products[2][1] ),
    .B(\products[4][1] ));
 sg13g2_xor2_1 _3273_ (.B(_2686_),
    .A(\products[3][1] ),
    .X(_2687_));
 sg13g2_nor2_1 _3274_ (.A(\products[2][0] ),
    .B(\products[4][0] ),
    .Y(_2688_));
 sg13g2_a21oi_1 _3275_ (.A1(\products[2][0] ),
    .A2(\products[4][0] ),
    .Y(_2689_),
    .B1(\products[3][0] ));
 sg13g2_nor2_2 _3276_ (.A(_2688_),
    .B(_2689_),
    .Y(_2690_));
 sg13g2_xnor2_1 _3277_ (.Y(_2691_),
    .A(\products[5][1] ),
    .B(\products[7][1] ));
 sg13g2_xnor2_1 _3278_ (.Y(_2692_),
    .A(\products[6][1] ),
    .B(_2691_));
 sg13g2_xnor2_1 _3279_ (.Y(_2693_),
    .A(_2690_),
    .B(_2692_));
 sg13g2_nand3_1 _3280_ (.B(_2687_),
    .C(_2693_),
    .A(_2685_),
    .Y(_2694_));
 sg13g2_xnor2_1 _3281_ (.Y(_2695_),
    .A(\products[3][1] ),
    .B(_2686_));
 sg13g2_nand3b_1 _3282_ (.B(_2695_),
    .C(_2685_),
    .Y(_2696_),
    .A_N(_2693_));
 sg13g2_nand3_1 _3283_ (.B(_2626_),
    .C(_2687_),
    .A(_2624_),
    .Y(_2697_));
 sg13g2_nand3_1 _3284_ (.B(_2626_),
    .C(_2695_),
    .A(_2624_),
    .Y(_2698_));
 sg13g2_mux2_1 _3285_ (.A0(_2697_),
    .A1(_2698_),
    .S(_2693_),
    .X(_2699_));
 sg13g2_and3_1 _3286_ (.X(_2700_),
    .A(_2694_),
    .B(_2696_),
    .C(_2699_));
 sg13g2_buf_1 _3287_ (.A(_2700_),
    .X(_2701_));
 sg13g2_xnor2_1 _3288_ (.Y(_2702_),
    .A(_2684_),
    .B(_2701_));
 sg13g2_xor2_1 _3289_ (.B(_2702_),
    .A(_2682_),
    .X(_2703_));
 sg13g2_buf_2 _3290_ (.A(_2703_),
    .X(_2704_));
 sg13g2_nand2_1 _3291_ (.Y(_2705_),
    .A(\products[8][0] ),
    .B(\products[9][0] ));
 sg13g2_nor2_1 _3292_ (.A(\products[5][0] ),
    .B(\products[7][0] ),
    .Y(_2706_));
 sg13g2_a21oi_1 _3293_ (.A1(\products[5][0] ),
    .A2(\products[7][0] ),
    .Y(_2707_),
    .B1(\products[6][0] ));
 sg13g2_nor2_1 _3294_ (.A(_2706_),
    .B(_2707_),
    .Y(_2708_));
 sg13g2_xnor2_1 _3295_ (.Y(_2709_),
    .A(\products[8][1] ),
    .B(\products[9][1] ));
 sg13g2_xnor2_1 _3296_ (.Y(_2710_),
    .A(_2708_),
    .B(_2709_));
 sg13g2_xor2_1 _3297_ (.B(_2710_),
    .A(_2705_),
    .X(_2711_));
 sg13g2_nand2_2 _3298_ (.Y(_2712_),
    .A(_2622_),
    .B(_2627_));
 sg13g2_nand2_1 _3299_ (.Y(_2713_),
    .A(_2613_),
    .B(_2628_));
 sg13g2_and2_1 _3300_ (.A(_2712_),
    .B(_2713_),
    .X(_2714_));
 sg13g2_buf_1 _3301_ (.A(_2714_),
    .X(_2715_));
 sg13g2_xnor2_1 _3302_ (.Y(_2716_),
    .A(_2711_),
    .B(_2715_));
 sg13g2_xnor2_1 _3303_ (.Y(_2717_),
    .A(_2704_),
    .B(_2716_));
 sg13g2_nand2_1 _3304_ (.Y(_2718_),
    .A(net4),
    .B(_2647_));
 sg13g2_o21ai_1 _3305_ (.B1(_2718_),
    .Y(_2719_),
    .A1(_2647_),
    .A2(_2717_));
 sg13g2_buf_1 _3306_ (.A(_2719_),
    .X(_2720_));
 sg13g2_buf_1 _3307_ (.A(net45),
    .X(_2721_));
 sg13g2_buf_1 _3308_ (.A(\mem[0][1] ),
    .X(_2722_));
 sg13g2_mux2_1 _3309_ (.A0(net44),
    .A1(net174),
    .S(_2645_),
    .X(_0002_));
 sg13g2_xnor2_1 _3310_ (.Y(_2723_),
    .A(\products[5][2] ),
    .B(\products[7][2] ));
 sg13g2_xnor2_1 _3311_ (.Y(_2724_),
    .A(\products[6][2] ),
    .B(_2723_));
 sg13g2_nor2_1 _3312_ (.A(\products[2][1] ),
    .B(\products[4][1] ),
    .Y(_2725_));
 sg13g2_a21oi_1 _3313_ (.A1(\products[2][1] ),
    .A2(\products[4][1] ),
    .Y(_2726_),
    .B1(\products[3][1] ));
 sg13g2_nor2_1 _3314_ (.A(_2725_),
    .B(_2726_),
    .Y(_2727_));
 sg13g2_xnor2_1 _3315_ (.Y(_2728_),
    .A(\products[2][2] ),
    .B(\products[4][2] ));
 sg13g2_xnor2_1 _3316_ (.Y(_2729_),
    .A(\products[3][2] ),
    .B(_2728_));
 sg13g2_xor2_1 _3317_ (.B(_2729_),
    .A(_2727_),
    .X(_2730_));
 sg13g2_xnor2_1 _3318_ (.Y(_2731_),
    .A(_2724_),
    .B(_2730_));
 sg13g2_nand2_1 _3319_ (.Y(_2732_),
    .A(_2651_),
    .B(_2652_));
 sg13g2_nand2_1 _3320_ (.Y(_2733_),
    .A(_2649_),
    .B(_2650_));
 sg13g2_o21ai_1 _3321_ (.B1(_2733_),
    .Y(_2734_),
    .A1(_2732_),
    .A2(_2658_));
 sg13g2_nand2_1 _3322_ (.Y(_2735_),
    .A(_2732_),
    .B(_2658_));
 sg13g2_a21o_1 _3323_ (.A2(_2695_),
    .A1(_2692_),
    .B1(_2690_),
    .X(_2736_));
 sg13g2_nand2b_1 _3324_ (.Y(_2737_),
    .B(_2687_),
    .A_N(_2692_));
 sg13g2_nand4_1 _3325_ (.B(_2735_),
    .C(_2736_),
    .A(_2734_),
    .Y(_2738_),
    .D(_2737_));
 sg13g2_nand2_1 _3326_ (.Y(_2739_),
    .A(_2690_),
    .B(_2692_));
 sg13g2_a21o_1 _3327_ (.A2(_2658_),
    .A1(_2733_),
    .B1(_2732_),
    .X(_2740_));
 sg13g2_or2_1 _3328_ (.X(_2741_),
    .B(_2658_),
    .A(_2733_));
 sg13g2_o21ai_1 _3329_ (.B1(_2695_),
    .Y(_2742_),
    .A1(_2690_),
    .A2(_2692_));
 sg13g2_nand4_1 _3330_ (.B(_2740_),
    .C(_2741_),
    .A(_2739_),
    .Y(_2743_),
    .D(_2742_));
 sg13g2_nand3_1 _3331_ (.B(_2738_),
    .C(_2743_),
    .A(_2731_),
    .Y(_2744_));
 sg13g2_buf_2 _3332_ (.A(_2744_),
    .X(_2745_));
 sg13g2_a21o_1 _3333_ (.A2(_2743_),
    .A1(_2738_),
    .B1(_2731_),
    .X(_2746_));
 sg13g2_buf_2 _3334_ (.A(_2746_),
    .X(_2747_));
 sg13g2_a21oi_2 _3335_ (.B1(_2680_),
    .Y(_2748_),
    .A2(_2663_),
    .A1(_2678_));
 sg13g2_a21oi_1 _3336_ (.A1(_2745_),
    .A2(_2747_),
    .Y(_2749_),
    .B1(_2748_));
 sg13g2_and3_1 _3337_ (.X(_2750_),
    .A(_2748_),
    .B(_2745_),
    .C(_2747_));
 sg13g2_xnor2_1 _3338_ (.Y(_2751_),
    .A(\products[11][2] ),
    .B(\products[13][2] ));
 sg13g2_xnor2_1 _3339_ (.Y(_2752_),
    .A(\products[12][2] ),
    .B(_2751_));
 sg13g2_nor2_1 _3340_ (.A(_2665_),
    .B(\products[10][1] ),
    .Y(_2753_));
 sg13g2_a21oi_1 _3341_ (.A1(_2665_),
    .A2(\products[10][1] ),
    .Y(_2754_),
    .B1(\products[0][1] ));
 sg13g2_nor2_1 _3342_ (.A(_2753_),
    .B(_2754_),
    .Y(_2755_));
 sg13g2_buf_2 _3343_ (.A(\prev_acc[2] ),
    .X(_2756_));
 sg13g2_xnor2_1 _3344_ (.Y(_2757_),
    .A(_2756_),
    .B(\products[10][2] ));
 sg13g2_xnor2_1 _3345_ (.Y(_2758_),
    .A(\products[0][2] ),
    .B(_2757_));
 sg13g2_xnor2_1 _3346_ (.Y(_2759_),
    .A(_2755_),
    .B(_2758_));
 sg13g2_xnor2_1 _3347_ (.Y(_2760_),
    .A(_2752_),
    .B(_2759_));
 sg13g2_or2_1 _3348_ (.X(_2761_),
    .B(_2667_),
    .A(_2670_));
 sg13g2_buf_1 _3349_ (.A(_2761_),
    .X(_2762_));
 sg13g2_a21o_1 _3350_ (.A2(_2667_),
    .A1(_2670_),
    .B1(_2674_),
    .X(_2763_));
 sg13g2_buf_8 _3351_ (.A(\products[14][2] ),
    .X(_2764_));
 sg13g2_buf_8 _3352_ (.A(\products[1][2] ),
    .X(_2765_));
 sg13g2_xnor2_1 _3353_ (.Y(_2766_),
    .A(_2764_),
    .B(_2765_));
 sg13g2_xnor2_1 _3354_ (.Y(_2767_),
    .A(\products[15][2] ),
    .B(_2766_));
 sg13g2_or2_1 _3355_ (.X(_2768_),
    .B(_2672_),
    .A(_2671_));
 sg13g2_a21o_1 _3356_ (.A2(_2672_),
    .A1(_2671_),
    .B1(\products[12][1] ),
    .X(_2769_));
 sg13g2_nand2_1 _3357_ (.Y(_2770_),
    .A(_2655_),
    .B(_2656_));
 sg13g2_o21ai_1 _3358_ (.B1(\products[15][1] ),
    .Y(_2771_),
    .A1(_2655_),
    .A2(_2656_));
 sg13g2_nand4_1 _3359_ (.B(_2769_),
    .C(_2770_),
    .A(_2768_),
    .Y(_2772_),
    .D(_2771_));
 sg13g2_nand2_1 _3360_ (.Y(_2773_),
    .A(_2671_),
    .B(_2672_));
 sg13g2_o21ai_1 _3361_ (.B1(\products[12][1] ),
    .Y(_2774_),
    .A1(_2671_),
    .A2(_2672_));
 sg13g2_or2_1 _3362_ (.X(_2775_),
    .B(_2656_),
    .A(_2655_));
 sg13g2_a21o_1 _3363_ (.A2(_2656_),
    .A1(_2655_),
    .B1(\products[15][1] ),
    .X(_2776_));
 sg13g2_nand4_1 _3364_ (.B(_2774_),
    .C(_2775_),
    .A(_2773_),
    .Y(_2777_),
    .D(_2776_));
 sg13g2_nand3_1 _3365_ (.B(_2772_),
    .C(_2777_),
    .A(_2767_),
    .Y(_2778_));
 sg13g2_a21o_1 _3366_ (.A2(_2777_),
    .A1(_2772_),
    .B1(_2767_),
    .X(_2779_));
 sg13g2_a22oi_1 _3367_ (.Y(_2780_),
    .B1(_2778_),
    .B2(_2779_),
    .A2(_2763_),
    .A1(_2762_));
 sg13g2_and4_1 _3368_ (.A(_2762_),
    .B(_2763_),
    .C(_2778_),
    .D(_2779_),
    .X(_2781_));
 sg13g2_or3_1 _3369_ (.A(_2760_),
    .B(_2780_),
    .C(_2781_),
    .X(_2782_));
 sg13g2_buf_2 _3370_ (.A(_2782_),
    .X(_2783_));
 sg13g2_o21ai_1 _3371_ (.B1(_2760_),
    .Y(_2784_),
    .A1(_2780_),
    .A2(_2781_));
 sg13g2_buf_2 _3372_ (.A(_2784_),
    .X(_2785_));
 sg13g2_nand2_2 _3373_ (.Y(_2786_),
    .A(_2783_),
    .B(_2785_));
 sg13g2_o21ai_1 _3374_ (.B1(_2786_),
    .Y(_2787_),
    .A1(_2749_),
    .A2(_2750_));
 sg13g2_and2_1 _3375_ (.A(_2783_),
    .B(_2785_),
    .X(_2788_));
 sg13g2_buf_2 _3376_ (.A(_2788_),
    .X(_2789_));
 sg13g2_a21o_1 _3377_ (.A2(_2747_),
    .A1(_2745_),
    .B1(_2748_),
    .X(_2790_));
 sg13g2_nand3_1 _3378_ (.B(_2745_),
    .C(_2747_),
    .A(_2748_),
    .Y(_2791_));
 sg13g2_nand3_1 _3379_ (.B(_2790_),
    .C(_2791_),
    .A(_2789_),
    .Y(_2792_));
 sg13g2_nor2_1 _3380_ (.A(\products[5][1] ),
    .B(\products[7][1] ),
    .Y(_2793_));
 sg13g2_a21oi_1 _3381_ (.A1(\products[5][1] ),
    .A2(\products[7][1] ),
    .Y(_2794_),
    .B1(\products[6][1] ));
 sg13g2_nor2_1 _3382_ (.A(_2793_),
    .B(_2794_),
    .Y(_0395_));
 sg13g2_xnor2_1 _3383_ (.Y(_0396_),
    .A(\products[8][2] ),
    .B(\products[9][2] ));
 sg13g2_xnor2_1 _3384_ (.Y(_0397_),
    .A(_0395_),
    .B(_0396_));
 sg13g2_or2_1 _3385_ (.X(_0398_),
    .B(\products[9][1] ),
    .A(\products[8][1] ));
 sg13g2_and2_1 _3386_ (.A(\products[8][1] ),
    .B(\products[9][1] ),
    .X(_0399_));
 sg13g2_a21oi_2 _3387_ (.B1(_0399_),
    .Y(_0400_),
    .A2(_0398_),
    .A1(_2708_));
 sg13g2_xor2_1 _3388_ (.B(_0400_),
    .A(_0397_),
    .X(_0401_));
 sg13g2_xnor2_1 _3389_ (.Y(_0402_),
    .A(_2699_),
    .B(_0401_));
 sg13g2_inv_1 _3390_ (.Y(_0403_),
    .A(_0402_));
 sg13g2_o21ai_1 _3391_ (.B1(_2701_),
    .Y(_0404_),
    .A1(_2677_),
    .A2(_2681_));
 sg13g2_buf_1 _3392_ (.A(_0404_),
    .X(_0405_));
 sg13g2_nor2_1 _3393_ (.A(_2683_),
    .B(_2676_),
    .Y(_0406_));
 sg13g2_nand2_1 _3394_ (.Y(_0407_),
    .A(_2663_),
    .B(_2664_));
 sg13g2_nor4_1 _3395_ (.A(_2683_),
    .B(_2678_),
    .C(_2679_),
    .D(_2680_),
    .Y(_0408_));
 sg13g2_a221oi_1 _3396_ (.B2(_0407_),
    .C1(_0408_),
    .B1(_0406_),
    .A1(_2684_),
    .Y(_0409_),
    .A2(_2701_));
 sg13g2_buf_2 _3397_ (.A(_0409_),
    .X(_0410_));
 sg13g2_nand3_1 _3398_ (.B(_0405_),
    .C(_0410_),
    .A(_0403_),
    .Y(_0411_));
 sg13g2_a21o_1 _3399_ (.A2(_0410_),
    .A1(_0405_),
    .B1(_0403_),
    .X(_0412_));
 sg13g2_and4_1 _3400_ (.A(_2787_),
    .B(_2792_),
    .C(_0411_),
    .D(_0412_),
    .X(_0413_));
 sg13g2_buf_1 _3401_ (.A(_0413_),
    .X(_0414_));
 sg13g2_a22oi_1 _3402_ (.Y(_0415_),
    .B1(_0411_),
    .B2(_0412_),
    .A2(_2792_),
    .A1(_2787_));
 sg13g2_nor2_2 _3403_ (.A(_0414_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_nor2b_2 _3404_ (.A(_2710_),
    .B_N(_2705_),
    .Y(_0417_));
 sg13g2_nand2b_1 _3405_ (.Y(_0418_),
    .B(_2710_),
    .A_N(_2705_));
 sg13g2_a21o_1 _3406_ (.A2(_0418_),
    .A1(_2715_),
    .B1(_0417_),
    .X(_0419_));
 sg13g2_nor3_1 _3407_ (.A(_2704_),
    .B(_2715_),
    .C(_0418_),
    .Y(_0420_));
 sg13g2_a221oi_1 _3408_ (.B2(_2704_),
    .C1(_0420_),
    .B1(_0419_),
    .A1(_2715_),
    .Y(_0421_),
    .A2(_0417_));
 sg13g2_xnor2_1 _3409_ (.Y(_0422_),
    .A(_0416_),
    .B(_0421_));
 sg13g2_nand2_1 _3410_ (.Y(_0423_),
    .A(net5),
    .B(_2647_));
 sg13g2_o21ai_1 _3411_ (.B1(_0423_),
    .Y(_0424_),
    .A1(_2647_),
    .A2(_0422_));
 sg13g2_buf_1 _3412_ (.A(_0424_),
    .X(_0425_));
 sg13g2_buf_1 _3413_ (.A(net38),
    .X(_0426_));
 sg13g2_buf_1 _3414_ (.A(\mem[0][2] ),
    .X(_0427_));
 sg13g2_mux2_1 _3415_ (.A0(net37),
    .A1(net173),
    .S(_2645_),
    .X(_0003_));
 sg13g2_nor2_1 _3416_ (.A(_2712_),
    .B(_2704_),
    .Y(_0428_));
 sg13g2_and2_1 _3417_ (.A(_2712_),
    .B(_2704_),
    .X(_0429_));
 sg13g2_mux2_1 _3418_ (.A0(_0428_),
    .A1(_0429_),
    .S(_0416_),
    .X(_0430_));
 sg13g2_nor2_1 _3419_ (.A(_2713_),
    .B(_2711_),
    .Y(_0431_));
 sg13g2_xnor2_1 _3420_ (.Y(_0432_),
    .A(_2712_),
    .B(_2704_));
 sg13g2_nor2_1 _3421_ (.A(_2713_),
    .B(_0432_),
    .Y(_0433_));
 sg13g2_nor2b_1 _3422_ (.A(_2705_),
    .B_N(_2710_),
    .Y(_0434_));
 sg13g2_mux2_1 _3423_ (.A0(_0434_),
    .A1(_0417_),
    .S(_0416_),
    .X(_0435_));
 sg13g2_a22oi_1 _3424_ (.Y(_0436_),
    .B1(_0433_),
    .B2(_0435_),
    .A2(_0431_),
    .A1(_0430_));
 sg13g2_o21ai_1 _3425_ (.B1(_0418_),
    .Y(_0437_),
    .A1(_0414_),
    .A2(_0415_));
 sg13g2_nor2_1 _3426_ (.A(_2712_),
    .B(_0417_),
    .Y(_0438_));
 sg13g2_xnor2_1 _3427_ (.Y(_0439_),
    .A(_2682_),
    .B(_2702_));
 sg13g2_inv_1 _3428_ (.Y(_0440_),
    .A(_0417_));
 sg13g2_a21oi_1 _3429_ (.A1(_0439_),
    .A2(_0440_),
    .Y(_0441_),
    .B1(_0434_));
 sg13g2_nor3_1 _3430_ (.A(_0414_),
    .B(_0415_),
    .C(_0441_),
    .Y(_0442_));
 sg13g2_a221oi_1 _3431_ (.B2(_0416_),
    .C1(_0442_),
    .B1(_0438_),
    .A1(_0428_),
    .Y(_0443_),
    .A2(_0437_));
 sg13g2_nand2_1 _3432_ (.Y(_0444_),
    .A(_2778_),
    .B(_2779_));
 sg13g2_a22oi_1 _3433_ (.Y(_0445_),
    .B1(_2760_),
    .B2(_0444_),
    .A2(_2763_),
    .A1(_2762_));
 sg13g2_nor2_1 _3434_ (.A(_2760_),
    .B(_0444_),
    .Y(_0446_));
 sg13g2_nor2_1 _3435_ (.A(_0445_),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_buf_2 _3436_ (.A(\products[14][3] ),
    .X(_0448_));
 sg13g2_buf_2 _3437_ (.A(\products[1][3] ),
    .X(_0449_));
 sg13g2_xnor2_1 _3438_ (.Y(_0450_),
    .A(_0448_),
    .B(_0449_));
 sg13g2_xnor2_1 _3439_ (.Y(_0451_),
    .A(\products[15][3] ),
    .B(_0450_));
 sg13g2_nand2_1 _3440_ (.Y(_0452_),
    .A(\products[11][2] ),
    .B(\products[13][2] ));
 sg13g2_o21ai_1 _3441_ (.B1(\products[12][2] ),
    .Y(_0453_),
    .A1(\products[11][2] ),
    .A2(\products[13][2] ));
 sg13g2_buf_1 _3442_ (.A(_0453_),
    .X(_0454_));
 sg13g2_or2_1 _3443_ (.X(_0455_),
    .B(_2765_),
    .A(_2764_));
 sg13g2_a21o_1 _3444_ (.A2(_2765_),
    .A1(_2764_),
    .B1(\products[15][2] ),
    .X(_0456_));
 sg13g2_a22oi_1 _3445_ (.Y(_0457_),
    .B1(_0455_),
    .B2(_0456_),
    .A2(_0454_),
    .A1(_0452_));
 sg13g2_and4_1 _3446_ (.A(_0452_),
    .B(_0454_),
    .C(_0455_),
    .D(_0456_),
    .X(_0458_));
 sg13g2_or3_1 _3447_ (.A(_0451_),
    .B(_0457_),
    .C(_0458_),
    .X(_0459_));
 sg13g2_o21ai_1 _3448_ (.B1(_0451_),
    .Y(_0460_),
    .A1(_0457_),
    .A2(_0458_));
 sg13g2_or2_1 _3449_ (.X(_0461_),
    .B(_2758_),
    .A(_2752_));
 sg13g2_buf_1 _3450_ (.A(_0461_),
    .X(_0462_));
 sg13g2_a21o_1 _3451_ (.A2(_2758_),
    .A1(_2752_),
    .B1(_2755_),
    .X(_0463_));
 sg13g2_and4_1 _3452_ (.A(_0459_),
    .B(_0460_),
    .C(_0462_),
    .D(_0463_),
    .X(_0464_));
 sg13g2_a22oi_1 _3453_ (.Y(_0465_),
    .B1(_0462_),
    .B2(_0463_),
    .A2(_0460_),
    .A1(_0459_));
 sg13g2_buf_2 _3454_ (.A(\products[11][3] ),
    .X(_0466_));
 sg13g2_buf_2 _3455_ (.A(\products[13][3] ),
    .X(_0467_));
 sg13g2_xnor2_1 _3456_ (.Y(_0468_),
    .A(_0466_),
    .B(_0467_));
 sg13g2_xnor2_1 _3457_ (.Y(_0469_),
    .A(\products[12][3] ),
    .B(_0468_));
 sg13g2_nor2_1 _3458_ (.A(_2756_),
    .B(\products[10][2] ),
    .Y(_0470_));
 sg13g2_a21oi_1 _3459_ (.A1(_2756_),
    .A2(\products[10][2] ),
    .Y(_0471_),
    .B1(\products[0][2] ));
 sg13g2_nor2_1 _3460_ (.A(_0470_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_buf_1 _3461_ (.A(\prev_acc[3] ),
    .X(_0473_));
 sg13g2_xnor2_1 _3462_ (.Y(_0474_),
    .A(_0473_),
    .B(\products[10][3] ));
 sg13g2_xnor2_1 _3463_ (.Y(_0475_),
    .A(\products[0][3] ),
    .B(_0474_));
 sg13g2_xor2_1 _3464_ (.B(_0475_),
    .A(_0472_),
    .X(_0476_));
 sg13g2_xor2_1 _3465_ (.B(_0476_),
    .A(_0469_),
    .X(_0477_));
 sg13g2_o21ai_1 _3466_ (.B1(_0477_),
    .Y(_0478_),
    .A1(_0464_),
    .A2(_0465_));
 sg13g2_xnor2_1 _3467_ (.Y(_0479_),
    .A(_0469_),
    .B(_0476_));
 sg13g2_nand4_1 _3468_ (.B(_0460_),
    .C(_0462_),
    .A(_0459_),
    .Y(_0480_),
    .D(_0463_));
 sg13g2_nand3b_1 _3469_ (.B(_0479_),
    .C(_0480_),
    .Y(_0481_),
    .A_N(_0465_));
 sg13g2_a22oi_1 _3470_ (.Y(_0482_),
    .B1(_2770_),
    .B2(_2771_),
    .A2(_2774_),
    .A1(_2773_));
 sg13g2_nand4_1 _3471_ (.B(_2774_),
    .C(_2770_),
    .A(_2773_),
    .Y(_0483_),
    .D(_2771_));
 sg13g2_o21ai_1 _3472_ (.B1(_0483_),
    .Y(_0484_),
    .A1(_2767_),
    .A2(_0482_));
 sg13g2_nand2_1 _3473_ (.Y(_0485_),
    .A(_2724_),
    .B(_2729_));
 sg13g2_o21ai_1 _3474_ (.B1(_2727_),
    .Y(_0486_),
    .A1(_2724_),
    .A2(_2729_));
 sg13g2_and3_1 _3475_ (.X(_0487_),
    .A(_0484_),
    .B(_0485_),
    .C(_0486_));
 sg13g2_a21oi_1 _3476_ (.A1(_0485_),
    .A2(_0486_),
    .Y(_0488_),
    .B1(_0484_));
 sg13g2_xnor2_1 _3477_ (.Y(_0489_),
    .A(\products[2][3] ),
    .B(\products[4][3] ));
 sg13g2_xnor2_1 _3478_ (.Y(_0490_),
    .A(\products[3][3] ),
    .B(_0489_));
 sg13g2_a21oi_1 _3479_ (.A1(\products[2][2] ),
    .A2(\products[4][2] ),
    .Y(_0491_),
    .B1(\products[3][2] ));
 sg13g2_nor2_1 _3480_ (.A(\products[2][2] ),
    .B(\products[4][2] ),
    .Y(_0492_));
 sg13g2_nor2_1 _3481_ (.A(_0491_),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_xnor2_1 _3482_ (.Y(_0494_),
    .A(\products[5][3] ),
    .B(\products[7][3] ));
 sg13g2_xnor2_1 _3483_ (.Y(_0495_),
    .A(\products[6][3] ),
    .B(_0494_));
 sg13g2_xnor2_1 _3484_ (.Y(_0496_),
    .A(_0493_),
    .B(_0495_));
 sg13g2_xnor2_1 _3485_ (.Y(_0497_),
    .A(_0490_),
    .B(_0496_));
 sg13g2_o21ai_1 _3486_ (.B1(_0497_),
    .Y(_0498_),
    .A1(_0487_),
    .A2(_0488_));
 sg13g2_or3_1 _3487_ (.A(_0497_),
    .B(_0487_),
    .C(_0488_),
    .X(_0499_));
 sg13g2_buf_1 _3488_ (.A(_0499_),
    .X(_0500_));
 sg13g2_a22oi_1 _3489_ (.Y(_0501_),
    .B1(_0498_),
    .B2(_0500_),
    .A2(_0481_),
    .A1(_0478_));
 sg13g2_and4_1 _3490_ (.A(_0478_),
    .B(_0481_),
    .C(_0498_),
    .D(_0500_),
    .X(_0502_));
 sg13g2_or3_1 _3491_ (.A(_0447_),
    .B(_0501_),
    .C(_0502_),
    .X(_0503_));
 sg13g2_o21ai_1 _3492_ (.B1(_0447_),
    .Y(_0504_),
    .A1(_0501_),
    .A2(_0502_));
 sg13g2_and2_1 _3493_ (.A(_0503_),
    .B(_0504_),
    .X(_0505_));
 sg13g2_nand4_1 _3494_ (.B(_2785_),
    .C(_2745_),
    .A(_2783_),
    .Y(_0506_),
    .D(_2747_));
 sg13g2_a22oi_1 _3495_ (.Y(_0507_),
    .B1(_2745_),
    .B2(_2747_),
    .A2(_2785_),
    .A1(_2783_));
 sg13g2_a21oi_1 _3496_ (.A1(_2748_),
    .A2(_0506_),
    .Y(_0508_),
    .B1(_0507_));
 sg13g2_xor2_1 _3497_ (.B(_2730_),
    .A(_2724_),
    .X(_0509_));
 sg13g2_nand4_1 _3498_ (.B(_2734_),
    .C(_2735_),
    .A(_2739_),
    .Y(_0510_),
    .D(_2742_));
 sg13g2_a22oi_1 _3499_ (.Y(_0511_),
    .B1(_2742_),
    .B2(_2739_),
    .A2(_2735_),
    .A1(_2734_));
 sg13g2_a21oi_1 _3500_ (.A1(_0509_),
    .A2(_0510_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_nor2_1 _3501_ (.A(\products[5][2] ),
    .B(\products[7][2] ),
    .Y(_0513_));
 sg13g2_a21oi_1 _3502_ (.A1(\products[5][2] ),
    .A2(\products[7][2] ),
    .Y(_0514_),
    .B1(\products[6][2] ));
 sg13g2_nor2_1 _3503_ (.A(_0513_),
    .B(_0514_),
    .Y(_0515_));
 sg13g2_xnor2_1 _3504_ (.Y(_0516_),
    .A(\products[8][3] ),
    .B(\products[9][3] ));
 sg13g2_xnor2_1 _3505_ (.Y(_0517_),
    .A(_0515_),
    .B(_0516_));
 sg13g2_inv_1 _3506_ (.Y(_0518_),
    .A(_0517_));
 sg13g2_a21o_1 _3507_ (.A2(\products[9][2] ),
    .A1(\products[8][2] ),
    .B1(_0395_),
    .X(_0519_));
 sg13g2_o21ai_1 _3508_ (.B1(_0519_),
    .Y(_0520_),
    .A1(\products[8][2] ),
    .A2(\products[9][2] ));
 sg13g2_xnor2_1 _3509_ (.Y(_0521_),
    .A(_0518_),
    .B(_0520_));
 sg13g2_xnor2_1 _3510_ (.Y(_0522_),
    .A(_0512_),
    .B(_0521_));
 sg13g2_xnor2_1 _3511_ (.Y(_0523_),
    .A(_0508_),
    .B(_0522_));
 sg13g2_xnor2_1 _3512_ (.Y(_0524_),
    .A(_0505_),
    .B(_0523_));
 sg13g2_nand2_1 _3513_ (.Y(_0525_),
    .A(_2790_),
    .B(_2791_));
 sg13g2_and2_1 _3514_ (.A(_0405_),
    .B(_0410_),
    .X(_0526_));
 sg13g2_nor2b_1 _3515_ (.A(_0397_),
    .B_N(_0400_),
    .Y(_0527_));
 sg13g2_nand2b_1 _3516_ (.Y(_0528_),
    .B(_0397_),
    .A_N(_0400_));
 sg13g2_o21ai_1 _3517_ (.B1(_0528_),
    .Y(_0529_),
    .A1(_2699_),
    .A2(_0527_));
 sg13g2_buf_2 _3518_ (.A(_0529_),
    .X(_0530_));
 sg13g2_nand4_1 _3519_ (.B(_0525_),
    .C(_0526_),
    .A(_2789_),
    .Y(_0531_),
    .D(_0530_));
 sg13g2_nor2_1 _3520_ (.A(_2749_),
    .B(_2750_),
    .Y(_0532_));
 sg13g2_nand4_1 _3521_ (.B(_0532_),
    .C(_0526_),
    .A(_2786_),
    .Y(_0533_),
    .D(_0530_));
 sg13g2_nand2_1 _3522_ (.Y(_0534_),
    .A(_0402_),
    .B(_0530_));
 sg13g2_inv_1 _3523_ (.Y(_0535_),
    .A(_0534_));
 sg13g2_nor2_1 _3524_ (.A(_2786_),
    .B(_0534_),
    .Y(_0536_));
 sg13g2_a22oi_1 _3525_ (.Y(_0537_),
    .B1(_0536_),
    .B2(_0525_),
    .A2(_0535_),
    .A1(_0526_));
 sg13g2_nor2_1 _3526_ (.A(_2789_),
    .B(_0534_),
    .Y(_0538_));
 sg13g2_nor2_1 _3527_ (.A(_0402_),
    .B(_0530_),
    .Y(_0539_));
 sg13g2_nand2_2 _3528_ (.Y(_0540_),
    .A(_0405_),
    .B(_0410_));
 sg13g2_a22oi_1 _3529_ (.Y(_0541_),
    .B1(_0539_),
    .B2(_0540_),
    .A2(_0538_),
    .A1(_0532_));
 sg13g2_nand4_1 _3530_ (.B(_0533_),
    .C(_0537_),
    .A(_0531_),
    .Y(_0542_),
    .D(_0541_));
 sg13g2_inv_1 _3531_ (.Y(_0543_),
    .A(_0530_));
 sg13g2_nand4_1 _3532_ (.B(_0525_),
    .C(_0540_),
    .A(_2786_),
    .Y(_0544_),
    .D(_0543_));
 sg13g2_nand4_1 _3533_ (.B(_0532_),
    .C(_0540_),
    .A(_2789_),
    .Y(_0545_),
    .D(_0543_));
 sg13g2_nand3_1 _3534_ (.B(_0525_),
    .C(_0539_),
    .A(_2786_),
    .Y(_0546_));
 sg13g2_nand3_1 _3535_ (.B(_0532_),
    .C(_0539_),
    .A(_2789_),
    .Y(_0547_));
 sg13g2_nand4_1 _3536_ (.B(_0545_),
    .C(_0546_),
    .A(_0544_),
    .Y(_0548_),
    .D(_0547_));
 sg13g2_or3_1 _3537_ (.A(_0524_),
    .B(_0542_),
    .C(_0548_),
    .X(_0549_));
 sg13g2_o21ai_1 _3538_ (.B1(_0524_),
    .Y(_0550_),
    .A1(_0542_),
    .A2(_0548_));
 sg13g2_and2_1 _3539_ (.A(_0549_),
    .B(_0550_),
    .X(_0551_));
 sg13g2_xor2_1 _3540_ (.B(_0551_),
    .A(_0443_),
    .X(_0552_));
 sg13g2_xor2_1 _3541_ (.B(_0552_),
    .A(_0436_),
    .X(_0553_));
 sg13g2_mux2_1 _3542_ (.A0(net6),
    .A1(_0553_),
    .S(net58),
    .X(_0554_));
 sg13g2_buf_8 _3543_ (.A(_0554_),
    .X(_0555_));
 sg13g2_buf_8 _3544_ (.A(net31),
    .X(_0556_));
 sg13g2_buf_1 _3545_ (.A(\mem[0][3] ),
    .X(_0557_));
 sg13g2_buf_1 _3546_ (.A(_0557_),
    .X(_0558_));
 sg13g2_mux2_1 _3547_ (.A0(net30),
    .A1(net81),
    .S(_2645_),
    .X(_0004_));
 sg13g2_buf_1 _3548_ (.A(\mem[10][0] ),
    .X(_0559_));
 sg13g2_inv_1 _3549_ (.Y(_0560_),
    .A(_2636_));
 sg13g2_nor4_1 _3550_ (.A(_2635_),
    .B(_0560_),
    .C(_2637_),
    .D(_2611_),
    .Y(_0561_));
 sg13g2_buf_4 _3551_ (.X(_0562_),
    .A(_0561_));
 sg13g2_buf_1 _3552_ (.A(_2640_),
    .X(_0563_));
 sg13g2_nand2b_1 _3553_ (.Y(_0564_),
    .B(net171),
    .A_N(_2641_));
 sg13g2_nor3_1 _3554_ (.A(_2642_),
    .B(net58),
    .C(_0564_),
    .Y(_0565_));
 sg13g2_buf_4 _3555_ (.X(_0566_),
    .A(_0565_));
 sg13g2_nand2_2 _3556_ (.Y(_0567_),
    .A(_0562_),
    .B(_0566_));
 sg13g2_mux2_1 _3557_ (.A0(net51),
    .A1(net172),
    .S(_0567_),
    .X(_0005_));
 sg13g2_buf_1 _3558_ (.A(\mem[10][1] ),
    .X(_0568_));
 sg13g2_mux2_1 _3559_ (.A0(net44),
    .A1(_0568_),
    .S(_0567_),
    .X(_0006_));
 sg13g2_buf_1 _3560_ (.A(\mem[10][2] ),
    .X(_0569_));
 sg13g2_mux2_1 _3561_ (.A0(net37),
    .A1(net170),
    .S(_0567_),
    .X(_0007_));
 sg13g2_buf_2 _3562_ (.A(\mem[10][3] ),
    .X(_0570_));
 sg13g2_mux2_1 _3563_ (.A0(net30),
    .A1(_0570_),
    .S(_0567_),
    .X(_0008_));
 sg13g2_buf_1 _3564_ (.A(\mem[11][0] ),
    .X(_0571_));
 sg13g2_inv_1 _3565_ (.Y(_0572_),
    .A(_0571_));
 sg13g2_inv_1 _3566_ (.Y(_0573_),
    .A(_2635_));
 sg13g2_buf_1 _3567_ (.A(_2637_),
    .X(_0574_));
 sg13g2_nor4_1 _3568_ (.A(_0573_),
    .B(_0560_),
    .C(_0574_),
    .D(net58),
    .Y(_0575_));
 sg13g2_buf_4 _3569_ (.X(_0576_),
    .A(_0575_));
 sg13g2_nand2_2 _3570_ (.Y(_0577_),
    .A(_0566_),
    .B(_0576_));
 sg13g2_nor2_1 _3571_ (.A(net52),
    .B(_0577_),
    .Y(_0578_));
 sg13g2_a21oi_1 _3572_ (.A1(_0572_),
    .A2(_0577_),
    .Y(_0009_),
    .B1(_0578_));
 sg13g2_buf_1 _3573_ (.A(\mem[11][1] ),
    .X(_0579_));
 sg13g2_buf_1 _3574_ (.A(_0579_),
    .X(_0580_));
 sg13g2_mux2_1 _3575_ (.A0(net44),
    .A1(net80),
    .S(_0577_),
    .X(_0010_));
 sg13g2_buf_1 _3576_ (.A(\mem[11][2] ),
    .X(_0581_));
 sg13g2_buf_1 _3577_ (.A(_0581_),
    .X(_0582_));
 sg13g2_buf_1 _3578_ (.A(net79),
    .X(_0583_));
 sg13g2_mux2_1 _3579_ (.A0(net37),
    .A1(net63),
    .S(_0577_),
    .X(_0011_));
 sg13g2_buf_1 _3580_ (.A(\mem[11][3] ),
    .X(_0584_));
 sg13g2_mux2_1 _3581_ (.A0(net30),
    .A1(net168),
    .S(_0577_),
    .X(_0012_));
 sg13g2_buf_1 _3582_ (.A(\mem[12][0] ),
    .X(_0585_));
 sg13g2_buf_1 _3583_ (.A(_2635_),
    .X(_0586_));
 sg13g2_nand2_2 _3584_ (.Y(_0587_),
    .A(_2637_),
    .B(_2647_));
 sg13g2_nor3_1 _3585_ (.A(_0586_),
    .B(_2636_),
    .C(_0587_),
    .Y(_0588_));
 sg13g2_buf_4 _3586_ (.X(_0589_),
    .A(_0588_));
 sg13g2_nand2_2 _3587_ (.Y(_0590_),
    .A(_0566_),
    .B(_0589_));
 sg13g2_mux2_1 _3588_ (.A0(net51),
    .A1(net167),
    .S(_0590_),
    .X(_0013_));
 sg13g2_buf_2 _3589_ (.A(\mem[12][1] ),
    .X(_0591_));
 sg13g2_mux2_1 _3590_ (.A0(net44),
    .A1(_0591_),
    .S(_0590_),
    .X(_0014_));
 sg13g2_buf_1 _3591_ (.A(\mem[12][2] ),
    .X(_0592_));
 sg13g2_mux2_1 _3592_ (.A0(net37),
    .A1(net165),
    .S(_0590_),
    .X(_0015_));
 sg13g2_buf_2 _3593_ (.A(\mem[12][3] ),
    .X(_0593_));
 sg13g2_mux2_1 _3594_ (.A0(net30),
    .A1(_0593_),
    .S(_0590_),
    .X(_0016_));
 sg13g2_buf_1 _3595_ (.A(\mem[13][0] ),
    .X(_0594_));
 sg13g2_nand2_2 _3596_ (.Y(_0595_),
    .A(_2635_),
    .B(_0560_));
 sg13g2_nor2_1 _3597_ (.A(_0587_),
    .B(_0595_),
    .Y(_0596_));
 sg13g2_buf_4 _3598_ (.X(_0597_),
    .A(_0596_));
 sg13g2_nand2_2 _3599_ (.Y(_0598_),
    .A(_0566_),
    .B(_0597_));
 sg13g2_mux2_1 _3600_ (.A0(_2633_),
    .A1(net164),
    .S(_0598_),
    .X(_0017_));
 sg13g2_buf_2 _3601_ (.A(\mem[13][1] ),
    .X(_0599_));
 sg13g2_mux2_1 _3602_ (.A0(_2721_),
    .A1(_0599_),
    .S(_0598_),
    .X(_0018_));
 sg13g2_buf_1 _3603_ (.A(\mem[13][2] ),
    .X(_0600_));
 sg13g2_mux2_1 _3604_ (.A0(net37),
    .A1(net163),
    .S(_0598_),
    .X(_0019_));
 sg13g2_buf_2 _3605_ (.A(\mem[13][3] ),
    .X(_0601_));
 sg13g2_mux2_1 _3606_ (.A0(_0556_),
    .A1(_0601_),
    .S(_0598_),
    .X(_0020_));
 sg13g2_buf_1 _3607_ (.A(\mem[14][0] ),
    .X(_0602_));
 sg13g2_nor3_1 _3608_ (.A(net166),
    .B(_0560_),
    .C(_0587_),
    .Y(_0603_));
 sg13g2_buf_4 _3609_ (.X(_0604_),
    .A(_0603_));
 sg13g2_nand2_2 _3610_ (.Y(_0605_),
    .A(_0566_),
    .B(_0604_));
 sg13g2_mux2_1 _3611_ (.A0(net51),
    .A1(net162),
    .S(_0605_),
    .X(_0021_));
 sg13g2_buf_2 _3612_ (.A(\mem[14][1] ),
    .X(_0606_));
 sg13g2_mux2_1 _3613_ (.A0(net44),
    .A1(_0606_),
    .S(_0605_),
    .X(_0022_));
 sg13g2_buf_1 _3614_ (.A(\mem[14][2] ),
    .X(_0607_));
 sg13g2_mux2_1 _3615_ (.A0(net37),
    .A1(net161),
    .S(_0605_),
    .X(_0023_));
 sg13g2_buf_2 _3616_ (.A(\mem[14][3] ),
    .X(_0608_));
 sg13g2_mux2_1 _3617_ (.A0(net30),
    .A1(_0608_),
    .S(_0605_),
    .X(_0024_));
 sg13g2_buf_1 _3618_ (.A(\mem[15][0] ),
    .X(_0609_));
 sg13g2_nor3_1 _3619_ (.A(_0573_),
    .B(_0560_),
    .C(_0587_),
    .Y(_0610_));
 sg13g2_buf_4 _3620_ (.X(_0611_),
    .A(_0610_));
 sg13g2_nand2_2 _3621_ (.Y(_0612_),
    .A(_0566_),
    .B(_0611_));
 sg13g2_mux2_1 _3622_ (.A0(net51),
    .A1(net160),
    .S(_0612_),
    .X(_0025_));
 sg13g2_buf_2 _3623_ (.A(\mem[15][1] ),
    .X(_0613_));
 sg13g2_mux2_1 _3624_ (.A0(net44),
    .A1(_0613_),
    .S(_0612_),
    .X(_0026_));
 sg13g2_buf_1 _3625_ (.A(\mem[15][2] ),
    .X(_0614_));
 sg13g2_mux2_1 _3626_ (.A0(net37),
    .A1(net159),
    .S(_0612_),
    .X(_0027_));
 sg13g2_buf_2 _3627_ (.A(\mem[15][3] ),
    .X(_0615_));
 sg13g2_mux2_1 _3628_ (.A0(net30),
    .A1(_0615_),
    .S(_0612_),
    .X(_0028_));
 sg13g2_buf_1 _3629_ (.A(\mem[16][0] ),
    .X(_0616_));
 sg13g2_nand2b_1 _3630_ (.Y(_0617_),
    .B(net177),
    .A_N(net171));
 sg13g2_nor3_1 _3631_ (.A(net176),
    .B(net58),
    .C(_0617_),
    .Y(_0618_));
 sg13g2_buf_4 _3632_ (.X(_0619_),
    .A(_0618_));
 sg13g2_nand2_2 _3633_ (.Y(_0620_),
    .A(_2639_),
    .B(_0619_));
 sg13g2_mux2_1 _3634_ (.A0(net51),
    .A1(net158),
    .S(_0620_),
    .X(_0029_));
 sg13g2_buf_2 _3635_ (.A(\mem[16][1] ),
    .X(_0621_));
 sg13g2_mux2_1 _3636_ (.A0(net44),
    .A1(_0621_),
    .S(_0620_),
    .X(_0030_));
 sg13g2_buf_1 _3637_ (.A(\mem[16][2] ),
    .X(_0622_));
 sg13g2_mux2_1 _3638_ (.A0(net37),
    .A1(net157),
    .S(_0620_),
    .X(_0031_));
 sg13g2_buf_2 _3639_ (.A(\mem[16][3] ),
    .X(_0623_));
 sg13g2_mux2_1 _3640_ (.A0(net30),
    .A1(_0623_),
    .S(_0620_),
    .X(_0032_));
 sg13g2_buf_1 _3641_ (.A(\mem[17][0] ),
    .X(_0624_));
 sg13g2_nand3_1 _3642_ (.B(_2608_),
    .C(_2606_),
    .A(_2607_),
    .Y(_0625_));
 sg13g2_buf_1 _3643_ (.A(_0625_),
    .X(_0626_));
 sg13g2_or3_1 _3644_ (.A(_0574_),
    .B(net58),
    .C(_0595_),
    .X(_0627_));
 sg13g2_nand2_1 _3645_ (.Y(_0628_),
    .A(net62),
    .B(_0627_));
 sg13g2_buf_2 _3646_ (.A(_0628_),
    .X(_0629_));
 sg13g2_nand2_2 _3647_ (.Y(_0630_),
    .A(_0619_),
    .B(_0629_));
 sg13g2_mux2_1 _3648_ (.A0(_2633_),
    .A1(net156),
    .S(_0630_),
    .X(_0033_));
 sg13g2_buf_1 _3649_ (.A(\mem[17][1] ),
    .X(_0631_));
 sg13g2_inv_1 _3650_ (.Y(_0632_),
    .A(net155));
 sg13g2_buf_1 _3651_ (.A(net45),
    .X(_0633_));
 sg13g2_nor2_1 _3652_ (.A(_0633_),
    .B(_0630_),
    .Y(_0634_));
 sg13g2_a21oi_1 _3653_ (.A1(_0632_),
    .A2(_0630_),
    .Y(_0034_),
    .B1(_0634_));
 sg13g2_buf_1 _3654_ (.A(\mem[17][2] ),
    .X(_0635_));
 sg13g2_mux2_1 _3655_ (.A0(_0426_),
    .A1(net154),
    .S(_0630_),
    .X(_0035_));
 sg13g2_buf_1 _3656_ (.A(\mem[17][3] ),
    .X(_0636_));
 sg13g2_mux2_1 _3657_ (.A0(_0556_),
    .A1(net153),
    .S(_0630_),
    .X(_0036_));
 sg13g2_buf_1 _3658_ (.A(\mem[18][0] ),
    .X(_0637_));
 sg13g2_nand2_2 _3659_ (.Y(_0638_),
    .A(_0562_),
    .B(_0619_));
 sg13g2_mux2_1 _3660_ (.A0(net51),
    .A1(net152),
    .S(_0638_),
    .X(_0037_));
 sg13g2_buf_1 _3661_ (.A(\mem[18][1] ),
    .X(_0639_));
 sg13g2_inv_1 _3662_ (.Y(_0640_),
    .A(net151));
 sg13g2_nor2_1 _3663_ (.A(net43),
    .B(_0638_),
    .Y(_0641_));
 sg13g2_a21oi_1 _3664_ (.A1(_0640_),
    .A2(_0638_),
    .Y(_0038_),
    .B1(_0641_));
 sg13g2_buf_1 _3665_ (.A(\mem[18][2] ),
    .X(_0642_));
 sg13g2_mux2_1 _3666_ (.A0(_0426_),
    .A1(net150),
    .S(_0638_),
    .X(_0039_));
 sg13g2_buf_1 _3667_ (.A(\mem[18][3] ),
    .X(_0643_));
 sg13g2_mux2_1 _3668_ (.A0(net30),
    .A1(net149),
    .S(_0638_),
    .X(_0040_));
 sg13g2_buf_1 _3669_ (.A(\mem[19][0] ),
    .X(_0644_));
 sg13g2_nand2_2 _3670_ (.Y(_0645_),
    .A(_0576_),
    .B(_0619_));
 sg13g2_mux2_1 _3671_ (.A0(net51),
    .A1(net148),
    .S(_0645_),
    .X(_0041_));
 sg13g2_buf_1 _3672_ (.A(\mem[19][1] ),
    .X(_0646_));
 sg13g2_inv_1 _3673_ (.Y(_0647_),
    .A(net147));
 sg13g2_buf_1 _3674_ (.A(net45),
    .X(_0648_));
 sg13g2_nor2_1 _3675_ (.A(net42),
    .B(_0645_),
    .Y(_0649_));
 sg13g2_a21oi_1 _3676_ (.A1(_0647_),
    .A2(_0645_),
    .Y(_0042_),
    .B1(_0649_));
 sg13g2_buf_1 _3677_ (.A(_0425_),
    .X(_0650_));
 sg13g2_buf_1 _3678_ (.A(\mem[19][2] ),
    .X(_0651_));
 sg13g2_mux2_1 _3679_ (.A0(_0650_),
    .A1(net146),
    .S(_0645_),
    .X(_0043_));
 sg13g2_buf_8 _3680_ (.A(net31),
    .X(_0652_));
 sg13g2_buf_1 _3681_ (.A(\mem[19][3] ),
    .X(_0653_));
 sg13g2_mux2_1 _3682_ (.A0(_0652_),
    .A1(net145),
    .S(_0645_),
    .X(_0044_));
 sg13g2_buf_1 _3683_ (.A(\mem[1][0] ),
    .X(_0654_));
 sg13g2_buf_1 _3684_ (.A(net52),
    .X(_0655_));
 sg13g2_o21ai_1 _3685_ (.B1(_2647_),
    .Y(_0656_),
    .A1(net169),
    .A2(_0595_));
 sg13g2_and2_1 _3686_ (.A(_2644_),
    .B(_0656_),
    .X(_0657_));
 sg13g2_buf_2 _3687_ (.A(_0657_),
    .X(_0658_));
 sg13g2_mux2_1 _3688_ (.A0(net144),
    .A1(net50),
    .S(_0658_),
    .X(_0045_));
 sg13g2_buf_2 _3689_ (.A(\mem[1][1] ),
    .X(_0659_));
 sg13g2_mux2_1 _3690_ (.A0(_0659_),
    .A1(_0633_),
    .S(_0658_),
    .X(_0046_));
 sg13g2_buf_1 _3691_ (.A(\mem[1][2] ),
    .X(_0660_));
 sg13g2_buf_1 _3692_ (.A(net38),
    .X(_0661_));
 sg13g2_mux2_1 _3693_ (.A0(net143),
    .A1(net35),
    .S(_0658_),
    .X(_0047_));
 sg13g2_buf_2 _3694_ (.A(\mem[1][3] ),
    .X(_0662_));
 sg13g2_buf_8 _3695_ (.A(net31),
    .X(_0663_));
 sg13g2_mux2_1 _3696_ (.A0(_0662_),
    .A1(net28),
    .S(_0658_),
    .X(_0048_));
 sg13g2_buf_1 _3697_ (.A(net52),
    .X(_0664_));
 sg13g2_buf_1 _3698_ (.A(\mem[20][0] ),
    .X(_0665_));
 sg13g2_nand2_2 _3699_ (.Y(_0666_),
    .A(_0589_),
    .B(_0619_));
 sg13g2_mux2_1 _3700_ (.A0(net49),
    .A1(net142),
    .S(_0666_),
    .X(_0049_));
 sg13g2_buf_1 _3701_ (.A(\mem[20][1] ),
    .X(_0667_));
 sg13g2_inv_1 _3702_ (.Y(_0668_),
    .A(net141));
 sg13g2_nor2_1 _3703_ (.A(net42),
    .B(_0666_),
    .Y(_0669_));
 sg13g2_a21oi_1 _3704_ (.A1(_0668_),
    .A2(_0666_),
    .Y(_0050_),
    .B1(_0669_));
 sg13g2_buf_1 _3705_ (.A(\mem[20][2] ),
    .X(_0670_));
 sg13g2_mux2_1 _3706_ (.A0(net36),
    .A1(net140),
    .S(_0666_),
    .X(_0051_));
 sg13g2_buf_1 _3707_ (.A(\mem[20][3] ),
    .X(_0671_));
 sg13g2_mux2_1 _3708_ (.A0(net29),
    .A1(net139),
    .S(_0666_),
    .X(_0052_));
 sg13g2_buf_1 _3709_ (.A(\mem[21][0] ),
    .X(_0672_));
 sg13g2_nand2_2 _3710_ (.Y(_0673_),
    .A(_0597_),
    .B(_0619_));
 sg13g2_mux2_1 _3711_ (.A0(net49),
    .A1(_0672_),
    .S(_0673_),
    .X(_0053_));
 sg13g2_buf_1 _3712_ (.A(\mem[21][1] ),
    .X(_0674_));
 sg13g2_inv_1 _3713_ (.Y(_0675_),
    .A(net137));
 sg13g2_nor2_1 _3714_ (.A(net42),
    .B(_0673_),
    .Y(_0676_));
 sg13g2_a21oi_1 _3715_ (.A1(_0675_),
    .A2(_0673_),
    .Y(_0054_),
    .B1(_0676_));
 sg13g2_buf_1 _3716_ (.A(\mem[21][2] ),
    .X(_0677_));
 sg13g2_mux2_1 _3717_ (.A0(net36),
    .A1(net136),
    .S(_0673_),
    .X(_0055_));
 sg13g2_buf_1 _3718_ (.A(\mem[21][3] ),
    .X(_0678_));
 sg13g2_mux2_1 _3719_ (.A0(net29),
    .A1(net135),
    .S(_0673_),
    .X(_0056_));
 sg13g2_buf_1 _3720_ (.A(\mem[22][0] ),
    .X(_0679_));
 sg13g2_nand2_2 _3721_ (.Y(_0680_),
    .A(_0604_),
    .B(_0619_));
 sg13g2_mux2_1 _3722_ (.A0(net49),
    .A1(_0679_),
    .S(_0680_),
    .X(_0057_));
 sg13g2_buf_1 _3723_ (.A(\mem[22][1] ),
    .X(_0681_));
 sg13g2_inv_1 _3724_ (.Y(_0682_),
    .A(net133));
 sg13g2_nor2_1 _3725_ (.A(net42),
    .B(_0680_),
    .Y(_0683_));
 sg13g2_a21oi_1 _3726_ (.A1(_0682_),
    .A2(_0680_),
    .Y(_0058_),
    .B1(_0683_));
 sg13g2_buf_1 _3727_ (.A(\mem[22][2] ),
    .X(_0684_));
 sg13g2_mux2_1 _3728_ (.A0(net36),
    .A1(net132),
    .S(_0680_),
    .X(_0059_));
 sg13g2_buf_1 _3729_ (.A(\mem[22][3] ),
    .X(_0685_));
 sg13g2_mux2_1 _3730_ (.A0(net29),
    .A1(net131),
    .S(_0680_),
    .X(_0060_));
 sg13g2_buf_1 _3731_ (.A(\mem[23][0] ),
    .X(_0686_));
 sg13g2_nand2_2 _3732_ (.Y(_0687_),
    .A(_0611_),
    .B(_0619_));
 sg13g2_mux2_1 _3733_ (.A0(net49),
    .A1(_0686_),
    .S(_0687_),
    .X(_0061_));
 sg13g2_buf_2 _3734_ (.A(\mem[23][1] ),
    .X(_0688_));
 sg13g2_inv_1 _3735_ (.Y(_0689_),
    .A(_0688_));
 sg13g2_nor2_1 _3736_ (.A(net42),
    .B(_0687_),
    .Y(_0690_));
 sg13g2_a21oi_1 _3737_ (.A1(_0689_),
    .A2(_0687_),
    .Y(_0062_),
    .B1(_0690_));
 sg13g2_buf_1 _3738_ (.A(\mem[23][2] ),
    .X(_0691_));
 sg13g2_mux2_1 _3739_ (.A0(_0650_),
    .A1(net129),
    .S(_0687_),
    .X(_0063_));
 sg13g2_buf_1 _3740_ (.A(\mem[23][3] ),
    .X(_0692_));
 sg13g2_mux2_1 _3741_ (.A0(_0652_),
    .A1(_0692_),
    .S(_0687_),
    .X(_0064_));
 sg13g2_buf_1 _3742_ (.A(\mem[24][0] ),
    .X(_0693_));
 sg13g2_nand2_1 _3743_ (.Y(_0694_),
    .A(net171),
    .B(net177));
 sg13g2_nor3_1 _3744_ (.A(net176),
    .B(net58),
    .C(_0694_),
    .Y(_0695_));
 sg13g2_buf_4 _3745_ (.X(_0696_),
    .A(_0695_));
 sg13g2_nand2_2 _3746_ (.Y(_0697_),
    .A(_2639_),
    .B(_0696_));
 sg13g2_mux2_1 _3747_ (.A0(net49),
    .A1(net127),
    .S(_0697_),
    .X(_0065_));
 sg13g2_buf_2 _3748_ (.A(\mem[24][1] ),
    .X(_0698_));
 sg13g2_inv_1 _3749_ (.Y(_0699_),
    .A(_0698_));
 sg13g2_nor2_1 _3750_ (.A(net42),
    .B(_0697_),
    .Y(_0700_));
 sg13g2_a21oi_1 _3751_ (.A1(_0699_),
    .A2(_0697_),
    .Y(_0066_),
    .B1(_0700_));
 sg13g2_buf_2 _3752_ (.A(\mem[24][2] ),
    .X(_0701_));
 sg13g2_mux2_1 _3753_ (.A0(net36),
    .A1(_0701_),
    .S(_0697_),
    .X(_0067_));
 sg13g2_buf_1 _3754_ (.A(\mem[24][3] ),
    .X(_0702_));
 sg13g2_mux2_1 _3755_ (.A0(net29),
    .A1(net126),
    .S(_0697_),
    .X(_0068_));
 sg13g2_buf_1 _3756_ (.A(\mem[25][0] ),
    .X(_0703_));
 sg13g2_nand2_2 _3757_ (.Y(_0704_),
    .A(_0629_),
    .B(_0696_));
 sg13g2_mux2_1 _3758_ (.A0(net49),
    .A1(net125),
    .S(_0704_),
    .X(_0069_));
 sg13g2_buf_2 _3759_ (.A(\mem[25][1] ),
    .X(_0705_));
 sg13g2_inv_1 _3760_ (.Y(_0706_),
    .A(_0705_));
 sg13g2_nor2_1 _3761_ (.A(_0648_),
    .B(_0704_),
    .Y(_0707_));
 sg13g2_a21oi_1 _3762_ (.A1(_0706_),
    .A2(_0704_),
    .Y(_0070_),
    .B1(_0707_));
 sg13g2_buf_2 _3763_ (.A(\mem[25][2] ),
    .X(_0708_));
 sg13g2_mux2_1 _3764_ (.A0(net36),
    .A1(_0708_),
    .S(_0704_),
    .X(_0071_));
 sg13g2_buf_1 _3765_ (.A(\mem[25][3] ),
    .X(_0709_));
 sg13g2_mux2_1 _3766_ (.A0(net29),
    .A1(net124),
    .S(_0704_),
    .X(_0072_));
 sg13g2_buf_1 _3767_ (.A(\mem[26][0] ),
    .X(_0710_));
 sg13g2_nand2_2 _3768_ (.Y(_0711_),
    .A(_0562_),
    .B(_0696_));
 sg13g2_mux2_1 _3769_ (.A0(net49),
    .A1(net123),
    .S(_0711_),
    .X(_0073_));
 sg13g2_buf_2 _3770_ (.A(\mem[26][1] ),
    .X(_0712_));
 sg13g2_inv_1 _3771_ (.Y(_0713_),
    .A(_0712_));
 sg13g2_nor2_1 _3772_ (.A(net42),
    .B(_0711_),
    .Y(_0714_));
 sg13g2_a21oi_1 _3773_ (.A1(_0713_),
    .A2(_0711_),
    .Y(_0074_),
    .B1(_0714_));
 sg13g2_buf_2 _3774_ (.A(\mem[26][2] ),
    .X(_0715_));
 sg13g2_mux2_1 _3775_ (.A0(net36),
    .A1(_0715_),
    .S(_0711_),
    .X(_0075_));
 sg13g2_buf_1 _3776_ (.A(\mem[26][3] ),
    .X(_0716_));
 sg13g2_mux2_1 _3777_ (.A0(net29),
    .A1(net122),
    .S(_0711_),
    .X(_0076_));
 sg13g2_buf_2 _3778_ (.A(\mem[27][0] ),
    .X(_0717_));
 sg13g2_inv_1 _3779_ (.Y(_0718_),
    .A(_0717_));
 sg13g2_nand2_2 _3780_ (.Y(_0719_),
    .A(_0576_),
    .B(_0696_));
 sg13g2_nor2_1 _3781_ (.A(_2632_),
    .B(_0719_),
    .Y(_0720_));
 sg13g2_a21oi_1 _3782_ (.A1(_0718_),
    .A2(_0719_),
    .Y(_0077_),
    .B1(_0720_));
 sg13g2_buf_2 _3783_ (.A(\mem[27][1] ),
    .X(_0721_));
 sg13g2_inv_1 _3784_ (.Y(_0722_),
    .A(_0721_));
 sg13g2_nor2_1 _3785_ (.A(net42),
    .B(_0719_),
    .Y(_0723_));
 sg13g2_a21oi_1 _3786_ (.A1(_0722_),
    .A2(_0719_),
    .Y(_0078_),
    .B1(_0723_));
 sg13g2_buf_1 _3787_ (.A(\mem[27][2] ),
    .X(_0724_));
 sg13g2_buf_1 _3788_ (.A(net121),
    .X(_0725_));
 sg13g2_mux2_1 _3789_ (.A0(net36),
    .A1(net78),
    .S(_0719_),
    .X(_0079_));
 sg13g2_buf_1 _3790_ (.A(\mem[27][3] ),
    .X(_0726_));
 sg13g2_buf_1 _3791_ (.A(_0726_),
    .X(_0727_));
 sg13g2_mux2_1 _3792_ (.A0(net29),
    .A1(net77),
    .S(_0719_),
    .X(_0080_));
 sg13g2_buf_1 _3793_ (.A(\mem[28][0] ),
    .X(_0728_));
 sg13g2_nand2_2 _3794_ (.Y(_0729_),
    .A(_0589_),
    .B(_0696_));
 sg13g2_mux2_1 _3795_ (.A0(_0664_),
    .A1(net120),
    .S(_0729_),
    .X(_0081_));
 sg13g2_buf_1 _3796_ (.A(\mem[28][1] ),
    .X(_0730_));
 sg13g2_inv_1 _3797_ (.Y(_0731_),
    .A(net119));
 sg13g2_nor2_1 _3798_ (.A(_0648_),
    .B(_0729_),
    .Y(_0732_));
 sg13g2_a21oi_1 _3799_ (.A1(_0731_),
    .A2(_0729_),
    .Y(_0082_),
    .B1(_0732_));
 sg13g2_buf_1 _3800_ (.A(\mem[28][2] ),
    .X(_0733_));
 sg13g2_mux2_1 _3801_ (.A0(net36),
    .A1(net118),
    .S(_0729_),
    .X(_0083_));
 sg13g2_buf_1 _3802_ (.A(\mem[28][3] ),
    .X(_0734_));
 sg13g2_mux2_1 _3803_ (.A0(net29),
    .A1(net117),
    .S(_0729_),
    .X(_0084_));
 sg13g2_buf_1 _3804_ (.A(\mem[29][0] ),
    .X(_0735_));
 sg13g2_nand2_2 _3805_ (.Y(_0736_),
    .A(_0597_),
    .B(_0696_));
 sg13g2_mux2_1 _3806_ (.A0(_0664_),
    .A1(net116),
    .S(_0736_),
    .X(_0085_));
 sg13g2_buf_2 _3807_ (.A(\mem[29][1] ),
    .X(_0737_));
 sg13g2_inv_1 _3808_ (.Y(_0738_),
    .A(_0737_));
 sg13g2_nor2_1 _3809_ (.A(net45),
    .B(_0736_),
    .Y(_0739_));
 sg13g2_a21oi_1 _3810_ (.A1(_0738_),
    .A2(_0736_),
    .Y(_0086_),
    .B1(_0739_));
 sg13g2_buf_1 _3811_ (.A(net38),
    .X(_0740_));
 sg13g2_buf_2 _3812_ (.A(\mem[29][2] ),
    .X(_0741_));
 sg13g2_mux2_1 _3813_ (.A0(net34),
    .A1(_0741_),
    .S(_0736_),
    .X(_0087_));
 sg13g2_buf_8 _3814_ (.A(net31),
    .X(_0742_));
 sg13g2_buf_1 _3815_ (.A(\mem[29][3] ),
    .X(_0743_));
 sg13g2_mux2_1 _3816_ (.A0(net27),
    .A1(net115),
    .S(_0736_),
    .X(_0088_));
 sg13g2_buf_1 _3817_ (.A(\mem[2][0] ),
    .X(_0744_));
 sg13g2_nand2_2 _3818_ (.Y(_0745_),
    .A(_2644_),
    .B(_0562_));
 sg13g2_mux2_1 _3819_ (.A0(net49),
    .A1(net114),
    .S(_0745_),
    .X(_0089_));
 sg13g2_buf_2 _3820_ (.A(\mem[2][1] ),
    .X(_0746_));
 sg13g2_mux2_1 _3821_ (.A0(net44),
    .A1(_0746_),
    .S(_0745_),
    .X(_0090_));
 sg13g2_buf_1 _3822_ (.A(\mem[2][2] ),
    .X(_0747_));
 sg13g2_mux2_1 _3823_ (.A0(net34),
    .A1(net113),
    .S(_0745_),
    .X(_0091_));
 sg13g2_buf_2 _3824_ (.A(\mem[2][3] ),
    .X(_0748_));
 sg13g2_mux2_1 _3825_ (.A0(net27),
    .A1(_0748_),
    .S(_0745_),
    .X(_0092_));
 sg13g2_buf_1 _3826_ (.A(net52),
    .X(_0749_));
 sg13g2_buf_1 _3827_ (.A(\mem[30][0] ),
    .X(_0750_));
 sg13g2_nand2_2 _3828_ (.Y(_0751_),
    .A(_0604_),
    .B(_0696_));
 sg13g2_mux2_1 _3829_ (.A0(_0749_),
    .A1(net112),
    .S(_0751_),
    .X(_0093_));
 sg13g2_buf_1 _3830_ (.A(\mem[30][1] ),
    .X(_0752_));
 sg13g2_inv_1 _3831_ (.Y(_0753_),
    .A(net111));
 sg13g2_nor2_1 _3832_ (.A(net45),
    .B(_0751_),
    .Y(_0754_));
 sg13g2_a21oi_1 _3833_ (.A1(_0753_),
    .A2(_0751_),
    .Y(_0094_),
    .B1(_0754_));
 sg13g2_buf_1 _3834_ (.A(\mem[30][2] ),
    .X(_0755_));
 sg13g2_mux2_1 _3835_ (.A0(_0740_),
    .A1(net110),
    .S(_0751_),
    .X(_0095_));
 sg13g2_buf_1 _3836_ (.A(\mem[30][3] ),
    .X(_0756_));
 sg13g2_mux2_1 _3837_ (.A0(_0742_),
    .A1(net109),
    .S(_0751_),
    .X(_0096_));
 sg13g2_buf_1 _3838_ (.A(\mem[31][0] ),
    .X(_0757_));
 sg13g2_nand2_2 _3839_ (.Y(_0758_),
    .A(_0611_),
    .B(_0696_));
 sg13g2_mux2_1 _3840_ (.A0(_0749_),
    .A1(net108),
    .S(_0758_),
    .X(_0097_));
 sg13g2_buf_1 _3841_ (.A(\mem[31][1] ),
    .X(_0759_));
 sg13g2_inv_1 _3842_ (.Y(_0760_),
    .A(net107));
 sg13g2_nor2_1 _3843_ (.A(_2720_),
    .B(_0758_),
    .Y(_0761_));
 sg13g2_a21oi_1 _3844_ (.A1(_0760_),
    .A2(_0758_),
    .Y(_0098_),
    .B1(_0761_));
 sg13g2_buf_1 _3845_ (.A(\mem[31][2] ),
    .X(_0762_));
 sg13g2_mux2_1 _3846_ (.A0(_0740_),
    .A1(net106),
    .S(_0758_),
    .X(_0099_));
 sg13g2_buf_1 _3847_ (.A(\mem[31][3] ),
    .X(_0763_));
 sg13g2_mux2_1 _3848_ (.A0(_0742_),
    .A1(net105),
    .S(_0758_),
    .X(_0100_));
 sg13g2_buf_1 _3849_ (.A(\mem[32][0] ),
    .X(_0764_));
 sg13g2_nor2_1 _3850_ (.A(_2640_),
    .B(net177),
    .Y(_0765_));
 sg13g2_a21oi_1 _3851_ (.A1(net176),
    .A2(_0765_),
    .Y(_0766_),
    .B1(_2611_));
 sg13g2_buf_2 _3852_ (.A(_0766_),
    .X(_0767_));
 sg13g2_nor2b_1 _3853_ (.A(_0767_),
    .B_N(_2639_),
    .Y(_0768_));
 sg13g2_buf_2 _3854_ (.A(_0768_),
    .X(_0769_));
 sg13g2_mux2_1 _3855_ (.A0(net104),
    .A1(net50),
    .S(_0769_),
    .X(_0101_));
 sg13g2_buf_1 _3856_ (.A(\mem[32][1] ),
    .X(_0770_));
 sg13g2_inv_1 _3857_ (.Y(_0771_),
    .A(net103));
 sg13g2_nand2_1 _3858_ (.Y(_0772_),
    .A(net43),
    .B(_0769_));
 sg13g2_o21ai_1 _3859_ (.B1(_0772_),
    .Y(_0102_),
    .A1(_0771_),
    .A2(_0769_));
 sg13g2_buf_1 _3860_ (.A(\mem[32][2] ),
    .X(_0773_));
 sg13g2_mux2_1 _3861_ (.A0(net102),
    .A1(net35),
    .S(_0769_),
    .X(_0103_));
 sg13g2_buf_1 _3862_ (.A(\mem[32][3] ),
    .X(_0774_));
 sg13g2_mux2_1 _3863_ (.A0(net101),
    .A1(net28),
    .S(_0769_),
    .X(_0104_));
 sg13g2_a21oi_2 _3864_ (.B1(_0767_),
    .Y(_0775_),
    .A2(_0627_),
    .A1(net62));
 sg13g2_mux2_1 _3865_ (.A0(net17),
    .A1(net50),
    .S(_0775_),
    .X(_0105_));
 sg13g2_mux2_1 _3866_ (.A0(net18),
    .A1(net43),
    .S(_0775_),
    .X(_0106_));
 sg13g2_mux2_1 _3867_ (.A0(net19),
    .A1(net35),
    .S(_0775_),
    .X(_0107_));
 sg13g2_mux2_1 _3868_ (.A0(net20),
    .A1(net28),
    .S(_0775_),
    .X(_0108_));
 sg13g2_nand3b_1 _3869_ (.B(_0549_),
    .C(_0550_),
    .Y(_0776_),
    .A_N(_0443_));
 sg13g2_a21o_1 _3870_ (.A2(_0438_),
    .A1(_0416_),
    .B1(_0442_),
    .X(_0777_));
 sg13g2_a221oi_1 _3871_ (.B2(_0550_),
    .C1(_0777_),
    .B1(_0549_),
    .A1(_0428_),
    .Y(_0778_),
    .A2(_0437_));
 sg13g2_a21oi_2 _3872_ (.B1(_0778_),
    .Y(_0779_),
    .A2(_0776_),
    .A1(_0436_));
 sg13g2_nand2_1 _3873_ (.Y(_0780_),
    .A(_2787_),
    .B(_2792_));
 sg13g2_nor2_1 _3874_ (.A(_0780_),
    .B(_0540_),
    .Y(_0781_));
 sg13g2_a21oi_1 _3875_ (.A1(_0780_),
    .A2(_0540_),
    .Y(_0782_),
    .B1(_0403_));
 sg13g2_nor2_1 _3876_ (.A(_0781_),
    .B(_0782_),
    .Y(_0783_));
 sg13g2_o21ai_1 _3877_ (.B1(_0783_),
    .Y(_0784_),
    .A1(_0524_),
    .A2(_0530_));
 sg13g2_nand2_1 _3878_ (.Y(_0785_),
    .A(_0524_),
    .B(_0530_));
 sg13g2_nor2_1 _3879_ (.A(_0518_),
    .B(_0520_),
    .Y(_0786_));
 sg13g2_a21oi_1 _3880_ (.A1(_0518_),
    .A2(_0520_),
    .Y(_0787_),
    .B1(_0512_));
 sg13g2_or2_1 _3881_ (.X(_0788_),
    .B(_0787_),
    .A(_0786_));
 sg13g2_buf_1 _3882_ (.A(_0788_),
    .X(_0789_));
 sg13g2_inv_1 _3883_ (.Y(_0790_),
    .A(_0789_));
 sg13g2_nand2_1 _3884_ (.Y(_0791_),
    .A(_0469_),
    .B(_0475_));
 sg13g2_o21ai_1 _3885_ (.B1(_0472_),
    .Y(_0792_),
    .A1(_0469_),
    .A2(_0475_));
 sg13g2_xnor2_1 _3886_ (.Y(_0793_),
    .A(\products[14][4] ),
    .B(\products[1][4] ));
 sg13g2_xnor2_1 _3887_ (.Y(_0794_),
    .A(\products[15][4] ),
    .B(_0793_));
 sg13g2_or2_1 _3888_ (.X(_0795_),
    .B(_0467_),
    .A(_0466_));
 sg13g2_a21o_1 _3889_ (.A2(_0467_),
    .A1(_0466_),
    .B1(\products[12][3] ),
    .X(_0796_));
 sg13g2_nand2_1 _3890_ (.Y(_0797_),
    .A(_0448_),
    .B(_0449_));
 sg13g2_o21ai_1 _3891_ (.B1(\products[15][3] ),
    .Y(_0798_),
    .A1(_0448_),
    .A2(_0449_));
 sg13g2_nand4_1 _3892_ (.B(_0796_),
    .C(_0797_),
    .A(_0795_),
    .Y(_0799_),
    .D(_0798_));
 sg13g2_nand2_1 _3893_ (.Y(_0800_),
    .A(_0466_),
    .B(_0467_));
 sg13g2_o21ai_1 _3894_ (.B1(\products[12][3] ),
    .Y(_0801_),
    .A1(_0466_),
    .A2(_0467_));
 sg13g2_or2_1 _3895_ (.X(_0802_),
    .B(_0449_),
    .A(_0448_));
 sg13g2_a21o_1 _3896_ (.A2(_0449_),
    .A1(_0448_),
    .B1(\products[15][3] ),
    .X(_0803_));
 sg13g2_nand4_1 _3897_ (.B(_0801_),
    .C(_0802_),
    .A(_0800_),
    .Y(_0804_),
    .D(_0803_));
 sg13g2_nand3_1 _3898_ (.B(_0799_),
    .C(_0804_),
    .A(_0794_),
    .Y(_0805_));
 sg13g2_a21o_1 _3899_ (.A2(_0804_),
    .A1(_0799_),
    .B1(_0794_),
    .X(_0806_));
 sg13g2_a22oi_1 _3900_ (.Y(_0807_),
    .B1(_0805_),
    .B2(_0806_),
    .A2(_0792_),
    .A1(_0791_));
 sg13g2_and4_1 _3901_ (.A(_0791_),
    .B(_0792_),
    .C(_0805_),
    .D(_0806_),
    .X(_0808_));
 sg13g2_buf_1 _3902_ (.A(_0808_),
    .X(_0809_));
 sg13g2_xnor2_1 _3903_ (.Y(_0810_),
    .A(\products[11][4] ),
    .B(\products[13][4] ));
 sg13g2_xnor2_1 _3904_ (.Y(_0811_),
    .A(\products[12][4] ),
    .B(_0810_));
 sg13g2_a21o_1 _3905_ (.A2(\products[10][3] ),
    .A1(_0473_),
    .B1(\products[0][3] ),
    .X(_0812_));
 sg13g2_o21ai_1 _3906_ (.B1(_0812_),
    .Y(_0813_),
    .A1(_0473_),
    .A2(\products[10][3] ));
 sg13g2_buf_1 _3907_ (.A(\prev_acc[4] ),
    .X(_0814_));
 sg13g2_xnor2_1 _3908_ (.Y(_0815_),
    .A(_0814_),
    .B(\products[10][4] ));
 sg13g2_xnor2_1 _3909_ (.Y(_0816_),
    .A(\products[0][4] ),
    .B(_0815_));
 sg13g2_xnor2_1 _3910_ (.Y(_0817_),
    .A(_0813_),
    .B(_0816_));
 sg13g2_xnor2_1 _3911_ (.Y(_0818_),
    .A(_0811_),
    .B(_0817_));
 sg13g2_o21ai_1 _3912_ (.B1(_0818_),
    .Y(_0819_),
    .A1(_0807_),
    .A2(_0809_));
 sg13g2_or3_1 _3913_ (.A(_0818_),
    .B(_0807_),
    .C(_0809_),
    .X(_0820_));
 sg13g2_buf_1 _3914_ (.A(_0820_),
    .X(_0821_));
 sg13g2_nand2_1 _3915_ (.Y(_0822_),
    .A(_0819_),
    .B(_0821_));
 sg13g2_a21o_1 _3916_ (.A2(_0480_),
    .A1(_0479_),
    .B1(_0465_),
    .X(_0823_));
 sg13g2_nand2_1 _3917_ (.Y(_0824_),
    .A(_0490_),
    .B(_0495_));
 sg13g2_o21ai_1 _3918_ (.B1(_0493_),
    .Y(_0825_),
    .A1(_0490_),
    .A2(_0495_));
 sg13g2_nand2_1 _3919_ (.Y(_0826_),
    .A(_2764_),
    .B(_2765_));
 sg13g2_o21ai_1 _3920_ (.B1(\products[15][2] ),
    .Y(_0827_),
    .A1(_2764_),
    .A2(_2765_));
 sg13g2_a22oi_1 _3921_ (.Y(_0828_),
    .B1(_0826_),
    .B2(_0827_),
    .A2(_0454_),
    .A1(_0452_));
 sg13g2_nand4_1 _3922_ (.B(_0454_),
    .C(_0826_),
    .A(_0452_),
    .Y(_0829_),
    .D(_0827_));
 sg13g2_o21ai_1 _3923_ (.B1(_0829_),
    .Y(_0830_),
    .A1(_0451_),
    .A2(_0828_));
 sg13g2_a21o_1 _3924_ (.A2(_0825_),
    .A1(_0824_),
    .B1(_0830_),
    .X(_0831_));
 sg13g2_nand3_1 _3925_ (.B(_0824_),
    .C(_0825_),
    .A(_0830_),
    .Y(_0832_));
 sg13g2_xnor2_1 _3926_ (.Y(_0833_),
    .A(\products[2][4] ),
    .B(\products[4][4] ));
 sg13g2_xnor2_1 _3927_ (.Y(_0834_),
    .A(\products[3][4] ),
    .B(_0833_));
 sg13g2_nor2_1 _3928_ (.A(\products[2][3] ),
    .B(\products[4][3] ),
    .Y(_0835_));
 sg13g2_a21oi_1 _3929_ (.A1(\products[2][3] ),
    .A2(\products[4][3] ),
    .Y(_0836_),
    .B1(\products[3][3] ));
 sg13g2_nor2_1 _3930_ (.A(_0835_),
    .B(_0836_),
    .Y(_0837_));
 sg13g2_xnor2_1 _3931_ (.Y(_0838_),
    .A(\products[5][4] ),
    .B(\products[7][4] ));
 sg13g2_xnor2_1 _3932_ (.Y(_0839_),
    .A(\products[6][4] ),
    .B(_0838_));
 sg13g2_xnor2_1 _3933_ (.Y(_0840_),
    .A(_0837_),
    .B(_0839_));
 sg13g2_xnor2_1 _3934_ (.Y(_0841_),
    .A(_0834_),
    .B(_0840_));
 sg13g2_a21o_1 _3935_ (.A2(_0832_),
    .A1(_0831_),
    .B1(_0841_),
    .X(_0842_));
 sg13g2_nand3_1 _3936_ (.B(_0831_),
    .C(_0832_),
    .A(_0841_),
    .Y(_0843_));
 sg13g2_nand2_1 _3937_ (.Y(_0844_),
    .A(_0842_),
    .B(_0843_));
 sg13g2_xor2_1 _3938_ (.B(_0844_),
    .A(_0823_),
    .X(_0845_));
 sg13g2_xnor2_1 _3939_ (.Y(_0846_),
    .A(_0822_),
    .B(_0845_));
 sg13g2_nand4_1 _3940_ (.B(_0481_),
    .C(_0498_),
    .A(_0478_),
    .Y(_0847_),
    .D(_0500_));
 sg13g2_a21oi_1 _3941_ (.A1(_0447_),
    .A2(_0847_),
    .Y(_0848_),
    .B1(_0501_));
 sg13g2_nand2_1 _3942_ (.Y(_0849_),
    .A(_0485_),
    .B(_0486_));
 sg13g2_nand2_1 _3943_ (.Y(_0850_),
    .A(_0497_),
    .B(_0849_));
 sg13g2_nor2_1 _3944_ (.A(_0497_),
    .B(_0849_),
    .Y(_0851_));
 sg13g2_a21oi_1 _3945_ (.A1(_0484_),
    .A2(_0850_),
    .Y(_0852_),
    .B1(_0851_));
 sg13g2_nor2_1 _3946_ (.A(\products[5][3] ),
    .B(\products[7][3] ),
    .Y(_0853_));
 sg13g2_a21oi_1 _3947_ (.A1(\products[5][3] ),
    .A2(\products[7][3] ),
    .Y(_0854_),
    .B1(\products[6][3] ));
 sg13g2_nor2_1 _3948_ (.A(_0853_),
    .B(_0854_),
    .Y(_0855_));
 sg13g2_xnor2_1 _3949_ (.Y(_0856_),
    .A(\products[8][4] ),
    .B(\products[9][4] ));
 sg13g2_xnor2_1 _3950_ (.Y(_0857_),
    .A(_0855_),
    .B(_0856_));
 sg13g2_inv_1 _3951_ (.Y(_0858_),
    .A(_0857_));
 sg13g2_a21o_1 _3952_ (.A2(\products[9][3] ),
    .A1(\products[8][3] ),
    .B1(_0515_),
    .X(_0859_));
 sg13g2_o21ai_1 _3953_ (.B1(_0859_),
    .Y(_0860_),
    .A1(\products[8][3] ),
    .A2(\products[9][3] ));
 sg13g2_xnor2_1 _3954_ (.Y(_0861_),
    .A(_0858_),
    .B(_0860_));
 sg13g2_xnor2_1 _3955_ (.Y(_0862_),
    .A(_0852_),
    .B(_0861_));
 sg13g2_xnor2_1 _3956_ (.Y(_0863_),
    .A(_0848_),
    .B(_0862_));
 sg13g2_xnor2_1 _3957_ (.Y(_0864_),
    .A(_0846_),
    .B(_0863_));
 sg13g2_xnor2_1 _3958_ (.Y(_0865_),
    .A(_0790_),
    .B(_0864_));
 sg13g2_nand3_1 _3959_ (.B(_0504_),
    .C(_0522_),
    .A(_0503_),
    .Y(_0866_));
 sg13g2_a21oi_1 _3960_ (.A1(_0503_),
    .A2(_0504_),
    .Y(_0867_),
    .B1(_0522_));
 sg13g2_a21oi_1 _3961_ (.A1(_0508_),
    .A2(_0866_),
    .Y(_0868_),
    .B1(_0867_));
 sg13g2_xnor2_1 _3962_ (.Y(_0869_),
    .A(_0865_),
    .B(_0868_));
 sg13g2_a21oi_1 _3963_ (.A1(_0784_),
    .A2(_0785_),
    .Y(_0870_),
    .B1(_0869_));
 sg13g2_nand3_1 _3964_ (.B(_0785_),
    .C(_0869_),
    .A(_0784_),
    .Y(_0871_));
 sg13g2_nor2b_1 _3965_ (.A(_0870_),
    .B_N(_0871_),
    .Y(_0872_));
 sg13g2_xnor2_1 _3966_ (.Y(_0873_),
    .A(_0779_),
    .B(_0872_));
 sg13g2_nor2b_1 _3967_ (.A(_0767_),
    .B_N(_0562_),
    .Y(_0874_));
 sg13g2_buf_1 _3968_ (.A(_0874_),
    .X(_0875_));
 sg13g2_inv_1 _3969_ (.Y(_0876_),
    .A(_0626_));
 sg13g2_nor2_1 _3970_ (.A(_0876_),
    .B(_0875_),
    .Y(_0877_));
 sg13g2_a22oi_1 _3971_ (.Y(_0878_),
    .B1(_0877_),
    .B2(net21),
    .A2(_0875_),
    .A1(_2632_));
 sg13g2_o21ai_1 _3972_ (.B1(_0878_),
    .Y(_0109_),
    .A1(net62),
    .A2(_0873_));
 sg13g2_a21oi_1 _3973_ (.A1(_0779_),
    .A2(_0871_),
    .Y(_0879_),
    .B1(_0870_));
 sg13g2_nor2_1 _3974_ (.A(_0862_),
    .B(_0846_),
    .Y(_0880_));
 sg13g2_nand2_1 _3975_ (.Y(_0881_),
    .A(_0862_),
    .B(_0846_));
 sg13g2_o21ai_1 _3976_ (.B1(_0881_),
    .Y(_0882_),
    .A1(_0848_),
    .A2(_0880_));
 sg13g2_nor2_1 _3977_ (.A(_0818_),
    .B(_0809_),
    .Y(_0883_));
 sg13g2_nor2_1 _3978_ (.A(_0807_),
    .B(_0883_),
    .Y(_0884_));
 sg13g2_xnor2_1 _3979_ (.Y(_0885_),
    .A(\products[2][5] ),
    .B(\products[4][5] ));
 sg13g2_xnor2_1 _3980_ (.Y(_0886_),
    .A(\products[3][5] ),
    .B(_0885_));
 sg13g2_nor2_1 _3981_ (.A(\products[2][4] ),
    .B(\products[4][4] ),
    .Y(_0887_));
 sg13g2_a21oi_1 _3982_ (.A1(\products[2][4] ),
    .A2(\products[4][4] ),
    .Y(_0888_),
    .B1(\products[3][4] ));
 sg13g2_nor2_1 _3983_ (.A(_0887_),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_xnor2_1 _3984_ (.Y(_0890_),
    .A(\products[5][5] ),
    .B(\products[7][5] ));
 sg13g2_xnor2_1 _3985_ (.Y(_0891_),
    .A(\products[6][5] ),
    .B(_0890_));
 sg13g2_xor2_1 _3986_ (.B(_0891_),
    .A(_0889_),
    .X(_0892_));
 sg13g2_xnor2_1 _3987_ (.Y(_0893_),
    .A(_0886_),
    .B(_0892_));
 sg13g2_a22oi_1 _3988_ (.Y(_0894_),
    .B1(_0797_),
    .B2(_0798_),
    .A2(_0801_),
    .A1(_0800_));
 sg13g2_nand4_1 _3989_ (.B(_0801_),
    .C(_0797_),
    .A(_0800_),
    .Y(_0895_),
    .D(_0798_));
 sg13g2_o21ai_1 _3990_ (.B1(_0895_),
    .Y(_0896_),
    .A1(_0794_),
    .A2(_0894_));
 sg13g2_a21o_1 _3991_ (.A2(_0839_),
    .A1(_0834_),
    .B1(_0837_),
    .X(_0897_));
 sg13g2_o21ai_1 _3992_ (.B1(_0897_),
    .Y(_0898_),
    .A1(_0834_),
    .A2(_0839_));
 sg13g2_xnor2_1 _3993_ (.Y(_0899_),
    .A(_0896_),
    .B(_0898_));
 sg13g2_xnor2_1 _3994_ (.Y(_0900_),
    .A(_0893_),
    .B(_0899_));
 sg13g2_xnor2_1 _3995_ (.Y(_0901_),
    .A(\products[11][5] ),
    .B(\products[13][5] ));
 sg13g2_xnor2_1 _3996_ (.Y(_0902_),
    .A(\products[12][5] ),
    .B(_0901_));
 sg13g2_a21o_1 _3997_ (.A2(\products[10][4] ),
    .A1(_0814_),
    .B1(\products[0][4] ),
    .X(_0903_));
 sg13g2_o21ai_1 _3998_ (.B1(_0903_),
    .Y(_0904_),
    .A1(_0814_),
    .A2(\products[10][4] ));
 sg13g2_buf_1 _3999_ (.A(\prev_acc[5] ),
    .X(_0905_));
 sg13g2_xnor2_1 _4000_ (.Y(_0906_),
    .A(_0905_),
    .B(\products[10][5] ));
 sg13g2_xnor2_1 _4001_ (.Y(_0907_),
    .A(\products[0][5] ),
    .B(_0906_));
 sg13g2_xnor2_1 _4002_ (.Y(_0908_),
    .A(_0904_),
    .B(_0907_));
 sg13g2_xor2_1 _4003_ (.B(_0908_),
    .A(_0902_),
    .X(_0909_));
 sg13g2_nor2_1 _4004_ (.A(_0811_),
    .B(_0816_),
    .Y(_0910_));
 sg13g2_nand2_1 _4005_ (.Y(_0911_),
    .A(_0811_),
    .B(_0816_));
 sg13g2_o21ai_1 _4006_ (.B1(_0911_),
    .Y(_0912_),
    .A1(_0813_),
    .A2(_0910_));
 sg13g2_xnor2_1 _4007_ (.Y(_0913_),
    .A(\products[14][5] ),
    .B(\products[1][5] ));
 sg13g2_xnor2_1 _4008_ (.Y(_0914_),
    .A(\products[15][5] ),
    .B(_0913_));
 sg13g2_nor2_1 _4009_ (.A(\products[11][4] ),
    .B(\products[13][4] ),
    .Y(_0915_));
 sg13g2_a21oi_1 _4010_ (.A1(\products[11][4] ),
    .A2(\products[13][4] ),
    .Y(_0916_),
    .B1(\products[12][4] ));
 sg13g2_nor2_1 _4011_ (.A(_0915_),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_nor2_1 _4012_ (.A(\products[14][4] ),
    .B(\products[1][4] ),
    .Y(_0918_));
 sg13g2_a21oi_1 _4013_ (.A1(\products[14][4] ),
    .A2(\products[1][4] ),
    .Y(_0919_),
    .B1(\products[15][4] ));
 sg13g2_nor2_1 _4014_ (.A(_0918_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_xnor2_1 _4015_ (.Y(_0921_),
    .A(_0917_),
    .B(_0920_));
 sg13g2_xnor2_1 _4016_ (.Y(_0922_),
    .A(_0914_),
    .B(_0921_));
 sg13g2_xnor2_1 _4017_ (.Y(_0923_),
    .A(_0912_),
    .B(_0922_));
 sg13g2_xnor2_1 _4018_ (.Y(_0924_),
    .A(_0909_),
    .B(_0923_));
 sg13g2_xnor2_1 _4019_ (.Y(_0925_),
    .A(_0900_),
    .B(_0924_));
 sg13g2_xnor2_1 _4020_ (.Y(_0926_),
    .A(_0884_),
    .B(_0925_));
 sg13g2_a22oi_1 _4021_ (.Y(_0927_),
    .B1(_0842_),
    .B2(_0843_),
    .A2(_0821_),
    .A1(_0819_));
 sg13g2_nand4_1 _4022_ (.B(_0821_),
    .C(_0842_),
    .A(_0819_),
    .Y(_0928_),
    .D(_0843_));
 sg13g2_o21ai_1 _4023_ (.B1(_0928_),
    .Y(_0929_),
    .A1(_0823_),
    .A2(_0927_));
 sg13g2_nand2_1 _4024_ (.Y(_0930_),
    .A(_0824_),
    .B(_0825_));
 sg13g2_nor2_1 _4025_ (.A(_0841_),
    .B(_0930_),
    .Y(_0931_));
 sg13g2_nand2_1 _4026_ (.Y(_0932_),
    .A(_0841_),
    .B(_0930_));
 sg13g2_o21ai_1 _4027_ (.B1(_0932_),
    .Y(_0933_),
    .A1(_0830_),
    .A2(_0931_));
 sg13g2_nor2_1 _4028_ (.A(\products[5][4] ),
    .B(\products[7][4] ),
    .Y(_0934_));
 sg13g2_a21oi_1 _4029_ (.A1(\products[5][4] ),
    .A2(\products[7][4] ),
    .Y(_0935_),
    .B1(\products[6][4] ));
 sg13g2_nor2_1 _4030_ (.A(_0934_),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_xnor2_1 _4031_ (.Y(_0937_),
    .A(\products[8][5] ),
    .B(\products[9][5] ));
 sg13g2_xnor2_1 _4032_ (.Y(_0938_),
    .A(_0936_),
    .B(_0937_));
 sg13g2_a21o_1 _4033_ (.A2(\products[9][4] ),
    .A1(\products[8][4] ),
    .B1(_0855_),
    .X(_0939_));
 sg13g2_o21ai_1 _4034_ (.B1(_0939_),
    .Y(_0940_),
    .A1(\products[8][4] ),
    .A2(\products[9][4] ));
 sg13g2_xor2_1 _4035_ (.B(_0940_),
    .A(_0938_),
    .X(_0941_));
 sg13g2_xnor2_1 _4036_ (.Y(_0942_),
    .A(_0933_),
    .B(_0941_));
 sg13g2_xnor2_1 _4037_ (.Y(_0943_),
    .A(_0929_),
    .B(_0942_));
 sg13g2_xnor2_1 _4038_ (.Y(_0944_),
    .A(_0926_),
    .B(_0943_));
 sg13g2_inv_1 _4039_ (.Y(_0945_),
    .A(_0860_));
 sg13g2_a21oi_1 _4040_ (.A1(_0857_),
    .A2(_0945_),
    .Y(_0946_),
    .B1(_0852_));
 sg13g2_a21oi_1 _4041_ (.A1(_0858_),
    .A2(_0860_),
    .Y(_0947_),
    .B1(_0946_));
 sg13g2_xnor2_1 _4042_ (.Y(_0948_),
    .A(_0944_),
    .B(_0947_));
 sg13g2_xnor2_1 _4043_ (.Y(_0949_),
    .A(_0882_),
    .B(_0948_));
 sg13g2_xor2_1 _4044_ (.B(_0863_),
    .A(_0846_),
    .X(_0950_));
 sg13g2_a21oi_1 _4045_ (.A1(_0790_),
    .A2(_0864_),
    .Y(_0951_),
    .B1(_0868_));
 sg13g2_a21o_1 _4046_ (.A2(_0950_),
    .A1(_0789_),
    .B1(_0951_),
    .X(_0952_));
 sg13g2_nor2_1 _4047_ (.A(_0949_),
    .B(_0952_),
    .Y(_0953_));
 sg13g2_nand2_1 _4048_ (.Y(_0954_),
    .A(_0949_),
    .B(_0952_));
 sg13g2_nand2b_1 _4049_ (.Y(_0955_),
    .B(_0954_),
    .A_N(_0953_));
 sg13g2_xnor2_1 _4050_ (.Y(_0956_),
    .A(_0879_),
    .B(_0955_));
 sg13g2_a22oi_1 _4051_ (.Y(_0957_),
    .B1(_0877_),
    .B2(net22),
    .A2(_0875_),
    .A1(_2720_));
 sg13g2_o21ai_1 _4052_ (.B1(_0957_),
    .Y(_0110_),
    .A1(net62),
    .A2(_0956_));
 sg13g2_a21oi_1 _4053_ (.A1(_0879_),
    .A2(_0954_),
    .Y(_0958_),
    .B1(_0953_));
 sg13g2_and2_1 _4054_ (.A(_0944_),
    .B(_0947_),
    .X(_0959_));
 sg13g2_or2_1 _4055_ (.X(_0960_),
    .B(_0947_),
    .A(_0944_));
 sg13g2_o21ai_1 _4056_ (.B1(_0960_),
    .Y(_0961_),
    .A1(_0882_),
    .A2(_0959_));
 sg13g2_buf_1 _4057_ (.A(_0961_),
    .X(_0962_));
 sg13g2_o21ai_1 _4058_ (.B1(_0929_),
    .Y(_0963_),
    .A1(_0926_),
    .A2(_0942_));
 sg13g2_nand2_1 _4059_ (.Y(_0964_),
    .A(_0926_),
    .B(_0942_));
 sg13g2_and2_1 _4060_ (.A(_0963_),
    .B(_0964_),
    .X(_0965_));
 sg13g2_buf_1 _4061_ (.A(_0965_),
    .X(_0966_));
 sg13g2_a21o_1 _4062_ (.A2(_0922_),
    .A1(_0912_),
    .B1(_0909_),
    .X(_0967_));
 sg13g2_o21ai_1 _4063_ (.B1(_0967_),
    .Y(_0968_),
    .A1(_0912_),
    .A2(_0922_));
 sg13g2_nor2_1 _4064_ (.A(_0902_),
    .B(_0907_),
    .Y(_0969_));
 sg13g2_nand2_1 _4065_ (.Y(_0970_),
    .A(_0902_),
    .B(_0907_));
 sg13g2_o21ai_1 _4066_ (.B1(_0970_),
    .Y(_0971_),
    .A1(_0904_),
    .A2(_0969_));
 sg13g2_xnor2_1 _4067_ (.Y(_0972_),
    .A(\products[14][6] ),
    .B(\products[1][6] ));
 sg13g2_xnor2_1 _4068_ (.Y(_0973_),
    .A(\products[15][6] ),
    .B(_0972_));
 sg13g2_nor2_1 _4069_ (.A(\products[11][5] ),
    .B(\products[13][5] ),
    .Y(_0974_));
 sg13g2_a21oi_1 _4070_ (.A1(\products[11][5] ),
    .A2(\products[13][5] ),
    .Y(_0975_),
    .B1(\products[12][5] ));
 sg13g2_nor2_1 _4071_ (.A(_0974_),
    .B(_0975_),
    .Y(_0976_));
 sg13g2_nor2_1 _4072_ (.A(\products[14][5] ),
    .B(\products[1][5] ),
    .Y(_0977_));
 sg13g2_a21oi_1 _4073_ (.A1(\products[14][5] ),
    .A2(\products[1][5] ),
    .Y(_0978_),
    .B1(\products[15][5] ));
 sg13g2_nor2_1 _4074_ (.A(_0977_),
    .B(_0978_),
    .Y(_0979_));
 sg13g2_xnor2_1 _4075_ (.Y(_0980_),
    .A(_0976_),
    .B(_0979_));
 sg13g2_xor2_1 _4076_ (.B(_0980_),
    .A(_0973_),
    .X(_0981_));
 sg13g2_xnor2_1 _4077_ (.Y(_0982_),
    .A(_0971_),
    .B(_0981_));
 sg13g2_xor2_1 _4078_ (.B(\products[13][6] ),
    .A(\products[11][6] ),
    .X(_0983_));
 sg13g2_xnor2_1 _4079_ (.Y(_0984_),
    .A(\products[12][6] ),
    .B(_0983_));
 sg13g2_a21o_1 _4080_ (.A2(\products[10][5] ),
    .A1(_0905_),
    .B1(\products[0][5] ),
    .X(_0985_));
 sg13g2_o21ai_1 _4081_ (.B1(_0985_),
    .Y(_0986_),
    .A1(_0905_),
    .A2(\products[10][5] ));
 sg13g2_buf_1 _4082_ (.A(\prev_acc[6] ),
    .X(_0987_));
 sg13g2_xnor2_1 _4083_ (.Y(_0988_),
    .A(_0987_),
    .B(\products[10][6] ));
 sg13g2_xnor2_1 _4084_ (.Y(_0989_),
    .A(\products[0][6] ),
    .B(_0988_));
 sg13g2_xor2_1 _4085_ (.B(_0989_),
    .A(_0986_),
    .X(_0990_));
 sg13g2_xnor2_1 _4086_ (.Y(_0991_),
    .A(_0984_),
    .B(_0990_));
 sg13g2_xnor2_1 _4087_ (.Y(_0992_),
    .A(_0982_),
    .B(_0991_));
 sg13g2_xnor2_1 _4088_ (.Y(_0993_),
    .A(\products[5][6] ),
    .B(\products[7][6] ));
 sg13g2_xnor2_1 _4089_ (.Y(_0994_),
    .A(\products[6][6] ),
    .B(_0993_));
 sg13g2_a21o_1 _4090_ (.A2(\products[4][5] ),
    .A1(\products[2][5] ),
    .B1(\products[3][5] ),
    .X(_0995_));
 sg13g2_o21ai_1 _4091_ (.B1(_0995_),
    .Y(_0996_),
    .A1(\products[2][5] ),
    .A2(\products[4][5] ));
 sg13g2_xnor2_1 _4092_ (.Y(_0997_),
    .A(\products[2][6] ),
    .B(\products[4][6] ));
 sg13g2_xnor2_1 _4093_ (.Y(_0998_),
    .A(\products[3][6] ),
    .B(_0997_));
 sg13g2_xor2_1 _4094_ (.B(_0998_),
    .A(_0996_),
    .X(_0999_));
 sg13g2_xnor2_1 _4095_ (.Y(_1000_),
    .A(_0994_),
    .B(_0999_));
 sg13g2_a21o_1 _4096_ (.A2(_0920_),
    .A1(_0917_),
    .B1(_0914_),
    .X(_1001_));
 sg13g2_o21ai_1 _4097_ (.B1(_1001_),
    .Y(_1002_),
    .A1(_0917_),
    .A2(_0920_));
 sg13g2_nor2_1 _4098_ (.A(_0886_),
    .B(_0891_),
    .Y(_1003_));
 sg13g2_a21oi_1 _4099_ (.A1(_0886_),
    .A2(_0891_),
    .Y(_1004_),
    .B1(_0889_));
 sg13g2_nor2_1 _4100_ (.A(_1003_),
    .B(_1004_),
    .Y(_1005_));
 sg13g2_xnor2_1 _4101_ (.Y(_1006_),
    .A(_1002_),
    .B(_1005_));
 sg13g2_xnor2_1 _4102_ (.Y(_1007_),
    .A(_1000_),
    .B(_1006_));
 sg13g2_xnor2_1 _4103_ (.Y(_1008_),
    .A(_0992_),
    .B(_1007_));
 sg13g2_xnor2_1 _4104_ (.Y(_1009_),
    .A(_0968_),
    .B(_1008_));
 sg13g2_nor2b_1 _4105_ (.A(_0924_),
    .B_N(_0900_),
    .Y(_1010_));
 sg13g2_nand2b_1 _4106_ (.Y(_1011_),
    .B(_0924_),
    .A_N(_0900_));
 sg13g2_o21ai_1 _4107_ (.B1(_1011_),
    .Y(_1012_),
    .A1(_0884_),
    .A2(_1010_));
 sg13g2_nand2b_1 _4108_ (.Y(_1013_),
    .B(_0940_),
    .A_N(_0938_));
 sg13g2_nor2b_1 _4109_ (.A(_0940_),
    .B_N(_0938_),
    .Y(_1014_));
 sg13g2_a21o_1 _4110_ (.A2(_1013_),
    .A1(_0933_),
    .B1(_1014_),
    .X(_1015_));
 sg13g2_buf_1 _4111_ (.A(_1015_),
    .X(_1016_));
 sg13g2_nor2_1 _4112_ (.A(_0893_),
    .B(_0898_),
    .Y(_1017_));
 sg13g2_a21oi_1 _4113_ (.A1(_0893_),
    .A2(_0898_),
    .Y(_1018_),
    .B1(_0896_));
 sg13g2_nor2_1 _4114_ (.A(_1017_),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_nor2_1 _4115_ (.A(\products[5][5] ),
    .B(\products[7][5] ),
    .Y(_1020_));
 sg13g2_a21oi_1 _4116_ (.A1(\products[5][5] ),
    .A2(\products[7][5] ),
    .Y(_1021_),
    .B1(\products[6][5] ));
 sg13g2_nor2_1 _4117_ (.A(_1020_),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_xnor2_1 _4118_ (.Y(_1023_),
    .A(\products[8][6] ),
    .B(\products[9][6] ));
 sg13g2_xnor2_1 _4119_ (.Y(_1024_),
    .A(_1022_),
    .B(_1023_));
 sg13g2_nor2_1 _4120_ (.A(\products[8][5] ),
    .B(\products[9][5] ),
    .Y(_1025_));
 sg13g2_a21oi_1 _4121_ (.A1(\products[8][5] ),
    .A2(\products[9][5] ),
    .Y(_1026_),
    .B1(_0936_));
 sg13g2_nor2_1 _4122_ (.A(_1025_),
    .B(_1026_),
    .Y(_1027_));
 sg13g2_nor2_1 _4123_ (.A(_1024_),
    .B(_1027_),
    .Y(_1028_));
 sg13g2_nand2_1 _4124_ (.Y(_1029_),
    .A(_1024_),
    .B(_1027_));
 sg13g2_nor2b_1 _4125_ (.A(_1028_),
    .B_N(_1029_),
    .Y(_1030_));
 sg13g2_xnor2_1 _4126_ (.Y(_1031_),
    .A(_1019_),
    .B(_1030_));
 sg13g2_xnor2_1 _4127_ (.Y(_1032_),
    .A(_1016_),
    .B(_1031_));
 sg13g2_xnor2_1 _4128_ (.Y(_1033_),
    .A(_1012_),
    .B(_1032_));
 sg13g2_xnor2_1 _4129_ (.Y(_1034_),
    .A(_1009_),
    .B(_1033_));
 sg13g2_xnor2_1 _4130_ (.Y(_1035_),
    .A(_0966_),
    .B(_1034_));
 sg13g2_xor2_1 _4131_ (.B(_1035_),
    .A(_0962_),
    .X(_1036_));
 sg13g2_xnor2_1 _4132_ (.Y(_1037_),
    .A(_0958_),
    .B(_1036_));
 sg13g2_mux2_1 _4133_ (.A0(net23),
    .A1(net5),
    .S(_0875_),
    .X(_1038_));
 sg13g2_nand2_1 _4134_ (.Y(_1039_),
    .A(net62),
    .B(_1038_));
 sg13g2_o21ai_1 _4135_ (.B1(_1039_),
    .Y(_0111_),
    .A1(net62),
    .A2(_1037_));
 sg13g2_xor2_1 _4136_ (.B(_0948_),
    .A(_0882_),
    .X(_1040_));
 sg13g2_a21oi_1 _4137_ (.A1(_0789_),
    .A2(_0950_),
    .Y(_1041_),
    .B1(_0951_));
 sg13g2_o21ai_1 _4138_ (.B1(_1035_),
    .Y(_1042_),
    .A1(_1040_),
    .A2(_1041_));
 sg13g2_o21ai_1 _4139_ (.B1(_0962_),
    .Y(_1043_),
    .A1(_1040_),
    .A2(_1041_));
 sg13g2_a221oi_1 _4140_ (.B2(_1043_),
    .C1(_0870_),
    .B1(_1042_),
    .A1(_0779_),
    .Y(_1044_),
    .A2(_0871_));
 sg13g2_nand2_1 _4141_ (.Y(_1045_),
    .A(_0962_),
    .B(_1035_));
 sg13g2_o21ai_1 _4142_ (.B1(_0953_),
    .Y(_1046_),
    .A1(_0962_),
    .A2(_1035_));
 sg13g2_nand3b_1 _4143_ (.B(_1045_),
    .C(_1046_),
    .Y(_1047_),
    .A_N(_1044_));
 sg13g2_nand2b_1 _4144_ (.Y(_1048_),
    .B(_0971_),
    .A_N(_0981_));
 sg13g2_nor2_1 _4145_ (.A(_1048_),
    .B(_0984_),
    .Y(_1049_));
 sg13g2_nor2b_1 _4146_ (.A(_0971_),
    .B_N(_0981_),
    .Y(_1050_));
 sg13g2_a21oi_1 _4147_ (.A1(_1048_),
    .A2(_0984_),
    .Y(_1051_),
    .B1(_1050_));
 sg13g2_a21oi_1 _4148_ (.A1(_0989_),
    .A2(_1051_),
    .Y(_1052_),
    .B1(_1049_));
 sg13g2_nand2b_1 _4149_ (.Y(_1053_),
    .B(_1052_),
    .A_N(_0986_));
 sg13g2_nand2_1 _4150_ (.Y(_1054_),
    .A(_1050_),
    .B(_0984_));
 sg13g2_o21ai_1 _4151_ (.B1(_1054_),
    .Y(_1055_),
    .A1(_0989_),
    .A2(_1051_));
 sg13g2_nand2b_1 _4152_ (.Y(_1056_),
    .B(_0986_),
    .A_N(_1055_));
 sg13g2_nor2_1 _4153_ (.A(_0989_),
    .B(_1054_),
    .Y(_1057_));
 sg13g2_a221oi_1 _4154_ (.B2(_1056_),
    .C1(_1057_),
    .B1(_1053_),
    .A1(_0989_),
    .Y(_1058_),
    .A2(_1049_));
 sg13g2_nor2b_1 _4155_ (.A(_0992_),
    .B_N(_1007_),
    .Y(_1059_));
 sg13g2_nand2b_1 _4156_ (.Y(_1060_),
    .B(_0992_),
    .A_N(_1007_));
 sg13g2_o21ai_1 _4157_ (.B1(_1060_),
    .Y(_1061_),
    .A1(_0968_),
    .A2(_1059_));
 sg13g2_o21ai_1 _4158_ (.B1(_1029_),
    .Y(_1062_),
    .A1(_1019_),
    .A2(_1028_));
 sg13g2_xnor2_1 _4159_ (.Y(_1063_),
    .A(_1061_),
    .B(_1062_));
 sg13g2_xnor2_1 _4160_ (.Y(_1064_),
    .A(\products[14][7] ),
    .B(\products[6][7] ));
 sg13g2_a21o_1 _4161_ (.A2(\products[10][6] ),
    .A1(_0987_),
    .B1(\products[0][6] ),
    .X(_1065_));
 sg13g2_o21ai_1 _4162_ (.B1(_1065_),
    .Y(_1066_),
    .A1(_0987_),
    .A2(\products[10][6] ));
 sg13g2_xnor2_1 _4163_ (.Y(_1067_),
    .A(_1064_),
    .B(_1066_));
 sg13g2_a21o_1 _4164_ (.A2(\products[9][6] ),
    .A1(\products[8][6] ),
    .B1(_1022_),
    .X(_1068_));
 sg13g2_o21ai_1 _4165_ (.B1(_1068_),
    .Y(_1069_),
    .A1(\products[8][6] ),
    .A2(\products[9][6] ));
 sg13g2_xnor2_1 _4166_ (.Y(_1070_),
    .A(_1067_),
    .B(_1069_));
 sg13g2_xnor2_1 _4167_ (.Y(_1071_),
    .A(\products[2][7] ),
    .B(\products[4][7] ));
 sg13g2_xnor2_1 _4168_ (.Y(_1072_),
    .A(\products[1][7] ),
    .B(\products[3][7] ));
 sg13g2_xnor2_1 _4169_ (.Y(_1073_),
    .A(_1071_),
    .B(_1072_));
 sg13g2_xnor2_1 _4170_ (.Y(_1074_),
    .A(\products[15][7] ),
    .B(\products[5][7] ));
 sg13g2_xnor2_1 _4171_ (.Y(_1075_),
    .A(\products[11][7] ),
    .B(\products[13][7] ));
 sg13g2_xnor2_1 _4172_ (.Y(_1076_),
    .A(_1074_),
    .B(_1075_));
 sg13g2_xnor2_1 _4173_ (.Y(_1077_),
    .A(_1073_),
    .B(_1076_));
 sg13g2_xor2_1 _4174_ (.B(\products[12][7] ),
    .A(\products[10][7] ),
    .X(_1078_));
 sg13g2_xnor2_1 _4175_ (.Y(_1079_),
    .A(\products[0][7] ),
    .B(\prev_acc[7] ));
 sg13g2_xnor2_1 _4176_ (.Y(_1080_),
    .A(_1078_),
    .B(_1079_));
 sg13g2_xor2_1 _4177_ (.B(\products[9][7] ),
    .A(\products[8][7] ),
    .X(_1081_));
 sg13g2_xnor2_1 _4178_ (.Y(_1082_),
    .A(\products[7][7] ),
    .B(_1081_));
 sg13g2_xnor2_1 _4179_ (.Y(_1083_),
    .A(_1080_),
    .B(_1082_));
 sg13g2_xnor2_1 _4180_ (.Y(_1084_),
    .A(_1077_),
    .B(_1083_));
 sg13g2_nor2_1 _4181_ (.A(_0994_),
    .B(_0998_),
    .Y(_1085_));
 sg13g2_nand2_1 _4182_ (.Y(_1086_),
    .A(_0994_),
    .B(_0998_));
 sg13g2_o21ai_1 _4183_ (.B1(_1086_),
    .Y(_1087_),
    .A1(_0996_),
    .A2(_1085_));
 sg13g2_xnor2_1 _4184_ (.Y(_1088_),
    .A(_1084_),
    .B(_1087_));
 sg13g2_xnor2_1 _4185_ (.Y(_1089_),
    .A(_1070_),
    .B(_1088_));
 sg13g2_a21o_1 _4186_ (.A2(\products[1][6] ),
    .A1(\products[14][6] ),
    .B1(\products[15][6] ),
    .X(_1090_));
 sg13g2_o21ai_1 _4187_ (.B1(_1090_),
    .Y(_1091_),
    .A1(\products[14][6] ),
    .A2(\products[1][6] ));
 sg13g2_a21o_1 _4188_ (.A2(\products[4][6] ),
    .A1(\products[2][6] ),
    .B1(\products[3][6] ),
    .X(_1092_));
 sg13g2_o21ai_1 _4189_ (.B1(_1092_),
    .Y(_1093_),
    .A1(\products[2][6] ),
    .A2(\products[4][6] ));
 sg13g2_xor2_1 _4190_ (.B(_1093_),
    .A(_1091_),
    .X(_1094_));
 sg13g2_a21o_1 _4191_ (.A2(\products[13][6] ),
    .A1(\products[11][6] ),
    .B1(\products[12][6] ),
    .X(_1095_));
 sg13g2_o21ai_1 _4192_ (.B1(_1095_),
    .Y(_1096_),
    .A1(\products[11][6] ),
    .A2(\products[13][6] ));
 sg13g2_a21o_1 _4193_ (.A2(\products[7][6] ),
    .A1(\products[5][6] ),
    .B1(\products[6][6] ),
    .X(_1097_));
 sg13g2_o21ai_1 _4194_ (.B1(_1097_),
    .Y(_1098_),
    .A1(\products[5][6] ),
    .A2(\products[7][6] ));
 sg13g2_xor2_1 _4195_ (.B(_1098_),
    .A(_1096_),
    .X(_1099_));
 sg13g2_xnor2_1 _4196_ (.Y(_1100_),
    .A(_1094_),
    .B(_1099_));
 sg13g2_a21o_1 _4197_ (.A2(_0979_),
    .A1(_0976_),
    .B1(_0973_),
    .X(_1101_));
 sg13g2_o21ai_1 _4198_ (.B1(_1101_),
    .Y(_1102_),
    .A1(_0976_),
    .A2(_0979_));
 sg13g2_xnor2_1 _4199_ (.Y(_1103_),
    .A(_1100_),
    .B(_1102_));
 sg13g2_xnor2_1 _4200_ (.Y(_1104_),
    .A(_1089_),
    .B(_1103_));
 sg13g2_nor2_1 _4201_ (.A(_1000_),
    .B(_1005_),
    .Y(_1105_));
 sg13g2_nor2_1 _4202_ (.A(_1002_),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_a21oi_1 _4203_ (.A1(_1000_),
    .A2(_1005_),
    .Y(_1107_),
    .B1(_1106_));
 sg13g2_xnor2_1 _4204_ (.Y(_1108_),
    .A(_1104_),
    .B(_1107_));
 sg13g2_xnor2_1 _4205_ (.Y(_1109_),
    .A(_1063_),
    .B(_1108_));
 sg13g2_xnor2_1 _4206_ (.Y(_1110_),
    .A(_1058_),
    .B(_1109_));
 sg13g2_inv_1 _4207_ (.Y(_1111_),
    .A(_1012_));
 sg13g2_nor2_1 _4208_ (.A(_1009_),
    .B(_1031_),
    .Y(_1112_));
 sg13g2_nand2_1 _4209_ (.Y(_1113_),
    .A(_1009_),
    .B(_1031_));
 sg13g2_o21ai_1 _4210_ (.B1(_1113_),
    .Y(_1114_),
    .A1(_1111_),
    .A2(_1112_));
 sg13g2_nor2_1 _4211_ (.A(_1111_),
    .B(_1113_),
    .Y(_1115_));
 sg13g2_a21oi_1 _4212_ (.A1(_1016_),
    .A2(_1114_),
    .Y(_1116_),
    .B1(_1115_));
 sg13g2_nor2_1 _4213_ (.A(_0966_),
    .B(_1116_),
    .Y(_1117_));
 sg13g2_nand2_1 _4214_ (.Y(_1118_),
    .A(_1111_),
    .B(_1112_));
 sg13g2_nand2_1 _4215_ (.Y(_1119_),
    .A(_1016_),
    .B(_1115_));
 sg13g2_o21ai_1 _4216_ (.B1(_1119_),
    .Y(_1120_),
    .A1(_1016_),
    .A2(_1118_));
 sg13g2_o21ai_1 _4217_ (.B1(_1118_),
    .Y(_1121_),
    .A1(_1016_),
    .A2(_1114_));
 sg13g2_and2_1 _4218_ (.A(_0966_),
    .B(_1121_),
    .X(_1122_));
 sg13g2_nor3_1 _4219_ (.A(_1117_),
    .B(_1120_),
    .C(_1122_),
    .Y(_1123_));
 sg13g2_xnor2_1 _4220_ (.Y(_1124_),
    .A(_1110_),
    .B(_1123_));
 sg13g2_xnor2_1 _4221_ (.Y(_1125_),
    .A(_1047_),
    .B(_1124_));
 sg13g2_mux2_1 _4222_ (.A0(net24),
    .A1(net6),
    .S(_0875_),
    .X(_1126_));
 sg13g2_nand2_1 _4223_ (.Y(_1127_),
    .A(net62),
    .B(_1126_));
 sg13g2_o21ai_1 _4224_ (.B1(_1127_),
    .Y(_0112_),
    .A1(net62),
    .A2(_1125_));
 sg13g2_nor2b_1 _4225_ (.A(_0767_),
    .B_N(_0576_),
    .Y(_1128_));
 sg13g2_buf_1 _4226_ (.A(_1128_),
    .X(_1129_));
 sg13g2_mux2_1 _4227_ (.A0(\mem[35][0] ),
    .A1(net50),
    .S(_1129_),
    .X(_0113_));
 sg13g2_mux2_1 _4228_ (.A0(\mem[35][1] ),
    .A1(net43),
    .S(_1129_),
    .X(_0114_));
 sg13g2_mux2_1 _4229_ (.A0(\mem[35][2] ),
    .A1(net35),
    .S(_1129_),
    .X(_0115_));
 sg13g2_mux2_1 _4230_ (.A0(\mem[35][3] ),
    .A1(_0663_),
    .S(_1129_),
    .X(_0116_));
 sg13g2_nor2b_1 _4231_ (.A(_0767_),
    .B_N(_0589_),
    .Y(_1130_));
 sg13g2_buf_1 _4232_ (.A(_1130_),
    .X(_1131_));
 sg13g2_mux2_1 _4233_ (.A0(\mem[36][0] ),
    .A1(net50),
    .S(_1131_),
    .X(_0117_));
 sg13g2_mux2_1 _4234_ (.A0(\mem[36][1] ),
    .A1(net43),
    .S(_1131_),
    .X(_0118_));
 sg13g2_mux2_1 _4235_ (.A0(\mem[36][2] ),
    .A1(_0661_),
    .S(_1131_),
    .X(_0119_));
 sg13g2_mux2_1 _4236_ (.A0(\mem[36][3] ),
    .A1(_0663_),
    .S(_1131_),
    .X(_0120_));
 sg13g2_nor3_2 _4237_ (.A(_0587_),
    .B(_0595_),
    .C(_0767_),
    .Y(_1132_));
 sg13g2_mux2_1 _4238_ (.A0(\mem[37][0] ),
    .A1(_0655_),
    .S(_1132_),
    .X(_0121_));
 sg13g2_mux2_1 _4239_ (.A0(\mem[37][1] ),
    .A1(net43),
    .S(_1132_),
    .X(_0122_));
 sg13g2_mux2_1 _4240_ (.A0(\mem[37][2] ),
    .A1(net38),
    .S(_1132_),
    .X(_0123_));
 sg13g2_mux2_1 _4241_ (.A0(\mem[37][3] ),
    .A1(net31),
    .S(_1132_),
    .X(_0124_));
 sg13g2_nor2b_1 _4242_ (.A(_0767_),
    .B_N(_0604_),
    .Y(_1133_));
 sg13g2_buf_2 _4243_ (.A(_1133_),
    .X(_1134_));
 sg13g2_mux2_1 _4244_ (.A0(\mem[38][0] ),
    .A1(_0655_),
    .S(_1134_),
    .X(_0125_));
 sg13g2_mux2_1 _4245_ (.A0(\mem[38][1] ),
    .A1(net43),
    .S(_1134_),
    .X(_0126_));
 sg13g2_mux2_1 _4246_ (.A0(\mem[38][2] ),
    .A1(net38),
    .S(_1134_),
    .X(_0127_));
 sg13g2_mux2_1 _4247_ (.A0(\mem[38][3] ),
    .A1(_0555_),
    .S(_1134_),
    .X(_0128_));
 sg13g2_nor2b_1 _4248_ (.A(_0767_),
    .B_N(_0611_),
    .Y(_1135_));
 sg13g2_buf_1 _4249_ (.A(_1135_),
    .X(_1136_));
 sg13g2_mux2_1 _4250_ (.A0(\mem[39][0] ),
    .A1(net52),
    .S(_1136_),
    .X(_0129_));
 sg13g2_mux2_1 _4251_ (.A0(\mem[39][1] ),
    .A1(net43),
    .S(_1136_),
    .X(_0130_));
 sg13g2_mux2_1 _4252_ (.A0(\mem[39][2] ),
    .A1(net38),
    .S(_1136_),
    .X(_0131_));
 sg13g2_mux2_1 _4253_ (.A0(\mem[39][3] ),
    .A1(net31),
    .S(_1136_),
    .X(_0132_));
 sg13g2_buf_1 _4254_ (.A(\mem[3][0] ),
    .X(_1137_));
 sg13g2_nand2_2 _4255_ (.Y(_1138_),
    .A(_2644_),
    .B(_0576_));
 sg13g2_mux2_1 _4256_ (.A0(net48),
    .A1(net100),
    .S(_1138_),
    .X(_0133_));
 sg13g2_buf_2 _4257_ (.A(\mem[3][1] ),
    .X(_1139_));
 sg13g2_mux2_1 _4258_ (.A0(_2721_),
    .A1(_1139_),
    .S(_1138_),
    .X(_0134_));
 sg13g2_buf_1 _4259_ (.A(\mem[3][2] ),
    .X(_1140_));
 sg13g2_mux2_1 _4260_ (.A0(net34),
    .A1(_1140_),
    .S(_1138_),
    .X(_0135_));
 sg13g2_buf_2 _4261_ (.A(\mem[3][3] ),
    .X(_1141_));
 sg13g2_mux2_1 _4262_ (.A0(net27),
    .A1(_1141_),
    .S(_1138_),
    .X(_0136_));
 sg13g2_nand2_1 _4263_ (.Y(_1142_),
    .A(_2642_),
    .B(_2647_));
 sg13g2_nor2_1 _4264_ (.A(_0564_),
    .B(_1142_),
    .Y(_1143_));
 sg13g2_buf_4 _4265_ (.X(_1144_),
    .A(_1143_));
 sg13g2_nand2_2 _4266_ (.Y(_1145_),
    .A(_2639_),
    .B(_1144_));
 sg13g2_mux2_1 _4267_ (.A0(net48),
    .A1(\mem[40][0] ),
    .S(_1145_),
    .X(_0137_));
 sg13g2_buf_1 _4268_ (.A(net45),
    .X(_1146_));
 sg13g2_mux2_1 _4269_ (.A0(net41),
    .A1(\mem[40][1] ),
    .S(_1145_),
    .X(_0138_));
 sg13g2_mux2_1 _4270_ (.A0(net34),
    .A1(\mem[40][2] ),
    .S(_1145_),
    .X(_0139_));
 sg13g2_mux2_1 _4271_ (.A0(net27),
    .A1(\mem[40][3] ),
    .S(_1145_),
    .X(_0140_));
 sg13g2_nand2_2 _4272_ (.Y(_1147_),
    .A(_0629_),
    .B(_1144_));
 sg13g2_mux2_1 _4273_ (.A0(net48),
    .A1(\mem[41][0] ),
    .S(_1147_),
    .X(_0141_));
 sg13g2_mux2_1 _4274_ (.A0(net41),
    .A1(\mem[41][1] ),
    .S(_1147_),
    .X(_0142_));
 sg13g2_mux2_1 _4275_ (.A0(net34),
    .A1(\mem[41][2] ),
    .S(_1147_),
    .X(_0143_));
 sg13g2_mux2_1 _4276_ (.A0(net27),
    .A1(\mem[41][3] ),
    .S(_1147_),
    .X(_0144_));
 sg13g2_nand2_2 _4277_ (.Y(_1148_),
    .A(_0562_),
    .B(_1144_));
 sg13g2_mux2_1 _4278_ (.A0(net48),
    .A1(\mem[42][0] ),
    .S(_1148_),
    .X(_0145_));
 sg13g2_mux2_1 _4279_ (.A0(_1146_),
    .A1(\mem[42][1] ),
    .S(_1148_),
    .X(_0146_));
 sg13g2_mux2_1 _4280_ (.A0(net34),
    .A1(\mem[42][2] ),
    .S(_1148_),
    .X(_0147_));
 sg13g2_mux2_1 _4281_ (.A0(net27),
    .A1(\mem[42][3] ),
    .S(_1148_),
    .X(_0148_));
 sg13g2_nand2_2 _4282_ (.Y(_1149_),
    .A(_0576_),
    .B(_1144_));
 sg13g2_mux2_1 _4283_ (.A0(net48),
    .A1(\mem[43][0] ),
    .S(_1149_),
    .X(_0149_));
 sg13g2_mux2_1 _4284_ (.A0(net41),
    .A1(\mem[43][1] ),
    .S(_1149_),
    .X(_0150_));
 sg13g2_mux2_1 _4285_ (.A0(net34),
    .A1(\mem[43][2] ),
    .S(_1149_),
    .X(_0151_));
 sg13g2_mux2_1 _4286_ (.A0(net27),
    .A1(\mem[43][3] ),
    .S(_1149_),
    .X(_0152_));
 sg13g2_nand2_2 _4287_ (.Y(_1150_),
    .A(_0589_),
    .B(_1144_));
 sg13g2_mux2_1 _4288_ (.A0(net48),
    .A1(\mem[44][0] ),
    .S(_1150_),
    .X(_0153_));
 sg13g2_mux2_1 _4289_ (.A0(_1146_),
    .A1(\mem[44][1] ),
    .S(_1150_),
    .X(_0154_));
 sg13g2_mux2_1 _4290_ (.A0(net34),
    .A1(\mem[44][2] ),
    .S(_1150_),
    .X(_0155_));
 sg13g2_mux2_1 _4291_ (.A0(net27),
    .A1(\mem[44][3] ),
    .S(_1150_),
    .X(_0156_));
 sg13g2_nand2_2 _4292_ (.Y(_1151_),
    .A(_0597_),
    .B(_1144_));
 sg13g2_mux2_1 _4293_ (.A0(net48),
    .A1(\mem[45][0] ),
    .S(_1151_),
    .X(_0157_));
 sg13g2_mux2_1 _4294_ (.A0(net41),
    .A1(\mem[45][1] ),
    .S(_1151_),
    .X(_0158_));
 sg13g2_buf_1 _4295_ (.A(net38),
    .X(_1152_));
 sg13g2_mux2_1 _4296_ (.A0(net33),
    .A1(\mem[45][2] ),
    .S(_1151_),
    .X(_0159_));
 sg13g2_buf_8 _4297_ (.A(net31),
    .X(_1153_));
 sg13g2_mux2_1 _4298_ (.A0(net26),
    .A1(\mem[45][3] ),
    .S(_1151_),
    .X(_0160_));
 sg13g2_nand2_2 _4299_ (.Y(_1154_),
    .A(_0604_),
    .B(_1144_));
 sg13g2_mux2_1 _4300_ (.A0(net48),
    .A1(\mem[46][0] ),
    .S(_1154_),
    .X(_0161_));
 sg13g2_mux2_1 _4301_ (.A0(net41),
    .A1(\mem[46][1] ),
    .S(_1154_),
    .X(_0162_));
 sg13g2_mux2_1 _4302_ (.A0(net33),
    .A1(\mem[46][2] ),
    .S(_1154_),
    .X(_0163_));
 sg13g2_mux2_1 _4303_ (.A0(net26),
    .A1(\mem[46][3] ),
    .S(_1154_),
    .X(_0164_));
 sg13g2_buf_1 _4304_ (.A(net52),
    .X(_1155_));
 sg13g2_nand2_2 _4305_ (.Y(_1156_),
    .A(_0611_),
    .B(_1144_));
 sg13g2_mux2_1 _4306_ (.A0(net47),
    .A1(\mem[47][0] ),
    .S(_1156_),
    .X(_0165_));
 sg13g2_mux2_1 _4307_ (.A0(net41),
    .A1(\mem[47][1] ),
    .S(_1156_),
    .X(_0166_));
 sg13g2_mux2_1 _4308_ (.A0(net33),
    .A1(\mem[47][2] ),
    .S(_1156_),
    .X(_0167_));
 sg13g2_mux2_1 _4309_ (.A0(net26),
    .A1(\mem[47][3] ),
    .S(_1156_),
    .X(_0168_));
 sg13g2_nor2_1 _4310_ (.A(_0617_),
    .B(_1142_),
    .Y(_1157_));
 sg13g2_buf_4 _4311_ (.X(_1158_),
    .A(_1157_));
 sg13g2_nand2_2 _4312_ (.Y(_1159_),
    .A(_2639_),
    .B(_1158_));
 sg13g2_mux2_1 _4313_ (.A0(net47),
    .A1(\mem[48][0] ),
    .S(_1159_),
    .X(_0169_));
 sg13g2_mux2_1 _4314_ (.A0(net41),
    .A1(\mem[48][1] ),
    .S(_1159_),
    .X(_0170_));
 sg13g2_mux2_1 _4315_ (.A0(net33),
    .A1(\mem[48][2] ),
    .S(_1159_),
    .X(_0171_));
 sg13g2_mux2_1 _4316_ (.A0(net26),
    .A1(\mem[48][3] ),
    .S(_1159_),
    .X(_0172_));
 sg13g2_nand2_2 _4317_ (.Y(_1160_),
    .A(_0629_),
    .B(_1158_));
 sg13g2_mux2_1 _4318_ (.A0(net47),
    .A1(\mem[49][0] ),
    .S(_1160_),
    .X(_0173_));
 sg13g2_mux2_1 _4319_ (.A0(net41),
    .A1(\mem[49][1] ),
    .S(_1160_),
    .X(_0174_));
 sg13g2_mux2_1 _4320_ (.A0(net33),
    .A1(\mem[49][2] ),
    .S(_1160_),
    .X(_0175_));
 sg13g2_mux2_1 _4321_ (.A0(net26),
    .A1(\mem[49][3] ),
    .S(_1160_),
    .X(_0176_));
 sg13g2_buf_1 _4322_ (.A(\mem[4][0] ),
    .X(_1161_));
 sg13g2_nand2_2 _4323_ (.Y(_1162_),
    .A(_2644_),
    .B(_0589_));
 sg13g2_mux2_1 _4324_ (.A0(net47),
    .A1(net98),
    .S(_1162_),
    .X(_0177_));
 sg13g2_buf_1 _4325_ (.A(net45),
    .X(_1163_));
 sg13g2_buf_2 _4326_ (.A(\mem[4][1] ),
    .X(_1164_));
 sg13g2_mux2_1 _4327_ (.A0(net40),
    .A1(_1164_),
    .S(_1162_),
    .X(_0178_));
 sg13g2_buf_1 _4328_ (.A(\mem[4][2] ),
    .X(_1165_));
 sg13g2_mux2_1 _4329_ (.A0(net33),
    .A1(_1165_),
    .S(_1162_),
    .X(_0179_));
 sg13g2_buf_2 _4330_ (.A(\mem[4][3] ),
    .X(_1166_));
 sg13g2_mux2_1 _4331_ (.A0(net26),
    .A1(_1166_),
    .S(_1162_),
    .X(_0180_));
 sg13g2_nand2_2 _4332_ (.Y(_1167_),
    .A(_0562_),
    .B(_1158_));
 sg13g2_mux2_1 _4333_ (.A0(_1155_),
    .A1(\mem[50][0] ),
    .S(_1167_),
    .X(_0181_));
 sg13g2_mux2_1 _4334_ (.A0(net40),
    .A1(\mem[50][1] ),
    .S(_1167_),
    .X(_0182_));
 sg13g2_mux2_1 _4335_ (.A0(_1152_),
    .A1(\mem[50][2] ),
    .S(_1167_),
    .X(_0183_));
 sg13g2_mux2_1 _4336_ (.A0(_1153_),
    .A1(\mem[50][3] ),
    .S(_1167_),
    .X(_0184_));
 sg13g2_nand2_2 _4337_ (.Y(_1168_),
    .A(_0576_),
    .B(_1158_));
 sg13g2_mux2_1 _4338_ (.A0(_1155_),
    .A1(\mem[51][0] ),
    .S(_1168_),
    .X(_0185_));
 sg13g2_mux2_1 _4339_ (.A0(_1163_),
    .A1(\mem[51][1] ),
    .S(_1168_),
    .X(_0186_));
 sg13g2_mux2_1 _4340_ (.A0(_1152_),
    .A1(\mem[51][2] ),
    .S(_1168_),
    .X(_0187_));
 sg13g2_mux2_1 _4341_ (.A0(_1153_),
    .A1(\mem[51][3] ),
    .S(_1168_),
    .X(_0188_));
 sg13g2_nand2_2 _4342_ (.Y(_1169_),
    .A(_0589_),
    .B(_1158_));
 sg13g2_mux2_1 _4343_ (.A0(net47),
    .A1(\mem[52][0] ),
    .S(_1169_),
    .X(_0189_));
 sg13g2_mux2_1 _4344_ (.A0(net40),
    .A1(\mem[52][1] ),
    .S(_1169_),
    .X(_0190_));
 sg13g2_mux2_1 _4345_ (.A0(net33),
    .A1(\mem[52][2] ),
    .S(_1169_),
    .X(_0191_));
 sg13g2_mux2_1 _4346_ (.A0(net26),
    .A1(\mem[52][3] ),
    .S(_1169_),
    .X(_0192_));
 sg13g2_nand2_2 _4347_ (.Y(_1170_),
    .A(_0597_),
    .B(_1158_));
 sg13g2_mux2_1 _4348_ (.A0(net47),
    .A1(\mem[53][0] ),
    .S(_1170_),
    .X(_0193_));
 sg13g2_mux2_1 _4349_ (.A0(net40),
    .A1(\mem[53][1] ),
    .S(_1170_),
    .X(_0194_));
 sg13g2_mux2_1 _4350_ (.A0(net33),
    .A1(\mem[53][2] ),
    .S(_1170_),
    .X(_0195_));
 sg13g2_mux2_1 _4351_ (.A0(net26),
    .A1(\mem[53][3] ),
    .S(_1170_),
    .X(_0196_));
 sg13g2_nand2_2 _4352_ (.Y(_1171_),
    .A(_0604_),
    .B(_1158_));
 sg13g2_mux2_1 _4353_ (.A0(net47),
    .A1(\mem[54][0] ),
    .S(_1171_),
    .X(_0197_));
 sg13g2_mux2_1 _4354_ (.A0(_1163_),
    .A1(\mem[54][1] ),
    .S(_1171_),
    .X(_0198_));
 sg13g2_buf_1 _4355_ (.A(net38),
    .X(_1172_));
 sg13g2_mux2_1 _4356_ (.A0(net32),
    .A1(\mem[54][2] ),
    .S(_1171_),
    .X(_0199_));
 sg13g2_buf_8 _4357_ (.A(net31),
    .X(_1173_));
 sg13g2_mux2_1 _4358_ (.A0(net25),
    .A1(\mem[54][3] ),
    .S(_1171_),
    .X(_0200_));
 sg13g2_nand2_2 _4359_ (.Y(_1174_),
    .A(_0611_),
    .B(_1158_));
 sg13g2_mux2_1 _4360_ (.A0(net47),
    .A1(\mem[55][0] ),
    .S(_1174_),
    .X(_0201_));
 sg13g2_mux2_1 _4361_ (.A0(net40),
    .A1(\mem[55][1] ),
    .S(_1174_),
    .X(_0202_));
 sg13g2_mux2_1 _4362_ (.A0(net32),
    .A1(\mem[55][2] ),
    .S(_1174_),
    .X(_0203_));
 sg13g2_mux2_1 _4363_ (.A0(net25),
    .A1(\mem[55][3] ),
    .S(_1174_),
    .X(_0204_));
 sg13g2_buf_1 _4364_ (.A(net52),
    .X(_1175_));
 sg13g2_nor2_1 _4365_ (.A(_0694_),
    .B(_1142_),
    .Y(_1176_));
 sg13g2_buf_4 _4366_ (.X(_1177_),
    .A(_1176_));
 sg13g2_nand2_2 _4367_ (.Y(_1178_),
    .A(_2639_),
    .B(_1177_));
 sg13g2_mux2_1 _4368_ (.A0(net46),
    .A1(\mem[56][0] ),
    .S(_1178_),
    .X(_0205_));
 sg13g2_mux2_1 _4369_ (.A0(net40),
    .A1(\mem[56][1] ),
    .S(_1178_),
    .X(_0206_));
 sg13g2_mux2_1 _4370_ (.A0(net32),
    .A1(\mem[56][2] ),
    .S(_1178_),
    .X(_0207_));
 sg13g2_mux2_1 _4371_ (.A0(net25),
    .A1(\mem[56][3] ),
    .S(_1178_),
    .X(_0208_));
 sg13g2_nand2_2 _4372_ (.Y(_1179_),
    .A(_0629_),
    .B(_1177_));
 sg13g2_mux2_1 _4373_ (.A0(net46),
    .A1(\mem[57][0] ),
    .S(_1179_),
    .X(_0209_));
 sg13g2_mux2_1 _4374_ (.A0(net40),
    .A1(\mem[57][1] ),
    .S(_1179_),
    .X(_0210_));
 sg13g2_mux2_1 _4375_ (.A0(net32),
    .A1(\mem[57][2] ),
    .S(_1179_),
    .X(_0211_));
 sg13g2_mux2_1 _4376_ (.A0(net25),
    .A1(\mem[57][3] ),
    .S(_1179_),
    .X(_0212_));
 sg13g2_nand2_2 _4377_ (.Y(_1180_),
    .A(_0562_),
    .B(_1177_));
 sg13g2_mux2_1 _4378_ (.A0(net46),
    .A1(\mem[58][0] ),
    .S(_1180_),
    .X(_0213_));
 sg13g2_mux2_1 _4379_ (.A0(net40),
    .A1(\mem[58][1] ),
    .S(_1180_),
    .X(_0214_));
 sg13g2_mux2_1 _4380_ (.A0(net32),
    .A1(\mem[58][2] ),
    .S(_1180_),
    .X(_0215_));
 sg13g2_mux2_1 _4381_ (.A0(net25),
    .A1(\mem[58][3] ),
    .S(_1180_),
    .X(_0216_));
 sg13g2_nand2_2 _4382_ (.Y(_1181_),
    .A(_0576_),
    .B(_1177_));
 sg13g2_mux2_1 _4383_ (.A0(net46),
    .A1(\mem[59][0] ),
    .S(_1181_),
    .X(_0217_));
 sg13g2_buf_1 _4384_ (.A(net45),
    .X(_1182_));
 sg13g2_mux2_1 _4385_ (.A0(net39),
    .A1(\mem[59][1] ),
    .S(_1181_),
    .X(_0218_));
 sg13g2_mux2_1 _4386_ (.A0(net32),
    .A1(\mem[59][2] ),
    .S(_1181_),
    .X(_0219_));
 sg13g2_mux2_1 _4387_ (.A0(net25),
    .A1(\mem[59][3] ),
    .S(_1181_),
    .X(_0220_));
 sg13g2_buf_1 _4388_ (.A(\mem[5][0] ),
    .X(_1183_));
 sg13g2_nand2_2 _4389_ (.Y(_1184_),
    .A(_2644_),
    .B(_0597_));
 sg13g2_mux2_1 _4390_ (.A0(_1175_),
    .A1(net96),
    .S(_1184_),
    .X(_0221_));
 sg13g2_buf_2 _4391_ (.A(\mem[5][1] ),
    .X(_1185_));
 sg13g2_mux2_1 _4392_ (.A0(_1182_),
    .A1(_1185_),
    .S(_1184_),
    .X(_0222_));
 sg13g2_buf_1 _4393_ (.A(\mem[5][2] ),
    .X(_1186_));
 sg13g2_mux2_1 _4394_ (.A0(net32),
    .A1(_1186_),
    .S(_1184_),
    .X(_0223_));
 sg13g2_buf_2 _4395_ (.A(\mem[5][3] ),
    .X(_1187_));
 sg13g2_mux2_1 _4396_ (.A0(net25),
    .A1(_1187_),
    .S(_1184_),
    .X(_0224_));
 sg13g2_nand2_2 _4397_ (.Y(_1188_),
    .A(_0589_),
    .B(_1177_));
 sg13g2_mux2_1 _4398_ (.A0(net46),
    .A1(\mem[60][0] ),
    .S(_1188_),
    .X(_0225_));
 sg13g2_mux2_1 _4399_ (.A0(net39),
    .A1(\mem[60][1] ),
    .S(_1188_),
    .X(_0226_));
 sg13g2_mux2_1 _4400_ (.A0(net32),
    .A1(\mem[60][2] ),
    .S(_1188_),
    .X(_0227_));
 sg13g2_mux2_1 _4401_ (.A0(net25),
    .A1(\mem[60][3] ),
    .S(_1188_),
    .X(_0228_));
 sg13g2_nand2_2 _4402_ (.Y(_1189_),
    .A(_0597_),
    .B(_1177_));
 sg13g2_mux2_1 _4403_ (.A0(net46),
    .A1(\mem[61][0] ),
    .S(_1189_),
    .X(_0229_));
 sg13g2_mux2_1 _4404_ (.A0(net39),
    .A1(\mem[61][1] ),
    .S(_1189_),
    .X(_0230_));
 sg13g2_mux2_1 _4405_ (.A0(_1172_),
    .A1(\mem[61][2] ),
    .S(_1189_),
    .X(_0231_));
 sg13g2_mux2_1 _4406_ (.A0(_1173_),
    .A1(\mem[61][3] ),
    .S(_1189_),
    .X(_0232_));
 sg13g2_nand2_2 _4407_ (.Y(_1190_),
    .A(_0604_),
    .B(_1177_));
 sg13g2_mux2_1 _4408_ (.A0(net46),
    .A1(\mem[62][0] ),
    .S(_1190_),
    .X(_0233_));
 sg13g2_mux2_1 _4409_ (.A0(net39),
    .A1(\mem[62][1] ),
    .S(_1190_),
    .X(_0234_));
 sg13g2_mux2_1 _4410_ (.A0(_1172_),
    .A1(\mem[62][2] ),
    .S(_1190_),
    .X(_0235_));
 sg13g2_mux2_1 _4411_ (.A0(_1173_),
    .A1(\mem[62][3] ),
    .S(_1190_),
    .X(_0236_));
 sg13g2_nand2_2 _4412_ (.Y(_1191_),
    .A(_0611_),
    .B(_1177_));
 sg13g2_mux2_1 _4413_ (.A0(net46),
    .A1(\mem[63][0] ),
    .S(_1191_),
    .X(_0237_));
 sg13g2_mux2_1 _4414_ (.A0(net39),
    .A1(\mem[63][1] ),
    .S(_1191_),
    .X(_0238_));
 sg13g2_mux2_1 _4415_ (.A0(_0661_),
    .A1(\mem[63][2] ),
    .S(_1191_),
    .X(_0239_));
 sg13g2_mux2_1 _4416_ (.A0(net28),
    .A1(\mem[63][3] ),
    .S(_1191_),
    .X(_0240_));
 sg13g2_buf_1 _4417_ (.A(\mem[6][0] ),
    .X(_1192_));
 sg13g2_nand2_2 _4418_ (.Y(_1193_),
    .A(_2644_),
    .B(_0604_));
 sg13g2_mux2_1 _4419_ (.A0(_1175_),
    .A1(net94),
    .S(_1193_),
    .X(_0241_));
 sg13g2_buf_2 _4420_ (.A(\mem[6][1] ),
    .X(_1194_));
 sg13g2_mux2_1 _4421_ (.A0(net39),
    .A1(_1194_),
    .S(_1193_),
    .X(_0242_));
 sg13g2_buf_1 _4422_ (.A(\mem[6][2] ),
    .X(_1195_));
 sg13g2_mux2_1 _4423_ (.A0(net35),
    .A1(net93),
    .S(_1193_),
    .X(_0243_));
 sg13g2_buf_2 _4424_ (.A(\mem[6][3] ),
    .X(_1196_));
 sg13g2_mux2_1 _4425_ (.A0(net28),
    .A1(_1196_),
    .S(_1193_),
    .X(_0244_));
 sg13g2_buf_1 _4426_ (.A(\mem[7][0] ),
    .X(_1197_));
 sg13g2_nand2_2 _4427_ (.Y(_1198_),
    .A(_2644_),
    .B(_0611_));
 sg13g2_mux2_1 _4428_ (.A0(net50),
    .A1(net92),
    .S(_1198_),
    .X(_0245_));
 sg13g2_buf_2 _4429_ (.A(\mem[7][1] ),
    .X(_1199_));
 sg13g2_mux2_1 _4430_ (.A0(_1182_),
    .A1(_1199_),
    .S(_1198_),
    .X(_0246_));
 sg13g2_buf_1 _4431_ (.A(\mem[7][2] ),
    .X(_1200_));
 sg13g2_mux2_1 _4432_ (.A0(net35),
    .A1(net91),
    .S(_1198_),
    .X(_0247_));
 sg13g2_buf_2 _4433_ (.A(\mem[7][3] ),
    .X(_1201_));
 sg13g2_mux2_1 _4434_ (.A0(net28),
    .A1(_1201_),
    .S(_1198_),
    .X(_0248_));
 sg13g2_buf_1 _4435_ (.A(\mem[8][0] ),
    .X(_1202_));
 sg13g2_nand2_2 _4436_ (.Y(_1203_),
    .A(_2639_),
    .B(_0566_));
 sg13g2_mux2_1 _4437_ (.A0(net50),
    .A1(net90),
    .S(_1203_),
    .X(_0249_));
 sg13g2_buf_2 _4438_ (.A(\mem[8][1] ),
    .X(_1204_));
 sg13g2_mux2_1 _4439_ (.A0(net39),
    .A1(_1204_),
    .S(_1203_),
    .X(_0250_));
 sg13g2_buf_1 _4440_ (.A(\mem[8][2] ),
    .X(_1205_));
 sg13g2_mux2_1 _4441_ (.A0(net35),
    .A1(net89),
    .S(_1203_),
    .X(_0251_));
 sg13g2_buf_2 _4442_ (.A(\mem[8][3] ),
    .X(_1206_));
 sg13g2_mux2_1 _4443_ (.A0(net28),
    .A1(_1206_),
    .S(_1203_),
    .X(_0252_));
 sg13g2_buf_1 _4444_ (.A(\mem[9][0] ),
    .X(_1207_));
 sg13g2_nand2_2 _4445_ (.Y(_1208_),
    .A(_0566_),
    .B(_0629_));
 sg13g2_mux2_1 _4446_ (.A0(net50),
    .A1(net88),
    .S(_1208_),
    .X(_0253_));
 sg13g2_buf_1 _4447_ (.A(\mem[9][1] ),
    .X(_1209_));
 sg13g2_mux2_1 _4448_ (.A0(net39),
    .A1(_1209_),
    .S(_1208_),
    .X(_0254_));
 sg13g2_buf_1 _4449_ (.A(\mem[9][2] ),
    .X(_1210_));
 sg13g2_mux2_1 _4450_ (.A0(net35),
    .A1(net87),
    .S(_1208_),
    .X(_0255_));
 sg13g2_buf_2 _4451_ (.A(\mem[9][3] ),
    .X(_1211_));
 sg13g2_mux2_1 _4452_ (.A0(net28),
    .A1(_1211_),
    .S(_1208_),
    .X(_0256_));
 sg13g2_o21ai_1 _4453_ (.B1(_2606_),
    .Y(_1212_),
    .A1(_2607_),
    .A2(_2608_));
 sg13g2_inv_1 _4454_ (.Y(_0394_),
    .A(_1212_));
 sg13g2_nor2b_1 _4455_ (.A(_2608_),
    .B_N(_2607_),
    .Y(_1213_));
 sg13g2_buf_1 _4456_ (.A(_1213_),
    .X(_1214_));
 sg13g2_buf_1 _4457_ (.A(net61),
    .X(_1215_));
 sg13g2_nand2_1 _4458_ (.Y(_1216_),
    .A(net17),
    .B(net59));
 sg13g2_nand2b_1 _4459_ (.Y(_1217_),
    .B(_2618_),
    .A_N(net59));
 sg13g2_inv_1 _4460_ (.Y(_1218_),
    .A(_2606_));
 sg13g2_a21oi_1 _4461_ (.A1(_1216_),
    .A2(_1217_),
    .Y(_0257_),
    .B1(net86));
 sg13g2_nand2_1 _4462_ (.Y(_1219_),
    .A(net18),
    .B(net59));
 sg13g2_nand2b_1 _4463_ (.Y(_1220_),
    .B(_2665_),
    .A_N(net59));
 sg13g2_a21oi_1 _4464_ (.A1(_1219_),
    .A2(_1220_),
    .Y(_0258_),
    .B1(net86));
 sg13g2_nand2_1 _4465_ (.Y(_1221_),
    .A(net19),
    .B(net59));
 sg13g2_nand2b_1 _4466_ (.Y(_1222_),
    .B(_2756_),
    .A_N(net61));
 sg13g2_a21oi_1 _4467_ (.A1(_1221_),
    .A2(_1222_),
    .Y(_0259_),
    .B1(net86));
 sg13g2_nand2_1 _4468_ (.Y(_1223_),
    .A(net20),
    .B(net59));
 sg13g2_nand2b_1 _4469_ (.Y(_1224_),
    .B(_0473_),
    .A_N(net61));
 sg13g2_a21oi_1 _4470_ (.A1(_1223_),
    .A2(_1224_),
    .Y(_0260_),
    .B1(net86));
 sg13g2_nand2_1 _4471_ (.Y(_1225_),
    .A(net21),
    .B(net59));
 sg13g2_nand2b_1 _4472_ (.Y(_1226_),
    .B(_0814_),
    .A_N(net61));
 sg13g2_a21oi_1 _4473_ (.A1(_1225_),
    .A2(_1226_),
    .Y(_0261_),
    .B1(net86));
 sg13g2_nand2_1 _4474_ (.Y(_1227_),
    .A(net22),
    .B(_1215_));
 sg13g2_nand2b_1 _4475_ (.Y(_1228_),
    .B(_0905_),
    .A_N(net61));
 sg13g2_a21oi_1 _4476_ (.A1(_1227_),
    .A2(_1228_),
    .Y(_0262_),
    .B1(net86));
 sg13g2_nand2_1 _4477_ (.Y(_1229_),
    .A(net23),
    .B(_1215_));
 sg13g2_nand2b_1 _4478_ (.Y(_1230_),
    .B(_0987_),
    .A_N(_1214_));
 sg13g2_a21oi_1 _4479_ (.A1(_1229_),
    .A2(_1230_),
    .Y(_0263_),
    .B1(_1218_));
 sg13g2_nand2_1 _4480_ (.Y(_1231_),
    .A(net24),
    .B(net59));
 sg13g2_nand2b_1 _4481_ (.Y(_1232_),
    .B(\prev_acc[7] ),
    .A_N(net61));
 sg13g2_a21oi_1 _4482_ (.A1(_1231_),
    .A2(_1232_),
    .Y(_0264_),
    .B1(net86));
 sg13g2_nand2_1 _4483_ (.Y(_1233_),
    .A(_2606_),
    .B(net61));
 sg13g2_buf_2 _4484_ (.A(_1233_),
    .X(_1234_));
 sg13g2_nand2_1 _4485_ (.Y(_1235_),
    .A(net144),
    .B(net156));
 sg13g2_nor2_1 _4486_ (.A(_1234_),
    .B(_1235_),
    .Y(_0265_));
 sg13g2_nand2_1 _4487_ (.Y(_1236_),
    .A(net144),
    .B(net155));
 sg13g2_nand2_1 _4488_ (.Y(_1237_),
    .A(net156),
    .B(_0659_));
 sg13g2_xnor2_1 _4489_ (.Y(_1238_),
    .A(_1236_),
    .B(_1237_));
 sg13g2_nor2_1 _4490_ (.A(_1234_),
    .B(_1238_),
    .Y(_0266_));
 sg13g2_nand2_1 _4491_ (.Y(_1239_),
    .A(_0659_),
    .B(net155));
 sg13g2_nand2_1 _4492_ (.Y(_1240_),
    .A(net143),
    .B(_1239_));
 sg13g2_xor2_1 _4493_ (.B(net154),
    .A(net143),
    .X(_1241_));
 sg13g2_nand2_1 _4494_ (.Y(_1242_),
    .A(net144),
    .B(_1241_));
 sg13g2_o21ai_1 _4495_ (.B1(_1242_),
    .Y(_1243_),
    .A1(net144),
    .A2(_1240_));
 sg13g2_a21o_1 _4496_ (.A2(net143),
    .A1(net156),
    .B1(net144),
    .X(_1244_));
 sg13g2_o21ai_1 _4497_ (.B1(_1244_),
    .Y(_1245_),
    .A1(net156),
    .A2(net154));
 sg13g2_and2_1 _4498_ (.A(_0659_),
    .B(net155),
    .X(_1246_));
 sg13g2_buf_1 _4499_ (.A(_1246_),
    .X(_1247_));
 sg13g2_nand2_1 _4500_ (.Y(_1248_),
    .A(net144),
    .B(net154));
 sg13g2_nor3_1 _4501_ (.A(net156),
    .B(_1247_),
    .C(_1248_),
    .Y(_1249_));
 sg13g2_a221oi_1 _4502_ (.B2(_1247_),
    .C1(_1249_),
    .B1(_1245_),
    .A1(net156),
    .Y(_1250_),
    .A2(_1243_));
 sg13g2_nor2_1 _4503_ (.A(_1234_),
    .B(_1250_),
    .Y(_0267_));
 sg13g2_nand2_1 _4504_ (.Y(_1251_),
    .A(\mem[17][0] ),
    .B(_0662_));
 sg13g2_nand2_1 _4505_ (.Y(_1252_),
    .A(net155),
    .B(\mem[1][2] ));
 sg13g2_nand2_1 _4506_ (.Y(_1253_),
    .A(_0659_),
    .B(net154));
 sg13g2_xor2_1 _4507_ (.B(_1253_),
    .A(_1252_),
    .X(_1254_));
 sg13g2_xnor2_1 _4508_ (.Y(_1255_),
    .A(_1251_),
    .B(_1254_));
 sg13g2_buf_2 _4509_ (.A(_1255_),
    .X(_1256_));
 sg13g2_a21oi_1 _4510_ (.A1(_0624_),
    .A2(net143),
    .Y(_1257_),
    .B1(_1247_));
 sg13g2_nand3_1 _4511_ (.B(net143),
    .C(_1247_),
    .A(_0624_),
    .Y(_1258_));
 sg13g2_o21ai_1 _4512_ (.B1(_1258_),
    .Y(_1259_),
    .A1(_1248_),
    .A2(_1257_));
 sg13g2_buf_1 _4513_ (.A(_1259_),
    .X(_1260_));
 sg13g2_nand2_2 _4514_ (.Y(_1261_),
    .A(_0654_),
    .B(net153));
 sg13g2_nor3_2 _4515_ (.A(_1235_),
    .B(_1241_),
    .C(_1239_),
    .Y(_1262_));
 sg13g2_xor2_1 _4516_ (.B(_1262_),
    .A(_1261_),
    .X(_1263_));
 sg13g2_xnor2_1 _4517_ (.Y(_1264_),
    .A(_1260_),
    .B(_1263_));
 sg13g2_xnor2_1 _4518_ (.Y(_1265_),
    .A(_1256_),
    .B(_1264_));
 sg13g2_nor2_1 _4519_ (.A(_1234_),
    .B(_1265_),
    .Y(_0268_));
 sg13g2_and2_1 _4520_ (.A(_1252_),
    .B(_1253_),
    .X(_1266_));
 sg13g2_or2_1 _4521_ (.X(_1267_),
    .B(_1253_),
    .A(_1252_));
 sg13g2_o21ai_1 _4522_ (.B1(_1267_),
    .Y(_1268_),
    .A1(_1251_),
    .A2(_1266_));
 sg13g2_nand2_2 _4523_ (.Y(_1269_),
    .A(net143),
    .B(net154));
 sg13g2_nand2_1 _4524_ (.Y(_1270_),
    .A(net155),
    .B(_0662_));
 sg13g2_xor2_1 _4525_ (.B(_1270_),
    .A(_1269_),
    .X(_1271_));
 sg13g2_nand2_1 _4526_ (.Y(_1272_),
    .A(_0659_),
    .B(\mem[17][3] ));
 sg13g2_xor2_1 _4527_ (.B(_1272_),
    .A(_1271_),
    .X(_1273_));
 sg13g2_xnor2_1 _4528_ (.Y(_1274_),
    .A(_1268_),
    .B(_1273_));
 sg13g2_nand2_1 _4529_ (.Y(_1275_),
    .A(_1260_),
    .B(_1256_));
 sg13g2_nor2_1 _4530_ (.A(_1260_),
    .B(_1256_),
    .Y(_1276_));
 sg13g2_a21oi_1 _4531_ (.A1(_1261_),
    .A2(_1275_),
    .Y(_1277_),
    .B1(_1276_));
 sg13g2_inv_1 _4532_ (.Y(_1278_),
    .A(_1262_));
 sg13g2_nor3_1 _4533_ (.A(_1261_),
    .B(_1278_),
    .C(_1275_),
    .Y(_1279_));
 sg13g2_a21oi_1 _4534_ (.A1(_1261_),
    .A2(_1276_),
    .Y(_1280_),
    .B1(_1279_));
 sg13g2_o21ai_1 _4535_ (.B1(_1280_),
    .Y(_1281_),
    .A1(_1262_),
    .A2(_1277_));
 sg13g2_xor2_1 _4536_ (.B(_1281_),
    .A(_1274_),
    .X(_1282_));
 sg13g2_nor2_1 _4537_ (.A(_1234_),
    .B(_1282_),
    .Y(_0269_));
 sg13g2_and2_1 _4538_ (.A(_1256_),
    .B(_1262_),
    .X(_1283_));
 sg13g2_o21ai_1 _4539_ (.B1(_1260_),
    .Y(_1284_),
    .A1(_1256_),
    .A2(_1262_));
 sg13g2_nand2b_1 _4540_ (.Y(_1285_),
    .B(_1284_),
    .A_N(_1283_));
 sg13g2_o21ai_1 _4541_ (.B1(_1260_),
    .Y(_1286_),
    .A1(_1274_),
    .A2(_1283_));
 sg13g2_o21ai_1 _4542_ (.B1(_1274_),
    .Y(_1287_),
    .A1(_1256_),
    .A2(_1262_));
 sg13g2_a21oi_1 _4543_ (.A1(_1286_),
    .A2(_1287_),
    .Y(_1288_),
    .B1(_1261_));
 sg13g2_a21oi_1 _4544_ (.A1(_1274_),
    .A2(_1285_),
    .Y(_1289_),
    .B1(_1288_));
 sg13g2_nor2_1 _4545_ (.A(_1268_),
    .B(_1271_),
    .Y(_1290_));
 sg13g2_a22oi_1 _4546_ (.Y(_1291_),
    .B1(_1268_),
    .B2(_1271_),
    .A2(net153),
    .A1(_0659_));
 sg13g2_nor2_1 _4547_ (.A(_1290_),
    .B(_1291_),
    .Y(_1292_));
 sg13g2_o21ai_1 _4548_ (.B1(_0660_),
    .Y(_1293_),
    .A1(net155),
    .A2(net153));
 sg13g2_nand3_1 _4549_ (.B(_0662_),
    .C(_1293_),
    .A(net154),
    .Y(_1294_));
 sg13g2_nand3_1 _4550_ (.B(_0635_),
    .C(_0662_),
    .A(_0632_),
    .Y(_1295_));
 sg13g2_nand3_1 _4551_ (.B(_0636_),
    .C(_1295_),
    .A(_0660_),
    .Y(_1296_));
 sg13g2_and2_1 _4552_ (.A(_1294_),
    .B(_1296_),
    .X(_1297_));
 sg13g2_nor2b_1 _4553_ (.A(_1292_),
    .B_N(_1297_),
    .Y(_1298_));
 sg13g2_or3_1 _4554_ (.A(_1290_),
    .B(_1291_),
    .C(_1297_),
    .X(_1299_));
 sg13g2_nand2b_1 _4555_ (.Y(_1300_),
    .B(_1299_),
    .A_N(_1298_));
 sg13g2_xnor2_1 _4556_ (.Y(_1301_),
    .A(_1289_),
    .B(_1300_));
 sg13g2_nor2_1 _4557_ (.A(_1234_),
    .B(_1301_),
    .Y(_0270_));
 sg13g2_a21oi_2 _4558_ (.B1(_1298_),
    .Y(_1302_),
    .A2(_1299_),
    .A1(_1289_));
 sg13g2_nor3_1 _4559_ (.A(_0632_),
    .B(net153),
    .C(_1269_),
    .Y(_1303_));
 sg13g2_a21oi_1 _4560_ (.A1(net153),
    .A2(_1269_),
    .Y(_1304_),
    .B1(_1303_));
 sg13g2_nor2b_1 _4561_ (.A(_1304_),
    .B_N(_0662_),
    .Y(_1305_));
 sg13g2_xnor2_1 _4562_ (.Y(_1306_),
    .A(_1302_),
    .B(_1305_));
 sg13g2_nor2_1 _4563_ (.A(_1234_),
    .B(_1306_),
    .Y(_0271_));
 sg13g2_and2_1 _4564_ (.A(_2606_),
    .B(net61),
    .X(_1307_));
 sg13g2_buf_1 _4565_ (.A(_1307_),
    .X(_1308_));
 sg13g2_buf_1 _4566_ (.A(_1308_),
    .X(_1309_));
 sg13g2_a21oi_1 _4567_ (.A1(_0631_),
    .A2(_1302_),
    .Y(_1310_),
    .B1(net153));
 sg13g2_nand2_1 _4568_ (.Y(_1311_),
    .A(net153),
    .B(_1302_));
 sg13g2_o21ai_1 _4569_ (.B1(_1311_),
    .Y(_1312_),
    .A1(_1269_),
    .A2(_1310_));
 sg13g2_and3_1 _4570_ (.X(_0272_),
    .A(_0662_),
    .B(_1309_),
    .C(_1312_));
 sg13g2_buf_1 _4571_ (.A(_0000_),
    .X(_1313_));
 sg13g2_nand2_1 _4572_ (.Y(_1314_),
    .A(net81),
    .B(_1313_));
 sg13g2_nand2b_1 _4573_ (.Y(_1315_),
    .B(net174),
    .A_N(net175));
 sg13g2_a21oi_1 _4574_ (.A1(_1314_),
    .A2(_1315_),
    .Y(_1316_),
    .B1(net173));
 sg13g2_nor2_1 _4575_ (.A(net175),
    .B(net173),
    .Y(_1317_));
 sg13g2_o21ai_1 _4576_ (.B1(net57),
    .Y(_1318_),
    .A1(net81),
    .A2(_1317_));
 sg13g2_or2_1 _4577_ (.X(_1319_),
    .B(_1318_),
    .A(_1316_));
 sg13g2_buf_2 _4578_ (.A(_1319_),
    .X(_1320_));
 sg13g2_nor3_1 _4579_ (.A(_0572_),
    .B(_0718_),
    .C(_1320_),
    .Y(_0273_));
 sg13g2_buf_1 _4580_ (.A(_0571_),
    .X(_1321_));
 sg13g2_buf_1 _4581_ (.A(_0721_),
    .X(_1322_));
 sg13g2_nand2_1 _4582_ (.Y(_1323_),
    .A(net76),
    .B(net75));
 sg13g2_nand2_1 _4583_ (.Y(_1324_),
    .A(_0717_),
    .B(net80));
 sg13g2_xnor2_1 _4584_ (.Y(_1325_),
    .A(_1323_),
    .B(_1324_));
 sg13g2_nor2_1 _4585_ (.A(_1320_),
    .B(_1325_),
    .Y(_0274_));
 sg13g2_nand2_1 _4586_ (.Y(_1326_),
    .A(net80),
    .B(net75));
 sg13g2_nor2b_1 _4587_ (.A(net76),
    .B_N(net63),
    .Y(_1327_));
 sg13g2_xor2_1 _4588_ (.B(net78),
    .A(net63),
    .X(_1328_));
 sg13g2_a22oi_1 _4589_ (.Y(_1329_),
    .B1(_1328_),
    .B2(net76),
    .A2(_1327_),
    .A1(_1326_));
 sg13g2_nand2b_1 _4590_ (.Y(_1330_),
    .B(_0717_),
    .A_N(_1329_));
 sg13g2_a21oi_1 _4591_ (.A1(_0717_),
    .A2(net63),
    .Y(_1331_),
    .B1(net76));
 sg13g2_nor2_1 _4592_ (.A(_0717_),
    .B(net78),
    .Y(_1332_));
 sg13g2_and2_1 _4593_ (.A(net80),
    .B(net75),
    .X(_1333_));
 sg13g2_o21ai_1 _4594_ (.B1(_1333_),
    .Y(_1334_),
    .A1(_1331_),
    .A2(_1332_));
 sg13g2_nand4_1 _4595_ (.B(_0718_),
    .C(net78),
    .A(net76),
    .Y(_1335_),
    .D(_1326_));
 sg13g2_nand3_1 _4596_ (.B(_1334_),
    .C(_1335_),
    .A(_1330_),
    .Y(_1336_));
 sg13g2_nor2b_1 _4597_ (.A(_1320_),
    .B_N(_1336_),
    .Y(_0275_));
 sg13g2_nand2_1 _4598_ (.Y(_1337_),
    .A(_0581_),
    .B(net121));
 sg13g2_o21ai_1 _4599_ (.B1(_1337_),
    .Y(_1338_),
    .A1(net121),
    .A2(_1326_));
 sg13g2_a22oi_1 _4600_ (.Y(_1339_),
    .B1(_1338_),
    .B2(net76),
    .A2(_1333_),
    .A1(net63));
 sg13g2_nand2b_1 _4601_ (.Y(_1340_),
    .B(_0717_),
    .A_N(_1339_));
 sg13g2_nand2_1 _4602_ (.Y(_1341_),
    .A(_0717_),
    .B(net168));
 sg13g2_xor2_1 _4603_ (.B(_0726_),
    .A(_0581_),
    .X(_1342_));
 sg13g2_nand4_1 _4604_ (.B(_0579_),
    .C(net79),
    .A(_0572_),
    .Y(_1343_),
    .D(net121));
 sg13g2_o21ai_1 _4605_ (.B1(_1343_),
    .Y(_1344_),
    .A1(_0572_),
    .A2(_1342_));
 sg13g2_a21o_1 _4606_ (.A2(net79),
    .A1(_0721_),
    .B1(_0571_),
    .X(_1345_));
 sg13g2_o21ai_1 _4607_ (.B1(_1345_),
    .Y(_1346_),
    .A1(net75),
    .A2(net77));
 sg13g2_nand2_1 _4608_ (.Y(_1347_),
    .A(_0579_),
    .B(net121));
 sg13g2_buf_1 _4609_ (.A(_1347_),
    .X(_1348_));
 sg13g2_nand2_1 _4610_ (.Y(_1349_),
    .A(net76),
    .B(_0726_));
 sg13g2_nor3_1 _4611_ (.A(net75),
    .B(net60),
    .C(_1349_),
    .Y(_1350_));
 sg13g2_a221oi_1 _4612_ (.B2(net60),
    .C1(_1350_),
    .B1(_1346_),
    .A1(net75),
    .Y(_1351_),
    .A2(_1344_));
 sg13g2_xnor2_1 _4613_ (.Y(_1352_),
    .A(_1341_),
    .B(_1351_));
 sg13g2_nor2b_2 _4614_ (.A(_1340_),
    .B_N(_1352_),
    .Y(_1353_));
 sg13g2_nor2b_1 _4615_ (.A(_1352_),
    .B_N(_1340_),
    .Y(_1354_));
 sg13g2_nor3_1 _4616_ (.A(_1320_),
    .B(_1353_),
    .C(_1354_),
    .Y(_0276_));
 sg13g2_nand2_1 _4617_ (.Y(_1355_),
    .A(_0721_),
    .B(\mem[11][3] ));
 sg13g2_nand2_1 _4618_ (.Y(_1356_),
    .A(_0579_),
    .B(_0726_));
 sg13g2_xnor2_1 _4619_ (.Y(_1357_),
    .A(_1355_),
    .B(_1356_));
 sg13g2_xnor2_1 _4620_ (.Y(_1358_),
    .A(_1337_),
    .B(_1357_));
 sg13g2_nand4_1 _4621_ (.B(_0721_),
    .C(net79),
    .A(net80),
    .Y(_1359_),
    .D(net121));
 sg13g2_a22oi_1 _4622_ (.Y(_1360_),
    .B1(net121),
    .B2(net80),
    .A2(net79),
    .A1(_0721_));
 sg13g2_a21oi_1 _4623_ (.A1(_1349_),
    .A2(_1359_),
    .Y(_1361_),
    .B1(_1360_));
 sg13g2_xor2_1 _4624_ (.B(_1361_),
    .A(_1358_),
    .X(_1362_));
 sg13g2_nand3_1 _4625_ (.B(net79),
    .C(net60),
    .A(_0721_),
    .Y(_1363_));
 sg13g2_o21ai_1 _4626_ (.B1(_1363_),
    .Y(_1364_),
    .A1(net79),
    .A2(net60));
 sg13g2_nand2_1 _4627_ (.Y(_1365_),
    .A(_0572_),
    .B(_1364_));
 sg13g2_nand3_1 _4628_ (.B(_0726_),
    .C(net60),
    .A(_0571_),
    .Y(_1366_));
 sg13g2_o21ai_1 _4629_ (.B1(_1366_),
    .Y(_1367_),
    .A1(net76),
    .A2(net60));
 sg13g2_nand2_1 _4630_ (.Y(_1368_),
    .A(_0721_),
    .B(_1342_));
 sg13g2_o21ai_1 _4631_ (.B1(_1368_),
    .Y(_1369_),
    .A1(net77),
    .A2(_1348_));
 sg13g2_a22oi_1 _4632_ (.Y(_1370_),
    .B1(_1369_),
    .B2(_1321_),
    .A2(_1367_),
    .A1(_0722_));
 sg13g2_a21oi_1 _4633_ (.A1(_1365_),
    .A2(_1370_),
    .Y(_1371_),
    .B1(_1341_));
 sg13g2_nor3_1 _4634_ (.A(_1323_),
    .B(_1342_),
    .C(net60),
    .Y(_1372_));
 sg13g2_nor2_1 _4635_ (.A(_1371_),
    .B(_1372_),
    .Y(_1373_));
 sg13g2_xor2_1 _4636_ (.B(_1373_),
    .A(_1362_),
    .X(_1374_));
 sg13g2_xnor2_1 _4637_ (.Y(_1375_),
    .A(_1353_),
    .B(_1374_));
 sg13g2_nor2_1 _4638_ (.A(_1320_),
    .B(_1375_),
    .Y(_0277_));
 sg13g2_nor2_1 _4639_ (.A(_1362_),
    .B(_1373_),
    .Y(_1376_));
 sg13g2_a21oi_2 _4640_ (.B1(_1376_),
    .Y(_1377_),
    .A2(_1374_),
    .A1(_1353_));
 sg13g2_nand2b_1 _4641_ (.Y(_1378_),
    .B(_1361_),
    .A_N(_1358_));
 sg13g2_inv_1 _4642_ (.Y(_1379_),
    .A(net77));
 sg13g2_nand2_1 _4643_ (.Y(_1380_),
    .A(net78),
    .B(net77));
 sg13g2_nand3b_1 _4644_ (.B(net168),
    .C(net79),
    .Y(_1381_),
    .A_N(net78));
 sg13g2_o21ai_1 _4645_ (.B1(_1381_),
    .Y(_1382_),
    .A1(net63),
    .A2(_1380_));
 sg13g2_a22oi_1 _4646_ (.Y(_1383_),
    .B1(_1382_),
    .B2(net80),
    .A2(_1379_),
    .A1(net63));
 sg13g2_o21ai_1 _4647_ (.B1(net168),
    .Y(_1384_),
    .A1(net75),
    .A2(_0725_));
 sg13g2_nor2b_1 _4648_ (.A(_0583_),
    .B_N(_1384_),
    .Y(_1385_));
 sg13g2_nor2_1 _4649_ (.A(_0725_),
    .B(net77),
    .Y(_1386_));
 sg13g2_a21oi_1 _4650_ (.A1(net77),
    .A2(net60),
    .Y(_1387_),
    .B1(net168));
 sg13g2_and3_1 _4651_ (.X(_1388_),
    .A(_0582_),
    .B(net121),
    .C(_0727_));
 sg13g2_nor2b_1 _4652_ (.A(net75),
    .B_N(net168),
    .Y(_1389_));
 sg13g2_nor2_1 _4653_ (.A(_0582_),
    .B(_0724_),
    .Y(_1390_));
 sg13g2_a21oi_1 _4654_ (.A1(_1388_),
    .A2(_1389_),
    .Y(_1391_),
    .B1(_1390_));
 sg13g2_nor2_1 _4655_ (.A(net80),
    .B(_1391_),
    .Y(_1392_));
 sg13g2_nor4_1 _4656_ (.A(_1385_),
    .B(_1386_),
    .C(_1387_),
    .D(_1392_),
    .Y(_1393_));
 sg13g2_o21ai_1 _4657_ (.B1(_1393_),
    .Y(_1394_),
    .A1(_0722_),
    .A2(_1383_));
 sg13g2_xnor2_1 _4658_ (.Y(_1395_),
    .A(_1378_),
    .B(_1394_));
 sg13g2_xnor2_1 _4659_ (.Y(_1396_),
    .A(_1377_),
    .B(_1395_));
 sg13g2_nor2_1 _4660_ (.A(_1320_),
    .B(_1396_),
    .Y(_0278_));
 sg13g2_nand2_1 _4661_ (.Y(_1397_),
    .A(_1377_),
    .B(_1394_));
 sg13g2_o21ai_1 _4662_ (.B1(_1378_),
    .Y(_1398_),
    .A1(_1377_),
    .A2(_1394_));
 sg13g2_nand2_1 _4663_ (.Y(_1399_),
    .A(_1397_),
    .B(_1398_));
 sg13g2_a21oi_1 _4664_ (.A1(_1326_),
    .A2(_1337_),
    .Y(_1400_),
    .B1(_1390_));
 sg13g2_nand4_1 _4665_ (.B(net63),
    .C(net78),
    .A(_1322_),
    .Y(_1401_),
    .D(_1379_));
 sg13g2_o21ai_1 _4666_ (.B1(_1401_),
    .Y(_1402_),
    .A1(_1379_),
    .A2(_1400_));
 sg13g2_nor2b_1 _4667_ (.A(net168),
    .B_N(_0580_),
    .Y(_1403_));
 sg13g2_a22oi_1 _4668_ (.Y(_1404_),
    .B1(_1403_),
    .B2(_1388_),
    .A2(_1402_),
    .A1(net168));
 sg13g2_xnor2_1 _4669_ (.Y(_1405_),
    .A(_1399_),
    .B(_1404_));
 sg13g2_nor2_1 _4670_ (.A(_1320_),
    .B(_1405_),
    .Y(_0279_));
 sg13g2_nand3_1 _4671_ (.B(_0727_),
    .C(_1400_),
    .A(_0584_),
    .Y(_1406_));
 sg13g2_o21ai_1 _4672_ (.B1(_1406_),
    .Y(_1407_),
    .A1(_1399_),
    .A2(_1404_));
 sg13g2_nor2b_1 _4673_ (.A(_1320_),
    .B_N(_1407_),
    .Y(_0280_));
 sg13g2_nor3_2 _4674_ (.A(net175),
    .B(net174),
    .C(\mem[0][2] ),
    .Y(_1408_));
 sg13g2_nor2b_1 _4675_ (.A(_0557_),
    .B_N(_1408_),
    .Y(_1409_));
 sg13g2_nand2_1 _4676_ (.Y(_1410_),
    .A(\mem[0][2] ),
    .B(_0557_));
 sg13g2_nand2b_1 _4677_ (.Y(_1411_),
    .B(_1410_),
    .A_N(_1409_));
 sg13g2_nand2_1 _4678_ (.Y(_1412_),
    .A(net57),
    .B(_1411_));
 sg13g2_buf_1 _4679_ (.A(_1412_),
    .X(_1413_));
 sg13g2_nand2_1 _4680_ (.Y(_1414_),
    .A(net167),
    .B(net120));
 sg13g2_nor2_1 _4681_ (.A(net53),
    .B(_1414_),
    .Y(_0281_));
 sg13g2_nand2_1 _4682_ (.Y(_1415_),
    .A(net167),
    .B(net119));
 sg13g2_nand2_1 _4683_ (.Y(_1416_),
    .A(net120),
    .B(_0591_));
 sg13g2_xnor2_1 _4684_ (.Y(_1417_),
    .A(_1415_),
    .B(_1416_));
 sg13g2_nor2_1 _4685_ (.A(net53),
    .B(_1417_),
    .Y(_0282_));
 sg13g2_nand2_1 _4686_ (.Y(_1418_),
    .A(_0591_),
    .B(net119));
 sg13g2_nand2_1 _4687_ (.Y(_1419_),
    .A(net165),
    .B(_1418_));
 sg13g2_xor2_1 _4688_ (.B(net118),
    .A(net165),
    .X(_1420_));
 sg13g2_nand2_1 _4689_ (.Y(_1421_),
    .A(net167),
    .B(_1420_));
 sg13g2_o21ai_1 _4690_ (.B1(_1421_),
    .Y(_1422_),
    .A1(net167),
    .A2(_1419_));
 sg13g2_a21o_1 _4691_ (.A2(net165),
    .A1(net120),
    .B1(net167),
    .X(_1423_));
 sg13g2_o21ai_1 _4692_ (.B1(_1423_),
    .Y(_1424_),
    .A1(net120),
    .A2(net118));
 sg13g2_and2_1 _4693_ (.A(_0591_),
    .B(_0730_),
    .X(_1425_));
 sg13g2_buf_1 _4694_ (.A(_1425_),
    .X(_1426_));
 sg13g2_nand2_1 _4695_ (.Y(_1427_),
    .A(net167),
    .B(net118));
 sg13g2_nor3_1 _4696_ (.A(net120),
    .B(_1426_),
    .C(_1427_),
    .Y(_1428_));
 sg13g2_a221oi_1 _4697_ (.B2(_1426_),
    .C1(_1428_),
    .B1(_1424_),
    .A1(net120),
    .Y(_1429_),
    .A2(_1422_));
 sg13g2_nor2_1 _4698_ (.A(net53),
    .B(_1429_),
    .Y(_0283_));
 sg13g2_nand2_1 _4699_ (.Y(_1430_),
    .A(\mem[28][0] ),
    .B(_0593_));
 sg13g2_nand2_1 _4700_ (.Y(_1431_),
    .A(net119),
    .B(\mem[12][2] ));
 sg13g2_nand2_1 _4701_ (.Y(_1432_),
    .A(_0591_),
    .B(net118));
 sg13g2_xor2_1 _4702_ (.B(_1432_),
    .A(_1431_),
    .X(_1433_));
 sg13g2_xnor2_1 _4703_ (.Y(_1434_),
    .A(_1430_),
    .B(_1433_));
 sg13g2_buf_1 _4704_ (.A(_1434_),
    .X(_1435_));
 sg13g2_a21oi_1 _4705_ (.A1(_0728_),
    .A2(_0592_),
    .Y(_1436_),
    .B1(_1426_));
 sg13g2_nand3_1 _4706_ (.B(_0592_),
    .C(_1426_),
    .A(_0728_),
    .Y(_1437_));
 sg13g2_o21ai_1 _4707_ (.B1(_1437_),
    .Y(_1438_),
    .A1(_1427_),
    .A2(_1436_));
 sg13g2_buf_1 _4708_ (.A(_1438_),
    .X(_1439_));
 sg13g2_nand2_2 _4709_ (.Y(_1440_),
    .A(_0585_),
    .B(net117));
 sg13g2_nor3_2 _4710_ (.A(_1414_),
    .B(_1420_),
    .C(_1418_),
    .Y(_1441_));
 sg13g2_xor2_1 _4711_ (.B(_1441_),
    .A(_1440_),
    .X(_1442_));
 sg13g2_xnor2_1 _4712_ (.Y(_1443_),
    .A(_1439_),
    .B(_1442_));
 sg13g2_xnor2_1 _4713_ (.Y(_1444_),
    .A(_1435_),
    .B(_1443_));
 sg13g2_nor2_1 _4714_ (.A(net53),
    .B(_1444_),
    .Y(_0284_));
 sg13g2_and2_1 _4715_ (.A(_1431_),
    .B(_1432_),
    .X(_1445_));
 sg13g2_or2_1 _4716_ (.X(_1446_),
    .B(_1432_),
    .A(_1431_));
 sg13g2_o21ai_1 _4717_ (.B1(_1446_),
    .Y(_1447_),
    .A1(_1430_),
    .A2(_1445_));
 sg13g2_nand2_2 _4718_ (.Y(_1448_),
    .A(net165),
    .B(_0733_));
 sg13g2_nand2_1 _4719_ (.Y(_1449_),
    .A(net119),
    .B(_0593_));
 sg13g2_xor2_1 _4720_ (.B(_1449_),
    .A(_1448_),
    .X(_1450_));
 sg13g2_nand2_1 _4721_ (.Y(_1451_),
    .A(_0591_),
    .B(\mem[28][3] ));
 sg13g2_xor2_1 _4722_ (.B(_1451_),
    .A(_1450_),
    .X(_1452_));
 sg13g2_xnor2_1 _4723_ (.Y(_1453_),
    .A(_1447_),
    .B(_1452_));
 sg13g2_nand2_1 _4724_ (.Y(_1454_),
    .A(_1439_),
    .B(_1435_));
 sg13g2_nor2_1 _4725_ (.A(_1439_),
    .B(_1435_),
    .Y(_1455_));
 sg13g2_a21oi_1 _4726_ (.A1(_1440_),
    .A2(_1454_),
    .Y(_1456_),
    .B1(_1455_));
 sg13g2_inv_1 _4727_ (.Y(_1457_),
    .A(_1441_));
 sg13g2_nor3_1 _4728_ (.A(_1440_),
    .B(_1457_),
    .C(_1454_),
    .Y(_1458_));
 sg13g2_a21oi_1 _4729_ (.A1(_1440_),
    .A2(_1455_),
    .Y(_1459_),
    .B1(_1458_));
 sg13g2_o21ai_1 _4730_ (.B1(_1459_),
    .Y(_1460_),
    .A1(_1441_),
    .A2(_1456_));
 sg13g2_xor2_1 _4731_ (.B(_1460_),
    .A(_1453_),
    .X(_1461_));
 sg13g2_nor2_1 _4732_ (.A(net53),
    .B(_1461_),
    .Y(_0285_));
 sg13g2_and2_1 _4733_ (.A(_1435_),
    .B(_1441_),
    .X(_1462_));
 sg13g2_o21ai_1 _4734_ (.B1(_1439_),
    .Y(_1463_),
    .A1(_1435_),
    .A2(_1441_));
 sg13g2_nand2b_1 _4735_ (.Y(_1464_),
    .B(_1463_),
    .A_N(_1462_));
 sg13g2_o21ai_1 _4736_ (.B1(_1439_),
    .Y(_1465_),
    .A1(_1453_),
    .A2(_1462_));
 sg13g2_o21ai_1 _4737_ (.B1(_1453_),
    .Y(_1466_),
    .A1(_1435_),
    .A2(_1441_));
 sg13g2_a21oi_1 _4738_ (.A1(_1465_),
    .A2(_1466_),
    .Y(_1467_),
    .B1(_1440_));
 sg13g2_a21oi_1 _4739_ (.A1(_1453_),
    .A2(_1464_),
    .Y(_1468_),
    .B1(_1467_));
 sg13g2_nor2_1 _4740_ (.A(_1447_),
    .B(_1450_),
    .Y(_1469_));
 sg13g2_a22oi_1 _4741_ (.Y(_1470_),
    .B1(_1447_),
    .B2(_1450_),
    .A2(net117),
    .A1(_0591_));
 sg13g2_nor2_1 _4742_ (.A(_1469_),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_o21ai_1 _4743_ (.B1(net165),
    .Y(_1472_),
    .A1(net119),
    .A2(net117));
 sg13g2_nand3_1 _4744_ (.B(_0593_),
    .C(_1472_),
    .A(net118),
    .Y(_1473_));
 sg13g2_nand3_1 _4745_ (.B(net118),
    .C(_0593_),
    .A(_0731_),
    .Y(_1474_));
 sg13g2_nand3_1 _4746_ (.B(net117),
    .C(_1474_),
    .A(net165),
    .Y(_1475_));
 sg13g2_and2_1 _4747_ (.A(_1473_),
    .B(_1475_),
    .X(_1476_));
 sg13g2_nor2b_1 _4748_ (.A(_1471_),
    .B_N(_1476_),
    .Y(_1477_));
 sg13g2_or3_1 _4749_ (.A(_1469_),
    .B(_1470_),
    .C(_1476_),
    .X(_1478_));
 sg13g2_nand2b_1 _4750_ (.Y(_1479_),
    .B(_1478_),
    .A_N(_1477_));
 sg13g2_xnor2_1 _4751_ (.Y(_1480_),
    .A(_1468_),
    .B(_1479_));
 sg13g2_nor2_1 _4752_ (.A(net53),
    .B(_1480_),
    .Y(_0286_));
 sg13g2_a21oi_2 _4753_ (.B1(_1477_),
    .Y(_1481_),
    .A2(_1478_),
    .A1(_1468_));
 sg13g2_inv_1 _4754_ (.Y(_1482_),
    .A(_0593_));
 sg13g2_nor3_1 _4755_ (.A(_0731_),
    .B(net117),
    .C(_1448_),
    .Y(_1483_));
 sg13g2_a21oi_1 _4756_ (.A1(net117),
    .A2(_1448_),
    .Y(_1484_),
    .B1(_1483_));
 sg13g2_nor2_1 _4757_ (.A(_1482_),
    .B(_1484_),
    .Y(_1485_));
 sg13g2_xnor2_1 _4758_ (.Y(_1486_),
    .A(_1481_),
    .B(_1485_));
 sg13g2_nor2_1 _4759_ (.A(_1413_),
    .B(_1486_),
    .Y(_0287_));
 sg13g2_a21oi_1 _4760_ (.A1(net119),
    .A2(_1481_),
    .Y(_1487_),
    .B1(_0734_));
 sg13g2_nor2_1 _4761_ (.A(_1448_),
    .B(_1487_),
    .Y(_1488_));
 sg13g2_a21oi_1 _4762_ (.A1(_0734_),
    .A2(_1481_),
    .Y(_1489_),
    .B1(_1488_));
 sg13g2_nor3_1 _4763_ (.A(_1482_),
    .B(net53),
    .C(_1489_),
    .Y(_0288_));
 sg13g2_nor2_1 _4764_ (.A(net175),
    .B(net174),
    .Y(_1490_));
 sg13g2_nand2_1 _4765_ (.Y(_1491_),
    .A(_1308_),
    .B(_1409_));
 sg13g2_buf_1 _4766_ (.A(_1491_),
    .X(_1492_));
 sg13g2_a21o_1 _4767_ (.A2(_1492_),
    .A1(_1490_),
    .B1(net53),
    .X(_1493_));
 sg13g2_buf_2 _4768_ (.A(_1493_),
    .X(_1494_));
 sg13g2_nand2_1 _4769_ (.Y(_1495_),
    .A(net116),
    .B(net164));
 sg13g2_nor2_1 _4770_ (.A(_1494_),
    .B(_1495_),
    .Y(_0289_));
 sg13g2_nand2_1 _4771_ (.Y(_1496_),
    .A(_0737_),
    .B(net164));
 sg13g2_nand2_1 _4772_ (.Y(_1497_),
    .A(net116),
    .B(_0599_));
 sg13g2_xnor2_1 _4773_ (.Y(_1498_),
    .A(_1496_),
    .B(_1497_));
 sg13g2_nor2_1 _4774_ (.A(_1494_),
    .B(_1498_),
    .Y(_0290_));
 sg13g2_nand2_1 _4775_ (.Y(_1499_),
    .A(_0599_),
    .B(_0737_));
 sg13g2_buf_2 _4776_ (.A(_1499_),
    .X(_1500_));
 sg13g2_nand2_1 _4777_ (.Y(_1501_),
    .A(net163),
    .B(_1500_));
 sg13g2_xor2_1 _4778_ (.B(_0741_),
    .A(net163),
    .X(_1502_));
 sg13g2_nand2_1 _4779_ (.Y(_1503_),
    .A(net164),
    .B(_1502_));
 sg13g2_o21ai_1 _4780_ (.B1(_1503_),
    .Y(_1504_),
    .A1(net164),
    .A2(_1501_));
 sg13g2_nand2_2 _4781_ (.Y(_1505_),
    .A(net164),
    .B(_0741_));
 sg13g2_nor2_1 _4782_ (.A(net116),
    .B(_1505_),
    .Y(_1506_));
 sg13g2_nand2b_1 _4783_ (.Y(_1507_),
    .B(_1505_),
    .A_N(net116));
 sg13g2_or2_1 _4784_ (.X(_1508_),
    .B(net163),
    .A(net164));
 sg13g2_a21oi_1 _4785_ (.A1(_1507_),
    .A2(_1508_),
    .Y(_1509_),
    .B1(_1500_));
 sg13g2_a221oi_1 _4786_ (.B2(_1500_),
    .C1(_1509_),
    .B1(_1506_),
    .A1(net116),
    .Y(_1510_),
    .A2(_1504_));
 sg13g2_nor2_1 _4787_ (.A(_1494_),
    .B(_1510_),
    .Y(_0291_));
 sg13g2_nand2_1 _4788_ (.Y(_1511_),
    .A(net116),
    .B(_0601_));
 sg13g2_nand2_1 _4789_ (.Y(_1512_),
    .A(_0737_),
    .B(net163));
 sg13g2_nand2_1 _4790_ (.Y(_1513_),
    .A(_0599_),
    .B(_0741_));
 sg13g2_xor2_1 _4791_ (.B(_1513_),
    .A(_1512_),
    .X(_1514_));
 sg13g2_xnor2_1 _4792_ (.Y(_1515_),
    .A(_1511_),
    .B(_1514_));
 sg13g2_buf_1 _4793_ (.A(_1515_),
    .X(_1516_));
 sg13g2_nor2_1 _4794_ (.A(_1500_),
    .B(_1505_),
    .Y(_1517_));
 sg13g2_a21oi_1 _4795_ (.A1(_0735_),
    .A2(net163),
    .Y(_1518_),
    .B1(_1517_));
 sg13g2_a21oi_2 _4796_ (.B1(_1518_),
    .Y(_1519_),
    .A2(_1505_),
    .A1(_1500_));
 sg13g2_nand2_2 _4797_ (.Y(_1520_),
    .A(_0594_),
    .B(net115));
 sg13g2_nor3_2 _4798_ (.A(_1495_),
    .B(_1502_),
    .C(_1500_),
    .Y(_1521_));
 sg13g2_xor2_1 _4799_ (.B(_1521_),
    .A(_1520_),
    .X(_1522_));
 sg13g2_xnor2_1 _4800_ (.Y(_1523_),
    .A(_1519_),
    .B(_1522_));
 sg13g2_xnor2_1 _4801_ (.Y(_1524_),
    .A(_1516_),
    .B(_1523_));
 sg13g2_nor2_1 _4802_ (.A(_1494_),
    .B(_1524_),
    .Y(_0292_));
 sg13g2_and2_1 _4803_ (.A(_1512_),
    .B(_1513_),
    .X(_1525_));
 sg13g2_or2_1 _4804_ (.X(_1526_),
    .B(_1513_),
    .A(_1512_));
 sg13g2_o21ai_1 _4805_ (.B1(_1526_),
    .Y(_1527_),
    .A1(_1511_),
    .A2(_1525_));
 sg13g2_nand2_2 _4806_ (.Y(_1528_),
    .A(net163),
    .B(_0741_));
 sg13g2_nand2_1 _4807_ (.Y(_1529_),
    .A(_0737_),
    .B(_0601_));
 sg13g2_xor2_1 _4808_ (.B(_1529_),
    .A(_1528_),
    .X(_1530_));
 sg13g2_nand2_1 _4809_ (.Y(_1531_),
    .A(_0599_),
    .B(\mem[29][3] ));
 sg13g2_xor2_1 _4810_ (.B(_1531_),
    .A(_1530_),
    .X(_1532_));
 sg13g2_xnor2_1 _4811_ (.Y(_1533_),
    .A(_1527_),
    .B(_1532_));
 sg13g2_nand2_1 _4812_ (.Y(_1534_),
    .A(_1519_),
    .B(_1516_));
 sg13g2_nor2_1 _4813_ (.A(_1519_),
    .B(_1516_),
    .Y(_1535_));
 sg13g2_a21oi_1 _4814_ (.A1(_1520_),
    .A2(_1534_),
    .Y(_1536_),
    .B1(_1535_));
 sg13g2_inv_1 _4815_ (.Y(_1537_),
    .A(_1521_));
 sg13g2_nor3_1 _4816_ (.A(_1520_),
    .B(_1537_),
    .C(_1534_),
    .Y(_1538_));
 sg13g2_a21oi_1 _4817_ (.A1(_1520_),
    .A2(_1535_),
    .Y(_1539_),
    .B1(_1538_));
 sg13g2_o21ai_1 _4818_ (.B1(_1539_),
    .Y(_1540_),
    .A1(_1521_),
    .A2(_1536_));
 sg13g2_xor2_1 _4819_ (.B(_1540_),
    .A(_1533_),
    .X(_1541_));
 sg13g2_nor2_1 _4820_ (.A(_1494_),
    .B(_1541_),
    .Y(_0293_));
 sg13g2_and2_1 _4821_ (.A(_1516_),
    .B(_1521_),
    .X(_1542_));
 sg13g2_o21ai_1 _4822_ (.B1(_1519_),
    .Y(_1543_),
    .A1(_1516_),
    .A2(_1521_));
 sg13g2_nand2b_1 _4823_ (.Y(_1544_),
    .B(_1543_),
    .A_N(_1542_));
 sg13g2_o21ai_1 _4824_ (.B1(_1519_),
    .Y(_1545_),
    .A1(_1533_),
    .A2(_1542_));
 sg13g2_o21ai_1 _4825_ (.B1(_1533_),
    .Y(_1546_),
    .A1(_1516_),
    .A2(_1521_));
 sg13g2_a21oi_1 _4826_ (.A1(_1545_),
    .A2(_1546_),
    .Y(_1547_),
    .B1(_1520_));
 sg13g2_a21oi_1 _4827_ (.A1(_1533_),
    .A2(_1544_),
    .Y(_1548_),
    .B1(_1547_));
 sg13g2_nor2_1 _4828_ (.A(_1527_),
    .B(_1530_),
    .Y(_1549_));
 sg13g2_a22oi_1 _4829_ (.Y(_1550_),
    .B1(_1527_),
    .B2(_1530_),
    .A2(net115),
    .A1(_0599_));
 sg13g2_nor2_1 _4830_ (.A(_1549_),
    .B(_1550_),
    .Y(_1551_));
 sg13g2_o21ai_1 _4831_ (.B1(_0600_),
    .Y(_1552_),
    .A1(_0737_),
    .A2(_0743_));
 sg13g2_nand3_1 _4832_ (.B(_0601_),
    .C(_1552_),
    .A(_0741_),
    .Y(_1553_));
 sg13g2_nand3_1 _4833_ (.B(_0741_),
    .C(_0601_),
    .A(_0738_),
    .Y(_1554_));
 sg13g2_nand3_1 _4834_ (.B(_0743_),
    .C(_1554_),
    .A(_0600_),
    .Y(_1555_));
 sg13g2_and2_1 _4835_ (.A(_1553_),
    .B(_1555_),
    .X(_1556_));
 sg13g2_nor2b_1 _4836_ (.A(_1551_),
    .B_N(_1556_),
    .Y(_1557_));
 sg13g2_or3_1 _4837_ (.A(_1549_),
    .B(_1550_),
    .C(_1556_),
    .X(_1558_));
 sg13g2_nand2b_1 _4838_ (.Y(_1559_),
    .B(_1558_),
    .A_N(_1557_));
 sg13g2_xnor2_1 _4839_ (.Y(_1560_),
    .A(_1548_),
    .B(_1559_));
 sg13g2_nor2_1 _4840_ (.A(_1494_),
    .B(_1560_),
    .Y(_0294_));
 sg13g2_a21oi_2 _4841_ (.B1(_1557_),
    .Y(_1561_),
    .A2(_1558_),
    .A1(_1548_));
 sg13g2_inv_1 _4842_ (.Y(_1562_),
    .A(_0601_));
 sg13g2_nor3_1 _4843_ (.A(_0738_),
    .B(net115),
    .C(_1528_),
    .Y(_1563_));
 sg13g2_a21oi_1 _4844_ (.A1(net115),
    .A2(_1528_),
    .Y(_1564_),
    .B1(_1563_));
 sg13g2_nor2_1 _4845_ (.A(_1562_),
    .B(_1564_),
    .Y(_1565_));
 sg13g2_xnor2_1 _4846_ (.Y(_1566_),
    .A(_1561_),
    .B(_1565_));
 sg13g2_nor2_1 _4847_ (.A(_1494_),
    .B(_1566_),
    .Y(_0295_));
 sg13g2_a21oi_1 _4848_ (.A1(_0737_),
    .A2(_1561_),
    .Y(_1567_),
    .B1(net115));
 sg13g2_nor2_1 _4849_ (.A(_1528_),
    .B(_1567_),
    .Y(_1568_));
 sg13g2_a21oi_1 _4850_ (.A1(net115),
    .A2(_1561_),
    .Y(_1569_),
    .B1(_1568_));
 sg13g2_nor3_1 _4851_ (.A(_1562_),
    .B(_1494_),
    .C(_1569_),
    .Y(_0296_));
 sg13g2_and3_1 _4852_ (.X(_1570_),
    .A(net174),
    .B(_0427_),
    .C(_0558_));
 sg13g2_o21ai_1 _4853_ (.B1(_1309_),
    .Y(_1571_),
    .A1(_1409_),
    .A2(_1570_));
 sg13g2_buf_2 _4854_ (.A(_1571_),
    .X(_1572_));
 sg13g2_nand2_1 _4855_ (.Y(_1573_),
    .A(net162),
    .B(net112));
 sg13g2_nor2_1 _4856_ (.A(_1572_),
    .B(_1573_),
    .Y(_0297_));
 sg13g2_nand2_1 _4857_ (.Y(_1574_),
    .A(net162),
    .B(net111));
 sg13g2_nand2_1 _4858_ (.Y(_1575_),
    .A(net112),
    .B(_0606_));
 sg13g2_xnor2_1 _4859_ (.Y(_1576_),
    .A(_1574_),
    .B(_1575_));
 sg13g2_nor2_1 _4860_ (.A(_1572_),
    .B(_1576_),
    .Y(_0298_));
 sg13g2_nand2_1 _4861_ (.Y(_1577_),
    .A(_0606_),
    .B(net111));
 sg13g2_nand2_1 _4862_ (.Y(_1578_),
    .A(net161),
    .B(_1577_));
 sg13g2_xor2_1 _4863_ (.B(net110),
    .A(net161),
    .X(_1579_));
 sg13g2_nand2_1 _4864_ (.Y(_1580_),
    .A(net162),
    .B(_1579_));
 sg13g2_o21ai_1 _4865_ (.B1(_1580_),
    .Y(_1581_),
    .A1(net162),
    .A2(_1578_));
 sg13g2_a21o_1 _4866_ (.A2(net161),
    .A1(net112),
    .B1(net162),
    .X(_1582_));
 sg13g2_o21ai_1 _4867_ (.B1(_1582_),
    .Y(_1583_),
    .A1(net112),
    .A2(net110));
 sg13g2_and2_1 _4868_ (.A(_0606_),
    .B(net111),
    .X(_1584_));
 sg13g2_buf_1 _4869_ (.A(_1584_),
    .X(_1585_));
 sg13g2_nand2_1 _4870_ (.Y(_1586_),
    .A(net162),
    .B(net110));
 sg13g2_nor3_1 _4871_ (.A(net112),
    .B(_1585_),
    .C(_1586_),
    .Y(_1587_));
 sg13g2_a221oi_1 _4872_ (.B2(_1585_),
    .C1(_1587_),
    .B1(_1583_),
    .A1(net112),
    .Y(_1588_),
    .A2(_1581_));
 sg13g2_nor2_1 _4873_ (.A(_1572_),
    .B(_1588_),
    .Y(_0299_));
 sg13g2_nand2_1 _4874_ (.Y(_1589_),
    .A(\mem[30][0] ),
    .B(_0608_));
 sg13g2_nand2_1 _4875_ (.Y(_1590_),
    .A(net111),
    .B(\mem[14][2] ));
 sg13g2_nand2_1 _4876_ (.Y(_1591_),
    .A(_0606_),
    .B(net110));
 sg13g2_xor2_1 _4877_ (.B(_1591_),
    .A(_1590_),
    .X(_1592_));
 sg13g2_xnor2_1 _4878_ (.Y(_1593_),
    .A(_1589_),
    .B(_1592_));
 sg13g2_buf_1 _4879_ (.A(_1593_),
    .X(_1594_));
 sg13g2_a21oi_1 _4880_ (.A1(_0750_),
    .A2(net161),
    .Y(_1595_),
    .B1(_1585_));
 sg13g2_nand3_1 _4881_ (.B(net161),
    .C(_1585_),
    .A(_0750_),
    .Y(_1596_));
 sg13g2_o21ai_1 _4882_ (.B1(_1596_),
    .Y(_1597_),
    .A1(_1586_),
    .A2(_1595_));
 sg13g2_buf_1 _4883_ (.A(_1597_),
    .X(_1598_));
 sg13g2_nand2_2 _4884_ (.Y(_1599_),
    .A(_0602_),
    .B(net109));
 sg13g2_nor3_2 _4885_ (.A(_1573_),
    .B(_1579_),
    .C(_1577_),
    .Y(_1600_));
 sg13g2_xor2_1 _4886_ (.B(_1600_),
    .A(_1599_),
    .X(_1601_));
 sg13g2_xnor2_1 _4887_ (.Y(_1602_),
    .A(_1598_),
    .B(_1601_));
 sg13g2_xnor2_1 _4888_ (.Y(_1603_),
    .A(_1594_),
    .B(_1602_));
 sg13g2_nor2_1 _4889_ (.A(_1572_),
    .B(_1603_),
    .Y(_0300_));
 sg13g2_and2_1 _4890_ (.A(_1590_),
    .B(_1591_),
    .X(_1604_));
 sg13g2_or2_1 _4891_ (.X(_1605_),
    .B(_1591_),
    .A(_1590_));
 sg13g2_o21ai_1 _4892_ (.B1(_1605_),
    .Y(_1606_),
    .A1(_1589_),
    .A2(_1604_));
 sg13g2_nand2_2 _4893_ (.Y(_1607_),
    .A(net161),
    .B(net110));
 sg13g2_nand2_1 _4894_ (.Y(_1608_),
    .A(net111),
    .B(_0608_));
 sg13g2_xor2_1 _4895_ (.B(_1608_),
    .A(_1607_),
    .X(_1609_));
 sg13g2_nand2_1 _4896_ (.Y(_1610_),
    .A(_0606_),
    .B(\mem[30][3] ));
 sg13g2_xor2_1 _4897_ (.B(_1610_),
    .A(_1609_),
    .X(_1611_));
 sg13g2_xnor2_1 _4898_ (.Y(_1612_),
    .A(_1606_),
    .B(_1611_));
 sg13g2_nand2_1 _4899_ (.Y(_1613_),
    .A(_1598_),
    .B(_1594_));
 sg13g2_nor2_1 _4900_ (.A(_1598_),
    .B(_1594_),
    .Y(_1614_));
 sg13g2_a21oi_1 _4901_ (.A1(_1599_),
    .A2(_1613_),
    .Y(_1615_),
    .B1(_1614_));
 sg13g2_inv_1 _4902_ (.Y(_1616_),
    .A(_1600_));
 sg13g2_nor3_1 _4903_ (.A(_1599_),
    .B(_1616_),
    .C(_1613_),
    .Y(_1617_));
 sg13g2_a21oi_1 _4904_ (.A1(_1599_),
    .A2(_1614_),
    .Y(_1618_),
    .B1(_1617_));
 sg13g2_o21ai_1 _4905_ (.B1(_1618_),
    .Y(_1619_),
    .A1(_1600_),
    .A2(_1615_));
 sg13g2_xor2_1 _4906_ (.B(_1619_),
    .A(_1612_),
    .X(_1620_));
 sg13g2_nor2_1 _4907_ (.A(_1572_),
    .B(_1620_),
    .Y(_0301_));
 sg13g2_and2_1 _4908_ (.A(_1594_),
    .B(_1600_),
    .X(_1621_));
 sg13g2_o21ai_1 _4909_ (.B1(_1598_),
    .Y(_1622_),
    .A1(_1594_),
    .A2(_1600_));
 sg13g2_nand2b_1 _4910_ (.Y(_1623_),
    .B(_1622_),
    .A_N(_1621_));
 sg13g2_o21ai_1 _4911_ (.B1(_1598_),
    .Y(_1624_),
    .A1(_1612_),
    .A2(_1621_));
 sg13g2_o21ai_1 _4912_ (.B1(_1612_),
    .Y(_1625_),
    .A1(_1594_),
    .A2(_1600_));
 sg13g2_a21oi_1 _4913_ (.A1(_1624_),
    .A2(_1625_),
    .Y(_1626_),
    .B1(_1599_));
 sg13g2_a21oi_1 _4914_ (.A1(_1612_),
    .A2(_1623_),
    .Y(_1627_),
    .B1(_1626_));
 sg13g2_nor2_1 _4915_ (.A(_1606_),
    .B(_1609_),
    .Y(_1628_));
 sg13g2_a22oi_1 _4916_ (.Y(_1629_),
    .B1(_1606_),
    .B2(_1609_),
    .A2(net109),
    .A1(_0606_));
 sg13g2_nor2_1 _4917_ (.A(_1628_),
    .B(_1629_),
    .Y(_1630_));
 sg13g2_o21ai_1 _4918_ (.B1(_0607_),
    .Y(_1631_),
    .A1(net111),
    .A2(net109));
 sg13g2_nand3_1 _4919_ (.B(_0608_),
    .C(_1631_),
    .A(net110),
    .Y(_1632_));
 sg13g2_nand3_1 _4920_ (.B(_0755_),
    .C(_0608_),
    .A(_0753_),
    .Y(_1633_));
 sg13g2_nand3_1 _4921_ (.B(net109),
    .C(_1633_),
    .A(_0607_),
    .Y(_1634_));
 sg13g2_and2_1 _4922_ (.A(_1632_),
    .B(_1634_),
    .X(_1635_));
 sg13g2_nor2b_1 _4923_ (.A(_1630_),
    .B_N(_1635_),
    .Y(_1636_));
 sg13g2_or3_1 _4924_ (.A(_1628_),
    .B(_1629_),
    .C(_1635_),
    .X(_1637_));
 sg13g2_nand2b_1 _4925_ (.Y(_1638_),
    .B(_1637_),
    .A_N(_1636_));
 sg13g2_xnor2_1 _4926_ (.Y(_1639_),
    .A(_1627_),
    .B(_1638_));
 sg13g2_nor2_1 _4927_ (.A(_1572_),
    .B(_1639_),
    .Y(_0302_));
 sg13g2_a21oi_2 _4928_ (.B1(_1636_),
    .Y(_1640_),
    .A2(_1637_),
    .A1(_1627_));
 sg13g2_inv_1 _4929_ (.Y(_1641_),
    .A(_0608_));
 sg13g2_nor3_1 _4930_ (.A(_0753_),
    .B(net109),
    .C(_1607_),
    .Y(_1642_));
 sg13g2_a21oi_1 _4931_ (.A1(net109),
    .A2(_1607_),
    .Y(_1643_),
    .B1(_1642_));
 sg13g2_nor2_1 _4932_ (.A(_1641_),
    .B(_1643_),
    .Y(_1644_));
 sg13g2_xnor2_1 _4933_ (.Y(_1645_),
    .A(_1640_),
    .B(_1644_));
 sg13g2_nor2_1 _4934_ (.A(_1572_),
    .B(_1645_),
    .Y(_0303_));
 sg13g2_a21oi_1 _4935_ (.A1(_0752_),
    .A2(_1640_),
    .Y(_1646_),
    .B1(_0756_));
 sg13g2_nor2_1 _4936_ (.A(_1607_),
    .B(_1646_),
    .Y(_1647_));
 sg13g2_a21oi_1 _4937_ (.A1(_0756_),
    .A2(_1640_),
    .Y(_1648_),
    .B1(_1647_));
 sg13g2_nor3_1 _4938_ (.A(_1641_),
    .B(_1572_),
    .C(_1648_),
    .Y(_0304_));
 sg13g2_or2_1 _4939_ (.X(_1649_),
    .B(_0557_),
    .A(net173));
 sg13g2_o21ai_1 _4940_ (.B1(_1649_),
    .Y(_1650_),
    .A1(_1313_),
    .A2(_1410_));
 sg13g2_o21ai_1 _4941_ (.B1(net175),
    .Y(_1651_),
    .A1(_1313_),
    .A2(_1410_));
 sg13g2_nand4_1 _4942_ (.B(_1315_),
    .C(_1650_),
    .A(net57),
    .Y(_1652_),
    .D(_1651_));
 sg13g2_buf_2 _4943_ (.A(_1652_),
    .X(_1653_));
 sg13g2_nand2_1 _4944_ (.Y(_1654_),
    .A(net160),
    .B(net108));
 sg13g2_nor2_1 _4945_ (.A(_1653_),
    .B(_1654_),
    .Y(_0305_));
 sg13g2_nand2_1 _4946_ (.Y(_1655_),
    .A(net160),
    .B(net107));
 sg13g2_nand2_1 _4947_ (.Y(_1656_),
    .A(net108),
    .B(_0613_));
 sg13g2_xnor2_1 _4948_ (.Y(_1657_),
    .A(_1655_),
    .B(_1656_));
 sg13g2_nor2_1 _4949_ (.A(_1653_),
    .B(_1657_),
    .Y(_0306_));
 sg13g2_nand2_1 _4950_ (.Y(_1658_),
    .A(_0613_),
    .B(net107));
 sg13g2_nand2_1 _4951_ (.Y(_1659_),
    .A(net159),
    .B(_1658_));
 sg13g2_xor2_1 _4952_ (.B(net106),
    .A(net159),
    .X(_1660_));
 sg13g2_nand2_1 _4953_ (.Y(_1661_),
    .A(net160),
    .B(_1660_));
 sg13g2_o21ai_1 _4954_ (.B1(_1661_),
    .Y(_1662_),
    .A1(net160),
    .A2(_1659_));
 sg13g2_a21o_1 _4955_ (.A2(net159),
    .A1(net108),
    .B1(net160),
    .X(_1663_));
 sg13g2_o21ai_1 _4956_ (.B1(_1663_),
    .Y(_1664_),
    .A1(net108),
    .A2(net106));
 sg13g2_and2_1 _4957_ (.A(_0613_),
    .B(net107),
    .X(_1665_));
 sg13g2_buf_1 _4958_ (.A(_1665_),
    .X(_1666_));
 sg13g2_nand2_1 _4959_ (.Y(_1667_),
    .A(net160),
    .B(_0762_));
 sg13g2_nor3_1 _4960_ (.A(net108),
    .B(_1666_),
    .C(_1667_),
    .Y(_1668_));
 sg13g2_a221oi_1 _4961_ (.B2(_1666_),
    .C1(_1668_),
    .B1(_1664_),
    .A1(net108),
    .Y(_1669_),
    .A2(_1662_));
 sg13g2_nor2_1 _4962_ (.A(_1653_),
    .B(_1669_),
    .Y(_0307_));
 sg13g2_nand2_1 _4963_ (.Y(_1670_),
    .A(\mem[31][0] ),
    .B(_0615_));
 sg13g2_nand2_1 _4964_ (.Y(_1671_),
    .A(net107),
    .B(\mem[15][2] ));
 sg13g2_nand2_1 _4965_ (.Y(_1672_),
    .A(_0613_),
    .B(net106));
 sg13g2_xor2_1 _4966_ (.B(_1672_),
    .A(_1671_),
    .X(_1673_));
 sg13g2_xnor2_1 _4967_ (.Y(_1674_),
    .A(_1670_),
    .B(_1673_));
 sg13g2_buf_1 _4968_ (.A(_1674_),
    .X(_1675_));
 sg13g2_a21oi_1 _4969_ (.A1(_0757_),
    .A2(_0614_),
    .Y(_1676_),
    .B1(_1666_));
 sg13g2_nand3_1 _4970_ (.B(_0614_),
    .C(_1666_),
    .A(_0757_),
    .Y(_1677_));
 sg13g2_o21ai_1 _4971_ (.B1(_1677_),
    .Y(_1678_),
    .A1(_1667_),
    .A2(_1676_));
 sg13g2_buf_1 _4972_ (.A(_1678_),
    .X(_1679_));
 sg13g2_nand2_2 _4973_ (.Y(_1680_),
    .A(_0609_),
    .B(_0763_));
 sg13g2_nor3_2 _4974_ (.A(_1654_),
    .B(_1660_),
    .C(_1658_),
    .Y(_1681_));
 sg13g2_xor2_1 _4975_ (.B(_1681_),
    .A(_1680_),
    .X(_1682_));
 sg13g2_xnor2_1 _4976_ (.Y(_1683_),
    .A(_1679_),
    .B(_1682_));
 sg13g2_xnor2_1 _4977_ (.Y(_1684_),
    .A(_1675_),
    .B(_1683_));
 sg13g2_nor2_1 _4978_ (.A(_1653_),
    .B(_1684_),
    .Y(_0308_));
 sg13g2_and2_1 _4979_ (.A(_1671_),
    .B(_1672_),
    .X(_1685_));
 sg13g2_or2_1 _4980_ (.X(_1686_),
    .B(_1672_),
    .A(_1671_));
 sg13g2_o21ai_1 _4981_ (.B1(_1686_),
    .Y(_1687_),
    .A1(_1670_),
    .A2(_1685_));
 sg13g2_nand2_2 _4982_ (.Y(_1688_),
    .A(net159),
    .B(net106));
 sg13g2_nand2_1 _4983_ (.Y(_1689_),
    .A(net107),
    .B(_0615_));
 sg13g2_xor2_1 _4984_ (.B(_1689_),
    .A(_1688_),
    .X(_1690_));
 sg13g2_nand2_1 _4985_ (.Y(_1691_),
    .A(_0613_),
    .B(\mem[31][3] ));
 sg13g2_xor2_1 _4986_ (.B(_1691_),
    .A(_1690_),
    .X(_1692_));
 sg13g2_xnor2_1 _4987_ (.Y(_1693_),
    .A(_1687_),
    .B(_1692_));
 sg13g2_nand2_1 _4988_ (.Y(_1694_),
    .A(_1679_),
    .B(_1675_));
 sg13g2_nor2_1 _4989_ (.A(_1679_),
    .B(_1675_),
    .Y(_1695_));
 sg13g2_a21oi_1 _4990_ (.A1(_1680_),
    .A2(_1694_),
    .Y(_1696_),
    .B1(_1695_));
 sg13g2_inv_1 _4991_ (.Y(_1697_),
    .A(_1681_));
 sg13g2_nor3_1 _4992_ (.A(_1680_),
    .B(_1697_),
    .C(_1694_),
    .Y(_1698_));
 sg13g2_a21oi_1 _4993_ (.A1(_1680_),
    .A2(_1695_),
    .Y(_1699_),
    .B1(_1698_));
 sg13g2_o21ai_1 _4994_ (.B1(_1699_),
    .Y(_1700_),
    .A1(_1681_),
    .A2(_1696_));
 sg13g2_xor2_1 _4995_ (.B(_1700_),
    .A(_1693_),
    .X(_1701_));
 sg13g2_nor2_1 _4996_ (.A(_1653_),
    .B(_1701_),
    .Y(_0309_));
 sg13g2_and2_1 _4997_ (.A(_1675_),
    .B(_1681_),
    .X(_1702_));
 sg13g2_o21ai_1 _4998_ (.B1(_1679_),
    .Y(_1703_),
    .A1(_1675_),
    .A2(_1681_));
 sg13g2_nand2b_1 _4999_ (.Y(_1704_),
    .B(_1703_),
    .A_N(_1702_));
 sg13g2_o21ai_1 _5000_ (.B1(_1679_),
    .Y(_1705_),
    .A1(_1693_),
    .A2(_1702_));
 sg13g2_o21ai_1 _5001_ (.B1(_1693_),
    .Y(_1706_),
    .A1(_1675_),
    .A2(_1681_));
 sg13g2_a21oi_1 _5002_ (.A1(_1705_),
    .A2(_1706_),
    .Y(_1707_),
    .B1(_1680_));
 sg13g2_a21oi_1 _5003_ (.A1(_1693_),
    .A2(_1704_),
    .Y(_1708_),
    .B1(_1707_));
 sg13g2_nor2_1 _5004_ (.A(_1687_),
    .B(_1690_),
    .Y(_1709_));
 sg13g2_a22oi_1 _5005_ (.Y(_1710_),
    .B1(_1687_),
    .B2(_1690_),
    .A2(net105),
    .A1(_0613_));
 sg13g2_nor2_1 _5006_ (.A(_1709_),
    .B(_1710_),
    .Y(_1711_));
 sg13g2_o21ai_1 _5007_ (.B1(net159),
    .Y(_1712_),
    .A1(net107),
    .A2(net105));
 sg13g2_nand3_1 _5008_ (.B(_0615_),
    .C(_1712_),
    .A(net106),
    .Y(_1713_));
 sg13g2_nand3_1 _5009_ (.B(net106),
    .C(_0615_),
    .A(_0760_),
    .Y(_1714_));
 sg13g2_nand3_1 _5010_ (.B(net105),
    .C(_1714_),
    .A(net159),
    .Y(_1715_));
 sg13g2_and2_1 _5011_ (.A(_1713_),
    .B(_1715_),
    .X(_1716_));
 sg13g2_nor2b_1 _5012_ (.A(_1711_),
    .B_N(_1716_),
    .Y(_1717_));
 sg13g2_or3_1 _5013_ (.A(_1709_),
    .B(_1710_),
    .C(_1716_),
    .X(_1718_));
 sg13g2_nand2b_1 _5014_ (.Y(_1719_),
    .B(_1718_),
    .A_N(_1717_));
 sg13g2_xnor2_1 _5015_ (.Y(_1720_),
    .A(_1708_),
    .B(_1719_));
 sg13g2_nor2_1 _5016_ (.A(_1653_),
    .B(_1720_),
    .Y(_0310_));
 sg13g2_a21oi_2 _5017_ (.B1(_1717_),
    .Y(_1721_),
    .A2(_1718_),
    .A1(_1708_));
 sg13g2_inv_1 _5018_ (.Y(_1722_),
    .A(_0615_));
 sg13g2_nor3_1 _5019_ (.A(_0760_),
    .B(net105),
    .C(_1688_),
    .Y(_1723_));
 sg13g2_a21oi_1 _5020_ (.A1(net105),
    .A2(_1688_),
    .Y(_1724_),
    .B1(_1723_));
 sg13g2_nor2_1 _5021_ (.A(_1722_),
    .B(_1724_),
    .Y(_1725_));
 sg13g2_xnor2_1 _5022_ (.Y(_1726_),
    .A(_1721_),
    .B(_1725_));
 sg13g2_nor2_1 _5023_ (.A(_1653_),
    .B(_1726_),
    .Y(_0311_));
 sg13g2_a21oi_1 _5024_ (.A1(net107),
    .A2(_1721_),
    .Y(_1727_),
    .B1(net105));
 sg13g2_nor2_1 _5025_ (.A(_1688_),
    .B(_1727_),
    .Y(_1728_));
 sg13g2_a21oi_1 _5026_ (.A1(net105),
    .A2(_1721_),
    .Y(_1729_),
    .B1(_1728_));
 sg13g2_nor3_1 _5027_ (.A(_1722_),
    .B(_1653_),
    .C(_1729_),
    .Y(_0312_));
 sg13g2_nand2_1 _5028_ (.Y(_1730_),
    .A(net158),
    .B(net104));
 sg13g2_nor2_1 _5029_ (.A(net56),
    .B(_1730_),
    .Y(_0313_));
 sg13g2_nand2_1 _5030_ (.Y(_1731_),
    .A(net158),
    .B(net103));
 sg13g2_nand2_1 _5031_ (.Y(_1732_),
    .A(net104),
    .B(_0621_));
 sg13g2_xnor2_1 _5032_ (.Y(_1733_),
    .A(_1731_),
    .B(_1732_));
 sg13g2_nor2_1 _5033_ (.A(net56),
    .B(_1733_),
    .Y(_0314_));
 sg13g2_nand2_1 _5034_ (.Y(_1734_),
    .A(_0621_),
    .B(net103));
 sg13g2_nand2_1 _5035_ (.Y(_1735_),
    .A(_0622_),
    .B(_1734_));
 sg13g2_xor2_1 _5036_ (.B(net102),
    .A(net157),
    .X(_1736_));
 sg13g2_nand2_1 _5037_ (.Y(_1737_),
    .A(net158),
    .B(_1736_));
 sg13g2_o21ai_1 _5038_ (.B1(_1737_),
    .Y(_1738_),
    .A1(net158),
    .A2(_1735_));
 sg13g2_a21o_1 _5039_ (.A2(_0622_),
    .A1(net104),
    .B1(net158),
    .X(_1739_));
 sg13g2_o21ai_1 _5040_ (.B1(_1739_),
    .Y(_1740_),
    .A1(net104),
    .A2(net102));
 sg13g2_and2_1 _5041_ (.A(_0621_),
    .B(net103),
    .X(_1741_));
 sg13g2_buf_1 _5042_ (.A(_1741_),
    .X(_1742_));
 sg13g2_nand2_1 _5043_ (.Y(_1743_),
    .A(net158),
    .B(net102));
 sg13g2_nor3_1 _5044_ (.A(net104),
    .B(_1742_),
    .C(_1743_),
    .Y(_1744_));
 sg13g2_a221oi_1 _5045_ (.B2(_1742_),
    .C1(_1744_),
    .B1(_1740_),
    .A1(net104),
    .Y(_1745_),
    .A2(_1738_));
 sg13g2_nor2_1 _5046_ (.A(net56),
    .B(_1745_),
    .Y(_0315_));
 sg13g2_nand2_1 _5047_ (.Y(_1746_),
    .A(\mem[32][0] ),
    .B(_0623_));
 sg13g2_nand2_1 _5048_ (.Y(_1747_),
    .A(net103),
    .B(\mem[16][2] ));
 sg13g2_nand2_1 _5049_ (.Y(_1748_),
    .A(_0621_),
    .B(net102));
 sg13g2_xor2_1 _5050_ (.B(_1748_),
    .A(_1747_),
    .X(_1749_));
 sg13g2_xnor2_1 _5051_ (.Y(_1750_),
    .A(_1746_),
    .B(_1749_));
 sg13g2_buf_1 _5052_ (.A(_1750_),
    .X(_1751_));
 sg13g2_a21oi_1 _5053_ (.A1(_0764_),
    .A2(net157),
    .Y(_1752_),
    .B1(_1742_));
 sg13g2_nand3_1 _5054_ (.B(net157),
    .C(_1742_),
    .A(_0764_),
    .Y(_1753_));
 sg13g2_o21ai_1 _5055_ (.B1(_1753_),
    .Y(_1754_),
    .A1(_1743_),
    .A2(_1752_));
 sg13g2_buf_1 _5056_ (.A(_1754_),
    .X(_1755_));
 sg13g2_nand2_2 _5057_ (.Y(_1756_),
    .A(_0616_),
    .B(net101));
 sg13g2_nor3_2 _5058_ (.A(_1730_),
    .B(_1736_),
    .C(_1734_),
    .Y(_1757_));
 sg13g2_xor2_1 _5059_ (.B(_1757_),
    .A(_1756_),
    .X(_1758_));
 sg13g2_xnor2_1 _5060_ (.Y(_1759_),
    .A(_1755_),
    .B(_1758_));
 sg13g2_xnor2_1 _5061_ (.Y(_1760_),
    .A(_1751_),
    .B(_1759_));
 sg13g2_nor2_1 _5062_ (.A(net56),
    .B(_1760_),
    .Y(_0316_));
 sg13g2_and2_1 _5063_ (.A(_1747_),
    .B(_1748_),
    .X(_1761_));
 sg13g2_or2_1 _5064_ (.X(_1762_),
    .B(_1748_),
    .A(_1747_));
 sg13g2_o21ai_1 _5065_ (.B1(_1762_),
    .Y(_1763_),
    .A1(_1746_),
    .A2(_1761_));
 sg13g2_nand2_2 _5066_ (.Y(_1764_),
    .A(net157),
    .B(net102));
 sg13g2_nand2_1 _5067_ (.Y(_1765_),
    .A(net103),
    .B(_0623_));
 sg13g2_xor2_1 _5068_ (.B(_1765_),
    .A(_1764_),
    .X(_1766_));
 sg13g2_nand2_1 _5069_ (.Y(_1767_),
    .A(_0621_),
    .B(\mem[32][3] ));
 sg13g2_xor2_1 _5070_ (.B(_1767_),
    .A(_1766_),
    .X(_1768_));
 sg13g2_xnor2_1 _5071_ (.Y(_1769_),
    .A(_1763_),
    .B(_1768_));
 sg13g2_nand2_1 _5072_ (.Y(_1770_),
    .A(_1755_),
    .B(_1751_));
 sg13g2_nor2_1 _5073_ (.A(_1755_),
    .B(_1751_),
    .Y(_1771_));
 sg13g2_a21oi_1 _5074_ (.A1(_1756_),
    .A2(_1770_),
    .Y(_1772_),
    .B1(_1771_));
 sg13g2_inv_1 _5075_ (.Y(_1773_),
    .A(_1757_));
 sg13g2_nor3_1 _5076_ (.A(_1756_),
    .B(_1773_),
    .C(_1770_),
    .Y(_1774_));
 sg13g2_a21oi_1 _5077_ (.A1(_1756_),
    .A2(_1771_),
    .Y(_1775_),
    .B1(_1774_));
 sg13g2_o21ai_1 _5078_ (.B1(_1775_),
    .Y(_1776_),
    .A1(_1757_),
    .A2(_1772_));
 sg13g2_xor2_1 _5079_ (.B(_1776_),
    .A(_1769_),
    .X(_1777_));
 sg13g2_nor2_1 _5080_ (.A(net56),
    .B(_1777_),
    .Y(_0317_));
 sg13g2_and2_1 _5081_ (.A(_1751_),
    .B(_1757_),
    .X(_1778_));
 sg13g2_o21ai_1 _5082_ (.B1(_1755_),
    .Y(_1779_),
    .A1(_1751_),
    .A2(_1757_));
 sg13g2_nand2b_1 _5083_ (.Y(_1780_),
    .B(_1779_),
    .A_N(_1778_));
 sg13g2_o21ai_1 _5084_ (.B1(_1755_),
    .Y(_1781_),
    .A1(_1769_),
    .A2(_1778_));
 sg13g2_o21ai_1 _5085_ (.B1(_1769_),
    .Y(_1782_),
    .A1(_1751_),
    .A2(_1757_));
 sg13g2_a21oi_1 _5086_ (.A1(_1781_),
    .A2(_1782_),
    .Y(_1783_),
    .B1(_1756_));
 sg13g2_a21oi_1 _5087_ (.A1(_1769_),
    .A2(_1780_),
    .Y(_1784_),
    .B1(_1783_));
 sg13g2_nor2_1 _5088_ (.A(_1763_),
    .B(_1766_),
    .Y(_1785_));
 sg13g2_a22oi_1 _5089_ (.Y(_1786_),
    .B1(_1763_),
    .B2(_1766_),
    .A2(net101),
    .A1(_0621_));
 sg13g2_nor2_1 _5090_ (.A(_1785_),
    .B(_1786_),
    .Y(_1787_));
 sg13g2_o21ai_1 _5091_ (.B1(net157),
    .Y(_1788_),
    .A1(net103),
    .A2(net101));
 sg13g2_nand3_1 _5092_ (.B(_0623_),
    .C(_1788_),
    .A(net102),
    .Y(_1789_));
 sg13g2_nand3_1 _5093_ (.B(_0773_),
    .C(_0623_),
    .A(_0771_),
    .Y(_1790_));
 sg13g2_nand3_1 _5094_ (.B(net101),
    .C(_1790_),
    .A(net157),
    .Y(_1791_));
 sg13g2_and2_1 _5095_ (.A(_1789_),
    .B(_1791_),
    .X(_1792_));
 sg13g2_nor2b_1 _5096_ (.A(_1787_),
    .B_N(_1792_),
    .Y(_1793_));
 sg13g2_or3_1 _5097_ (.A(_1785_),
    .B(_1786_),
    .C(_1792_),
    .X(_1794_));
 sg13g2_nand2b_1 _5098_ (.Y(_1795_),
    .B(_1794_),
    .A_N(_1793_));
 sg13g2_xnor2_1 _5099_ (.Y(_1796_),
    .A(_1784_),
    .B(_1795_));
 sg13g2_nor2_1 _5100_ (.A(net56),
    .B(_1796_),
    .Y(_0318_));
 sg13g2_a21oi_2 _5101_ (.B1(_1793_),
    .Y(_1797_),
    .A2(_1794_),
    .A1(_1784_));
 sg13g2_inv_1 _5102_ (.Y(_1798_),
    .A(_0623_));
 sg13g2_nor3_1 _5103_ (.A(_0771_),
    .B(net101),
    .C(_1764_),
    .Y(_1799_));
 sg13g2_a21oi_1 _5104_ (.A1(net101),
    .A2(_1764_),
    .Y(_1800_),
    .B1(_1799_));
 sg13g2_nor2_1 _5105_ (.A(_1798_),
    .B(_1800_),
    .Y(_1801_));
 sg13g2_xnor2_1 _5106_ (.Y(_1802_),
    .A(_1797_),
    .B(_1801_));
 sg13g2_nor2_1 _5107_ (.A(net56),
    .B(_1802_),
    .Y(_0319_));
 sg13g2_a21oi_1 _5108_ (.A1(_0770_),
    .A2(_1797_),
    .Y(_1803_),
    .B1(_0774_));
 sg13g2_nor2_1 _5109_ (.A(_1764_),
    .B(_1803_),
    .Y(_1804_));
 sg13g2_a21oi_1 _5110_ (.A1(_0774_),
    .A2(_1797_),
    .Y(_1805_),
    .B1(_1804_));
 sg13g2_nor3_1 _5111_ (.A(_1798_),
    .B(net56),
    .C(_1805_),
    .Y(_0320_));
 sg13g2_o21ai_1 _5112_ (.B1(_1308_),
    .Y(_1806_),
    .A1(_1490_),
    .A2(_1649_));
 sg13g2_buf_1 _5113_ (.A(_1806_),
    .X(_1807_));
 sg13g2_nand2b_1 _5114_ (.Y(_1808_),
    .B(net57),
    .A_N(_1313_));
 sg13g2_and2_1 _5115_ (.A(net55),
    .B(_1808_),
    .X(_1809_));
 sg13g2_buf_2 _5116_ (.A(_1809_),
    .X(_1810_));
 sg13g2_nand2_1 _5117_ (.Y(_1811_),
    .A(net114),
    .B(net152));
 sg13g2_nor2_1 _5118_ (.A(_1810_),
    .B(_1811_),
    .Y(_0321_));
 sg13g2_nand2_1 _5119_ (.Y(_1812_),
    .A(net114),
    .B(net151));
 sg13g2_nand2_1 _5120_ (.Y(_1813_),
    .A(net152),
    .B(_0746_));
 sg13g2_xnor2_1 _5121_ (.Y(_1814_),
    .A(_1812_),
    .B(_1813_));
 sg13g2_nor2_1 _5122_ (.A(_1810_),
    .B(_1814_),
    .Y(_0322_));
 sg13g2_nand2_1 _5123_ (.Y(_1815_),
    .A(_0746_),
    .B(net151));
 sg13g2_nand2_1 _5124_ (.Y(_1816_),
    .A(net113),
    .B(_1815_));
 sg13g2_xor2_1 _5125_ (.B(net150),
    .A(net113),
    .X(_1817_));
 sg13g2_nand2_1 _5126_ (.Y(_1818_),
    .A(net114),
    .B(_1817_));
 sg13g2_o21ai_1 _5127_ (.B1(_1818_),
    .Y(_1819_),
    .A1(net114),
    .A2(_1816_));
 sg13g2_a21o_1 _5128_ (.A2(net113),
    .A1(net152),
    .B1(net114),
    .X(_1820_));
 sg13g2_o21ai_1 _5129_ (.B1(_1820_),
    .Y(_1821_),
    .A1(net152),
    .A2(net150));
 sg13g2_and2_1 _5130_ (.A(_0746_),
    .B(net151),
    .X(_1822_));
 sg13g2_buf_1 _5131_ (.A(_1822_),
    .X(_1823_));
 sg13g2_nand2_1 _5132_ (.Y(_1824_),
    .A(net114),
    .B(net150));
 sg13g2_nor3_1 _5133_ (.A(net152),
    .B(_1823_),
    .C(_1824_),
    .Y(_1825_));
 sg13g2_a221oi_1 _5134_ (.B2(_1823_),
    .C1(_1825_),
    .B1(_1821_),
    .A1(net152),
    .Y(_1826_),
    .A2(_1819_));
 sg13g2_nor2_1 _5135_ (.A(_1810_),
    .B(_1826_),
    .Y(_0323_));
 sg13g2_nand2_1 _5136_ (.Y(_1827_),
    .A(\mem[18][0] ),
    .B(_0748_));
 sg13g2_nand2_1 _5137_ (.Y(_1828_),
    .A(net151),
    .B(\mem[2][2] ));
 sg13g2_nand2_1 _5138_ (.Y(_1829_),
    .A(_0746_),
    .B(net150));
 sg13g2_xor2_1 _5139_ (.B(_1829_),
    .A(_1828_),
    .X(_1830_));
 sg13g2_xnor2_1 _5140_ (.Y(_1831_),
    .A(_1827_),
    .B(_1830_));
 sg13g2_buf_1 _5141_ (.A(_1831_),
    .X(_1832_));
 sg13g2_a21oi_1 _5142_ (.A1(_0637_),
    .A2(net113),
    .Y(_1833_),
    .B1(_1823_));
 sg13g2_nand3_1 _5143_ (.B(net113),
    .C(_1823_),
    .A(_0637_),
    .Y(_1834_));
 sg13g2_o21ai_1 _5144_ (.B1(_1834_),
    .Y(_1835_),
    .A1(_1824_),
    .A2(_1833_));
 sg13g2_buf_1 _5145_ (.A(_1835_),
    .X(_1836_));
 sg13g2_nand2_2 _5146_ (.Y(_1837_),
    .A(_0744_),
    .B(net149));
 sg13g2_nor3_2 _5147_ (.A(_1811_),
    .B(_1817_),
    .C(_1815_),
    .Y(_1838_));
 sg13g2_xor2_1 _5148_ (.B(_1838_),
    .A(_1837_),
    .X(_1839_));
 sg13g2_xnor2_1 _5149_ (.Y(_1840_),
    .A(_1836_),
    .B(_1839_));
 sg13g2_xnor2_1 _5150_ (.Y(_1841_),
    .A(_1832_),
    .B(_1840_));
 sg13g2_nor2_1 _5151_ (.A(_1810_),
    .B(_1841_),
    .Y(_0324_));
 sg13g2_and2_1 _5152_ (.A(_1828_),
    .B(_1829_),
    .X(_1842_));
 sg13g2_or2_1 _5153_ (.X(_1843_),
    .B(_1829_),
    .A(_1828_));
 sg13g2_o21ai_1 _5154_ (.B1(_1843_),
    .Y(_1844_),
    .A1(_1827_),
    .A2(_1842_));
 sg13g2_nand2_2 _5155_ (.Y(_1845_),
    .A(_0747_),
    .B(_0642_));
 sg13g2_nand2_1 _5156_ (.Y(_1846_),
    .A(net151),
    .B(_0748_));
 sg13g2_xor2_1 _5157_ (.B(_1846_),
    .A(_1845_),
    .X(_1847_));
 sg13g2_nand2_1 _5158_ (.Y(_1848_),
    .A(_0746_),
    .B(\mem[18][3] ));
 sg13g2_xor2_1 _5159_ (.B(_1848_),
    .A(_1847_),
    .X(_1849_));
 sg13g2_xnor2_1 _5160_ (.Y(_1850_),
    .A(_1844_),
    .B(_1849_));
 sg13g2_nand2_1 _5161_ (.Y(_1851_),
    .A(_1836_),
    .B(_1832_));
 sg13g2_nor2_1 _5162_ (.A(_1836_),
    .B(_1832_),
    .Y(_1852_));
 sg13g2_a21oi_1 _5163_ (.A1(_1837_),
    .A2(_1851_),
    .Y(_1853_),
    .B1(_1852_));
 sg13g2_inv_1 _5164_ (.Y(_1854_),
    .A(_1838_));
 sg13g2_nor3_1 _5165_ (.A(_1837_),
    .B(_1854_),
    .C(_1851_),
    .Y(_1855_));
 sg13g2_a21oi_1 _5166_ (.A1(_1837_),
    .A2(_1852_),
    .Y(_1856_),
    .B1(_1855_));
 sg13g2_o21ai_1 _5167_ (.B1(_1856_),
    .Y(_1857_),
    .A1(_1838_),
    .A2(_1853_));
 sg13g2_xor2_1 _5168_ (.B(_1857_),
    .A(_1850_),
    .X(_1858_));
 sg13g2_nor2_1 _5169_ (.A(_1810_),
    .B(_1858_),
    .Y(_0325_));
 sg13g2_and2_1 _5170_ (.A(_1832_),
    .B(_1838_),
    .X(_1859_));
 sg13g2_o21ai_1 _5171_ (.B1(_1836_),
    .Y(_1860_),
    .A1(_1832_),
    .A2(_1838_));
 sg13g2_nand2b_1 _5172_ (.Y(_1861_),
    .B(_1860_),
    .A_N(_1859_));
 sg13g2_o21ai_1 _5173_ (.B1(_1836_),
    .Y(_1862_),
    .A1(_1850_),
    .A2(_1859_));
 sg13g2_o21ai_1 _5174_ (.B1(_1850_),
    .Y(_1863_),
    .A1(_1832_),
    .A2(_1838_));
 sg13g2_a21oi_1 _5175_ (.A1(_1862_),
    .A2(_1863_),
    .Y(_1864_),
    .B1(_1837_));
 sg13g2_a21oi_1 _5176_ (.A1(_1850_),
    .A2(_1861_),
    .Y(_1865_),
    .B1(_1864_));
 sg13g2_nor2_1 _5177_ (.A(_1844_),
    .B(_1847_),
    .Y(_1866_));
 sg13g2_a22oi_1 _5178_ (.Y(_1867_),
    .B1(_1844_),
    .B2(_1847_),
    .A2(net149),
    .A1(_0746_));
 sg13g2_nor2_1 _5179_ (.A(_1866_),
    .B(_1867_),
    .Y(_1868_));
 sg13g2_o21ai_1 _5180_ (.B1(_0747_),
    .Y(_1869_),
    .A1(net151),
    .A2(net149));
 sg13g2_nand3_1 _5181_ (.B(_0748_),
    .C(_1869_),
    .A(net150),
    .Y(_1870_));
 sg13g2_nand3_1 _5182_ (.B(net150),
    .C(_0748_),
    .A(_0640_),
    .Y(_1871_));
 sg13g2_nand3_1 _5183_ (.B(net149),
    .C(_1871_),
    .A(net113),
    .Y(_1872_));
 sg13g2_and2_1 _5184_ (.A(_1870_),
    .B(_1872_),
    .X(_1873_));
 sg13g2_nor2b_1 _5185_ (.A(_1868_),
    .B_N(_1873_),
    .Y(_1874_));
 sg13g2_or3_1 _5186_ (.A(_1866_),
    .B(_1867_),
    .C(_1873_),
    .X(_1875_));
 sg13g2_nand2b_1 _5187_ (.Y(_1876_),
    .B(_1875_),
    .A_N(_1874_));
 sg13g2_xnor2_1 _5188_ (.Y(_1877_),
    .A(_1865_),
    .B(_1876_));
 sg13g2_nor2_1 _5189_ (.A(_1810_),
    .B(_1877_),
    .Y(_0326_));
 sg13g2_a21oi_2 _5190_ (.B1(_1874_),
    .Y(_1878_),
    .A2(_1875_),
    .A1(_1865_));
 sg13g2_inv_1 _5191_ (.Y(_1879_),
    .A(_0748_));
 sg13g2_nor3_1 _5192_ (.A(_0640_),
    .B(net149),
    .C(_1845_),
    .Y(_1880_));
 sg13g2_a21oi_1 _5193_ (.A1(net149),
    .A2(_1845_),
    .Y(_1881_),
    .B1(_1880_));
 sg13g2_nor2_1 _5194_ (.A(_1879_),
    .B(_1881_),
    .Y(_1882_));
 sg13g2_xnor2_1 _5195_ (.Y(_1883_),
    .A(_1878_),
    .B(_1882_));
 sg13g2_nor2_1 _5196_ (.A(_1810_),
    .B(_1883_),
    .Y(_0327_));
 sg13g2_a21oi_1 _5197_ (.A1(_0639_),
    .A2(_1878_),
    .Y(_1884_),
    .B1(_0643_));
 sg13g2_nor2_1 _5198_ (.A(_1845_),
    .B(_1884_),
    .Y(_1885_));
 sg13g2_a21oi_1 _5199_ (.A1(_0643_),
    .A2(_1878_),
    .Y(_1886_),
    .B1(_1885_));
 sg13g2_nor3_1 _5200_ (.A(_1879_),
    .B(_1810_),
    .C(_1886_),
    .Y(_0328_));
 sg13g2_nand3_1 _5201_ (.B(net174),
    .C(net57),
    .A(net175),
    .Y(_1887_));
 sg13g2_and2_1 _5202_ (.A(_1806_),
    .B(_1887_),
    .X(_1888_));
 sg13g2_buf_2 _5203_ (.A(_1888_),
    .X(_1889_));
 sg13g2_nand2_1 _5204_ (.Y(_1890_),
    .A(net100),
    .B(net148));
 sg13g2_nor2_1 _5205_ (.A(_1889_),
    .B(_1890_),
    .Y(_0329_));
 sg13g2_nand2_1 _5206_ (.Y(_1891_),
    .A(net100),
    .B(net147));
 sg13g2_nand2_1 _5207_ (.Y(_1892_),
    .A(net148),
    .B(_1139_));
 sg13g2_xnor2_1 _5208_ (.Y(_1893_),
    .A(_1891_),
    .B(_1892_));
 sg13g2_nor2_1 _5209_ (.A(_1889_),
    .B(_1893_),
    .Y(_0330_));
 sg13g2_nand2_1 _5210_ (.Y(_1894_),
    .A(_1139_),
    .B(net147));
 sg13g2_nand2_1 _5211_ (.Y(_1895_),
    .A(net99),
    .B(_1894_));
 sg13g2_xor2_1 _5212_ (.B(net146),
    .A(net99),
    .X(_1896_));
 sg13g2_nand2_1 _5213_ (.Y(_1897_),
    .A(net100),
    .B(_1896_));
 sg13g2_o21ai_1 _5214_ (.B1(_1897_),
    .Y(_1898_),
    .A1(net100),
    .A2(_1895_));
 sg13g2_a21o_1 _5215_ (.A2(net99),
    .A1(net148),
    .B1(net100),
    .X(_1899_));
 sg13g2_o21ai_1 _5216_ (.B1(_1899_),
    .Y(_1900_),
    .A1(net148),
    .A2(net146));
 sg13g2_and2_1 _5217_ (.A(_1139_),
    .B(net147),
    .X(_1901_));
 sg13g2_buf_1 _5218_ (.A(_1901_),
    .X(_1902_));
 sg13g2_nand2_1 _5219_ (.Y(_1903_),
    .A(net100),
    .B(net146));
 sg13g2_nor3_1 _5220_ (.A(net148),
    .B(_1902_),
    .C(_1903_),
    .Y(_1904_));
 sg13g2_a221oi_1 _5221_ (.B2(_1902_),
    .C1(_1904_),
    .B1(_1900_),
    .A1(net148),
    .Y(_1905_),
    .A2(_1898_));
 sg13g2_nor2_1 _5222_ (.A(_1889_),
    .B(_1905_),
    .Y(_0331_));
 sg13g2_nand2_1 _5223_ (.Y(_1906_),
    .A(\mem[19][0] ),
    .B(_1141_));
 sg13g2_nand2_1 _5224_ (.Y(_1907_),
    .A(net147),
    .B(\mem[3][2] ));
 sg13g2_nand2_1 _5225_ (.Y(_1908_),
    .A(_1139_),
    .B(net146));
 sg13g2_xor2_1 _5226_ (.B(_1908_),
    .A(_1907_),
    .X(_1909_));
 sg13g2_xnor2_1 _5227_ (.Y(_1910_),
    .A(_1906_),
    .B(_1909_));
 sg13g2_buf_2 _5228_ (.A(_1910_),
    .X(_1911_));
 sg13g2_a21oi_1 _5229_ (.A1(net148),
    .A2(net99),
    .Y(_1912_),
    .B1(_1902_));
 sg13g2_nand3_1 _5230_ (.B(net99),
    .C(_1902_),
    .A(_0644_),
    .Y(_1913_));
 sg13g2_o21ai_1 _5231_ (.B1(_1913_),
    .Y(_1914_),
    .A1(_1903_),
    .A2(_1912_));
 sg13g2_buf_1 _5232_ (.A(_1914_),
    .X(_1915_));
 sg13g2_nand2_2 _5233_ (.Y(_1916_),
    .A(_1137_),
    .B(net145));
 sg13g2_nor3_2 _5234_ (.A(_1890_),
    .B(_1896_),
    .C(_1894_),
    .Y(_1917_));
 sg13g2_xor2_1 _5235_ (.B(_1917_),
    .A(_1916_),
    .X(_1918_));
 sg13g2_xnor2_1 _5236_ (.Y(_1919_),
    .A(_1915_),
    .B(_1918_));
 sg13g2_xnor2_1 _5237_ (.Y(_1920_),
    .A(_1911_),
    .B(_1919_));
 sg13g2_nor2_1 _5238_ (.A(_1889_),
    .B(_1920_),
    .Y(_0332_));
 sg13g2_and2_1 _5239_ (.A(_1907_),
    .B(_1908_),
    .X(_1921_));
 sg13g2_or2_1 _5240_ (.X(_1922_),
    .B(_1908_),
    .A(_1907_));
 sg13g2_o21ai_1 _5241_ (.B1(_1922_),
    .Y(_1923_),
    .A1(_1906_),
    .A2(_1921_));
 sg13g2_nand2_2 _5242_ (.Y(_1924_),
    .A(net99),
    .B(net146));
 sg13g2_nand2_1 _5243_ (.Y(_1925_),
    .A(net147),
    .B(_1141_));
 sg13g2_xor2_1 _5244_ (.B(_1925_),
    .A(_1924_),
    .X(_1926_));
 sg13g2_nand2_1 _5245_ (.Y(_1927_),
    .A(_1139_),
    .B(\mem[19][3] ));
 sg13g2_xor2_1 _5246_ (.B(_1927_),
    .A(_1926_),
    .X(_1928_));
 sg13g2_xnor2_1 _5247_ (.Y(_1929_),
    .A(_1923_),
    .B(_1928_));
 sg13g2_nand2_1 _5248_ (.Y(_1930_),
    .A(_1915_),
    .B(_1911_));
 sg13g2_nor2_1 _5249_ (.A(_1915_),
    .B(_1911_),
    .Y(_1931_));
 sg13g2_a21oi_1 _5250_ (.A1(_1916_),
    .A2(_1930_),
    .Y(_1932_),
    .B1(_1931_));
 sg13g2_inv_1 _5251_ (.Y(_1933_),
    .A(_1917_));
 sg13g2_nor3_1 _5252_ (.A(_1916_),
    .B(_1933_),
    .C(_1930_),
    .Y(_1934_));
 sg13g2_a21oi_1 _5253_ (.A1(_1916_),
    .A2(_1931_),
    .Y(_1935_),
    .B1(_1934_));
 sg13g2_o21ai_1 _5254_ (.B1(_1935_),
    .Y(_1936_),
    .A1(_1917_),
    .A2(_1932_));
 sg13g2_xor2_1 _5255_ (.B(_1936_),
    .A(_1929_),
    .X(_1937_));
 sg13g2_nor2_1 _5256_ (.A(_1889_),
    .B(_1937_),
    .Y(_0333_));
 sg13g2_and2_1 _5257_ (.A(_1911_),
    .B(_1917_),
    .X(_1938_));
 sg13g2_o21ai_1 _5258_ (.B1(_1915_),
    .Y(_1939_),
    .A1(_1911_),
    .A2(_1917_));
 sg13g2_nand2b_1 _5259_ (.Y(_1940_),
    .B(_1939_),
    .A_N(_1938_));
 sg13g2_o21ai_1 _5260_ (.B1(_1915_),
    .Y(_1941_),
    .A1(_1929_),
    .A2(_1938_));
 sg13g2_o21ai_1 _5261_ (.B1(_1929_),
    .Y(_1942_),
    .A1(_1911_),
    .A2(_1917_));
 sg13g2_a21oi_1 _5262_ (.A1(_1941_),
    .A2(_1942_),
    .Y(_1943_),
    .B1(_1916_));
 sg13g2_a21oi_1 _5263_ (.A1(_1929_),
    .A2(_1940_),
    .Y(_1944_),
    .B1(_1943_));
 sg13g2_nor2_1 _5264_ (.A(_1923_),
    .B(_1926_),
    .Y(_1945_));
 sg13g2_a22oi_1 _5265_ (.Y(_1946_),
    .B1(_1923_),
    .B2(_1926_),
    .A2(_0653_),
    .A1(_1139_));
 sg13g2_nor2_1 _5266_ (.A(_1945_),
    .B(_1946_),
    .Y(_1947_));
 sg13g2_o21ai_1 _5267_ (.B1(net99),
    .Y(_1948_),
    .A1(net147),
    .A2(net145));
 sg13g2_nand3_1 _5268_ (.B(_1141_),
    .C(_1948_),
    .A(net146),
    .Y(_1949_));
 sg13g2_nand3_1 _5269_ (.B(net146),
    .C(_1141_),
    .A(_0647_),
    .Y(_1950_));
 sg13g2_nand3_1 _5270_ (.B(net145),
    .C(_1950_),
    .A(net99),
    .Y(_1951_));
 sg13g2_and2_1 _5271_ (.A(_1949_),
    .B(_1951_),
    .X(_1952_));
 sg13g2_nor2b_1 _5272_ (.A(_1947_),
    .B_N(_1952_),
    .Y(_1953_));
 sg13g2_or3_1 _5273_ (.A(_1945_),
    .B(_1946_),
    .C(_1952_),
    .X(_1954_));
 sg13g2_nand2b_1 _5274_ (.Y(_1955_),
    .B(_1954_),
    .A_N(_1953_));
 sg13g2_xnor2_1 _5275_ (.Y(_1956_),
    .A(_1944_),
    .B(_1955_));
 sg13g2_nor2_1 _5276_ (.A(_1889_),
    .B(_1956_),
    .Y(_0334_));
 sg13g2_a21oi_2 _5277_ (.B1(_1953_),
    .Y(_1957_),
    .A2(_1954_),
    .A1(_1944_));
 sg13g2_inv_1 _5278_ (.Y(_1958_),
    .A(_1141_));
 sg13g2_nor3_1 _5279_ (.A(_0647_),
    .B(net145),
    .C(_1924_),
    .Y(_1959_));
 sg13g2_a21oi_1 _5280_ (.A1(net145),
    .A2(_1924_),
    .Y(_1960_),
    .B1(_1959_));
 sg13g2_nor2_1 _5281_ (.A(_1958_),
    .B(_1960_),
    .Y(_1961_));
 sg13g2_xnor2_1 _5282_ (.Y(_1962_),
    .A(_1957_),
    .B(_1961_));
 sg13g2_nor2_1 _5283_ (.A(_1889_),
    .B(_1962_),
    .Y(_0335_));
 sg13g2_a21oi_1 _5284_ (.A1(net147),
    .A2(_1957_),
    .Y(_1963_),
    .B1(net145));
 sg13g2_nor2_1 _5285_ (.A(_1924_),
    .B(_1963_),
    .Y(_1964_));
 sg13g2_a21oi_1 _5286_ (.A1(net145),
    .A2(_1957_),
    .Y(_1965_),
    .B1(_1964_));
 sg13g2_nor3_1 _5287_ (.A(_1958_),
    .B(_1889_),
    .C(_1965_),
    .Y(_0336_));
 sg13g2_nand2_1 _5288_ (.Y(_1966_),
    .A(net98),
    .B(_0665_));
 sg13g2_nor2_1 _5289_ (.A(net55),
    .B(_1966_),
    .Y(_0337_));
 sg13g2_nand2_1 _5290_ (.Y(_1967_),
    .A(net98),
    .B(net141));
 sg13g2_nand2_1 _5291_ (.Y(_1968_),
    .A(net142),
    .B(_1164_));
 sg13g2_xnor2_1 _5292_ (.Y(_1969_),
    .A(_1967_),
    .B(_1968_));
 sg13g2_nor2_1 _5293_ (.A(_1807_),
    .B(_1969_),
    .Y(_0338_));
 sg13g2_nand2_1 _5294_ (.Y(_1970_),
    .A(_1164_),
    .B(net141));
 sg13g2_nand2_1 _5295_ (.Y(_1971_),
    .A(net97),
    .B(_1970_));
 sg13g2_xor2_1 _5296_ (.B(net140),
    .A(net97),
    .X(_1972_));
 sg13g2_nand2_1 _5297_ (.Y(_1973_),
    .A(net98),
    .B(_1972_));
 sg13g2_o21ai_1 _5298_ (.B1(_1973_),
    .Y(_1974_),
    .A1(net98),
    .A2(_1971_));
 sg13g2_a21o_1 _5299_ (.A2(net97),
    .A1(net142),
    .B1(net98),
    .X(_1975_));
 sg13g2_o21ai_1 _5300_ (.B1(_1975_),
    .Y(_1976_),
    .A1(net142),
    .A2(net140));
 sg13g2_and2_1 _5301_ (.A(_1164_),
    .B(_0667_),
    .X(_1977_));
 sg13g2_buf_1 _5302_ (.A(_1977_),
    .X(_1978_));
 sg13g2_nand2_1 _5303_ (.Y(_1979_),
    .A(net98),
    .B(net140));
 sg13g2_nor3_1 _5304_ (.A(net142),
    .B(_1978_),
    .C(_1979_),
    .Y(_1980_));
 sg13g2_a221oi_1 _5305_ (.B2(_1978_),
    .C1(_1980_),
    .B1(_1976_),
    .A1(_0665_),
    .Y(_1981_),
    .A2(_1974_));
 sg13g2_nor2_1 _5306_ (.A(net55),
    .B(_1981_),
    .Y(_0339_));
 sg13g2_nand2_1 _5307_ (.Y(_1982_),
    .A(\mem[20][0] ),
    .B(_1166_));
 sg13g2_nand2_1 _5308_ (.Y(_1983_),
    .A(net141),
    .B(\mem[4][2] ));
 sg13g2_nand2_1 _5309_ (.Y(_1984_),
    .A(_1164_),
    .B(_0670_));
 sg13g2_xor2_1 _5310_ (.B(_1984_),
    .A(_1983_),
    .X(_1985_));
 sg13g2_xnor2_1 _5311_ (.Y(_1986_),
    .A(_1982_),
    .B(_1985_));
 sg13g2_buf_1 _5312_ (.A(_1986_),
    .X(_1987_));
 sg13g2_a21oi_1 _5313_ (.A1(net142),
    .A2(net97),
    .Y(_1988_),
    .B1(_1978_));
 sg13g2_nand3_1 _5314_ (.B(net97),
    .C(_1978_),
    .A(net142),
    .Y(_1989_));
 sg13g2_o21ai_1 _5315_ (.B1(_1989_),
    .Y(_1990_),
    .A1(_1979_),
    .A2(_1988_));
 sg13g2_buf_1 _5316_ (.A(_1990_),
    .X(_1991_));
 sg13g2_nand2_2 _5317_ (.Y(_1992_),
    .A(_1161_),
    .B(_0671_));
 sg13g2_nor3_2 _5318_ (.A(_1966_),
    .B(_1972_),
    .C(_1970_),
    .Y(_1993_));
 sg13g2_xor2_1 _5319_ (.B(_1993_),
    .A(_1992_),
    .X(_1994_));
 sg13g2_xnor2_1 _5320_ (.Y(_1995_),
    .A(_1991_),
    .B(_1994_));
 sg13g2_xnor2_1 _5321_ (.Y(_1996_),
    .A(_1987_),
    .B(_1995_));
 sg13g2_nor2_1 _5322_ (.A(net55),
    .B(_1996_),
    .Y(_0340_));
 sg13g2_and2_1 _5323_ (.A(_1983_),
    .B(_1984_),
    .X(_1997_));
 sg13g2_or2_1 _5324_ (.X(_1998_),
    .B(_1984_),
    .A(_1983_));
 sg13g2_o21ai_1 _5325_ (.B1(_1998_),
    .Y(_1999_),
    .A1(_1982_),
    .A2(_1997_));
 sg13g2_nand2_2 _5326_ (.Y(_2000_),
    .A(net97),
    .B(net140));
 sg13g2_nand2_1 _5327_ (.Y(_2001_),
    .A(net141),
    .B(_1166_));
 sg13g2_xor2_1 _5328_ (.B(_2001_),
    .A(_2000_),
    .X(_2002_));
 sg13g2_nand2_1 _5329_ (.Y(_2003_),
    .A(_1164_),
    .B(\mem[20][3] ));
 sg13g2_xor2_1 _5330_ (.B(_2003_),
    .A(_2002_),
    .X(_2004_));
 sg13g2_xnor2_1 _5331_ (.Y(_2005_),
    .A(_1999_),
    .B(_2004_));
 sg13g2_nand2_1 _5332_ (.Y(_2006_),
    .A(_1991_),
    .B(_1987_));
 sg13g2_nor2_1 _5333_ (.A(_1991_),
    .B(_1987_),
    .Y(_2007_));
 sg13g2_a21oi_1 _5334_ (.A1(_1992_),
    .A2(_2006_),
    .Y(_2008_),
    .B1(_2007_));
 sg13g2_inv_1 _5335_ (.Y(_2009_),
    .A(_1993_));
 sg13g2_nor3_1 _5336_ (.A(_1992_),
    .B(_2009_),
    .C(_2006_),
    .Y(_2010_));
 sg13g2_a21oi_1 _5337_ (.A1(_1992_),
    .A2(_2007_),
    .Y(_2011_),
    .B1(_2010_));
 sg13g2_o21ai_1 _5338_ (.B1(_2011_),
    .Y(_2012_),
    .A1(_1993_),
    .A2(_2008_));
 sg13g2_xor2_1 _5339_ (.B(_2012_),
    .A(_2005_),
    .X(_2013_));
 sg13g2_nor2_1 _5340_ (.A(net55),
    .B(_2013_),
    .Y(_0341_));
 sg13g2_and2_1 _5341_ (.A(_1987_),
    .B(_1993_),
    .X(_2014_));
 sg13g2_o21ai_1 _5342_ (.B1(_1991_),
    .Y(_2015_),
    .A1(_1987_),
    .A2(_1993_));
 sg13g2_nand2b_1 _5343_ (.Y(_2016_),
    .B(_2015_),
    .A_N(_2014_));
 sg13g2_o21ai_1 _5344_ (.B1(_1991_),
    .Y(_2017_),
    .A1(_2005_),
    .A2(_2014_));
 sg13g2_o21ai_1 _5345_ (.B1(_2005_),
    .Y(_2018_),
    .A1(_1987_),
    .A2(_1993_));
 sg13g2_a21oi_1 _5346_ (.A1(_2017_),
    .A2(_2018_),
    .Y(_2019_),
    .B1(_1992_));
 sg13g2_a21oi_1 _5347_ (.A1(_2005_),
    .A2(_2016_),
    .Y(_2020_),
    .B1(_2019_));
 sg13g2_nor2_1 _5348_ (.A(_1999_),
    .B(_2002_),
    .Y(_2021_));
 sg13g2_a22oi_1 _5349_ (.Y(_2022_),
    .B1(_1999_),
    .B2(_2002_),
    .A2(net139),
    .A1(_1164_));
 sg13g2_nor2_1 _5350_ (.A(_2021_),
    .B(_2022_),
    .Y(_2023_));
 sg13g2_o21ai_1 _5351_ (.B1(net97),
    .Y(_2024_),
    .A1(net141),
    .A2(net139));
 sg13g2_nand3_1 _5352_ (.B(_1166_),
    .C(_2024_),
    .A(net140),
    .Y(_2025_));
 sg13g2_nand3_1 _5353_ (.B(net140),
    .C(_1166_),
    .A(_0668_),
    .Y(_2026_));
 sg13g2_nand3_1 _5354_ (.B(net139),
    .C(_2026_),
    .A(_1165_),
    .Y(_2027_));
 sg13g2_and2_1 _5355_ (.A(_2025_),
    .B(_2027_),
    .X(_2028_));
 sg13g2_nor2b_1 _5356_ (.A(_2023_),
    .B_N(_2028_),
    .Y(_2029_));
 sg13g2_or3_1 _5357_ (.A(_2021_),
    .B(_2022_),
    .C(_2028_),
    .X(_2030_));
 sg13g2_nand2b_1 _5358_ (.Y(_2031_),
    .B(_2030_),
    .A_N(_2029_));
 sg13g2_xnor2_1 _5359_ (.Y(_2032_),
    .A(_2020_),
    .B(_2031_));
 sg13g2_nor2_1 _5360_ (.A(net55),
    .B(_2032_),
    .Y(_0342_));
 sg13g2_a21oi_2 _5361_ (.B1(_2029_),
    .Y(_2033_),
    .A2(_2030_),
    .A1(_2020_));
 sg13g2_inv_1 _5362_ (.Y(_2034_),
    .A(_1166_));
 sg13g2_nor3_1 _5363_ (.A(_0668_),
    .B(net139),
    .C(_2000_),
    .Y(_2035_));
 sg13g2_a21oi_1 _5364_ (.A1(net139),
    .A2(_2000_),
    .Y(_2036_),
    .B1(_2035_));
 sg13g2_nor2_1 _5365_ (.A(_2034_),
    .B(_2036_),
    .Y(_2037_));
 sg13g2_xnor2_1 _5366_ (.Y(_2038_),
    .A(_2033_),
    .B(_2037_));
 sg13g2_nor2_1 _5367_ (.A(net55),
    .B(_2038_),
    .Y(_0343_));
 sg13g2_a21oi_1 _5368_ (.A1(net141),
    .A2(_2033_),
    .Y(_2039_),
    .B1(net139));
 sg13g2_nor2_1 _5369_ (.A(_2000_),
    .B(_2039_),
    .Y(_2040_));
 sg13g2_a21oi_1 _5370_ (.A1(net139),
    .A2(_2033_),
    .Y(_2041_),
    .B1(_2040_));
 sg13g2_nor3_1 _5371_ (.A(_2034_),
    .B(net55),
    .C(_2041_),
    .Y(_0344_));
 sg13g2_xor2_1 _5372_ (.B(_1490_),
    .A(net173),
    .X(_2042_));
 sg13g2_o21ai_1 _5373_ (.B1(net57),
    .Y(_2043_),
    .A1(net81),
    .A2(_2042_));
 sg13g2_buf_2 _5374_ (.A(_2043_),
    .X(_2044_));
 sg13g2_nand2_1 _5375_ (.Y(_2045_),
    .A(net96),
    .B(net138));
 sg13g2_nor2_1 _5376_ (.A(_2044_),
    .B(_2045_),
    .Y(_0345_));
 sg13g2_nand2_1 _5377_ (.Y(_2046_),
    .A(net96),
    .B(net137));
 sg13g2_nand2_1 _5378_ (.Y(_2047_),
    .A(net138),
    .B(_1185_));
 sg13g2_xnor2_1 _5379_ (.Y(_2048_),
    .A(_2046_),
    .B(_2047_));
 sg13g2_nor2_1 _5380_ (.A(_2044_),
    .B(_2048_),
    .Y(_0346_));
 sg13g2_nand2_1 _5381_ (.Y(_2049_),
    .A(_1185_),
    .B(net137));
 sg13g2_nand2_1 _5382_ (.Y(_2050_),
    .A(net95),
    .B(_2049_));
 sg13g2_xor2_1 _5383_ (.B(net136),
    .A(net95),
    .X(_2051_));
 sg13g2_nand2_1 _5384_ (.Y(_2052_),
    .A(net96),
    .B(_2051_));
 sg13g2_o21ai_1 _5385_ (.B1(_2052_),
    .Y(_2053_),
    .A1(net96),
    .A2(_2050_));
 sg13g2_a21o_1 _5386_ (.A2(net95),
    .A1(net138),
    .B1(net96),
    .X(_2054_));
 sg13g2_o21ai_1 _5387_ (.B1(_2054_),
    .Y(_2055_),
    .A1(net138),
    .A2(_0677_));
 sg13g2_and2_1 _5388_ (.A(_1185_),
    .B(net137),
    .X(_2056_));
 sg13g2_buf_1 _5389_ (.A(_2056_),
    .X(_2057_));
 sg13g2_nand2_1 _5390_ (.Y(_2058_),
    .A(net96),
    .B(net136));
 sg13g2_nor3_1 _5391_ (.A(net138),
    .B(_2057_),
    .C(_2058_),
    .Y(_2059_));
 sg13g2_a221oi_1 _5392_ (.B2(_2057_),
    .C1(_2059_),
    .B1(_2055_),
    .A1(net138),
    .Y(_2060_),
    .A2(_2053_));
 sg13g2_nor2_1 _5393_ (.A(_2044_),
    .B(_2060_),
    .Y(_0347_));
 sg13g2_nand2_1 _5394_ (.Y(_2061_),
    .A(\mem[21][0] ),
    .B(_1187_));
 sg13g2_nand2_1 _5395_ (.Y(_2062_),
    .A(net137),
    .B(\mem[5][2] ));
 sg13g2_nand2_1 _5396_ (.Y(_2063_),
    .A(_1185_),
    .B(net136));
 sg13g2_xor2_1 _5397_ (.B(_2063_),
    .A(_2062_),
    .X(_2064_));
 sg13g2_xnor2_1 _5398_ (.Y(_2065_),
    .A(_2061_),
    .B(_2064_));
 sg13g2_buf_2 _5399_ (.A(_2065_),
    .X(_2066_));
 sg13g2_a21oi_1 _5400_ (.A1(net138),
    .A2(net95),
    .Y(_2067_),
    .B1(_2057_));
 sg13g2_nand3_1 _5401_ (.B(net95),
    .C(_2057_),
    .A(net138),
    .Y(_2068_));
 sg13g2_o21ai_1 _5402_ (.B1(_2068_),
    .Y(_2069_),
    .A1(_2058_),
    .A2(_2067_));
 sg13g2_buf_1 _5403_ (.A(_2069_),
    .X(_2070_));
 sg13g2_nand2_2 _5404_ (.Y(_2071_),
    .A(_1183_),
    .B(net135));
 sg13g2_nor3_2 _5405_ (.A(_2045_),
    .B(_2051_),
    .C(_2049_),
    .Y(_2072_));
 sg13g2_xor2_1 _5406_ (.B(_2072_),
    .A(_2071_),
    .X(_2073_));
 sg13g2_xnor2_1 _5407_ (.Y(_2074_),
    .A(_2070_),
    .B(_2073_));
 sg13g2_xnor2_1 _5408_ (.Y(_2075_),
    .A(_2066_),
    .B(_2074_));
 sg13g2_nor2_1 _5409_ (.A(_2044_),
    .B(_2075_),
    .Y(_0348_));
 sg13g2_and2_1 _5410_ (.A(_2062_),
    .B(_2063_),
    .X(_2076_));
 sg13g2_or2_1 _5411_ (.X(_2077_),
    .B(_2063_),
    .A(_2062_));
 sg13g2_o21ai_1 _5412_ (.B1(_2077_),
    .Y(_2078_),
    .A1(_2061_),
    .A2(_2076_));
 sg13g2_nand2_2 _5413_ (.Y(_2079_),
    .A(net95),
    .B(net136));
 sg13g2_nand2_1 _5414_ (.Y(_2080_),
    .A(net137),
    .B(_1187_));
 sg13g2_xor2_1 _5415_ (.B(_2080_),
    .A(_2079_),
    .X(_2081_));
 sg13g2_nand2_1 _5416_ (.Y(_2082_),
    .A(_1185_),
    .B(\mem[21][3] ));
 sg13g2_xor2_1 _5417_ (.B(_2082_),
    .A(_2081_),
    .X(_2083_));
 sg13g2_xnor2_1 _5418_ (.Y(_2084_),
    .A(_2078_),
    .B(_2083_));
 sg13g2_nand2_1 _5419_ (.Y(_2085_),
    .A(_2070_),
    .B(_2066_));
 sg13g2_nor2_1 _5420_ (.A(_2070_),
    .B(_2066_),
    .Y(_2086_));
 sg13g2_a21oi_1 _5421_ (.A1(_2071_),
    .A2(_2085_),
    .Y(_2087_),
    .B1(_2086_));
 sg13g2_inv_1 _5422_ (.Y(_2088_),
    .A(_2072_));
 sg13g2_nor3_1 _5423_ (.A(_2071_),
    .B(_2088_),
    .C(_2085_),
    .Y(_2089_));
 sg13g2_a21oi_1 _5424_ (.A1(_2071_),
    .A2(_2086_),
    .Y(_2090_),
    .B1(_2089_));
 sg13g2_o21ai_1 _5425_ (.B1(_2090_),
    .Y(_2091_),
    .A1(_2072_),
    .A2(_2087_));
 sg13g2_xor2_1 _5426_ (.B(_2091_),
    .A(_2084_),
    .X(_2092_));
 sg13g2_nor2_1 _5427_ (.A(_2044_),
    .B(_2092_),
    .Y(_0349_));
 sg13g2_and2_1 _5428_ (.A(_2066_),
    .B(_2072_),
    .X(_2093_));
 sg13g2_o21ai_1 _5429_ (.B1(_2070_),
    .Y(_2094_),
    .A1(_2066_),
    .A2(_2072_));
 sg13g2_nand2b_1 _5430_ (.Y(_2095_),
    .B(_2094_),
    .A_N(_2093_));
 sg13g2_o21ai_1 _5431_ (.B1(_2070_),
    .Y(_2096_),
    .A1(_2084_),
    .A2(_2093_));
 sg13g2_o21ai_1 _5432_ (.B1(_2084_),
    .Y(_2097_),
    .A1(_2066_),
    .A2(_2072_));
 sg13g2_a21oi_1 _5433_ (.A1(_2096_),
    .A2(_2097_),
    .Y(_2098_),
    .B1(_2071_));
 sg13g2_a21oi_1 _5434_ (.A1(_2084_),
    .A2(_2095_),
    .Y(_2099_),
    .B1(_2098_));
 sg13g2_nor2_1 _5435_ (.A(_2078_),
    .B(_2081_),
    .Y(_2100_));
 sg13g2_a22oi_1 _5436_ (.Y(_2101_),
    .B1(_2078_),
    .B2(_2081_),
    .A2(net135),
    .A1(_1185_));
 sg13g2_nor2_1 _5437_ (.A(_2100_),
    .B(_2101_),
    .Y(_2102_));
 sg13g2_o21ai_1 _5438_ (.B1(net95),
    .Y(_2103_),
    .A1(net137),
    .A2(net135));
 sg13g2_nand3_1 _5439_ (.B(_1187_),
    .C(_2103_),
    .A(net136),
    .Y(_2104_));
 sg13g2_nand3_1 _5440_ (.B(net136),
    .C(_1187_),
    .A(_0675_),
    .Y(_2105_));
 sg13g2_nand3_1 _5441_ (.B(net135),
    .C(_2105_),
    .A(net95),
    .Y(_2106_));
 sg13g2_and2_1 _5442_ (.A(_2104_),
    .B(_2106_),
    .X(_2107_));
 sg13g2_nor2b_1 _5443_ (.A(_2102_),
    .B_N(_2107_),
    .Y(_2108_));
 sg13g2_or3_1 _5444_ (.A(_2100_),
    .B(_2101_),
    .C(_2107_),
    .X(_2109_));
 sg13g2_nand2b_1 _5445_ (.Y(_2110_),
    .B(_2109_),
    .A_N(_2108_));
 sg13g2_xnor2_1 _5446_ (.Y(_2111_),
    .A(_2099_),
    .B(_2110_));
 sg13g2_nor2_1 _5447_ (.A(_2044_),
    .B(_2111_),
    .Y(_0350_));
 sg13g2_a21oi_1 _5448_ (.A1(_2099_),
    .A2(_2109_),
    .Y(_2112_),
    .B1(_2108_));
 sg13g2_inv_1 _5449_ (.Y(_2113_),
    .A(_1187_));
 sg13g2_nor3_1 _5450_ (.A(_0675_),
    .B(net135),
    .C(_2079_),
    .Y(_2114_));
 sg13g2_a21oi_1 _5451_ (.A1(net135),
    .A2(_2079_),
    .Y(_2115_),
    .B1(_2114_));
 sg13g2_nor2_1 _5452_ (.A(_2113_),
    .B(_2115_),
    .Y(_2116_));
 sg13g2_xnor2_1 _5453_ (.Y(_2117_),
    .A(_2112_),
    .B(_2116_));
 sg13g2_nor2_1 _5454_ (.A(_2044_),
    .B(_2117_),
    .Y(_0351_));
 sg13g2_a21oi_1 _5455_ (.A1(net137),
    .A2(_2112_),
    .Y(_2118_),
    .B1(_0678_));
 sg13g2_nor2_1 _5456_ (.A(_2079_),
    .B(_2118_),
    .Y(_2119_));
 sg13g2_a21oi_1 _5457_ (.A1(_0678_),
    .A2(_2112_),
    .Y(_2120_),
    .B1(_2119_));
 sg13g2_nor3_1 _5458_ (.A(_2113_),
    .B(_2044_),
    .C(_2120_),
    .Y(_0352_));
 sg13g2_nand3b_1 _5459_ (.B(_1313_),
    .C(net173),
    .Y(_2121_),
    .A_N(net81));
 sg13g2_nand2b_1 _5460_ (.Y(_2122_),
    .B(_2121_),
    .A_N(_1807_));
 sg13g2_buf_2 _5461_ (.A(_2122_),
    .X(_2123_));
 sg13g2_nand2_1 _5462_ (.Y(_2124_),
    .A(net94),
    .B(_0679_));
 sg13g2_nor2_1 _5463_ (.A(_2123_),
    .B(_2124_),
    .Y(_0353_));
 sg13g2_nand2_1 _5464_ (.Y(_2125_),
    .A(net94),
    .B(net133));
 sg13g2_nand2_1 _5465_ (.Y(_2126_),
    .A(net134),
    .B(_1194_));
 sg13g2_xnor2_1 _5466_ (.Y(_2127_),
    .A(_2125_),
    .B(_2126_));
 sg13g2_nor2_1 _5467_ (.A(_2123_),
    .B(_2127_),
    .Y(_0354_));
 sg13g2_nand2_1 _5468_ (.Y(_2128_),
    .A(_1194_),
    .B(net133));
 sg13g2_nand2_1 _5469_ (.Y(_2129_),
    .A(net93),
    .B(_2128_));
 sg13g2_xor2_1 _5470_ (.B(net132),
    .A(net93),
    .X(_2130_));
 sg13g2_nand2_1 _5471_ (.Y(_2131_),
    .A(net94),
    .B(_2130_));
 sg13g2_o21ai_1 _5472_ (.B1(_2131_),
    .Y(_2132_),
    .A1(net94),
    .A2(_2129_));
 sg13g2_a21o_1 _5473_ (.A2(net93),
    .A1(net134),
    .B1(net94),
    .X(_2133_));
 sg13g2_o21ai_1 _5474_ (.B1(_2133_),
    .Y(_2134_),
    .A1(net134),
    .A2(net132));
 sg13g2_and2_1 _5475_ (.A(_1194_),
    .B(net133),
    .X(_2135_));
 sg13g2_buf_1 _5476_ (.A(_2135_),
    .X(_2136_));
 sg13g2_nand2_1 _5477_ (.Y(_2137_),
    .A(net94),
    .B(_0684_));
 sg13g2_nor3_1 _5478_ (.A(net134),
    .B(_2136_),
    .C(_2137_),
    .Y(_2138_));
 sg13g2_a221oi_1 _5479_ (.B2(_2136_),
    .C1(_2138_),
    .B1(_2134_),
    .A1(net134),
    .Y(_2139_),
    .A2(_2132_));
 sg13g2_nor2_1 _5480_ (.A(_2123_),
    .B(_2139_),
    .Y(_0355_));
 sg13g2_nand2_1 _5481_ (.Y(_2140_),
    .A(\mem[22][0] ),
    .B(_1196_));
 sg13g2_nand2_1 _5482_ (.Y(_2141_),
    .A(net133),
    .B(\mem[6][2] ));
 sg13g2_nand2_1 _5483_ (.Y(_2142_),
    .A(_1194_),
    .B(net132));
 sg13g2_xor2_1 _5484_ (.B(_2142_),
    .A(_2141_),
    .X(_2143_));
 sg13g2_xnor2_1 _5485_ (.Y(_2144_),
    .A(_2140_),
    .B(_2143_));
 sg13g2_buf_1 _5486_ (.A(_2144_),
    .X(_2145_));
 sg13g2_a21oi_1 _5487_ (.A1(net134),
    .A2(net93),
    .Y(_2146_),
    .B1(_2136_));
 sg13g2_nand3_1 _5488_ (.B(_1195_),
    .C(_2136_),
    .A(net134),
    .Y(_2147_));
 sg13g2_o21ai_1 _5489_ (.B1(_2147_),
    .Y(_2148_),
    .A1(_2137_),
    .A2(_2146_));
 sg13g2_buf_1 _5490_ (.A(_2148_),
    .X(_2149_));
 sg13g2_nand2_2 _5491_ (.Y(_2150_),
    .A(net94),
    .B(_0685_));
 sg13g2_nor3_2 _5492_ (.A(_2124_),
    .B(_2130_),
    .C(_2128_),
    .Y(_2151_));
 sg13g2_xor2_1 _5493_ (.B(_2151_),
    .A(_2150_),
    .X(_2152_));
 sg13g2_xnor2_1 _5494_ (.Y(_2153_),
    .A(_2149_),
    .B(_2152_));
 sg13g2_xnor2_1 _5495_ (.Y(_2154_),
    .A(_2145_),
    .B(_2153_));
 sg13g2_nor2_1 _5496_ (.A(_2123_),
    .B(_2154_),
    .Y(_0356_));
 sg13g2_and2_1 _5497_ (.A(_2141_),
    .B(_2142_),
    .X(_2155_));
 sg13g2_or2_1 _5498_ (.X(_2156_),
    .B(_2142_),
    .A(_2141_));
 sg13g2_o21ai_1 _5499_ (.B1(_2156_),
    .Y(_2157_),
    .A1(_2140_),
    .A2(_2155_));
 sg13g2_nand2_2 _5500_ (.Y(_2158_),
    .A(net93),
    .B(net132));
 sg13g2_nand2_1 _5501_ (.Y(_2159_),
    .A(net133),
    .B(_1196_));
 sg13g2_xor2_1 _5502_ (.B(_2159_),
    .A(_2158_),
    .X(_2160_));
 sg13g2_nand2_1 _5503_ (.Y(_2161_),
    .A(_1194_),
    .B(\mem[22][3] ));
 sg13g2_xor2_1 _5504_ (.B(_2161_),
    .A(_2160_),
    .X(_2162_));
 sg13g2_xnor2_1 _5505_ (.Y(_2163_),
    .A(_2157_),
    .B(_2162_));
 sg13g2_nand2_1 _5506_ (.Y(_2164_),
    .A(_2149_),
    .B(_2145_));
 sg13g2_nor2_1 _5507_ (.A(_2149_),
    .B(_2145_),
    .Y(_2165_));
 sg13g2_a21oi_1 _5508_ (.A1(_2150_),
    .A2(_2164_),
    .Y(_2166_),
    .B1(_2165_));
 sg13g2_inv_1 _5509_ (.Y(_2167_),
    .A(_2151_));
 sg13g2_nor3_1 _5510_ (.A(_2150_),
    .B(_2167_),
    .C(_2164_),
    .Y(_2168_));
 sg13g2_a21oi_1 _5511_ (.A1(_2150_),
    .A2(_2165_),
    .Y(_2169_),
    .B1(_2168_));
 sg13g2_o21ai_1 _5512_ (.B1(_2169_),
    .Y(_2170_),
    .A1(_2151_),
    .A2(_2166_));
 sg13g2_xor2_1 _5513_ (.B(_2170_),
    .A(_2163_),
    .X(_2171_));
 sg13g2_nor2_1 _5514_ (.A(_2123_),
    .B(_2171_),
    .Y(_0357_));
 sg13g2_and2_1 _5515_ (.A(_2145_),
    .B(_2151_),
    .X(_2172_));
 sg13g2_o21ai_1 _5516_ (.B1(_2149_),
    .Y(_2173_),
    .A1(_2145_),
    .A2(_2151_));
 sg13g2_nand2b_1 _5517_ (.Y(_2174_),
    .B(_2173_),
    .A_N(_2172_));
 sg13g2_o21ai_1 _5518_ (.B1(_2149_),
    .Y(_2175_),
    .A1(_2163_),
    .A2(_2172_));
 sg13g2_o21ai_1 _5519_ (.B1(_2163_),
    .Y(_2176_),
    .A1(_2145_),
    .A2(_2151_));
 sg13g2_a21oi_1 _5520_ (.A1(_2175_),
    .A2(_2176_),
    .Y(_2177_),
    .B1(_2150_));
 sg13g2_a21oi_1 _5521_ (.A1(_2163_),
    .A2(_2174_),
    .Y(_2178_),
    .B1(_2177_));
 sg13g2_nor2_1 _5522_ (.A(_2157_),
    .B(_2160_),
    .Y(_2179_));
 sg13g2_a22oi_1 _5523_ (.Y(_2180_),
    .B1(_2157_),
    .B2(_2160_),
    .A2(net131),
    .A1(_1194_));
 sg13g2_nor2_1 _5524_ (.A(_2179_),
    .B(_2180_),
    .Y(_2181_));
 sg13g2_o21ai_1 _5525_ (.B1(net93),
    .Y(_2182_),
    .A1(net133),
    .A2(net131));
 sg13g2_nand3_1 _5526_ (.B(_1196_),
    .C(_2182_),
    .A(net132),
    .Y(_2183_));
 sg13g2_nand3_1 _5527_ (.B(net132),
    .C(_1196_),
    .A(_0682_),
    .Y(_2184_));
 sg13g2_nand3_1 _5528_ (.B(net131),
    .C(_2184_),
    .A(net93),
    .Y(_2185_));
 sg13g2_and2_1 _5529_ (.A(_2183_),
    .B(_2185_),
    .X(_2186_));
 sg13g2_nor2b_1 _5530_ (.A(_2181_),
    .B_N(_2186_),
    .Y(_2187_));
 sg13g2_or3_1 _5531_ (.A(_2179_),
    .B(_2180_),
    .C(_2186_),
    .X(_2188_));
 sg13g2_nand2b_1 _5532_ (.Y(_2189_),
    .B(_2188_),
    .A_N(_2187_));
 sg13g2_xnor2_1 _5533_ (.Y(_2190_),
    .A(_2178_),
    .B(_2189_));
 sg13g2_nor2_1 _5534_ (.A(_2123_),
    .B(_2190_),
    .Y(_0358_));
 sg13g2_a21oi_2 _5535_ (.B1(_2187_),
    .Y(_2191_),
    .A2(_2188_),
    .A1(_2178_));
 sg13g2_inv_1 _5536_ (.Y(_2192_),
    .A(_1196_));
 sg13g2_nor3_1 _5537_ (.A(_0682_),
    .B(net131),
    .C(_2158_),
    .Y(_2193_));
 sg13g2_a21oi_1 _5538_ (.A1(net131),
    .A2(_2158_),
    .Y(_2194_),
    .B1(_2193_));
 sg13g2_nor2_1 _5539_ (.A(_2192_),
    .B(_2194_),
    .Y(_2195_));
 sg13g2_xnor2_1 _5540_ (.Y(_2196_),
    .A(_2191_),
    .B(_2195_));
 sg13g2_nor2_1 _5541_ (.A(_2123_),
    .B(_2196_),
    .Y(_0359_));
 sg13g2_a21oi_1 _5542_ (.A1(net133),
    .A2(_2191_),
    .Y(_2197_),
    .B1(net131));
 sg13g2_nor2_1 _5543_ (.A(_2158_),
    .B(_2197_),
    .Y(_2198_));
 sg13g2_a21oi_1 _5544_ (.A1(net131),
    .A2(_2191_),
    .Y(_2199_),
    .B1(_2198_));
 sg13g2_nor3_1 _5545_ (.A(_2192_),
    .B(_2123_),
    .C(_2199_),
    .Y(_0360_));
 sg13g2_nand3_1 _5546_ (.B(net174),
    .C(net173),
    .A(_2634_),
    .Y(_2200_));
 sg13g2_nand2b_1 _5547_ (.Y(_2201_),
    .B(_2200_),
    .A_N(_1408_));
 sg13g2_o21ai_1 _5548_ (.B1(net57),
    .Y(_2202_),
    .A1(net81),
    .A2(_2201_));
 sg13g2_buf_2 _5549_ (.A(_2202_),
    .X(_2203_));
 sg13g2_nand2_1 _5550_ (.Y(_2204_),
    .A(net92),
    .B(net130));
 sg13g2_nor2_1 _5551_ (.A(_2203_),
    .B(_2204_),
    .Y(_0361_));
 sg13g2_nand2_1 _5552_ (.Y(_2205_),
    .A(net130),
    .B(_1199_));
 sg13g2_nand2_1 _5553_ (.Y(_2206_),
    .A(net92),
    .B(_0688_));
 sg13g2_xnor2_1 _5554_ (.Y(_2207_),
    .A(_2205_),
    .B(_2206_));
 sg13g2_nor2_1 _5555_ (.A(_2203_),
    .B(_2207_),
    .Y(_0362_));
 sg13g2_nand2_2 _5556_ (.Y(_2208_),
    .A(net130),
    .B(net91));
 sg13g2_and2_1 _5557_ (.A(_0688_),
    .B(_1199_),
    .X(_2209_));
 sg13g2_buf_1 _5558_ (.A(_2209_),
    .X(_2210_));
 sg13g2_nand2b_1 _5559_ (.Y(_2211_),
    .B(_2210_),
    .A_N(net130));
 sg13g2_nand3_1 _5560_ (.B(_2211_),
    .C(_2208_),
    .A(net129),
    .Y(_2212_));
 sg13g2_o21ai_1 _5561_ (.B1(_2212_),
    .Y(_2213_),
    .A1(net129),
    .A2(_2208_));
 sg13g2_nand2b_1 _5562_ (.Y(_2214_),
    .B(_2208_),
    .A_N(net92));
 sg13g2_o21ai_1 _5563_ (.B1(_2214_),
    .Y(_2215_),
    .A1(net129),
    .A2(net130));
 sg13g2_nor3_1 _5564_ (.A(net92),
    .B(_2210_),
    .C(_2208_),
    .Y(_2216_));
 sg13g2_a221oi_1 _5565_ (.B2(_2210_),
    .C1(_2216_),
    .B1(_2215_),
    .A1(net92),
    .Y(_2217_),
    .A2(_2213_));
 sg13g2_nor2_1 _5566_ (.A(_2203_),
    .B(_2217_),
    .Y(_0363_));
 sg13g2_nand2_1 _5567_ (.Y(_2218_),
    .A(\mem[23][2] ),
    .B(_1199_));
 sg13g2_nand2_1 _5568_ (.Y(_2219_),
    .A(_0688_),
    .B(net91));
 sg13g2_nand2_1 _5569_ (.Y(_2220_),
    .A(net130),
    .B(_1201_));
 sg13g2_xor2_1 _5570_ (.B(_2220_),
    .A(_2219_),
    .X(_2221_));
 sg13g2_xnor2_1 _5571_ (.Y(_2222_),
    .A(_2218_),
    .B(_2221_));
 sg13g2_nand2_1 _5572_ (.Y(_2223_),
    .A(_0688_),
    .B(_1199_));
 sg13g2_inv_1 _5573_ (.Y(_2224_),
    .A(_2208_));
 sg13g2_a22oi_1 _5574_ (.Y(_2225_),
    .B1(_2210_),
    .B2(_2224_),
    .A2(net92),
    .A1(net129));
 sg13g2_a21oi_2 _5575_ (.B1(_2225_),
    .Y(_2226_),
    .A2(_2208_),
    .A1(_2223_));
 sg13g2_nand2_2 _5576_ (.Y(_2227_),
    .A(_1197_),
    .B(net128));
 sg13g2_xnor2_1 _5577_ (.Y(_2228_),
    .A(net129),
    .B(net91));
 sg13g2_nand4_1 _5578_ (.B(net130),
    .C(_2210_),
    .A(_1197_),
    .Y(_2229_),
    .D(_2228_));
 sg13g2_buf_1 _5579_ (.A(_2229_),
    .X(_2230_));
 sg13g2_xnor2_1 _5580_ (.Y(_2231_),
    .A(_2227_),
    .B(_2230_));
 sg13g2_xnor2_1 _5581_ (.Y(_2232_),
    .A(_2226_),
    .B(_2231_));
 sg13g2_xnor2_1 _5582_ (.Y(_2233_),
    .A(_2222_),
    .B(_2232_));
 sg13g2_nor2_1 _5583_ (.A(_2203_),
    .B(_2233_),
    .Y(_0364_));
 sg13g2_and2_1 _5584_ (.A(_2219_),
    .B(_2220_),
    .X(_2234_));
 sg13g2_or2_1 _5585_ (.X(_2235_),
    .B(_2220_),
    .A(_2219_));
 sg13g2_o21ai_1 _5586_ (.B1(_2235_),
    .Y(_2236_),
    .A1(_2218_),
    .A2(_2234_));
 sg13g2_nand2_1 _5587_ (.Y(_2237_),
    .A(\mem[23][2] ),
    .B(net91));
 sg13g2_nand2_1 _5588_ (.Y(_2238_),
    .A(_1201_),
    .B(_0688_));
 sg13g2_xor2_1 _5589_ (.B(_2238_),
    .A(_2237_),
    .X(_2239_));
 sg13g2_nand2_1 _5590_ (.Y(_2240_),
    .A(_1199_),
    .B(net128));
 sg13g2_xor2_1 _5591_ (.B(_2240_),
    .A(_2239_),
    .X(_2241_));
 sg13g2_xnor2_1 _5592_ (.Y(_2242_),
    .A(_2236_),
    .B(_2241_));
 sg13g2_nor2_1 _5593_ (.A(_2226_),
    .B(_2222_),
    .Y(_2243_));
 sg13g2_nand2_1 _5594_ (.Y(_2244_),
    .A(_2226_),
    .B(_2222_));
 sg13g2_a21o_1 _5595_ (.A2(_2244_),
    .A1(_2227_),
    .B1(_2243_),
    .X(_2245_));
 sg13g2_nor3_1 _5596_ (.A(_2227_),
    .B(_2230_),
    .C(_2244_),
    .Y(_2246_));
 sg13g2_a221oi_1 _5597_ (.B2(_2230_),
    .C1(_2246_),
    .B1(_2245_),
    .A1(_2227_),
    .Y(_2247_),
    .A2(_2243_));
 sg13g2_xnor2_1 _5598_ (.Y(_2248_),
    .A(_2242_),
    .B(_2247_));
 sg13g2_nor2_1 _5599_ (.A(_2203_),
    .B(_2248_),
    .Y(_0365_));
 sg13g2_nand2b_1 _5600_ (.Y(_2249_),
    .B(_2230_),
    .A_N(_2222_));
 sg13g2_nor2b_1 _5601_ (.A(_2230_),
    .B_N(_2222_),
    .Y(_2250_));
 sg13g2_a21o_1 _5602_ (.A2(_2249_),
    .A1(_2226_),
    .B1(_2250_),
    .X(_2251_));
 sg13g2_o21ai_1 _5603_ (.B1(_2226_),
    .Y(_2252_),
    .A1(_2242_),
    .A2(_2250_));
 sg13g2_nand2_1 _5604_ (.Y(_2253_),
    .A(_2242_),
    .B(_2249_));
 sg13g2_a21oi_1 _5605_ (.A1(_2252_),
    .A2(_2253_),
    .Y(_2254_),
    .B1(_2227_));
 sg13g2_a21oi_1 _5606_ (.A1(_2242_),
    .A2(_2251_),
    .Y(_2255_),
    .B1(_2254_));
 sg13g2_nor2_1 _5607_ (.A(_2236_),
    .B(_2239_),
    .Y(_2256_));
 sg13g2_nand2_1 _5608_ (.Y(_2257_),
    .A(_2236_),
    .B(_2239_));
 sg13g2_o21ai_1 _5609_ (.B1(_2257_),
    .Y(_2258_),
    .A1(_2240_),
    .A2(_2256_));
 sg13g2_nand4_1 _5610_ (.B(_1201_),
    .C(_0689_),
    .A(net129),
    .Y(_2259_),
    .D(net128));
 sg13g2_nand2b_1 _5611_ (.Y(_2260_),
    .B(_0688_),
    .A_N(net128));
 sg13g2_nand2_1 _5612_ (.Y(_2261_),
    .A(_2259_),
    .B(_2260_));
 sg13g2_a22oi_1 _5613_ (.Y(_2262_),
    .B1(net91),
    .B2(net128),
    .A2(_1201_),
    .A1(net129));
 sg13g2_a21oi_1 _5614_ (.A1(net91),
    .A2(_2261_),
    .Y(_2263_),
    .B1(_2262_));
 sg13g2_nor2_1 _5615_ (.A(_2258_),
    .B(_2263_),
    .Y(_2264_));
 sg13g2_nand2_1 _5616_ (.Y(_2265_),
    .A(_2258_),
    .B(_2263_));
 sg13g2_nand2b_1 _5617_ (.Y(_2266_),
    .B(_2265_),
    .A_N(_2264_));
 sg13g2_xnor2_1 _5618_ (.Y(_2267_),
    .A(_2255_),
    .B(_2266_));
 sg13g2_nor2_1 _5619_ (.A(_2203_),
    .B(_2267_),
    .Y(_0366_));
 sg13g2_nand2_1 _5620_ (.Y(_2268_),
    .A(net128),
    .B(_2237_));
 sg13g2_o21ai_1 _5621_ (.B1(_2268_),
    .Y(_2269_),
    .A1(_2237_),
    .A2(_2260_));
 sg13g2_nand2_1 _5622_ (.Y(_2270_),
    .A(_1201_),
    .B(_2269_));
 sg13g2_a21oi_1 _5623_ (.A1(_2255_),
    .A2(_2265_),
    .Y(_2271_),
    .B1(_2264_));
 sg13g2_xor2_1 _5624_ (.B(_2271_),
    .A(_2270_),
    .X(_2272_));
 sg13g2_nor2_1 _5625_ (.A(_2203_),
    .B(_2272_),
    .Y(_0367_));
 sg13g2_nand2b_1 _5626_ (.Y(_2273_),
    .B(_2271_),
    .A_N(_2270_));
 sg13g2_nand4_1 _5627_ (.B(_1201_),
    .C(_1200_),
    .A(_0691_),
    .Y(_2274_),
    .D(net128));
 sg13g2_a21oi_1 _5628_ (.A1(_2273_),
    .A2(_2274_),
    .Y(_0368_),
    .B1(_2203_));
 sg13g2_o21ai_1 _5629_ (.B1(_1308_),
    .Y(_2275_),
    .A1(_0557_),
    .A2(_1408_));
 sg13g2_buf_1 _5630_ (.A(_2275_),
    .X(_2276_));
 sg13g2_nand2_1 _5631_ (.Y(_2277_),
    .A(net127),
    .B(net90));
 sg13g2_nor2_1 _5632_ (.A(net54),
    .B(_2277_),
    .Y(_0369_));
 sg13g2_nand2_1 _5633_ (.Y(_2278_),
    .A(_0698_),
    .B(net90));
 sg13g2_nand2_1 _5634_ (.Y(_2279_),
    .A(net127),
    .B(_1204_));
 sg13g2_xnor2_1 _5635_ (.Y(_2280_),
    .A(_2278_),
    .B(_2279_));
 sg13g2_nor2_1 _5636_ (.A(_2276_),
    .B(_2280_),
    .Y(_0370_));
 sg13g2_nand2_1 _5637_ (.Y(_2281_),
    .A(_1204_),
    .B(_0698_));
 sg13g2_buf_2 _5638_ (.A(_2281_),
    .X(_2282_));
 sg13g2_nand2_1 _5639_ (.Y(_2283_),
    .A(net89),
    .B(_2282_));
 sg13g2_xor2_1 _5640_ (.B(_0701_),
    .A(net89),
    .X(_2284_));
 sg13g2_nand2_1 _5641_ (.Y(_2285_),
    .A(net90),
    .B(_2284_));
 sg13g2_o21ai_1 _5642_ (.B1(_2285_),
    .Y(_2286_),
    .A1(net90),
    .A2(_2283_));
 sg13g2_nand2_2 _5643_ (.Y(_2287_),
    .A(net90),
    .B(_0701_));
 sg13g2_nor2_1 _5644_ (.A(net127),
    .B(_2287_),
    .Y(_2288_));
 sg13g2_nand2b_1 _5645_ (.Y(_2289_),
    .B(_2287_),
    .A_N(net127));
 sg13g2_or2_1 _5646_ (.X(_2290_),
    .B(net89),
    .A(net90));
 sg13g2_a21oi_1 _5647_ (.A1(_2289_),
    .A2(_2290_),
    .Y(_2291_),
    .B1(_2282_));
 sg13g2_a221oi_1 _5648_ (.B2(_2282_),
    .C1(_2291_),
    .B1(_2288_),
    .A1(net127),
    .Y(_2292_),
    .A2(_2286_));
 sg13g2_nor2_1 _5649_ (.A(net54),
    .B(_2292_),
    .Y(_0371_));
 sg13g2_nand2_1 _5650_ (.Y(_2293_),
    .A(net127),
    .B(_1206_));
 sg13g2_nand2_1 _5651_ (.Y(_2294_),
    .A(_0698_),
    .B(net89));
 sg13g2_nand2_1 _5652_ (.Y(_2295_),
    .A(_1204_),
    .B(_0701_));
 sg13g2_xor2_1 _5653_ (.B(_2295_),
    .A(_2294_),
    .X(_2296_));
 sg13g2_xnor2_1 _5654_ (.Y(_2297_),
    .A(_2293_),
    .B(_2296_));
 sg13g2_buf_2 _5655_ (.A(_2297_),
    .X(_2298_));
 sg13g2_nor2_1 _5656_ (.A(_2282_),
    .B(_2287_),
    .Y(_2299_));
 sg13g2_a21oi_1 _5657_ (.A1(net127),
    .A2(_1205_),
    .Y(_2300_),
    .B1(_2299_));
 sg13g2_a21oi_2 _5658_ (.B1(_2300_),
    .Y(_2301_),
    .A2(_2287_),
    .A1(_2282_));
 sg13g2_nand2_2 _5659_ (.Y(_2302_),
    .A(_1202_),
    .B(net126));
 sg13g2_nor3_2 _5660_ (.A(_2277_),
    .B(_2284_),
    .C(_2282_),
    .Y(_2303_));
 sg13g2_xor2_1 _5661_ (.B(_2303_),
    .A(_2302_),
    .X(_2304_));
 sg13g2_xnor2_1 _5662_ (.Y(_2305_),
    .A(_2301_),
    .B(_2304_));
 sg13g2_xnor2_1 _5663_ (.Y(_2306_),
    .A(_2298_),
    .B(_2305_));
 sg13g2_nor2_1 _5664_ (.A(net54),
    .B(_2306_),
    .Y(_0372_));
 sg13g2_and2_1 _5665_ (.A(_2294_),
    .B(_2295_),
    .X(_2307_));
 sg13g2_or2_1 _5666_ (.X(_2308_),
    .B(_2295_),
    .A(_2294_));
 sg13g2_o21ai_1 _5667_ (.B1(_2308_),
    .Y(_2309_),
    .A1(_2293_),
    .A2(_2307_));
 sg13g2_nand2_2 _5668_ (.Y(_2310_),
    .A(net89),
    .B(_0701_));
 sg13g2_nand2_1 _5669_ (.Y(_2311_),
    .A(_0698_),
    .B(_1206_));
 sg13g2_xor2_1 _5670_ (.B(_2311_),
    .A(_2310_),
    .X(_2312_));
 sg13g2_nand2_1 _5671_ (.Y(_2313_),
    .A(_1204_),
    .B(\mem[24][3] ));
 sg13g2_xor2_1 _5672_ (.B(_2313_),
    .A(_2312_),
    .X(_2314_));
 sg13g2_xnor2_1 _5673_ (.Y(_2315_),
    .A(_2309_),
    .B(_2314_));
 sg13g2_nand2_1 _5674_ (.Y(_2316_),
    .A(_2301_),
    .B(_2298_));
 sg13g2_nor2_1 _5675_ (.A(_2301_),
    .B(_2298_),
    .Y(_2317_));
 sg13g2_a21oi_1 _5676_ (.A1(_2302_),
    .A2(_2316_),
    .Y(_2318_),
    .B1(_2317_));
 sg13g2_inv_1 _5677_ (.Y(_2319_),
    .A(_2303_));
 sg13g2_nor3_1 _5678_ (.A(_2302_),
    .B(_2319_),
    .C(_2316_),
    .Y(_2320_));
 sg13g2_a21oi_1 _5679_ (.A1(_2302_),
    .A2(_2317_),
    .Y(_2321_),
    .B1(_2320_));
 sg13g2_o21ai_1 _5680_ (.B1(_2321_),
    .Y(_2322_),
    .A1(_2303_),
    .A2(_2318_));
 sg13g2_xor2_1 _5681_ (.B(_2322_),
    .A(_2315_),
    .X(_2323_));
 sg13g2_nor2_1 _5682_ (.A(net54),
    .B(_2323_),
    .Y(_0373_));
 sg13g2_and2_1 _5683_ (.A(_2298_),
    .B(_2303_),
    .X(_2324_));
 sg13g2_o21ai_1 _5684_ (.B1(_2301_),
    .Y(_2325_),
    .A1(_2298_),
    .A2(_2303_));
 sg13g2_nand2b_1 _5685_ (.Y(_2326_),
    .B(_2325_),
    .A_N(_2324_));
 sg13g2_o21ai_1 _5686_ (.B1(_2301_),
    .Y(_2327_),
    .A1(_2315_),
    .A2(_2324_));
 sg13g2_o21ai_1 _5687_ (.B1(_2315_),
    .Y(_2328_),
    .A1(_2298_),
    .A2(_2303_));
 sg13g2_a21oi_1 _5688_ (.A1(_2327_),
    .A2(_2328_),
    .Y(_2329_),
    .B1(_2302_));
 sg13g2_a21oi_1 _5689_ (.A1(_2315_),
    .A2(_2326_),
    .Y(_2330_),
    .B1(_2329_));
 sg13g2_nor2_1 _5690_ (.A(_2309_),
    .B(_2312_),
    .Y(_2331_));
 sg13g2_a22oi_1 _5691_ (.Y(_2332_),
    .B1(_2309_),
    .B2(_2312_),
    .A2(net126),
    .A1(_1204_));
 sg13g2_nor2_1 _5692_ (.A(_2331_),
    .B(_2332_),
    .Y(_2333_));
 sg13g2_o21ai_1 _5693_ (.B1(net89),
    .Y(_2334_),
    .A1(_0698_),
    .A2(net126));
 sg13g2_nand3_1 _5694_ (.B(_1206_),
    .C(_2334_),
    .A(_0701_),
    .Y(_2335_));
 sg13g2_nand3_1 _5695_ (.B(_0701_),
    .C(_1206_),
    .A(_0699_),
    .Y(_2336_));
 sg13g2_nand3_1 _5696_ (.B(net126),
    .C(_2336_),
    .A(_1205_),
    .Y(_2337_));
 sg13g2_and2_1 _5697_ (.A(_2335_),
    .B(_2337_),
    .X(_2338_));
 sg13g2_nor2b_1 _5698_ (.A(_2333_),
    .B_N(_2338_),
    .Y(_2339_));
 sg13g2_or3_1 _5699_ (.A(_2331_),
    .B(_2332_),
    .C(_2338_),
    .X(_2340_));
 sg13g2_nand2b_1 _5700_ (.Y(_2341_),
    .B(_2340_),
    .A_N(_2339_));
 sg13g2_xnor2_1 _5701_ (.Y(_2342_),
    .A(_2330_),
    .B(_2341_));
 sg13g2_nor2_1 _5702_ (.A(net54),
    .B(_2342_),
    .Y(_0374_));
 sg13g2_a21oi_2 _5703_ (.B1(_2339_),
    .Y(_2343_),
    .A2(_2340_),
    .A1(_2330_));
 sg13g2_inv_1 _5704_ (.Y(_2344_),
    .A(_1206_));
 sg13g2_nor3_1 _5705_ (.A(_0699_),
    .B(net126),
    .C(_2310_),
    .Y(_2345_));
 sg13g2_a21oi_1 _5706_ (.A1(net126),
    .A2(_2310_),
    .Y(_2346_),
    .B1(_2345_));
 sg13g2_nor2_1 _5707_ (.A(_2344_),
    .B(_2346_),
    .Y(_2347_));
 sg13g2_xnor2_1 _5708_ (.Y(_2348_),
    .A(_2343_),
    .B(_2347_));
 sg13g2_nor2_1 _5709_ (.A(net54),
    .B(_2348_),
    .Y(_0375_));
 sg13g2_a21oi_1 _5710_ (.A1(_0698_),
    .A2(_2343_),
    .Y(_2349_),
    .B1(net126));
 sg13g2_nor2_1 _5711_ (.A(_2310_),
    .B(_2349_),
    .Y(_2350_));
 sg13g2_a21oi_1 _5712_ (.A1(_0702_),
    .A2(_2343_),
    .Y(_2351_),
    .B1(_2350_));
 sg13g2_nor3_1 _5713_ (.A(_2344_),
    .B(net54),
    .C(_2351_),
    .Y(_0376_));
 sg13g2_nor2b_1 _5714_ (.A(_1408_),
    .B_N(net81),
    .Y(_2352_));
 sg13g2_o21ai_1 _5715_ (.B1(net57),
    .Y(_2353_),
    .A1(_1409_),
    .A2(_2352_));
 sg13g2_buf_2 _5716_ (.A(_2353_),
    .X(_2354_));
 sg13g2_nand2_1 _5717_ (.Y(_2355_),
    .A(net125),
    .B(net88));
 sg13g2_nor2_1 _5718_ (.A(_2354_),
    .B(_2355_),
    .Y(_0377_));
 sg13g2_nand2_1 _5719_ (.Y(_2356_),
    .A(_0705_),
    .B(net88));
 sg13g2_nand2_1 _5720_ (.Y(_2357_),
    .A(net125),
    .B(_1209_));
 sg13g2_xnor2_1 _5721_ (.Y(_2358_),
    .A(_2356_),
    .B(_2357_));
 sg13g2_nor2_1 _5722_ (.A(_2354_),
    .B(_2358_),
    .Y(_0378_));
 sg13g2_nand2_1 _5723_ (.Y(_2359_),
    .A(_1209_),
    .B(_0705_));
 sg13g2_buf_2 _5724_ (.A(_2359_),
    .X(_2360_));
 sg13g2_nand2_1 _5725_ (.Y(_2361_),
    .A(net87),
    .B(_2360_));
 sg13g2_xor2_1 _5726_ (.B(_0708_),
    .A(net87),
    .X(_2362_));
 sg13g2_nand2_1 _5727_ (.Y(_2363_),
    .A(net88),
    .B(_2362_));
 sg13g2_o21ai_1 _5728_ (.B1(_2363_),
    .Y(_2364_),
    .A1(net88),
    .A2(_2361_));
 sg13g2_nand2_2 _5729_ (.Y(_2365_),
    .A(net88),
    .B(_0708_));
 sg13g2_nor2_1 _5730_ (.A(net125),
    .B(_2365_),
    .Y(_2366_));
 sg13g2_nand2b_1 _5731_ (.Y(_2367_),
    .B(_2365_),
    .A_N(net125));
 sg13g2_or2_1 _5732_ (.X(_2368_),
    .B(_1210_),
    .A(net88));
 sg13g2_a21oi_1 _5733_ (.A1(_2367_),
    .A2(_2368_),
    .Y(_2369_),
    .B1(_2360_));
 sg13g2_a221oi_1 _5734_ (.B2(_2360_),
    .C1(_2369_),
    .B1(_2366_),
    .A1(net125),
    .Y(_2370_),
    .A2(_2364_));
 sg13g2_nor2_1 _5735_ (.A(_2354_),
    .B(_2370_),
    .Y(_0379_));
 sg13g2_nand2_1 _5736_ (.Y(_2371_),
    .A(net125),
    .B(_1211_));
 sg13g2_nand2_1 _5737_ (.Y(_2372_),
    .A(_0705_),
    .B(net87));
 sg13g2_nand2_1 _5738_ (.Y(_2373_),
    .A(_1209_),
    .B(_0708_));
 sg13g2_xor2_1 _5739_ (.B(_2373_),
    .A(_2372_),
    .X(_2374_));
 sg13g2_xnor2_1 _5740_ (.Y(_2375_),
    .A(_2371_),
    .B(_2374_));
 sg13g2_buf_1 _5741_ (.A(_2375_),
    .X(_2376_));
 sg13g2_nor2_1 _5742_ (.A(_2360_),
    .B(_2365_),
    .Y(_2377_));
 sg13g2_a21oi_1 _5743_ (.A1(net125),
    .A2(_1210_),
    .Y(_2378_),
    .B1(_2377_));
 sg13g2_a21oi_2 _5744_ (.B1(_2378_),
    .Y(_2379_),
    .A2(_2365_),
    .A1(_2360_));
 sg13g2_nand2_2 _5745_ (.Y(_2380_),
    .A(_1207_),
    .B(_0709_));
 sg13g2_nor3_2 _5746_ (.A(_2355_),
    .B(_2362_),
    .C(_2360_),
    .Y(_2381_));
 sg13g2_xor2_1 _5747_ (.B(_2381_),
    .A(_2380_),
    .X(_2382_));
 sg13g2_xnor2_1 _5748_ (.Y(_2383_),
    .A(_2379_),
    .B(_2382_));
 sg13g2_xnor2_1 _5749_ (.Y(_2384_),
    .A(_2376_),
    .B(_2383_));
 sg13g2_nor2_1 _5750_ (.A(_2354_),
    .B(_2384_),
    .Y(_0380_));
 sg13g2_and2_1 _5751_ (.A(_2372_),
    .B(_2373_),
    .X(_2385_));
 sg13g2_or2_1 _5752_ (.X(_2386_),
    .B(_2373_),
    .A(_2372_));
 sg13g2_o21ai_1 _5753_ (.B1(_2386_),
    .Y(_2387_),
    .A1(_2371_),
    .A2(_2385_));
 sg13g2_nand2_2 _5754_ (.Y(_2388_),
    .A(net87),
    .B(_0708_));
 sg13g2_nand2_1 _5755_ (.Y(_2389_),
    .A(_0705_),
    .B(_1211_));
 sg13g2_xor2_1 _5756_ (.B(_2389_),
    .A(_2388_),
    .X(_2390_));
 sg13g2_nand2_1 _5757_ (.Y(_2391_),
    .A(_1209_),
    .B(\mem[25][3] ));
 sg13g2_xor2_1 _5758_ (.B(_2391_),
    .A(_2390_),
    .X(_2392_));
 sg13g2_xnor2_1 _5759_ (.Y(_2393_),
    .A(_2387_),
    .B(_2392_));
 sg13g2_nand2_1 _5760_ (.Y(_2394_),
    .A(_2379_),
    .B(_2376_));
 sg13g2_nor2_1 _5761_ (.A(_2379_),
    .B(_2376_),
    .Y(_2395_));
 sg13g2_a21oi_1 _5762_ (.A1(_2380_),
    .A2(_2394_),
    .Y(_2396_),
    .B1(_2395_));
 sg13g2_inv_1 _5763_ (.Y(_2397_),
    .A(_2381_));
 sg13g2_nor3_1 _5764_ (.A(_2380_),
    .B(_2397_),
    .C(_2394_),
    .Y(_2398_));
 sg13g2_a21oi_1 _5765_ (.A1(_2380_),
    .A2(_2395_),
    .Y(_2399_),
    .B1(_2398_));
 sg13g2_o21ai_1 _5766_ (.B1(_2399_),
    .Y(_2400_),
    .A1(_2381_),
    .A2(_2396_));
 sg13g2_xor2_1 _5767_ (.B(_2400_),
    .A(_2393_),
    .X(_2401_));
 sg13g2_nor2_1 _5768_ (.A(_2354_),
    .B(_2401_),
    .Y(_0381_));
 sg13g2_and2_1 _5769_ (.A(_2376_),
    .B(_2381_),
    .X(_2402_));
 sg13g2_o21ai_1 _5770_ (.B1(_2379_),
    .Y(_2403_),
    .A1(_2376_),
    .A2(_2381_));
 sg13g2_nand2b_1 _5771_ (.Y(_2404_),
    .B(_2403_),
    .A_N(_2402_));
 sg13g2_o21ai_1 _5772_ (.B1(_2379_),
    .Y(_2405_),
    .A1(_2393_),
    .A2(_2402_));
 sg13g2_o21ai_1 _5773_ (.B1(_2393_),
    .Y(_2406_),
    .A1(_2376_),
    .A2(_2381_));
 sg13g2_a21oi_1 _5774_ (.A1(_2405_),
    .A2(_2406_),
    .Y(_2407_),
    .B1(_2380_));
 sg13g2_a21oi_1 _5775_ (.A1(_2393_),
    .A2(_2404_),
    .Y(_2408_),
    .B1(_2407_));
 sg13g2_nor2_1 _5776_ (.A(_2387_),
    .B(_2390_),
    .Y(_2409_));
 sg13g2_a22oi_1 _5777_ (.Y(_2410_),
    .B1(_2387_),
    .B2(_2390_),
    .A2(net124),
    .A1(_1209_));
 sg13g2_nor2_1 _5778_ (.A(_2409_),
    .B(_2410_),
    .Y(_2411_));
 sg13g2_o21ai_1 _5779_ (.B1(net87),
    .Y(_2412_),
    .A1(_0705_),
    .A2(net124));
 sg13g2_nand3_1 _5780_ (.B(_1211_),
    .C(_2412_),
    .A(_0708_),
    .Y(_2413_));
 sg13g2_nand3_1 _5781_ (.B(_0708_),
    .C(_1211_),
    .A(_0706_),
    .Y(_2414_));
 sg13g2_nand3_1 _5782_ (.B(net124),
    .C(_2414_),
    .A(net87),
    .Y(_2415_));
 sg13g2_and2_1 _5783_ (.A(_2413_),
    .B(_2415_),
    .X(_2416_));
 sg13g2_nor2b_1 _5784_ (.A(_2411_),
    .B_N(_2416_),
    .Y(_2417_));
 sg13g2_or3_1 _5785_ (.A(_2409_),
    .B(_2410_),
    .C(_2416_),
    .X(_2418_));
 sg13g2_nand2b_1 _5786_ (.Y(_2419_),
    .B(_2418_),
    .A_N(_2417_));
 sg13g2_xnor2_1 _5787_ (.Y(_2420_),
    .A(_2408_),
    .B(_2419_));
 sg13g2_nor2_1 _5788_ (.A(_2354_),
    .B(_2420_),
    .Y(_0382_));
 sg13g2_a21oi_2 _5789_ (.B1(_2417_),
    .Y(_2421_),
    .A2(_2418_),
    .A1(_2408_));
 sg13g2_inv_1 _5790_ (.Y(_2422_),
    .A(_1211_));
 sg13g2_nor3_1 _5791_ (.A(_0706_),
    .B(net124),
    .C(_2388_),
    .Y(_2423_));
 sg13g2_a21oi_1 _5792_ (.A1(net124),
    .A2(_2388_),
    .Y(_2424_),
    .B1(_2423_));
 sg13g2_nor2_1 _5793_ (.A(_2422_),
    .B(_2424_),
    .Y(_2425_));
 sg13g2_xnor2_1 _5794_ (.Y(_2426_),
    .A(_2421_),
    .B(_2425_));
 sg13g2_nor2_1 _5795_ (.A(_2354_),
    .B(_2426_),
    .Y(_0383_));
 sg13g2_a21oi_1 _5796_ (.A1(_0705_),
    .A2(_2421_),
    .Y(_2427_),
    .B1(net124));
 sg13g2_nor2_1 _5797_ (.A(_2388_),
    .B(_2427_),
    .Y(_2428_));
 sg13g2_a21oi_1 _5798_ (.A1(net124),
    .A2(_2421_),
    .Y(_2429_),
    .B1(_2428_));
 sg13g2_nor3_1 _5799_ (.A(_2422_),
    .B(_2354_),
    .C(_2429_),
    .Y(_0384_));
 sg13g2_nor2_1 _5800_ (.A(net174),
    .B(net173),
    .Y(_2430_));
 sg13g2_a21o_1 _5801_ (.A2(_2430_),
    .A1(net81),
    .B1(net54),
    .X(_2431_));
 sg13g2_buf_2 _5802_ (.A(_2431_),
    .X(_2432_));
 sg13g2_nand2_1 _5803_ (.Y(_2433_),
    .A(net123),
    .B(net172));
 sg13g2_nor2_1 _5804_ (.A(_2432_),
    .B(_2433_),
    .Y(_0385_));
 sg13g2_nand2_1 _5805_ (.Y(_2434_),
    .A(_0712_),
    .B(net172));
 sg13g2_nand2_1 _5806_ (.Y(_2435_),
    .A(net123),
    .B(_0568_));
 sg13g2_xnor2_1 _5807_ (.Y(_2436_),
    .A(_2434_),
    .B(_2435_));
 sg13g2_nor2_1 _5808_ (.A(_2432_),
    .B(_2436_),
    .Y(_0386_));
 sg13g2_nand2_1 _5809_ (.Y(_2437_),
    .A(_0568_),
    .B(_0712_));
 sg13g2_buf_2 _5810_ (.A(_2437_),
    .X(_2438_));
 sg13g2_nand2_1 _5811_ (.Y(_2439_),
    .A(net170),
    .B(_2438_));
 sg13g2_xor2_1 _5812_ (.B(_0715_),
    .A(net170),
    .X(_2440_));
 sg13g2_nand2_1 _5813_ (.Y(_2441_),
    .A(net172),
    .B(_2440_));
 sg13g2_o21ai_1 _5814_ (.B1(_2441_),
    .Y(_2442_),
    .A1(net172),
    .A2(_2439_));
 sg13g2_nand2_2 _5815_ (.Y(_2443_),
    .A(net172),
    .B(_0715_));
 sg13g2_nor2_1 _5816_ (.A(net123),
    .B(_2443_),
    .Y(_2444_));
 sg13g2_nand2b_1 _5817_ (.Y(_2445_),
    .B(_2443_),
    .A_N(net123));
 sg13g2_or2_1 _5818_ (.X(_2446_),
    .B(_0569_),
    .A(net172));
 sg13g2_a21oi_1 _5819_ (.A1(_2445_),
    .A2(_2446_),
    .Y(_2447_),
    .B1(_2438_));
 sg13g2_a221oi_1 _5820_ (.B2(_2438_),
    .C1(_2447_),
    .B1(_2444_),
    .A1(net123),
    .Y(_2448_),
    .A2(_2442_));
 sg13g2_nor2_1 _5821_ (.A(_2432_),
    .B(_2448_),
    .Y(_0387_));
 sg13g2_nand2_1 _5822_ (.Y(_2449_),
    .A(net123),
    .B(_0570_));
 sg13g2_nand2_1 _5823_ (.Y(_2450_),
    .A(_0712_),
    .B(net170));
 sg13g2_nand2_1 _5824_ (.Y(_2451_),
    .A(_0568_),
    .B(_0715_));
 sg13g2_xor2_1 _5825_ (.B(_2451_),
    .A(_2450_),
    .X(_2452_));
 sg13g2_xnor2_1 _5826_ (.Y(_2453_),
    .A(_2449_),
    .B(_2452_));
 sg13g2_buf_1 _5827_ (.A(_2453_),
    .X(_2454_));
 sg13g2_nor2_1 _5828_ (.A(_2438_),
    .B(_2443_),
    .Y(_2455_));
 sg13g2_a21oi_1 _5829_ (.A1(_0710_),
    .A2(_0569_),
    .Y(_2456_),
    .B1(_2455_));
 sg13g2_a21oi_2 _5830_ (.B1(_2456_),
    .Y(_2457_),
    .A2(_2443_),
    .A1(_2438_));
 sg13g2_nand2_2 _5831_ (.Y(_2458_),
    .A(_0559_),
    .B(net122));
 sg13g2_nor3_2 _5832_ (.A(_2433_),
    .B(_2440_),
    .C(_2438_),
    .Y(_2459_));
 sg13g2_xor2_1 _5833_ (.B(_2459_),
    .A(_2458_),
    .X(_2460_));
 sg13g2_xnor2_1 _5834_ (.Y(_2461_),
    .A(_2457_),
    .B(_2460_));
 sg13g2_xnor2_1 _5835_ (.Y(_2462_),
    .A(_2454_),
    .B(_2461_));
 sg13g2_nor2_1 _5836_ (.A(_2432_),
    .B(_2462_),
    .Y(_0388_));
 sg13g2_and2_1 _5837_ (.A(_2450_),
    .B(_2451_),
    .X(_2463_));
 sg13g2_or2_1 _5838_ (.X(_2464_),
    .B(_2451_),
    .A(_2450_));
 sg13g2_o21ai_1 _5839_ (.B1(_2464_),
    .Y(_2465_),
    .A1(_2449_),
    .A2(_2463_));
 sg13g2_nand2_2 _5840_ (.Y(_2466_),
    .A(net170),
    .B(_0715_));
 sg13g2_nand2_1 _5841_ (.Y(_2467_),
    .A(_0712_),
    .B(_0570_));
 sg13g2_xor2_1 _5842_ (.B(_2467_),
    .A(_2466_),
    .X(_2468_));
 sg13g2_nand2_1 _5843_ (.Y(_2469_),
    .A(_0568_),
    .B(\mem[26][3] ));
 sg13g2_xor2_1 _5844_ (.B(_2469_),
    .A(_2468_),
    .X(_2470_));
 sg13g2_xnor2_1 _5845_ (.Y(_2471_),
    .A(_2465_),
    .B(_2470_));
 sg13g2_nand2_1 _5846_ (.Y(_2472_),
    .A(_2457_),
    .B(_2454_));
 sg13g2_nor2_1 _5847_ (.A(_2457_),
    .B(_2454_),
    .Y(_2473_));
 sg13g2_a21oi_1 _5848_ (.A1(_2458_),
    .A2(_2472_),
    .Y(_2474_),
    .B1(_2473_));
 sg13g2_inv_1 _5849_ (.Y(_2475_),
    .A(_2459_));
 sg13g2_nor3_1 _5850_ (.A(_2458_),
    .B(_2475_),
    .C(_2472_),
    .Y(_2476_));
 sg13g2_a21oi_1 _5851_ (.A1(_2458_),
    .A2(_2473_),
    .Y(_2477_),
    .B1(_2476_));
 sg13g2_o21ai_1 _5852_ (.B1(_2477_),
    .Y(_2478_),
    .A1(_2459_),
    .A2(_2474_));
 sg13g2_xor2_1 _5853_ (.B(_2478_),
    .A(_2471_),
    .X(_2479_));
 sg13g2_nor2_1 _5854_ (.A(_2432_),
    .B(_2479_),
    .Y(_0389_));
 sg13g2_and2_1 _5855_ (.A(_2454_),
    .B(_2459_),
    .X(_2480_));
 sg13g2_o21ai_1 _5856_ (.B1(_2457_),
    .Y(_2481_),
    .A1(_2454_),
    .A2(_2459_));
 sg13g2_nand2b_1 _5857_ (.Y(_2482_),
    .B(_2481_),
    .A_N(_2480_));
 sg13g2_o21ai_1 _5858_ (.B1(_2457_),
    .Y(_2483_),
    .A1(_2471_),
    .A2(_2480_));
 sg13g2_o21ai_1 _5859_ (.B1(_2471_),
    .Y(_2484_),
    .A1(_2454_),
    .A2(_2459_));
 sg13g2_a21oi_1 _5860_ (.A1(_2483_),
    .A2(_2484_),
    .Y(_2485_),
    .B1(_2458_));
 sg13g2_a21oi_1 _5861_ (.A1(_2471_),
    .A2(_2482_),
    .Y(_2486_),
    .B1(_2485_));
 sg13g2_nor2_1 _5862_ (.A(_2465_),
    .B(_2468_),
    .Y(_2487_));
 sg13g2_a22oi_1 _5863_ (.Y(_2488_),
    .B1(_2465_),
    .B2(_2468_),
    .A2(net122),
    .A1(_0568_));
 sg13g2_nor2_1 _5864_ (.A(_2487_),
    .B(_2488_),
    .Y(_2489_));
 sg13g2_o21ai_1 _5865_ (.B1(net170),
    .Y(_2490_),
    .A1(_0712_),
    .A2(net122));
 sg13g2_nand3_1 _5866_ (.B(_0570_),
    .C(_2490_),
    .A(_0715_),
    .Y(_2491_));
 sg13g2_nand3_1 _5867_ (.B(_0715_),
    .C(_0570_),
    .A(_0713_),
    .Y(_2492_));
 sg13g2_nand3_1 _5868_ (.B(net122),
    .C(_2492_),
    .A(net170),
    .Y(_2493_));
 sg13g2_and2_1 _5869_ (.A(_2491_),
    .B(_2493_),
    .X(_2494_));
 sg13g2_nor2b_1 _5870_ (.A(_2489_),
    .B_N(_2494_),
    .Y(_2495_));
 sg13g2_or3_1 _5871_ (.A(_2487_),
    .B(_2488_),
    .C(_2494_),
    .X(_2496_));
 sg13g2_nand2b_1 _5872_ (.Y(_2497_),
    .B(_2496_),
    .A_N(_2495_));
 sg13g2_xnor2_1 _5873_ (.Y(_2498_),
    .A(_2486_),
    .B(_2497_));
 sg13g2_nor2_1 _5874_ (.A(_2432_),
    .B(_2498_),
    .Y(_0390_));
 sg13g2_a21oi_2 _5875_ (.B1(_2495_),
    .Y(_2499_),
    .A2(_2496_),
    .A1(_2486_));
 sg13g2_inv_1 _5876_ (.Y(_2500_),
    .A(_0570_));
 sg13g2_nor3_1 _5877_ (.A(_0713_),
    .B(net122),
    .C(_2466_),
    .Y(_2501_));
 sg13g2_a21oi_1 _5878_ (.A1(net122),
    .A2(_2466_),
    .Y(_2502_),
    .B1(_2501_));
 sg13g2_nor2_1 _5879_ (.A(_2500_),
    .B(_2502_),
    .Y(_2503_));
 sg13g2_xnor2_1 _5880_ (.Y(_2504_),
    .A(_2499_),
    .B(_2503_));
 sg13g2_nor2_1 _5881_ (.A(_2432_),
    .B(_2504_),
    .Y(_0391_));
 sg13g2_a21oi_1 _5882_ (.A1(_0712_),
    .A2(_2499_),
    .Y(_2505_),
    .B1(net122));
 sg13g2_nor2_1 _5883_ (.A(_2466_),
    .B(_2505_),
    .Y(_2506_));
 sg13g2_a21oi_1 _5884_ (.A1(_0716_),
    .A2(_2499_),
    .Y(_2507_),
    .B1(_2506_));
 sg13g2_nor3_1 _5885_ (.A(_2500_),
    .B(_2432_),
    .C(_2507_),
    .Y(_0392_));
 sg13g2_inv_1 _5886_ (.Y(_2508_),
    .A(net1));
 sg13g2_a21oi_1 _5887_ (.A1(_2508_),
    .A2(net2),
    .Y(_2509_),
    .B1(_2607_));
 sg13g2_nor3_1 _5888_ (.A(_2608_),
    .B(net86),
    .C(_2509_),
    .Y(_0393_));
 sg13g2_nor2_1 _5889_ (.A(net1),
    .B(net2),
    .Y(read_operation));
 sg13g2_buf_2 _5890_ (.A(net166),
    .X(_2510_));
 sg13g2_buf_1 _5891_ (.A(_2636_),
    .X(_2511_));
 sg13g2_buf_1 _5892_ (.A(net85),
    .X(_2512_));
 sg13g2_mux4_1 _5893_ (.S0(net74),
    .A0(net175),
    .A1(net144),
    .A2(net114),
    .A3(net100),
    .S1(net73),
    .X(_2513_));
 sg13g2_buf_2 _5894_ (.A(net166),
    .X(_2514_));
 sg13g2_buf_1 _5895_ (.A(net85),
    .X(_2515_));
 sg13g2_mux4_1 _5896_ (.S0(net72),
    .A0(net98),
    .A1(net96),
    .A2(_1192_),
    .A3(net92),
    .S1(net71),
    .X(_2516_));
 sg13g2_buf_2 _5897_ (.A(_2635_),
    .X(_2517_));
 sg13g2_buf_1 _5898_ (.A(net85),
    .X(_2518_));
 sg13g2_mux4_1 _5899_ (.S0(net84),
    .A0(net90),
    .A1(net88),
    .A2(net172),
    .A3(_1321_),
    .S1(net70),
    .X(_2519_));
 sg13g2_buf_1 _5900_ (.A(net166),
    .X(_2520_));
 sg13g2_mux4_1 _5901_ (.S0(net85),
    .A0(net167),
    .A1(net162),
    .A2(net164),
    .A3(net160),
    .S1(net69),
    .X(_2521_));
 sg13g2_buf_2 _5902_ (.A(net169),
    .X(_2522_));
 sg13g2_buf_1 _5903_ (.A(net171),
    .X(_2523_));
 sg13g2_mux4_1 _5904_ (.S0(net68),
    .A0(_2513_),
    .A1(_2516_),
    .A2(_2519_),
    .A3(_2521_),
    .S1(net67),
    .X(_2524_));
 sg13g2_mux4_1 _5905_ (.S0(net72),
    .A0(net158),
    .A1(net156),
    .A2(net152),
    .A3(_0644_),
    .S1(_2515_),
    .X(_2525_));
 sg13g2_mux4_1 _5906_ (.S0(net69),
    .A0(net142),
    .A1(_0672_),
    .A2(net134),
    .A3(net130),
    .S1(net71),
    .X(_2526_));
 sg13g2_buf_1 _5907_ (.A(net85),
    .X(_2527_));
 sg13g2_mux4_1 _5908_ (.S0(net74),
    .A0(_0693_),
    .A1(_0703_),
    .A2(net123),
    .A3(_0717_),
    .S1(net66),
    .X(_2528_));
 sg13g2_buf_2 _5909_ (.A(_2636_),
    .X(_2529_));
 sg13g2_mux4_1 _5910_ (.S0(net83),
    .A0(net120),
    .A1(net112),
    .A2(net116),
    .A3(net108),
    .S1(net69),
    .X(_2530_));
 sg13g2_mux4_1 _5911_ (.S0(net68),
    .A0(_2525_),
    .A1(_2526_),
    .A2(_2528_),
    .A3(_2530_),
    .S1(net67),
    .X(_2531_));
 sg13g2_mux4_1 _5912_ (.S0(_2517_),
    .A0(net104),
    .A1(net17),
    .A2(net21),
    .A3(\mem[35][0] ),
    .S1(net70),
    .X(_2532_));
 sg13g2_buf_2 _5913_ (.A(_0586_),
    .X(_2533_));
 sg13g2_mux4_1 _5914_ (.S0(net65),
    .A0(\mem[36][0] ),
    .A1(\mem[37][0] ),
    .A2(\mem[38][0] ),
    .A3(\mem[39][0] ),
    .S1(net66),
    .X(_2534_));
 sg13g2_mux4_1 _5915_ (.S0(net166),
    .A0(\mem[40][0] ),
    .A1(\mem[41][0] ),
    .A2(\mem[42][0] ),
    .A3(\mem[43][0] ),
    .S1(net83),
    .X(_2535_));
 sg13g2_buf_2 _5916_ (.A(_2635_),
    .X(_2536_));
 sg13g2_buf_1 _5917_ (.A(net85),
    .X(_2537_));
 sg13g2_mux4_1 _5918_ (.S0(net82),
    .A0(\mem[44][0] ),
    .A1(\mem[45][0] ),
    .A2(\mem[46][0] ),
    .A3(\mem[47][0] ),
    .S1(net64),
    .X(_2538_));
 sg13g2_mux4_1 _5919_ (.S0(net169),
    .A0(_2532_),
    .A1(_2534_),
    .A2(_2535_),
    .A3(_2538_),
    .S1(net171),
    .X(_2539_));
 sg13g2_mux4_1 _5920_ (.S0(net65),
    .A0(\mem[48][0] ),
    .A1(\mem[49][0] ),
    .A2(\mem[50][0] ),
    .A3(\mem[51][0] ),
    .S1(net66),
    .X(_2540_));
 sg13g2_mux4_1 _5921_ (.S0(net74),
    .A0(\mem[52][0] ),
    .A1(\mem[53][0] ),
    .A2(\mem[54][0] ),
    .A3(\mem[55][0] ),
    .S1(net73),
    .X(_2541_));
 sg13g2_mux4_1 _5922_ (.S0(net82),
    .A0(\mem[56][0] ),
    .A1(\mem[57][0] ),
    .A2(\mem[58][0] ),
    .A3(\mem[59][0] ),
    .S1(net64),
    .X(_2542_));
 sg13g2_mux4_1 _5923_ (.S0(net84),
    .A0(\mem[60][0] ),
    .A1(\mem[61][0] ),
    .A2(\mem[62][0] ),
    .A3(\mem[63][0] ),
    .S1(net64),
    .X(_2543_));
 sg13g2_mux4_1 _5924_ (.S0(net68),
    .A0(_2540_),
    .A1(_2541_),
    .A2(_2542_),
    .A3(_2543_),
    .S1(net67),
    .X(_2544_));
 sg13g2_mux4_1 _5925_ (.S0(net177),
    .A0(_2524_),
    .A1(_2531_),
    .A2(_2539_),
    .A3(_2544_),
    .S1(net176),
    .X(net11));
 sg13g2_mux4_1 _5926_ (.S0(net74),
    .A0(_2722_),
    .A1(_0659_),
    .A2(_0746_),
    .A3(_1139_),
    .S1(net73),
    .X(_2545_));
 sg13g2_mux4_1 _5927_ (.S0(net72),
    .A0(_1164_),
    .A1(_1185_),
    .A2(_1194_),
    .A3(_1199_),
    .S1(net71),
    .X(_2546_));
 sg13g2_mux4_1 _5928_ (.S0(net84),
    .A0(_1204_),
    .A1(_1209_),
    .A2(_0568_),
    .A3(_0580_),
    .S1(net70),
    .X(_2547_));
 sg13g2_mux4_1 _5929_ (.S0(net85),
    .A0(_0591_),
    .A1(_0606_),
    .A2(_0599_),
    .A3(_0613_),
    .S1(net69),
    .X(_2548_));
 sg13g2_mux4_1 _5930_ (.S0(net68),
    .A0(_2545_),
    .A1(_2546_),
    .A2(_2547_),
    .A3(_2548_),
    .S1(net67),
    .X(_2549_));
 sg13g2_mux4_1 _5931_ (.S0(net72),
    .A0(_0621_),
    .A1(net155),
    .A2(net151),
    .A3(_0646_),
    .S1(_2515_),
    .X(_2550_));
 sg13g2_mux4_1 _5932_ (.S0(net69),
    .A0(net141),
    .A1(_0674_),
    .A2(_0681_),
    .A3(_0688_),
    .S1(net71),
    .X(_2551_));
 sg13g2_mux4_1 _5933_ (.S0(net74),
    .A0(_0698_),
    .A1(_0705_),
    .A2(_0712_),
    .A3(_1322_),
    .S1(net66),
    .X(_2552_));
 sg13g2_mux4_1 _5934_ (.S0(net83),
    .A0(net119),
    .A1(net111),
    .A2(_0737_),
    .A3(_0759_),
    .S1(net69),
    .X(_2553_));
 sg13g2_mux4_1 _5935_ (.S0(net68),
    .A0(_2550_),
    .A1(_2551_),
    .A2(_2552_),
    .A3(_2553_),
    .S1(net67),
    .X(_2554_));
 sg13g2_mux4_1 _5936_ (.S0(_2517_),
    .A0(net103),
    .A1(net18),
    .A2(net22),
    .A3(\mem[35][1] ),
    .S1(net70),
    .X(_2555_));
 sg13g2_mux4_1 _5937_ (.S0(net65),
    .A0(\mem[36][1] ),
    .A1(\mem[37][1] ),
    .A2(\mem[38][1] ),
    .A3(\mem[39][1] ),
    .S1(net66),
    .X(_2556_));
 sg13g2_mux4_1 _5938_ (.S0(net166),
    .A0(\mem[40][1] ),
    .A1(\mem[41][1] ),
    .A2(\mem[42][1] ),
    .A3(\mem[43][1] ),
    .S1(net83),
    .X(_2557_));
 sg13g2_mux4_1 _5939_ (.S0(net82),
    .A0(\mem[44][1] ),
    .A1(\mem[45][1] ),
    .A2(\mem[46][1] ),
    .A3(\mem[47][1] ),
    .S1(net64),
    .X(_2558_));
 sg13g2_mux4_1 _5940_ (.S0(net169),
    .A0(_2555_),
    .A1(_2556_),
    .A2(_2557_),
    .A3(_2558_),
    .S1(net171),
    .X(_2559_));
 sg13g2_mux4_1 _5941_ (.S0(net65),
    .A0(\mem[48][1] ),
    .A1(\mem[49][1] ),
    .A2(\mem[50][1] ),
    .A3(\mem[51][1] ),
    .S1(net66),
    .X(_2560_));
 sg13g2_mux4_1 _5942_ (.S0(net74),
    .A0(\mem[52][1] ),
    .A1(\mem[53][1] ),
    .A2(\mem[54][1] ),
    .A3(\mem[55][1] ),
    .S1(net73),
    .X(_2561_));
 sg13g2_mux4_1 _5943_ (.S0(net82),
    .A0(\mem[56][1] ),
    .A1(\mem[57][1] ),
    .A2(\mem[58][1] ),
    .A3(\mem[59][1] ),
    .S1(net64),
    .X(_2562_));
 sg13g2_mux4_1 _5944_ (.S0(net84),
    .A0(\mem[60][1] ),
    .A1(\mem[61][1] ),
    .A2(\mem[62][1] ),
    .A3(\mem[63][1] ),
    .S1(net64),
    .X(_2563_));
 sg13g2_mux4_1 _5945_ (.S0(net68),
    .A0(_2560_),
    .A1(_2561_),
    .A2(_2562_),
    .A3(_2563_),
    .S1(net67),
    .X(_2564_));
 sg13g2_mux4_1 _5946_ (.S0(net177),
    .A0(_2549_),
    .A1(_2554_),
    .A2(_2559_),
    .A3(_2564_),
    .S1(net176),
    .X(net12));
 sg13g2_mux4_1 _5947_ (.S0(_2510_),
    .A0(_0427_),
    .A1(net143),
    .A2(net113),
    .A3(_1140_),
    .S1(net73),
    .X(_2565_));
 sg13g2_mux4_1 _5948_ (.S0(net72),
    .A0(net97),
    .A1(_1186_),
    .A2(_1195_),
    .A3(net91),
    .S1(net71),
    .X(_2566_));
 sg13g2_mux4_1 _5949_ (.S0(net84),
    .A0(net89),
    .A1(net87),
    .A2(net170),
    .A3(_0583_),
    .S1(_2518_),
    .X(_2567_));
 sg13g2_mux4_1 _5950_ (.S0(net85),
    .A0(net165),
    .A1(net161),
    .A2(net163),
    .A3(net159),
    .S1(net69),
    .X(_2568_));
 sg13g2_mux4_1 _5951_ (.S0(net68),
    .A0(_2565_),
    .A1(_2566_),
    .A2(_2567_),
    .A3(_2568_),
    .S1(net67),
    .X(_2569_));
 sg13g2_mux4_1 _5952_ (.S0(_2514_),
    .A0(net157),
    .A1(net154),
    .A2(net150),
    .A3(_0651_),
    .S1(net73),
    .X(_2570_));
 sg13g2_mux4_1 _5953_ (.S0(net72),
    .A0(net140),
    .A1(net136),
    .A2(net132),
    .A3(_0691_),
    .S1(net71),
    .X(_2571_));
 sg13g2_mux4_1 _5954_ (.S0(_2533_),
    .A0(_0701_),
    .A1(_0708_),
    .A2(_0715_),
    .A3(net78),
    .S1(_2527_),
    .X(_2572_));
 sg13g2_mux4_1 _5955_ (.S0(_2529_),
    .A0(net118),
    .A1(net110),
    .A2(_0741_),
    .A3(net106),
    .S1(net69),
    .X(_2573_));
 sg13g2_mux4_1 _5956_ (.S0(net68),
    .A0(_2570_),
    .A1(_2571_),
    .A2(_2572_),
    .A3(_2573_),
    .S1(net67),
    .X(_2574_));
 sg13g2_mux4_1 _5957_ (.S0(net84),
    .A0(net102),
    .A1(net19),
    .A2(net23),
    .A3(\mem[35][2] ),
    .S1(net70),
    .X(_2575_));
 sg13g2_mux4_1 _5958_ (.S0(net65),
    .A0(\mem[36][2] ),
    .A1(\mem[37][2] ),
    .A2(\mem[38][2] ),
    .A3(\mem[39][2] ),
    .S1(net66),
    .X(_2576_));
 sg13g2_mux4_1 _5959_ (.S0(net166),
    .A0(\mem[40][2] ),
    .A1(\mem[41][2] ),
    .A2(\mem[42][2] ),
    .A3(\mem[43][2] ),
    .S1(net83),
    .X(_2577_));
 sg13g2_mux4_1 _5960_ (.S0(net82),
    .A0(\mem[44][2] ),
    .A1(\mem[45][2] ),
    .A2(\mem[46][2] ),
    .A3(\mem[47][2] ),
    .S1(net64),
    .X(_2578_));
 sg13g2_mux4_1 _5961_ (.S0(net169),
    .A0(_2575_),
    .A1(_2576_),
    .A2(_2577_),
    .A3(_2578_),
    .S1(_0563_),
    .X(_2579_));
 sg13g2_mux4_1 _5962_ (.S0(net65),
    .A0(\mem[48][2] ),
    .A1(\mem[49][2] ),
    .A2(\mem[50][2] ),
    .A3(\mem[51][2] ),
    .S1(net70),
    .X(_2580_));
 sg13g2_mux4_1 _5963_ (.S0(net74),
    .A0(\mem[52][2] ),
    .A1(\mem[53][2] ),
    .A2(\mem[54][2] ),
    .A3(\mem[55][2] ),
    .S1(net73),
    .X(_2581_));
 sg13g2_mux4_1 _5964_ (.S0(net82),
    .A0(\mem[56][2] ),
    .A1(\mem[57][2] ),
    .A2(\mem[58][2] ),
    .A3(\mem[59][2] ),
    .S1(net83),
    .X(_2582_));
 sg13g2_mux4_1 _5965_ (.S0(_2536_),
    .A0(\mem[60][2] ),
    .A1(\mem[61][2] ),
    .A2(\mem[62][2] ),
    .A3(\mem[63][2] ),
    .S1(_2537_),
    .X(_2583_));
 sg13g2_mux4_1 _5966_ (.S0(net169),
    .A0(_2580_),
    .A1(_2581_),
    .A2(_2582_),
    .A3(_2583_),
    .S1(net171),
    .X(_2584_));
 sg13g2_mux4_1 _5967_ (.S0(net177),
    .A0(_2569_),
    .A1(_2574_),
    .A2(_2579_),
    .A3(_2584_),
    .S1(net176),
    .X(net13));
 sg13g2_mux4_1 _5968_ (.S0(_2510_),
    .A0(_0558_),
    .A1(_0662_),
    .A2(_0748_),
    .A3(_1141_),
    .S1(_2512_),
    .X(_2585_));
 sg13g2_mux4_1 _5969_ (.S0(net72),
    .A0(_1166_),
    .A1(_1187_),
    .A2(_1196_),
    .A3(_1201_),
    .S1(net71),
    .X(_2586_));
 sg13g2_mux4_1 _5970_ (.S0(net84),
    .A0(_1206_),
    .A1(_1211_),
    .A2(_0570_),
    .A3(_0584_),
    .S1(_2518_),
    .X(_2587_));
 sg13g2_mux4_1 _5971_ (.S0(_2511_),
    .A0(_0593_),
    .A1(_0608_),
    .A2(_0601_),
    .A3(_0615_),
    .S1(_2520_),
    .X(_2588_));
 sg13g2_mux4_1 _5972_ (.S0(_2522_),
    .A0(_2585_),
    .A1(_2586_),
    .A2(_2587_),
    .A3(_2588_),
    .S1(_2523_),
    .X(_2589_));
 sg13g2_mux4_1 _5973_ (.S0(_2514_),
    .A0(_0623_),
    .A1(_0636_),
    .A2(net149),
    .A3(_0653_),
    .S1(_2512_),
    .X(_2590_));
 sg13g2_mux4_1 _5974_ (.S0(net72),
    .A0(_0671_),
    .A1(net135),
    .A2(_0685_),
    .A3(net128),
    .S1(net71),
    .X(_2591_));
 sg13g2_mux4_1 _5975_ (.S0(_2533_),
    .A0(_0702_),
    .A1(_0709_),
    .A2(_0716_),
    .A3(net77),
    .S1(_2527_),
    .X(_2592_));
 sg13g2_mux4_1 _5976_ (.S0(_2529_),
    .A0(net117),
    .A1(net109),
    .A2(net115),
    .A3(_0763_),
    .S1(_2520_),
    .X(_2593_));
 sg13g2_mux4_1 _5977_ (.S0(_2522_),
    .A0(_2590_),
    .A1(_2591_),
    .A2(_2592_),
    .A3(_2593_),
    .S1(_2523_),
    .X(_2594_));
 sg13g2_mux4_1 _5978_ (.S0(net84),
    .A0(net101),
    .A1(net20),
    .A2(net24),
    .A3(\mem[35][3] ),
    .S1(net70),
    .X(_2595_));
 sg13g2_mux4_1 _5979_ (.S0(net65),
    .A0(\mem[36][3] ),
    .A1(\mem[37][3] ),
    .A2(\mem[38][3] ),
    .A3(\mem[39][3] ),
    .S1(net66),
    .X(_2596_));
 sg13g2_mux4_1 _5980_ (.S0(net166),
    .A0(\mem[40][3] ),
    .A1(\mem[41][3] ),
    .A2(\mem[42][3] ),
    .A3(\mem[43][3] ),
    .S1(net83),
    .X(_2597_));
 sg13g2_mux4_1 _5981_ (.S0(net82),
    .A0(\mem[44][3] ),
    .A1(\mem[45][3] ),
    .A2(\mem[46][3] ),
    .A3(\mem[47][3] ),
    .S1(net64),
    .X(_2598_));
 sg13g2_mux4_1 _5982_ (.S0(net169),
    .A0(_2595_),
    .A1(_2596_),
    .A2(_2597_),
    .A3(_2598_),
    .S1(_0563_),
    .X(_2599_));
 sg13g2_mux4_1 _5983_ (.S0(net65),
    .A0(\mem[48][3] ),
    .A1(\mem[49][3] ),
    .A2(\mem[50][3] ),
    .A3(\mem[51][3] ),
    .S1(net70),
    .X(_2600_));
 sg13g2_mux4_1 _5984_ (.S0(net74),
    .A0(\mem[52][3] ),
    .A1(\mem[53][3] ),
    .A2(\mem[54][3] ),
    .A3(\mem[55][3] ),
    .S1(net73),
    .X(_2601_));
 sg13g2_mux4_1 _5985_ (.S0(net82),
    .A0(\mem[56][3] ),
    .A1(\mem[57][3] ),
    .A2(\mem[58][3] ),
    .A3(\mem[59][3] ),
    .S1(net83),
    .X(_2602_));
 sg13g2_mux4_1 _5986_ (.S0(_2536_),
    .A0(\mem[60][3] ),
    .A1(\mem[61][3] ),
    .A2(\mem[62][3] ),
    .A3(\mem[63][3] ),
    .S1(_2537_),
    .X(_2603_));
 sg13g2_mux4_1 _5987_ (.S0(net169),
    .A0(_2600_),
    .A1(_2601_),
    .A2(_2602_),
    .A3(_2603_),
    .S1(net171),
    .X(_2604_));
 sg13g2_mux4_1 _5988_ (.S0(net177),
    .A0(_2589_),
    .A1(_2594_),
    .A2(_2599_),
    .A3(_2604_),
    .S1(net176),
    .X(net14));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_3_0__leaf_clk));
 sg13g2_tiehi _5995__182 (.L_HI(net182));
 sg13g2_buf_1 _5991_ (.A(read_operation),
    .X(net7));
 sg13g2_buf_1 _5992_ (.A(read_operation),
    .X(net8));
 sg13g2_buf_1 _5993_ (.A(read_operation),
    .X(net9));
 sg13g2_buf_1 _5994_ (.A(read_operation),
    .X(net10));
 sg13g2_buf_1 _5995_ (.A(net182),
    .X(uio_oe[4]));
 sg13g2_buf_1 _5996_ (.A(net183),
    .X(uio_oe[5]));
 sg13g2_buf_1 _5997_ (.A(net178),
    .X(uio_oe[6]));
 sg13g2_buf_1 _5998_ (.A(net179),
    .X(uio_oe[7]));
 sg13g2_buf_1 _5999_ (.A(net180),
    .X(uio_out[6]));
 sg13g2_buf_1 _6000_ (.A(net181),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \mem[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net184),
    .D(_0001_),
    .Q_N(_3187_),
    .Q(\mem[0][0] ));
 sg13g2_dfrbp_1 \mem[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net185),
    .D(_0002_),
    .Q_N(_0000_),
    .Q(\mem[0][1] ));
 sg13g2_dfrbp_1 \mem[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net186),
    .D(_0003_),
    .Q_N(_3186_),
    .Q(\mem[0][2] ));
 sg13g2_dfrbp_1 \mem[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net187),
    .D(_0004_),
    .Q_N(_3185_),
    .Q(\mem[0][3] ));
 sg13g2_dfrbp_1 \mem[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net188),
    .D(_0005_),
    .Q_N(_3184_),
    .Q(\mem[10][0] ));
 sg13g2_dfrbp_1 \mem[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net189),
    .D(_0006_),
    .Q_N(_3183_),
    .Q(\mem[10][1] ));
 sg13g2_dfrbp_1 \mem[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net190),
    .D(_0007_),
    .Q_N(_3182_),
    .Q(\mem[10][2] ));
 sg13g2_dfrbp_1 \mem[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net191),
    .D(_0008_),
    .Q_N(_3181_),
    .Q(\mem[10][3] ));
 sg13g2_dfrbp_1 \mem[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net192),
    .D(_0009_),
    .Q_N(_3180_),
    .Q(\mem[11][0] ));
 sg13g2_dfrbp_1 \mem[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net193),
    .D(_0010_),
    .Q_N(_3179_),
    .Q(\mem[11][1] ));
 sg13g2_dfrbp_1 \mem[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net194),
    .D(_0011_),
    .Q_N(_3178_),
    .Q(\mem[11][2] ));
 sg13g2_dfrbp_1 \mem[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net195),
    .D(_0012_),
    .Q_N(_3177_),
    .Q(\mem[11][3] ));
 sg13g2_dfrbp_1 \mem[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net196),
    .D(_0013_),
    .Q_N(_3176_),
    .Q(\mem[12][0] ));
 sg13g2_dfrbp_1 \mem[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net197),
    .D(_0014_),
    .Q_N(_3175_),
    .Q(\mem[12][1] ));
 sg13g2_dfrbp_1 \mem[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net198),
    .D(_0015_),
    .Q_N(_3174_),
    .Q(\mem[12][2] ));
 sg13g2_dfrbp_1 \mem[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net199),
    .D(_0016_),
    .Q_N(_3173_),
    .Q(\mem[12][3] ));
 sg13g2_dfrbp_1 \mem[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net200),
    .D(_0017_),
    .Q_N(_3172_),
    .Q(\mem[13][0] ));
 sg13g2_dfrbp_1 \mem[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net201),
    .D(_0018_),
    .Q_N(_3171_),
    .Q(\mem[13][1] ));
 sg13g2_dfrbp_1 \mem[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net202),
    .D(_0019_),
    .Q_N(_3170_),
    .Q(\mem[13][2] ));
 sg13g2_dfrbp_1 \mem[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net203),
    .D(_0020_),
    .Q_N(_3169_),
    .Q(\mem[13][3] ));
 sg13g2_dfrbp_1 \mem[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net204),
    .D(_0021_),
    .Q_N(_3168_),
    .Q(\mem[14][0] ));
 sg13g2_dfrbp_1 \mem[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net205),
    .D(_0022_),
    .Q_N(_3167_),
    .Q(\mem[14][1] ));
 sg13g2_dfrbp_1 \mem[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net206),
    .D(_0023_),
    .Q_N(_3166_),
    .Q(\mem[14][2] ));
 sg13g2_dfrbp_1 \mem[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net207),
    .D(_0024_),
    .Q_N(_3165_),
    .Q(\mem[14][3] ));
 sg13g2_dfrbp_1 \mem[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net208),
    .D(_0025_),
    .Q_N(_3164_),
    .Q(\mem[15][0] ));
 sg13g2_dfrbp_1 \mem[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net209),
    .D(_0026_),
    .Q_N(_3163_),
    .Q(\mem[15][1] ));
 sg13g2_dfrbp_1 \mem[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net210),
    .D(_0027_),
    .Q_N(_3162_),
    .Q(\mem[15][2] ));
 sg13g2_dfrbp_1 \mem[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net211),
    .D(_0028_),
    .Q_N(_3161_),
    .Q(\mem[15][3] ));
 sg13g2_dfrbp_1 \mem[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net212),
    .D(_0029_),
    .Q_N(_3160_),
    .Q(\mem[16][0] ));
 sg13g2_dfrbp_1 \mem[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net213),
    .D(_0030_),
    .Q_N(_3159_),
    .Q(\mem[16][1] ));
 sg13g2_dfrbp_1 \mem[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net214),
    .D(_0031_),
    .Q_N(_3158_),
    .Q(\mem[16][2] ));
 sg13g2_dfrbp_1 \mem[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net215),
    .D(_0032_),
    .Q_N(_3157_),
    .Q(\mem[16][3] ));
 sg13g2_dfrbp_1 \mem[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net216),
    .D(_0033_),
    .Q_N(_3156_),
    .Q(\mem[17][0] ));
 sg13g2_dfrbp_1 \mem[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net217),
    .D(_0034_),
    .Q_N(_3155_),
    .Q(\mem[17][1] ));
 sg13g2_dfrbp_1 \mem[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net218),
    .D(_0035_),
    .Q_N(_3154_),
    .Q(\mem[17][2] ));
 sg13g2_dfrbp_1 \mem[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net219),
    .D(_0036_),
    .Q_N(_3153_),
    .Q(\mem[17][3] ));
 sg13g2_dfrbp_1 \mem[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net220),
    .D(_0037_),
    .Q_N(_3152_),
    .Q(\mem[18][0] ));
 sg13g2_dfrbp_1 \mem[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net221),
    .D(_0038_),
    .Q_N(_3151_),
    .Q(\mem[18][1] ));
 sg13g2_dfrbp_1 \mem[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net222),
    .D(_0039_),
    .Q_N(_3150_),
    .Q(\mem[18][2] ));
 sg13g2_dfrbp_1 \mem[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net223),
    .D(_0040_),
    .Q_N(_3149_),
    .Q(\mem[18][3] ));
 sg13g2_dfrbp_1 \mem[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net224),
    .D(_0041_),
    .Q_N(_3148_),
    .Q(\mem[19][0] ));
 sg13g2_dfrbp_1 \mem[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net225),
    .D(_0042_),
    .Q_N(_3147_),
    .Q(\mem[19][1] ));
 sg13g2_dfrbp_1 \mem[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net226),
    .D(_0043_),
    .Q_N(_3146_),
    .Q(\mem[19][2] ));
 sg13g2_dfrbp_1 \mem[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net227),
    .D(_0044_),
    .Q_N(_3145_),
    .Q(\mem[19][3] ));
 sg13g2_dfrbp_1 \mem[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net228),
    .D(_0045_),
    .Q_N(_3144_),
    .Q(\mem[1][0] ));
 sg13g2_dfrbp_1 \mem[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net229),
    .D(_0046_),
    .Q_N(_3143_),
    .Q(\mem[1][1] ));
 sg13g2_dfrbp_1 \mem[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net230),
    .D(_0047_),
    .Q_N(_3142_),
    .Q(\mem[1][2] ));
 sg13g2_dfrbp_1 \mem[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net231),
    .D(_0048_),
    .Q_N(_3141_),
    .Q(\mem[1][3] ));
 sg13g2_dfrbp_1 \mem[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net232),
    .D(_0049_),
    .Q_N(_3140_),
    .Q(\mem[20][0] ));
 sg13g2_dfrbp_1 \mem[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net233),
    .D(_0050_),
    .Q_N(_3139_),
    .Q(\mem[20][1] ));
 sg13g2_dfrbp_1 \mem[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net234),
    .D(_0051_),
    .Q_N(_3138_),
    .Q(\mem[20][2] ));
 sg13g2_dfrbp_1 \mem[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net235),
    .D(_0052_),
    .Q_N(_3137_),
    .Q(\mem[20][3] ));
 sg13g2_dfrbp_1 \mem[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net236),
    .D(_0053_),
    .Q_N(_3136_),
    .Q(\mem[21][0] ));
 sg13g2_dfrbp_1 \mem[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net237),
    .D(_0054_),
    .Q_N(_3135_),
    .Q(\mem[21][1] ));
 sg13g2_dfrbp_1 \mem[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net238),
    .D(_0055_),
    .Q_N(_3134_),
    .Q(\mem[21][2] ));
 sg13g2_dfrbp_1 \mem[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net239),
    .D(_0056_),
    .Q_N(_3133_),
    .Q(\mem[21][3] ));
 sg13g2_dfrbp_1 \mem[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net240),
    .D(_0057_),
    .Q_N(_3132_),
    .Q(\mem[22][0] ));
 sg13g2_dfrbp_1 \mem[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net241),
    .D(_0058_),
    .Q_N(_3131_),
    .Q(\mem[22][1] ));
 sg13g2_dfrbp_1 \mem[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net242),
    .D(_0059_),
    .Q_N(_3130_),
    .Q(\mem[22][2] ));
 sg13g2_dfrbp_1 \mem[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net243),
    .D(_0060_),
    .Q_N(_3129_),
    .Q(\mem[22][3] ));
 sg13g2_dfrbp_1 \mem[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net244),
    .D(_0061_),
    .Q_N(_3128_),
    .Q(\mem[23][0] ));
 sg13g2_dfrbp_1 \mem[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net245),
    .D(_0062_),
    .Q_N(_3127_),
    .Q(\mem[23][1] ));
 sg13g2_dfrbp_1 \mem[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net246),
    .D(_0063_),
    .Q_N(_3126_),
    .Q(\mem[23][2] ));
 sg13g2_dfrbp_1 \mem[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net247),
    .D(_0064_),
    .Q_N(_3125_),
    .Q(\mem[23][3] ));
 sg13g2_dfrbp_1 \mem[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net248),
    .D(_0065_),
    .Q_N(_3124_),
    .Q(\mem[24][0] ));
 sg13g2_dfrbp_1 \mem[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net249),
    .D(_0066_),
    .Q_N(_3123_),
    .Q(\mem[24][1] ));
 sg13g2_dfrbp_1 \mem[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net250),
    .D(_0067_),
    .Q_N(_3122_),
    .Q(\mem[24][2] ));
 sg13g2_dfrbp_1 \mem[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net251),
    .D(_0068_),
    .Q_N(_3121_),
    .Q(\mem[24][3] ));
 sg13g2_dfrbp_1 \mem[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net252),
    .D(_0069_),
    .Q_N(_3120_),
    .Q(\mem[25][0] ));
 sg13g2_dfrbp_1 \mem[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net253),
    .D(_0070_),
    .Q_N(_3119_),
    .Q(\mem[25][1] ));
 sg13g2_dfrbp_1 \mem[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net254),
    .D(_0071_),
    .Q_N(_3118_),
    .Q(\mem[25][2] ));
 sg13g2_dfrbp_1 \mem[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net255),
    .D(_0072_),
    .Q_N(_3117_),
    .Q(\mem[25][3] ));
 sg13g2_dfrbp_1 \mem[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net256),
    .D(_0073_),
    .Q_N(_3116_),
    .Q(\mem[26][0] ));
 sg13g2_dfrbp_1 \mem[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net257),
    .D(_0074_),
    .Q_N(_3115_),
    .Q(\mem[26][1] ));
 sg13g2_dfrbp_1 \mem[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net258),
    .D(_0075_),
    .Q_N(_3114_),
    .Q(\mem[26][2] ));
 sg13g2_dfrbp_1 \mem[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net259),
    .D(_0076_),
    .Q_N(_3113_),
    .Q(\mem[26][3] ));
 sg13g2_dfrbp_1 \mem[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net260),
    .D(_0077_),
    .Q_N(_3112_),
    .Q(\mem[27][0] ));
 sg13g2_dfrbp_1 \mem[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net261),
    .D(_0078_),
    .Q_N(_3111_),
    .Q(\mem[27][1] ));
 sg13g2_dfrbp_1 \mem[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net262),
    .D(_0079_),
    .Q_N(_3110_),
    .Q(\mem[27][2] ));
 sg13g2_dfrbp_1 \mem[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net263),
    .D(_0080_),
    .Q_N(_3109_),
    .Q(\mem[27][3] ));
 sg13g2_dfrbp_1 \mem[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net264),
    .D(_0081_),
    .Q_N(_3108_),
    .Q(\mem[28][0] ));
 sg13g2_dfrbp_1 \mem[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net265),
    .D(_0082_),
    .Q_N(_3107_),
    .Q(\mem[28][1] ));
 sg13g2_dfrbp_1 \mem[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net266),
    .D(_0083_),
    .Q_N(_3106_),
    .Q(\mem[28][2] ));
 sg13g2_dfrbp_1 \mem[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net267),
    .D(_0084_),
    .Q_N(_3105_),
    .Q(\mem[28][3] ));
 sg13g2_dfrbp_1 \mem[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net268),
    .D(_0085_),
    .Q_N(_3104_),
    .Q(\mem[29][0] ));
 sg13g2_dfrbp_1 \mem[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net269),
    .D(_0086_),
    .Q_N(_3103_),
    .Q(\mem[29][1] ));
 sg13g2_dfrbp_1 \mem[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net270),
    .D(_0087_),
    .Q_N(_3102_),
    .Q(\mem[29][2] ));
 sg13g2_dfrbp_1 \mem[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net271),
    .D(_0088_),
    .Q_N(_3101_),
    .Q(\mem[29][3] ));
 sg13g2_dfrbp_1 \mem[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net272),
    .D(_0089_),
    .Q_N(_3100_),
    .Q(\mem[2][0] ));
 sg13g2_dfrbp_1 \mem[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net273),
    .D(_0090_),
    .Q_N(_3099_),
    .Q(\mem[2][1] ));
 sg13g2_dfrbp_1 \mem[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net274),
    .D(_0091_),
    .Q_N(_3098_),
    .Q(\mem[2][2] ));
 sg13g2_dfrbp_1 \mem[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net275),
    .D(_0092_),
    .Q_N(_3097_),
    .Q(\mem[2][3] ));
 sg13g2_dfrbp_1 \mem[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net276),
    .D(_0093_),
    .Q_N(_3096_),
    .Q(\mem[30][0] ));
 sg13g2_dfrbp_1 \mem[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net277),
    .D(_0094_),
    .Q_N(_3095_),
    .Q(\mem[30][1] ));
 sg13g2_dfrbp_1 \mem[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net278),
    .D(_0095_),
    .Q_N(_3094_),
    .Q(\mem[30][2] ));
 sg13g2_dfrbp_1 \mem[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net279),
    .D(_0096_),
    .Q_N(_3093_),
    .Q(\mem[30][3] ));
 sg13g2_dfrbp_1 \mem[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net280),
    .D(_0097_),
    .Q_N(_3092_),
    .Q(\mem[31][0] ));
 sg13g2_dfrbp_1 \mem[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net281),
    .D(_0098_),
    .Q_N(_3091_),
    .Q(\mem[31][1] ));
 sg13g2_dfrbp_1 \mem[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net282),
    .D(_0099_),
    .Q_N(_3090_),
    .Q(\mem[31][2] ));
 sg13g2_dfrbp_1 \mem[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net283),
    .D(_0100_),
    .Q_N(_3089_),
    .Q(\mem[31][3] ));
 sg13g2_dfrbp_1 \mem[32][0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net284),
    .D(_0101_),
    .Q_N(_3088_),
    .Q(\mem[32][0] ));
 sg13g2_dfrbp_1 \mem[32][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net285),
    .D(_0102_),
    .Q_N(_3087_),
    .Q(\mem[32][1] ));
 sg13g2_dfrbp_1 \mem[32][2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net286),
    .D(_0103_),
    .Q_N(_3086_),
    .Q(\mem[32][2] ));
 sg13g2_dfrbp_1 \mem[32][3]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net287),
    .D(_0104_),
    .Q_N(_3085_),
    .Q(\mem[32][3] ));
 sg13g2_dfrbp_1 \mem[33][0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net288),
    .D(_0105_),
    .Q_N(_3084_),
    .Q(net17));
 sg13g2_dfrbp_1 \mem[33][1]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net289),
    .D(_0106_),
    .Q_N(_3083_),
    .Q(net18));
 sg13g2_dfrbp_1 \mem[33][2]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net290),
    .D(_0107_),
    .Q_N(_3082_),
    .Q(net19));
 sg13g2_dfrbp_1 \mem[33][3]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net291),
    .D(_0108_),
    .Q_N(_3081_),
    .Q(net20));
 sg13g2_dfrbp_1 \mem[34][0]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net292),
    .D(_0109_),
    .Q_N(_3080_),
    .Q(net21));
 sg13g2_dfrbp_1 \mem[34][1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net293),
    .D(_0110_),
    .Q_N(_3079_),
    .Q(net22));
 sg13g2_dfrbp_1 \mem[34][2]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net294),
    .D(_0111_),
    .Q_N(_3078_),
    .Q(net23));
 sg13g2_dfrbp_1 \mem[34][3]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net295),
    .D(_0112_),
    .Q_N(_3077_),
    .Q(net24));
 sg13g2_dfrbp_1 \mem[35][0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net296),
    .D(_0113_),
    .Q_N(_3076_),
    .Q(\mem[35][0] ));
 sg13g2_dfrbp_1 \mem[35][1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net297),
    .D(_0114_),
    .Q_N(_3075_),
    .Q(\mem[35][1] ));
 sg13g2_dfrbp_1 \mem[35][2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net298),
    .D(_0115_),
    .Q_N(_3074_),
    .Q(\mem[35][2] ));
 sg13g2_dfrbp_1 \mem[35][3]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net299),
    .D(_0116_),
    .Q_N(_3073_),
    .Q(\mem[35][3] ));
 sg13g2_dfrbp_1 \mem[36][0]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net300),
    .D(_0117_),
    .Q_N(_3072_),
    .Q(\mem[36][0] ));
 sg13g2_dfrbp_1 \mem[36][1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net301),
    .D(_0118_),
    .Q_N(_3071_),
    .Q(\mem[36][1] ));
 sg13g2_dfrbp_1 \mem[36][2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net302),
    .D(_0119_),
    .Q_N(_3070_),
    .Q(\mem[36][2] ));
 sg13g2_dfrbp_1 \mem[36][3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net303),
    .D(_0120_),
    .Q_N(_3069_),
    .Q(\mem[36][3] ));
 sg13g2_dfrbp_1 \mem[37][0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net304),
    .D(_0121_),
    .Q_N(_3068_),
    .Q(\mem[37][0] ));
 sg13g2_dfrbp_1 \mem[37][1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net305),
    .D(_0122_),
    .Q_N(_3067_),
    .Q(\mem[37][1] ));
 sg13g2_dfrbp_1 \mem[37][2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net306),
    .D(_0123_),
    .Q_N(_3066_),
    .Q(\mem[37][2] ));
 sg13g2_dfrbp_1 \mem[37][3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net307),
    .D(_0124_),
    .Q_N(_3065_),
    .Q(\mem[37][3] ));
 sg13g2_dfrbp_1 \mem[38][0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net308),
    .D(_0125_),
    .Q_N(_3064_),
    .Q(\mem[38][0] ));
 sg13g2_dfrbp_1 \mem[38][1]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net309),
    .D(_0126_),
    .Q_N(_3063_),
    .Q(\mem[38][1] ));
 sg13g2_dfrbp_1 \mem[38][2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net310),
    .D(_0127_),
    .Q_N(_3062_),
    .Q(\mem[38][2] ));
 sg13g2_dfrbp_1 \mem[38][3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net311),
    .D(_0128_),
    .Q_N(_3061_),
    .Q(\mem[38][3] ));
 sg13g2_dfrbp_1 \mem[39][0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net312),
    .D(_0129_),
    .Q_N(_3060_),
    .Q(\mem[39][0] ));
 sg13g2_dfrbp_1 \mem[39][1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net313),
    .D(_0130_),
    .Q_N(_3059_),
    .Q(\mem[39][1] ));
 sg13g2_dfrbp_1 \mem[39][2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net314),
    .D(_0131_),
    .Q_N(_3058_),
    .Q(\mem[39][2] ));
 sg13g2_dfrbp_1 \mem[39][3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net315),
    .D(_0132_),
    .Q_N(_3057_),
    .Q(\mem[39][3] ));
 sg13g2_dfrbp_1 \mem[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net316),
    .D(_0133_),
    .Q_N(_3056_),
    .Q(\mem[3][0] ));
 sg13g2_dfrbp_1 \mem[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net317),
    .D(_0134_),
    .Q_N(_3055_),
    .Q(\mem[3][1] ));
 sg13g2_dfrbp_1 \mem[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net318),
    .D(_0135_),
    .Q_N(_3054_),
    .Q(\mem[3][2] ));
 sg13g2_dfrbp_1 \mem[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net319),
    .D(_0136_),
    .Q_N(_3053_),
    .Q(\mem[3][3] ));
 sg13g2_dfrbp_1 \mem[40][0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net320),
    .D(_0137_),
    .Q_N(_3052_),
    .Q(\mem[40][0] ));
 sg13g2_dfrbp_1 \mem[40][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net321),
    .D(_0138_),
    .Q_N(_3051_),
    .Q(\mem[40][1] ));
 sg13g2_dfrbp_1 \mem[40][2]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net322),
    .D(_0139_),
    .Q_N(_3050_),
    .Q(\mem[40][2] ));
 sg13g2_dfrbp_1 \mem[40][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net323),
    .D(_0140_),
    .Q_N(_3049_),
    .Q(\mem[40][3] ));
 sg13g2_dfrbp_1 \mem[41][0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net324),
    .D(_0141_),
    .Q_N(_3048_),
    .Q(\mem[41][0] ));
 sg13g2_dfrbp_1 \mem[41][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net325),
    .D(_0142_),
    .Q_N(_3047_),
    .Q(\mem[41][1] ));
 sg13g2_dfrbp_1 \mem[41][2]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net326),
    .D(_0143_),
    .Q_N(_3046_),
    .Q(\mem[41][2] ));
 sg13g2_dfrbp_1 \mem[41][3]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net327),
    .D(_0144_),
    .Q_N(_3045_),
    .Q(\mem[41][3] ));
 sg13g2_dfrbp_1 \mem[42][0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net328),
    .D(_0145_),
    .Q_N(_3044_),
    .Q(\mem[42][0] ));
 sg13g2_dfrbp_1 \mem[42][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net329),
    .D(_0146_),
    .Q_N(_3043_),
    .Q(\mem[42][1] ));
 sg13g2_dfrbp_1 \mem[42][2]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net330),
    .D(_0147_),
    .Q_N(_3042_),
    .Q(\mem[42][2] ));
 sg13g2_dfrbp_1 \mem[42][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net331),
    .D(_0148_),
    .Q_N(_3041_),
    .Q(\mem[42][3] ));
 sg13g2_dfrbp_1 \mem[43][0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net332),
    .D(_0149_),
    .Q_N(_3040_),
    .Q(\mem[43][0] ));
 sg13g2_dfrbp_1 \mem[43][1]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net333),
    .D(_0150_),
    .Q_N(_3039_),
    .Q(\mem[43][1] ));
 sg13g2_dfrbp_1 \mem[43][2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net334),
    .D(_0151_),
    .Q_N(_3038_),
    .Q(\mem[43][2] ));
 sg13g2_dfrbp_1 \mem[43][3]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net335),
    .D(_0152_),
    .Q_N(_3037_),
    .Q(\mem[43][3] ));
 sg13g2_dfrbp_1 \mem[44][0]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net336),
    .D(_0153_),
    .Q_N(_3036_),
    .Q(\mem[44][0] ));
 sg13g2_dfrbp_1 \mem[44][1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net337),
    .D(_0154_),
    .Q_N(_3035_),
    .Q(\mem[44][1] ));
 sg13g2_dfrbp_1 \mem[44][2]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net338),
    .D(_0155_),
    .Q_N(_3034_),
    .Q(\mem[44][2] ));
 sg13g2_dfrbp_1 \mem[44][3]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net339),
    .D(_0156_),
    .Q_N(_3033_),
    .Q(\mem[44][3] ));
 sg13g2_dfrbp_1 \mem[45][0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net340),
    .D(_0157_),
    .Q_N(_3032_),
    .Q(\mem[45][0] ));
 sg13g2_dfrbp_1 \mem[45][1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net341),
    .D(_0158_),
    .Q_N(_3031_),
    .Q(\mem[45][1] ));
 sg13g2_dfrbp_1 \mem[45][2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net342),
    .D(_0159_),
    .Q_N(_3030_),
    .Q(\mem[45][2] ));
 sg13g2_dfrbp_1 \mem[45][3]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net343),
    .D(_0160_),
    .Q_N(_3029_),
    .Q(\mem[45][3] ));
 sg13g2_dfrbp_1 \mem[46][0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net344),
    .D(_0161_),
    .Q_N(_3028_),
    .Q(\mem[46][0] ));
 sg13g2_dfrbp_1 \mem[46][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net345),
    .D(_0162_),
    .Q_N(_3027_),
    .Q(\mem[46][1] ));
 sg13g2_dfrbp_1 \mem[46][2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net346),
    .D(_0163_),
    .Q_N(_3026_),
    .Q(\mem[46][2] ));
 sg13g2_dfrbp_1 \mem[46][3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net347),
    .D(_0164_),
    .Q_N(_3025_),
    .Q(\mem[46][3] ));
 sg13g2_dfrbp_1 \mem[47][0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net348),
    .D(_0165_),
    .Q_N(_3024_),
    .Q(\mem[47][0] ));
 sg13g2_dfrbp_1 \mem[47][1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net349),
    .D(_0166_),
    .Q_N(_3023_),
    .Q(\mem[47][1] ));
 sg13g2_dfrbp_1 \mem[47][2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net350),
    .D(_0167_),
    .Q_N(_3022_),
    .Q(\mem[47][2] ));
 sg13g2_dfrbp_1 \mem[47][3]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net351),
    .D(_0168_),
    .Q_N(_3021_),
    .Q(\mem[47][3] ));
 sg13g2_dfrbp_1 \mem[48][0]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net352),
    .D(_0169_),
    .Q_N(_3020_),
    .Q(\mem[48][0] ));
 sg13g2_dfrbp_1 \mem[48][1]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net353),
    .D(_0170_),
    .Q_N(_3019_),
    .Q(\mem[48][1] ));
 sg13g2_dfrbp_1 \mem[48][2]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net354),
    .D(_0171_),
    .Q_N(_3018_),
    .Q(\mem[48][2] ));
 sg13g2_dfrbp_1 \mem[48][3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net355),
    .D(_0172_),
    .Q_N(_3017_),
    .Q(\mem[48][3] ));
 sg13g2_dfrbp_1 \mem[49][0]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net356),
    .D(_0173_),
    .Q_N(_3016_),
    .Q(\mem[49][0] ));
 sg13g2_dfrbp_1 \mem[49][1]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net357),
    .D(_0174_),
    .Q_N(_3015_),
    .Q(\mem[49][1] ));
 sg13g2_dfrbp_1 \mem[49][2]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net358),
    .D(_0175_),
    .Q_N(_3014_),
    .Q(\mem[49][2] ));
 sg13g2_dfrbp_1 \mem[49][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net359),
    .D(_0176_),
    .Q_N(_3013_),
    .Q(\mem[49][3] ));
 sg13g2_dfrbp_1 \mem[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net360),
    .D(_0177_),
    .Q_N(_3012_),
    .Q(\mem[4][0] ));
 sg13g2_dfrbp_1 \mem[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net361),
    .D(_0178_),
    .Q_N(_3011_),
    .Q(\mem[4][1] ));
 sg13g2_dfrbp_1 \mem[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net362),
    .D(_0179_),
    .Q_N(_3010_),
    .Q(\mem[4][2] ));
 sg13g2_dfrbp_1 \mem[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net363),
    .D(_0180_),
    .Q_N(_3009_),
    .Q(\mem[4][3] ));
 sg13g2_dfrbp_1 \mem[50][0]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net364),
    .D(_0181_),
    .Q_N(_3008_),
    .Q(\mem[50][0] ));
 sg13g2_dfrbp_1 \mem[50][1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net365),
    .D(_0182_),
    .Q_N(_3007_),
    .Q(\mem[50][1] ));
 sg13g2_dfrbp_1 \mem[50][2]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net366),
    .D(_0183_),
    .Q_N(_3006_),
    .Q(\mem[50][2] ));
 sg13g2_dfrbp_1 \mem[50][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net367),
    .D(_0184_),
    .Q_N(_3005_),
    .Q(\mem[50][3] ));
 sg13g2_dfrbp_1 \mem[51][0]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net368),
    .D(_0185_),
    .Q_N(_3004_),
    .Q(\mem[51][0] ));
 sg13g2_dfrbp_1 \mem[51][1]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net369),
    .D(_0186_),
    .Q_N(_3003_),
    .Q(\mem[51][1] ));
 sg13g2_dfrbp_1 \mem[51][2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net370),
    .D(_0187_),
    .Q_N(_3002_),
    .Q(\mem[51][2] ));
 sg13g2_dfrbp_1 \mem[51][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net371),
    .D(_0188_),
    .Q_N(_3001_),
    .Q(\mem[51][3] ));
 sg13g2_dfrbp_1 \mem[52][0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net372),
    .D(_0189_),
    .Q_N(_3000_),
    .Q(\mem[52][0] ));
 sg13g2_dfrbp_1 \mem[52][1]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net373),
    .D(_0190_),
    .Q_N(_2999_),
    .Q(\mem[52][1] ));
 sg13g2_dfrbp_1 \mem[52][2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net374),
    .D(_0191_),
    .Q_N(_2998_),
    .Q(\mem[52][2] ));
 sg13g2_dfrbp_1 \mem[52][3]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net375),
    .D(_0192_),
    .Q_N(_2997_),
    .Q(\mem[52][3] ));
 sg13g2_dfrbp_1 \mem[53][0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net376),
    .D(_0193_),
    .Q_N(_2996_),
    .Q(\mem[53][0] ));
 sg13g2_dfrbp_1 \mem[53][1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net377),
    .D(_0194_),
    .Q_N(_2995_),
    .Q(\mem[53][1] ));
 sg13g2_dfrbp_1 \mem[53][2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net378),
    .D(_0195_),
    .Q_N(_2994_),
    .Q(\mem[53][2] ));
 sg13g2_dfrbp_1 \mem[53][3]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net379),
    .D(_0196_),
    .Q_N(_2993_),
    .Q(\mem[53][3] ));
 sg13g2_dfrbp_1 \mem[54][0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net380),
    .D(_0197_),
    .Q_N(_2992_),
    .Q(\mem[54][0] ));
 sg13g2_dfrbp_1 \mem[54][1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net381),
    .D(_0198_),
    .Q_N(_2991_),
    .Q(\mem[54][1] ));
 sg13g2_dfrbp_1 \mem[54][2]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net382),
    .D(_0199_),
    .Q_N(_2990_),
    .Q(\mem[54][2] ));
 sg13g2_dfrbp_1 \mem[54][3]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net383),
    .D(_0200_),
    .Q_N(_2989_),
    .Q(\mem[54][3] ));
 sg13g2_dfrbp_1 \mem[55][0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net384),
    .D(_0201_),
    .Q_N(_2988_),
    .Q(\mem[55][0] ));
 sg13g2_dfrbp_1 \mem[55][1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net385),
    .D(_0202_),
    .Q_N(_2987_),
    .Q(\mem[55][1] ));
 sg13g2_dfrbp_1 \mem[55][2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net386),
    .D(_0203_),
    .Q_N(_2986_),
    .Q(\mem[55][2] ));
 sg13g2_dfrbp_1 \mem[55][3]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net387),
    .D(_0204_),
    .Q_N(_2985_),
    .Q(\mem[55][3] ));
 sg13g2_dfrbp_1 \mem[56][0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net388),
    .D(_0205_),
    .Q_N(_2984_),
    .Q(\mem[56][0] ));
 sg13g2_dfrbp_1 \mem[56][1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net389),
    .D(_0206_),
    .Q_N(_2983_),
    .Q(\mem[56][1] ));
 sg13g2_dfrbp_1 \mem[56][2]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net390),
    .D(_0207_),
    .Q_N(_2982_),
    .Q(\mem[56][2] ));
 sg13g2_dfrbp_1 \mem[56][3]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net391),
    .D(_0208_),
    .Q_N(_2981_),
    .Q(\mem[56][3] ));
 sg13g2_dfrbp_1 \mem[57][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net392),
    .D(_0209_),
    .Q_N(_2980_),
    .Q(\mem[57][0] ));
 sg13g2_dfrbp_1 \mem[57][1]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net393),
    .D(_0210_),
    .Q_N(_2979_),
    .Q(\mem[57][1] ));
 sg13g2_dfrbp_1 \mem[57][2]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net394),
    .D(_0211_),
    .Q_N(_2978_),
    .Q(\mem[57][2] ));
 sg13g2_dfrbp_1 \mem[57][3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net395),
    .D(_0212_),
    .Q_N(_2977_),
    .Q(\mem[57][3] ));
 sg13g2_dfrbp_1 \mem[58][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net396),
    .D(_0213_),
    .Q_N(_2976_),
    .Q(\mem[58][0] ));
 sg13g2_dfrbp_1 \mem[58][1]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net397),
    .D(_0214_),
    .Q_N(_2975_),
    .Q(\mem[58][1] ));
 sg13g2_dfrbp_1 \mem[58][2]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net398),
    .D(_0215_),
    .Q_N(_2974_),
    .Q(\mem[58][2] ));
 sg13g2_dfrbp_1 \mem[58][3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net399),
    .D(_0216_),
    .Q_N(_2973_),
    .Q(\mem[58][3] ));
 sg13g2_dfrbp_1 \mem[59][0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net400),
    .D(_0217_),
    .Q_N(_2972_),
    .Q(\mem[59][0] ));
 sg13g2_dfrbp_1 \mem[59][1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net401),
    .D(_0218_),
    .Q_N(_2971_),
    .Q(\mem[59][1] ));
 sg13g2_dfrbp_1 \mem[59][2]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net402),
    .D(_0219_),
    .Q_N(_2970_),
    .Q(\mem[59][2] ));
 sg13g2_dfrbp_1 \mem[59][3]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net403),
    .D(_0220_),
    .Q_N(_2969_),
    .Q(\mem[59][3] ));
 sg13g2_dfrbp_1 \mem[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net404),
    .D(_0221_),
    .Q_N(_2968_),
    .Q(\mem[5][0] ));
 sg13g2_dfrbp_1 \mem[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net405),
    .D(_0222_),
    .Q_N(_2967_),
    .Q(\mem[5][1] ));
 sg13g2_dfrbp_1 \mem[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net406),
    .D(_0223_),
    .Q_N(_2966_),
    .Q(\mem[5][2] ));
 sg13g2_dfrbp_1 \mem[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net407),
    .D(_0224_),
    .Q_N(_2965_),
    .Q(\mem[5][3] ));
 sg13g2_dfrbp_1 \mem[60][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net408),
    .D(_0225_),
    .Q_N(_2964_),
    .Q(\mem[60][0] ));
 sg13g2_dfrbp_1 \mem[60][1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net409),
    .D(_0226_),
    .Q_N(_2963_),
    .Q(\mem[60][1] ));
 sg13g2_dfrbp_1 \mem[60][2]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net410),
    .D(_0227_),
    .Q_N(_2962_),
    .Q(\mem[60][2] ));
 sg13g2_dfrbp_1 \mem[60][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net411),
    .D(_0228_),
    .Q_N(_2961_),
    .Q(\mem[60][3] ));
 sg13g2_dfrbp_1 \mem[61][0]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net412),
    .D(_0229_),
    .Q_N(_2960_),
    .Q(\mem[61][0] ));
 sg13g2_dfrbp_1 \mem[61][1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net413),
    .D(_0230_),
    .Q_N(_2959_),
    .Q(\mem[61][1] ));
 sg13g2_dfrbp_1 \mem[61][2]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net414),
    .D(_0231_),
    .Q_N(_2958_),
    .Q(\mem[61][2] ));
 sg13g2_dfrbp_1 \mem[61][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net415),
    .D(_0232_),
    .Q_N(_2957_),
    .Q(\mem[61][3] ));
 sg13g2_dfrbp_1 \mem[62][0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net416),
    .D(_0233_),
    .Q_N(_2956_),
    .Q(\mem[62][0] ));
 sg13g2_dfrbp_1 \mem[62][1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net417),
    .D(_0234_),
    .Q_N(_2955_),
    .Q(\mem[62][1] ));
 sg13g2_dfrbp_1 \mem[62][2]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net418),
    .D(_0235_),
    .Q_N(_2954_),
    .Q(\mem[62][2] ));
 sg13g2_dfrbp_1 \mem[62][3]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net419),
    .D(_0236_),
    .Q_N(_2953_),
    .Q(\mem[62][3] ));
 sg13g2_dfrbp_1 \mem[63][0]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net420),
    .D(_0237_),
    .Q_N(_2952_),
    .Q(\mem[63][0] ));
 sg13g2_dfrbp_1 \mem[63][1]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net421),
    .D(_0238_),
    .Q_N(_2951_),
    .Q(\mem[63][1] ));
 sg13g2_dfrbp_1 \mem[63][2]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net422),
    .D(_0239_),
    .Q_N(_2950_),
    .Q(\mem[63][2] ));
 sg13g2_dfrbp_1 \mem[63][3]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net423),
    .D(_0240_),
    .Q_N(_2949_),
    .Q(\mem[63][3] ));
 sg13g2_dfrbp_1 \mem[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net424),
    .D(_0241_),
    .Q_N(_2948_),
    .Q(\mem[6][0] ));
 sg13g2_dfrbp_1 \mem[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net425),
    .D(_0242_),
    .Q_N(_2947_),
    .Q(\mem[6][1] ));
 sg13g2_dfrbp_1 \mem[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net426),
    .D(_0243_),
    .Q_N(_2946_),
    .Q(\mem[6][2] ));
 sg13g2_dfrbp_1 \mem[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net427),
    .D(_0244_),
    .Q_N(_2945_),
    .Q(\mem[6][3] ));
 sg13g2_dfrbp_1 \mem[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net428),
    .D(_0245_),
    .Q_N(_2944_),
    .Q(\mem[7][0] ));
 sg13g2_dfrbp_1 \mem[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net429),
    .D(_0246_),
    .Q_N(_2943_),
    .Q(\mem[7][1] ));
 sg13g2_dfrbp_1 \mem[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net430),
    .D(_0247_),
    .Q_N(_2942_),
    .Q(\mem[7][2] ));
 sg13g2_dfrbp_1 \mem[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net431),
    .D(_0248_),
    .Q_N(_2941_),
    .Q(\mem[7][3] ));
 sg13g2_dfrbp_1 \mem[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net432),
    .D(_0249_),
    .Q_N(_2940_),
    .Q(\mem[8][0] ));
 sg13g2_dfrbp_1 \mem[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net433),
    .D(_0250_),
    .Q_N(_2939_),
    .Q(\mem[8][1] ));
 sg13g2_dfrbp_1 \mem[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net434),
    .D(_0251_),
    .Q_N(_2938_),
    .Q(\mem[8][2] ));
 sg13g2_dfrbp_1 \mem[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net435),
    .D(_0252_),
    .Q_N(_2937_),
    .Q(\mem[8][3] ));
 sg13g2_dfrbp_1 \mem[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net436),
    .D(_0253_),
    .Q_N(_2936_),
    .Q(\mem[9][0] ));
 sg13g2_dfrbp_1 \mem[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net437),
    .D(_0254_),
    .Q_N(_2935_),
    .Q(\mem[9][1] ));
 sg13g2_dfrbp_1 \mem[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net438),
    .D(_0255_),
    .Q_N(_2934_),
    .Q(\mem[9][2] ));
 sg13g2_dfrbp_1 \mem[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net439),
    .D(_0256_),
    .Q_N(_2933_),
    .Q(\mem[9][3] ));
 sg13g2_dfrbp_1 \prev_acc[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net440),
    .D(_0257_),
    .Q_N(_2932_),
    .Q(\prev_acc[0] ));
 sg13g2_dfrbp_1 \prev_acc[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net441),
    .D(_0258_),
    .Q_N(_2931_),
    .Q(\prev_acc[1] ));
 sg13g2_dfrbp_1 \prev_acc[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net442),
    .D(_0259_),
    .Q_N(_2930_),
    .Q(\prev_acc[2] ));
 sg13g2_dfrbp_1 \prev_acc[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net443),
    .D(_0260_),
    .Q_N(_2929_),
    .Q(\prev_acc[3] ));
 sg13g2_dfrbp_1 \prev_acc[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net444),
    .D(_0261_),
    .Q_N(_2928_),
    .Q(\prev_acc[4] ));
 sg13g2_dfrbp_1 \prev_acc[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net445),
    .D(_0262_),
    .Q_N(_2927_),
    .Q(\prev_acc[5] ));
 sg13g2_dfrbp_1 \prev_acc[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net446),
    .D(_0263_),
    .Q_N(_2926_),
    .Q(\prev_acc[6] ));
 sg13g2_dfrbp_1 \prev_acc[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net447),
    .D(_0264_),
    .Q_N(_2925_),
    .Q(\prev_acc[7] ));
 sg13g2_dfrbp_1 \products[0][0]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net448),
    .D(_0265_),
    .Q_N(_2924_),
    .Q(\products[0][0] ));
 sg13g2_dfrbp_1 \products[0][1]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net449),
    .D(_0266_),
    .Q_N(_2923_),
    .Q(\products[0][1] ));
 sg13g2_dfrbp_1 \products[0][2]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net450),
    .D(_0267_),
    .Q_N(_2922_),
    .Q(\products[0][2] ));
 sg13g2_dfrbp_1 \products[0][3]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net451),
    .D(_0268_),
    .Q_N(_2921_),
    .Q(\products[0][3] ));
 sg13g2_dfrbp_1 \products[0][4]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net452),
    .D(_0269_),
    .Q_N(_2920_),
    .Q(\products[0][4] ));
 sg13g2_dfrbp_1 \products[0][5]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net453),
    .D(_0270_),
    .Q_N(_2919_),
    .Q(\products[0][5] ));
 sg13g2_dfrbp_1 \products[0][6]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net454),
    .D(_0271_),
    .Q_N(_2918_),
    .Q(\products[0][6] ));
 sg13g2_dfrbp_1 \products[0][7]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net455),
    .D(_0272_),
    .Q_N(_2917_),
    .Q(\products[0][7] ));
 sg13g2_dfrbp_1 \products[10][0]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net456),
    .D(_0273_),
    .Q_N(_2916_),
    .Q(\products[10][0] ));
 sg13g2_dfrbp_1 \products[10][1]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net457),
    .D(_0274_),
    .Q_N(_2915_),
    .Q(\products[10][1] ));
 sg13g2_dfrbp_1 \products[10][2]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net458),
    .D(_0275_),
    .Q_N(_2914_),
    .Q(\products[10][2] ));
 sg13g2_dfrbp_1 \products[10][3]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net459),
    .D(_0276_),
    .Q_N(_2913_),
    .Q(\products[10][3] ));
 sg13g2_dfrbp_1 \products[10][4]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net460),
    .D(_0277_),
    .Q_N(_2912_),
    .Q(\products[10][4] ));
 sg13g2_dfrbp_1 \products[10][5]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net461),
    .D(_0278_),
    .Q_N(_2911_),
    .Q(\products[10][5] ));
 sg13g2_dfrbp_1 \products[10][6]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net462),
    .D(_0279_),
    .Q_N(_2910_),
    .Q(\products[10][6] ));
 sg13g2_dfrbp_1 \products[10][7]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net463),
    .D(_0280_),
    .Q_N(_2909_),
    .Q(\products[10][7] ));
 sg13g2_dfrbp_1 \products[11][0]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net464),
    .D(_0281_),
    .Q_N(_2908_),
    .Q(\products[11][0] ));
 sg13g2_dfrbp_1 \products[11][1]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net465),
    .D(_0282_),
    .Q_N(_2907_),
    .Q(\products[11][1] ));
 sg13g2_dfrbp_1 \products[11][2]$_SDFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net466),
    .D(_0283_),
    .Q_N(_2906_),
    .Q(\products[11][2] ));
 sg13g2_dfrbp_1 \products[11][3]$_SDFF_PN0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net467),
    .D(_0284_),
    .Q_N(_2905_),
    .Q(\products[11][3] ));
 sg13g2_dfrbp_1 \products[11][4]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net468),
    .D(_0285_),
    .Q_N(_2904_),
    .Q(\products[11][4] ));
 sg13g2_dfrbp_1 \products[11][5]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net469),
    .D(_0286_),
    .Q_N(_2903_),
    .Q(\products[11][5] ));
 sg13g2_dfrbp_1 \products[11][6]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net470),
    .D(_0287_),
    .Q_N(_2902_),
    .Q(\products[11][6] ));
 sg13g2_dfrbp_1 \products[11][7]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net471),
    .D(_0288_),
    .Q_N(_2901_),
    .Q(\products[11][7] ));
 sg13g2_dfrbp_1 \products[12][0]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net472),
    .D(_0289_),
    .Q_N(_2900_),
    .Q(\products[12][0] ));
 sg13g2_dfrbp_1 \products[12][1]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net473),
    .D(_0290_),
    .Q_N(_2899_),
    .Q(\products[12][1] ));
 sg13g2_dfrbp_1 \products[12][2]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net474),
    .D(_0291_),
    .Q_N(_2898_),
    .Q(\products[12][2] ));
 sg13g2_dfrbp_1 \products[12][3]$_SDFF_PN0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net475),
    .D(_0292_),
    .Q_N(_2897_),
    .Q(\products[12][3] ));
 sg13g2_dfrbp_1 \products[12][4]$_SDFF_PN0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net476),
    .D(_0293_),
    .Q_N(_2896_),
    .Q(\products[12][4] ));
 sg13g2_dfrbp_1 \products[12][5]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net477),
    .D(_0294_),
    .Q_N(_2895_),
    .Q(\products[12][5] ));
 sg13g2_dfrbp_1 \products[12][6]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net478),
    .D(_0295_),
    .Q_N(_2894_),
    .Q(\products[12][6] ));
 sg13g2_dfrbp_1 \products[12][7]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net479),
    .D(_0296_),
    .Q_N(_2893_),
    .Q(\products[12][7] ));
 sg13g2_dfrbp_1 \products[13][0]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net480),
    .D(_0297_),
    .Q_N(_2892_),
    .Q(\products[13][0] ));
 sg13g2_dfrbp_1 \products[13][1]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net481),
    .D(_0298_),
    .Q_N(_2891_),
    .Q(\products[13][1] ));
 sg13g2_dfrbp_1 \products[13][2]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net482),
    .D(_0299_),
    .Q_N(_2890_),
    .Q(\products[13][2] ));
 sg13g2_dfrbp_1 \products[13][3]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net483),
    .D(_0300_),
    .Q_N(_2889_),
    .Q(\products[13][3] ));
 sg13g2_dfrbp_1 \products[13][4]$_SDFF_PN0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net484),
    .D(_0301_),
    .Q_N(_2888_),
    .Q(\products[13][4] ));
 sg13g2_dfrbp_1 \products[13][5]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net485),
    .D(_0302_),
    .Q_N(_2887_),
    .Q(\products[13][5] ));
 sg13g2_dfrbp_1 \products[13][6]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net486),
    .D(_0303_),
    .Q_N(_2886_),
    .Q(\products[13][6] ));
 sg13g2_dfrbp_1 \products[13][7]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net487),
    .D(_0304_),
    .Q_N(_2885_),
    .Q(\products[13][7] ));
 sg13g2_dfrbp_1 \products[14][0]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net488),
    .D(_0305_),
    .Q_N(_2884_),
    .Q(\products[14][0] ));
 sg13g2_dfrbp_1 \products[14][1]$_SDFF_PN0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net489),
    .D(_0306_),
    .Q_N(_2883_),
    .Q(\products[14][1] ));
 sg13g2_dfrbp_1 \products[14][2]$_SDFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net490),
    .D(_0307_),
    .Q_N(_2882_),
    .Q(\products[14][2] ));
 sg13g2_dfrbp_1 \products[14][3]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net491),
    .D(_0308_),
    .Q_N(_2881_),
    .Q(\products[14][3] ));
 sg13g2_dfrbp_1 \products[14][4]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net492),
    .D(_0309_),
    .Q_N(_2880_),
    .Q(\products[14][4] ));
 sg13g2_dfrbp_1 \products[14][5]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net493),
    .D(_0310_),
    .Q_N(_2879_),
    .Q(\products[14][5] ));
 sg13g2_dfrbp_1 \products[14][6]$_SDFF_PN0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net494),
    .D(_0311_),
    .Q_N(_2878_),
    .Q(\products[14][6] ));
 sg13g2_dfrbp_1 \products[14][7]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net495),
    .D(_0312_),
    .Q_N(_2877_),
    .Q(\products[14][7] ));
 sg13g2_dfrbp_1 \products[15][0]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net496),
    .D(_0313_),
    .Q_N(_2876_),
    .Q(\products[15][0] ));
 sg13g2_dfrbp_1 \products[15][1]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net497),
    .D(_0314_),
    .Q_N(_2875_),
    .Q(\products[15][1] ));
 sg13g2_dfrbp_1 \products[15][2]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net498),
    .D(_0315_),
    .Q_N(_2874_),
    .Q(\products[15][2] ));
 sg13g2_dfrbp_1 \products[15][3]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net499),
    .D(_0316_),
    .Q_N(_2873_),
    .Q(\products[15][3] ));
 sg13g2_dfrbp_1 \products[15][4]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net500),
    .D(_0317_),
    .Q_N(_2872_),
    .Q(\products[15][4] ));
 sg13g2_dfrbp_1 \products[15][5]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net501),
    .D(_0318_),
    .Q_N(_2871_),
    .Q(\products[15][5] ));
 sg13g2_dfrbp_1 \products[15][6]$_SDFF_PN0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net502),
    .D(_0319_),
    .Q_N(_2870_),
    .Q(\products[15][6] ));
 sg13g2_dfrbp_1 \products[15][7]$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net503),
    .D(_0320_),
    .Q_N(_2869_),
    .Q(\products[15][7] ));
 sg13g2_dfrbp_1 \products[1][0]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net504),
    .D(_0321_),
    .Q_N(_2868_),
    .Q(\products[1][0] ));
 sg13g2_dfrbp_1 \products[1][1]$_SDFF_PN0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net505),
    .D(_0322_),
    .Q_N(_2867_),
    .Q(\products[1][1] ));
 sg13g2_dfrbp_1 \products[1][2]$_SDFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net506),
    .D(_0323_),
    .Q_N(_2866_),
    .Q(\products[1][2] ));
 sg13g2_dfrbp_1 \products[1][3]$_SDFF_PN0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net507),
    .D(_0324_),
    .Q_N(_2865_),
    .Q(\products[1][3] ));
 sg13g2_dfrbp_1 \products[1][4]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net508),
    .D(_0325_),
    .Q_N(_2864_),
    .Q(\products[1][4] ));
 sg13g2_dfrbp_1 \products[1][5]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net509),
    .D(_0326_),
    .Q_N(_2863_),
    .Q(\products[1][5] ));
 sg13g2_dfrbp_1 \products[1][6]$_SDFF_PN0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net510),
    .D(_0327_),
    .Q_N(_2862_),
    .Q(\products[1][6] ));
 sg13g2_dfrbp_1 \products[1][7]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net511),
    .D(_0328_),
    .Q_N(_2861_),
    .Q(\products[1][7] ));
 sg13g2_dfrbp_1 \products[2][0]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net512),
    .D(_0329_),
    .Q_N(_2860_),
    .Q(\products[2][0] ));
 sg13g2_dfrbp_1 \products[2][1]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net513),
    .D(_0330_),
    .Q_N(_2859_),
    .Q(\products[2][1] ));
 sg13g2_dfrbp_1 \products[2][2]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net514),
    .D(_0331_),
    .Q_N(_2858_),
    .Q(\products[2][2] ));
 sg13g2_dfrbp_1 \products[2][3]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net515),
    .D(_0332_),
    .Q_N(_2857_),
    .Q(\products[2][3] ));
 sg13g2_dfrbp_1 \products[2][4]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net516),
    .D(_0333_),
    .Q_N(_2856_),
    .Q(\products[2][4] ));
 sg13g2_dfrbp_1 \products[2][5]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net517),
    .D(_0334_),
    .Q_N(_2855_),
    .Q(\products[2][5] ));
 sg13g2_dfrbp_1 \products[2][6]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net518),
    .D(_0335_),
    .Q_N(_2854_),
    .Q(\products[2][6] ));
 sg13g2_dfrbp_1 \products[2][7]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net519),
    .D(_0336_),
    .Q_N(_2853_),
    .Q(\products[2][7] ));
 sg13g2_dfrbp_1 \products[3][0]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net520),
    .D(_0337_),
    .Q_N(_2852_),
    .Q(\products[3][0] ));
 sg13g2_dfrbp_1 \products[3][1]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net521),
    .D(_0338_),
    .Q_N(_2851_),
    .Q(\products[3][1] ));
 sg13g2_dfrbp_1 \products[3][2]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net522),
    .D(_0339_),
    .Q_N(_2850_),
    .Q(\products[3][2] ));
 sg13g2_dfrbp_1 \products[3][3]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net523),
    .D(_0340_),
    .Q_N(_2849_),
    .Q(\products[3][3] ));
 sg13g2_dfrbp_1 \products[3][4]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net524),
    .D(_0341_),
    .Q_N(_2848_),
    .Q(\products[3][4] ));
 sg13g2_dfrbp_1 \products[3][5]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net525),
    .D(_0342_),
    .Q_N(_2847_),
    .Q(\products[3][5] ));
 sg13g2_dfrbp_1 \products[3][6]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net526),
    .D(_0343_),
    .Q_N(_2846_),
    .Q(\products[3][6] ));
 sg13g2_dfrbp_1 \products[3][7]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net527),
    .D(_0344_),
    .Q_N(_2845_),
    .Q(\products[3][7] ));
 sg13g2_dfrbp_1 \products[4][0]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net528),
    .D(_0345_),
    .Q_N(_2844_),
    .Q(\products[4][0] ));
 sg13g2_dfrbp_1 \products[4][1]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net529),
    .D(_0346_),
    .Q_N(_2843_),
    .Q(\products[4][1] ));
 sg13g2_dfrbp_1 \products[4][2]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net530),
    .D(_0347_),
    .Q_N(_2842_),
    .Q(\products[4][2] ));
 sg13g2_dfrbp_1 \products[4][3]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net531),
    .D(_0348_),
    .Q_N(_2841_),
    .Q(\products[4][3] ));
 sg13g2_dfrbp_1 \products[4][4]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net532),
    .D(_0349_),
    .Q_N(_2840_),
    .Q(\products[4][4] ));
 sg13g2_dfrbp_1 \products[4][5]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net533),
    .D(_0350_),
    .Q_N(_2839_),
    .Q(\products[4][5] ));
 sg13g2_dfrbp_1 \products[4][6]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net534),
    .D(_0351_),
    .Q_N(_2838_),
    .Q(\products[4][6] ));
 sg13g2_dfrbp_1 \products[4][7]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net535),
    .D(_0352_),
    .Q_N(_2837_),
    .Q(\products[4][7] ));
 sg13g2_dfrbp_1 \products[5][0]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net536),
    .D(_0353_),
    .Q_N(_2836_),
    .Q(\products[5][0] ));
 sg13g2_dfrbp_1 \products[5][1]$_SDFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net537),
    .D(_0354_),
    .Q_N(_2835_),
    .Q(\products[5][1] ));
 sg13g2_dfrbp_1 \products[5][2]$_SDFF_PN0_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net538),
    .D(_0355_),
    .Q_N(_2834_),
    .Q(\products[5][2] ));
 sg13g2_dfrbp_1 \products[5][3]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net539),
    .D(_0356_),
    .Q_N(_2833_),
    .Q(\products[5][3] ));
 sg13g2_dfrbp_1 \products[5][4]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net540),
    .D(_0357_),
    .Q_N(_2832_),
    .Q(\products[5][4] ));
 sg13g2_dfrbp_1 \products[5][5]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net541),
    .D(_0358_),
    .Q_N(_2831_),
    .Q(\products[5][5] ));
 sg13g2_dfrbp_1 \products[5][6]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net542),
    .D(_0359_),
    .Q_N(_2830_),
    .Q(\products[5][6] ));
 sg13g2_dfrbp_1 \products[5][7]$_SDFF_PN0_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net543),
    .D(_0360_),
    .Q_N(_2829_),
    .Q(\products[5][7] ));
 sg13g2_dfrbp_1 \products[6][0]$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net544),
    .D(_0361_),
    .Q_N(_2828_),
    .Q(\products[6][0] ));
 sg13g2_dfrbp_1 \products[6][1]$_SDFF_PN0_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net545),
    .D(_0362_),
    .Q_N(_2827_),
    .Q(\products[6][1] ));
 sg13g2_dfrbp_1 \products[6][2]$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net546),
    .D(_0363_),
    .Q_N(_2826_),
    .Q(\products[6][2] ));
 sg13g2_dfrbp_1 \products[6][3]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net547),
    .D(_0364_),
    .Q_N(_2825_),
    .Q(\products[6][3] ));
 sg13g2_dfrbp_1 \products[6][4]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net548),
    .D(_0365_),
    .Q_N(_2824_),
    .Q(\products[6][4] ));
 sg13g2_dfrbp_1 \products[6][5]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net549),
    .D(_0366_),
    .Q_N(_2823_),
    .Q(\products[6][5] ));
 sg13g2_dfrbp_1 \products[6][6]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net550),
    .D(_0367_),
    .Q_N(_2822_),
    .Q(\products[6][6] ));
 sg13g2_dfrbp_1 \products[6][7]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net551),
    .D(_0368_),
    .Q_N(_2821_),
    .Q(\products[6][7] ));
 sg13g2_dfrbp_1 \products[7][0]$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net552),
    .D(_0369_),
    .Q_N(_2820_),
    .Q(\products[7][0] ));
 sg13g2_dfrbp_1 \products[7][1]$_SDFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net553),
    .D(_0370_),
    .Q_N(_2819_),
    .Q(\products[7][1] ));
 sg13g2_dfrbp_1 \products[7][2]$_SDFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net554),
    .D(_0371_),
    .Q_N(_2818_),
    .Q(\products[7][2] ));
 sg13g2_dfrbp_1 \products[7][3]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net555),
    .D(_0372_),
    .Q_N(_2817_),
    .Q(\products[7][3] ));
 sg13g2_dfrbp_1 \products[7][4]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net556),
    .D(_0373_),
    .Q_N(_2816_),
    .Q(\products[7][4] ));
 sg13g2_dfrbp_1 \products[7][5]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net557),
    .D(_0374_),
    .Q_N(_2815_),
    .Q(\products[7][5] ));
 sg13g2_dfrbp_1 \products[7][6]$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net558),
    .D(_0375_),
    .Q_N(_2814_),
    .Q(\products[7][6] ));
 sg13g2_dfrbp_1 \products[7][7]$_SDFF_PN0_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net559),
    .D(_0376_),
    .Q_N(_2813_),
    .Q(\products[7][7] ));
 sg13g2_dfrbp_1 \products[8][0]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net560),
    .D(_0377_),
    .Q_N(_2812_),
    .Q(\products[8][0] ));
 sg13g2_dfrbp_1 \products[8][1]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net561),
    .D(_0378_),
    .Q_N(_2811_),
    .Q(\products[8][1] ));
 sg13g2_dfrbp_1 \products[8][2]$_SDFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net562),
    .D(_0379_),
    .Q_N(_2810_),
    .Q(\products[8][2] ));
 sg13g2_dfrbp_1 \products[8][3]$_SDFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net563),
    .D(_0380_),
    .Q_N(_2809_),
    .Q(\products[8][3] ));
 sg13g2_dfrbp_1 \products[8][4]$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net564),
    .D(_0381_),
    .Q_N(_2808_),
    .Q(\products[8][4] ));
 sg13g2_dfrbp_1 \products[8][5]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net565),
    .D(_0382_),
    .Q_N(_2807_),
    .Q(\products[8][5] ));
 sg13g2_dfrbp_1 \products[8][6]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net566),
    .D(_0383_),
    .Q_N(_2806_),
    .Q(\products[8][6] ));
 sg13g2_dfrbp_1 \products[8][7]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net567),
    .D(_0384_),
    .Q_N(_2805_),
    .Q(\products[8][7] ));
 sg13g2_dfrbp_1 \products[9][0]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net568),
    .D(_0385_),
    .Q_N(_2804_),
    .Q(\products[9][0] ));
 sg13g2_dfrbp_1 \products[9][1]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net569),
    .D(_0386_),
    .Q_N(_2803_),
    .Q(\products[9][1] ));
 sg13g2_dfrbp_1 \products[9][2]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net570),
    .D(_0387_),
    .Q_N(_2802_),
    .Q(\products[9][2] ));
 sg13g2_dfrbp_1 \products[9][3]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net571),
    .D(_0388_),
    .Q_N(_2801_),
    .Q(\products[9][3] ));
 sg13g2_dfrbp_1 \products[9][4]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net572),
    .D(_0389_),
    .Q_N(_2800_),
    .Q(\products[9][4] ));
 sg13g2_dfrbp_1 \products[9][5]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net573),
    .D(_0390_),
    .Q_N(_2799_),
    .Q(\products[9][5] ));
 sg13g2_dfrbp_1 \products[9][6]$_SDFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net574),
    .D(_0391_),
    .Q_N(_2798_),
    .Q(\products[9][6] ));
 sg13g2_dfrbp_1 \products[9][7]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net575),
    .D(_0392_),
    .Q_N(_2797_),
    .Q(\products[9][7] ));
 sg13g2_dfrbp_1 \state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net576),
    .D(_0393_),
    .Q_N(_2796_),
    .Q(net15));
 sg13g2_dfrbp_1 \state[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net577),
    .D(_0394_),
    .Q_N(_2795_),
    .Q(net16));
 sg13g2_buf_1 input1 (.A(ui_in[6]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[7]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[0]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[2]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[3]),
    .X(net6));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[0]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[1]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[2]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[3]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout25 (.A(_1173_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1153_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0742_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0663_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0652_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0556_),
    .X(net30));
 sg13g2_buf_4 fanout31 (.X(net31),
    .A(_0555_));
 sg13g2_buf_2 fanout32 (.A(_1172_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1152_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0740_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0661_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0650_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0426_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0425_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1182_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1163_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1146_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0648_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0633_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_2721_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_2720_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1175_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1155_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0749_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0664_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0655_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_2633_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_2632_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1413_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2276_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1807_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1492_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1309_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2612_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1215_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1348_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1214_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0626_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0583_),
    .X(net63));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(_2537_));
 sg13g2_buf_4 fanout65 (.X(net65),
    .A(_2533_));
 sg13g2_buf_4 fanout66 (.X(net66),
    .A(_2527_));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(_2523_));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(_2522_));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(_2520_));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(_2518_));
 sg13g2_buf_4 fanout71 (.X(net71),
    .A(_2515_));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_2514_));
 sg13g2_buf_4 fanout73 (.X(net73),
    .A(_2512_));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(_2510_));
 sg13g2_buf_2 fanout75 (.A(_1322_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1321_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0727_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0725_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0582_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0580_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0558_),
    .X(net81));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_2536_));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_2529_));
 sg13g2_buf_8 fanout84 (.A(_2517_),
    .X(net84));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(_2511_));
 sg13g2_buf_2 fanout86 (.A(_1218_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1210_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1207_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1205_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1202_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1200_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_1197_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1195_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_1192_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_1186_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_1183_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1165_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1161_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_1140_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1137_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0774_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0773_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0770_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0764_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0763_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0762_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0759_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0757_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0756_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_0755_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0752_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0750_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0747_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0744_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0743_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0735_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0734_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0733_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0730_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0728_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0724_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0716_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_0710_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_0709_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0703_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_0702_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_0693_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_0692_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_0691_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0686_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_0685_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_0684_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_0681_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_0679_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_0678_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_0677_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_0674_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_0672_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_0671_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_0670_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_0667_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_0665_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0660_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_0654_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_0653_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_0651_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0646_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_0644_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_0643_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_0642_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_0639_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0637_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_0636_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_0635_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0631_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_0624_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_0622_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_0616_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_0614_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_0609_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_0607_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_0602_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_0600_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_0594_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_0592_),
    .X(net165));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(_0586_));
 sg13g2_buf_2 fanout167 (.A(_0585_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_0584_),
    .X(net168));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(_0574_));
 sg13g2_buf_2 fanout170 (.A(_0569_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_0563_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0559_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_0427_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_2722_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_2634_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_2642_),
    .X(net176));
 sg13g2_buf_4 fanout177 (.X(net177),
    .A(_2641_));
 sg13g2_tielo _5997__178 (.L_LO(net178));
 sg13g2_tielo _5998__179 (.L_LO(net179));
 sg13g2_tielo _5999__180 (.L_LO(net180));
 sg13g2_tielo _6000__181 (.L_LO(net181));
 sg13g2_tiehi _5996__183 (.L_HI(net183));
 sg13g2_tiehi \mem[0][0]$_DFFE_PP__184  (.L_HI(net184));
 sg13g2_tiehi \mem[0][1]$_DFFE_PP__185  (.L_HI(net185));
 sg13g2_tiehi \mem[0][2]$_DFFE_PP__186  (.L_HI(net186));
 sg13g2_tiehi \mem[0][3]$_DFFE_PP__187  (.L_HI(net187));
 sg13g2_tiehi \mem[10][0]$_DFFE_PP__188  (.L_HI(net188));
 sg13g2_tiehi \mem[10][1]$_DFFE_PP__189  (.L_HI(net189));
 sg13g2_tiehi \mem[10][2]$_DFFE_PP__190  (.L_HI(net190));
 sg13g2_tiehi \mem[10][3]$_DFFE_PP__191  (.L_HI(net191));
 sg13g2_tiehi \mem[11][0]$_DFFE_PP__192  (.L_HI(net192));
 sg13g2_tiehi \mem[11][1]$_DFFE_PP__193  (.L_HI(net193));
 sg13g2_tiehi \mem[11][2]$_DFFE_PP__194  (.L_HI(net194));
 sg13g2_tiehi \mem[11][3]$_DFFE_PP__195  (.L_HI(net195));
 sg13g2_tiehi \mem[12][0]$_DFFE_PP__196  (.L_HI(net196));
 sg13g2_tiehi \mem[12][1]$_DFFE_PP__197  (.L_HI(net197));
 sg13g2_tiehi \mem[12][2]$_DFFE_PP__198  (.L_HI(net198));
 sg13g2_tiehi \mem[12][3]$_DFFE_PP__199  (.L_HI(net199));
 sg13g2_tiehi \mem[13][0]$_DFFE_PP__200  (.L_HI(net200));
 sg13g2_tiehi \mem[13][1]$_DFFE_PP__201  (.L_HI(net201));
 sg13g2_tiehi \mem[13][2]$_DFFE_PP__202  (.L_HI(net202));
 sg13g2_tiehi \mem[13][3]$_DFFE_PP__203  (.L_HI(net203));
 sg13g2_tiehi \mem[14][0]$_DFFE_PP__204  (.L_HI(net204));
 sg13g2_tiehi \mem[14][1]$_DFFE_PP__205  (.L_HI(net205));
 sg13g2_tiehi \mem[14][2]$_DFFE_PP__206  (.L_HI(net206));
 sg13g2_tiehi \mem[14][3]$_DFFE_PP__207  (.L_HI(net207));
 sg13g2_tiehi \mem[15][0]$_DFFE_PP__208  (.L_HI(net208));
 sg13g2_tiehi \mem[15][1]$_DFFE_PP__209  (.L_HI(net209));
 sg13g2_tiehi \mem[15][2]$_DFFE_PP__210  (.L_HI(net210));
 sg13g2_tiehi \mem[15][3]$_DFFE_PP__211  (.L_HI(net211));
 sg13g2_tiehi \mem[16][0]$_DFFE_PP__212  (.L_HI(net212));
 sg13g2_tiehi \mem[16][1]$_DFFE_PP__213  (.L_HI(net213));
 sg13g2_tiehi \mem[16][2]$_DFFE_PP__214  (.L_HI(net214));
 sg13g2_tiehi \mem[16][3]$_DFFE_PP__215  (.L_HI(net215));
 sg13g2_tiehi \mem[17][0]$_DFFE_PP__216  (.L_HI(net216));
 sg13g2_tiehi \mem[17][1]$_DFFE_PP__217  (.L_HI(net217));
 sg13g2_tiehi \mem[17][2]$_DFFE_PP__218  (.L_HI(net218));
 sg13g2_tiehi \mem[17][3]$_DFFE_PP__219  (.L_HI(net219));
 sg13g2_tiehi \mem[18][0]$_DFFE_PP__220  (.L_HI(net220));
 sg13g2_tiehi \mem[18][1]$_DFFE_PP__221  (.L_HI(net221));
 sg13g2_tiehi \mem[18][2]$_DFFE_PP__222  (.L_HI(net222));
 sg13g2_tiehi \mem[18][3]$_DFFE_PP__223  (.L_HI(net223));
 sg13g2_tiehi \mem[19][0]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \mem[19][1]$_DFFE_PP__225  (.L_HI(net225));
 sg13g2_tiehi \mem[19][2]$_DFFE_PP__226  (.L_HI(net226));
 sg13g2_tiehi \mem[19][3]$_DFFE_PP__227  (.L_HI(net227));
 sg13g2_tiehi \mem[1][0]$_DFFE_PP__228  (.L_HI(net228));
 sg13g2_tiehi \mem[1][1]$_DFFE_PP__229  (.L_HI(net229));
 sg13g2_tiehi \mem[1][2]$_DFFE_PP__230  (.L_HI(net230));
 sg13g2_tiehi \mem[1][3]$_DFFE_PP__231  (.L_HI(net231));
 sg13g2_tiehi \mem[20][0]$_DFFE_PP__232  (.L_HI(net232));
 sg13g2_tiehi \mem[20][1]$_DFFE_PP__233  (.L_HI(net233));
 sg13g2_tiehi \mem[20][2]$_DFFE_PP__234  (.L_HI(net234));
 sg13g2_tiehi \mem[20][3]$_DFFE_PP__235  (.L_HI(net235));
 sg13g2_tiehi \mem[21][0]$_DFFE_PP__236  (.L_HI(net236));
 sg13g2_tiehi \mem[21][1]$_DFFE_PP__237  (.L_HI(net237));
 sg13g2_tiehi \mem[21][2]$_DFFE_PP__238  (.L_HI(net238));
 sg13g2_tiehi \mem[21][3]$_DFFE_PP__239  (.L_HI(net239));
 sg13g2_tiehi \mem[22][0]$_DFFE_PP__240  (.L_HI(net240));
 sg13g2_tiehi \mem[22][1]$_DFFE_PP__241  (.L_HI(net241));
 sg13g2_tiehi \mem[22][2]$_DFFE_PP__242  (.L_HI(net242));
 sg13g2_tiehi \mem[22][3]$_DFFE_PP__243  (.L_HI(net243));
 sg13g2_tiehi \mem[23][0]$_DFFE_PP__244  (.L_HI(net244));
 sg13g2_tiehi \mem[23][1]$_DFFE_PP__245  (.L_HI(net245));
 sg13g2_tiehi \mem[23][2]$_DFFE_PP__246  (.L_HI(net246));
 sg13g2_tiehi \mem[23][3]$_DFFE_PP__247  (.L_HI(net247));
 sg13g2_tiehi \mem[24][0]$_DFFE_PP__248  (.L_HI(net248));
 sg13g2_tiehi \mem[24][1]$_DFFE_PP__249  (.L_HI(net249));
 sg13g2_tiehi \mem[24][2]$_DFFE_PP__250  (.L_HI(net250));
 sg13g2_tiehi \mem[24][3]$_DFFE_PP__251  (.L_HI(net251));
 sg13g2_tiehi \mem[25][0]$_DFFE_PP__252  (.L_HI(net252));
 sg13g2_tiehi \mem[25][1]$_DFFE_PP__253  (.L_HI(net253));
 sg13g2_tiehi \mem[25][2]$_DFFE_PP__254  (.L_HI(net254));
 sg13g2_tiehi \mem[25][3]$_DFFE_PP__255  (.L_HI(net255));
 sg13g2_tiehi \mem[26][0]$_DFFE_PP__256  (.L_HI(net256));
 sg13g2_tiehi \mem[26][1]$_DFFE_PP__257  (.L_HI(net257));
 sg13g2_tiehi \mem[26][2]$_DFFE_PP__258  (.L_HI(net258));
 sg13g2_tiehi \mem[26][3]$_DFFE_PP__259  (.L_HI(net259));
 sg13g2_tiehi \mem[27][0]$_DFFE_PP__260  (.L_HI(net260));
 sg13g2_tiehi \mem[27][1]$_DFFE_PP__261  (.L_HI(net261));
 sg13g2_tiehi \mem[27][2]$_DFFE_PP__262  (.L_HI(net262));
 sg13g2_tiehi \mem[27][3]$_DFFE_PP__263  (.L_HI(net263));
 sg13g2_tiehi \mem[28][0]$_DFFE_PP__264  (.L_HI(net264));
 sg13g2_tiehi \mem[28][1]$_DFFE_PP__265  (.L_HI(net265));
 sg13g2_tiehi \mem[28][2]$_DFFE_PP__266  (.L_HI(net266));
 sg13g2_tiehi \mem[28][3]$_DFFE_PP__267  (.L_HI(net267));
 sg13g2_tiehi \mem[29][0]$_DFFE_PP__268  (.L_HI(net268));
 sg13g2_tiehi \mem[29][1]$_DFFE_PP__269  (.L_HI(net269));
 sg13g2_tiehi \mem[29][2]$_DFFE_PP__270  (.L_HI(net270));
 sg13g2_tiehi \mem[29][3]$_DFFE_PP__271  (.L_HI(net271));
 sg13g2_tiehi \mem[2][0]$_DFFE_PP__272  (.L_HI(net272));
 sg13g2_tiehi \mem[2][1]$_DFFE_PP__273  (.L_HI(net273));
 sg13g2_tiehi \mem[2][2]$_DFFE_PP__274  (.L_HI(net274));
 sg13g2_tiehi \mem[2][3]$_DFFE_PP__275  (.L_HI(net275));
 sg13g2_tiehi \mem[30][0]$_DFFE_PP__276  (.L_HI(net276));
 sg13g2_tiehi \mem[30][1]$_DFFE_PP__277  (.L_HI(net277));
 sg13g2_tiehi \mem[30][2]$_DFFE_PP__278  (.L_HI(net278));
 sg13g2_tiehi \mem[30][3]$_DFFE_PP__279  (.L_HI(net279));
 sg13g2_tiehi \mem[31][0]$_DFFE_PP__280  (.L_HI(net280));
 sg13g2_tiehi \mem[31][1]$_DFFE_PP__281  (.L_HI(net281));
 sg13g2_tiehi \mem[31][2]$_DFFE_PP__282  (.L_HI(net282));
 sg13g2_tiehi \mem[31][3]$_DFFE_PP__283  (.L_HI(net283));
 sg13g2_tiehi \mem[32][0]$_DFFE_PP__284  (.L_HI(net284));
 sg13g2_tiehi \mem[32][1]$_DFFE_PP__285  (.L_HI(net285));
 sg13g2_tiehi \mem[32][2]$_DFFE_PP__286  (.L_HI(net286));
 sg13g2_tiehi \mem[32][3]$_DFFE_PP__287  (.L_HI(net287));
 sg13g2_tiehi \mem[33][0]$_DFFE_PP__288  (.L_HI(net288));
 sg13g2_tiehi \mem[33][1]$_DFFE_PP__289  (.L_HI(net289));
 sg13g2_tiehi \mem[33][2]$_DFFE_PP__290  (.L_HI(net290));
 sg13g2_tiehi \mem[33][3]$_DFFE_PP__291  (.L_HI(net291));
 sg13g2_tiehi \mem[34][0]$_DFFE_PP__292  (.L_HI(net292));
 sg13g2_tiehi \mem[34][1]$_DFFE_PP__293  (.L_HI(net293));
 sg13g2_tiehi \mem[34][2]$_DFFE_PP__294  (.L_HI(net294));
 sg13g2_tiehi \mem[34][3]$_DFFE_PP__295  (.L_HI(net295));
 sg13g2_tiehi \mem[35][0]$_DFFE_PP__296  (.L_HI(net296));
 sg13g2_tiehi \mem[35][1]$_DFFE_PP__297  (.L_HI(net297));
 sg13g2_tiehi \mem[35][2]$_DFFE_PP__298  (.L_HI(net298));
 sg13g2_tiehi \mem[35][3]$_DFFE_PP__299  (.L_HI(net299));
 sg13g2_tiehi \mem[36][0]$_DFFE_PP__300  (.L_HI(net300));
 sg13g2_tiehi \mem[36][1]$_DFFE_PP__301  (.L_HI(net301));
 sg13g2_tiehi \mem[36][2]$_DFFE_PP__302  (.L_HI(net302));
 sg13g2_tiehi \mem[36][3]$_DFFE_PP__303  (.L_HI(net303));
 sg13g2_tiehi \mem[37][0]$_DFFE_PP__304  (.L_HI(net304));
 sg13g2_tiehi \mem[37][1]$_DFFE_PP__305  (.L_HI(net305));
 sg13g2_tiehi \mem[37][2]$_DFFE_PP__306  (.L_HI(net306));
 sg13g2_tiehi \mem[37][3]$_DFFE_PP__307  (.L_HI(net307));
 sg13g2_tiehi \mem[38][0]$_DFFE_PP__308  (.L_HI(net308));
 sg13g2_tiehi \mem[38][1]$_DFFE_PP__309  (.L_HI(net309));
 sg13g2_tiehi \mem[38][2]$_DFFE_PP__310  (.L_HI(net310));
 sg13g2_tiehi \mem[38][3]$_DFFE_PP__311  (.L_HI(net311));
 sg13g2_tiehi \mem[39][0]$_DFFE_PP__312  (.L_HI(net312));
 sg13g2_tiehi \mem[39][1]$_DFFE_PP__313  (.L_HI(net313));
 sg13g2_tiehi \mem[39][2]$_DFFE_PP__314  (.L_HI(net314));
 sg13g2_tiehi \mem[39][3]$_DFFE_PP__315  (.L_HI(net315));
 sg13g2_tiehi \mem[3][0]$_DFFE_PP__316  (.L_HI(net316));
 sg13g2_tiehi \mem[3][1]$_DFFE_PP__317  (.L_HI(net317));
 sg13g2_tiehi \mem[3][2]$_DFFE_PP__318  (.L_HI(net318));
 sg13g2_tiehi \mem[3][3]$_DFFE_PP__319  (.L_HI(net319));
 sg13g2_tiehi \mem[40][0]$_DFFE_PP__320  (.L_HI(net320));
 sg13g2_tiehi \mem[40][1]$_DFFE_PP__321  (.L_HI(net321));
 sg13g2_tiehi \mem[40][2]$_DFFE_PP__322  (.L_HI(net322));
 sg13g2_tiehi \mem[40][3]$_DFFE_PP__323  (.L_HI(net323));
 sg13g2_tiehi \mem[41][0]$_DFFE_PP__324  (.L_HI(net324));
 sg13g2_tiehi \mem[41][1]$_DFFE_PP__325  (.L_HI(net325));
 sg13g2_tiehi \mem[41][2]$_DFFE_PP__326  (.L_HI(net326));
 sg13g2_tiehi \mem[41][3]$_DFFE_PP__327  (.L_HI(net327));
 sg13g2_tiehi \mem[42][0]$_DFFE_PP__328  (.L_HI(net328));
 sg13g2_tiehi \mem[42][1]$_DFFE_PP__329  (.L_HI(net329));
 sg13g2_tiehi \mem[42][2]$_DFFE_PP__330  (.L_HI(net330));
 sg13g2_tiehi \mem[42][3]$_DFFE_PP__331  (.L_HI(net331));
 sg13g2_tiehi \mem[43][0]$_DFFE_PP__332  (.L_HI(net332));
 sg13g2_tiehi \mem[43][1]$_DFFE_PP__333  (.L_HI(net333));
 sg13g2_tiehi \mem[43][2]$_DFFE_PP__334  (.L_HI(net334));
 sg13g2_tiehi \mem[43][3]$_DFFE_PP__335  (.L_HI(net335));
 sg13g2_tiehi \mem[44][0]$_DFFE_PP__336  (.L_HI(net336));
 sg13g2_tiehi \mem[44][1]$_DFFE_PP__337  (.L_HI(net337));
 sg13g2_tiehi \mem[44][2]$_DFFE_PP__338  (.L_HI(net338));
 sg13g2_tiehi \mem[44][3]$_DFFE_PP__339  (.L_HI(net339));
 sg13g2_tiehi \mem[45][0]$_DFFE_PP__340  (.L_HI(net340));
 sg13g2_tiehi \mem[45][1]$_DFFE_PP__341  (.L_HI(net341));
 sg13g2_tiehi \mem[45][2]$_DFFE_PP__342  (.L_HI(net342));
 sg13g2_tiehi \mem[45][3]$_DFFE_PP__343  (.L_HI(net343));
 sg13g2_tiehi \mem[46][0]$_DFFE_PP__344  (.L_HI(net344));
 sg13g2_tiehi \mem[46][1]$_DFFE_PP__345  (.L_HI(net345));
 sg13g2_tiehi \mem[46][2]$_DFFE_PP__346  (.L_HI(net346));
 sg13g2_tiehi \mem[46][3]$_DFFE_PP__347  (.L_HI(net347));
 sg13g2_tiehi \mem[47][0]$_DFFE_PP__348  (.L_HI(net348));
 sg13g2_tiehi \mem[47][1]$_DFFE_PP__349  (.L_HI(net349));
 sg13g2_tiehi \mem[47][2]$_DFFE_PP__350  (.L_HI(net350));
 sg13g2_tiehi \mem[47][3]$_DFFE_PP__351  (.L_HI(net351));
 sg13g2_tiehi \mem[48][0]$_DFFE_PP__352  (.L_HI(net352));
 sg13g2_tiehi \mem[48][1]$_DFFE_PP__353  (.L_HI(net353));
 sg13g2_tiehi \mem[48][2]$_DFFE_PP__354  (.L_HI(net354));
 sg13g2_tiehi \mem[48][3]$_DFFE_PP__355  (.L_HI(net355));
 sg13g2_tiehi \mem[49][0]$_DFFE_PP__356  (.L_HI(net356));
 sg13g2_tiehi \mem[49][1]$_DFFE_PP__357  (.L_HI(net357));
 sg13g2_tiehi \mem[49][2]$_DFFE_PP__358  (.L_HI(net358));
 sg13g2_tiehi \mem[49][3]$_DFFE_PP__359  (.L_HI(net359));
 sg13g2_tiehi \mem[4][0]$_DFFE_PP__360  (.L_HI(net360));
 sg13g2_tiehi \mem[4][1]$_DFFE_PP__361  (.L_HI(net361));
 sg13g2_tiehi \mem[4][2]$_DFFE_PP__362  (.L_HI(net362));
 sg13g2_tiehi \mem[4][3]$_DFFE_PP__363  (.L_HI(net363));
 sg13g2_tiehi \mem[50][0]$_DFFE_PP__364  (.L_HI(net364));
 sg13g2_tiehi \mem[50][1]$_DFFE_PP__365  (.L_HI(net365));
 sg13g2_tiehi \mem[50][2]$_DFFE_PP__366  (.L_HI(net366));
 sg13g2_tiehi \mem[50][3]$_DFFE_PP__367  (.L_HI(net367));
 sg13g2_tiehi \mem[51][0]$_DFFE_PP__368  (.L_HI(net368));
 sg13g2_tiehi \mem[51][1]$_DFFE_PP__369  (.L_HI(net369));
 sg13g2_tiehi \mem[51][2]$_DFFE_PP__370  (.L_HI(net370));
 sg13g2_tiehi \mem[51][3]$_DFFE_PP__371  (.L_HI(net371));
 sg13g2_tiehi \mem[52][0]$_DFFE_PP__372  (.L_HI(net372));
 sg13g2_tiehi \mem[52][1]$_DFFE_PP__373  (.L_HI(net373));
 sg13g2_tiehi \mem[52][2]$_DFFE_PP__374  (.L_HI(net374));
 sg13g2_tiehi \mem[52][3]$_DFFE_PP__375  (.L_HI(net375));
 sg13g2_tiehi \mem[53][0]$_DFFE_PP__376  (.L_HI(net376));
 sg13g2_tiehi \mem[53][1]$_DFFE_PP__377  (.L_HI(net377));
 sg13g2_tiehi \mem[53][2]$_DFFE_PP__378  (.L_HI(net378));
 sg13g2_tiehi \mem[53][3]$_DFFE_PP__379  (.L_HI(net379));
 sg13g2_tiehi \mem[54][0]$_DFFE_PP__380  (.L_HI(net380));
 sg13g2_tiehi \mem[54][1]$_DFFE_PP__381  (.L_HI(net381));
 sg13g2_tiehi \mem[54][2]$_DFFE_PP__382  (.L_HI(net382));
 sg13g2_tiehi \mem[54][3]$_DFFE_PP__383  (.L_HI(net383));
 sg13g2_tiehi \mem[55][0]$_DFFE_PP__384  (.L_HI(net384));
 sg13g2_tiehi \mem[55][1]$_DFFE_PP__385  (.L_HI(net385));
 sg13g2_tiehi \mem[55][2]$_DFFE_PP__386  (.L_HI(net386));
 sg13g2_tiehi \mem[55][3]$_DFFE_PP__387  (.L_HI(net387));
 sg13g2_tiehi \mem[56][0]$_DFFE_PP__388  (.L_HI(net388));
 sg13g2_tiehi \mem[56][1]$_DFFE_PP__389  (.L_HI(net389));
 sg13g2_tiehi \mem[56][2]$_DFFE_PP__390  (.L_HI(net390));
 sg13g2_tiehi \mem[56][3]$_DFFE_PP__391  (.L_HI(net391));
 sg13g2_tiehi \mem[57][0]$_DFFE_PP__392  (.L_HI(net392));
 sg13g2_tiehi \mem[57][1]$_DFFE_PP__393  (.L_HI(net393));
 sg13g2_tiehi \mem[57][2]$_DFFE_PP__394  (.L_HI(net394));
 sg13g2_tiehi \mem[57][3]$_DFFE_PP__395  (.L_HI(net395));
 sg13g2_tiehi \mem[58][0]$_DFFE_PP__396  (.L_HI(net396));
 sg13g2_tiehi \mem[58][1]$_DFFE_PP__397  (.L_HI(net397));
 sg13g2_tiehi \mem[58][2]$_DFFE_PP__398  (.L_HI(net398));
 sg13g2_tiehi \mem[58][3]$_DFFE_PP__399  (.L_HI(net399));
 sg13g2_tiehi \mem[59][0]$_DFFE_PP__400  (.L_HI(net400));
 sg13g2_tiehi \mem[59][1]$_DFFE_PP__401  (.L_HI(net401));
 sg13g2_tiehi \mem[59][2]$_DFFE_PP__402  (.L_HI(net402));
 sg13g2_tiehi \mem[59][3]$_DFFE_PP__403  (.L_HI(net403));
 sg13g2_tiehi \mem[5][0]$_DFFE_PP__404  (.L_HI(net404));
 sg13g2_tiehi \mem[5][1]$_DFFE_PP__405  (.L_HI(net405));
 sg13g2_tiehi \mem[5][2]$_DFFE_PP__406  (.L_HI(net406));
 sg13g2_tiehi \mem[5][3]$_DFFE_PP__407  (.L_HI(net407));
 sg13g2_tiehi \mem[60][0]$_DFFE_PP__408  (.L_HI(net408));
 sg13g2_tiehi \mem[60][1]$_DFFE_PP__409  (.L_HI(net409));
 sg13g2_tiehi \mem[60][2]$_DFFE_PP__410  (.L_HI(net410));
 sg13g2_tiehi \mem[60][3]$_DFFE_PP__411  (.L_HI(net411));
 sg13g2_tiehi \mem[61][0]$_DFFE_PP__412  (.L_HI(net412));
 sg13g2_tiehi \mem[61][1]$_DFFE_PP__413  (.L_HI(net413));
 sg13g2_tiehi \mem[61][2]$_DFFE_PP__414  (.L_HI(net414));
 sg13g2_tiehi \mem[61][3]$_DFFE_PP__415  (.L_HI(net415));
 sg13g2_tiehi \mem[62][0]$_DFFE_PP__416  (.L_HI(net416));
 sg13g2_tiehi \mem[62][1]$_DFFE_PP__417  (.L_HI(net417));
 sg13g2_tiehi \mem[62][2]$_DFFE_PP__418  (.L_HI(net418));
 sg13g2_tiehi \mem[62][3]$_DFFE_PP__419  (.L_HI(net419));
 sg13g2_tiehi \mem[63][0]$_DFFE_PP__420  (.L_HI(net420));
 sg13g2_tiehi \mem[63][1]$_DFFE_PP__421  (.L_HI(net421));
 sg13g2_tiehi \mem[63][2]$_DFFE_PP__422  (.L_HI(net422));
 sg13g2_tiehi \mem[63][3]$_DFFE_PP__423  (.L_HI(net423));
 sg13g2_tiehi \mem[6][0]$_DFFE_PP__424  (.L_HI(net424));
 sg13g2_tiehi \mem[6][1]$_DFFE_PP__425  (.L_HI(net425));
 sg13g2_tiehi \mem[6][2]$_DFFE_PP__426  (.L_HI(net426));
 sg13g2_tiehi \mem[6][3]$_DFFE_PP__427  (.L_HI(net427));
 sg13g2_tiehi \mem[7][0]$_DFFE_PP__428  (.L_HI(net428));
 sg13g2_tiehi \mem[7][1]$_DFFE_PP__429  (.L_HI(net429));
 sg13g2_tiehi \mem[7][2]$_DFFE_PP__430  (.L_HI(net430));
 sg13g2_tiehi \mem[7][3]$_DFFE_PP__431  (.L_HI(net431));
 sg13g2_tiehi \mem[8][0]$_DFFE_PP__432  (.L_HI(net432));
 sg13g2_tiehi \mem[8][1]$_DFFE_PP__433  (.L_HI(net433));
 sg13g2_tiehi \mem[8][2]$_DFFE_PP__434  (.L_HI(net434));
 sg13g2_tiehi \mem[8][3]$_DFFE_PP__435  (.L_HI(net435));
 sg13g2_tiehi \mem[9][0]$_DFFE_PP__436  (.L_HI(net436));
 sg13g2_tiehi \mem[9][1]$_DFFE_PP__437  (.L_HI(net437));
 sg13g2_tiehi \mem[9][2]$_DFFE_PP__438  (.L_HI(net438));
 sg13g2_tiehi \mem[9][3]$_DFFE_PP__439  (.L_HI(net439));
 sg13g2_tiehi \prev_acc[0]$_SDFFE_PN0P__440  (.L_HI(net440));
 sg13g2_tiehi \prev_acc[1]$_SDFFE_PN0P__441  (.L_HI(net441));
 sg13g2_tiehi \prev_acc[2]$_SDFFE_PN0P__442  (.L_HI(net442));
 sg13g2_tiehi \prev_acc[3]$_SDFFE_PN0P__443  (.L_HI(net443));
 sg13g2_tiehi \prev_acc[4]$_SDFFE_PN0P__444  (.L_HI(net444));
 sg13g2_tiehi \prev_acc[5]$_SDFFE_PN0P__445  (.L_HI(net445));
 sg13g2_tiehi \prev_acc[6]$_SDFFE_PN0P__446  (.L_HI(net446));
 sg13g2_tiehi \prev_acc[7]$_SDFFE_PN0P__447  (.L_HI(net447));
 sg13g2_tiehi \products[0][0]$_SDFF_PN0__448  (.L_HI(net448));
 sg13g2_tiehi \products[0][1]$_SDFF_PN0__449  (.L_HI(net449));
 sg13g2_tiehi \products[0][2]$_SDFF_PN0__450  (.L_HI(net450));
 sg13g2_tiehi \products[0][3]$_SDFF_PN0__451  (.L_HI(net451));
 sg13g2_tiehi \products[0][4]$_SDFF_PN0__452  (.L_HI(net452));
 sg13g2_tiehi \products[0][5]$_SDFF_PN0__453  (.L_HI(net453));
 sg13g2_tiehi \products[0][6]$_SDFF_PN0__454  (.L_HI(net454));
 sg13g2_tiehi \products[0][7]$_SDFF_PN0__455  (.L_HI(net455));
 sg13g2_tiehi \products[10][0]$_SDFF_PN0__456  (.L_HI(net456));
 sg13g2_tiehi \products[10][1]$_SDFF_PN0__457  (.L_HI(net457));
 sg13g2_tiehi \products[10][2]$_SDFF_PN0__458  (.L_HI(net458));
 sg13g2_tiehi \products[10][3]$_SDFF_PN0__459  (.L_HI(net459));
 sg13g2_tiehi \products[10][4]$_SDFF_PN0__460  (.L_HI(net460));
 sg13g2_tiehi \products[10][5]$_SDFF_PN0__461  (.L_HI(net461));
 sg13g2_tiehi \products[10][6]$_SDFF_PN0__462  (.L_HI(net462));
 sg13g2_tiehi \products[10][7]$_SDFF_PN0__463  (.L_HI(net463));
 sg13g2_tiehi \products[11][0]$_SDFF_PN0__464  (.L_HI(net464));
 sg13g2_tiehi \products[11][1]$_SDFF_PN0__465  (.L_HI(net465));
 sg13g2_tiehi \products[11][2]$_SDFF_PN0__466  (.L_HI(net466));
 sg13g2_tiehi \products[11][3]$_SDFF_PN0__467  (.L_HI(net467));
 sg13g2_tiehi \products[11][4]$_SDFF_PN0__468  (.L_HI(net468));
 sg13g2_tiehi \products[11][5]$_SDFF_PN0__469  (.L_HI(net469));
 sg13g2_tiehi \products[11][6]$_SDFF_PN0__470  (.L_HI(net470));
 sg13g2_tiehi \products[11][7]$_SDFF_PN0__471  (.L_HI(net471));
 sg13g2_tiehi \products[12][0]$_SDFF_PN0__472  (.L_HI(net472));
 sg13g2_tiehi \products[12][1]$_SDFF_PN0__473  (.L_HI(net473));
 sg13g2_tiehi \products[12][2]$_SDFF_PN0__474  (.L_HI(net474));
 sg13g2_tiehi \products[12][3]$_SDFF_PN0__475  (.L_HI(net475));
 sg13g2_tiehi \products[12][4]$_SDFF_PN0__476  (.L_HI(net476));
 sg13g2_tiehi \products[12][5]$_SDFF_PN0__477  (.L_HI(net477));
 sg13g2_tiehi \products[12][6]$_SDFF_PN0__478  (.L_HI(net478));
 sg13g2_tiehi \products[12][7]$_SDFF_PN0__479  (.L_HI(net479));
 sg13g2_tiehi \products[13][0]$_SDFF_PN0__480  (.L_HI(net480));
 sg13g2_tiehi \products[13][1]$_SDFF_PN0__481  (.L_HI(net481));
 sg13g2_tiehi \products[13][2]$_SDFF_PN0__482  (.L_HI(net482));
 sg13g2_tiehi \products[13][3]$_SDFF_PN0__483  (.L_HI(net483));
 sg13g2_tiehi \products[13][4]$_SDFF_PN0__484  (.L_HI(net484));
 sg13g2_tiehi \products[13][5]$_SDFF_PN0__485  (.L_HI(net485));
 sg13g2_tiehi \products[13][6]$_SDFF_PN0__486  (.L_HI(net486));
 sg13g2_tiehi \products[13][7]$_SDFF_PN0__487  (.L_HI(net487));
 sg13g2_tiehi \products[14][0]$_SDFF_PN0__488  (.L_HI(net488));
 sg13g2_tiehi \products[14][1]$_SDFF_PN0__489  (.L_HI(net489));
 sg13g2_tiehi \products[14][2]$_SDFF_PN0__490  (.L_HI(net490));
 sg13g2_tiehi \products[14][3]$_SDFF_PN0__491  (.L_HI(net491));
 sg13g2_tiehi \products[14][4]$_SDFF_PN0__492  (.L_HI(net492));
 sg13g2_tiehi \products[14][5]$_SDFF_PN0__493  (.L_HI(net493));
 sg13g2_tiehi \products[14][6]$_SDFF_PN0__494  (.L_HI(net494));
 sg13g2_tiehi \products[14][7]$_SDFF_PN0__495  (.L_HI(net495));
 sg13g2_tiehi \products[15][0]$_SDFF_PN0__496  (.L_HI(net496));
 sg13g2_tiehi \products[15][1]$_SDFF_PN0__497  (.L_HI(net497));
 sg13g2_tiehi \products[15][2]$_SDFF_PN0__498  (.L_HI(net498));
 sg13g2_tiehi \products[15][3]$_SDFF_PN0__499  (.L_HI(net499));
 sg13g2_tiehi \products[15][4]$_SDFF_PN0__500  (.L_HI(net500));
 sg13g2_tiehi \products[15][5]$_SDFF_PN0__501  (.L_HI(net501));
 sg13g2_tiehi \products[15][6]$_SDFF_PN0__502  (.L_HI(net502));
 sg13g2_tiehi \products[15][7]$_SDFF_PN0__503  (.L_HI(net503));
 sg13g2_tiehi \products[1][0]$_SDFF_PN0__504  (.L_HI(net504));
 sg13g2_tiehi \products[1][1]$_SDFF_PN0__505  (.L_HI(net505));
 sg13g2_tiehi \products[1][2]$_SDFF_PN0__506  (.L_HI(net506));
 sg13g2_tiehi \products[1][3]$_SDFF_PN0__507  (.L_HI(net507));
 sg13g2_tiehi \products[1][4]$_SDFF_PN0__508  (.L_HI(net508));
 sg13g2_tiehi \products[1][5]$_SDFF_PN0__509  (.L_HI(net509));
 sg13g2_tiehi \products[1][6]$_SDFF_PN0__510  (.L_HI(net510));
 sg13g2_tiehi \products[1][7]$_SDFF_PN0__511  (.L_HI(net511));
 sg13g2_tiehi \products[2][0]$_SDFF_PN0__512  (.L_HI(net512));
 sg13g2_tiehi \products[2][1]$_SDFF_PN0__513  (.L_HI(net513));
 sg13g2_tiehi \products[2][2]$_SDFF_PN0__514  (.L_HI(net514));
 sg13g2_tiehi \products[2][3]$_SDFF_PN0__515  (.L_HI(net515));
 sg13g2_tiehi \products[2][4]$_SDFF_PN0__516  (.L_HI(net516));
 sg13g2_tiehi \products[2][5]$_SDFF_PN0__517  (.L_HI(net517));
 sg13g2_tiehi \products[2][6]$_SDFF_PN0__518  (.L_HI(net518));
 sg13g2_tiehi \products[2][7]$_SDFF_PN0__519  (.L_HI(net519));
 sg13g2_tiehi \products[3][0]$_SDFF_PN0__520  (.L_HI(net520));
 sg13g2_tiehi \products[3][1]$_SDFF_PN0__521  (.L_HI(net521));
 sg13g2_tiehi \products[3][2]$_SDFF_PN0__522  (.L_HI(net522));
 sg13g2_tiehi \products[3][3]$_SDFF_PN0__523  (.L_HI(net523));
 sg13g2_tiehi \products[3][4]$_SDFF_PN0__524  (.L_HI(net524));
 sg13g2_tiehi \products[3][5]$_SDFF_PN0__525  (.L_HI(net525));
 sg13g2_tiehi \products[3][6]$_SDFF_PN0__526  (.L_HI(net526));
 sg13g2_tiehi \products[3][7]$_SDFF_PN0__527  (.L_HI(net527));
 sg13g2_tiehi \products[4][0]$_SDFF_PN0__528  (.L_HI(net528));
 sg13g2_tiehi \products[4][1]$_SDFF_PN0__529  (.L_HI(net529));
 sg13g2_tiehi \products[4][2]$_SDFF_PN0__530  (.L_HI(net530));
 sg13g2_tiehi \products[4][3]$_SDFF_PN0__531  (.L_HI(net531));
 sg13g2_tiehi \products[4][4]$_SDFF_PN0__532  (.L_HI(net532));
 sg13g2_tiehi \products[4][5]$_SDFF_PN0__533  (.L_HI(net533));
 sg13g2_tiehi \products[4][6]$_SDFF_PN0__534  (.L_HI(net534));
 sg13g2_tiehi \products[4][7]$_SDFF_PN0__535  (.L_HI(net535));
 sg13g2_tiehi \products[5][0]$_SDFF_PN0__536  (.L_HI(net536));
 sg13g2_tiehi \products[5][1]$_SDFF_PN0__537  (.L_HI(net537));
 sg13g2_tiehi \products[5][2]$_SDFF_PN0__538  (.L_HI(net538));
 sg13g2_tiehi \products[5][3]$_SDFF_PN0__539  (.L_HI(net539));
 sg13g2_tiehi \products[5][4]$_SDFF_PN0__540  (.L_HI(net540));
 sg13g2_tiehi \products[5][5]$_SDFF_PN0__541  (.L_HI(net541));
 sg13g2_tiehi \products[5][6]$_SDFF_PN0__542  (.L_HI(net542));
 sg13g2_tiehi \products[5][7]$_SDFF_PN0__543  (.L_HI(net543));
 sg13g2_tiehi \products[6][0]$_SDFF_PN0__544  (.L_HI(net544));
 sg13g2_tiehi \products[6][1]$_SDFF_PN0__545  (.L_HI(net545));
 sg13g2_tiehi \products[6][2]$_SDFF_PN0__546  (.L_HI(net546));
 sg13g2_tiehi \products[6][3]$_SDFF_PN0__547  (.L_HI(net547));
 sg13g2_tiehi \products[6][4]$_SDFF_PN0__548  (.L_HI(net548));
 sg13g2_tiehi \products[6][5]$_SDFF_PN0__549  (.L_HI(net549));
 sg13g2_tiehi \products[6][6]$_SDFF_PN0__550  (.L_HI(net550));
 sg13g2_tiehi \products[6][7]$_SDFF_PN0__551  (.L_HI(net551));
 sg13g2_tiehi \products[7][0]$_SDFF_PN0__552  (.L_HI(net552));
 sg13g2_tiehi \products[7][1]$_SDFF_PN0__553  (.L_HI(net553));
 sg13g2_tiehi \products[7][2]$_SDFF_PN0__554  (.L_HI(net554));
 sg13g2_tiehi \products[7][3]$_SDFF_PN0__555  (.L_HI(net555));
 sg13g2_tiehi \products[7][4]$_SDFF_PN0__556  (.L_HI(net556));
 sg13g2_tiehi \products[7][5]$_SDFF_PN0__557  (.L_HI(net557));
 sg13g2_tiehi \products[7][6]$_SDFF_PN0__558  (.L_HI(net558));
 sg13g2_tiehi \products[7][7]$_SDFF_PN0__559  (.L_HI(net559));
 sg13g2_tiehi \products[8][0]$_SDFF_PN0__560  (.L_HI(net560));
 sg13g2_tiehi \products[8][1]$_SDFF_PN0__561  (.L_HI(net561));
 sg13g2_tiehi \products[8][2]$_SDFF_PN0__562  (.L_HI(net562));
 sg13g2_tiehi \products[8][3]$_SDFF_PN0__563  (.L_HI(net563));
 sg13g2_tiehi \products[8][4]$_SDFF_PN0__564  (.L_HI(net564));
 sg13g2_tiehi \products[8][5]$_SDFF_PN0__565  (.L_HI(net565));
 sg13g2_tiehi \products[8][6]$_SDFF_PN0__566  (.L_HI(net566));
 sg13g2_tiehi \products[8][7]$_SDFF_PN0__567  (.L_HI(net567));
 sg13g2_tiehi \products[9][0]$_SDFF_PN0__568  (.L_HI(net568));
 sg13g2_tiehi \products[9][1]$_SDFF_PN0__569  (.L_HI(net569));
 sg13g2_tiehi \products[9][2]$_SDFF_PN0__570  (.L_HI(net570));
 sg13g2_tiehi \products[9][3]$_SDFF_PN0__571  (.L_HI(net571));
 sg13g2_tiehi \products[9][4]$_SDFF_PN0__572  (.L_HI(net572));
 sg13g2_tiehi \products[9][5]$_SDFF_PN0__573  (.L_HI(net573));
 sg13g2_tiehi \products[9][6]$_SDFF_PN0__574  (.L_HI(net574));
 sg13g2_tiehi \products[9][7]$_SDFF_PN0__575  (.L_HI(net575));
 sg13g2_tiehi \state[0]$_SDFFE_PN0P__576  (.L_HI(net576));
 sg13g2_tiehi \state[1]$_SDFFE_PP0P__577  (.L_HI(net577));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_3_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_3_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_3_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_3_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_3_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_3_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_3_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_3_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_3_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_3_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_3_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_3_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_3_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_3_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_3_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_3_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_3_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_3_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_3_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_3_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_3_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_3_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_3_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_3_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_3_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_3_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_3_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_3_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_3_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_3_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_3_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_3_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_3_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_3_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_3_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_3_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_3_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_3_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_3_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_3_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_3_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_3_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_3_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_3_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_3_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_3_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_3_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_3_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_3_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_2 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_2 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_2 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_4 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_4 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_4_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_leaf_50_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_47_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_18_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_42_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_37_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_leaf_31_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0273_));
 sg13g2_antennanp ANTENNA_2 (.A(_0273_));
 sg13g2_antennanp ANTENNA_3 (.A(_0275_));
 sg13g2_antennanp ANTENNA_4 (.A(_0275_));
 sg13g2_antennanp ANTENNA_5 (.A(_0313_));
 sg13g2_antennanp ANTENNA_6 (.A(_0313_));
 sg13g2_antennanp ANTENNA_7 (.A(_0314_));
 sg13g2_antennanp ANTENNA_8 (.A(_0314_));
 sg13g2_antennanp ANTENNA_9 (.A(_0321_));
 sg13g2_antennanp ANTENNA_10 (.A(_0322_));
 sg13g2_antennanp ANTENNA_11 (.A(_0322_));
 sg13g2_antennanp ANTENNA_12 (.A(_0337_));
 sg13g2_antennanp ANTENNA_13 (.A(_0337_));
 sg13g2_antennanp ANTENNA_14 (.A(_0338_));
 sg13g2_antennanp ANTENNA_15 (.A(_0338_));
 sg13g2_antennanp ANTENNA_16 (.A(_0339_));
 sg13g2_antennanp ANTENNA_17 (.A(_0339_));
 sg13g2_antennanp ANTENNA_18 (.A(_0345_));
 sg13g2_antennanp ANTENNA_19 (.A(_0345_));
 sg13g2_antennanp ANTENNA_20 (.A(_0346_));
 sg13g2_antennanp ANTENNA_21 (.A(_0346_));
 sg13g2_antennanp ANTENNA_22 (.A(_0348_));
 sg13g2_antennanp ANTENNA_23 (.A(_0348_));
 sg13g2_antennanp ANTENNA_24 (.A(_0356_));
 sg13g2_antennanp ANTENNA_25 (.A(_0356_));
 sg13g2_antennanp ANTENNA_26 (.A(_0357_));
 sg13g2_antennanp ANTENNA_27 (.A(_0357_));
 sg13g2_antennanp ANTENNA_28 (.A(_0358_));
 sg13g2_antennanp ANTENNA_29 (.A(_0358_));
 sg13g2_antennanp ANTENNA_30 (.A(_0372_));
 sg13g2_antennanp ANTENNA_31 (.A(_0372_));
 sg13g2_antennanp ANTENNA_32 (.A(_0373_));
 sg13g2_antennanp ANTENNA_33 (.A(_0373_));
 sg13g2_antennanp ANTENNA_34 (.A(_0374_));
 sg13g2_antennanp ANTENNA_35 (.A(_0377_));
 sg13g2_antennanp ANTENNA_36 (.A(_0377_));
 sg13g2_antennanp ANTENNA_37 (.A(_0382_));
 sg13g2_antennanp ANTENNA_38 (.A(_0382_));
 sg13g2_antennanp ANTENNA_39 (.A(_0383_));
 sg13g2_antennanp ANTENNA_40 (.A(_0383_));
 sg13g2_antennanp ANTENNA_41 (.A(_0385_));
 sg13g2_antennanp ANTENNA_42 (.A(_0385_));
 sg13g2_antennanp ANTENNA_43 (.A(_0389_));
 sg13g2_antennanp ANTENNA_44 (.A(_0390_));
 sg13g2_antennanp ANTENNA_45 (.A(_0390_));
 sg13g2_antennanp ANTENNA_46 (.A(_0391_));
 sg13g2_antennanp ANTENNA_47 (.A(_0391_));
 sg13g2_antennanp ANTENNA_48 (.A(_0873_));
 sg13g2_antennanp ANTENNA_49 (.A(net45));
 sg13g2_antennanp ANTENNA_50 (.A(net45));
 sg13g2_antennanp ANTENNA_51 (.A(net45));
 sg13g2_antennanp ANTENNA_52 (.A(net45));
 sg13g2_antennanp ANTENNA_53 (.A(net45));
 sg13g2_antennanp ANTENNA_54 (.A(net45));
 sg13g2_antennanp ANTENNA_55 (.A(net45));
 sg13g2_antennanp ANTENNA_56 (.A(net45));
 sg13g2_antennanp ANTENNA_57 (.A(_0273_));
 sg13g2_antennanp ANTENNA_58 (.A(_0273_));
 sg13g2_antennanp ANTENNA_59 (.A(_0275_));
 sg13g2_antennanp ANTENNA_60 (.A(_0275_));
 sg13g2_antennanp ANTENNA_61 (.A(_0321_));
 sg13g2_antennanp ANTENNA_62 (.A(_0337_));
 sg13g2_antennanp ANTENNA_63 (.A(_0337_));
 sg13g2_antennanp ANTENNA_64 (.A(_0338_));
 sg13g2_antennanp ANTENNA_65 (.A(_0338_));
 sg13g2_antennanp ANTENNA_66 (.A(_0339_));
 sg13g2_antennanp ANTENNA_67 (.A(_0339_));
 sg13g2_antennanp ANTENNA_68 (.A(_0356_));
 sg13g2_antennanp ANTENNA_69 (.A(_0356_));
 sg13g2_antennanp ANTENNA_70 (.A(_0357_));
 sg13g2_antennanp ANTENNA_71 (.A(_0357_));
 sg13g2_antennanp ANTENNA_72 (.A(_0358_));
 sg13g2_antennanp ANTENNA_73 (.A(_0358_));
 sg13g2_antennanp ANTENNA_74 (.A(_0372_));
 sg13g2_antennanp ANTENNA_75 (.A(_0372_));
 sg13g2_antennanp ANTENNA_76 (.A(_0374_));
 sg13g2_antennanp ANTENNA_77 (.A(_0374_));
 sg13g2_antennanp ANTENNA_78 (.A(_0377_));
 sg13g2_antennanp ANTENNA_79 (.A(_0385_));
 sg13g2_antennanp ANTENNA_80 (.A(_0385_));
 sg13g2_antennanp ANTENNA_81 (.A(_0873_));
 sg13g2_antennanp ANTENNA_82 (.A(_0273_));
 sg13g2_antennanp ANTENNA_83 (.A(_0273_));
 sg13g2_antennanp ANTENNA_84 (.A(_0275_));
 sg13g2_antennanp ANTENNA_85 (.A(_0275_));
 sg13g2_antennanp ANTENNA_86 (.A(_0337_));
 sg13g2_antennanp ANTENNA_87 (.A(_0337_));
 sg13g2_antennanp ANTENNA_88 (.A(_0338_));
 sg13g2_antennanp ANTENNA_89 (.A(_0338_));
 sg13g2_antennanp ANTENNA_90 (.A(_0339_));
 sg13g2_antennanp ANTENNA_91 (.A(_0339_));
 sg13g2_antennanp ANTENNA_92 (.A(_0356_));
 sg13g2_antennanp ANTENNA_93 (.A(_0356_));
 sg13g2_antennanp ANTENNA_94 (.A(_0357_));
 sg13g2_antennanp ANTENNA_95 (.A(_0357_));
 sg13g2_antennanp ANTENNA_96 (.A(_0358_));
 sg13g2_antennanp ANTENNA_97 (.A(_0358_));
 sg13g2_antennanp ANTENNA_98 (.A(_0372_));
 sg13g2_antennanp ANTENNA_99 (.A(_0372_));
 sg13g2_antennanp ANTENNA_100 (.A(_0377_));
 sg13g2_antennanp ANTENNA_101 (.A(_0385_));
 sg13g2_antennanp ANTENNA_102 (.A(_0385_));
 sg13g2_antennanp ANTENNA_103 (.A(_0873_));
 sg13g2_antennanp ANTENNA_104 (.A(_0273_));
 sg13g2_antennanp ANTENNA_105 (.A(_0273_));
 sg13g2_antennanp ANTENNA_106 (.A(_0275_));
 sg13g2_antennanp ANTENNA_107 (.A(_0275_));
 sg13g2_antennanp ANTENNA_108 (.A(_0337_));
 sg13g2_antennanp ANTENNA_109 (.A(_0337_));
 sg13g2_antennanp ANTENNA_110 (.A(_0338_));
 sg13g2_antennanp ANTENNA_111 (.A(_0338_));
 sg13g2_antennanp ANTENNA_112 (.A(_0339_));
 sg13g2_antennanp ANTENNA_113 (.A(_0339_));
 sg13g2_antennanp ANTENNA_114 (.A(_0356_));
 sg13g2_antennanp ANTENNA_115 (.A(_0356_));
 sg13g2_antennanp ANTENNA_116 (.A(_0357_));
 sg13g2_antennanp ANTENNA_117 (.A(_0357_));
 sg13g2_antennanp ANTENNA_118 (.A(_0358_));
 sg13g2_antennanp ANTENNA_119 (.A(_0358_));
 sg13g2_antennanp ANTENNA_120 (.A(_0372_));
 sg13g2_antennanp ANTENNA_121 (.A(_0372_));
 sg13g2_antennanp ANTENNA_122 (.A(_0377_));
 sg13g2_antennanp ANTENNA_123 (.A(_0385_));
 sg13g2_antennanp ANTENNA_124 (.A(_0385_));
 sg13g2_antennanp ANTENNA_125 (.A(_0273_));
 sg13g2_antennanp ANTENNA_126 (.A(_0273_));
 sg13g2_antennanp ANTENNA_127 (.A(_0275_));
 sg13g2_antennanp ANTENNA_128 (.A(_0275_));
 sg13g2_antennanp ANTENNA_129 (.A(_0337_));
 sg13g2_antennanp ANTENNA_130 (.A(_0337_));
 sg13g2_antennanp ANTENNA_131 (.A(_0338_));
 sg13g2_antennanp ANTENNA_132 (.A(_0338_));
 sg13g2_antennanp ANTENNA_133 (.A(_0339_));
 sg13g2_antennanp ANTENNA_134 (.A(_0339_));
 sg13g2_antennanp ANTENNA_135 (.A(_0356_));
 sg13g2_antennanp ANTENNA_136 (.A(_0356_));
 sg13g2_antennanp ANTENNA_137 (.A(_0357_));
 sg13g2_antennanp ANTENNA_138 (.A(_0357_));
 sg13g2_antennanp ANTENNA_139 (.A(_0358_));
 sg13g2_antennanp ANTENNA_140 (.A(_0358_));
 sg13g2_antennanp ANTENNA_141 (.A(_0372_));
 sg13g2_antennanp ANTENNA_142 (.A(_0372_));
 sg13g2_antennanp ANTENNA_143 (.A(_0377_));
 sg13g2_antennanp ANTENNA_144 (.A(_0385_));
 sg13g2_antennanp ANTENNA_145 (.A(_0385_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_fill_2 FILLER_0_875 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_fill_2 FILLER_1_875 ();
 sg13g2_fill_1 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_fill_2 FILLER_2_875 ();
 sg13g2_fill_1 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_fill_2 FILLER_3_875 ();
 sg13g2_fill_1 FILLER_3_877 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_fill_2 FILLER_4_875 ();
 sg13g2_fill_1 FILLER_4_877 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_decap_8 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_5_868 ();
 sg13g2_fill_2 FILLER_5_875 ();
 sg13g2_fill_1 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_decap_8 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_6_868 ();
 sg13g2_fill_2 FILLER_6_875 ();
 sg13g2_fill_1 FILLER_6_877 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_fill_2 FILLER_7_875 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_fill_2 FILLER_8_875 ();
 sg13g2_fill_1 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_fill_2 FILLER_9_875 ();
 sg13g2_fill_1 FILLER_9_877 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_868 ();
 sg13g2_fill_2 FILLER_10_875 ();
 sg13g2_fill_1 FILLER_10_877 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_decap_8 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_11_868 ();
 sg13g2_fill_2 FILLER_11_875 ();
 sg13g2_fill_1 FILLER_11_877 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_decap_8 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_12_868 ();
 sg13g2_fill_2 FILLER_12_875 ();
 sg13g2_fill_1 FILLER_12_877 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_decap_8 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_13_868 ();
 sg13g2_fill_2 FILLER_13_875 ();
 sg13g2_fill_1 FILLER_13_877 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_decap_8 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_14_868 ();
 sg13g2_fill_2 FILLER_14_875 ();
 sg13g2_fill_1 FILLER_14_877 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_decap_8 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_15_868 ();
 sg13g2_fill_2 FILLER_15_875 ();
 sg13g2_fill_1 FILLER_15_877 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_decap_8 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_16_868 ();
 sg13g2_fill_2 FILLER_16_875 ();
 sg13g2_fill_1 FILLER_16_877 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_fill_2 FILLER_17_875 ();
 sg13g2_fill_1 FILLER_17_877 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_decap_8 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_18_868 ();
 sg13g2_fill_2 FILLER_18_875 ();
 sg13g2_fill_1 FILLER_18_877 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_decap_8 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_19_868 ();
 sg13g2_fill_2 FILLER_19_875 ();
 sg13g2_fill_1 FILLER_19_877 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_decap_8 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_20_868 ();
 sg13g2_fill_2 FILLER_20_875 ();
 sg13g2_fill_1 FILLER_20_877 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_21_868 ();
 sg13g2_fill_2 FILLER_21_875 ();
 sg13g2_fill_1 FILLER_21_877 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_decap_8 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_22_868 ();
 sg13g2_fill_2 FILLER_22_875 ();
 sg13g2_fill_1 FILLER_22_877 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_decap_8 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_fill_2 FILLER_23_875 ();
 sg13g2_fill_1 FILLER_23_877 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_decap_8 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_24_868 ();
 sg13g2_fill_2 FILLER_24_875 ();
 sg13g2_fill_1 FILLER_24_877 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_decap_8 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_581 ();
 sg13g2_decap_8 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_decap_8 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_fill_2 FILLER_25_875 ();
 sg13g2_fill_1 FILLER_25_877 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_8 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_decap_8 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_26_868 ();
 sg13g2_fill_2 FILLER_26_875 ();
 sg13g2_fill_1 FILLER_26_877 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_fill_2 FILLER_27_875 ();
 sg13g2_fill_1 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_decap_8 FILLER_28_427 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_decap_8 FILLER_28_441 ();
 sg13g2_decap_8 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_462 ();
 sg13g2_decap_8 FILLER_28_469 ();
 sg13g2_decap_8 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_483 ();
 sg13g2_decap_8 FILLER_28_490 ();
 sg13g2_decap_8 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_504 ();
 sg13g2_decap_8 FILLER_28_511 ();
 sg13g2_decap_8 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_decap_8 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_546 ();
 sg13g2_decap_8 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_560 ();
 sg13g2_decap_8 FILLER_28_567 ();
 sg13g2_decap_8 FILLER_28_574 ();
 sg13g2_decap_8 FILLER_28_581 ();
 sg13g2_decap_8 FILLER_28_588 ();
 sg13g2_decap_8 FILLER_28_595 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_decap_8 FILLER_28_609 ();
 sg13g2_decap_8 FILLER_28_616 ();
 sg13g2_decap_8 FILLER_28_623 ();
 sg13g2_decap_8 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_decap_8 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_decap_8 FILLER_28_679 ();
 sg13g2_decap_8 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_693 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_decap_8 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_28_868 ();
 sg13g2_fill_2 FILLER_28_875 ();
 sg13g2_fill_1 FILLER_28_877 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_490 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_decap_8 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_525 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_8 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_8 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_decap_8 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_29_868 ();
 sg13g2_fill_2 FILLER_29_875 ();
 sg13g2_fill_1 FILLER_29_877 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_fill_2 FILLER_30_322 ();
 sg13g2_fill_2 FILLER_30_329 ();
 sg13g2_fill_1 FILLER_30_331 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_8 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_349 ();
 sg13g2_fill_2 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_fill_2 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_8 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_30_410 ();
 sg13g2_decap_8 FILLER_30_417 ();
 sg13g2_decap_8 FILLER_30_424 ();
 sg13g2_decap_8 FILLER_30_431 ();
 sg13g2_decap_8 FILLER_30_438 ();
 sg13g2_decap_8 FILLER_30_445 ();
 sg13g2_decap_8 FILLER_30_452 ();
 sg13g2_decap_8 FILLER_30_459 ();
 sg13g2_decap_8 FILLER_30_466 ();
 sg13g2_decap_8 FILLER_30_473 ();
 sg13g2_decap_8 FILLER_30_480 ();
 sg13g2_decap_8 FILLER_30_487 ();
 sg13g2_decap_8 FILLER_30_494 ();
 sg13g2_decap_8 FILLER_30_501 ();
 sg13g2_decap_8 FILLER_30_508 ();
 sg13g2_decap_8 FILLER_30_515 ();
 sg13g2_decap_8 FILLER_30_522 ();
 sg13g2_decap_8 FILLER_30_529 ();
 sg13g2_decap_8 FILLER_30_536 ();
 sg13g2_decap_8 FILLER_30_543 ();
 sg13g2_decap_8 FILLER_30_550 ();
 sg13g2_decap_8 FILLER_30_557 ();
 sg13g2_decap_8 FILLER_30_564 ();
 sg13g2_decap_8 FILLER_30_571 ();
 sg13g2_decap_8 FILLER_30_578 ();
 sg13g2_decap_8 FILLER_30_585 ();
 sg13g2_decap_8 FILLER_30_592 ();
 sg13g2_decap_8 FILLER_30_599 ();
 sg13g2_decap_8 FILLER_30_606 ();
 sg13g2_decap_8 FILLER_30_613 ();
 sg13g2_decap_8 FILLER_30_620 ();
 sg13g2_decap_8 FILLER_30_627 ();
 sg13g2_decap_8 FILLER_30_634 ();
 sg13g2_decap_8 FILLER_30_641 ();
 sg13g2_decap_8 FILLER_30_648 ();
 sg13g2_decap_8 FILLER_30_655 ();
 sg13g2_decap_8 FILLER_30_662 ();
 sg13g2_decap_8 FILLER_30_669 ();
 sg13g2_decap_8 FILLER_30_676 ();
 sg13g2_decap_8 FILLER_30_683 ();
 sg13g2_decap_8 FILLER_30_690 ();
 sg13g2_decap_8 FILLER_30_697 ();
 sg13g2_decap_8 FILLER_30_704 ();
 sg13g2_decap_8 FILLER_30_711 ();
 sg13g2_decap_8 FILLER_30_718 ();
 sg13g2_decap_8 FILLER_30_725 ();
 sg13g2_decap_8 FILLER_30_732 ();
 sg13g2_decap_8 FILLER_30_739 ();
 sg13g2_decap_8 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_decap_8 FILLER_30_767 ();
 sg13g2_decap_8 FILLER_30_774 ();
 sg13g2_decap_8 FILLER_30_781 ();
 sg13g2_decap_8 FILLER_30_788 ();
 sg13g2_decap_8 FILLER_30_795 ();
 sg13g2_decap_8 FILLER_30_802 ();
 sg13g2_decap_8 FILLER_30_809 ();
 sg13g2_decap_8 FILLER_30_816 ();
 sg13g2_decap_8 FILLER_30_823 ();
 sg13g2_decap_8 FILLER_30_830 ();
 sg13g2_decap_8 FILLER_30_837 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_8 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_30_865 ();
 sg13g2_decap_4 FILLER_30_872 ();
 sg13g2_fill_2 FILLER_30_876 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_fill_2 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_361 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_413 ();
 sg13g2_decap_4 FILLER_31_418 ();
 sg13g2_fill_2 FILLER_31_422 ();
 sg13g2_decap_8 FILLER_31_450 ();
 sg13g2_decap_8 FILLER_31_457 ();
 sg13g2_decap_4 FILLER_31_464 ();
 sg13g2_fill_1 FILLER_31_468 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_4 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_505 ();
 sg13g2_decap_8 FILLER_31_512 ();
 sg13g2_decap_8 FILLER_31_519 ();
 sg13g2_fill_1 FILLER_31_526 ();
 sg13g2_decap_8 FILLER_31_557 ();
 sg13g2_decap_8 FILLER_31_564 ();
 sg13g2_decap_8 FILLER_31_571 ();
 sg13g2_decap_8 FILLER_31_578 ();
 sg13g2_decap_8 FILLER_31_585 ();
 sg13g2_decap_8 FILLER_31_592 ();
 sg13g2_decap_8 FILLER_31_599 ();
 sg13g2_decap_8 FILLER_31_606 ();
 sg13g2_decap_8 FILLER_31_613 ();
 sg13g2_decap_8 FILLER_31_620 ();
 sg13g2_decap_8 FILLER_31_627 ();
 sg13g2_decap_8 FILLER_31_634 ();
 sg13g2_decap_8 FILLER_31_641 ();
 sg13g2_decap_8 FILLER_31_648 ();
 sg13g2_decap_8 FILLER_31_655 ();
 sg13g2_decap_8 FILLER_31_662 ();
 sg13g2_decap_8 FILLER_31_669 ();
 sg13g2_decap_8 FILLER_31_676 ();
 sg13g2_decap_8 FILLER_31_683 ();
 sg13g2_decap_8 FILLER_31_690 ();
 sg13g2_decap_8 FILLER_31_697 ();
 sg13g2_decap_8 FILLER_31_704 ();
 sg13g2_decap_8 FILLER_31_711 ();
 sg13g2_decap_8 FILLER_31_718 ();
 sg13g2_decap_8 FILLER_31_725 ();
 sg13g2_decap_8 FILLER_31_732 ();
 sg13g2_decap_8 FILLER_31_739 ();
 sg13g2_decap_8 FILLER_31_746 ();
 sg13g2_decap_8 FILLER_31_753 ();
 sg13g2_decap_8 FILLER_31_760 ();
 sg13g2_decap_8 FILLER_31_767 ();
 sg13g2_decap_8 FILLER_31_774 ();
 sg13g2_decap_8 FILLER_31_781 ();
 sg13g2_decap_8 FILLER_31_788 ();
 sg13g2_decap_8 FILLER_31_795 ();
 sg13g2_decap_8 FILLER_31_802 ();
 sg13g2_decap_8 FILLER_31_809 ();
 sg13g2_decap_8 FILLER_31_816 ();
 sg13g2_decap_8 FILLER_31_823 ();
 sg13g2_decap_8 FILLER_31_830 ();
 sg13g2_decap_8 FILLER_31_837 ();
 sg13g2_decap_8 FILLER_31_844 ();
 sg13g2_decap_8 FILLER_31_851 ();
 sg13g2_decap_8 FILLER_31_858 ();
 sg13g2_decap_8 FILLER_31_865 ();
 sg13g2_decap_4 FILLER_31_872 ();
 sg13g2_fill_2 FILLER_31_876 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_4 FILLER_32_287 ();
 sg13g2_fill_2 FILLER_32_291 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_decap_4 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_346 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_fill_2 FILLER_32_401 ();
 sg13g2_decap_4 FILLER_32_416 ();
 sg13g2_fill_1 FILLER_32_420 ();
 sg13g2_fill_1 FILLER_32_455 ();
 sg13g2_fill_1 FILLER_32_464 ();
 sg13g2_fill_1 FILLER_32_491 ();
 sg13g2_fill_2 FILLER_32_518 ();
 sg13g2_decap_8 FILLER_32_528 ();
 sg13g2_fill_2 FILLER_32_535 ();
 sg13g2_decap_4 FILLER_32_568 ();
 sg13g2_fill_1 FILLER_32_572 ();
 sg13g2_decap_8 FILLER_32_581 ();
 sg13g2_decap_8 FILLER_32_588 ();
 sg13g2_decap_4 FILLER_32_595 ();
 sg13g2_decap_8 FILLER_32_625 ();
 sg13g2_decap_8 FILLER_32_632 ();
 sg13g2_decap_4 FILLER_32_639 ();
 sg13g2_fill_1 FILLER_32_643 ();
 sg13g2_decap_8 FILLER_32_647 ();
 sg13g2_decap_8 FILLER_32_654 ();
 sg13g2_decap_8 FILLER_32_661 ();
 sg13g2_decap_8 FILLER_32_668 ();
 sg13g2_decap_8 FILLER_32_675 ();
 sg13g2_decap_8 FILLER_32_682 ();
 sg13g2_decap_8 FILLER_32_689 ();
 sg13g2_decap_8 FILLER_32_696 ();
 sg13g2_decap_8 FILLER_32_703 ();
 sg13g2_decap_8 FILLER_32_710 ();
 sg13g2_decap_8 FILLER_32_717 ();
 sg13g2_decap_8 FILLER_32_724 ();
 sg13g2_decap_8 FILLER_32_731 ();
 sg13g2_decap_8 FILLER_32_738 ();
 sg13g2_decap_8 FILLER_32_745 ();
 sg13g2_decap_8 FILLER_32_752 ();
 sg13g2_decap_8 FILLER_32_759 ();
 sg13g2_decap_8 FILLER_32_766 ();
 sg13g2_decap_8 FILLER_32_773 ();
 sg13g2_decap_8 FILLER_32_780 ();
 sg13g2_decap_8 FILLER_32_787 ();
 sg13g2_decap_8 FILLER_32_794 ();
 sg13g2_decap_8 FILLER_32_801 ();
 sg13g2_decap_8 FILLER_32_808 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_decap_8 FILLER_32_822 ();
 sg13g2_decap_8 FILLER_32_829 ();
 sg13g2_decap_8 FILLER_32_836 ();
 sg13g2_decap_8 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_850 ();
 sg13g2_decap_8 FILLER_32_857 ();
 sg13g2_decap_8 FILLER_32_864 ();
 sg13g2_decap_8 FILLER_32_871 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_fill_1 FILLER_33_383 ();
 sg13g2_fill_2 FILLER_33_392 ();
 sg13g2_fill_1 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_33_398 ();
 sg13g2_fill_1 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_409 ();
 sg13g2_fill_2 FILLER_33_432 ();
 sg13g2_fill_1 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_439 ();
 sg13g2_decap_4 FILLER_33_446 ();
 sg13g2_fill_1 FILLER_33_458 ();
 sg13g2_fill_2 FILLER_33_501 ();
 sg13g2_fill_1 FILLER_33_503 ();
 sg13g2_fill_2 FILLER_33_508 ();
 sg13g2_fill_2 FILLER_33_522 ();
 sg13g2_fill_1 FILLER_33_524 ();
 sg13g2_fill_2 FILLER_33_533 ();
 sg13g2_fill_1 FILLER_33_535 ();
 sg13g2_fill_2 FILLER_33_569 ();
 sg13g2_fill_1 FILLER_33_571 ();
 sg13g2_fill_1 FILLER_33_580 ();
 sg13g2_fill_1 FILLER_33_590 ();
 sg13g2_fill_2 FILLER_33_601 ();
 sg13g2_fill_1 FILLER_33_606 ();
 sg13g2_decap_8 FILLER_33_611 ();
 sg13g2_decap_8 FILLER_33_618 ();
 sg13g2_decap_8 FILLER_33_625 ();
 sg13g2_decap_4 FILLER_33_632 ();
 sg13g2_fill_1 FILLER_33_636 ();
 sg13g2_decap_8 FILLER_33_670 ();
 sg13g2_decap_8 FILLER_33_677 ();
 sg13g2_decap_8 FILLER_33_684 ();
 sg13g2_decap_8 FILLER_33_691 ();
 sg13g2_decap_8 FILLER_33_698 ();
 sg13g2_decap_8 FILLER_33_705 ();
 sg13g2_decap_8 FILLER_33_712 ();
 sg13g2_decap_8 FILLER_33_719 ();
 sg13g2_decap_8 FILLER_33_726 ();
 sg13g2_decap_8 FILLER_33_733 ();
 sg13g2_decap_8 FILLER_33_740 ();
 sg13g2_decap_8 FILLER_33_747 ();
 sg13g2_decap_8 FILLER_33_754 ();
 sg13g2_decap_8 FILLER_33_761 ();
 sg13g2_decap_8 FILLER_33_768 ();
 sg13g2_decap_8 FILLER_33_775 ();
 sg13g2_decap_8 FILLER_33_782 ();
 sg13g2_decap_8 FILLER_33_789 ();
 sg13g2_decap_8 FILLER_33_796 ();
 sg13g2_decap_8 FILLER_33_803 ();
 sg13g2_decap_8 FILLER_33_810 ();
 sg13g2_decap_8 FILLER_33_817 ();
 sg13g2_decap_8 FILLER_33_824 ();
 sg13g2_decap_8 FILLER_33_831 ();
 sg13g2_decap_8 FILLER_33_838 ();
 sg13g2_decap_8 FILLER_33_845 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_decap_8 FILLER_33_859 ();
 sg13g2_decap_8 FILLER_33_866 ();
 sg13g2_decap_4 FILLER_33_873 ();
 sg13g2_fill_1 FILLER_33_877 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_decap_8 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_232 ();
 sg13g2_decap_8 FILLER_34_239 ();
 sg13g2_decap_8 FILLER_34_246 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_decap_4 FILLER_34_260 ();
 sg13g2_decap_4 FILLER_34_280 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_330 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_decap_4 FILLER_34_376 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_fill_2 FILLER_34_389 ();
 sg13g2_fill_1 FILLER_34_400 ();
 sg13g2_fill_1 FILLER_34_406 ();
 sg13g2_fill_2 FILLER_34_437 ();
 sg13g2_fill_2 FILLER_34_482 ();
 sg13g2_fill_2 FILLER_34_496 ();
 sg13g2_fill_1 FILLER_34_536 ();
 sg13g2_decap_8 FILLER_34_549 ();
 sg13g2_decap_8 FILLER_34_556 ();
 sg13g2_fill_1 FILLER_34_573 ();
 sg13g2_fill_2 FILLER_34_579 ();
 sg13g2_fill_2 FILLER_34_614 ();
 sg13g2_decap_8 FILLER_34_620 ();
 sg13g2_decap_4 FILLER_34_627 ();
 sg13g2_decap_8 FILLER_34_667 ();
 sg13g2_decap_8 FILLER_34_674 ();
 sg13g2_decap_8 FILLER_34_681 ();
 sg13g2_decap_4 FILLER_34_688 ();
 sg13g2_decap_8 FILLER_34_695 ();
 sg13g2_decap_8 FILLER_34_702 ();
 sg13g2_decap_8 FILLER_34_709 ();
 sg13g2_decap_8 FILLER_34_716 ();
 sg13g2_decap_8 FILLER_34_723 ();
 sg13g2_decap_8 FILLER_34_730 ();
 sg13g2_decap_8 FILLER_34_737 ();
 sg13g2_decap_8 FILLER_34_744 ();
 sg13g2_decap_8 FILLER_34_751 ();
 sg13g2_decap_8 FILLER_34_758 ();
 sg13g2_decap_8 FILLER_34_765 ();
 sg13g2_decap_8 FILLER_34_772 ();
 sg13g2_decap_8 FILLER_34_779 ();
 sg13g2_decap_8 FILLER_34_786 ();
 sg13g2_decap_8 FILLER_34_793 ();
 sg13g2_decap_8 FILLER_34_800 ();
 sg13g2_decap_8 FILLER_34_807 ();
 sg13g2_decap_8 FILLER_34_814 ();
 sg13g2_decap_8 FILLER_34_821 ();
 sg13g2_decap_8 FILLER_34_828 ();
 sg13g2_decap_8 FILLER_34_835 ();
 sg13g2_decap_8 FILLER_34_842 ();
 sg13g2_decap_8 FILLER_34_849 ();
 sg13g2_decap_8 FILLER_34_856 ();
 sg13g2_decap_8 FILLER_34_863 ();
 sg13g2_decap_8 FILLER_34_870 ();
 sg13g2_fill_1 FILLER_34_877 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_4 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_decap_8 FILLER_35_253 ();
 sg13g2_decap_4 FILLER_35_260 ();
 sg13g2_fill_1 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_331 ();
 sg13g2_fill_1 FILLER_35_336 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_353 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_fill_2 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_372 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_395 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_fill_1 FILLER_35_430 ();
 sg13g2_fill_2 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_459 ();
 sg13g2_fill_2 FILLER_35_496 ();
 sg13g2_fill_1 FILLER_35_498 ();
 sg13g2_fill_2 FILLER_35_530 ();
 sg13g2_fill_1 FILLER_35_532 ();
 sg13g2_fill_2 FILLER_35_555 ();
 sg13g2_fill_2 FILLER_35_563 ();
 sg13g2_fill_2 FILLER_35_585 ();
 sg13g2_fill_1 FILLER_35_647 ();
 sg13g2_decap_8 FILLER_35_674 ();
 sg13g2_fill_1 FILLER_35_681 ();
 sg13g2_fill_1 FILLER_35_691 ();
 sg13g2_decap_8 FILLER_35_718 ();
 sg13g2_decap_8 FILLER_35_725 ();
 sg13g2_decap_8 FILLER_35_732 ();
 sg13g2_decap_8 FILLER_35_739 ();
 sg13g2_decap_8 FILLER_35_746 ();
 sg13g2_decap_8 FILLER_35_753 ();
 sg13g2_decap_8 FILLER_35_760 ();
 sg13g2_decap_8 FILLER_35_767 ();
 sg13g2_decap_8 FILLER_35_774 ();
 sg13g2_decap_8 FILLER_35_781 ();
 sg13g2_decap_8 FILLER_35_788 ();
 sg13g2_decap_8 FILLER_35_795 ();
 sg13g2_decap_8 FILLER_35_802 ();
 sg13g2_decap_8 FILLER_35_809 ();
 sg13g2_decap_8 FILLER_35_816 ();
 sg13g2_decap_8 FILLER_35_823 ();
 sg13g2_decap_8 FILLER_35_830 ();
 sg13g2_decap_8 FILLER_35_837 ();
 sg13g2_decap_8 FILLER_35_844 ();
 sg13g2_decap_8 FILLER_35_851 ();
 sg13g2_decap_8 FILLER_35_858 ();
 sg13g2_decap_8 FILLER_35_865 ();
 sg13g2_decap_4 FILLER_35_872 ();
 sg13g2_fill_2 FILLER_35_876 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_4 FILLER_36_231 ();
 sg13g2_fill_2 FILLER_36_265 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_fill_1 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_365 ();
 sg13g2_fill_1 FILLER_36_397 ();
 sg13g2_fill_1 FILLER_36_422 ();
 sg13g2_fill_1 FILLER_36_443 ();
 sg13g2_fill_2 FILLER_36_473 ();
 sg13g2_fill_1 FILLER_36_475 ();
 sg13g2_fill_2 FILLER_36_480 ();
 sg13g2_fill_1 FILLER_36_482 ();
 sg13g2_fill_1 FILLER_36_488 ();
 sg13g2_fill_1 FILLER_36_494 ();
 sg13g2_fill_1 FILLER_36_500 ();
 sg13g2_fill_1 FILLER_36_512 ();
 sg13g2_fill_2 FILLER_36_548 ();
 sg13g2_fill_2 FILLER_36_640 ();
 sg13g2_fill_1 FILLER_36_668 ();
 sg13g2_decap_8 FILLER_36_719 ();
 sg13g2_decap_8 FILLER_36_726 ();
 sg13g2_decap_8 FILLER_36_733 ();
 sg13g2_decap_8 FILLER_36_740 ();
 sg13g2_decap_8 FILLER_36_747 ();
 sg13g2_decap_8 FILLER_36_754 ();
 sg13g2_decap_8 FILLER_36_761 ();
 sg13g2_decap_8 FILLER_36_768 ();
 sg13g2_decap_8 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_782 ();
 sg13g2_decap_8 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_796 ();
 sg13g2_decap_8 FILLER_36_803 ();
 sg13g2_decap_8 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_8 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_838 ();
 sg13g2_decap_8 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_decap_8 FILLER_36_859 ();
 sg13g2_decap_8 FILLER_36_866 ();
 sg13g2_decap_4 FILLER_36_873 ();
 sg13g2_fill_1 FILLER_36_877 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_207 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_221 ();
 sg13g2_fill_1 FILLER_37_290 ();
 sg13g2_fill_2 FILLER_37_323 ();
 sg13g2_fill_1 FILLER_37_325 ();
 sg13g2_fill_2 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_341 ();
 sg13g2_fill_1 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_348 ();
 sg13g2_fill_2 FILLER_37_353 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_fill_1 FILLER_37_366 ();
 sg13g2_fill_2 FILLER_37_371 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_fill_1 FILLER_37_392 ();
 sg13g2_fill_1 FILLER_37_397 ();
 sg13g2_fill_1 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_411 ();
 sg13g2_fill_1 FILLER_37_416 ();
 sg13g2_decap_4 FILLER_37_435 ();
 sg13g2_fill_1 FILLER_37_461 ();
 sg13g2_fill_1 FILLER_37_466 ();
 sg13g2_fill_2 FILLER_37_479 ();
 sg13g2_decap_8 FILLER_37_503 ();
 sg13g2_fill_2 FILLER_37_541 ();
 sg13g2_fill_1 FILLER_37_548 ();
 sg13g2_fill_2 FILLER_37_553 ();
 sg13g2_fill_1 FILLER_37_560 ();
 sg13g2_fill_1 FILLER_37_614 ();
 sg13g2_fill_1 FILLER_37_690 ();
 sg13g2_decap_8 FILLER_37_720 ();
 sg13g2_fill_1 FILLER_37_727 ();
 sg13g2_decap_8 FILLER_37_732 ();
 sg13g2_decap_8 FILLER_37_739 ();
 sg13g2_decap_8 FILLER_37_746 ();
 sg13g2_decap_8 FILLER_37_753 ();
 sg13g2_decap_8 FILLER_37_760 ();
 sg13g2_decap_8 FILLER_37_767 ();
 sg13g2_decap_8 FILLER_37_774 ();
 sg13g2_decap_8 FILLER_37_781 ();
 sg13g2_decap_8 FILLER_37_788 ();
 sg13g2_decap_8 FILLER_37_795 ();
 sg13g2_decap_8 FILLER_37_802 ();
 sg13g2_decap_8 FILLER_37_809 ();
 sg13g2_decap_8 FILLER_37_816 ();
 sg13g2_decap_8 FILLER_37_823 ();
 sg13g2_decap_8 FILLER_37_830 ();
 sg13g2_decap_8 FILLER_37_837 ();
 sg13g2_decap_8 FILLER_37_844 ();
 sg13g2_decap_8 FILLER_37_851 ();
 sg13g2_decap_8 FILLER_37_858 ();
 sg13g2_decap_8 FILLER_37_865 ();
 sg13g2_decap_4 FILLER_37_872 ();
 sg13g2_fill_2 FILLER_37_876 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_261 ();
 sg13g2_fill_1 FILLER_38_287 ();
 sg13g2_decap_4 FILLER_38_354 ();
 sg13g2_fill_2 FILLER_38_358 ();
 sg13g2_decap_4 FILLER_38_417 ();
 sg13g2_fill_2 FILLER_38_430 ();
 sg13g2_fill_2 FILLER_38_436 ();
 sg13g2_fill_1 FILLER_38_438 ();
 sg13g2_fill_1 FILLER_38_443 ();
 sg13g2_fill_1 FILLER_38_454 ();
 sg13g2_fill_1 FILLER_38_481 ();
 sg13g2_fill_1 FILLER_38_508 ();
 sg13g2_fill_1 FILLER_38_535 ();
 sg13g2_fill_1 FILLER_38_540 ();
 sg13g2_fill_2 FILLER_38_603 ();
 sg13g2_fill_1 FILLER_38_634 ();
 sg13g2_fill_1 FILLER_38_647 ();
 sg13g2_fill_1 FILLER_38_683 ();
 sg13g2_fill_2 FILLER_38_717 ();
 sg13g2_decap_8 FILLER_38_732 ();
 sg13g2_decap_8 FILLER_38_739 ();
 sg13g2_decap_8 FILLER_38_746 ();
 sg13g2_decap_8 FILLER_38_753 ();
 sg13g2_decap_8 FILLER_38_760 ();
 sg13g2_decap_8 FILLER_38_767 ();
 sg13g2_decap_8 FILLER_38_774 ();
 sg13g2_decap_8 FILLER_38_781 ();
 sg13g2_decap_8 FILLER_38_788 ();
 sg13g2_decap_8 FILLER_38_795 ();
 sg13g2_decap_8 FILLER_38_802 ();
 sg13g2_decap_8 FILLER_38_809 ();
 sg13g2_decap_8 FILLER_38_816 ();
 sg13g2_decap_8 FILLER_38_823 ();
 sg13g2_decap_8 FILLER_38_830 ();
 sg13g2_decap_8 FILLER_38_837 ();
 sg13g2_decap_8 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_decap_8 FILLER_38_858 ();
 sg13g2_decap_8 FILLER_38_865 ();
 sg13g2_decap_4 FILLER_38_872 ();
 sg13g2_fill_2 FILLER_38_876 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_4 FILLER_39_189 ();
 sg13g2_fill_2 FILLER_39_193 ();
 sg13g2_decap_4 FILLER_39_200 ();
 sg13g2_fill_1 FILLER_39_204 ();
 sg13g2_fill_2 FILLER_39_239 ();
 sg13g2_fill_1 FILLER_39_257 ();
 sg13g2_fill_1 FILLER_39_264 ();
 sg13g2_fill_1 FILLER_39_272 ();
 sg13g2_fill_2 FILLER_39_278 ();
 sg13g2_fill_1 FILLER_39_285 ();
 sg13g2_fill_1 FILLER_39_294 ();
 sg13g2_fill_1 FILLER_39_299 ();
 sg13g2_fill_1 FILLER_39_305 ();
 sg13g2_fill_1 FILLER_39_311 ();
 sg13g2_fill_1 FILLER_39_316 ();
 sg13g2_fill_1 FILLER_39_338 ();
 sg13g2_fill_1 FILLER_39_420 ();
 sg13g2_fill_2 FILLER_39_425 ();
 sg13g2_decap_8 FILLER_39_431 ();
 sg13g2_fill_2 FILLER_39_438 ();
 sg13g2_fill_1 FILLER_39_444 ();
 sg13g2_fill_2 FILLER_39_471 ();
 sg13g2_fill_2 FILLER_39_477 ();
 sg13g2_fill_1 FILLER_39_489 ();
 sg13g2_decap_4 FILLER_39_495 ();
 sg13g2_fill_2 FILLER_39_499 ();
 sg13g2_fill_1 FILLER_39_523 ();
 sg13g2_fill_2 FILLER_39_529 ();
 sg13g2_fill_2 FILLER_39_535 ();
 sg13g2_fill_1 FILLER_39_537 ();
 sg13g2_fill_1 FILLER_39_583 ();
 sg13g2_fill_2 FILLER_39_621 ();
 sg13g2_fill_1 FILLER_39_683 ();
 sg13g2_fill_1 FILLER_39_689 ();
 sg13g2_decap_8 FILLER_39_715 ();
 sg13g2_decap_8 FILLER_39_736 ();
 sg13g2_decap_8 FILLER_39_743 ();
 sg13g2_decap_8 FILLER_39_750 ();
 sg13g2_decap_8 FILLER_39_757 ();
 sg13g2_decap_8 FILLER_39_764 ();
 sg13g2_decap_8 FILLER_39_771 ();
 sg13g2_decap_8 FILLER_39_778 ();
 sg13g2_decap_8 FILLER_39_785 ();
 sg13g2_decap_8 FILLER_39_792 ();
 sg13g2_decap_8 FILLER_39_799 ();
 sg13g2_decap_8 FILLER_39_806 ();
 sg13g2_decap_8 FILLER_39_813 ();
 sg13g2_decap_8 FILLER_39_820 ();
 sg13g2_decap_8 FILLER_39_827 ();
 sg13g2_decap_8 FILLER_39_834 ();
 sg13g2_decap_8 FILLER_39_841 ();
 sg13g2_decap_8 FILLER_39_848 ();
 sg13g2_decap_8 FILLER_39_855 ();
 sg13g2_decap_8 FILLER_39_862 ();
 sg13g2_decap_8 FILLER_39_869 ();
 sg13g2_fill_2 FILLER_39_876 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_4 FILLER_40_168 ();
 sg13g2_decap_4 FILLER_40_198 ();
 sg13g2_fill_1 FILLER_40_232 ();
 sg13g2_fill_2 FILLER_40_238 ();
 sg13g2_fill_2 FILLER_40_289 ();
 sg13g2_fill_2 FILLER_40_295 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_1 FILLER_40_309 ();
 sg13g2_fill_2 FILLER_40_315 ();
 sg13g2_fill_1 FILLER_40_325 ();
 sg13g2_fill_2 FILLER_40_335 ();
 sg13g2_fill_2 FILLER_40_358 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_fill_1 FILLER_40_365 ();
 sg13g2_fill_2 FILLER_40_370 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_2 FILLER_40_381 ();
 sg13g2_fill_1 FILLER_40_383 ();
 sg13g2_fill_2 FILLER_40_389 ();
 sg13g2_fill_1 FILLER_40_391 ();
 sg13g2_fill_2 FILLER_40_409 ();
 sg13g2_fill_1 FILLER_40_452 ();
 sg13g2_fill_1 FILLER_40_461 ();
 sg13g2_fill_1 FILLER_40_467 ();
 sg13g2_fill_2 FILLER_40_473 ();
 sg13g2_fill_2 FILLER_40_479 ();
 sg13g2_fill_1 FILLER_40_481 ();
 sg13g2_fill_1 FILLER_40_506 ();
 sg13g2_fill_2 FILLER_40_523 ();
 sg13g2_fill_2 FILLER_40_539 ();
 sg13g2_fill_1 FILLER_40_570 ();
 sg13g2_fill_1 FILLER_40_621 ();
 sg13g2_fill_1 FILLER_40_626 ();
 sg13g2_decap_4 FILLER_40_688 ();
 sg13g2_fill_1 FILLER_40_692 ();
 sg13g2_fill_2 FILLER_40_705 ();
 sg13g2_fill_2 FILLER_40_711 ();
 sg13g2_fill_2 FILLER_40_725 ();
 sg13g2_fill_2 FILLER_40_730 ();
 sg13g2_decap_8 FILLER_40_745 ();
 sg13g2_decap_8 FILLER_40_752 ();
 sg13g2_decap_8 FILLER_40_759 ();
 sg13g2_decap_8 FILLER_40_766 ();
 sg13g2_decap_8 FILLER_40_773 ();
 sg13g2_decap_8 FILLER_40_780 ();
 sg13g2_decap_8 FILLER_40_787 ();
 sg13g2_decap_8 FILLER_40_794 ();
 sg13g2_decap_8 FILLER_40_801 ();
 sg13g2_decap_8 FILLER_40_808 ();
 sg13g2_decap_8 FILLER_40_815 ();
 sg13g2_decap_8 FILLER_40_822 ();
 sg13g2_decap_8 FILLER_40_829 ();
 sg13g2_decap_8 FILLER_40_836 ();
 sg13g2_decap_8 FILLER_40_843 ();
 sg13g2_decap_8 FILLER_40_850 ();
 sg13g2_decap_8 FILLER_40_857 ();
 sg13g2_decap_8 FILLER_40_864 ();
 sg13g2_decap_8 FILLER_40_871 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_4 FILLER_41_161 ();
 sg13g2_fill_1 FILLER_41_165 ();
 sg13g2_decap_4 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_184 ();
 sg13g2_fill_2 FILLER_41_195 ();
 sg13g2_fill_1 FILLER_41_207 ();
 sg13g2_fill_2 FILLER_41_216 ();
 sg13g2_fill_1 FILLER_41_222 ();
 sg13g2_fill_2 FILLER_41_258 ();
 sg13g2_fill_1 FILLER_41_260 ();
 sg13g2_fill_2 FILLER_41_286 ();
 sg13g2_fill_1 FILLER_41_293 ();
 sg13g2_fill_2 FILLER_41_355 ();
 sg13g2_fill_1 FILLER_41_378 ();
 sg13g2_fill_1 FILLER_41_405 ();
 sg13g2_fill_1 FILLER_41_410 ();
 sg13g2_fill_1 FILLER_41_416 ();
 sg13g2_fill_1 FILLER_41_427 ();
 sg13g2_decap_4 FILLER_41_438 ();
 sg13g2_fill_1 FILLER_41_451 ();
 sg13g2_fill_1 FILLER_41_458 ();
 sg13g2_fill_1 FILLER_41_462 ();
 sg13g2_fill_1 FILLER_41_479 ();
 sg13g2_fill_1 FILLER_41_485 ();
 sg13g2_fill_1 FILLER_41_494 ();
 sg13g2_decap_4 FILLER_41_499 ();
 sg13g2_fill_1 FILLER_41_503 ();
 sg13g2_fill_1 FILLER_41_538 ();
 sg13g2_fill_2 FILLER_41_558 ();
 sg13g2_fill_2 FILLER_41_575 ();
 sg13g2_fill_2 FILLER_41_585 ();
 sg13g2_fill_2 FILLER_41_591 ();
 sg13g2_fill_2 FILLER_41_626 ();
 sg13g2_fill_1 FILLER_41_633 ();
 sg13g2_fill_2 FILLER_41_649 ();
 sg13g2_fill_1 FILLER_41_651 ();
 sg13g2_fill_1 FILLER_41_665 ();
 sg13g2_decap_4 FILLER_41_690 ();
 sg13g2_fill_2 FILLER_41_694 ();
 sg13g2_decap_4 FILLER_41_704 ();
 sg13g2_fill_2 FILLER_41_708 ();
 sg13g2_fill_2 FILLER_41_714 ();
 sg13g2_fill_1 FILLER_41_721 ();
 sg13g2_fill_2 FILLER_41_725 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_decap_8 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_fill_2 FILLER_41_875 ();
 sg13g2_fill_1 FILLER_41_877 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_4 FILLER_42_140 ();
 sg13g2_fill_2 FILLER_42_175 ();
 sg13g2_fill_1 FILLER_42_181 ();
 sg13g2_fill_2 FILLER_42_192 ();
 sg13g2_fill_1 FILLER_42_235 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_fill_2 FILLER_42_273 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_fill_1 FILLER_42_301 ();
 sg13g2_fill_1 FILLER_42_307 ();
 sg13g2_fill_2 FILLER_42_316 ();
 sg13g2_decap_4 FILLER_42_326 ();
 sg13g2_decap_8 FILLER_42_334 ();
 sg13g2_fill_2 FILLER_42_346 ();
 sg13g2_fill_2 FILLER_42_369 ();
 sg13g2_fill_1 FILLER_42_371 ();
 sg13g2_fill_1 FILLER_42_394 ();
 sg13g2_fill_1 FILLER_42_415 ();
 sg13g2_decap_4 FILLER_42_443 ();
 sg13g2_decap_4 FILLER_42_463 ();
 sg13g2_fill_1 FILLER_42_467 ();
 sg13g2_fill_1 FILLER_42_488 ();
 sg13g2_fill_2 FILLER_42_498 ();
 sg13g2_fill_1 FILLER_42_500 ();
 sg13g2_fill_1 FILLER_42_506 ();
 sg13g2_fill_2 FILLER_42_511 ();
 sg13g2_fill_2 FILLER_42_518 ();
 sg13g2_fill_2 FILLER_42_524 ();
 sg13g2_fill_1 FILLER_42_526 ();
 sg13g2_fill_1 FILLER_42_550 ();
 sg13g2_fill_2 FILLER_42_555 ();
 sg13g2_fill_2 FILLER_42_598 ();
 sg13g2_fill_2 FILLER_42_626 ();
 sg13g2_fill_2 FILLER_42_673 ();
 sg13g2_fill_1 FILLER_42_675 ();
 sg13g2_fill_2 FILLER_42_709 ();
 sg13g2_fill_1 FILLER_42_711 ();
 sg13g2_decap_8 FILLER_42_759 ();
 sg13g2_decap_8 FILLER_42_766 ();
 sg13g2_decap_8 FILLER_42_773 ();
 sg13g2_decap_8 FILLER_42_780 ();
 sg13g2_decap_8 FILLER_42_787 ();
 sg13g2_decap_8 FILLER_42_794 ();
 sg13g2_decap_8 FILLER_42_801 ();
 sg13g2_decap_8 FILLER_42_808 ();
 sg13g2_decap_8 FILLER_42_815 ();
 sg13g2_decap_8 FILLER_42_822 ();
 sg13g2_decap_8 FILLER_42_829 ();
 sg13g2_decap_8 FILLER_42_836 ();
 sg13g2_decap_8 FILLER_42_843 ();
 sg13g2_decap_8 FILLER_42_850 ();
 sg13g2_decap_8 FILLER_42_857 ();
 sg13g2_decap_8 FILLER_42_864 ();
 sg13g2_decap_8 FILLER_42_871 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_fill_2 FILLER_43_133 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_decap_4 FILLER_43_146 ();
 sg13g2_decap_4 FILLER_43_154 ();
 sg13g2_fill_2 FILLER_43_158 ();
 sg13g2_fill_1 FILLER_43_278 ();
 sg13g2_fill_2 FILLER_43_297 ();
 sg13g2_fill_2 FILLER_43_303 ();
 sg13g2_fill_2 FILLER_43_309 ();
 sg13g2_fill_2 FILLER_43_315 ();
 sg13g2_fill_2 FILLER_43_373 ();
 sg13g2_fill_1 FILLER_43_383 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_414 ();
 sg13g2_fill_2 FILLER_43_434 ();
 sg13g2_decap_4 FILLER_43_442 ();
 sg13g2_fill_2 FILLER_43_446 ();
 sg13g2_fill_1 FILLER_43_478 ();
 sg13g2_fill_2 FILLER_43_488 ();
 sg13g2_fill_1 FILLER_43_498 ();
 sg13g2_fill_2 FILLER_43_512 ();
 sg13g2_decap_4 FILLER_43_540 ();
 sg13g2_fill_2 FILLER_43_574 ();
 sg13g2_fill_1 FILLER_43_584 ();
 sg13g2_fill_2 FILLER_43_654 ();
 sg13g2_fill_1 FILLER_43_656 ();
 sg13g2_fill_2 FILLER_43_679 ();
 sg13g2_fill_2 FILLER_43_697 ();
 sg13g2_fill_1 FILLER_43_746 ();
 sg13g2_fill_2 FILLER_43_755 ();
 sg13g2_decap_4 FILLER_43_765 ();
 sg13g2_fill_1 FILLER_43_769 ();
 sg13g2_decap_8 FILLER_43_786 ();
 sg13g2_decap_8 FILLER_43_793 ();
 sg13g2_decap_8 FILLER_43_800 ();
 sg13g2_decap_8 FILLER_43_807 ();
 sg13g2_decap_8 FILLER_43_814 ();
 sg13g2_decap_8 FILLER_43_821 ();
 sg13g2_decap_8 FILLER_43_828 ();
 sg13g2_decap_8 FILLER_43_835 ();
 sg13g2_decap_8 FILLER_43_842 ();
 sg13g2_decap_8 FILLER_43_849 ();
 sg13g2_decap_8 FILLER_43_856 ();
 sg13g2_decap_8 FILLER_43_863 ();
 sg13g2_decap_8 FILLER_43_870 ();
 sg13g2_fill_1 FILLER_43_877 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_fill_1 FILLER_44_171 ();
 sg13g2_fill_1 FILLER_44_178 ();
 sg13g2_fill_1 FILLER_44_189 ();
 sg13g2_fill_1 FILLER_44_200 ();
 sg13g2_fill_1 FILLER_44_207 ();
 sg13g2_decap_4 FILLER_44_223 ();
 sg13g2_fill_1 FILLER_44_227 ();
 sg13g2_decap_4 FILLER_44_233 ();
 sg13g2_decap_4 FILLER_44_247 ();
 sg13g2_fill_2 FILLER_44_277 ();
 sg13g2_fill_1 FILLER_44_279 ();
 sg13g2_fill_2 FILLER_44_285 ();
 sg13g2_fill_1 FILLER_44_295 ();
 sg13g2_fill_2 FILLER_44_301 ();
 sg13g2_fill_2 FILLER_44_307 ();
 sg13g2_fill_2 FILLER_44_317 ();
 sg13g2_fill_1 FILLER_44_319 ();
 sg13g2_fill_1 FILLER_44_324 ();
 sg13g2_fill_2 FILLER_44_346 ();
 sg13g2_fill_1 FILLER_44_358 ();
 sg13g2_fill_2 FILLER_44_367 ();
 sg13g2_fill_1 FILLER_44_379 ();
 sg13g2_fill_1 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_437 ();
 sg13g2_fill_1 FILLER_44_464 ();
 sg13g2_fill_2 FILLER_44_525 ();
 sg13g2_fill_1 FILLER_44_534 ();
 sg13g2_fill_2 FILLER_44_543 ();
 sg13g2_fill_1 FILLER_44_545 ();
 sg13g2_fill_1 FILLER_44_550 ();
 sg13g2_decap_4 FILLER_44_567 ();
 sg13g2_fill_1 FILLER_44_571 ();
 sg13g2_fill_1 FILLER_44_608 ();
 sg13g2_fill_1 FILLER_44_623 ();
 sg13g2_fill_2 FILLER_44_686 ();
 sg13g2_fill_1 FILLER_44_703 ();
 sg13g2_fill_2 FILLER_44_746 ();
 sg13g2_fill_2 FILLER_44_753 ();
 sg13g2_fill_1 FILLER_44_755 ();
 sg13g2_fill_2 FILLER_44_764 ();
 sg13g2_decap_8 FILLER_44_788 ();
 sg13g2_decap_8 FILLER_44_795 ();
 sg13g2_decap_8 FILLER_44_802 ();
 sg13g2_decap_8 FILLER_44_809 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_8 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_8 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_44_865 ();
 sg13g2_decap_4 FILLER_44_872 ();
 sg13g2_fill_2 FILLER_44_876 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_fill_2 FILLER_45_126 ();
 sg13g2_fill_2 FILLER_45_227 ();
 sg13g2_fill_1 FILLER_45_229 ();
 sg13g2_fill_2 FILLER_45_272 ();
 sg13g2_fill_1 FILLER_45_274 ();
 sg13g2_fill_2 FILLER_45_320 ();
 sg13g2_fill_2 FILLER_45_351 ();
 sg13g2_fill_1 FILLER_45_353 ();
 sg13g2_fill_1 FILLER_45_380 ();
 sg13g2_fill_1 FILLER_45_449 ();
 sg13g2_fill_1 FILLER_45_455 ();
 sg13g2_fill_2 FILLER_45_460 ();
 sg13g2_fill_1 FILLER_45_462 ();
 sg13g2_fill_2 FILLER_45_471 ();
 sg13g2_fill_1 FILLER_45_473 ();
 sg13g2_fill_2 FILLER_45_512 ();
 sg13g2_fill_1 FILLER_45_514 ();
 sg13g2_fill_1 FILLER_45_546 ();
 sg13g2_decap_4 FILLER_45_564 ();
 sg13g2_fill_1 FILLER_45_568 ();
 sg13g2_fill_1 FILLER_45_598 ();
 sg13g2_fill_1 FILLER_45_607 ();
 sg13g2_fill_1 FILLER_45_616 ();
 sg13g2_fill_2 FILLER_45_632 ();
 sg13g2_fill_1 FILLER_45_650 ();
 sg13g2_fill_2 FILLER_45_659 ();
 sg13g2_fill_1 FILLER_45_661 ();
 sg13g2_fill_2 FILLER_45_678 ();
 sg13g2_fill_2 FILLER_45_688 ();
 sg13g2_fill_1 FILLER_45_690 ();
 sg13g2_fill_1 FILLER_45_710 ();
 sg13g2_fill_2 FILLER_45_736 ();
 sg13g2_fill_1 FILLER_45_738 ();
 sg13g2_decap_8 FILLER_45_755 ();
 sg13g2_fill_2 FILLER_45_762 ();
 sg13g2_fill_2 FILLER_45_777 ();
 sg13g2_decap_8 FILLER_45_792 ();
 sg13g2_decap_8 FILLER_45_799 ();
 sg13g2_decap_8 FILLER_45_806 ();
 sg13g2_decap_8 FILLER_45_813 ();
 sg13g2_decap_8 FILLER_45_820 ();
 sg13g2_decap_8 FILLER_45_827 ();
 sg13g2_decap_8 FILLER_45_834 ();
 sg13g2_decap_8 FILLER_45_841 ();
 sg13g2_decap_8 FILLER_45_848 ();
 sg13g2_decap_8 FILLER_45_855 ();
 sg13g2_decap_8 FILLER_45_862 ();
 sg13g2_decap_8 FILLER_45_869 ();
 sg13g2_fill_2 FILLER_45_876 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_4 FILLER_46_112 ();
 sg13g2_fill_1 FILLER_46_116 ();
 sg13g2_decap_8 FILLER_46_121 ();
 sg13g2_fill_1 FILLER_46_128 ();
 sg13g2_fill_2 FILLER_46_143 ();
 sg13g2_fill_1 FILLER_46_162 ();
 sg13g2_fill_1 FILLER_46_167 ();
 sg13g2_fill_1 FILLER_46_174 ();
 sg13g2_fill_1 FILLER_46_180 ();
 sg13g2_fill_2 FILLER_46_185 ();
 sg13g2_fill_1 FILLER_46_197 ();
 sg13g2_fill_2 FILLER_46_224 ();
 sg13g2_fill_1 FILLER_46_249 ();
 sg13g2_fill_2 FILLER_46_276 ();
 sg13g2_fill_2 FILLER_46_291 ();
 sg13g2_fill_2 FILLER_46_297 ();
 sg13g2_fill_2 FILLER_46_332 ();
 sg13g2_fill_1 FILLER_46_334 ();
 sg13g2_fill_1 FILLER_46_361 ();
 sg13g2_fill_1 FILLER_46_366 ();
 sg13g2_fill_1 FILLER_46_371 ();
 sg13g2_fill_2 FILLER_46_402 ();
 sg13g2_fill_2 FILLER_46_420 ();
 sg13g2_fill_1 FILLER_46_422 ();
 sg13g2_decap_4 FILLER_46_427 ();
 sg13g2_fill_1 FILLER_46_431 ();
 sg13g2_fill_2 FILLER_46_458 ();
 sg13g2_fill_2 FILLER_46_472 ();
 sg13g2_fill_1 FILLER_46_474 ();
 sg13g2_fill_2 FILLER_46_519 ();
 sg13g2_decap_4 FILLER_46_525 ();
 sg13g2_fill_1 FILLER_46_540 ();
 sg13g2_fill_2 FILLER_46_545 ();
 sg13g2_fill_1 FILLER_46_602 ();
 sg13g2_fill_2 FILLER_46_651 ();
 sg13g2_fill_1 FILLER_46_653 ();
 sg13g2_fill_1 FILLER_46_659 ();
 sg13g2_fill_1 FILLER_46_665 ();
 sg13g2_fill_1 FILLER_46_671 ();
 sg13g2_fill_1 FILLER_46_680 ();
 sg13g2_fill_2 FILLER_46_689 ();
 sg13g2_decap_4 FILLER_46_696 ();
 sg13g2_fill_1 FILLER_46_705 ();
 sg13g2_decap_4 FILLER_46_717 ();
 sg13g2_decap_8 FILLER_46_739 ();
 sg13g2_fill_2 FILLER_46_754 ();
 sg13g2_decap_8 FILLER_46_792 ();
 sg13g2_decap_8 FILLER_46_799 ();
 sg13g2_decap_8 FILLER_46_806 ();
 sg13g2_decap_8 FILLER_46_813 ();
 sg13g2_decap_8 FILLER_46_820 ();
 sg13g2_decap_8 FILLER_46_827 ();
 sg13g2_decap_8 FILLER_46_834 ();
 sg13g2_decap_8 FILLER_46_841 ();
 sg13g2_decap_8 FILLER_46_848 ();
 sg13g2_decap_8 FILLER_46_855 ();
 sg13g2_decap_8 FILLER_46_862 ();
 sg13g2_decap_8 FILLER_46_869 ();
 sg13g2_fill_2 FILLER_46_876 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_4 FILLER_47_105 ();
 sg13g2_fill_1 FILLER_47_109 ();
 sg13g2_decap_4 FILLER_47_136 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_fill_2 FILLER_47_217 ();
 sg13g2_fill_1 FILLER_47_246 ();
 sg13g2_fill_2 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_258 ();
 sg13g2_decap_8 FILLER_47_286 ();
 sg13g2_fill_2 FILLER_47_293 ();
 sg13g2_fill_2 FILLER_47_303 ();
 sg13g2_fill_1 FILLER_47_310 ();
 sg13g2_fill_1 FILLER_47_315 ();
 sg13g2_fill_1 FILLER_47_325 ();
 sg13g2_decap_8 FILLER_47_330 ();
 sg13g2_fill_1 FILLER_47_337 ();
 sg13g2_fill_1 FILLER_47_342 ();
 sg13g2_decap_4 FILLER_47_386 ();
 sg13g2_fill_1 FILLER_47_390 ();
 sg13g2_fill_2 FILLER_47_408 ();
 sg13g2_fill_2 FILLER_47_415 ();
 sg13g2_fill_1 FILLER_47_417 ();
 sg13g2_fill_2 FILLER_47_431 ();
 sg13g2_fill_2 FILLER_47_467 ();
 sg13g2_fill_1 FILLER_47_469 ();
 sg13g2_fill_2 FILLER_47_526 ();
 sg13g2_fill_1 FILLER_47_528 ();
 sg13g2_fill_1 FILLER_47_555 ();
 sg13g2_decap_4 FILLER_47_572 ();
 sg13g2_fill_2 FILLER_47_613 ();
 sg13g2_fill_1 FILLER_47_615 ();
 sg13g2_fill_2 FILLER_47_655 ();
 sg13g2_decap_8 FILLER_47_669 ();
 sg13g2_fill_1 FILLER_47_676 ();
 sg13g2_fill_2 FILLER_47_685 ();
 sg13g2_fill_2 FILLER_47_695 ();
 sg13g2_fill_1 FILLER_47_697 ();
 sg13g2_fill_1 FILLER_47_703 ();
 sg13g2_decap_4 FILLER_47_712 ();
 sg13g2_fill_1 FILLER_47_726 ();
 sg13g2_fill_1 FILLER_47_740 ();
 sg13g2_fill_2 FILLER_47_750 ();
 sg13g2_fill_2 FILLER_47_763 ();
 sg13g2_fill_1 FILLER_47_765 ();
 sg13g2_fill_2 FILLER_47_788 ();
 sg13g2_fill_1 FILLER_47_797 ();
 sg13g2_decap_8 FILLER_47_811 ();
 sg13g2_decap_8 FILLER_47_828 ();
 sg13g2_decap_8 FILLER_47_835 ();
 sg13g2_decap_8 FILLER_47_842 ();
 sg13g2_decap_8 FILLER_47_849 ();
 sg13g2_decap_8 FILLER_47_856 ();
 sg13g2_decap_8 FILLER_47_863 ();
 sg13g2_decap_8 FILLER_47_870 ();
 sg13g2_fill_1 FILLER_47_877 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_fill_2 FILLER_48_98 ();
 sg13g2_fill_2 FILLER_48_140 ();
 sg13g2_fill_2 FILLER_48_152 ();
 sg13g2_fill_1 FILLER_48_154 ();
 sg13g2_fill_1 FILLER_48_181 ();
 sg13g2_fill_2 FILLER_48_230 ();
 sg13g2_fill_1 FILLER_48_232 ();
 sg13g2_fill_1 FILLER_48_280 ();
 sg13g2_fill_2 FILLER_48_285 ();
 sg13g2_decap_8 FILLER_48_292 ();
 sg13g2_fill_1 FILLER_48_308 ();
 sg13g2_fill_1 FILLER_48_320 ();
 sg13g2_fill_1 FILLER_48_329 ();
 sg13g2_fill_1 FILLER_48_370 ();
 sg13g2_fill_1 FILLER_48_375 ();
 sg13g2_fill_1 FILLER_48_380 ();
 sg13g2_fill_2 FILLER_48_390 ();
 sg13g2_fill_1 FILLER_48_392 ();
 sg13g2_fill_2 FILLER_48_417 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_fill_1 FILLER_48_434 ();
 sg13g2_fill_1 FILLER_48_440 ();
 sg13g2_decap_8 FILLER_48_445 ();
 sg13g2_fill_1 FILLER_48_452 ();
 sg13g2_fill_2 FILLER_48_458 ();
 sg13g2_fill_1 FILLER_48_460 ();
 sg13g2_fill_2 FILLER_48_469 ();
 sg13g2_fill_2 FILLER_48_476 ();
 sg13g2_fill_2 FILLER_48_482 ();
 sg13g2_fill_1 FILLER_48_484 ();
 sg13g2_fill_1 FILLER_48_536 ();
 sg13g2_fill_2 FILLER_48_553 ();
 sg13g2_fill_2 FILLER_48_563 ();
 sg13g2_fill_1 FILLER_48_565 ();
 sg13g2_fill_2 FILLER_48_574 ();
 sg13g2_fill_1 FILLER_48_576 ();
 sg13g2_fill_2 FILLER_48_634 ();
 sg13g2_fill_1 FILLER_48_636 ();
 sg13g2_fill_2 FILLER_48_642 ();
 sg13g2_decap_4 FILLER_48_652 ();
 sg13g2_fill_1 FILLER_48_656 ();
 sg13g2_fill_1 FILLER_48_670 ();
 sg13g2_fill_1 FILLER_48_676 ();
 sg13g2_fill_1 FILLER_48_684 ();
 sg13g2_fill_1 FILLER_48_693 ();
 sg13g2_fill_2 FILLER_48_702 ();
 sg13g2_fill_1 FILLER_48_728 ();
 sg13g2_decap_4 FILLER_48_737 ();
 sg13g2_fill_2 FILLER_48_741 ();
 sg13g2_fill_1 FILLER_48_754 ();
 sg13g2_decap_4 FILLER_48_787 ();
 sg13g2_fill_2 FILLER_48_791 ();
 sg13g2_fill_1 FILLER_48_801 ();
 sg13g2_decap_4 FILLER_48_807 ();
 sg13g2_fill_1 FILLER_48_811 ();
 sg13g2_decap_8 FILLER_48_837 ();
 sg13g2_decap_8 FILLER_48_844 ();
 sg13g2_decap_8 FILLER_48_851 ();
 sg13g2_decap_8 FILLER_48_858 ();
 sg13g2_decap_8 FILLER_48_865 ();
 sg13g2_decap_4 FILLER_48_872 ();
 sg13g2_fill_2 FILLER_48_876 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_4 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_118 ();
 sg13g2_fill_1 FILLER_49_135 ();
 sg13g2_fill_1 FILLER_49_142 ();
 sg13g2_fill_1 FILLER_49_179 ();
 sg13g2_fill_1 FILLER_49_194 ();
 sg13g2_fill_2 FILLER_49_270 ();
 sg13g2_fill_1 FILLER_49_329 ();
 sg13g2_fill_2 FILLER_49_334 ();
 sg13g2_fill_1 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_341 ();
 sg13g2_fill_1 FILLER_49_348 ();
 sg13g2_fill_1 FILLER_49_356 ();
 sg13g2_fill_2 FILLER_49_392 ();
 sg13g2_fill_1 FILLER_49_410 ();
 sg13g2_decap_4 FILLER_49_418 ();
 sg13g2_fill_2 FILLER_49_422 ();
 sg13g2_fill_1 FILLER_49_444 ();
 sg13g2_fill_1 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_507 ();
 sg13g2_fill_1 FILLER_49_514 ();
 sg13g2_decap_4 FILLER_49_575 ();
 sg13g2_fill_1 FILLER_49_591 ();
 sg13g2_fill_2 FILLER_49_623 ();
 sg13g2_fill_2 FILLER_49_641 ();
 sg13g2_fill_1 FILLER_49_643 ();
 sg13g2_fill_2 FILLER_49_652 ();
 sg13g2_fill_1 FILLER_49_654 ();
 sg13g2_decap_8 FILLER_49_671 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_fill_2 FILLER_49_726 ();
 sg13g2_fill_1 FILLER_49_728 ();
 sg13g2_decap_4 FILLER_49_736 ();
 sg13g2_fill_2 FILLER_49_740 ();
 sg13g2_fill_1 FILLER_49_746 ();
 sg13g2_fill_2 FILLER_49_769 ();
 sg13g2_decap_4 FILLER_49_774 ();
 sg13g2_decap_8 FILLER_49_783 ();
 sg13g2_fill_2 FILLER_49_790 ();
 sg13g2_fill_1 FILLER_49_808 ();
 sg13g2_fill_2 FILLER_49_822 ();
 sg13g2_decap_8 FILLER_49_836 ();
 sg13g2_decap_8 FILLER_49_843 ();
 sg13g2_decap_8 FILLER_49_850 ();
 sg13g2_decap_8 FILLER_49_857 ();
 sg13g2_decap_8 FILLER_49_864 ();
 sg13g2_decap_8 FILLER_49_871 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_fill_2 FILLER_50_56 ();
 sg13g2_fill_1 FILLER_50_84 ();
 sg13g2_fill_1 FILLER_50_111 ();
 sg13g2_fill_2 FILLER_50_138 ();
 sg13g2_fill_2 FILLER_50_166 ();
 sg13g2_fill_1 FILLER_50_194 ();
 sg13g2_fill_2 FILLER_50_244 ();
 sg13g2_fill_1 FILLER_50_255 ();
 sg13g2_decap_4 FILLER_50_268 ();
 sg13g2_fill_2 FILLER_50_272 ();
 sg13g2_decap_4 FILLER_50_282 ();
 sg13g2_fill_2 FILLER_50_286 ();
 sg13g2_decap_4 FILLER_50_292 ();
 sg13g2_fill_1 FILLER_50_296 ();
 sg13g2_decap_4 FILLER_50_313 ();
 sg13g2_fill_1 FILLER_50_400 ();
 sg13g2_fill_1 FILLER_50_405 ();
 sg13g2_fill_1 FILLER_50_411 ();
 sg13g2_fill_1 FILLER_50_416 ();
 sg13g2_fill_2 FILLER_50_427 ();
 sg13g2_decap_4 FILLER_50_442 ();
 sg13g2_fill_1 FILLER_50_446 ();
 sg13g2_fill_2 FILLER_50_452 ();
 sg13g2_fill_2 FILLER_50_480 ();
 sg13g2_fill_1 FILLER_50_496 ();
 sg13g2_fill_1 FILLER_50_502 ();
 sg13g2_fill_2 FILLER_50_529 ();
 sg13g2_fill_1 FILLER_50_536 ();
 sg13g2_fill_2 FILLER_50_545 ();
 sg13g2_fill_2 FILLER_50_591 ();
 sg13g2_fill_1 FILLER_50_605 ();
 sg13g2_decap_8 FILLER_50_610 ();
 sg13g2_fill_2 FILLER_50_617 ();
 sg13g2_fill_1 FILLER_50_619 ();
 sg13g2_fill_2 FILLER_50_624 ();
 sg13g2_fill_1 FILLER_50_664 ();
 sg13g2_fill_1 FILLER_50_701 ();
 sg13g2_fill_1 FILLER_50_714 ();
 sg13g2_fill_2 FILLER_50_719 ();
 sg13g2_fill_2 FILLER_50_726 ();
 sg13g2_decap_4 FILLER_50_736 ();
 sg13g2_fill_1 FILLER_50_752 ();
 sg13g2_fill_2 FILLER_50_760 ();
 sg13g2_fill_2 FILLER_50_772 ();
 sg13g2_decap_4 FILLER_50_787 ();
 sg13g2_fill_1 FILLER_50_838 ();
 sg13g2_fill_2 FILLER_50_843 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_8 FILLER_50_856 ();
 sg13g2_decap_8 FILLER_50_863 ();
 sg13g2_decap_8 FILLER_50_870 ();
 sg13g2_fill_1 FILLER_50_877 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_4 FILLER_51_49 ();
 sg13g2_fill_2 FILLER_51_53 ();
 sg13g2_fill_1 FILLER_51_111 ();
 sg13g2_fill_1 FILLER_51_162 ();
 sg13g2_fill_1 FILLER_51_184 ();
 sg13g2_fill_1 FILLER_51_225 ();
 sg13g2_fill_2 FILLER_51_256 ();
 sg13g2_fill_1 FILLER_51_284 ();
 sg13g2_fill_2 FILLER_51_311 ();
 sg13g2_fill_2 FILLER_51_317 ();
 sg13g2_fill_2 FILLER_51_327 ();
 sg13g2_fill_2 FILLER_51_333 ();
 sg13g2_fill_1 FILLER_51_335 ();
 sg13g2_fill_1 FILLER_51_345 ();
 sg13g2_fill_1 FILLER_51_364 ();
 sg13g2_fill_2 FILLER_51_371 ();
 sg13g2_fill_1 FILLER_51_399 ();
 sg13g2_fill_1 FILLER_51_404 ();
 sg13g2_fill_1 FILLER_51_409 ();
 sg13g2_fill_2 FILLER_51_415 ();
 sg13g2_fill_2 FILLER_51_446 ();
 sg13g2_decap_4 FILLER_51_467 ();
 sg13g2_fill_1 FILLER_51_471 ();
 sg13g2_fill_1 FILLER_51_498 ();
 sg13g2_fill_1 FILLER_51_504 ();
 sg13g2_fill_1 FILLER_51_509 ();
 sg13g2_fill_1 FILLER_51_536 ();
 sg13g2_fill_2 FILLER_51_601 ();
 sg13g2_fill_2 FILLER_51_629 ();
 sg13g2_fill_1 FILLER_51_631 ();
 sg13g2_fill_1 FILLER_51_675 ();
 sg13g2_decap_4 FILLER_51_680 ();
 sg13g2_decap_8 FILLER_51_717 ();
 sg13g2_fill_1 FILLER_51_724 ();
 sg13g2_fill_2 FILLER_51_746 ();
 sg13g2_fill_2 FILLER_51_752 ();
 sg13g2_fill_1 FILLER_51_754 ();
 sg13g2_decap_4 FILLER_51_769 ();
 sg13g2_fill_2 FILLER_51_773 ();
 sg13g2_fill_1 FILLER_51_808 ();
 sg13g2_decap_4 FILLER_51_817 ();
 sg13g2_fill_1 FILLER_51_821 ();
 sg13g2_fill_2 FILLER_51_843 ();
 sg13g2_fill_1 FILLER_51_845 ();
 sg13g2_decap_8 FILLER_51_851 ();
 sg13g2_decap_8 FILLER_51_858 ();
 sg13g2_decap_8 FILLER_51_865 ();
 sg13g2_decap_4 FILLER_51_872 ();
 sg13g2_fill_2 FILLER_51_876 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_fill_2 FILLER_52_53 ();
 sg13g2_fill_1 FILLER_52_63 ();
 sg13g2_fill_1 FILLER_52_78 ();
 sg13g2_fill_1 FILLER_52_83 ();
 sg13g2_fill_2 FILLER_52_120 ();
 sg13g2_fill_1 FILLER_52_122 ();
 sg13g2_fill_1 FILLER_52_195 ();
 sg13g2_fill_1 FILLER_52_202 ();
 sg13g2_fill_2 FILLER_52_213 ();
 sg13g2_fill_2 FILLER_52_246 ();
 sg13g2_fill_1 FILLER_52_253 ();
 sg13g2_fill_2 FILLER_52_284 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_fill_1 FILLER_52_314 ();
 sg13g2_fill_1 FILLER_52_326 ();
 sg13g2_fill_1 FILLER_52_332 ();
 sg13g2_fill_2 FILLER_52_341 ();
 sg13g2_fill_1 FILLER_52_343 ();
 sg13g2_fill_1 FILLER_52_389 ();
 sg13g2_fill_1 FILLER_52_394 ();
 sg13g2_fill_1 FILLER_52_400 ();
 sg13g2_fill_1 FILLER_52_410 ();
 sg13g2_fill_1 FILLER_52_415 ();
 sg13g2_fill_2 FILLER_52_421 ();
 sg13g2_decap_4 FILLER_52_442 ();
 sg13g2_fill_2 FILLER_52_490 ();
 sg13g2_fill_2 FILLER_52_506 ();
 sg13g2_fill_1 FILLER_52_508 ();
 sg13g2_fill_1 FILLER_52_534 ();
 sg13g2_fill_2 FILLER_52_590 ();
 sg13g2_decap_4 FILLER_52_600 ();
 sg13g2_decap_4 FILLER_52_618 ();
 sg13g2_fill_2 FILLER_52_663 ();
 sg13g2_fill_1 FILLER_52_665 ();
 sg13g2_fill_2 FILLER_52_691 ();
 sg13g2_fill_2 FILLER_52_733 ();
 sg13g2_decap_8 FILLER_52_764 ();
 sg13g2_fill_1 FILLER_52_771 ();
 sg13g2_decap_4 FILLER_52_816 ();
 sg13g2_fill_1 FILLER_52_820 ();
 sg13g2_decap_8 FILLER_52_849 ();
 sg13g2_decap_8 FILLER_52_856 ();
 sg13g2_decap_8 FILLER_52_863 ();
 sg13g2_decap_8 FILLER_52_870 ();
 sg13g2_fill_1 FILLER_52_877 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_98 ();
 sg13g2_fill_1 FILLER_53_106 ();
 sg13g2_fill_1 FILLER_53_137 ();
 sg13g2_fill_1 FILLER_53_159 ();
 sg13g2_fill_2 FILLER_53_168 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_fill_2 FILLER_53_231 ();
 sg13g2_fill_1 FILLER_53_255 ();
 sg13g2_fill_1 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_272 ();
 sg13g2_fill_1 FILLER_53_294 ();
 sg13g2_fill_2 FILLER_53_333 ();
 sg13g2_fill_2 FILLER_53_423 ();
 sg13g2_fill_1 FILLER_53_444 ();
 sg13g2_fill_2 FILLER_53_491 ();
 sg13g2_fill_2 FILLER_53_647 ();
 sg13g2_fill_1 FILLER_53_679 ();
 sg13g2_decap_8 FILLER_53_685 ();
 sg13g2_fill_2 FILLER_53_692 ();
 sg13g2_fill_1 FILLER_53_714 ();
 sg13g2_fill_1 FILLER_53_725 ();
 sg13g2_fill_1 FILLER_53_813 ();
 sg13g2_decap_4 FILLER_53_819 ();
 sg13g2_fill_2 FILLER_53_828 ();
 sg13g2_decap_8 FILLER_53_834 ();
 sg13g2_decap_8 FILLER_53_841 ();
 sg13g2_fill_1 FILLER_53_848 ();
 sg13g2_decap_8 FILLER_53_852 ();
 sg13g2_decap_8 FILLER_53_859 ();
 sg13g2_decap_8 FILLER_53_866 ();
 sg13g2_decap_4 FILLER_53_873 ();
 sg13g2_fill_1 FILLER_53_877 ();
 sg13g2_decap_8 FILLER_54_26 ();
 sg13g2_decap_4 FILLER_54_33 ();
 sg13g2_fill_2 FILLER_54_37 ();
 sg13g2_fill_2 FILLER_54_65 ();
 sg13g2_fill_2 FILLER_54_77 ();
 sg13g2_fill_1 FILLER_54_103 ();
 sg13g2_fill_2 FILLER_54_128 ();
 sg13g2_fill_2 FILLER_54_156 ();
 sg13g2_fill_1 FILLER_54_194 ();
 sg13g2_decap_4 FILLER_54_199 ();
 sg13g2_fill_2 FILLER_54_248 ();
 sg13g2_fill_1 FILLER_54_284 ();
 sg13g2_fill_1 FILLER_54_299 ();
 sg13g2_fill_1 FILLER_54_304 ();
 sg13g2_fill_1 FILLER_54_313 ();
 sg13g2_fill_1 FILLER_54_319 ();
 sg13g2_fill_2 FILLER_54_325 ();
 sg13g2_fill_2 FILLER_54_340 ();
 sg13g2_fill_1 FILLER_54_346 ();
 sg13g2_fill_1 FILLER_54_357 ();
 sg13g2_fill_1 FILLER_54_363 ();
 sg13g2_fill_1 FILLER_54_368 ();
 sg13g2_fill_1 FILLER_54_405 ();
 sg13g2_fill_1 FILLER_54_411 ();
 sg13g2_fill_1 FILLER_54_417 ();
 sg13g2_fill_1 FILLER_54_423 ();
 sg13g2_fill_1 FILLER_54_428 ();
 sg13g2_fill_2 FILLER_54_486 ();
 sg13g2_fill_2 FILLER_54_494 ();
 sg13g2_fill_1 FILLER_54_496 ();
 sg13g2_fill_2 FILLER_54_507 ();
 sg13g2_fill_1 FILLER_54_509 ();
 sg13g2_fill_2 FILLER_54_514 ();
 sg13g2_fill_1 FILLER_54_516 ();
 sg13g2_fill_1 FILLER_54_543 ();
 sg13g2_fill_2 FILLER_54_553 ();
 sg13g2_fill_1 FILLER_54_598 ();
 sg13g2_fill_1 FILLER_54_608 ();
 sg13g2_fill_2 FILLER_54_622 ();
 sg13g2_fill_2 FILLER_54_645 ();
 sg13g2_fill_2 FILLER_54_693 ();
 sg13g2_fill_2 FILLER_54_734 ();
 sg13g2_decap_4 FILLER_54_775 ();
 sg13g2_decap_8 FILLER_54_787 ();
 sg13g2_fill_2 FILLER_54_794 ();
 sg13g2_fill_2 FILLER_54_821 ();
 sg13g2_fill_1 FILLER_54_823 ();
 sg13g2_decap_8 FILLER_54_857 ();
 sg13g2_decap_8 FILLER_54_864 ();
 sg13g2_decap_8 FILLER_54_871 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_11 ();
 sg13g2_fill_1 FILLER_55_18 ();
 sg13g2_fill_1 FILLER_55_45 ();
 sg13g2_decap_4 FILLER_55_80 ();
 sg13g2_fill_2 FILLER_55_121 ();
 sg13g2_decap_4 FILLER_55_149 ();
 sg13g2_fill_1 FILLER_55_167 ();
 sg13g2_fill_2 FILLER_55_194 ();
 sg13g2_fill_1 FILLER_55_315 ();
 sg13g2_fill_1 FILLER_55_320 ();
 sg13g2_fill_2 FILLER_55_334 ();
 sg13g2_fill_2 FILLER_55_366 ();
 sg13g2_fill_1 FILLER_55_404 ();
 sg13g2_fill_1 FILLER_55_409 ();
 sg13g2_fill_1 FILLER_55_418 ();
 sg13g2_fill_1 FILLER_55_459 ();
 sg13g2_fill_2 FILLER_55_474 ();
 sg13g2_fill_2 FILLER_55_489 ();
 sg13g2_decap_4 FILLER_55_495 ();
 sg13g2_fill_2 FILLER_55_499 ();
 sg13g2_fill_1 FILLER_55_531 ();
 sg13g2_fill_2 FILLER_55_536 ();
 sg13g2_fill_1 FILLER_55_538 ();
 sg13g2_fill_2 FILLER_55_543 ();
 sg13g2_fill_1 FILLER_55_545 ();
 sg13g2_fill_2 FILLER_55_572 ();
 sg13g2_fill_1 FILLER_55_574 ();
 sg13g2_fill_2 FILLER_55_584 ();
 sg13g2_fill_1 FILLER_55_594 ();
 sg13g2_fill_1 FILLER_55_603 ();
 sg13g2_fill_1 FILLER_55_613 ();
 sg13g2_fill_1 FILLER_55_652 ();
 sg13g2_fill_2 FILLER_55_724 ();
 sg13g2_decap_8 FILLER_55_751 ();
 sg13g2_decap_4 FILLER_55_758 ();
 sg13g2_fill_1 FILLER_55_762 ();
 sg13g2_decap_8 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_791 ();
 sg13g2_fill_2 FILLER_55_851 ();
 sg13g2_decap_8 FILLER_55_859 ();
 sg13g2_decap_8 FILLER_55_866 ();
 sg13g2_decap_4 FILLER_55_873 ();
 sg13g2_fill_1 FILLER_55_877 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_4 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_fill_2 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_58 ();
 sg13g2_fill_2 FILLER_56_88 ();
 sg13g2_fill_1 FILLER_56_116 ();
 sg13g2_fill_2 FILLER_56_174 ();
 sg13g2_fill_1 FILLER_56_176 ();
 sg13g2_decap_4 FILLER_56_217 ();
 sg13g2_fill_1 FILLER_56_221 ();
 sg13g2_fill_1 FILLER_56_241 ();
 sg13g2_fill_2 FILLER_56_278 ();
 sg13g2_decap_4 FILLER_56_297 ();
 sg13g2_fill_1 FILLER_56_301 ();
 sg13g2_fill_2 FILLER_56_328 ();
 sg13g2_fill_1 FILLER_56_355 ();
 sg13g2_fill_2 FILLER_56_435 ();
 sg13g2_fill_1 FILLER_56_449 ();
 sg13g2_fill_2 FILLER_56_484 ();
 sg13g2_fill_1 FILLER_56_491 ();
 sg13g2_fill_2 FILLER_56_504 ();
 sg13g2_fill_1 FILLER_56_506 ();
 sg13g2_fill_2 FILLER_56_511 ();
 sg13g2_fill_2 FILLER_56_523 ();
 sg13g2_decap_4 FILLER_56_530 ();
 sg13g2_fill_1 FILLER_56_557 ();
 sg13g2_fill_1 FILLER_56_584 ();
 sg13g2_fill_2 FILLER_56_633 ();
 sg13g2_fill_1 FILLER_56_635 ();
 sg13g2_fill_2 FILLER_56_653 ();
 sg13g2_fill_1 FILLER_56_671 ();
 sg13g2_fill_2 FILLER_56_676 ();
 sg13g2_fill_1 FILLER_56_678 ();
 sg13g2_fill_2 FILLER_56_684 ();
 sg13g2_decap_8 FILLER_56_690 ();
 sg13g2_fill_2 FILLER_56_697 ();
 sg13g2_fill_1 FILLER_56_731 ();
 sg13g2_fill_2 FILLER_56_758 ();
 sg13g2_fill_1 FILLER_56_760 ();
 sg13g2_fill_1 FILLER_56_770 ();
 sg13g2_decap_8 FILLER_56_778 ();
 sg13g2_fill_2 FILLER_56_795 ();
 sg13g2_fill_1 FILLER_56_797 ();
 sg13g2_decap_4 FILLER_56_808 ();
 sg13g2_fill_1 FILLER_56_817 ();
 sg13g2_fill_1 FILLER_56_822 ();
 sg13g2_fill_1 FILLER_56_827 ();
 sg13g2_fill_1 FILLER_56_831 ();
 sg13g2_fill_1 FILLER_56_838 ();
 sg13g2_fill_1 FILLER_56_842 ();
 sg13g2_fill_2 FILLER_56_848 ();
 sg13g2_decap_8 FILLER_56_856 ();
 sg13g2_decap_8 FILLER_56_863 ();
 sg13g2_decap_8 FILLER_56_870 ();
 sg13g2_fill_1 FILLER_56_877 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_38 ();
 sg13g2_fill_1 FILLER_57_87 ();
 sg13g2_fill_1 FILLER_57_102 ();
 sg13g2_fill_1 FILLER_57_108 ();
 sg13g2_fill_2 FILLER_57_139 ();
 sg13g2_fill_2 FILLER_57_145 ();
 sg13g2_fill_2 FILLER_57_188 ();
 sg13g2_fill_2 FILLER_57_224 ();
 sg13g2_fill_1 FILLER_57_226 ();
 sg13g2_fill_2 FILLER_57_265 ();
 sg13g2_fill_1 FILLER_57_267 ();
 sg13g2_fill_2 FILLER_57_286 ();
 sg13g2_fill_2 FILLER_57_297 ();
 sg13g2_fill_2 FILLER_57_320 ();
 sg13g2_fill_2 FILLER_57_339 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_fill_1 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_368 ();
 sg13g2_fill_1 FILLER_57_394 ();
 sg13g2_fill_1 FILLER_57_435 ();
 sg13g2_fill_1 FILLER_57_451 ();
 sg13g2_fill_1 FILLER_57_468 ();
 sg13g2_fill_2 FILLER_57_490 ();
 sg13g2_fill_1 FILLER_57_571 ();
 sg13g2_decap_4 FILLER_57_582 ();
 sg13g2_fill_2 FILLER_57_586 ();
 sg13g2_fill_2 FILLER_57_619 ();
 sg13g2_decap_4 FILLER_57_626 ();
 sg13g2_fill_1 FILLER_57_630 ();
 sg13g2_fill_1 FILLER_57_653 ();
 sg13g2_fill_1 FILLER_57_688 ();
 sg13g2_fill_2 FILLER_57_750 ();
 sg13g2_fill_1 FILLER_57_782 ();
 sg13g2_decap_4 FILLER_57_813 ();
 sg13g2_fill_2 FILLER_57_817 ();
 sg13g2_decap_8 FILLER_57_850 ();
 sg13g2_decap_8 FILLER_57_857 ();
 sg13g2_decap_8 FILLER_57_864 ();
 sg13g2_decap_8 FILLER_57_871 ();
 sg13g2_fill_1 FILLER_58_26 ();
 sg13g2_fill_2 FILLER_58_84 ();
 sg13g2_fill_1 FILLER_58_86 ();
 sg13g2_fill_2 FILLER_58_117 ();
 sg13g2_decap_8 FILLER_58_155 ();
 sg13g2_fill_2 FILLER_58_162 ();
 sg13g2_fill_1 FILLER_58_164 ();
 sg13g2_fill_2 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_224 ();
 sg13g2_fill_2 FILLER_58_231 ();
 sg13g2_fill_2 FILLER_58_304 ();
 sg13g2_fill_1 FILLER_58_306 ();
 sg13g2_fill_1 FILLER_58_336 ();
 sg13g2_fill_1 FILLER_58_358 ();
 sg13g2_fill_2 FILLER_58_365 ();
 sg13g2_fill_1 FILLER_58_388 ();
 sg13g2_fill_1 FILLER_58_393 ();
 sg13g2_fill_1 FILLER_58_404 ();
 sg13g2_fill_2 FILLER_58_412 ();
 sg13g2_fill_2 FILLER_58_424 ();
 sg13g2_fill_1 FILLER_58_431 ();
 sg13g2_fill_1 FILLER_58_437 ();
 sg13g2_fill_1 FILLER_58_443 ();
 sg13g2_fill_1 FILLER_58_448 ();
 sg13g2_fill_2 FILLER_58_453 ();
 sg13g2_fill_1 FILLER_58_474 ();
 sg13g2_fill_1 FILLER_58_480 ();
 sg13g2_fill_1 FILLER_58_487 ();
 sg13g2_fill_2 FILLER_58_498 ();
 sg13g2_fill_1 FILLER_58_504 ();
 sg13g2_fill_1 FILLER_58_515 ();
 sg13g2_fill_2 FILLER_58_546 ();
 sg13g2_decap_8 FILLER_58_574 ();
 sg13g2_fill_2 FILLER_58_581 ();
 sg13g2_fill_1 FILLER_58_583 ();
 sg13g2_decap_8 FILLER_58_600 ();
 sg13g2_decap_4 FILLER_58_607 ();
 sg13g2_fill_1 FILLER_58_615 ();
 sg13g2_fill_2 FILLER_58_642 ();
 sg13g2_fill_2 FILLER_58_664 ();
 sg13g2_fill_1 FILLER_58_692 ();
 sg13g2_fill_1 FILLER_58_706 ();
 sg13g2_fill_1 FILLER_58_760 ();
 sg13g2_fill_1 FILLER_58_772 ();
 sg13g2_fill_1 FILLER_58_780 ();
 sg13g2_fill_1 FILLER_58_786 ();
 sg13g2_fill_2 FILLER_58_798 ();
 sg13g2_fill_1 FILLER_58_800 ();
 sg13g2_decap_4 FILLER_58_805 ();
 sg13g2_decap_8 FILLER_58_840 ();
 sg13g2_decap_8 FILLER_58_847 ();
 sg13g2_decap_8 FILLER_58_854 ();
 sg13g2_decap_8 FILLER_58_861 ();
 sg13g2_decap_8 FILLER_58_868 ();
 sg13g2_fill_2 FILLER_58_875 ();
 sg13g2_fill_1 FILLER_58_877 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_8 ();
 sg13g2_fill_2 FILLER_59_14 ();
 sg13g2_fill_1 FILLER_59_16 ();
 sg13g2_fill_2 FILLER_59_27 ();
 sg13g2_fill_1 FILLER_59_29 ();
 sg13g2_fill_2 FILLER_59_40 ();
 sg13g2_fill_1 FILLER_59_70 ();
 sg13g2_fill_2 FILLER_59_77 ();
 sg13g2_fill_1 FILLER_59_95 ();
 sg13g2_fill_2 FILLER_59_130 ();
 sg13g2_fill_1 FILLER_59_136 ();
 sg13g2_fill_1 FILLER_59_158 ();
 sg13g2_fill_2 FILLER_59_203 ();
 sg13g2_fill_2 FILLER_59_217 ();
 sg13g2_fill_2 FILLER_59_260 ();
 sg13g2_fill_1 FILLER_59_262 ();
 sg13g2_fill_2 FILLER_59_267 ();
 sg13g2_fill_2 FILLER_59_302 ();
 sg13g2_fill_1 FILLER_59_304 ();
 sg13g2_decap_8 FILLER_59_326 ();
 sg13g2_decap_8 FILLER_59_337 ();
 sg13g2_fill_2 FILLER_59_344 ();
 sg13g2_fill_1 FILLER_59_346 ();
 sg13g2_fill_2 FILLER_59_368 ();
 sg13g2_fill_2 FILLER_59_391 ();
 sg13g2_fill_1 FILLER_59_414 ();
 sg13g2_fill_1 FILLER_59_419 ();
 sg13g2_fill_1 FILLER_59_446 ();
 sg13g2_fill_1 FILLER_59_452 ();
 sg13g2_fill_1 FILLER_59_487 ();
 sg13g2_fill_1 FILLER_59_530 ();
 sg13g2_fill_2 FILLER_59_541 ();
 sg13g2_decap_4 FILLER_59_552 ();
 sg13g2_fill_2 FILLER_59_574 ();
 sg13g2_fill_2 FILLER_59_580 ();
 sg13g2_fill_1 FILLER_59_619 ();
 sg13g2_fill_2 FILLER_59_625 ();
 sg13g2_fill_2 FILLER_59_632 ();
 sg13g2_fill_1 FILLER_59_652 ();
 sg13g2_fill_2 FILLER_59_682 ();
 sg13g2_fill_1 FILLER_59_710 ();
 sg13g2_fill_2 FILLER_59_719 ();
 sg13g2_fill_2 FILLER_59_763 ();
 sg13g2_decap_4 FILLER_59_781 ();
 sg13g2_fill_2 FILLER_59_785 ();
 sg13g2_decap_8 FILLER_59_800 ();
 sg13g2_fill_2 FILLER_59_807 ();
 sg13g2_fill_1 FILLER_59_809 ();
 sg13g2_fill_1 FILLER_59_814 ();
 sg13g2_fill_1 FILLER_59_819 ();
 sg13g2_decap_8 FILLER_59_824 ();
 sg13g2_decap_8 FILLER_59_831 ();
 sg13g2_decap_8 FILLER_59_838 ();
 sg13g2_decap_8 FILLER_59_845 ();
 sg13g2_decap_8 FILLER_59_852 ();
 sg13g2_decap_8 FILLER_59_859 ();
 sg13g2_decap_8 FILLER_59_866 ();
 sg13g2_decap_4 FILLER_59_873 ();
 sg13g2_fill_1 FILLER_59_877 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_28 ();
 sg13g2_fill_1 FILLER_60_30 ();
 sg13g2_fill_2 FILLER_60_65 ();
 sg13g2_fill_2 FILLER_60_79 ();
 sg13g2_fill_1 FILLER_60_183 ();
 sg13g2_fill_1 FILLER_60_224 ();
 sg13g2_fill_2 FILLER_60_238 ();
 sg13g2_fill_1 FILLER_60_240 ();
 sg13g2_fill_2 FILLER_60_246 ();
 sg13g2_fill_1 FILLER_60_272 ();
 sg13g2_fill_1 FILLER_60_281 ();
 sg13g2_fill_1 FILLER_60_291 ();
 sg13g2_fill_1 FILLER_60_297 ();
 sg13g2_fill_1 FILLER_60_361 ();
 sg13g2_fill_2 FILLER_60_395 ();
 sg13g2_fill_2 FILLER_60_418 ();
 sg13g2_fill_2 FILLER_60_425 ();
 sg13g2_fill_2 FILLER_60_464 ();
 sg13g2_decap_4 FILLER_60_470 ();
 sg13g2_fill_1 FILLER_60_474 ();
 sg13g2_fill_1 FILLER_60_480 ();
 sg13g2_fill_2 FILLER_60_486 ();
 sg13g2_fill_2 FILLER_60_509 ();
 sg13g2_fill_2 FILLER_60_532 ();
 sg13g2_fill_1 FILLER_60_534 ();
 sg13g2_fill_2 FILLER_60_556 ();
 sg13g2_fill_1 FILLER_60_573 ();
 sg13g2_fill_2 FILLER_60_578 ();
 sg13g2_fill_1 FILLER_60_580 ();
 sg13g2_fill_2 FILLER_60_584 ();
 sg13g2_decap_8 FILLER_60_617 ();
 sg13g2_decap_4 FILLER_60_624 ();
 sg13g2_fill_1 FILLER_60_637 ();
 sg13g2_fill_1 FILLER_60_668 ();
 sg13g2_fill_2 FILLER_60_678 ();
 sg13g2_decap_4 FILLER_60_688 ();
 sg13g2_fill_2 FILLER_60_696 ();
 sg13g2_fill_1 FILLER_60_706 ();
 sg13g2_decap_4 FILLER_60_753 ();
 sg13g2_decap_4 FILLER_60_761 ();
 sg13g2_decap_8 FILLER_60_774 ();
 sg13g2_decap_4 FILLER_60_781 ();
 sg13g2_fill_1 FILLER_60_785 ();
 sg13g2_fill_2 FILLER_60_815 ();
 sg13g2_decap_8 FILLER_60_822 ();
 sg13g2_fill_1 FILLER_60_829 ();
 sg13g2_decap_8 FILLER_60_838 ();
 sg13g2_decap_8 FILLER_60_845 ();
 sg13g2_decap_8 FILLER_60_852 ();
 sg13g2_decap_8 FILLER_60_859 ();
 sg13g2_decap_8 FILLER_60_866 ();
 sg13g2_decap_4 FILLER_60_873 ();
 sg13g2_fill_1 FILLER_60_877 ();
 sg13g2_fill_1 FILLER_61_42 ();
 sg13g2_fill_2 FILLER_61_95 ();
 sg13g2_fill_2 FILLER_61_111 ();
 sg13g2_fill_2 FILLER_61_139 ();
 sg13g2_fill_2 FILLER_61_162 ();
 sg13g2_fill_1 FILLER_61_164 ();
 sg13g2_fill_2 FILLER_61_169 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_fill_2 FILLER_61_177 ();
 sg13g2_fill_1 FILLER_61_179 ();
 sg13g2_fill_1 FILLER_61_201 ();
 sg13g2_fill_1 FILLER_61_223 ();
 sg13g2_fill_1 FILLER_61_238 ();
 sg13g2_fill_1 FILLER_61_271 ();
 sg13g2_fill_2 FILLER_61_279 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_fill_2 FILLER_61_357 ();
 sg13g2_decap_8 FILLER_61_380 ();
 sg13g2_fill_1 FILLER_61_387 ();
 sg13g2_decap_4 FILLER_61_447 ();
 sg13g2_decap_8 FILLER_61_458 ();
 sg13g2_fill_2 FILLER_61_487 ();
 sg13g2_fill_1 FILLER_61_489 ();
 sg13g2_decap_4 FILLER_61_494 ();
 sg13g2_fill_2 FILLER_61_498 ();
 sg13g2_decap_4 FILLER_61_505 ();
 sg13g2_fill_1 FILLER_61_509 ();
 sg13g2_fill_1 FILLER_61_514 ();
 sg13g2_fill_1 FILLER_61_519 ();
 sg13g2_fill_1 FILLER_61_525 ();
 sg13g2_fill_1 FILLER_61_531 ();
 sg13g2_fill_1 FILLER_61_536 ();
 sg13g2_fill_2 FILLER_61_567 ();
 sg13g2_fill_1 FILLER_61_569 ();
 sg13g2_decap_4 FILLER_61_638 ();
 sg13g2_fill_1 FILLER_61_647 ();
 sg13g2_fill_2 FILLER_61_653 ();
 sg13g2_fill_1 FILLER_61_655 ();
 sg13g2_fill_1 FILLER_61_669 ();
 sg13g2_decap_4 FILLER_61_708 ();
 sg13g2_fill_2 FILLER_61_712 ();
 sg13g2_fill_2 FILLER_61_777 ();
 sg13g2_fill_1 FILLER_61_784 ();
 sg13g2_fill_1 FILLER_61_789 ();
 sg13g2_fill_1 FILLER_61_802 ();
 sg13g2_fill_1 FILLER_61_809 ();
 sg13g2_fill_2 FILLER_61_823 ();
 sg13g2_fill_1 FILLER_61_825 ();
 sg13g2_decap_8 FILLER_61_834 ();
 sg13g2_decap_8 FILLER_61_841 ();
 sg13g2_decap_8 FILLER_61_848 ();
 sg13g2_decap_8 FILLER_61_855 ();
 sg13g2_decap_8 FILLER_61_862 ();
 sg13g2_decap_8 FILLER_61_869 ();
 sg13g2_fill_2 FILLER_61_876 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_1 FILLER_62_29 ();
 sg13g2_fill_2 FILLER_62_51 ();
 sg13g2_fill_1 FILLER_62_53 ();
 sg13g2_fill_2 FILLER_62_79 ();
 sg13g2_fill_1 FILLER_62_85 ();
 sg13g2_fill_2 FILLER_62_112 ();
 sg13g2_fill_1 FILLER_62_128 ();
 sg13g2_fill_1 FILLER_62_150 ();
 sg13g2_decap_8 FILLER_62_202 ();
 sg13g2_fill_2 FILLER_62_209 ();
 sg13g2_fill_1 FILLER_62_211 ();
 sg13g2_decap_4 FILLER_62_217 ();
 sg13g2_fill_1 FILLER_62_253 ();
 sg13g2_fill_1 FILLER_62_278 ();
 sg13g2_fill_2 FILLER_62_303 ();
 sg13g2_fill_1 FILLER_62_305 ();
 sg13g2_fill_1 FILLER_62_327 ();
 sg13g2_fill_2 FILLER_62_332 ();
 sg13g2_decap_8 FILLER_62_388 ();
 sg13g2_fill_1 FILLER_62_395 ();
 sg13g2_fill_1 FILLER_62_421 ();
 sg13g2_fill_1 FILLER_62_448 ();
 sg13g2_fill_1 FILLER_62_485 ();
 sg13g2_fill_2 FILLER_62_507 ();
 sg13g2_fill_1 FILLER_62_535 ();
 sg13g2_fill_2 FILLER_62_557 ();
 sg13g2_fill_1 FILLER_62_559 ();
 sg13g2_fill_2 FILLER_62_564 ();
 sg13g2_decap_4 FILLER_62_571 ();
 sg13g2_fill_1 FILLER_62_579 ();
 sg13g2_fill_2 FILLER_62_596 ();
 sg13g2_fill_1 FILLER_62_602 ();
 sg13g2_fill_1 FILLER_62_608 ();
 sg13g2_fill_2 FILLER_62_613 ();
 sg13g2_fill_2 FILLER_62_620 ();
 sg13g2_fill_1 FILLER_62_626 ();
 sg13g2_fill_1 FILLER_62_640 ();
 sg13g2_fill_1 FILLER_62_653 ();
 sg13g2_decap_8 FILLER_62_689 ();
 sg13g2_decap_4 FILLER_62_696 ();
 sg13g2_decap_8 FILLER_62_704 ();
 sg13g2_fill_2 FILLER_62_711 ();
 sg13g2_fill_1 FILLER_62_713 ();
 sg13g2_fill_2 FILLER_62_751 ();
 sg13g2_decap_4 FILLER_62_765 ();
 sg13g2_fill_2 FILLER_62_800 ();
 sg13g2_fill_1 FILLER_62_811 ();
 sg13g2_decap_8 FILLER_62_835 ();
 sg13g2_decap_8 FILLER_62_842 ();
 sg13g2_decap_8 FILLER_62_849 ();
 sg13g2_decap_8 FILLER_62_856 ();
 sg13g2_decap_8 FILLER_62_863 ();
 sg13g2_decap_8 FILLER_62_870 ();
 sg13g2_fill_1 FILLER_62_877 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_27 ();
 sg13g2_fill_2 FILLER_63_38 ();
 sg13g2_fill_2 FILLER_63_66 ();
 sg13g2_fill_2 FILLER_63_94 ();
 sg13g2_fill_1 FILLER_63_96 ();
 sg13g2_decap_4 FILLER_63_101 ();
 sg13g2_fill_2 FILLER_63_131 ();
 sg13g2_fill_1 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_138 ();
 sg13g2_fill_2 FILLER_63_145 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_fill_1 FILLER_63_182 ();
 sg13g2_fill_2 FILLER_63_265 ();
 sg13g2_fill_1 FILLER_63_282 ();
 sg13g2_fill_2 FILLER_63_318 ();
 sg13g2_fill_1 FILLER_63_324 ();
 sg13g2_fill_1 FILLER_63_334 ();
 sg13g2_fill_2 FILLER_63_339 ();
 sg13g2_fill_1 FILLER_63_341 ();
 sg13g2_decap_8 FILLER_63_346 ();
 sg13g2_fill_2 FILLER_63_358 ();
 sg13g2_fill_2 FILLER_63_364 ();
 sg13g2_fill_1 FILLER_63_366 ();
 sg13g2_fill_2 FILLER_63_393 ();
 sg13g2_fill_1 FILLER_63_395 ();
 sg13g2_fill_2 FILLER_63_401 ();
 sg13g2_fill_1 FILLER_63_421 ();
 sg13g2_fill_2 FILLER_63_450 ();
 sg13g2_fill_2 FILLER_63_470 ();
 sg13g2_fill_2 FILLER_63_476 ();
 sg13g2_fill_1 FILLER_63_478 ();
 sg13g2_fill_1 FILLER_63_523 ();
 sg13g2_fill_1 FILLER_63_529 ();
 sg13g2_decap_4 FILLER_63_570 ();
 sg13g2_fill_1 FILLER_63_574 ();
 sg13g2_fill_2 FILLER_63_605 ();
 sg13g2_fill_1 FILLER_63_631 ();
 sg13g2_fill_2 FILLER_63_652 ();
 sg13g2_fill_1 FILLER_63_654 ();
 sg13g2_fill_2 FILLER_63_663 ();
 sg13g2_fill_1 FILLER_63_665 ();
 sg13g2_fill_2 FILLER_63_678 ();
 sg13g2_fill_2 FILLER_63_688 ();
 sg13g2_fill_1 FILLER_63_690 ();
 sg13g2_fill_1 FILLER_63_728 ();
 sg13g2_fill_1 FILLER_63_791 ();
 sg13g2_decap_4 FILLER_63_796 ();
 sg13g2_fill_1 FILLER_63_800 ();
 sg13g2_fill_1 FILLER_63_806 ();
 sg13g2_decap_4 FILLER_63_831 ();
 sg13g2_fill_2 FILLER_63_835 ();
 sg13g2_decap_8 FILLER_63_844 ();
 sg13g2_decap_8 FILLER_63_851 ();
 sg13g2_decap_8 FILLER_63_858 ();
 sg13g2_decap_8 FILLER_63_865 ();
 sg13g2_decap_4 FILLER_63_872 ();
 sg13g2_fill_2 FILLER_63_876 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_2 ();
 sg13g2_fill_2 FILLER_64_39 ();
 sg13g2_fill_1 FILLER_64_41 ();
 sg13g2_fill_2 FILLER_64_52 ();
 sg13g2_fill_1 FILLER_64_54 ();
 sg13g2_fill_2 FILLER_64_91 ();
 sg13g2_decap_4 FILLER_64_97 ();
 sg13g2_fill_2 FILLER_64_101 ();
 sg13g2_fill_2 FILLER_64_153 ();
 sg13g2_fill_2 FILLER_64_219 ();
 sg13g2_fill_2 FILLER_64_268 ();
 sg13g2_decap_4 FILLER_64_302 ();
 sg13g2_fill_2 FILLER_64_328 ();
 sg13g2_fill_2 FILLER_64_343 ();
 sg13g2_decap_4 FILLER_64_371 ();
 sg13g2_decap_8 FILLER_64_383 ();
 sg13g2_decap_4 FILLER_64_390 ();
 sg13g2_fill_1 FILLER_64_394 ();
 sg13g2_fill_1 FILLER_64_449 ();
 sg13g2_decap_4 FILLER_64_493 ();
 sg13g2_fill_2 FILLER_64_533 ();
 sg13g2_fill_1 FILLER_64_535 ();
 sg13g2_fill_1 FILLER_64_569 ();
 sg13g2_fill_2 FILLER_64_627 ();
 sg13g2_fill_1 FILLER_64_629 ();
 sg13g2_fill_1 FILLER_64_655 ();
 sg13g2_fill_2 FILLER_64_674 ();
 sg13g2_decap_4 FILLER_64_790 ();
 sg13g2_fill_2 FILLER_64_806 ();
 sg13g2_decap_8 FILLER_64_853 ();
 sg13g2_decap_8 FILLER_64_860 ();
 sg13g2_decap_8 FILLER_64_867 ();
 sg13g2_decap_4 FILLER_64_874 ();
 sg13g2_fill_1 FILLER_65_4 ();
 sg13g2_fill_2 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_173 ();
 sg13g2_fill_1 FILLER_65_178 ();
 sg13g2_fill_1 FILLER_65_189 ();
 sg13g2_fill_2 FILLER_65_194 ();
 sg13g2_fill_2 FILLER_65_200 ();
 sg13g2_fill_1 FILLER_65_259 ();
 sg13g2_fill_1 FILLER_65_345 ();
 sg13g2_fill_1 FILLER_65_351 ();
 sg13g2_fill_2 FILLER_65_356 ();
 sg13g2_fill_1 FILLER_65_372 ();
 sg13g2_fill_2 FILLER_65_399 ();
 sg13g2_fill_2 FILLER_65_439 ();
 sg13g2_fill_1 FILLER_65_454 ();
 sg13g2_fill_2 FILLER_65_481 ();
 sg13g2_fill_1 FILLER_65_483 ();
 sg13g2_fill_2 FILLER_65_530 ();
 sg13g2_fill_1 FILLER_65_570 ();
 sg13g2_fill_1 FILLER_65_593 ();
 sg13g2_fill_1 FILLER_65_599 ();
 sg13g2_fill_1 FILLER_65_612 ();
 sg13g2_fill_2 FILLER_65_619 ();
 sg13g2_fill_1 FILLER_65_621 ();
 sg13g2_fill_1 FILLER_65_634 ();
 sg13g2_fill_2 FILLER_65_639 ();
 sg13g2_fill_2 FILLER_65_645 ();
 sg13g2_fill_2 FILLER_65_652 ();
 sg13g2_fill_1 FILLER_65_689 ();
 sg13g2_fill_1 FILLER_65_694 ();
 sg13g2_decap_8 FILLER_65_782 ();
 sg13g2_fill_2 FILLER_65_789 ();
 sg13g2_fill_1 FILLER_65_791 ();
 sg13g2_fill_1 FILLER_65_800 ();
 sg13g2_fill_1 FILLER_65_808 ();
 sg13g2_fill_1 FILLER_65_819 ();
 sg13g2_fill_1 FILLER_65_826 ();
 sg13g2_decap_4 FILLER_65_839 ();
 sg13g2_decap_8 FILLER_65_851 ();
 sg13g2_decap_8 FILLER_65_858 ();
 sg13g2_decap_8 FILLER_65_865 ();
 sg13g2_decap_4 FILLER_65_872 ();
 sg13g2_fill_2 FILLER_65_876 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_22 ();
 sg13g2_fill_2 FILLER_66_31 ();
 sg13g2_fill_1 FILLER_66_37 ();
 sg13g2_fill_2 FILLER_66_98 ();
 sg13g2_fill_1 FILLER_66_100 ();
 sg13g2_fill_2 FILLER_66_111 ();
 sg13g2_fill_1 FILLER_66_123 ();
 sg13g2_fill_2 FILLER_66_150 ();
 sg13g2_fill_1 FILLER_66_162 ();
 sg13g2_fill_1 FILLER_66_173 ();
 sg13g2_fill_2 FILLER_66_188 ();
 sg13g2_fill_1 FILLER_66_194 ();
 sg13g2_fill_1 FILLER_66_199 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_fill_2 FILLER_66_266 ();
 sg13g2_fill_1 FILLER_66_278 ();
 sg13g2_fill_1 FILLER_66_305 ();
 sg13g2_fill_1 FILLER_66_320 ();
 sg13g2_fill_1 FILLER_66_325 ();
 sg13g2_fill_2 FILLER_66_331 ();
 sg13g2_fill_1 FILLER_66_369 ();
 sg13g2_fill_1 FILLER_66_411 ();
 sg13g2_fill_1 FILLER_66_417 ();
 sg13g2_fill_1 FILLER_66_439 ();
 sg13g2_fill_1 FILLER_66_449 ();
 sg13g2_decap_4 FILLER_66_455 ();
 sg13g2_fill_1 FILLER_66_474 ();
 sg13g2_fill_2 FILLER_66_487 ();
 sg13g2_fill_1 FILLER_66_493 ();
 sg13g2_fill_1 FILLER_66_504 ();
 sg13g2_fill_1 FILLER_66_531 ();
 sg13g2_fill_2 FILLER_66_563 ();
 sg13g2_decap_4 FILLER_66_601 ();
 sg13g2_fill_1 FILLER_66_605 ();
 sg13g2_fill_1 FILLER_66_710 ();
 sg13g2_fill_2 FILLER_66_741 ();
 sg13g2_fill_2 FILLER_66_756 ();
 sg13g2_decap_4 FILLER_66_765 ();
 sg13g2_fill_1 FILLER_66_769 ();
 sg13g2_fill_1 FILLER_66_778 ();
 sg13g2_fill_1 FILLER_66_783 ();
 sg13g2_fill_1 FILLER_66_801 ();
 sg13g2_fill_2 FILLER_66_810 ();
 sg13g2_fill_1 FILLER_66_816 ();
 sg13g2_fill_2 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_833 ();
 sg13g2_decap_8 FILLER_66_840 ();
 sg13g2_decap_8 FILLER_66_847 ();
 sg13g2_decap_8 FILLER_66_854 ();
 sg13g2_decap_8 FILLER_66_861 ();
 sg13g2_decap_8 FILLER_66_868 ();
 sg13g2_fill_2 FILLER_66_875 ();
 sg13g2_fill_1 FILLER_66_877 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_5 ();
 sg13g2_fill_1 FILLER_67_11 ();
 sg13g2_fill_1 FILLER_67_46 ();
 sg13g2_fill_1 FILLER_67_57 ();
 sg13g2_fill_1 FILLER_67_72 ();
 sg13g2_fill_2 FILLER_67_87 ();
 sg13g2_fill_2 FILLER_67_115 ();
 sg13g2_fill_2 FILLER_67_149 ();
 sg13g2_fill_1 FILLER_67_212 ();
 sg13g2_fill_1 FILLER_67_226 ();
 sg13g2_fill_1 FILLER_67_278 ();
 sg13g2_fill_1 FILLER_67_323 ();
 sg13g2_fill_1 FILLER_67_350 ();
 sg13g2_fill_1 FILLER_67_355 ();
 sg13g2_fill_1 FILLER_67_362 ();
 sg13g2_fill_1 FILLER_67_373 ();
 sg13g2_fill_1 FILLER_67_414 ();
 sg13g2_fill_2 FILLER_67_420 ();
 sg13g2_fill_2 FILLER_67_478 ();
 sg13g2_fill_2 FILLER_67_531 ();
 sg13g2_fill_1 FILLER_67_533 ();
 sg13g2_fill_2 FILLER_67_537 ();
 sg13g2_fill_2 FILLER_67_559 ();
 sg13g2_fill_1 FILLER_67_561 ();
 sg13g2_fill_2 FILLER_67_627 ();
 sg13g2_decap_4 FILLER_67_638 ();
 sg13g2_decap_4 FILLER_67_676 ();
 sg13g2_fill_1 FILLER_67_680 ();
 sg13g2_decap_8 FILLER_67_762 ();
 sg13g2_decap_8 FILLER_67_769 ();
 sg13g2_decap_8 FILLER_67_776 ();
 sg13g2_decap_8 FILLER_67_783 ();
 sg13g2_fill_2 FILLER_67_790 ();
 sg13g2_fill_2 FILLER_67_821 ();
 sg13g2_decap_8 FILLER_67_828 ();
 sg13g2_decap_8 FILLER_67_835 ();
 sg13g2_decap_8 FILLER_67_842 ();
 sg13g2_decap_8 FILLER_67_849 ();
 sg13g2_decap_8 FILLER_67_856 ();
 sg13g2_decap_8 FILLER_67_863 ();
 sg13g2_decap_8 FILLER_67_870 ();
 sg13g2_fill_1 FILLER_67_877 ();
 sg13g2_decap_4 FILLER_68_82 ();
 sg13g2_fill_1 FILLER_68_86 ();
 sg13g2_fill_2 FILLER_68_127 ();
 sg13g2_fill_1 FILLER_68_129 ();
 sg13g2_fill_2 FILLER_68_164 ();
 sg13g2_fill_2 FILLER_68_211 ();
 sg13g2_fill_1 FILLER_68_221 ();
 sg13g2_fill_1 FILLER_68_235 ();
 sg13g2_fill_1 FILLER_68_241 ();
 sg13g2_fill_1 FILLER_68_268 ();
 sg13g2_fill_2 FILLER_68_299 ();
 sg13g2_fill_1 FILLER_68_301 ();
 sg13g2_fill_1 FILLER_68_308 ();
 sg13g2_fill_2 FILLER_68_319 ();
 sg13g2_fill_2 FILLER_68_335 ();
 sg13g2_fill_2 FILLER_68_363 ();
 sg13g2_fill_1 FILLER_68_365 ();
 sg13g2_fill_1 FILLER_68_376 ();
 sg13g2_fill_1 FILLER_68_381 ();
 sg13g2_fill_2 FILLER_68_386 ();
 sg13g2_fill_2 FILLER_68_401 ();
 sg13g2_fill_1 FILLER_68_403 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_fill_1 FILLER_68_422 ();
 sg13g2_fill_1 FILLER_68_427 ();
 sg13g2_fill_2 FILLER_68_434 ();
 sg13g2_fill_1 FILLER_68_459 ();
 sg13g2_fill_2 FILLER_68_489 ();
 sg13g2_fill_2 FILLER_68_501 ();
 sg13g2_fill_1 FILLER_68_548 ();
 sg13g2_fill_2 FILLER_68_634 ();
 sg13g2_fill_1 FILLER_68_649 ();
 sg13g2_fill_2 FILLER_68_676 ();
 sg13g2_fill_1 FILLER_68_686 ();
 sg13g2_fill_2 FILLER_68_695 ();
 sg13g2_fill_2 FILLER_68_705 ();
 sg13g2_fill_1 FILLER_68_727 ();
 sg13g2_decap_8 FILLER_68_762 ();
 sg13g2_decap_8 FILLER_68_769 ();
 sg13g2_decap_8 FILLER_68_776 ();
 sg13g2_decap_8 FILLER_68_783 ();
 sg13g2_decap_8 FILLER_68_790 ();
 sg13g2_decap_8 FILLER_68_797 ();
 sg13g2_decap_8 FILLER_68_804 ();
 sg13g2_decap_8 FILLER_68_811 ();
 sg13g2_decap_8 FILLER_68_818 ();
 sg13g2_decap_8 FILLER_68_825 ();
 sg13g2_decap_8 FILLER_68_832 ();
 sg13g2_decap_8 FILLER_68_839 ();
 sg13g2_decap_8 FILLER_68_846 ();
 sg13g2_decap_8 FILLER_68_853 ();
 sg13g2_decap_8 FILLER_68_860 ();
 sg13g2_decap_8 FILLER_68_867 ();
 sg13g2_decap_4 FILLER_68_874 ();
 sg13g2_fill_1 FILLER_69_36 ();
 sg13g2_fill_2 FILLER_69_91 ();
 sg13g2_fill_2 FILLER_69_196 ();
 sg13g2_fill_2 FILLER_69_203 ();
 sg13g2_fill_1 FILLER_69_223 ();
 sg13g2_fill_2 FILLER_69_239 ();
 sg13g2_fill_2 FILLER_69_250 ();
 sg13g2_fill_2 FILLER_69_265 ();
 sg13g2_fill_1 FILLER_69_267 ();
 sg13g2_fill_1 FILLER_69_278 ();
 sg13g2_fill_1 FILLER_69_284 ();
 sg13g2_fill_2 FILLER_69_294 ();
 sg13g2_fill_1 FILLER_69_301 ();
 sg13g2_fill_1 FILLER_69_316 ();
 sg13g2_fill_1 FILLER_69_343 ();
 sg13g2_fill_2 FILLER_69_348 ();
 sg13g2_fill_2 FILLER_69_354 ();
 sg13g2_fill_1 FILLER_69_356 ();
 sg13g2_decap_4 FILLER_69_362 ();
 sg13g2_fill_1 FILLER_69_396 ();
 sg13g2_fill_1 FILLER_69_402 ();
 sg13g2_fill_1 FILLER_69_411 ();
 sg13g2_fill_1 FILLER_69_417 ();
 sg13g2_fill_2 FILLER_69_423 ();
 sg13g2_fill_1 FILLER_69_449 ();
 sg13g2_fill_2 FILLER_69_453 ();
 sg13g2_fill_2 FILLER_69_485 ();
 sg13g2_fill_1 FILLER_69_518 ();
 sg13g2_fill_1 FILLER_69_575 ();
 sg13g2_fill_2 FILLER_69_581 ();
 sg13g2_fill_1 FILLER_69_588 ();
 sg13g2_fill_2 FILLER_69_593 ();
 sg13g2_fill_2 FILLER_69_599 ();
 sg13g2_fill_1 FILLER_69_601 ();
 sg13g2_fill_2 FILLER_69_606 ();
 sg13g2_fill_1 FILLER_69_608 ();
 sg13g2_fill_2 FILLER_69_613 ();
 sg13g2_decap_8 FILLER_69_622 ();
 sg13g2_decap_4 FILLER_69_629 ();
 sg13g2_fill_1 FILLER_69_633 ();
 sg13g2_fill_1 FILLER_69_656 ();
 sg13g2_fill_2 FILLER_69_699 ();
 sg13g2_fill_2 FILLER_69_706 ();
 sg13g2_fill_1 FILLER_69_708 ();
 sg13g2_decap_8 FILLER_69_747 ();
 sg13g2_decap_8 FILLER_69_754 ();
 sg13g2_decap_8 FILLER_69_761 ();
 sg13g2_decap_8 FILLER_69_768 ();
 sg13g2_decap_8 FILLER_69_775 ();
 sg13g2_decap_8 FILLER_69_782 ();
 sg13g2_decap_8 FILLER_69_789 ();
 sg13g2_decap_8 FILLER_69_796 ();
 sg13g2_decap_8 FILLER_69_803 ();
 sg13g2_decap_8 FILLER_69_810 ();
 sg13g2_decap_8 FILLER_69_817 ();
 sg13g2_decap_8 FILLER_69_824 ();
 sg13g2_decap_8 FILLER_69_831 ();
 sg13g2_decap_8 FILLER_69_838 ();
 sg13g2_decap_8 FILLER_69_845 ();
 sg13g2_decap_8 FILLER_69_852 ();
 sg13g2_decap_8 FILLER_69_859 ();
 sg13g2_decap_8 FILLER_69_866 ();
 sg13g2_decap_4 FILLER_69_873 ();
 sg13g2_fill_1 FILLER_69_877 ();
 sg13g2_fill_2 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_56 ();
 sg13g2_fill_2 FILLER_70_78 ();
 sg13g2_fill_1 FILLER_70_145 ();
 sg13g2_fill_2 FILLER_70_208 ();
 sg13g2_fill_1 FILLER_70_263 ();
 sg13g2_fill_1 FILLER_70_274 ();
 sg13g2_fill_1 FILLER_70_301 ();
 sg13g2_fill_2 FILLER_70_350 ();
 sg13g2_decap_4 FILLER_70_415 ();
 sg13g2_fill_2 FILLER_70_419 ();
 sg13g2_fill_2 FILLER_70_447 ();
 sg13g2_fill_1 FILLER_70_449 ();
 sg13g2_fill_1 FILLER_70_464 ();
 sg13g2_fill_1 FILLER_70_469 ();
 sg13g2_fill_2 FILLER_70_480 ();
 sg13g2_fill_2 FILLER_70_587 ();
 sg13g2_decap_4 FILLER_70_624 ();
 sg13g2_fill_1 FILLER_70_628 ();
 sg13g2_fill_1 FILLER_70_667 ();
 sg13g2_fill_2 FILLER_70_682 ();
 sg13g2_decap_8 FILLER_70_739 ();
 sg13g2_decap_8 FILLER_70_746 ();
 sg13g2_decap_8 FILLER_70_753 ();
 sg13g2_decap_8 FILLER_70_760 ();
 sg13g2_decap_8 FILLER_70_767 ();
 sg13g2_decap_8 FILLER_70_774 ();
 sg13g2_decap_8 FILLER_70_781 ();
 sg13g2_decap_8 FILLER_70_788 ();
 sg13g2_decap_8 FILLER_70_795 ();
 sg13g2_decap_8 FILLER_70_802 ();
 sg13g2_decap_8 FILLER_70_809 ();
 sg13g2_decap_8 FILLER_70_816 ();
 sg13g2_decap_8 FILLER_70_823 ();
 sg13g2_decap_8 FILLER_70_830 ();
 sg13g2_decap_8 FILLER_70_837 ();
 sg13g2_decap_8 FILLER_70_844 ();
 sg13g2_decap_8 FILLER_70_851 ();
 sg13g2_decap_8 FILLER_70_858 ();
 sg13g2_decap_8 FILLER_70_865 ();
 sg13g2_decap_4 FILLER_70_872 ();
 sg13g2_fill_2 FILLER_70_876 ();
 sg13g2_fill_1 FILLER_71_70 ();
 sg13g2_fill_1 FILLER_71_77 ();
 sg13g2_fill_1 FILLER_71_151 ();
 sg13g2_fill_2 FILLER_71_178 ();
 sg13g2_fill_2 FILLER_71_183 ();
 sg13g2_fill_2 FILLER_71_275 ();
 sg13g2_fill_2 FILLER_71_282 ();
 sg13g2_fill_1 FILLER_71_284 ();
 sg13g2_fill_1 FILLER_71_289 ();
 sg13g2_fill_1 FILLER_71_328 ();
 sg13g2_fill_2 FILLER_71_333 ();
 sg13g2_fill_1 FILLER_71_339 ();
 sg13g2_fill_1 FILLER_71_348 ();
 sg13g2_fill_2 FILLER_71_374 ();
 sg13g2_fill_2 FILLER_71_385 ();
 sg13g2_fill_1 FILLER_71_387 ();
 sg13g2_fill_1 FILLER_71_423 ();
 sg13g2_decap_8 FILLER_71_433 ();
 sg13g2_fill_1 FILLER_71_445 ();
 sg13g2_decap_4 FILLER_71_458 ();
 sg13g2_decap_4 FILLER_71_522 ();
 sg13g2_fill_1 FILLER_71_526 ();
 sg13g2_fill_1 FILLER_71_604 ();
 sg13g2_decap_4 FILLER_71_620 ();
 sg13g2_fill_1 FILLER_71_624 ();
 sg13g2_fill_1 FILLER_71_634 ();
 sg13g2_fill_1 FILLER_71_639 ();
 sg13g2_fill_1 FILLER_71_647 ();
 sg13g2_fill_2 FILLER_71_680 ();
 sg13g2_fill_2 FILLER_71_692 ();
 sg13g2_fill_2 FILLER_71_716 ();
 sg13g2_fill_1 FILLER_71_726 ();
 sg13g2_decap_8 FILLER_71_735 ();
 sg13g2_decap_8 FILLER_71_742 ();
 sg13g2_decap_8 FILLER_71_749 ();
 sg13g2_decap_8 FILLER_71_756 ();
 sg13g2_decap_8 FILLER_71_763 ();
 sg13g2_decap_8 FILLER_71_770 ();
 sg13g2_decap_8 FILLER_71_777 ();
 sg13g2_decap_8 FILLER_71_784 ();
 sg13g2_decap_8 FILLER_71_791 ();
 sg13g2_decap_8 FILLER_71_798 ();
 sg13g2_decap_8 FILLER_71_805 ();
 sg13g2_decap_8 FILLER_71_812 ();
 sg13g2_decap_8 FILLER_71_819 ();
 sg13g2_decap_8 FILLER_71_826 ();
 sg13g2_decap_8 FILLER_71_833 ();
 sg13g2_decap_8 FILLER_71_840 ();
 sg13g2_decap_8 FILLER_71_847 ();
 sg13g2_decap_8 FILLER_71_854 ();
 sg13g2_decap_8 FILLER_71_861 ();
 sg13g2_decap_8 FILLER_71_868 ();
 sg13g2_fill_2 FILLER_71_875 ();
 sg13g2_fill_1 FILLER_71_877 ();
 sg13g2_fill_2 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_6 ();
 sg13g2_fill_1 FILLER_72_8 ();
 sg13g2_fill_1 FILLER_72_19 ();
 sg13g2_fill_2 FILLER_72_46 ();
 sg13g2_fill_1 FILLER_72_48 ();
 sg13g2_fill_2 FILLER_72_70 ();
 sg13g2_fill_1 FILLER_72_72 ();
 sg13g2_fill_2 FILLER_72_99 ();
 sg13g2_fill_1 FILLER_72_101 ();
 sg13g2_fill_2 FILLER_72_192 ();
 sg13g2_fill_1 FILLER_72_194 ();
 sg13g2_fill_1 FILLER_72_221 ();
 sg13g2_fill_1 FILLER_72_265 ();
 sg13g2_fill_2 FILLER_72_287 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_fill_1 FILLER_72_365 ();
 sg13g2_fill_2 FILLER_72_410 ();
 sg13g2_fill_1 FILLER_72_417 ();
 sg13g2_fill_1 FILLER_72_423 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_fill_2 FILLER_72_466 ();
 sg13g2_fill_1 FILLER_72_468 ();
 sg13g2_fill_2 FILLER_72_495 ();
 sg13g2_fill_1 FILLER_72_497 ();
 sg13g2_decap_8 FILLER_72_502 ();
 sg13g2_fill_2 FILLER_72_509 ();
 sg13g2_fill_1 FILLER_72_516 ();
 sg13g2_fill_2 FILLER_72_524 ();
 sg13g2_fill_1 FILLER_72_526 ();
 sg13g2_fill_2 FILLER_72_531 ();
 sg13g2_fill_1 FILLER_72_560 ();
 sg13g2_fill_2 FILLER_72_587 ();
 sg13g2_fill_1 FILLER_72_614 ();
 sg13g2_fill_1 FILLER_72_654 ();
 sg13g2_fill_2 FILLER_72_676 ();
 sg13g2_fill_2 FILLER_72_682 ();
 sg13g2_fill_1 FILLER_72_712 ();
 sg13g2_decap_8 FILLER_72_729 ();
 sg13g2_decap_8 FILLER_72_736 ();
 sg13g2_decap_8 FILLER_72_743 ();
 sg13g2_decap_8 FILLER_72_750 ();
 sg13g2_decap_8 FILLER_72_757 ();
 sg13g2_decap_8 FILLER_72_764 ();
 sg13g2_decap_8 FILLER_72_771 ();
 sg13g2_decap_8 FILLER_72_778 ();
 sg13g2_decap_8 FILLER_72_785 ();
 sg13g2_decap_8 FILLER_72_792 ();
 sg13g2_decap_8 FILLER_72_799 ();
 sg13g2_decap_8 FILLER_72_806 ();
 sg13g2_decap_8 FILLER_72_813 ();
 sg13g2_decap_8 FILLER_72_820 ();
 sg13g2_decap_8 FILLER_72_827 ();
 sg13g2_decap_8 FILLER_72_834 ();
 sg13g2_decap_8 FILLER_72_841 ();
 sg13g2_decap_8 FILLER_72_848 ();
 sg13g2_decap_8 FILLER_72_855 ();
 sg13g2_decap_8 FILLER_72_862 ();
 sg13g2_decap_8 FILLER_72_869 ();
 sg13g2_fill_2 FILLER_72_876 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_27 ();
 sg13g2_fill_1 FILLER_73_58 ();
 sg13g2_fill_2 FILLER_73_121 ();
 sg13g2_fill_2 FILLER_73_203 ();
 sg13g2_fill_1 FILLER_73_210 ();
 sg13g2_fill_1 FILLER_73_304 ();
 sg13g2_fill_1 FILLER_73_310 ();
 sg13g2_fill_1 FILLER_73_315 ();
 sg13g2_fill_1 FILLER_73_321 ();
 sg13g2_fill_1 FILLER_73_359 ();
 sg13g2_fill_1 FILLER_73_365 ();
 sg13g2_fill_1 FILLER_73_375 ();
 sg13g2_fill_2 FILLER_73_391 ();
 sg13g2_fill_1 FILLER_73_404 ();
 sg13g2_fill_2 FILLER_73_427 ();
 sg13g2_decap_8 FILLER_73_444 ();
 sg13g2_decap_4 FILLER_73_451 ();
 sg13g2_fill_1 FILLER_73_455 ();
 sg13g2_fill_1 FILLER_73_471 ();
 sg13g2_fill_2 FILLER_73_476 ();
 sg13g2_fill_1 FILLER_73_482 ();
 sg13g2_fill_2 FILLER_73_488 ();
 sg13g2_fill_1 FILLER_73_502 ();
 sg13g2_fill_1 FILLER_73_527 ();
 sg13g2_fill_1 FILLER_73_541 ();
 sg13g2_fill_2 FILLER_73_562 ();
 sg13g2_fill_1 FILLER_73_590 ();
 sg13g2_fill_1 FILLER_73_596 ();
 sg13g2_fill_2 FILLER_73_607 ();
 sg13g2_fill_1 FILLER_73_609 ();
 sg13g2_fill_1 FILLER_73_622 ();
 sg13g2_fill_2 FILLER_73_639 ();
 sg13g2_fill_1 FILLER_73_650 ();
 sg13g2_fill_1 FILLER_73_655 ();
 sg13g2_fill_1 FILLER_73_680 ();
 sg13g2_fill_2 FILLER_73_715 ();
 sg13g2_decap_8 FILLER_73_729 ();
 sg13g2_decap_8 FILLER_73_736 ();
 sg13g2_decap_8 FILLER_73_743 ();
 sg13g2_decap_8 FILLER_73_750 ();
 sg13g2_decap_8 FILLER_73_757 ();
 sg13g2_decap_8 FILLER_73_764 ();
 sg13g2_decap_8 FILLER_73_771 ();
 sg13g2_decap_8 FILLER_73_778 ();
 sg13g2_decap_8 FILLER_73_785 ();
 sg13g2_decap_8 FILLER_73_792 ();
 sg13g2_decap_8 FILLER_73_799 ();
 sg13g2_decap_8 FILLER_73_806 ();
 sg13g2_decap_8 FILLER_73_813 ();
 sg13g2_decap_8 FILLER_73_820 ();
 sg13g2_decap_8 FILLER_73_827 ();
 sg13g2_decap_8 FILLER_73_834 ();
 sg13g2_decap_8 FILLER_73_841 ();
 sg13g2_decap_8 FILLER_73_848 ();
 sg13g2_decap_8 FILLER_73_855 ();
 sg13g2_decap_8 FILLER_73_862 ();
 sg13g2_decap_8 FILLER_73_869 ();
 sg13g2_fill_2 FILLER_73_876 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_15 ();
 sg13g2_fill_1 FILLER_74_26 ();
 sg13g2_fill_1 FILLER_74_37 ();
 sg13g2_fill_1 FILLER_74_42 ();
 sg13g2_fill_1 FILLER_74_53 ();
 sg13g2_fill_1 FILLER_74_80 ();
 sg13g2_fill_1 FILLER_74_91 ();
 sg13g2_fill_1 FILLER_74_156 ();
 sg13g2_fill_2 FILLER_74_225 ();
 sg13g2_fill_1 FILLER_74_365 ();
 sg13g2_fill_1 FILLER_74_371 ();
 sg13g2_fill_1 FILLER_74_381 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_2 FILLER_74_410 ();
 sg13g2_decap_4 FILLER_74_421 ();
 sg13g2_fill_2 FILLER_74_428 ();
 sg13g2_fill_1 FILLER_74_435 ();
 sg13g2_fill_1 FILLER_74_440 ();
 sg13g2_fill_1 FILLER_74_471 ();
 sg13g2_fill_2 FILLER_74_476 ();
 sg13g2_fill_1 FILLER_74_486 ();
 sg13g2_fill_2 FILLER_74_511 ();
 sg13g2_fill_2 FILLER_74_544 ();
 sg13g2_fill_2 FILLER_74_554 ();
 sg13g2_fill_1 FILLER_74_556 ();
 sg13g2_fill_2 FILLER_74_581 ();
 sg13g2_fill_1 FILLER_74_583 ();
 sg13g2_decap_4 FILLER_74_610 ();
 sg13g2_fill_1 FILLER_74_614 ();
 sg13g2_fill_2 FILLER_74_711 ();
 sg13g2_decap_8 FILLER_74_730 ();
 sg13g2_decap_8 FILLER_74_737 ();
 sg13g2_decap_8 FILLER_74_744 ();
 sg13g2_decap_8 FILLER_74_751 ();
 sg13g2_decap_8 FILLER_74_758 ();
 sg13g2_decap_8 FILLER_74_765 ();
 sg13g2_decap_8 FILLER_74_772 ();
 sg13g2_decap_8 FILLER_74_779 ();
 sg13g2_decap_8 FILLER_74_786 ();
 sg13g2_decap_8 FILLER_74_793 ();
 sg13g2_decap_8 FILLER_74_800 ();
 sg13g2_decap_8 FILLER_74_807 ();
 sg13g2_decap_8 FILLER_74_814 ();
 sg13g2_decap_8 FILLER_74_821 ();
 sg13g2_decap_8 FILLER_74_828 ();
 sg13g2_decap_8 FILLER_74_835 ();
 sg13g2_decap_8 FILLER_74_842 ();
 sg13g2_decap_8 FILLER_74_849 ();
 sg13g2_decap_8 FILLER_74_856 ();
 sg13g2_decap_8 FILLER_74_863 ();
 sg13g2_decap_8 FILLER_74_870 ();
 sg13g2_fill_1 FILLER_74_877 ();
 sg13g2_fill_1 FILLER_75_14 ();
 sg13g2_fill_2 FILLER_75_103 ();
 sg13g2_fill_1 FILLER_75_152 ();
 sg13g2_fill_2 FILLER_75_215 ();
 sg13g2_fill_1 FILLER_75_235 ();
 sg13g2_fill_1 FILLER_75_241 ();
 sg13g2_fill_1 FILLER_75_260 ();
 sg13g2_fill_2 FILLER_75_324 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_fill_1 FILLER_75_337 ();
 sg13g2_fill_2 FILLER_75_371 ();
 sg13g2_fill_1 FILLER_75_373 ();
 sg13g2_fill_2 FILLER_75_387 ();
 sg13g2_fill_2 FILLER_75_394 ();
 sg13g2_fill_1 FILLER_75_402 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_fill_1 FILLER_75_414 ();
 sg13g2_fill_1 FILLER_75_420 ();
 sg13g2_fill_2 FILLER_75_437 ();
 sg13g2_fill_1 FILLER_75_439 ();
 sg13g2_fill_2 FILLER_75_445 ();
 sg13g2_fill_1 FILLER_75_447 ();
 sg13g2_decap_8 FILLER_75_452 ();
 sg13g2_fill_1 FILLER_75_459 ();
 sg13g2_fill_1 FILLER_75_488 ();
 sg13g2_fill_2 FILLER_75_512 ();
 sg13g2_fill_1 FILLER_75_514 ();
 sg13g2_fill_1 FILLER_75_528 ();
 sg13g2_fill_1 FILLER_75_554 ();
 sg13g2_fill_1 FILLER_75_563 ();
 sg13g2_fill_2 FILLER_75_569 ();
 sg13g2_fill_2 FILLER_75_609 ();
 sg13g2_fill_1 FILLER_75_611 ();
 sg13g2_fill_2 FILLER_75_617 ();
 sg13g2_fill_1 FILLER_75_660 ();
 sg13g2_fill_1 FILLER_75_673 ();
 sg13g2_fill_1 FILLER_75_679 ();
 sg13g2_decap_8 FILLER_75_700 ();
 sg13g2_decap_8 FILLER_75_707 ();
 sg13g2_decap_8 FILLER_75_714 ();
 sg13g2_decap_8 FILLER_75_721 ();
 sg13g2_decap_8 FILLER_75_728 ();
 sg13g2_decap_8 FILLER_75_735 ();
 sg13g2_decap_8 FILLER_75_742 ();
 sg13g2_decap_8 FILLER_75_749 ();
 sg13g2_decap_8 FILLER_75_756 ();
 sg13g2_decap_8 FILLER_75_763 ();
 sg13g2_decap_8 FILLER_75_770 ();
 sg13g2_decap_8 FILLER_75_777 ();
 sg13g2_decap_8 FILLER_75_784 ();
 sg13g2_decap_8 FILLER_75_791 ();
 sg13g2_decap_8 FILLER_75_798 ();
 sg13g2_decap_8 FILLER_75_805 ();
 sg13g2_decap_8 FILLER_75_812 ();
 sg13g2_decap_8 FILLER_75_819 ();
 sg13g2_decap_8 FILLER_75_826 ();
 sg13g2_decap_8 FILLER_75_833 ();
 sg13g2_decap_8 FILLER_75_840 ();
 sg13g2_decap_8 FILLER_75_847 ();
 sg13g2_decap_8 FILLER_75_854 ();
 sg13g2_decap_8 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_fill_2 FILLER_75_875 ();
 sg13g2_fill_1 FILLER_75_877 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_139 ();
 sg13g2_fill_2 FILLER_76_149 ();
 sg13g2_fill_1 FILLER_76_228 ();
 sg13g2_fill_1 FILLER_76_301 ();
 sg13g2_fill_1 FILLER_76_306 ();
 sg13g2_fill_1 FILLER_76_343 ();
 sg13g2_fill_1 FILLER_76_355 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_1 FILLER_76_406 ();
 sg13g2_fill_1 FILLER_76_412 ();
 sg13g2_fill_1 FILLER_76_425 ();
 sg13g2_fill_1 FILLER_76_434 ();
 sg13g2_fill_2 FILLER_76_439 ();
 sg13g2_fill_2 FILLER_76_467 ();
 sg13g2_fill_1 FILLER_76_479 ();
 sg13g2_fill_1 FILLER_76_489 ();
 sg13g2_fill_2 FILLER_76_498 ();
 sg13g2_decap_8 FILLER_76_514 ();
 sg13g2_decap_4 FILLER_76_521 ();
 sg13g2_fill_1 FILLER_76_525 ();
 sg13g2_fill_1 FILLER_76_578 ();
 sg13g2_fill_2 FILLER_76_583 ();
 sg13g2_fill_1 FILLER_76_585 ();
 sg13g2_fill_1 FILLER_76_612 ();
 sg13g2_decap_8 FILLER_76_676 ();
 sg13g2_decap_8 FILLER_76_683 ();
 sg13g2_decap_8 FILLER_76_690 ();
 sg13g2_decap_8 FILLER_76_697 ();
 sg13g2_decap_8 FILLER_76_704 ();
 sg13g2_decap_8 FILLER_76_711 ();
 sg13g2_decap_8 FILLER_76_718 ();
 sg13g2_decap_8 FILLER_76_725 ();
 sg13g2_decap_8 FILLER_76_732 ();
 sg13g2_decap_8 FILLER_76_739 ();
 sg13g2_decap_8 FILLER_76_746 ();
 sg13g2_decap_8 FILLER_76_753 ();
 sg13g2_decap_8 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_767 ();
 sg13g2_decap_8 FILLER_76_774 ();
 sg13g2_decap_8 FILLER_76_781 ();
 sg13g2_decap_8 FILLER_76_788 ();
 sg13g2_decap_8 FILLER_76_795 ();
 sg13g2_decap_8 FILLER_76_802 ();
 sg13g2_decap_8 FILLER_76_809 ();
 sg13g2_decap_8 FILLER_76_816 ();
 sg13g2_decap_8 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_830 ();
 sg13g2_decap_8 FILLER_76_837 ();
 sg13g2_decap_8 FILLER_76_844 ();
 sg13g2_decap_8 FILLER_76_851 ();
 sg13g2_decap_8 FILLER_76_858 ();
 sg13g2_decap_8 FILLER_76_865 ();
 sg13g2_decap_4 FILLER_76_872 ();
 sg13g2_fill_2 FILLER_76_876 ();
 sg13g2_fill_1 FILLER_77_38 ();
 sg13g2_fill_2 FILLER_77_78 ();
 sg13g2_fill_1 FILLER_77_103 ();
 sg13g2_fill_2 FILLER_77_216 ();
 sg13g2_fill_1 FILLER_77_218 ();
 sg13g2_fill_1 FILLER_77_245 ();
 sg13g2_fill_1 FILLER_77_280 ();
 sg13g2_fill_1 FILLER_77_300 ();
 sg13g2_fill_1 FILLER_77_311 ();
 sg13g2_fill_1 FILLER_77_320 ();
 sg13g2_fill_1 FILLER_77_352 ();
 sg13g2_fill_1 FILLER_77_361 ();
 sg13g2_fill_2 FILLER_77_388 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_decap_8 FILLER_77_449 ();
 sg13g2_fill_2 FILLER_77_456 ();
 sg13g2_fill_1 FILLER_77_458 ();
 sg13g2_fill_2 FILLER_77_509 ();
 sg13g2_fill_1 FILLER_77_519 ();
 sg13g2_fill_1 FILLER_77_528 ();
 sg13g2_fill_1 FILLER_77_534 ();
 sg13g2_fill_1 FILLER_77_540 ();
 sg13g2_fill_1 FILLER_77_579 ();
 sg13g2_fill_2 FILLER_77_610 ();
 sg13g2_fill_1 FILLER_77_612 ();
 sg13g2_fill_1 FILLER_77_621 ();
 sg13g2_fill_1 FILLER_77_626 ();
 sg13g2_decap_8 FILLER_77_661 ();
 sg13g2_decap_8 FILLER_77_668 ();
 sg13g2_decap_8 FILLER_77_675 ();
 sg13g2_decap_8 FILLER_77_682 ();
 sg13g2_decap_8 FILLER_77_689 ();
 sg13g2_decap_8 FILLER_77_696 ();
 sg13g2_decap_8 FILLER_77_703 ();
 sg13g2_decap_8 FILLER_77_710 ();
 sg13g2_decap_8 FILLER_77_717 ();
 sg13g2_decap_8 FILLER_77_724 ();
 sg13g2_decap_8 FILLER_77_731 ();
 sg13g2_decap_8 FILLER_77_738 ();
 sg13g2_decap_8 FILLER_77_745 ();
 sg13g2_decap_8 FILLER_77_752 ();
 sg13g2_decap_8 FILLER_77_759 ();
 sg13g2_decap_8 FILLER_77_766 ();
 sg13g2_decap_8 FILLER_77_773 ();
 sg13g2_decap_8 FILLER_77_780 ();
 sg13g2_decap_8 FILLER_77_787 ();
 sg13g2_decap_8 FILLER_77_794 ();
 sg13g2_decap_8 FILLER_77_801 ();
 sg13g2_decap_8 FILLER_77_808 ();
 sg13g2_decap_8 FILLER_77_815 ();
 sg13g2_decap_8 FILLER_77_822 ();
 sg13g2_decap_8 FILLER_77_829 ();
 sg13g2_decap_8 FILLER_77_836 ();
 sg13g2_decap_8 FILLER_77_843 ();
 sg13g2_decap_8 FILLER_77_850 ();
 sg13g2_decap_8 FILLER_77_857 ();
 sg13g2_decap_8 FILLER_77_864 ();
 sg13g2_decap_8 FILLER_77_871 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_54 ();
 sg13g2_fill_2 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_79 ();
 sg13g2_fill_1 FILLER_78_92 ();
 sg13g2_fill_1 FILLER_78_101 ();
 sg13g2_fill_1 FILLER_78_194 ();
 sg13g2_fill_2 FILLER_78_199 ();
 sg13g2_fill_2 FILLER_78_205 ();
 sg13g2_fill_1 FILLER_78_207 ();
 sg13g2_fill_2 FILLER_78_280 ();
 sg13g2_fill_2 FILLER_78_343 ();
 sg13g2_fill_1 FILLER_78_370 ();
 sg13g2_fill_1 FILLER_78_375 ();
 sg13g2_fill_1 FILLER_78_380 ();
 sg13g2_fill_1 FILLER_78_386 ();
 sg13g2_fill_1 FILLER_78_392 ();
 sg13g2_fill_2 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_411 ();
 sg13g2_fill_1 FILLER_78_415 ();
 sg13g2_decap_4 FILLER_78_493 ();
 sg13g2_fill_1 FILLER_78_501 ();
 sg13g2_fill_1 FILLER_78_506 ();
 sg13g2_fill_1 FILLER_78_516 ();
 sg13g2_fill_2 FILLER_78_522 ();
 sg13g2_fill_1 FILLER_78_586 ();
 sg13g2_fill_1 FILLER_78_651 ();
 sg13g2_decap_8 FILLER_78_668 ();
 sg13g2_decap_8 FILLER_78_675 ();
 sg13g2_decap_8 FILLER_78_682 ();
 sg13g2_decap_8 FILLER_78_689 ();
 sg13g2_decap_8 FILLER_78_696 ();
 sg13g2_decap_8 FILLER_78_703 ();
 sg13g2_decap_8 FILLER_78_710 ();
 sg13g2_decap_8 FILLER_78_717 ();
 sg13g2_decap_8 FILLER_78_724 ();
 sg13g2_decap_8 FILLER_78_731 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_decap_8 FILLER_78_745 ();
 sg13g2_decap_8 FILLER_78_752 ();
 sg13g2_decap_8 FILLER_78_759 ();
 sg13g2_decap_8 FILLER_78_766 ();
 sg13g2_decap_8 FILLER_78_773 ();
 sg13g2_decap_8 FILLER_78_780 ();
 sg13g2_decap_8 FILLER_78_787 ();
 sg13g2_decap_8 FILLER_78_794 ();
 sg13g2_decap_8 FILLER_78_801 ();
 sg13g2_decap_8 FILLER_78_808 ();
 sg13g2_decap_8 FILLER_78_815 ();
 sg13g2_decap_8 FILLER_78_822 ();
 sg13g2_decap_8 FILLER_78_829 ();
 sg13g2_decap_8 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_843 ();
 sg13g2_decap_8 FILLER_78_850 ();
 sg13g2_decap_8 FILLER_78_857 ();
 sg13g2_decap_8 FILLER_78_864 ();
 sg13g2_decap_8 FILLER_78_871 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_2 ();
 sg13g2_fill_1 FILLER_79_34 ();
 sg13g2_fill_1 FILLER_79_237 ();
 sg13g2_fill_2 FILLER_79_356 ();
 sg13g2_fill_2 FILLER_79_369 ();
 sg13g2_fill_1 FILLER_79_375 ();
 sg13g2_fill_1 FILLER_79_381 ();
 sg13g2_fill_1 FILLER_79_411 ();
 sg13g2_decap_4 FILLER_79_425 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_79_440 ();
 sg13g2_fill_2 FILLER_79_467 ();
 sg13g2_fill_1 FILLER_79_481 ();
 sg13g2_fill_1 FILLER_79_487 ();
 sg13g2_fill_1 FILLER_79_527 ();
 sg13g2_fill_1 FILLER_79_537 ();
 sg13g2_fill_1 FILLER_79_543 ();
 sg13g2_fill_1 FILLER_79_554 ();
 sg13g2_decap_4 FILLER_79_559 ();
 sg13g2_fill_1 FILLER_79_563 ();
 sg13g2_decap_8 FILLER_79_571 ();
 sg13g2_decap_4 FILLER_79_578 ();
 sg13g2_fill_2 FILLER_79_587 ();
 sg13g2_fill_1 FILLER_79_594 ();
 sg13g2_fill_1 FILLER_79_599 ();
 sg13g2_fill_2 FILLER_79_604 ();
 sg13g2_fill_1 FILLER_79_606 ();
 sg13g2_fill_2 FILLER_79_616 ();
 sg13g2_fill_1 FILLER_79_637 ();
 sg13g2_fill_2 FILLER_79_657 ();
 sg13g2_decap_8 FILLER_79_663 ();
 sg13g2_fill_2 FILLER_79_670 ();
 sg13g2_fill_1 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_678 ();
 sg13g2_decap_8 FILLER_79_685 ();
 sg13g2_decap_8 FILLER_79_692 ();
 sg13g2_decap_8 FILLER_79_699 ();
 sg13g2_decap_8 FILLER_79_706 ();
 sg13g2_decap_8 FILLER_79_713 ();
 sg13g2_decap_8 FILLER_79_720 ();
 sg13g2_decap_8 FILLER_79_727 ();
 sg13g2_decap_8 FILLER_79_734 ();
 sg13g2_decap_8 FILLER_79_741 ();
 sg13g2_decap_8 FILLER_79_748 ();
 sg13g2_decap_8 FILLER_79_755 ();
 sg13g2_decap_8 FILLER_79_762 ();
 sg13g2_decap_8 FILLER_79_769 ();
 sg13g2_decap_8 FILLER_79_776 ();
 sg13g2_decap_8 FILLER_79_783 ();
 sg13g2_decap_8 FILLER_79_790 ();
 sg13g2_decap_8 FILLER_79_797 ();
 sg13g2_decap_8 FILLER_79_804 ();
 sg13g2_decap_8 FILLER_79_811 ();
 sg13g2_decap_8 FILLER_79_818 ();
 sg13g2_decap_8 FILLER_79_825 ();
 sg13g2_decap_8 FILLER_79_832 ();
 sg13g2_decap_8 FILLER_79_839 ();
 sg13g2_decap_8 FILLER_79_846 ();
 sg13g2_decap_8 FILLER_79_853 ();
 sg13g2_decap_8 FILLER_79_860 ();
 sg13g2_decap_8 FILLER_79_867 ();
 sg13g2_decap_4 FILLER_79_874 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_20 ();
 sg13g2_fill_1 FILLER_80_79 ();
 sg13g2_fill_1 FILLER_80_202 ();
 sg13g2_fill_1 FILLER_80_269 ();
 sg13g2_fill_1 FILLER_80_308 ();
 sg13g2_fill_1 FILLER_80_366 ();
 sg13g2_decap_8 FILLER_80_423 ();
 sg13g2_decap_8 FILLER_80_430 ();
 sg13g2_decap_4 FILLER_80_437 ();
 sg13g2_fill_2 FILLER_80_441 ();
 sg13g2_fill_2 FILLER_80_508 ();
 sg13g2_fill_1 FILLER_80_510 ();
 sg13g2_fill_2 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_574 ();
 sg13g2_decap_4 FILLER_80_581 ();
 sg13g2_fill_2 FILLER_80_585 ();
 sg13g2_decap_4 FILLER_80_618 ();
 sg13g2_decap_8 FILLER_80_679 ();
 sg13g2_decap_8 FILLER_80_686 ();
 sg13g2_decap_8 FILLER_80_693 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_8 FILLER_80_707 ();
 sg13g2_decap_8 FILLER_80_714 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_decap_8 FILLER_80_770 ();
 sg13g2_decap_8 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_833 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_decap_8 FILLER_80_861 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_fill_2 FILLER_80_875 ();
 sg13g2_fill_1 FILLER_80_877 ();
endmodule
