module tt_um_urish_sram_test (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire clknet_0_clk;
 wire net77;
 wire \addr[6] ;
 wire \addr[7] ;
 wire \addr[8] ;
 wire \addr[9] ;
 wire \addr_high_reg[0] ;
 wire \addr_high_reg[1] ;
 wire \addr_high_reg[2] ;
 wire \addr_high_reg[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sg13g2_inv_1 _12_ (.Y(_01_),
    .A(net13));
 sg13g2_nor2_1 _13_ (.A(_01_),
    .B(net12),
    .Y(_00_));
 sg13g2_mux2_2 _14_ (.A0(net4),
    .A1(net14),
    .S(net12),
    .X(\addr[6] ));
 sg13g2_and2_1 _15_ (.A(net5),
    .B(\addr[6] ),
    .X(_02_));
 sg13g2_mux2_2 _16_ (.A0(net2),
    .A1(net15),
    .S(net12),
    .X(\addr[7] ));
 sg13g2_and2_1 _17_ (.A(net5),
    .B(\addr[7] ),
    .X(_03_));
 sg13g2_mux2_2 _18_ (.A0(net3),
    .A1(net16),
    .S(net12),
    .X(\addr[8] ));
 sg13g2_and2_1 _19_ (.A(net5),
    .B(\addr[8] ),
    .X(_04_));
 sg13g2_mux2_2 _20_ (.A0(net1),
    .A1(net17),
    .S(net12),
    .X(\addr[9] ));
 sg13g2_and2_1 _21_ (.A(net5),
    .B(\addr[9] ),
    .X(_05_));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \addr_high_reg[0]$_SDFF_PN0__73  (.L_HI(net77));
 sg13g2_buf_1 _24_ (.A(net30),
    .X(uio_oe[0]));
 sg13g2_buf_1 _25_ (.A(net31),
    .X(uio_oe[1]));
 sg13g2_buf_1 _26_ (.A(net32),
    .X(uio_oe[2]));
 sg13g2_buf_1 _27_ (.A(net33),
    .X(uio_oe[3]));
 sg13g2_buf_1 _28_ (.A(net34),
    .X(uio_oe[4]));
 sg13g2_buf_1 _29_ (.A(net35),
    .X(uio_oe[5]));
 sg13g2_buf_1 _30_ (.A(net36),
    .X(uio_oe[6]));
 sg13g2_buf_1 _31_ (.A(net37),
    .X(uio_oe[7]));
 sg13g2_buf_1 _32_ (.A(net38),
    .X(uio_out[0]));
 sg13g2_buf_1 _33_ (.A(net39),
    .X(uio_out[1]));
 sg13g2_buf_1 _34_ (.A(net40),
    .X(uio_out[2]));
 sg13g2_buf_1 _35_ (.A(net41),
    .X(uio_out[3]));
 sg13g2_buf_1 _36_ (.A(net42),
    .X(uio_out[4]));
 sg13g2_buf_1 _37_ (.A(net43),
    .X(uio_out[5]));
 sg13g2_buf_1 _38_ (.A(net44),
    .X(uio_out[6]));
 sg13g2_buf_1 _39_ (.A(net45),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \addr_high_reg[0]$_SDFF_PN0_  (.CLK(clknet_1_1__leaf_clk),
    .RESET_B(net77),
    .D(_02_),
    .Q_N(_09_),
    .Q(\addr_high_reg[0] ));
 sg13g2_dfrbp_1 \addr_high_reg[1]$_SDFF_PN0_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net78),
    .D(_03_),
    .Q_N(_08_),
    .Q(\addr_high_reg[1] ));
 sg13g2_dfrbp_1 \addr_high_reg[2]$_SDFF_PN0_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net79),
    .D(_04_),
    .Q_N(_07_),
    .Q(\addr_high_reg[2] ));
 sg13g2_dfrbp_1 \addr_high_reg[3]$_SDFF_PN0_  (.CLK(clknet_1_0__leaf_clk),
    .RESET_B(net80),
    .D(_05_),
    .Q_N(_06_),
    .Q(\addr_high_reg[3] ));
 RM_IHPSG13_1P_1024x8_c2_bm_bist sram (.A_CLK(clknet_1_1__leaf_clk),
    .A_REN(_01_),
    .A_WEN(_00_),
    .A_MEN(net5),
    .A_DLY(net89),
    .A_BIST_EN(net72),
    .A_BIST_CLK(net73),
    .A_BIST_REN(net74),
    .A_BIST_WEN(net75),
    .A_BIST_MEN(net76),
    .A_ADDR({\addr[9] ,
    \addr[8] ,
    \addr[7] ,
    \addr[6] ,
    net11,
    net10,
    net9,
    net8,
    net7,
    net6}),
    .A_BIST_ADDR({net71,
    net70,
    net69,
    net68,
    net67,
    net66,
    net65,
    net64,
    net63,
    net62}),
    .A_BIST_BM({net60,
    net56,
    net52,
    net48,
    net49,
    net53,
    net57,
    net61}),
    .A_BIST_DIN({net58,
    net54,
    net50,
    net46,
    net47,
    net51,
    net55,
    net59}),
    .A_BM({net87,
    net85,
    net83,
    net81,
    net82,
    net84,
    net86,
    net88}),
    .A_DIN({net21,
    net20,
    net19,
    net18,
    net17,
    net16,
    net15,
    net14}),
    .A_DOUT({net29,
    net28,
    net27,
    net26,
    net25,
    net24,
    net23,
    net22}));
 sg13g2_dlygate4sd3_1 hold1 (.A(\addr_high_reg[3] ),
    .X(net1));
 sg13g2_dlygate4sd3_1 hold2 (.A(\addr_high_reg[1] ),
    .X(net2));
 sg13g2_dlygate4sd3_1 hold3 (.A(\addr_high_reg[2] ),
    .X(net3));
 sg13g2_dlygate4sd3_1 hold4 (.A(\addr_high_reg[0] ),
    .X(net4));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net5));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net6));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net7));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net8));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net9));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net10));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net11));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net12));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net13));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net14));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net15));
 sg13g2_buf_1 input12 (.A(uio_in[2]),
    .X(net16));
 sg13g2_buf_1 input13 (.A(uio_in[3]),
    .X(net17));
 sg13g2_buf_1 input14 (.A(uio_in[4]),
    .X(net18));
 sg13g2_buf_1 input15 (.A(uio_in[5]),
    .X(net19));
 sg13g2_buf_1 input16 (.A(uio_in[6]),
    .X(net20));
 sg13g2_buf_1 input17 (.A(uio_in[7]),
    .X(net21));
 sg13g2_buf_1 output18 (.A(net22),
    .X(uo_out[0]));
 sg13g2_buf_1 output19 (.A(net23),
    .X(uo_out[1]));
 sg13g2_buf_1 output20 (.A(net24),
    .X(uo_out[2]));
 sg13g2_buf_1 output21 (.A(net25),
    .X(uo_out[3]));
 sg13g2_buf_1 output22 (.A(net26),
    .X(uo_out[4]));
 sg13g2_buf_1 output23 (.A(net27),
    .X(uo_out[5]));
 sg13g2_buf_1 output24 (.A(net28),
    .X(uo_out[6]));
 sg13g2_buf_1 output25 (.A(net29),
    .X(uo_out[7]));
 sg13g2_tielo _24__26 (.L_LO(net30));
 sg13g2_tielo _25__27 (.L_LO(net31));
 sg13g2_tielo _26__28 (.L_LO(net32));
 sg13g2_tielo _27__29 (.L_LO(net33));
 sg13g2_tielo _28__30 (.L_LO(net34));
 sg13g2_tielo _29__31 (.L_LO(net35));
 sg13g2_tielo _30__32 (.L_LO(net36));
 sg13g2_tielo _31__33 (.L_LO(net37));
 sg13g2_tielo _32__34 (.L_LO(net38));
 sg13g2_tielo _33__35 (.L_LO(net39));
 sg13g2_tielo _34__36 (.L_LO(net40));
 sg13g2_tielo _35__37 (.L_LO(net41));
 sg13g2_tielo _36__38 (.L_LO(net42));
 sg13g2_tielo _37__39 (.L_LO(net43));
 sg13g2_tielo _38__40 (.L_LO(net44));
 sg13g2_tielo _39__41 (.L_LO(net45));
 sg13g2_tielo sram_42 (.L_LO(net46));
 sg13g2_tielo sram_43 (.L_LO(net47));
 sg13g2_tielo sram_44 (.L_LO(net48));
 sg13g2_tielo sram_45 (.L_LO(net49));
 sg13g2_tielo sram_46 (.L_LO(net50));
 sg13g2_tielo sram_47 (.L_LO(net51));
 sg13g2_tielo sram_48 (.L_LO(net52));
 sg13g2_tielo sram_49 (.L_LO(net53));
 sg13g2_tielo sram_50 (.L_LO(net54));
 sg13g2_tielo sram_51 (.L_LO(net55));
 sg13g2_tielo sram_52 (.L_LO(net56));
 sg13g2_tielo sram_53 (.L_LO(net57));
 sg13g2_tielo sram_54 (.L_LO(net58));
 sg13g2_tielo sram_55 (.L_LO(net59));
 sg13g2_tielo sram_56 (.L_LO(net60));
 sg13g2_tielo sram_57 (.L_LO(net61));
 sg13g2_tielo sram_58 (.L_LO(net62));
 sg13g2_tielo sram_59 (.L_LO(net63));
 sg13g2_tielo sram_60 (.L_LO(net64));
 sg13g2_tielo sram_61 (.L_LO(net65));
 sg13g2_tielo sram_62 (.L_LO(net66));
 sg13g2_tielo sram_63 (.L_LO(net67));
 sg13g2_tielo sram_64 (.L_LO(net68));
 sg13g2_tielo sram_65 (.L_LO(net69));
 sg13g2_tielo sram_66 (.L_LO(net70));
 sg13g2_tielo sram_67 (.L_LO(net71));
 sg13g2_tielo sram_68 (.L_LO(net72));
 sg13g2_tielo sram_69 (.L_LO(net73));
 sg13g2_tielo sram_70 (.L_LO(net74));
 sg13g2_tielo sram_71 (.L_LO(net75));
 sg13g2_tielo sram_72 (.L_LO(net76));
 sg13g2_tiehi \addr_high_reg[1]$_SDFF_PN0__74  (.L_HI(net78));
 sg13g2_tiehi \addr_high_reg[2]$_SDFF_PN0__75  (.L_HI(net79));
 sg13g2_tiehi \addr_high_reg[3]$_SDFF_PN0__76  (.L_HI(net80));
 sg13g2_tiehi sram_77 (.L_HI(net81));
 sg13g2_tiehi sram_78 (.L_HI(net82));
 sg13g2_tiehi sram_79 (.L_HI(net83));
 sg13g2_tiehi sram_80 (.L_HI(net84));
 sg13g2_tiehi sram_81 (.L_HI(net85));
 sg13g2_tiehi sram_82 (.L_HI(net86));
 sg13g2_tiehi sram_83 (.L_HI(net87));
 sg13g2_tiehi sram_84 (.L_HI(net88));
 sg13g2_tiehi sram_85 (.L_HI(net89));
 sg13g2_buf_2 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_2 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_2 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_3 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_4 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_antennanp ANTENNA_7 (.A(clk));
 sg13g2_antennanp ANTENNA_8 (.A(net22));
 sg13g2_antennanp ANTENNA_9 (.A(net22));
 sg13g2_antennanp ANTENNA_10 (.A(net23));
 sg13g2_antennanp ANTENNA_11 (.A(net23));
 sg13g2_antennanp ANTENNA_12 (.A(net24));
 sg13g2_antennanp ANTENNA_13 (.A(net24));
 sg13g2_antennanp ANTENNA_14 (.A(net25));
 sg13g2_antennanp ANTENNA_15 (.A(net25));
 sg13g2_antennanp ANTENNA_16 (.A(net26));
 sg13g2_antennanp ANTENNA_17 (.A(net26));
 sg13g2_antennanp ANTENNA_18 (.A(net27));
 sg13g2_antennanp ANTENNA_19 (.A(net27));
 sg13g2_antennanp ANTENNA_20 (.A(net28));
 sg13g2_antennanp ANTENNA_21 (.A(net28));
 sg13g2_antennanp ANTENNA_22 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_23 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_24 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_25 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_26 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_27 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_28 (.A(clk));
 sg13g2_antennanp ANTENNA_29 (.A(clk));
 sg13g2_antennanp ANTENNA_30 (.A(clk));
 sg13g2_antennanp ANTENNA_31 (.A(net22));
 sg13g2_antennanp ANTENNA_32 (.A(net22));
 sg13g2_antennanp ANTENNA_33 (.A(net23));
 sg13g2_antennanp ANTENNA_34 (.A(net23));
 sg13g2_antennanp ANTENNA_35 (.A(net24));
 sg13g2_antennanp ANTENNA_36 (.A(net24));
 sg13g2_antennanp ANTENNA_37 (.A(net25));
 sg13g2_antennanp ANTENNA_38 (.A(net25));
 sg13g2_antennanp ANTENNA_39 (.A(net26));
 sg13g2_antennanp ANTENNA_40 (.A(net26));
 sg13g2_antennanp ANTENNA_41 (.A(net27));
 sg13g2_antennanp ANTENNA_42 (.A(net27));
 sg13g2_antennanp ANTENNA_43 (.A(net28));
 sg13g2_antennanp ANTENNA_44 (.A(net28));
 sg13g2_antennanp ANTENNA_45 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_46 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_47 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_48 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_49 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_50 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_51 (.A(clk));
 sg13g2_antennanp ANTENNA_52 (.A(clk));
 sg13g2_antennanp ANTENNA_53 (.A(clk));
 sg13g2_antennanp ANTENNA_54 (.A(net22));
 sg13g2_antennanp ANTENNA_55 (.A(net22));
 sg13g2_antennanp ANTENNA_56 (.A(net23));
 sg13g2_antennanp ANTENNA_57 (.A(net23));
 sg13g2_antennanp ANTENNA_58 (.A(net24));
 sg13g2_antennanp ANTENNA_59 (.A(net24));
 sg13g2_antennanp ANTENNA_60 (.A(net25));
 sg13g2_antennanp ANTENNA_61 (.A(net25));
 sg13g2_antennanp ANTENNA_62 (.A(net26));
 sg13g2_antennanp ANTENNA_63 (.A(net26));
 sg13g2_antennanp ANTENNA_64 (.A(net27));
 sg13g2_antennanp ANTENNA_65 (.A(net27));
 sg13g2_antennanp ANTENNA_66 (.A(net28));
 sg13g2_antennanp ANTENNA_67 (.A(net28));
 sg13g2_antennanp ANTENNA_68 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_69 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_70 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_71 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_72 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_73 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_74 (.A(clk));
 sg13g2_antennanp ANTENNA_75 (.A(clk));
 sg13g2_antennanp ANTENNA_76 (.A(clk));
 sg13g2_antennanp ANTENNA_77 (.A(net22));
 sg13g2_antennanp ANTENNA_78 (.A(net22));
 sg13g2_antennanp ANTENNA_79 (.A(net23));
 sg13g2_antennanp ANTENNA_80 (.A(net23));
 sg13g2_antennanp ANTENNA_81 (.A(net25));
 sg13g2_antennanp ANTENNA_82 (.A(net25));
 sg13g2_antennanp ANTENNA_83 (.A(net26));
 sg13g2_antennanp ANTENNA_84 (.A(net26));
 sg13g2_antennanp ANTENNA_85 (.A(net27));
 sg13g2_antennanp ANTENNA_86 (.A(net27));
 sg13g2_antennanp ANTENNA_87 (.A(net28));
 sg13g2_antennanp ANTENNA_88 (.A(net28));
 sg13g2_antennanp ANTENNA_89 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_90 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_91 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_92 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_93 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_94 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_95 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_96 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_97 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_98 (.A(clknet_0_clk));
 sg13g2_antennanp ANTENNA_99 (.A(clk));
 sg13g2_antennanp ANTENNA_100 (.A(clk));
 sg13g2_antennanp ANTENNA_101 (.A(clk));
 sg13g2_antennanp ANTENNA_102 (.A(net22));
 sg13g2_antennanp ANTENNA_103 (.A(net22));
 sg13g2_antennanp ANTENNA_104 (.A(net23));
 sg13g2_antennanp ANTENNA_105 (.A(net23));
 sg13g2_antennanp ANTENNA_106 (.A(net24));
 sg13g2_antennanp ANTENNA_107 (.A(net24));
 sg13g2_antennanp ANTENNA_108 (.A(net25));
 sg13g2_antennanp ANTENNA_109 (.A(net25));
 sg13g2_antennanp ANTENNA_110 (.A(net26));
 sg13g2_antennanp ANTENNA_111 (.A(net26));
 sg13g2_antennanp ANTENNA_112 (.A(net28));
 sg13g2_antennanp ANTENNA_113 (.A(net28));
 sg13g2_antennanp ANTENNA_114 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_115 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_116 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_117 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_118 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_119 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_120 (.A(clknet_1_1__leaf_clk));
 sg13g2_antennanp ANTENNA_121 (.A(clknet_1_1__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_fill_2 FILLER_0_875 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_fill_2 FILLER_1_875 ();
 sg13g2_fill_1 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_fill_2 FILLER_2_875 ();
 sg13g2_fill_1 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_fill_2 FILLER_3_875 ();
 sg13g2_fill_1 FILLER_3_877 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_fill_2 FILLER_4_875 ();
 sg13g2_fill_1 FILLER_4_877 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_decap_8 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_5_868 ();
 sg13g2_fill_2 FILLER_5_875 ();
 sg13g2_fill_1 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_decap_8 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_6_868 ();
 sg13g2_fill_2 FILLER_6_875 ();
 sg13g2_fill_1 FILLER_6_877 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_fill_2 FILLER_7_875 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_fill_2 FILLER_8_875 ();
 sg13g2_fill_1 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_fill_2 FILLER_9_875 ();
 sg13g2_fill_1 FILLER_9_877 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_decap_8 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_868 ();
 sg13g2_fill_2 FILLER_10_875 ();
 sg13g2_fill_1 FILLER_10_877 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_decap_8 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_11_868 ();
 sg13g2_fill_2 FILLER_11_875 ();
 sg13g2_fill_1 FILLER_11_877 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_decap_8 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_12_868 ();
 sg13g2_fill_2 FILLER_12_875 ();
 sg13g2_fill_1 FILLER_12_877 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_decap_8 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_13_868 ();
 sg13g2_fill_2 FILLER_13_875 ();
 sg13g2_fill_1 FILLER_13_877 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_decap_8 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_14_868 ();
 sg13g2_fill_2 FILLER_14_875 ();
 sg13g2_fill_1 FILLER_14_877 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_decap_8 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_15_868 ();
 sg13g2_fill_2 FILLER_15_875 ();
 sg13g2_fill_1 FILLER_15_877 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_decap_8 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_16_868 ();
 sg13g2_fill_2 FILLER_16_875 ();
 sg13g2_fill_1 FILLER_16_877 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_fill_2 FILLER_17_875 ();
 sg13g2_fill_1 FILLER_17_877 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_decap_8 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_18_868 ();
 sg13g2_fill_2 FILLER_18_875 ();
 sg13g2_fill_1 FILLER_18_877 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_decap_8 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_19_868 ();
 sg13g2_fill_2 FILLER_19_875 ();
 sg13g2_fill_1 FILLER_19_877 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_decap_8 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_20_868 ();
 sg13g2_fill_2 FILLER_20_875 ();
 sg13g2_fill_1 FILLER_20_877 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_21_868 ();
 sg13g2_fill_2 FILLER_21_875 ();
 sg13g2_fill_1 FILLER_21_877 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_8 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_22_847 ();
 sg13g2_decap_8 FILLER_22_854 ();
 sg13g2_decap_8 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_22_868 ();
 sg13g2_fill_2 FILLER_22_875 ();
 sg13g2_fill_1 FILLER_22_877 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_decap_8 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_fill_2 FILLER_23_875 ();
 sg13g2_fill_1 FILLER_23_877 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_decap_8 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_24_847 ();
 sg13g2_decap_8 FILLER_24_854 ();
 sg13g2_decap_8 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_24_868 ();
 sg13g2_fill_2 FILLER_24_875 ();
 sg13g2_fill_1 FILLER_24_877 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_decap_8 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_581 ();
 sg13g2_decap_8 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_decap_8 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_fill_2 FILLER_25_875 ();
 sg13g2_fill_1 FILLER_25_877 ();
 sg13g2_decap_8 FILLER_26_26 ();
 sg13g2_decap_8 FILLER_26_33 ();
 sg13g2_decap_8 FILLER_26_40 ();
 sg13g2_decap_8 FILLER_26_47 ();
 sg13g2_decap_8 FILLER_26_54 ();
 sg13g2_decap_8 FILLER_26_61 ();
 sg13g2_decap_8 FILLER_26_68 ();
 sg13g2_decap_8 FILLER_26_75 ();
 sg13g2_decap_8 FILLER_26_82 ();
 sg13g2_decap_8 FILLER_26_89 ();
 sg13g2_decap_8 FILLER_26_96 ();
 sg13g2_decap_8 FILLER_26_103 ();
 sg13g2_decap_8 FILLER_26_110 ();
 sg13g2_decap_8 FILLER_26_117 ();
 sg13g2_decap_8 FILLER_26_124 ();
 sg13g2_decap_8 FILLER_26_131 ();
 sg13g2_decap_8 FILLER_26_138 ();
 sg13g2_decap_8 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_159 ();
 sg13g2_decap_8 FILLER_26_166 ();
 sg13g2_decap_8 FILLER_26_173 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_decap_8 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_201 ();
 sg13g2_decap_8 FILLER_26_208 ();
 sg13g2_decap_8 FILLER_26_215 ();
 sg13g2_decap_8 FILLER_26_222 ();
 sg13g2_decap_8 FILLER_26_229 ();
 sg13g2_decap_8 FILLER_26_236 ();
 sg13g2_decap_8 FILLER_26_243 ();
 sg13g2_decap_8 FILLER_26_250 ();
 sg13g2_decap_8 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_264 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_decap_8 FILLER_26_278 ();
 sg13g2_decap_8 FILLER_26_285 ();
 sg13g2_decap_8 FILLER_26_292 ();
 sg13g2_decap_8 FILLER_26_299 ();
 sg13g2_decap_8 FILLER_26_306 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_decap_8 FILLER_26_320 ();
 sg13g2_decap_8 FILLER_26_327 ();
 sg13g2_decap_8 FILLER_26_334 ();
 sg13g2_decap_8 FILLER_26_341 ();
 sg13g2_decap_8 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_8 FILLER_26_404 ();
 sg13g2_decap_8 FILLER_26_411 ();
 sg13g2_decap_8 FILLER_26_418 ();
 sg13g2_decap_8 FILLER_26_425 ();
 sg13g2_decap_8 FILLER_26_432 ();
 sg13g2_decap_8 FILLER_26_439 ();
 sg13g2_decap_8 FILLER_26_446 ();
 sg13g2_decap_8 FILLER_26_453 ();
 sg13g2_decap_8 FILLER_26_460 ();
 sg13g2_decap_8 FILLER_26_467 ();
 sg13g2_decap_8 FILLER_26_474 ();
 sg13g2_decap_8 FILLER_26_481 ();
 sg13g2_decap_8 FILLER_26_488 ();
 sg13g2_decap_8 FILLER_26_495 ();
 sg13g2_decap_8 FILLER_26_502 ();
 sg13g2_decap_8 FILLER_26_509 ();
 sg13g2_decap_8 FILLER_26_516 ();
 sg13g2_decap_8 FILLER_26_523 ();
 sg13g2_decap_8 FILLER_26_530 ();
 sg13g2_decap_8 FILLER_26_537 ();
 sg13g2_decap_8 FILLER_26_544 ();
 sg13g2_decap_8 FILLER_26_551 ();
 sg13g2_decap_8 FILLER_26_558 ();
 sg13g2_decap_8 FILLER_26_565 ();
 sg13g2_decap_8 FILLER_26_572 ();
 sg13g2_decap_8 FILLER_26_579 ();
 sg13g2_decap_8 FILLER_26_586 ();
 sg13g2_decap_8 FILLER_26_593 ();
 sg13g2_decap_8 FILLER_26_600 ();
 sg13g2_decap_8 FILLER_26_607 ();
 sg13g2_decap_8 FILLER_26_614 ();
 sg13g2_decap_8 FILLER_26_621 ();
 sg13g2_decap_8 FILLER_26_628 ();
 sg13g2_decap_8 FILLER_26_635 ();
 sg13g2_decap_8 FILLER_26_642 ();
 sg13g2_decap_8 FILLER_26_649 ();
 sg13g2_decap_8 FILLER_26_656 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_684 ();
 sg13g2_decap_8 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_698 ();
 sg13g2_decap_8 FILLER_26_705 ();
 sg13g2_decap_8 FILLER_26_712 ();
 sg13g2_decap_8 FILLER_26_719 ();
 sg13g2_decap_8 FILLER_26_726 ();
 sg13g2_decap_8 FILLER_26_733 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_decap_8 FILLER_26_747 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_decap_8 FILLER_26_859 ();
 sg13g2_decap_8 FILLER_26_866 ();
 sg13g2_decap_4 FILLER_26_873 ();
 sg13g2_fill_1 FILLER_26_877 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_15 ();
 sg13g2_decap_8 FILLER_27_22 ();
 sg13g2_decap_8 FILLER_27_29 ();
 sg13g2_decap_8 FILLER_27_36 ();
 sg13g2_decap_8 FILLER_27_43 ();
 sg13g2_decap_8 FILLER_27_50 ();
 sg13g2_decap_8 FILLER_27_57 ();
 sg13g2_decap_8 FILLER_27_64 ();
 sg13g2_decap_8 FILLER_27_71 ();
 sg13g2_decap_8 FILLER_27_78 ();
 sg13g2_decap_8 FILLER_27_85 ();
 sg13g2_decap_8 FILLER_27_92 ();
 sg13g2_decap_8 FILLER_27_99 ();
 sg13g2_decap_8 FILLER_27_106 ();
 sg13g2_decap_8 FILLER_27_113 ();
 sg13g2_decap_8 FILLER_27_120 ();
 sg13g2_decap_8 FILLER_27_127 ();
 sg13g2_decap_8 FILLER_27_134 ();
 sg13g2_decap_8 FILLER_27_141 ();
 sg13g2_decap_8 FILLER_27_148 ();
 sg13g2_decap_8 FILLER_27_155 ();
 sg13g2_decap_8 FILLER_27_162 ();
 sg13g2_decap_8 FILLER_27_169 ();
 sg13g2_decap_8 FILLER_27_176 ();
 sg13g2_decap_8 FILLER_27_183 ();
 sg13g2_decap_8 FILLER_27_190 ();
 sg13g2_decap_8 FILLER_27_197 ();
 sg13g2_decap_8 FILLER_27_204 ();
 sg13g2_decap_8 FILLER_27_211 ();
 sg13g2_decap_8 FILLER_27_218 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_decap_8 FILLER_27_232 ();
 sg13g2_decap_8 FILLER_27_239 ();
 sg13g2_decap_8 FILLER_27_246 ();
 sg13g2_decap_8 FILLER_27_253 ();
 sg13g2_decap_8 FILLER_27_260 ();
 sg13g2_decap_4 FILLER_27_267 ();
 sg13g2_decap_8 FILLER_27_274 ();
 sg13g2_decap_8 FILLER_27_281 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_302 ();
 sg13g2_decap_8 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_8 FILLER_27_330 ();
 sg13g2_decap_8 FILLER_27_337 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_27_424 ();
 sg13g2_decap_8 FILLER_27_431 ();
 sg13g2_decap_8 FILLER_27_438 ();
 sg13g2_decap_8 FILLER_27_445 ();
 sg13g2_decap_8 FILLER_27_452 ();
 sg13g2_decap_8 FILLER_27_459 ();
 sg13g2_decap_8 FILLER_27_466 ();
 sg13g2_decap_8 FILLER_27_473 ();
 sg13g2_decap_8 FILLER_27_480 ();
 sg13g2_decap_8 FILLER_27_487 ();
 sg13g2_decap_8 FILLER_27_494 ();
 sg13g2_decap_8 FILLER_27_501 ();
 sg13g2_decap_8 FILLER_27_508 ();
 sg13g2_decap_8 FILLER_27_515 ();
 sg13g2_decap_8 FILLER_27_522 ();
 sg13g2_decap_8 FILLER_27_529 ();
 sg13g2_decap_8 FILLER_27_536 ();
 sg13g2_decap_8 FILLER_27_543 ();
 sg13g2_decap_8 FILLER_27_550 ();
 sg13g2_decap_8 FILLER_27_557 ();
 sg13g2_decap_8 FILLER_27_564 ();
 sg13g2_decap_8 FILLER_27_571 ();
 sg13g2_decap_8 FILLER_27_578 ();
 sg13g2_decap_8 FILLER_27_585 ();
 sg13g2_decap_8 FILLER_27_592 ();
 sg13g2_decap_8 FILLER_27_599 ();
 sg13g2_decap_8 FILLER_27_606 ();
 sg13g2_decap_8 FILLER_27_613 ();
 sg13g2_decap_8 FILLER_27_620 ();
 sg13g2_decap_8 FILLER_27_627 ();
 sg13g2_decap_8 FILLER_27_634 ();
 sg13g2_decap_8 FILLER_27_641 ();
 sg13g2_decap_8 FILLER_27_648 ();
 sg13g2_decap_8 FILLER_27_655 ();
 sg13g2_decap_8 FILLER_27_662 ();
 sg13g2_decap_8 FILLER_27_669 ();
 sg13g2_decap_8 FILLER_27_676 ();
 sg13g2_decap_8 FILLER_27_683 ();
 sg13g2_decap_8 FILLER_27_690 ();
 sg13g2_decap_8 FILLER_27_697 ();
 sg13g2_decap_8 FILLER_27_704 ();
 sg13g2_decap_8 FILLER_27_711 ();
 sg13g2_decap_8 FILLER_27_718 ();
 sg13g2_decap_8 FILLER_27_725 ();
 sg13g2_decap_8 FILLER_27_732 ();
 sg13g2_decap_8 FILLER_27_739 ();
 sg13g2_decap_8 FILLER_27_746 ();
 sg13g2_decap_8 FILLER_27_753 ();
 sg13g2_decap_8 FILLER_27_760 ();
 sg13g2_decap_8 FILLER_27_767 ();
 sg13g2_decap_8 FILLER_27_774 ();
 sg13g2_decap_8 FILLER_27_781 ();
 sg13g2_decap_8 FILLER_27_788 ();
 sg13g2_decap_8 FILLER_27_795 ();
 sg13g2_decap_8 FILLER_27_802 ();
 sg13g2_decap_8 FILLER_27_809 ();
 sg13g2_decap_8 FILLER_27_816 ();
 sg13g2_decap_8 FILLER_27_823 ();
 sg13g2_decap_8 FILLER_27_830 ();
 sg13g2_decap_8 FILLER_27_837 ();
 sg13g2_decap_8 FILLER_27_844 ();
 sg13g2_decap_8 FILLER_27_851 ();
 sg13g2_decap_8 FILLER_27_858 ();
 sg13g2_decap_8 FILLER_27_865 ();
 sg13g2_decap_4 FILLER_27_872 ();
 sg13g2_fill_2 FILLER_27_876 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_fill_2 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_290 ();
 sg13g2_decap_8 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_decap_8 FILLER_28_311 ();
 sg13g2_decap_8 FILLER_28_318 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_decap_8 FILLER_28_332 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_28_424 ();
 sg13g2_decap_8 FILLER_28_431 ();
 sg13g2_decap_8 FILLER_28_438 ();
 sg13g2_decap_8 FILLER_28_445 ();
 sg13g2_decap_8 FILLER_28_452 ();
 sg13g2_decap_8 FILLER_28_459 ();
 sg13g2_decap_8 FILLER_28_466 ();
 sg13g2_decap_8 FILLER_28_473 ();
 sg13g2_decap_8 FILLER_28_480 ();
 sg13g2_decap_8 FILLER_28_487 ();
 sg13g2_decap_8 FILLER_28_494 ();
 sg13g2_decap_8 FILLER_28_501 ();
 sg13g2_decap_8 FILLER_28_508 ();
 sg13g2_decap_8 FILLER_28_515 ();
 sg13g2_decap_8 FILLER_28_522 ();
 sg13g2_decap_8 FILLER_28_529 ();
 sg13g2_decap_8 FILLER_28_536 ();
 sg13g2_decap_8 FILLER_28_543 ();
 sg13g2_decap_8 FILLER_28_550 ();
 sg13g2_decap_8 FILLER_28_557 ();
 sg13g2_decap_8 FILLER_28_564 ();
 sg13g2_decap_8 FILLER_28_571 ();
 sg13g2_decap_8 FILLER_28_578 ();
 sg13g2_decap_8 FILLER_28_585 ();
 sg13g2_decap_8 FILLER_28_592 ();
 sg13g2_decap_8 FILLER_28_599 ();
 sg13g2_decap_8 FILLER_28_606 ();
 sg13g2_decap_8 FILLER_28_613 ();
 sg13g2_decap_8 FILLER_28_620 ();
 sg13g2_decap_8 FILLER_28_627 ();
 sg13g2_decap_8 FILLER_28_634 ();
 sg13g2_decap_8 FILLER_28_641 ();
 sg13g2_decap_8 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_655 ();
 sg13g2_decap_8 FILLER_28_662 ();
 sg13g2_decap_8 FILLER_28_669 ();
 sg13g2_decap_8 FILLER_28_676 ();
 sg13g2_decap_8 FILLER_28_683 ();
 sg13g2_decap_8 FILLER_28_690 ();
 sg13g2_decap_8 FILLER_28_697 ();
 sg13g2_decap_8 FILLER_28_704 ();
 sg13g2_decap_8 FILLER_28_711 ();
 sg13g2_decap_8 FILLER_28_718 ();
 sg13g2_decap_8 FILLER_28_725 ();
 sg13g2_decap_8 FILLER_28_732 ();
 sg13g2_decap_8 FILLER_28_739 ();
 sg13g2_decap_8 FILLER_28_746 ();
 sg13g2_decap_8 FILLER_28_753 ();
 sg13g2_decap_8 FILLER_28_760 ();
 sg13g2_decap_8 FILLER_28_767 ();
 sg13g2_decap_8 FILLER_28_774 ();
 sg13g2_decap_8 FILLER_28_781 ();
 sg13g2_decap_8 FILLER_28_788 ();
 sg13g2_decap_8 FILLER_28_795 ();
 sg13g2_decap_8 FILLER_28_802 ();
 sg13g2_decap_8 FILLER_28_809 ();
 sg13g2_decap_8 FILLER_28_816 ();
 sg13g2_decap_8 FILLER_28_823 ();
 sg13g2_decap_8 FILLER_28_830 ();
 sg13g2_decap_8 FILLER_28_837 ();
 sg13g2_decap_8 FILLER_28_844 ();
 sg13g2_decap_8 FILLER_28_851 ();
 sg13g2_decap_8 FILLER_28_858 ();
 sg13g2_decap_8 FILLER_28_865 ();
 sg13g2_decap_4 FILLER_28_872 ();
 sg13g2_fill_2 FILLER_28_876 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_4 FILLER_29_266 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_decap_8 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_290 ();
 sg13g2_decap_8 FILLER_29_297 ();
 sg13g2_decap_8 FILLER_29_304 ();
 sg13g2_decap_8 FILLER_29_311 ();
 sg13g2_decap_8 FILLER_29_318 ();
 sg13g2_decap_8 FILLER_29_325 ();
 sg13g2_decap_8 FILLER_29_332 ();
 sg13g2_decap_8 FILLER_29_339 ();
 sg13g2_decap_8 FILLER_29_346 ();
 sg13g2_decap_8 FILLER_29_353 ();
 sg13g2_decap_8 FILLER_29_360 ();
 sg13g2_decap_8 FILLER_29_367 ();
 sg13g2_decap_8 FILLER_29_374 ();
 sg13g2_decap_8 FILLER_29_381 ();
 sg13g2_decap_8 FILLER_29_388 ();
 sg13g2_decap_4 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_490 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_decap_8 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_525 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_8 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_8 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_decap_8 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_29_847 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_decap_8 FILLER_29_861 ();
 sg13g2_decap_8 FILLER_29_868 ();
 sg13g2_fill_2 FILLER_29_875 ();
 sg13g2_fill_1 FILLER_29_877 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_12 ();
 sg13g2_decap_8 FILLER_30_19 ();
 sg13g2_decap_8 FILLER_30_26 ();
 sg13g2_decap_8 FILLER_30_33 ();
 sg13g2_decap_8 FILLER_30_40 ();
 sg13g2_decap_8 FILLER_30_47 ();
 sg13g2_decap_8 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_61 ();
 sg13g2_decap_8 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_75 ();
 sg13g2_decap_8 FILLER_30_82 ();
 sg13g2_decap_8 FILLER_30_89 ();
 sg13g2_fill_1 FILLER_30_96 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_decap_8 FILLER_30_856 ();
 sg13g2_decap_8 FILLER_30_863 ();
 sg13g2_decap_8 FILLER_30_870 ();
 sg13g2_fill_1 FILLER_30_877 ();
 sg13g2_decap_8 FILLER_31_26 ();
 sg13g2_decap_8 FILLER_31_33 ();
 sg13g2_decap_8 FILLER_31_40 ();
 sg13g2_decap_8 FILLER_31_47 ();
 sg13g2_decap_8 FILLER_31_54 ();
 sg13g2_decap_8 FILLER_31_61 ();
 sg13g2_decap_8 FILLER_31_68 ();
 sg13g2_decap_8 FILLER_31_75 ();
 sg13g2_decap_8 FILLER_31_82 ();
 sg13g2_decap_8 FILLER_31_89 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_decap_8 FILLER_31_807 ();
 sg13g2_decap_8 FILLER_31_814 ();
 sg13g2_decap_8 FILLER_31_821 ();
 sg13g2_decap_8 FILLER_31_828 ();
 sg13g2_decap_8 FILLER_31_835 ();
 sg13g2_decap_8 FILLER_31_842 ();
 sg13g2_decap_8 FILLER_31_849 ();
 sg13g2_decap_8 FILLER_31_856 ();
 sg13g2_decap_8 FILLER_31_863 ();
 sg13g2_decap_8 FILLER_31_870 ();
 sg13g2_fill_1 FILLER_31_877 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_15 ();
 sg13g2_decap_8 FILLER_32_22 ();
 sg13g2_decap_8 FILLER_32_29 ();
 sg13g2_decap_8 FILLER_32_36 ();
 sg13g2_decap_8 FILLER_32_43 ();
 sg13g2_decap_8 FILLER_32_50 ();
 sg13g2_decap_8 FILLER_32_57 ();
 sg13g2_decap_8 FILLER_32_64 ();
 sg13g2_decap_8 FILLER_32_71 ();
 sg13g2_decap_8 FILLER_32_78 ();
 sg13g2_decap_8 FILLER_32_85 ();
 sg13g2_decap_4 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_96 ();
 sg13g2_decap_8 FILLER_32_811 ();
 sg13g2_decap_8 FILLER_32_818 ();
 sg13g2_decap_8 FILLER_32_825 ();
 sg13g2_decap_8 FILLER_32_832 ();
 sg13g2_decap_8 FILLER_32_839 ();
 sg13g2_decap_8 FILLER_32_846 ();
 sg13g2_decap_8 FILLER_32_853 ();
 sg13g2_decap_8 FILLER_32_860 ();
 sg13g2_decap_8 FILLER_32_867 ();
 sg13g2_decap_4 FILLER_32_874 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_4 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_95 ();
 sg13g2_decap_8 FILLER_33_811 ();
 sg13g2_decap_8 FILLER_33_818 ();
 sg13g2_decap_8 FILLER_33_825 ();
 sg13g2_decap_8 FILLER_33_832 ();
 sg13g2_decap_8 FILLER_33_839 ();
 sg13g2_decap_8 FILLER_33_846 ();
 sg13g2_decap_8 FILLER_33_853 ();
 sg13g2_decap_8 FILLER_33_860 ();
 sg13g2_decap_8 FILLER_33_867 ();
 sg13g2_decap_4 FILLER_33_874 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_12 ();
 sg13g2_decap_8 FILLER_34_19 ();
 sg13g2_decap_8 FILLER_34_26 ();
 sg13g2_decap_8 FILLER_34_33 ();
 sg13g2_decap_8 FILLER_34_40 ();
 sg13g2_decap_8 FILLER_34_47 ();
 sg13g2_decap_8 FILLER_34_54 ();
 sg13g2_decap_8 FILLER_34_61 ();
 sg13g2_decap_8 FILLER_34_68 ();
 sg13g2_decap_8 FILLER_34_75 ();
 sg13g2_decap_8 FILLER_34_82 ();
 sg13g2_decap_8 FILLER_34_89 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_811 ();
 sg13g2_decap_8 FILLER_34_818 ();
 sg13g2_decap_8 FILLER_34_825 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_decap_8 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_34_867 ();
 sg13g2_decap_4 FILLER_34_874 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_12 ();
 sg13g2_decap_8 FILLER_35_19 ();
 sg13g2_decap_8 FILLER_35_26 ();
 sg13g2_decap_8 FILLER_35_33 ();
 sg13g2_decap_8 FILLER_35_40 ();
 sg13g2_decap_8 FILLER_35_47 ();
 sg13g2_decap_8 FILLER_35_54 ();
 sg13g2_decap_8 FILLER_35_61 ();
 sg13g2_decap_8 FILLER_35_68 ();
 sg13g2_decap_8 FILLER_35_75 ();
 sg13g2_decap_8 FILLER_35_82 ();
 sg13g2_decap_8 FILLER_35_89 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_decap_8 FILLER_35_811 ();
 sg13g2_decap_8 FILLER_35_818 ();
 sg13g2_decap_8 FILLER_35_825 ();
 sg13g2_decap_8 FILLER_35_832 ();
 sg13g2_decap_8 FILLER_35_839 ();
 sg13g2_decap_8 FILLER_35_846 ();
 sg13g2_decap_8 FILLER_35_853 ();
 sg13g2_decap_8 FILLER_35_860 ();
 sg13g2_decap_8 FILLER_35_867 ();
 sg13g2_decap_4 FILLER_35_874 ();
 sg13g2_decap_8 FILLER_36_26 ();
 sg13g2_decap_8 FILLER_36_33 ();
 sg13g2_decap_8 FILLER_36_40 ();
 sg13g2_decap_8 FILLER_36_47 ();
 sg13g2_decap_8 FILLER_36_54 ();
 sg13g2_decap_8 FILLER_36_61 ();
 sg13g2_decap_8 FILLER_36_68 ();
 sg13g2_decap_8 FILLER_36_75 ();
 sg13g2_decap_8 FILLER_36_82 ();
 sg13g2_decap_8 FILLER_36_89 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_decap_8 FILLER_36_811 ();
 sg13g2_decap_8 FILLER_36_818 ();
 sg13g2_decap_8 FILLER_36_825 ();
 sg13g2_decap_8 FILLER_36_832 ();
 sg13g2_decap_8 FILLER_36_839 ();
 sg13g2_decap_8 FILLER_36_846 ();
 sg13g2_decap_8 FILLER_36_853 ();
 sg13g2_decap_8 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_36_867 ();
 sg13g2_decap_4 FILLER_36_874 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_4 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_15 ();
 sg13g2_decap_8 FILLER_37_22 ();
 sg13g2_decap_8 FILLER_37_29 ();
 sg13g2_decap_8 FILLER_37_36 ();
 sg13g2_decap_8 FILLER_37_43 ();
 sg13g2_decap_8 FILLER_37_50 ();
 sg13g2_decap_8 FILLER_37_57 ();
 sg13g2_decap_8 FILLER_37_64 ();
 sg13g2_decap_8 FILLER_37_71 ();
 sg13g2_decap_8 FILLER_37_78 ();
 sg13g2_decap_8 FILLER_37_85 ();
 sg13g2_decap_4 FILLER_37_92 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_decap_8 FILLER_37_811 ();
 sg13g2_decap_8 FILLER_37_818 ();
 sg13g2_decap_8 FILLER_37_825 ();
 sg13g2_decap_8 FILLER_37_832 ();
 sg13g2_decap_8 FILLER_37_839 ();
 sg13g2_decap_8 FILLER_37_846 ();
 sg13g2_decap_8 FILLER_37_853 ();
 sg13g2_decap_8 FILLER_37_860 ();
 sg13g2_decap_8 FILLER_37_867 ();
 sg13g2_decap_4 FILLER_37_874 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_95 ();
 sg13g2_decap_8 FILLER_38_811 ();
 sg13g2_decap_8 FILLER_38_818 ();
 sg13g2_decap_8 FILLER_38_825 ();
 sg13g2_decap_8 FILLER_38_832 ();
 sg13g2_decap_8 FILLER_38_839 ();
 sg13g2_decap_8 FILLER_38_846 ();
 sg13g2_decap_8 FILLER_38_853 ();
 sg13g2_decap_8 FILLER_38_860 ();
 sg13g2_decap_8 FILLER_38_867 ();
 sg13g2_decap_4 FILLER_38_874 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_4 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_4 FILLER_39_91 ();
 sg13g2_fill_2 FILLER_39_95 ();
 sg13g2_decap_8 FILLER_39_811 ();
 sg13g2_decap_8 FILLER_39_818 ();
 sg13g2_decap_8 FILLER_39_825 ();
 sg13g2_decap_8 FILLER_39_832 ();
 sg13g2_decap_8 FILLER_39_839 ();
 sg13g2_decap_8 FILLER_39_846 ();
 sg13g2_decap_8 FILLER_39_853 ();
 sg13g2_decap_8 FILLER_39_860 ();
 sg13g2_decap_8 FILLER_39_867 ();
 sg13g2_decap_4 FILLER_39_874 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_4 FILLER_40_91 ();
 sg13g2_fill_2 FILLER_40_95 ();
 sg13g2_decap_8 FILLER_40_811 ();
 sg13g2_decap_8 FILLER_40_818 ();
 sg13g2_decap_8 FILLER_40_825 ();
 sg13g2_decap_8 FILLER_40_832 ();
 sg13g2_decap_8 FILLER_40_839 ();
 sg13g2_decap_8 FILLER_40_846 ();
 sg13g2_decap_8 FILLER_40_853 ();
 sg13g2_decap_8 FILLER_40_860 ();
 sg13g2_decap_8 FILLER_40_867 ();
 sg13g2_decap_4 FILLER_40_874 ();
 sg13g2_fill_2 FILLER_41_3 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_4 FILLER_41_91 ();
 sg13g2_fill_2 FILLER_41_95 ();
 sg13g2_decap_8 FILLER_41_811 ();
 sg13g2_decap_8 FILLER_41_818 ();
 sg13g2_decap_8 FILLER_41_825 ();
 sg13g2_decap_8 FILLER_41_832 ();
 sg13g2_decap_8 FILLER_41_839 ();
 sg13g2_decap_8 FILLER_41_846 ();
 sg13g2_decap_8 FILLER_41_853 ();
 sg13g2_decap_8 FILLER_41_860 ();
 sg13g2_decap_8 FILLER_41_867 ();
 sg13g2_decap_4 FILLER_41_874 ();
 sg13g2_decap_8 FILLER_42_12 ();
 sg13g2_decap_8 FILLER_42_19 ();
 sg13g2_decap_8 FILLER_42_26 ();
 sg13g2_decap_8 FILLER_42_33 ();
 sg13g2_decap_8 FILLER_42_40 ();
 sg13g2_decap_8 FILLER_42_47 ();
 sg13g2_decap_8 FILLER_42_54 ();
 sg13g2_decap_8 FILLER_42_61 ();
 sg13g2_decap_8 FILLER_42_68 ();
 sg13g2_decap_8 FILLER_42_75 ();
 sg13g2_decap_8 FILLER_42_82 ();
 sg13g2_decap_8 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_96 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_846 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_decap_8 FILLER_42_860 ();
 sg13g2_decap_8 FILLER_42_867 ();
 sg13g2_decap_4 FILLER_42_874 ();
 sg13g2_decap_8 FILLER_43_32 ();
 sg13g2_decap_8 FILLER_43_39 ();
 sg13g2_decap_8 FILLER_43_46 ();
 sg13g2_decap_8 FILLER_43_53 ();
 sg13g2_decap_8 FILLER_43_60 ();
 sg13g2_decap_8 FILLER_43_67 ();
 sg13g2_decap_8 FILLER_43_74 ();
 sg13g2_decap_8 FILLER_43_81 ();
 sg13g2_decap_8 FILLER_43_88 ();
 sg13g2_fill_2 FILLER_43_95 ();
 sg13g2_decap_8 FILLER_43_811 ();
 sg13g2_decap_8 FILLER_43_818 ();
 sg13g2_decap_8 FILLER_43_825 ();
 sg13g2_decap_8 FILLER_43_832 ();
 sg13g2_decap_8 FILLER_43_839 ();
 sg13g2_decap_8 FILLER_43_846 ();
 sg13g2_decap_8 FILLER_43_853 ();
 sg13g2_decap_8 FILLER_43_860 ();
 sg13g2_decap_8 FILLER_43_867 ();
 sg13g2_decap_4 FILLER_43_874 ();
 sg13g2_decap_4 FILLER_44_6 ();
 sg13g2_fill_1 FILLER_44_10 ();
 sg13g2_decap_8 FILLER_44_15 ();
 sg13g2_decap_8 FILLER_44_22 ();
 sg13g2_decap_8 FILLER_44_29 ();
 sg13g2_decap_8 FILLER_44_36 ();
 sg13g2_decap_8 FILLER_44_43 ();
 sg13g2_decap_8 FILLER_44_50 ();
 sg13g2_decap_8 FILLER_44_57 ();
 sg13g2_decap_8 FILLER_44_64 ();
 sg13g2_decap_8 FILLER_44_71 ();
 sg13g2_decap_8 FILLER_44_78 ();
 sg13g2_decap_8 FILLER_44_85 ();
 sg13g2_decap_4 FILLER_44_92 ();
 sg13g2_fill_1 FILLER_44_96 ();
 sg13g2_decap_8 FILLER_44_807 ();
 sg13g2_decap_8 FILLER_44_814 ();
 sg13g2_decap_8 FILLER_44_821 ();
 sg13g2_decap_8 FILLER_44_828 ();
 sg13g2_decap_8 FILLER_44_835 ();
 sg13g2_decap_8 FILLER_44_842 ();
 sg13g2_decap_8 FILLER_44_849 ();
 sg13g2_decap_8 FILLER_44_856 ();
 sg13g2_decap_8 FILLER_44_863 ();
 sg13g2_decap_8 FILLER_44_870 ();
 sg13g2_fill_1 FILLER_44_877 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_4 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_4 FILLER_45_91 ();
 sg13g2_fill_2 FILLER_45_95 ();
 sg13g2_decap_8 FILLER_45_807 ();
 sg13g2_decap_8 FILLER_45_814 ();
 sg13g2_decap_8 FILLER_45_821 ();
 sg13g2_decap_8 FILLER_45_828 ();
 sg13g2_decap_8 FILLER_45_835 ();
 sg13g2_decap_8 FILLER_45_842 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_decap_8 FILLER_45_856 ();
 sg13g2_decap_8 FILLER_45_863 ();
 sg13g2_decap_8 FILLER_45_870 ();
 sg13g2_fill_1 FILLER_45_877 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_decap_8 FILLER_46_16 ();
 sg13g2_decap_8 FILLER_46_23 ();
 sg13g2_decap_8 FILLER_46_30 ();
 sg13g2_decap_8 FILLER_46_37 ();
 sg13g2_decap_8 FILLER_46_44 ();
 sg13g2_decap_8 FILLER_46_51 ();
 sg13g2_decap_8 FILLER_46_58 ();
 sg13g2_decap_8 FILLER_46_65 ();
 sg13g2_decap_8 FILLER_46_72 ();
 sg13g2_decap_8 FILLER_46_79 ();
 sg13g2_decap_8 FILLER_46_86 ();
 sg13g2_decap_4 FILLER_46_93 ();
 sg13g2_decap_8 FILLER_46_815 ();
 sg13g2_decap_8 FILLER_46_822 ();
 sg13g2_decap_8 FILLER_46_829 ();
 sg13g2_decap_8 FILLER_46_836 ();
 sg13g2_decap_8 FILLER_46_843 ();
 sg13g2_decap_8 FILLER_46_850 ();
 sg13g2_decap_8 FILLER_46_857 ();
 sg13g2_decap_8 FILLER_46_864 ();
 sg13g2_decap_8 FILLER_46_871 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_4 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_95 ();
 sg13g2_decap_8 FILLER_47_807 ();
 sg13g2_decap_8 FILLER_47_814 ();
 sg13g2_decap_8 FILLER_47_821 ();
 sg13g2_decap_8 FILLER_47_828 ();
 sg13g2_decap_8 FILLER_47_835 ();
 sg13g2_decap_8 FILLER_47_842 ();
 sg13g2_decap_8 FILLER_47_849 ();
 sg13g2_decap_8 FILLER_47_856 ();
 sg13g2_decap_8 FILLER_47_863 ();
 sg13g2_decap_8 FILLER_47_870 ();
 sg13g2_fill_1 FILLER_47_877 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_4 ();
 sg13g2_decap_8 FILLER_48_16 ();
 sg13g2_decap_8 FILLER_48_23 ();
 sg13g2_decap_8 FILLER_48_30 ();
 sg13g2_decap_8 FILLER_48_37 ();
 sg13g2_decap_8 FILLER_48_44 ();
 sg13g2_decap_8 FILLER_48_51 ();
 sg13g2_decap_8 FILLER_48_58 ();
 sg13g2_decap_8 FILLER_48_65 ();
 sg13g2_decap_8 FILLER_48_72 ();
 sg13g2_decap_8 FILLER_48_79 ();
 sg13g2_decap_8 FILLER_48_86 ();
 sg13g2_decap_4 FILLER_48_93 ();
 sg13g2_decap_8 FILLER_48_815 ();
 sg13g2_decap_8 FILLER_48_822 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_decap_8 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_850 ();
 sg13g2_decap_8 FILLER_48_857 ();
 sg13g2_decap_8 FILLER_48_864 ();
 sg13g2_decap_8 FILLER_48_871 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_4 FILLER_49_91 ();
 sg13g2_fill_2 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_814 ();
 sg13g2_decap_8 FILLER_49_821 ();
 sg13g2_decap_8 FILLER_49_828 ();
 sg13g2_decap_8 FILLER_49_835 ();
 sg13g2_decap_8 FILLER_49_842 ();
 sg13g2_decap_8 FILLER_49_849 ();
 sg13g2_decap_8 FILLER_49_856 ();
 sg13g2_decap_8 FILLER_49_863 ();
 sg13g2_decap_8 FILLER_49_870 ();
 sg13g2_fill_1 FILLER_49_877 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_4 FILLER_50_91 ();
 sg13g2_fill_2 FILLER_50_95 ();
 sg13g2_decap_8 FILLER_50_831 ();
 sg13g2_decap_8 FILLER_50_838 ();
 sg13g2_decap_8 FILLER_50_845 ();
 sg13g2_decap_8 FILLER_50_852 ();
 sg13g2_decap_8 FILLER_50_859 ();
 sg13g2_decap_8 FILLER_50_866 ();
 sg13g2_decap_4 FILLER_50_873 ();
 sg13g2_fill_1 FILLER_50_877 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_4 FILLER_51_91 ();
 sg13g2_fill_2 FILLER_51_95 ();
 sg13g2_decap_8 FILLER_51_819 ();
 sg13g2_decap_8 FILLER_51_826 ();
 sg13g2_decap_8 FILLER_51_833 ();
 sg13g2_decap_8 FILLER_51_840 ();
 sg13g2_decap_8 FILLER_51_847 ();
 sg13g2_decap_8 FILLER_51_854 ();
 sg13g2_decap_8 FILLER_51_861 ();
 sg13g2_decap_8 FILLER_51_868 ();
 sg13g2_fill_2 FILLER_51_875 ();
 sg13g2_fill_1 FILLER_51_877 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_4 FILLER_52_91 ();
 sg13g2_fill_2 FILLER_52_95 ();
 sg13g2_decap_8 FILLER_52_815 ();
 sg13g2_decap_8 FILLER_52_822 ();
 sg13g2_decap_8 FILLER_52_829 ();
 sg13g2_decap_8 FILLER_52_836 ();
 sg13g2_decap_8 FILLER_52_843 ();
 sg13g2_decap_8 FILLER_52_850 ();
 sg13g2_decap_8 FILLER_52_857 ();
 sg13g2_decap_8 FILLER_52_864 ();
 sg13g2_decap_8 FILLER_52_871 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_4 FILLER_53_91 ();
 sg13g2_fill_2 FILLER_53_95 ();
 sg13g2_decap_8 FILLER_53_811 ();
 sg13g2_decap_8 FILLER_53_818 ();
 sg13g2_decap_8 FILLER_53_825 ();
 sg13g2_decap_8 FILLER_53_832 ();
 sg13g2_decap_8 FILLER_53_839 ();
 sg13g2_decap_8 FILLER_53_846 ();
 sg13g2_decap_8 FILLER_53_853 ();
 sg13g2_decap_8 FILLER_53_860 ();
 sg13g2_decap_8 FILLER_53_867 ();
 sg13g2_decap_4 FILLER_53_874 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_4 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_95 ();
 sg13g2_decap_8 FILLER_54_815 ();
 sg13g2_decap_8 FILLER_54_822 ();
 sg13g2_decap_8 FILLER_54_829 ();
 sg13g2_decap_8 FILLER_54_836 ();
 sg13g2_decap_8 FILLER_54_843 ();
 sg13g2_decap_8 FILLER_54_850 ();
 sg13g2_decap_8 FILLER_54_857 ();
 sg13g2_decap_8 FILLER_54_864 ();
 sg13g2_decap_8 FILLER_54_871 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_4 FILLER_55_91 ();
 sg13g2_fill_2 FILLER_55_95 ();
 sg13g2_decap_8 FILLER_55_807 ();
 sg13g2_decap_8 FILLER_55_814 ();
 sg13g2_decap_8 FILLER_55_821 ();
 sg13g2_decap_8 FILLER_55_828 ();
 sg13g2_decap_8 FILLER_55_835 ();
 sg13g2_decap_8 FILLER_55_842 ();
 sg13g2_decap_8 FILLER_55_849 ();
 sg13g2_decap_8 FILLER_55_856 ();
 sg13g2_decap_8 FILLER_55_863 ();
 sg13g2_decap_8 FILLER_55_870 ();
 sg13g2_fill_1 FILLER_55_877 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_4 FILLER_56_91 ();
 sg13g2_fill_2 FILLER_56_95 ();
 sg13g2_decap_8 FILLER_56_807 ();
 sg13g2_decap_8 FILLER_56_814 ();
 sg13g2_decap_8 FILLER_56_821 ();
 sg13g2_decap_8 FILLER_56_828 ();
 sg13g2_decap_8 FILLER_56_835 ();
 sg13g2_decap_8 FILLER_56_842 ();
 sg13g2_decap_8 FILLER_56_849 ();
 sg13g2_decap_8 FILLER_56_856 ();
 sg13g2_decap_8 FILLER_56_863 ();
 sg13g2_decap_8 FILLER_56_870 ();
 sg13g2_fill_1 FILLER_56_877 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_4 FILLER_57_91 ();
 sg13g2_fill_2 FILLER_57_95 ();
 sg13g2_decap_8 FILLER_57_807 ();
 sg13g2_decap_8 FILLER_57_814 ();
 sg13g2_decap_8 FILLER_57_821 ();
 sg13g2_decap_8 FILLER_57_828 ();
 sg13g2_decap_8 FILLER_57_835 ();
 sg13g2_decap_8 FILLER_57_842 ();
 sg13g2_decap_8 FILLER_57_849 ();
 sg13g2_decap_8 FILLER_57_856 ();
 sg13g2_decap_8 FILLER_57_863 ();
 sg13g2_decap_8 FILLER_57_870 ();
 sg13g2_fill_1 FILLER_57_877 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_4 FILLER_58_91 ();
 sg13g2_fill_2 FILLER_58_95 ();
 sg13g2_decap_8 FILLER_58_815 ();
 sg13g2_decap_8 FILLER_58_822 ();
 sg13g2_decap_8 FILLER_58_829 ();
 sg13g2_decap_8 FILLER_58_836 ();
 sg13g2_decap_8 FILLER_58_843 ();
 sg13g2_decap_8 FILLER_58_850 ();
 sg13g2_decap_8 FILLER_58_857 ();
 sg13g2_decap_8 FILLER_58_864 ();
 sg13g2_decap_8 FILLER_58_871 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_4 FILLER_59_91 ();
 sg13g2_fill_2 FILLER_59_95 ();
 sg13g2_decap_8 FILLER_59_807 ();
 sg13g2_decap_8 FILLER_59_814 ();
 sg13g2_decap_8 FILLER_59_821 ();
 sg13g2_decap_8 FILLER_59_828 ();
 sg13g2_decap_8 FILLER_59_835 ();
 sg13g2_decap_8 FILLER_59_842 ();
 sg13g2_decap_8 FILLER_59_849 ();
 sg13g2_decap_8 FILLER_59_856 ();
 sg13g2_decap_8 FILLER_59_863 ();
 sg13g2_decap_8 FILLER_59_870 ();
 sg13g2_fill_1 FILLER_59_877 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_4 FILLER_60_91 ();
 sg13g2_fill_2 FILLER_60_95 ();
 sg13g2_decap_8 FILLER_60_811 ();
 sg13g2_decap_8 FILLER_60_818 ();
 sg13g2_decap_8 FILLER_60_825 ();
 sg13g2_decap_8 FILLER_60_832 ();
 sg13g2_decap_8 FILLER_60_839 ();
 sg13g2_decap_8 FILLER_60_846 ();
 sg13g2_decap_8 FILLER_60_853 ();
 sg13g2_decap_8 FILLER_60_860 ();
 sg13g2_decap_8 FILLER_60_867 ();
 sg13g2_decap_4 FILLER_60_874 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_11 ();
 sg13g2_decap_8 FILLER_61_18 ();
 sg13g2_decap_8 FILLER_61_25 ();
 sg13g2_decap_8 FILLER_61_32 ();
 sg13g2_decap_8 FILLER_61_39 ();
 sg13g2_decap_8 FILLER_61_46 ();
 sg13g2_decap_8 FILLER_61_53 ();
 sg13g2_decap_8 FILLER_61_60 ();
 sg13g2_decap_8 FILLER_61_67 ();
 sg13g2_decap_8 FILLER_61_74 ();
 sg13g2_decap_8 FILLER_61_81 ();
 sg13g2_decap_8 FILLER_61_88 ();
 sg13g2_fill_2 FILLER_61_95 ();
 sg13g2_decap_8 FILLER_61_815 ();
 sg13g2_decap_8 FILLER_61_822 ();
 sg13g2_decap_8 FILLER_61_829 ();
 sg13g2_decap_8 FILLER_61_836 ();
 sg13g2_decap_8 FILLER_61_843 ();
 sg13g2_decap_8 FILLER_61_850 ();
 sg13g2_decap_8 FILLER_61_857 ();
 sg13g2_decap_8 FILLER_61_864 ();
 sg13g2_decap_8 FILLER_61_871 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_4 FILLER_62_91 ();
 sg13g2_fill_2 FILLER_62_95 ();
 sg13g2_decap_8 FILLER_62_807 ();
 sg13g2_decap_8 FILLER_62_814 ();
 sg13g2_decap_8 FILLER_62_821 ();
 sg13g2_decap_8 FILLER_62_828 ();
 sg13g2_decap_8 FILLER_62_835 ();
 sg13g2_decap_8 FILLER_62_842 ();
 sg13g2_decap_8 FILLER_62_849 ();
 sg13g2_decap_8 FILLER_62_856 ();
 sg13g2_decap_8 FILLER_62_863 ();
 sg13g2_decap_8 FILLER_62_870 ();
 sg13g2_fill_1 FILLER_62_877 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_4 FILLER_63_91 ();
 sg13g2_fill_2 FILLER_63_95 ();
 sg13g2_decap_8 FILLER_63_811 ();
 sg13g2_decap_8 FILLER_63_818 ();
 sg13g2_decap_8 FILLER_63_825 ();
 sg13g2_decap_8 FILLER_63_832 ();
 sg13g2_decap_8 FILLER_63_839 ();
 sg13g2_decap_8 FILLER_63_846 ();
 sg13g2_decap_8 FILLER_63_853 ();
 sg13g2_decap_8 FILLER_63_860 ();
 sg13g2_decap_8 FILLER_63_867 ();
 sg13g2_decap_4 FILLER_63_874 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_4 FILLER_64_91 ();
 sg13g2_fill_2 FILLER_64_95 ();
 sg13g2_decap_8 FILLER_64_815 ();
 sg13g2_decap_8 FILLER_64_822 ();
 sg13g2_decap_8 FILLER_64_829 ();
 sg13g2_decap_8 FILLER_64_836 ();
 sg13g2_decap_8 FILLER_64_843 ();
 sg13g2_decap_8 FILLER_64_850 ();
 sg13g2_decap_8 FILLER_64_857 ();
 sg13g2_decap_8 FILLER_64_864 ();
 sg13g2_decap_8 FILLER_64_871 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_4 FILLER_65_91 ();
 sg13g2_fill_2 FILLER_65_95 ();
 sg13g2_decap_8 FILLER_65_811 ();
 sg13g2_decap_8 FILLER_65_818 ();
 sg13g2_decap_8 FILLER_65_825 ();
 sg13g2_decap_8 FILLER_65_832 ();
 sg13g2_decap_8 FILLER_65_839 ();
 sg13g2_decap_8 FILLER_65_846 ();
 sg13g2_decap_8 FILLER_65_853 ();
 sg13g2_decap_8 FILLER_65_860 ();
 sg13g2_decap_8 FILLER_65_867 ();
 sg13g2_decap_4 FILLER_65_874 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_4 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_95 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_8 FILLER_66_856 ();
 sg13g2_decap_8 FILLER_66_863 ();
 sg13g2_decap_8 FILLER_66_870 ();
 sg13g2_fill_1 FILLER_66_877 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_4 FILLER_67_91 ();
 sg13g2_fill_2 FILLER_67_95 ();
 sg13g2_decap_8 FILLER_67_815 ();
 sg13g2_decap_8 FILLER_67_822 ();
 sg13g2_decap_8 FILLER_67_829 ();
 sg13g2_decap_8 FILLER_67_836 ();
 sg13g2_decap_8 FILLER_67_843 ();
 sg13g2_decap_8 FILLER_67_850 ();
 sg13g2_decap_8 FILLER_67_857 ();
 sg13g2_decap_8 FILLER_67_864 ();
 sg13g2_decap_8 FILLER_67_871 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_4 FILLER_68_91 ();
 sg13g2_fill_2 FILLER_68_95 ();
 sg13g2_decap_8 FILLER_68_811 ();
 sg13g2_decap_8 FILLER_68_818 ();
 sg13g2_decap_8 FILLER_68_825 ();
 sg13g2_decap_8 FILLER_68_832 ();
 sg13g2_decap_8 FILLER_68_839 ();
 sg13g2_decap_8 FILLER_68_846 ();
 sg13g2_decap_8 FILLER_68_853 ();
 sg13g2_decap_8 FILLER_68_860 ();
 sg13g2_decap_8 FILLER_68_867 ();
 sg13g2_decap_4 FILLER_68_874 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_4 FILLER_69_91 ();
 sg13g2_fill_2 FILLER_69_95 ();
 sg13g2_decap_8 FILLER_69_807 ();
 sg13g2_decap_8 FILLER_69_814 ();
 sg13g2_decap_8 FILLER_69_821 ();
 sg13g2_decap_8 FILLER_69_828 ();
 sg13g2_decap_8 FILLER_69_835 ();
 sg13g2_decap_8 FILLER_69_842 ();
 sg13g2_decap_8 FILLER_69_849 ();
 sg13g2_decap_8 FILLER_69_856 ();
 sg13g2_decap_8 FILLER_69_863 ();
 sg13g2_decap_8 FILLER_69_870 ();
 sg13g2_fill_1 FILLER_69_877 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_4 FILLER_70_91 ();
 sg13g2_fill_2 FILLER_70_95 ();
 sg13g2_decap_8 FILLER_70_807 ();
 sg13g2_decap_8 FILLER_70_814 ();
 sg13g2_decap_8 FILLER_70_821 ();
 sg13g2_decap_8 FILLER_70_828 ();
 sg13g2_decap_8 FILLER_70_835 ();
 sg13g2_decap_8 FILLER_70_842 ();
 sg13g2_decap_8 FILLER_70_849 ();
 sg13g2_decap_8 FILLER_70_856 ();
 sg13g2_decap_8 FILLER_70_863 ();
 sg13g2_decap_8 FILLER_70_870 ();
 sg13g2_fill_1 FILLER_70_877 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_203 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_245 ();
 sg13g2_decap_8 FILLER_71_252 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_decap_8 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_273 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_decap_8 FILLER_71_315 ();
 sg13g2_decap_8 FILLER_71_322 ();
 sg13g2_decap_8 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_decap_8 FILLER_71_350 ();
 sg13g2_decap_8 FILLER_71_357 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_4 FILLER_71_385 ();
 sg13g2_fill_2 FILLER_71_389 ();
 sg13g2_decap_8 FILLER_71_436 ();
 sg13g2_decap_8 FILLER_71_443 ();
 sg13g2_decap_8 FILLER_71_450 ();
 sg13g2_decap_8 FILLER_71_457 ();
 sg13g2_decap_8 FILLER_71_464 ();
 sg13g2_decap_8 FILLER_71_471 ();
 sg13g2_decap_8 FILLER_71_478 ();
 sg13g2_decap_8 FILLER_71_485 ();
 sg13g2_decap_8 FILLER_71_492 ();
 sg13g2_decap_8 FILLER_71_499 ();
 sg13g2_decap_8 FILLER_71_506 ();
 sg13g2_decap_8 FILLER_71_513 ();
 sg13g2_decap_8 FILLER_71_520 ();
 sg13g2_decap_8 FILLER_71_527 ();
 sg13g2_decap_8 FILLER_71_534 ();
 sg13g2_decap_8 FILLER_71_541 ();
 sg13g2_decap_8 FILLER_71_548 ();
 sg13g2_decap_8 FILLER_71_555 ();
 sg13g2_decap_8 FILLER_71_562 ();
 sg13g2_decap_8 FILLER_71_569 ();
 sg13g2_decap_8 FILLER_71_576 ();
 sg13g2_decap_8 FILLER_71_583 ();
 sg13g2_decap_8 FILLER_71_590 ();
 sg13g2_decap_8 FILLER_71_597 ();
 sg13g2_decap_8 FILLER_71_604 ();
 sg13g2_decap_8 FILLER_71_611 ();
 sg13g2_decap_8 FILLER_71_618 ();
 sg13g2_decap_8 FILLER_71_625 ();
 sg13g2_decap_8 FILLER_71_632 ();
 sg13g2_decap_8 FILLER_71_639 ();
 sg13g2_decap_8 FILLER_71_646 ();
 sg13g2_decap_8 FILLER_71_653 ();
 sg13g2_decap_8 FILLER_71_660 ();
 sg13g2_decap_8 FILLER_71_667 ();
 sg13g2_decap_8 FILLER_71_674 ();
 sg13g2_decap_8 FILLER_71_681 ();
 sg13g2_decap_8 FILLER_71_688 ();
 sg13g2_decap_8 FILLER_71_695 ();
 sg13g2_decap_8 FILLER_71_702 ();
 sg13g2_decap_8 FILLER_71_709 ();
 sg13g2_decap_8 FILLER_71_716 ();
 sg13g2_decap_8 FILLER_71_723 ();
 sg13g2_decap_8 FILLER_71_730 ();
 sg13g2_decap_8 FILLER_71_737 ();
 sg13g2_decap_8 FILLER_71_744 ();
 sg13g2_decap_8 FILLER_71_751 ();
 sg13g2_decap_8 FILLER_71_758 ();
 sg13g2_decap_8 FILLER_71_765 ();
 sg13g2_decap_8 FILLER_71_772 ();
 sg13g2_decap_8 FILLER_71_779 ();
 sg13g2_decap_8 FILLER_71_786 ();
 sg13g2_decap_8 FILLER_71_793 ();
 sg13g2_decap_8 FILLER_71_800 ();
 sg13g2_decap_8 FILLER_71_807 ();
 sg13g2_decap_8 FILLER_71_814 ();
 sg13g2_decap_8 FILLER_71_821 ();
 sg13g2_decap_8 FILLER_71_828 ();
 sg13g2_decap_8 FILLER_71_835 ();
 sg13g2_decap_8 FILLER_71_842 ();
 sg13g2_decap_8 FILLER_71_849 ();
 sg13g2_decap_8 FILLER_71_856 ();
 sg13g2_decap_8 FILLER_71_863 ();
 sg13g2_decap_8 FILLER_71_870 ();
 sg13g2_fill_1 FILLER_71_877 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_252 ();
 sg13g2_decap_8 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_280 ();
 sg13g2_decap_8 FILLER_72_287 ();
 sg13g2_decap_8 FILLER_72_294 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_8 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_343 ();
 sg13g2_decap_8 FILLER_72_350 ();
 sg13g2_decap_8 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_fill_2 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_420 ();
 sg13g2_decap_8 FILLER_72_433 ();
 sg13g2_decap_8 FILLER_72_440 ();
 sg13g2_decap_8 FILLER_72_447 ();
 sg13g2_decap_8 FILLER_72_454 ();
 sg13g2_decap_8 FILLER_72_461 ();
 sg13g2_decap_8 FILLER_72_468 ();
 sg13g2_decap_8 FILLER_72_475 ();
 sg13g2_decap_8 FILLER_72_482 ();
 sg13g2_decap_8 FILLER_72_489 ();
 sg13g2_decap_8 FILLER_72_496 ();
 sg13g2_decap_8 FILLER_72_503 ();
 sg13g2_decap_8 FILLER_72_510 ();
 sg13g2_decap_8 FILLER_72_517 ();
 sg13g2_decap_8 FILLER_72_524 ();
 sg13g2_decap_8 FILLER_72_531 ();
 sg13g2_decap_8 FILLER_72_538 ();
 sg13g2_decap_8 FILLER_72_545 ();
 sg13g2_decap_8 FILLER_72_552 ();
 sg13g2_decap_8 FILLER_72_559 ();
 sg13g2_decap_8 FILLER_72_566 ();
 sg13g2_decap_8 FILLER_72_573 ();
 sg13g2_decap_8 FILLER_72_580 ();
 sg13g2_decap_8 FILLER_72_587 ();
 sg13g2_decap_8 FILLER_72_594 ();
 sg13g2_decap_8 FILLER_72_601 ();
 sg13g2_decap_8 FILLER_72_608 ();
 sg13g2_decap_8 FILLER_72_615 ();
 sg13g2_decap_8 FILLER_72_622 ();
 sg13g2_decap_8 FILLER_72_629 ();
 sg13g2_decap_8 FILLER_72_636 ();
 sg13g2_decap_8 FILLER_72_643 ();
 sg13g2_decap_8 FILLER_72_650 ();
 sg13g2_decap_8 FILLER_72_657 ();
 sg13g2_decap_8 FILLER_72_664 ();
 sg13g2_decap_8 FILLER_72_671 ();
 sg13g2_decap_8 FILLER_72_678 ();
 sg13g2_decap_8 FILLER_72_685 ();
 sg13g2_decap_8 FILLER_72_692 ();
 sg13g2_decap_8 FILLER_72_699 ();
 sg13g2_decap_8 FILLER_72_706 ();
 sg13g2_decap_8 FILLER_72_713 ();
 sg13g2_decap_8 FILLER_72_720 ();
 sg13g2_decap_8 FILLER_72_727 ();
 sg13g2_decap_8 FILLER_72_734 ();
 sg13g2_decap_8 FILLER_72_741 ();
 sg13g2_decap_8 FILLER_72_748 ();
 sg13g2_decap_8 FILLER_72_755 ();
 sg13g2_decap_8 FILLER_72_762 ();
 sg13g2_decap_8 FILLER_72_769 ();
 sg13g2_decap_8 FILLER_72_776 ();
 sg13g2_decap_8 FILLER_72_783 ();
 sg13g2_decap_8 FILLER_72_790 ();
 sg13g2_decap_8 FILLER_72_797 ();
 sg13g2_decap_8 FILLER_72_804 ();
 sg13g2_decap_8 FILLER_72_811 ();
 sg13g2_decap_8 FILLER_72_818 ();
 sg13g2_decap_8 FILLER_72_825 ();
 sg13g2_decap_8 FILLER_72_832 ();
 sg13g2_decap_8 FILLER_72_839 ();
 sg13g2_decap_8 FILLER_72_846 ();
 sg13g2_decap_8 FILLER_72_853 ();
 sg13g2_decap_8 FILLER_72_860 ();
 sg13g2_decap_8 FILLER_72_867 ();
 sg13g2_decap_4 FILLER_72_874 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_8 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_decap_8 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_245 ();
 sg13g2_decap_8 FILLER_73_252 ();
 sg13g2_decap_8 FILLER_73_259 ();
 sg13g2_decap_8 FILLER_73_266 ();
 sg13g2_decap_8 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_decap_8 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_322 ();
 sg13g2_decap_8 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_73_336 ();
 sg13g2_decap_8 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_350 ();
 sg13g2_decap_8 FILLER_73_357 ();
 sg13g2_decap_8 FILLER_73_364 ();
 sg13g2_decap_8 FILLER_73_371 ();
 sg13g2_decap_8 FILLER_73_378 ();
 sg13g2_decap_8 FILLER_73_385 ();
 sg13g2_decap_8 FILLER_73_392 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_decap_8 FILLER_73_427 ();
 sg13g2_decap_8 FILLER_73_434 ();
 sg13g2_decap_8 FILLER_73_441 ();
 sg13g2_decap_8 FILLER_73_448 ();
 sg13g2_decap_8 FILLER_73_455 ();
 sg13g2_decap_8 FILLER_73_462 ();
 sg13g2_decap_8 FILLER_73_469 ();
 sg13g2_decap_8 FILLER_73_476 ();
 sg13g2_decap_8 FILLER_73_483 ();
 sg13g2_decap_8 FILLER_73_490 ();
 sg13g2_decap_8 FILLER_73_497 ();
 sg13g2_decap_8 FILLER_73_504 ();
 sg13g2_decap_8 FILLER_73_511 ();
 sg13g2_decap_8 FILLER_73_518 ();
 sg13g2_decap_8 FILLER_73_525 ();
 sg13g2_decap_8 FILLER_73_532 ();
 sg13g2_decap_8 FILLER_73_539 ();
 sg13g2_decap_8 FILLER_73_546 ();
 sg13g2_decap_8 FILLER_73_553 ();
 sg13g2_decap_8 FILLER_73_560 ();
 sg13g2_decap_8 FILLER_73_567 ();
 sg13g2_decap_8 FILLER_73_574 ();
 sg13g2_decap_8 FILLER_73_581 ();
 sg13g2_decap_8 FILLER_73_588 ();
 sg13g2_decap_8 FILLER_73_595 ();
 sg13g2_decap_8 FILLER_73_602 ();
 sg13g2_decap_8 FILLER_73_609 ();
 sg13g2_decap_8 FILLER_73_616 ();
 sg13g2_decap_8 FILLER_73_623 ();
 sg13g2_decap_8 FILLER_73_630 ();
 sg13g2_decap_8 FILLER_73_637 ();
 sg13g2_decap_8 FILLER_73_644 ();
 sg13g2_decap_8 FILLER_73_651 ();
 sg13g2_decap_8 FILLER_73_658 ();
 sg13g2_decap_8 FILLER_73_665 ();
 sg13g2_decap_8 FILLER_73_672 ();
 sg13g2_decap_8 FILLER_73_679 ();
 sg13g2_decap_8 FILLER_73_686 ();
 sg13g2_decap_8 FILLER_73_693 ();
 sg13g2_decap_8 FILLER_73_700 ();
 sg13g2_decap_8 FILLER_73_707 ();
 sg13g2_decap_8 FILLER_73_714 ();
 sg13g2_decap_8 FILLER_73_721 ();
 sg13g2_decap_8 FILLER_73_728 ();
 sg13g2_decap_8 FILLER_73_735 ();
 sg13g2_decap_8 FILLER_73_742 ();
 sg13g2_decap_8 FILLER_73_749 ();
 sg13g2_decap_8 FILLER_73_756 ();
 sg13g2_decap_8 FILLER_73_763 ();
 sg13g2_decap_8 FILLER_73_770 ();
 sg13g2_decap_8 FILLER_73_777 ();
 sg13g2_decap_8 FILLER_73_784 ();
 sg13g2_decap_8 FILLER_73_791 ();
 sg13g2_decap_8 FILLER_73_798 ();
 sg13g2_decap_8 FILLER_73_805 ();
 sg13g2_decap_8 FILLER_73_812 ();
 sg13g2_decap_8 FILLER_73_819 ();
 sg13g2_decap_8 FILLER_73_826 ();
 sg13g2_decap_8 FILLER_73_833 ();
 sg13g2_decap_8 FILLER_73_840 ();
 sg13g2_decap_8 FILLER_73_847 ();
 sg13g2_decap_8 FILLER_73_854 ();
 sg13g2_decap_8 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_73_868 ();
 sg13g2_fill_2 FILLER_73_875 ();
 sg13g2_fill_1 FILLER_73_877 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_20 ();
 sg13g2_decap_8 FILLER_74_27 ();
 sg13g2_decap_8 FILLER_74_34 ();
 sg13g2_decap_8 FILLER_74_41 ();
 sg13g2_decap_8 FILLER_74_48 ();
 sg13g2_decap_8 FILLER_74_55 ();
 sg13g2_decap_8 FILLER_74_62 ();
 sg13g2_decap_8 FILLER_74_69 ();
 sg13g2_decap_8 FILLER_74_76 ();
 sg13g2_decap_8 FILLER_74_83 ();
 sg13g2_decap_8 FILLER_74_90 ();
 sg13g2_decap_8 FILLER_74_97 ();
 sg13g2_decap_8 FILLER_74_104 ();
 sg13g2_decap_8 FILLER_74_111 ();
 sg13g2_decap_8 FILLER_74_118 ();
 sg13g2_decap_8 FILLER_74_125 ();
 sg13g2_decap_8 FILLER_74_132 ();
 sg13g2_decap_8 FILLER_74_139 ();
 sg13g2_decap_8 FILLER_74_146 ();
 sg13g2_decap_8 FILLER_74_153 ();
 sg13g2_decap_8 FILLER_74_160 ();
 sg13g2_decap_8 FILLER_74_167 ();
 sg13g2_decap_8 FILLER_74_174 ();
 sg13g2_decap_8 FILLER_74_181 ();
 sg13g2_decap_8 FILLER_74_188 ();
 sg13g2_decap_8 FILLER_74_195 ();
 sg13g2_decap_8 FILLER_74_202 ();
 sg13g2_decap_8 FILLER_74_209 ();
 sg13g2_decap_8 FILLER_74_216 ();
 sg13g2_decap_8 FILLER_74_223 ();
 sg13g2_decap_8 FILLER_74_230 ();
 sg13g2_decap_8 FILLER_74_237 ();
 sg13g2_decap_8 FILLER_74_244 ();
 sg13g2_decap_8 FILLER_74_251 ();
 sg13g2_decap_8 FILLER_74_258 ();
 sg13g2_decap_8 FILLER_74_265 ();
 sg13g2_decap_8 FILLER_74_272 ();
 sg13g2_decap_8 FILLER_74_279 ();
 sg13g2_decap_8 FILLER_74_286 ();
 sg13g2_decap_8 FILLER_74_293 ();
 sg13g2_decap_8 FILLER_74_300 ();
 sg13g2_decap_8 FILLER_74_307 ();
 sg13g2_decap_8 FILLER_74_314 ();
 sg13g2_decap_8 FILLER_74_321 ();
 sg13g2_decap_8 FILLER_74_328 ();
 sg13g2_decap_8 FILLER_74_335 ();
 sg13g2_decap_8 FILLER_74_342 ();
 sg13g2_decap_8 FILLER_74_349 ();
 sg13g2_decap_8 FILLER_74_356 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_decap_8 FILLER_74_370 ();
 sg13g2_decap_8 FILLER_74_377 ();
 sg13g2_decap_8 FILLER_74_384 ();
 sg13g2_decap_8 FILLER_74_391 ();
 sg13g2_decap_8 FILLER_74_398 ();
 sg13g2_decap_8 FILLER_74_405 ();
 sg13g2_decap_8 FILLER_74_412 ();
 sg13g2_decap_8 FILLER_74_419 ();
 sg13g2_decap_8 FILLER_74_426 ();
 sg13g2_decap_8 FILLER_74_433 ();
 sg13g2_decap_8 FILLER_74_440 ();
 sg13g2_decap_8 FILLER_74_447 ();
 sg13g2_decap_8 FILLER_74_454 ();
 sg13g2_decap_8 FILLER_74_461 ();
 sg13g2_decap_8 FILLER_74_468 ();
 sg13g2_decap_8 FILLER_74_475 ();
 sg13g2_decap_8 FILLER_74_482 ();
 sg13g2_decap_8 FILLER_74_489 ();
 sg13g2_decap_8 FILLER_74_496 ();
 sg13g2_decap_8 FILLER_74_503 ();
 sg13g2_decap_8 FILLER_74_510 ();
 sg13g2_decap_8 FILLER_74_517 ();
 sg13g2_decap_8 FILLER_74_524 ();
 sg13g2_decap_8 FILLER_74_531 ();
 sg13g2_decap_8 FILLER_74_538 ();
 sg13g2_decap_8 FILLER_74_545 ();
 sg13g2_decap_8 FILLER_74_552 ();
 sg13g2_decap_8 FILLER_74_559 ();
 sg13g2_decap_8 FILLER_74_566 ();
 sg13g2_decap_8 FILLER_74_573 ();
 sg13g2_decap_8 FILLER_74_580 ();
 sg13g2_decap_8 FILLER_74_587 ();
 sg13g2_decap_8 FILLER_74_594 ();
 sg13g2_decap_8 FILLER_74_601 ();
 sg13g2_decap_8 FILLER_74_608 ();
 sg13g2_decap_8 FILLER_74_615 ();
 sg13g2_decap_8 FILLER_74_622 ();
 sg13g2_decap_8 FILLER_74_629 ();
 sg13g2_decap_8 FILLER_74_636 ();
 sg13g2_decap_8 FILLER_74_643 ();
 sg13g2_decap_8 FILLER_74_650 ();
 sg13g2_decap_8 FILLER_74_657 ();
 sg13g2_decap_8 FILLER_74_664 ();
 sg13g2_decap_8 FILLER_74_671 ();
 sg13g2_decap_8 FILLER_74_678 ();
 sg13g2_decap_8 FILLER_74_685 ();
 sg13g2_decap_8 FILLER_74_692 ();
 sg13g2_decap_8 FILLER_74_699 ();
 sg13g2_decap_8 FILLER_74_706 ();
 sg13g2_decap_8 FILLER_74_713 ();
 sg13g2_decap_8 FILLER_74_720 ();
 sg13g2_decap_8 FILLER_74_727 ();
 sg13g2_decap_8 FILLER_74_734 ();
 sg13g2_decap_8 FILLER_74_741 ();
 sg13g2_decap_8 FILLER_74_748 ();
 sg13g2_decap_8 FILLER_74_755 ();
 sg13g2_decap_8 FILLER_74_762 ();
 sg13g2_decap_8 FILLER_74_769 ();
 sg13g2_decap_8 FILLER_74_776 ();
 sg13g2_decap_8 FILLER_74_783 ();
 sg13g2_decap_8 FILLER_74_790 ();
 sg13g2_decap_8 FILLER_74_797 ();
 sg13g2_decap_8 FILLER_74_804 ();
 sg13g2_decap_8 FILLER_74_811 ();
 sg13g2_decap_8 FILLER_74_818 ();
 sg13g2_decap_8 FILLER_74_825 ();
 sg13g2_decap_8 FILLER_74_832 ();
 sg13g2_decap_8 FILLER_74_839 ();
 sg13g2_decap_8 FILLER_74_846 ();
 sg13g2_decap_8 FILLER_74_853 ();
 sg13g2_decap_8 FILLER_74_860 ();
 sg13g2_decap_8 FILLER_74_867 ();
 sg13g2_decap_4 FILLER_74_874 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_12 ();
 sg13g2_decap_8 FILLER_75_19 ();
 sg13g2_decap_8 FILLER_75_26 ();
 sg13g2_decap_8 FILLER_75_33 ();
 sg13g2_decap_8 FILLER_75_40 ();
 sg13g2_decap_8 FILLER_75_47 ();
 sg13g2_decap_8 FILLER_75_54 ();
 sg13g2_decap_8 FILLER_75_61 ();
 sg13g2_decap_8 FILLER_75_68 ();
 sg13g2_decap_8 FILLER_75_75 ();
 sg13g2_decap_8 FILLER_75_82 ();
 sg13g2_decap_8 FILLER_75_89 ();
 sg13g2_decap_8 FILLER_75_96 ();
 sg13g2_decap_8 FILLER_75_103 ();
 sg13g2_decap_8 FILLER_75_110 ();
 sg13g2_decap_8 FILLER_75_117 ();
 sg13g2_decap_8 FILLER_75_124 ();
 sg13g2_decap_8 FILLER_75_131 ();
 sg13g2_decap_8 FILLER_75_138 ();
 sg13g2_decap_8 FILLER_75_145 ();
 sg13g2_decap_8 FILLER_75_152 ();
 sg13g2_decap_8 FILLER_75_159 ();
 sg13g2_decap_8 FILLER_75_166 ();
 sg13g2_decap_8 FILLER_75_173 ();
 sg13g2_decap_8 FILLER_75_180 ();
 sg13g2_decap_8 FILLER_75_187 ();
 sg13g2_decap_8 FILLER_75_194 ();
 sg13g2_decap_8 FILLER_75_201 ();
 sg13g2_decap_8 FILLER_75_208 ();
 sg13g2_decap_8 FILLER_75_215 ();
 sg13g2_decap_8 FILLER_75_222 ();
 sg13g2_decap_8 FILLER_75_229 ();
 sg13g2_decap_8 FILLER_75_236 ();
 sg13g2_decap_8 FILLER_75_243 ();
 sg13g2_decap_8 FILLER_75_250 ();
 sg13g2_decap_8 FILLER_75_257 ();
 sg13g2_decap_8 FILLER_75_264 ();
 sg13g2_decap_8 FILLER_75_271 ();
 sg13g2_decap_8 FILLER_75_278 ();
 sg13g2_decap_8 FILLER_75_285 ();
 sg13g2_decap_8 FILLER_75_292 ();
 sg13g2_decap_8 FILLER_75_299 ();
 sg13g2_decap_8 FILLER_75_306 ();
 sg13g2_decap_8 FILLER_75_313 ();
 sg13g2_decap_8 FILLER_75_320 ();
 sg13g2_decap_8 FILLER_75_327 ();
 sg13g2_decap_8 FILLER_75_334 ();
 sg13g2_decap_8 FILLER_75_341 ();
 sg13g2_decap_8 FILLER_75_348 ();
 sg13g2_decap_8 FILLER_75_355 ();
 sg13g2_decap_8 FILLER_75_362 ();
 sg13g2_decap_8 FILLER_75_369 ();
 sg13g2_decap_8 FILLER_75_376 ();
 sg13g2_decap_8 FILLER_75_383 ();
 sg13g2_decap_8 FILLER_75_390 ();
 sg13g2_decap_8 FILLER_75_397 ();
 sg13g2_decap_8 FILLER_75_404 ();
 sg13g2_decap_8 FILLER_75_411 ();
 sg13g2_decap_8 FILLER_75_418 ();
 sg13g2_decap_8 FILLER_75_425 ();
 sg13g2_decap_8 FILLER_75_432 ();
 sg13g2_decap_8 FILLER_75_439 ();
 sg13g2_decap_8 FILLER_75_446 ();
 sg13g2_decap_8 FILLER_75_453 ();
 sg13g2_decap_8 FILLER_75_460 ();
 sg13g2_decap_8 FILLER_75_467 ();
 sg13g2_decap_8 FILLER_75_474 ();
 sg13g2_decap_8 FILLER_75_481 ();
 sg13g2_decap_8 FILLER_75_488 ();
 sg13g2_decap_8 FILLER_75_495 ();
 sg13g2_decap_8 FILLER_75_502 ();
 sg13g2_decap_8 FILLER_75_509 ();
 sg13g2_decap_8 FILLER_75_516 ();
 sg13g2_decap_8 FILLER_75_523 ();
 sg13g2_decap_8 FILLER_75_530 ();
 sg13g2_decap_8 FILLER_75_537 ();
 sg13g2_decap_8 FILLER_75_544 ();
 sg13g2_decap_8 FILLER_75_551 ();
 sg13g2_decap_8 FILLER_75_558 ();
 sg13g2_decap_8 FILLER_75_565 ();
 sg13g2_decap_8 FILLER_75_572 ();
 sg13g2_decap_8 FILLER_75_579 ();
 sg13g2_decap_8 FILLER_75_586 ();
 sg13g2_decap_8 FILLER_75_593 ();
 sg13g2_decap_8 FILLER_75_600 ();
 sg13g2_decap_8 FILLER_75_607 ();
 sg13g2_decap_8 FILLER_75_614 ();
 sg13g2_decap_8 FILLER_75_621 ();
 sg13g2_decap_8 FILLER_75_628 ();
 sg13g2_decap_8 FILLER_75_635 ();
 sg13g2_decap_8 FILLER_75_642 ();
 sg13g2_decap_8 FILLER_75_649 ();
 sg13g2_decap_8 FILLER_75_656 ();
 sg13g2_decap_8 FILLER_75_663 ();
 sg13g2_decap_8 FILLER_75_670 ();
 sg13g2_decap_8 FILLER_75_677 ();
 sg13g2_decap_8 FILLER_75_684 ();
 sg13g2_decap_8 FILLER_75_691 ();
 sg13g2_decap_8 FILLER_75_698 ();
 sg13g2_decap_8 FILLER_75_705 ();
 sg13g2_decap_8 FILLER_75_712 ();
 sg13g2_decap_8 FILLER_75_719 ();
 sg13g2_decap_8 FILLER_75_726 ();
 sg13g2_decap_8 FILLER_75_733 ();
 sg13g2_decap_8 FILLER_75_740 ();
 sg13g2_decap_8 FILLER_75_747 ();
 sg13g2_decap_8 FILLER_75_754 ();
 sg13g2_decap_8 FILLER_75_761 ();
 sg13g2_decap_8 FILLER_75_768 ();
 sg13g2_decap_8 FILLER_75_775 ();
 sg13g2_decap_8 FILLER_75_782 ();
 sg13g2_decap_8 FILLER_75_789 ();
 sg13g2_decap_8 FILLER_75_796 ();
 sg13g2_decap_8 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_810 ();
 sg13g2_decap_8 FILLER_75_817 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_decap_8 FILLER_75_859 ();
 sg13g2_decap_8 FILLER_75_866 ();
 sg13g2_decap_4 FILLER_75_873 ();
 sg13g2_fill_1 FILLER_75_877 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_413 ();
 sg13g2_decap_8 FILLER_76_420 ();
 sg13g2_decap_8 FILLER_76_427 ();
 sg13g2_decap_8 FILLER_76_434 ();
 sg13g2_decap_8 FILLER_76_441 ();
 sg13g2_decap_8 FILLER_76_448 ();
 sg13g2_decap_8 FILLER_76_455 ();
 sg13g2_decap_8 FILLER_76_462 ();
 sg13g2_decap_8 FILLER_76_469 ();
 sg13g2_decap_8 FILLER_76_476 ();
 sg13g2_decap_8 FILLER_76_483 ();
 sg13g2_decap_8 FILLER_76_490 ();
 sg13g2_decap_8 FILLER_76_497 ();
 sg13g2_decap_8 FILLER_76_504 ();
 sg13g2_decap_8 FILLER_76_511 ();
 sg13g2_decap_8 FILLER_76_518 ();
 sg13g2_decap_8 FILLER_76_525 ();
 sg13g2_decap_8 FILLER_76_532 ();
 sg13g2_decap_8 FILLER_76_539 ();
 sg13g2_decap_8 FILLER_76_546 ();
 sg13g2_decap_8 FILLER_76_553 ();
 sg13g2_decap_8 FILLER_76_560 ();
 sg13g2_decap_8 FILLER_76_567 ();
 sg13g2_decap_8 FILLER_76_574 ();
 sg13g2_decap_8 FILLER_76_581 ();
 sg13g2_decap_8 FILLER_76_588 ();
 sg13g2_decap_8 FILLER_76_595 ();
 sg13g2_decap_8 FILLER_76_602 ();
 sg13g2_decap_8 FILLER_76_609 ();
 sg13g2_decap_8 FILLER_76_616 ();
 sg13g2_decap_8 FILLER_76_623 ();
 sg13g2_decap_8 FILLER_76_630 ();
 sg13g2_decap_8 FILLER_76_637 ();
 sg13g2_decap_8 FILLER_76_644 ();
 sg13g2_decap_8 FILLER_76_651 ();
 sg13g2_decap_8 FILLER_76_658 ();
 sg13g2_decap_8 FILLER_76_665 ();
 sg13g2_decap_8 FILLER_76_672 ();
 sg13g2_decap_8 FILLER_76_679 ();
 sg13g2_decap_8 FILLER_76_686 ();
 sg13g2_decap_8 FILLER_76_693 ();
 sg13g2_decap_8 FILLER_76_700 ();
 sg13g2_decap_8 FILLER_76_707 ();
 sg13g2_decap_8 FILLER_76_714 ();
 sg13g2_decap_8 FILLER_76_721 ();
 sg13g2_decap_8 FILLER_76_728 ();
 sg13g2_decap_8 FILLER_76_735 ();
 sg13g2_decap_8 FILLER_76_742 ();
 sg13g2_decap_8 FILLER_76_749 ();
 sg13g2_decap_8 FILLER_76_756 ();
 sg13g2_decap_8 FILLER_76_763 ();
 sg13g2_decap_8 FILLER_76_770 ();
 sg13g2_decap_8 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_784 ();
 sg13g2_decap_8 FILLER_76_791 ();
 sg13g2_decap_8 FILLER_76_798 ();
 sg13g2_decap_8 FILLER_76_805 ();
 sg13g2_decap_8 FILLER_76_812 ();
 sg13g2_decap_8 FILLER_76_819 ();
 sg13g2_decap_8 FILLER_76_826 ();
 sg13g2_decap_8 FILLER_76_833 ();
 sg13g2_decap_8 FILLER_76_840 ();
 sg13g2_decap_8 FILLER_76_847 ();
 sg13g2_decap_8 FILLER_76_854 ();
 sg13g2_decap_8 FILLER_76_861 ();
 sg13g2_decap_8 FILLER_76_868 ();
 sg13g2_fill_2 FILLER_76_875 ();
 sg13g2_fill_1 FILLER_76_877 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_4 FILLER_77_224 ();
 sg13g2_fill_1 FILLER_77_228 ();
 sg13g2_decap_4 FILLER_77_232 ();
 sg13g2_fill_1 FILLER_77_236 ();
 sg13g2_fill_2 FILLER_77_243 ();
 sg13g2_fill_2 FILLER_77_251 ();
 sg13g2_decap_8 FILLER_77_256 ();
 sg13g2_decap_8 FILLER_77_263 ();
 sg13g2_decap_8 FILLER_77_270 ();
 sg13g2_decap_8 FILLER_77_277 ();
 sg13g2_decap_8 FILLER_77_284 ();
 sg13g2_decap_8 FILLER_77_291 ();
 sg13g2_decap_8 FILLER_77_298 ();
 sg13g2_decap_8 FILLER_77_305 ();
 sg13g2_decap_8 FILLER_77_312 ();
 sg13g2_decap_8 FILLER_77_319 ();
 sg13g2_decap_8 FILLER_77_326 ();
 sg13g2_decap_8 FILLER_77_333 ();
 sg13g2_decap_8 FILLER_77_340 ();
 sg13g2_decap_8 FILLER_77_347 ();
 sg13g2_decap_8 FILLER_77_354 ();
 sg13g2_decap_8 FILLER_77_361 ();
 sg13g2_decap_8 FILLER_77_368 ();
 sg13g2_decap_8 FILLER_77_375 ();
 sg13g2_decap_8 FILLER_77_382 ();
 sg13g2_decap_8 FILLER_77_389 ();
 sg13g2_decap_8 FILLER_77_396 ();
 sg13g2_decap_8 FILLER_77_403 ();
 sg13g2_decap_8 FILLER_77_410 ();
 sg13g2_decap_8 FILLER_77_417 ();
 sg13g2_decap_8 FILLER_77_424 ();
 sg13g2_decap_8 FILLER_77_431 ();
 sg13g2_decap_8 FILLER_77_438 ();
 sg13g2_decap_8 FILLER_77_445 ();
 sg13g2_decap_8 FILLER_77_452 ();
 sg13g2_decap_8 FILLER_77_459 ();
 sg13g2_decap_8 FILLER_77_466 ();
 sg13g2_decap_8 FILLER_77_473 ();
 sg13g2_decap_8 FILLER_77_480 ();
 sg13g2_decap_8 FILLER_77_487 ();
 sg13g2_decap_8 FILLER_77_494 ();
 sg13g2_decap_8 FILLER_77_501 ();
 sg13g2_decap_8 FILLER_77_508 ();
 sg13g2_decap_8 FILLER_77_515 ();
 sg13g2_decap_8 FILLER_77_522 ();
 sg13g2_decap_8 FILLER_77_529 ();
 sg13g2_decap_8 FILLER_77_536 ();
 sg13g2_decap_8 FILLER_77_543 ();
 sg13g2_decap_8 FILLER_77_550 ();
 sg13g2_decap_8 FILLER_77_557 ();
 sg13g2_decap_8 FILLER_77_564 ();
 sg13g2_decap_8 FILLER_77_571 ();
 sg13g2_decap_8 FILLER_77_578 ();
 sg13g2_decap_8 FILLER_77_585 ();
 sg13g2_decap_8 FILLER_77_592 ();
 sg13g2_decap_8 FILLER_77_599 ();
 sg13g2_decap_8 FILLER_77_606 ();
 sg13g2_decap_8 FILLER_77_613 ();
 sg13g2_decap_8 FILLER_77_620 ();
 sg13g2_decap_8 FILLER_77_627 ();
 sg13g2_decap_8 FILLER_77_634 ();
 sg13g2_decap_8 FILLER_77_641 ();
 sg13g2_decap_8 FILLER_77_648 ();
 sg13g2_decap_8 FILLER_77_655 ();
 sg13g2_decap_8 FILLER_77_662 ();
 sg13g2_decap_8 FILLER_77_669 ();
 sg13g2_decap_8 FILLER_77_676 ();
 sg13g2_decap_8 FILLER_77_683 ();
 sg13g2_decap_8 FILLER_77_690 ();
 sg13g2_decap_8 FILLER_77_697 ();
 sg13g2_decap_8 FILLER_77_704 ();
 sg13g2_decap_8 FILLER_77_711 ();
 sg13g2_decap_8 FILLER_77_718 ();
 sg13g2_decap_8 FILLER_77_725 ();
 sg13g2_decap_8 FILLER_77_732 ();
 sg13g2_decap_8 FILLER_77_739 ();
 sg13g2_decap_8 FILLER_77_746 ();
 sg13g2_decap_8 FILLER_77_753 ();
 sg13g2_decap_8 FILLER_77_760 ();
 sg13g2_decap_8 FILLER_77_767 ();
 sg13g2_decap_8 FILLER_77_774 ();
 sg13g2_decap_8 FILLER_77_781 ();
 sg13g2_decap_8 FILLER_77_788 ();
 sg13g2_decap_8 FILLER_77_795 ();
 sg13g2_decap_8 FILLER_77_802 ();
 sg13g2_decap_8 FILLER_77_809 ();
 sg13g2_decap_8 FILLER_77_816 ();
 sg13g2_decap_8 FILLER_77_823 ();
 sg13g2_decap_8 FILLER_77_830 ();
 sg13g2_decap_8 FILLER_77_837 ();
 sg13g2_decap_8 FILLER_77_844 ();
 sg13g2_decap_8 FILLER_77_851 ();
 sg13g2_decap_8 FILLER_77_858 ();
 sg13g2_decap_8 FILLER_77_865 ();
 sg13g2_decap_4 FILLER_77_872 ();
 sg13g2_fill_2 FILLER_77_876 ();
 sg13g2_decap_4 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_20 ();
 sg13g2_decap_8 FILLER_78_27 ();
 sg13g2_decap_8 FILLER_78_34 ();
 sg13g2_decap_8 FILLER_78_41 ();
 sg13g2_decap_8 FILLER_78_48 ();
 sg13g2_decap_8 FILLER_78_55 ();
 sg13g2_decap_8 FILLER_78_62 ();
 sg13g2_decap_8 FILLER_78_69 ();
 sg13g2_decap_8 FILLER_78_76 ();
 sg13g2_decap_8 FILLER_78_83 ();
 sg13g2_decap_8 FILLER_78_90 ();
 sg13g2_decap_8 FILLER_78_97 ();
 sg13g2_decap_8 FILLER_78_104 ();
 sg13g2_decap_8 FILLER_78_111 ();
 sg13g2_decap_8 FILLER_78_118 ();
 sg13g2_decap_8 FILLER_78_125 ();
 sg13g2_decap_8 FILLER_78_132 ();
 sg13g2_decap_8 FILLER_78_139 ();
 sg13g2_decap_8 FILLER_78_146 ();
 sg13g2_decap_8 FILLER_78_153 ();
 sg13g2_decap_8 FILLER_78_160 ();
 sg13g2_decap_8 FILLER_78_167 ();
 sg13g2_decap_8 FILLER_78_174 ();
 sg13g2_decap_8 FILLER_78_181 ();
 sg13g2_decap_8 FILLER_78_188 ();
 sg13g2_decap_8 FILLER_78_195 ();
 sg13g2_decap_4 FILLER_78_202 ();
 sg13g2_fill_1 FILLER_78_206 ();
 sg13g2_fill_2 FILLER_78_243 ();
 sg13g2_fill_2 FILLER_78_251 ();
 sg13g2_fill_2 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_270 ();
 sg13g2_decap_8 FILLER_78_277 ();
 sg13g2_decap_8 FILLER_78_284 ();
 sg13g2_decap_8 FILLER_78_291 ();
 sg13g2_decap_8 FILLER_78_298 ();
 sg13g2_decap_8 FILLER_78_305 ();
 sg13g2_decap_8 FILLER_78_312 ();
 sg13g2_decap_8 FILLER_78_319 ();
 sg13g2_decap_8 FILLER_78_326 ();
 sg13g2_decap_8 FILLER_78_333 ();
 sg13g2_decap_8 FILLER_78_340 ();
 sg13g2_decap_8 FILLER_78_347 ();
 sg13g2_decap_8 FILLER_78_354 ();
 sg13g2_decap_8 FILLER_78_361 ();
 sg13g2_decap_8 FILLER_78_368 ();
 sg13g2_decap_8 FILLER_78_375 ();
 sg13g2_decap_8 FILLER_78_382 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_8 FILLER_78_403 ();
 sg13g2_decap_8 FILLER_78_410 ();
 sg13g2_decap_8 FILLER_78_417 ();
 sg13g2_decap_8 FILLER_78_424 ();
 sg13g2_decap_8 FILLER_78_431 ();
 sg13g2_decap_8 FILLER_78_438 ();
 sg13g2_decap_8 FILLER_78_445 ();
 sg13g2_decap_8 FILLER_78_452 ();
 sg13g2_decap_8 FILLER_78_459 ();
 sg13g2_decap_8 FILLER_78_466 ();
 sg13g2_decap_8 FILLER_78_473 ();
 sg13g2_decap_8 FILLER_78_480 ();
 sg13g2_decap_8 FILLER_78_487 ();
 sg13g2_decap_8 FILLER_78_494 ();
 sg13g2_decap_8 FILLER_78_501 ();
 sg13g2_decap_8 FILLER_78_508 ();
 sg13g2_decap_8 FILLER_78_515 ();
 sg13g2_decap_8 FILLER_78_522 ();
 sg13g2_decap_8 FILLER_78_529 ();
 sg13g2_decap_8 FILLER_78_536 ();
 sg13g2_decap_8 FILLER_78_543 ();
 sg13g2_decap_8 FILLER_78_550 ();
 sg13g2_decap_8 FILLER_78_557 ();
 sg13g2_decap_8 FILLER_78_564 ();
 sg13g2_decap_8 FILLER_78_571 ();
 sg13g2_decap_8 FILLER_78_578 ();
 sg13g2_decap_8 FILLER_78_585 ();
 sg13g2_decap_8 FILLER_78_592 ();
 sg13g2_decap_8 FILLER_78_599 ();
 sg13g2_decap_8 FILLER_78_606 ();
 sg13g2_decap_8 FILLER_78_613 ();
 sg13g2_decap_8 FILLER_78_620 ();
 sg13g2_decap_8 FILLER_78_627 ();
 sg13g2_decap_8 FILLER_78_634 ();
 sg13g2_decap_8 FILLER_78_641 ();
 sg13g2_decap_8 FILLER_78_648 ();
 sg13g2_decap_8 FILLER_78_655 ();
 sg13g2_decap_8 FILLER_78_662 ();
 sg13g2_decap_8 FILLER_78_669 ();
 sg13g2_decap_8 FILLER_78_676 ();
 sg13g2_decap_8 FILLER_78_683 ();
 sg13g2_decap_8 FILLER_78_690 ();
 sg13g2_decap_8 FILLER_78_697 ();
 sg13g2_decap_8 FILLER_78_704 ();
 sg13g2_decap_8 FILLER_78_711 ();
 sg13g2_decap_8 FILLER_78_718 ();
 sg13g2_decap_8 FILLER_78_725 ();
 sg13g2_decap_8 FILLER_78_732 ();
 sg13g2_decap_8 FILLER_78_739 ();
 sg13g2_decap_8 FILLER_78_746 ();
 sg13g2_decap_8 FILLER_78_753 ();
 sg13g2_decap_8 FILLER_78_760 ();
 sg13g2_decap_8 FILLER_78_767 ();
 sg13g2_decap_8 FILLER_78_774 ();
 sg13g2_decap_8 FILLER_78_781 ();
 sg13g2_decap_8 FILLER_78_788 ();
 sg13g2_decap_8 FILLER_78_795 ();
 sg13g2_decap_8 FILLER_78_802 ();
 sg13g2_decap_8 FILLER_78_809 ();
 sg13g2_decap_8 FILLER_78_816 ();
 sg13g2_decap_8 FILLER_78_823 ();
 sg13g2_decap_8 FILLER_78_830 ();
 sg13g2_decap_8 FILLER_78_837 ();
 sg13g2_decap_8 FILLER_78_844 ();
 sg13g2_decap_8 FILLER_78_851 ();
 sg13g2_decap_8 FILLER_78_858 ();
 sg13g2_decap_8 FILLER_78_865 ();
 sg13g2_decap_4 FILLER_78_872 ();
 sg13g2_fill_2 FILLER_78_876 ();
 sg13g2_fill_1 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_4 FILLER_79_189 ();
 sg13g2_fill_2 FILLER_79_193 ();
 sg13g2_fill_1 FILLER_79_219 ();
 sg13g2_fill_2 FILLER_79_235 ();
 sg13g2_fill_2 FILLER_79_243 ();
 sg13g2_fill_2 FILLER_79_251 ();
 sg13g2_fill_2 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_276 ();
 sg13g2_decap_8 FILLER_79_283 ();
 sg13g2_decap_8 FILLER_79_290 ();
 sg13g2_decap_8 FILLER_79_297 ();
 sg13g2_decap_8 FILLER_79_304 ();
 sg13g2_decap_8 FILLER_79_311 ();
 sg13g2_decap_8 FILLER_79_318 ();
 sg13g2_decap_8 FILLER_79_325 ();
 sg13g2_decap_8 FILLER_79_332 ();
 sg13g2_decap_8 FILLER_79_339 ();
 sg13g2_decap_8 FILLER_79_346 ();
 sg13g2_decap_8 FILLER_79_353 ();
 sg13g2_decap_8 FILLER_79_360 ();
 sg13g2_decap_8 FILLER_79_367 ();
 sg13g2_decap_8 FILLER_79_374 ();
 sg13g2_decap_8 FILLER_79_381 ();
 sg13g2_decap_8 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_79_409 ();
 sg13g2_decap_8 FILLER_79_416 ();
 sg13g2_decap_8 FILLER_79_423 ();
 sg13g2_decap_8 FILLER_79_430 ();
 sg13g2_decap_8 FILLER_79_437 ();
 sg13g2_decap_8 FILLER_79_444 ();
 sg13g2_decap_8 FILLER_79_451 ();
 sg13g2_decap_8 FILLER_79_458 ();
 sg13g2_decap_8 FILLER_79_465 ();
 sg13g2_decap_8 FILLER_79_472 ();
 sg13g2_decap_8 FILLER_79_479 ();
 sg13g2_decap_8 FILLER_79_486 ();
 sg13g2_decap_8 FILLER_79_493 ();
 sg13g2_decap_8 FILLER_79_500 ();
 sg13g2_decap_8 FILLER_79_507 ();
 sg13g2_decap_8 FILLER_79_514 ();
 sg13g2_decap_8 FILLER_79_521 ();
 sg13g2_decap_8 FILLER_79_528 ();
 sg13g2_decap_8 FILLER_79_535 ();
 sg13g2_decap_8 FILLER_79_542 ();
 sg13g2_decap_8 FILLER_79_549 ();
 sg13g2_decap_8 FILLER_79_556 ();
 sg13g2_decap_8 FILLER_79_563 ();
 sg13g2_decap_8 FILLER_79_570 ();
 sg13g2_decap_8 FILLER_79_577 ();
 sg13g2_decap_8 FILLER_79_584 ();
 sg13g2_decap_8 FILLER_79_591 ();
 sg13g2_decap_8 FILLER_79_598 ();
 sg13g2_decap_8 FILLER_79_605 ();
 sg13g2_decap_8 FILLER_79_612 ();
 sg13g2_decap_8 FILLER_79_619 ();
 sg13g2_decap_8 FILLER_79_626 ();
 sg13g2_decap_8 FILLER_79_633 ();
 sg13g2_decap_8 FILLER_79_640 ();
 sg13g2_decap_8 FILLER_79_647 ();
 sg13g2_decap_8 FILLER_79_654 ();
 sg13g2_decap_8 FILLER_79_661 ();
 sg13g2_decap_8 FILLER_79_668 ();
 sg13g2_decap_8 FILLER_79_675 ();
 sg13g2_decap_8 FILLER_79_682 ();
 sg13g2_decap_8 FILLER_79_689 ();
 sg13g2_decap_8 FILLER_79_696 ();
 sg13g2_decap_8 FILLER_79_703 ();
 sg13g2_decap_8 FILLER_79_710 ();
 sg13g2_decap_8 FILLER_79_717 ();
 sg13g2_decap_8 FILLER_79_724 ();
 sg13g2_decap_8 FILLER_79_731 ();
 sg13g2_decap_8 FILLER_79_738 ();
 sg13g2_decap_8 FILLER_79_745 ();
 sg13g2_decap_8 FILLER_79_752 ();
 sg13g2_decap_8 FILLER_79_759 ();
 sg13g2_decap_8 FILLER_79_766 ();
 sg13g2_decap_8 FILLER_79_773 ();
 sg13g2_decap_8 FILLER_79_780 ();
 sg13g2_decap_8 FILLER_79_787 ();
 sg13g2_decap_8 FILLER_79_794 ();
 sg13g2_decap_8 FILLER_79_801 ();
 sg13g2_decap_8 FILLER_79_808 ();
 sg13g2_decap_8 FILLER_79_815 ();
 sg13g2_decap_8 FILLER_79_822 ();
 sg13g2_decap_8 FILLER_79_829 ();
 sg13g2_decap_8 FILLER_79_836 ();
 sg13g2_decap_8 FILLER_79_843 ();
 sg13g2_decap_8 FILLER_79_850 ();
 sg13g2_decap_8 FILLER_79_857 ();
 sg13g2_decap_8 FILLER_79_864 ();
 sg13g2_decap_8 FILLER_79_871 ();
 sg13g2_decap_8 FILLER_80_32 ();
 sg13g2_decap_8 FILLER_80_39 ();
 sg13g2_decap_8 FILLER_80_46 ();
 sg13g2_decap_8 FILLER_80_53 ();
 sg13g2_decap_8 FILLER_80_60 ();
 sg13g2_decap_8 FILLER_80_67 ();
 sg13g2_decap_8 FILLER_80_74 ();
 sg13g2_decap_8 FILLER_80_81 ();
 sg13g2_decap_8 FILLER_80_88 ();
 sg13g2_decap_8 FILLER_80_95 ();
 sg13g2_decap_8 FILLER_80_102 ();
 sg13g2_decap_8 FILLER_80_109 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_8 FILLER_80_123 ();
 sg13g2_decap_8 FILLER_80_130 ();
 sg13g2_decap_8 FILLER_80_137 ();
 sg13g2_decap_8 FILLER_80_144 ();
 sg13g2_decap_8 FILLER_80_151 ();
 sg13g2_decap_8 FILLER_80_158 ();
 sg13g2_decap_8 FILLER_80_165 ();
 sg13g2_decap_8 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_179 ();
 sg13g2_fill_1 FILLER_80_183 ();
 sg13g2_fill_1 FILLER_80_212 ();
 sg13g2_fill_1 FILLER_80_220 ();
 sg13g2_fill_1 FILLER_80_228 ();
 sg13g2_fill_1 FILLER_80_236 ();
 sg13g2_fill_1 FILLER_80_244 ();
 sg13g2_fill_1 FILLER_80_252 ();
 sg13g2_fill_1 FILLER_80_260 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_fill_1 FILLER_80_279 ();
 sg13g2_decap_4 FILLER_80_284 ();
 sg13g2_decap_4 FILLER_80_292 ();
 sg13g2_decap_4 FILLER_80_300 ();
 sg13g2_decap_4 FILLER_80_308 ();
 sg13g2_decap_4 FILLER_80_316 ();
 sg13g2_decap_4 FILLER_80_324 ();
 sg13g2_decap_4 FILLER_80_332 ();
 sg13g2_decap_4 FILLER_80_340 ();
 sg13g2_fill_2 FILLER_80_349 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_decap_4 FILLER_80_372 ();
 sg13g2_decap_4 FILLER_80_380 ();
 sg13g2_decap_4 FILLER_80_388 ();
 sg13g2_decap_4 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_412 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_8 FILLER_80_426 ();
 sg13g2_decap_8 FILLER_80_433 ();
 sg13g2_decap_8 FILLER_80_440 ();
 sg13g2_decap_8 FILLER_80_447 ();
 sg13g2_decap_8 FILLER_80_454 ();
 sg13g2_decap_8 FILLER_80_461 ();
 sg13g2_decap_8 FILLER_80_468 ();
 sg13g2_decap_8 FILLER_80_475 ();
 sg13g2_decap_8 FILLER_80_482 ();
 sg13g2_decap_8 FILLER_80_489 ();
 sg13g2_decap_8 FILLER_80_496 ();
 sg13g2_decap_8 FILLER_80_503 ();
 sg13g2_decap_8 FILLER_80_510 ();
 sg13g2_decap_8 FILLER_80_517 ();
 sg13g2_decap_8 FILLER_80_524 ();
 sg13g2_decap_8 FILLER_80_531 ();
 sg13g2_decap_8 FILLER_80_538 ();
 sg13g2_decap_8 FILLER_80_545 ();
 sg13g2_decap_8 FILLER_80_552 ();
 sg13g2_decap_8 FILLER_80_559 ();
 sg13g2_decap_8 FILLER_80_566 ();
 sg13g2_decap_8 FILLER_80_573 ();
 sg13g2_decap_8 FILLER_80_580 ();
 sg13g2_decap_8 FILLER_80_587 ();
 sg13g2_decap_8 FILLER_80_594 ();
 sg13g2_decap_8 FILLER_80_601 ();
 sg13g2_decap_8 FILLER_80_608 ();
 sg13g2_decap_8 FILLER_80_615 ();
 sg13g2_decap_8 FILLER_80_622 ();
 sg13g2_decap_8 FILLER_80_629 ();
 sg13g2_decap_8 FILLER_80_636 ();
 sg13g2_decap_8 FILLER_80_643 ();
 sg13g2_decap_8 FILLER_80_650 ();
 sg13g2_decap_8 FILLER_80_657 ();
 sg13g2_decap_8 FILLER_80_664 ();
 sg13g2_decap_8 FILLER_80_671 ();
 sg13g2_decap_8 FILLER_80_678 ();
 sg13g2_decap_8 FILLER_80_685 ();
 sg13g2_decap_8 FILLER_80_692 ();
 sg13g2_decap_8 FILLER_80_699 ();
 sg13g2_decap_8 FILLER_80_706 ();
 sg13g2_decap_8 FILLER_80_713 ();
 sg13g2_decap_8 FILLER_80_720 ();
 sg13g2_decap_8 FILLER_80_727 ();
 sg13g2_decap_8 FILLER_80_734 ();
 sg13g2_decap_8 FILLER_80_741 ();
 sg13g2_decap_8 FILLER_80_748 ();
 sg13g2_decap_8 FILLER_80_755 ();
 sg13g2_decap_8 FILLER_80_762 ();
 sg13g2_decap_8 FILLER_80_769 ();
 sg13g2_decap_8 FILLER_80_776 ();
 sg13g2_decap_8 FILLER_80_783 ();
 sg13g2_decap_8 FILLER_80_790 ();
 sg13g2_decap_8 FILLER_80_797 ();
 sg13g2_decap_8 FILLER_80_804 ();
 sg13g2_decap_8 FILLER_80_811 ();
 sg13g2_decap_8 FILLER_80_818 ();
 sg13g2_decap_8 FILLER_80_825 ();
 sg13g2_decap_8 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_846 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_decap_8 FILLER_80_860 ();
 sg13g2_decap_8 FILLER_80_867 ();
 sg13g2_decap_4 FILLER_80_874 ();
endmodule
