module tt_um_demosiine_sda (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire clknet_0_clk;
 wire net268;
 wire audio;
 wire \audio_engine_1.counter[0] ;
 wire \audio_engine_1.counter[10] ;
 wire \audio_engine_1.counter[11] ;
 wire \audio_engine_1.counter[12] ;
 wire \audio_engine_1.counter[13] ;
 wire \audio_engine_1.counter[14] ;
 wire \audio_engine_1.counter[15] ;
 wire \audio_engine_1.counter[16] ;
 wire \audio_engine_1.counter[17] ;
 wire \audio_engine_1.counter[1] ;
 wire \audio_engine_1.counter[2] ;
 wire \audio_engine_1.counter[3] ;
 wire \audio_engine_1.counter[4] ;
 wire \audio_engine_1.counter[5] ;
 wire \audio_engine_1.counter[6] ;
 wire \audio_engine_1.counter[7] ;
 wire \audio_engine_1.counter[8] ;
 wire \audio_engine_1.counter[9] ;
 wire \audio_engine_1.en_seq_clk ;
 wire \audio_engine_1.freq_synth1.audio_reg ;
 wire \audio_engine_1.freq_synth1.en_synth_clk ;
 wire \audio_engine_1.freq_synth1.hp_ctr[0] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[1] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[2] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[3] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[4] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[5] ;
 wire \audio_engine_1.freq_synth1.hp_ctr[6] ;
 wire \audio_engine_1.seq_ctr[0] ;
 wire \audio_engine_1.seq_ctr[1] ;
 wire \audio_engine_1.seq_ctr[2] ;
 wire \audio_engine_1.seq_ctr[3] ;
 wire \audio_engine_1.seq_ctr[4] ;
 wire \audio_engine_1.seq_time[0] ;
 wire \audio_engine_1.seq_time[1] ;
 wire \audio_engine_1.seq_time[2] ;
 wire \audio_engine_1.seq_time[3] ;
 wire \audio_engine_1.seq_time[4] ;
 wire \audio_engine_1.seq_time[5] ;
 wire \audio_engine_1.seq_time[6] ;
 wire \graphics_engine_1.anim_2x[0] ;
 wire \graphics_engine_1.ctr[0] ;
 wire \graphics_engine_1.ctr[1] ;
 wire \graphics_engine_1.ctr[2] ;
 wire \graphics_engine_1.ctr[3] ;
 wire \graphics_engine_1.ctr[4] ;
 wire \graphics_engine_1.ctr[5] ;
 wire \graphics_engine_1.ctr[6] ;
 wire \graphics_engine_1.ctr[7] ;
 wire \graphics_engine_1.ctr[8] ;
 wire \graphics_engine_1.en_v_sync ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_x[0] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[0] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[1] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[2] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[4] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[5] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[6] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[7] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[2] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[5] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[6] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ;
 wire \graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ;
 wire \graphics_engine_1.v_sync ;
 wire h_sync;
 wire \vga_controller_1.y[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _3089_ (.A(\vga_controller_1.y[9] ),
    .X(_1068_));
 sg13g2_buf_1 _3090_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ),
    .X(_1079_));
 sg13g2_buf_1 _3091_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ),
    .X(_1090_));
 sg13g2_buf_1 _3092_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[5] ),
    .X(_1101_));
 sg13g2_buf_1 _3093_ (.A(_1101_),
    .X(_1112_));
 sg13g2_buf_1 _3094_ (.A(_1112_),
    .X(_1123_));
 sg13g2_buf_2 _3095_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[6] ),
    .X(_1134_));
 sg13g2_buf_1 _3096_ (.A(_1134_),
    .X(_1145_));
 sg13g2_and2_1 _3097_ (.A(_1123_),
    .B(_1145_),
    .X(_1156_));
 sg13g2_buf_1 _3098_ (.A(_1156_),
    .X(_1167_));
 sg13g2_nand3_1 _3099_ (.B(net244),
    .C(_1167_),
    .A(net245),
    .Y(_1178_));
 sg13g2_buf_1 _3100_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[0] ),
    .X(_1189_));
 sg13g2_buf_1 _3101_ (.A(net243),
    .X(_1200_));
 sg13g2_buf_1 _3102_ (.A(net223),
    .X(_1211_));
 sg13g2_buf_1 _3103_ (.A(net193),
    .X(_1222_));
 sg13g2_buf_1 _3104_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[1] ),
    .X(_1233_));
 sg13g2_buf_1 _3105_ (.A(_1233_),
    .X(_1244_));
 sg13g2_buf_1 _3106_ (.A(net222),
    .X(_1255_));
 sg13g2_inv_2 _3107_ (.Y(_1266_),
    .A(net192));
 sg13g2_buf_1 _3108_ (.A(_1266_),
    .X(_1277_));
 sg13g2_nand2_2 _3109_ (.Y(_1288_),
    .A(_1222_),
    .B(net145));
 sg13g2_buf_1 _3110_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ),
    .X(_1299_));
 sg13g2_buf_1 _3111_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[2] ),
    .X(_1310_));
 sg13g2_buf_1 _3112_ (.A(_1310_),
    .X(_1321_));
 sg13g2_inv_2 _3113_ (.Y(_1332_),
    .A(net221));
 sg13g2_nand2_1 _3114_ (.Y(_1343_),
    .A(net242),
    .B(_1332_));
 sg13g2_nor4_1 _3115_ (.A(_1068_),
    .B(_1178_),
    .C(_1288_),
    .D(_1343_),
    .Y(_0005_));
 sg13g2_buf_1 _3116_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[6] ),
    .X(_1364_));
 sg13g2_buf_1 _3117_ (.A(net241),
    .X(_1375_));
 sg13g2_buf_2 _3118_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[5] ),
    .X(_1386_));
 sg13g2_buf_8 _3119_ (.A(_1386_),
    .X(_1397_));
 sg13g2_buf_1 _3120_ (.A(net219),
    .X(_1408_));
 sg13g2_buf_2 _3121_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[4] ),
    .X(_1419_));
 sg13g2_buf_8 _3122_ (.A(_1419_),
    .X(_1430_));
 sg13g2_buf_1 _3123_ (.A(_1430_),
    .X(_1441_));
 sg13g2_or2_1 _3124_ (.X(_1452_),
    .B(net190),
    .A(_1408_));
 sg13g2_buf_2 _3125_ (.A(_1452_),
    .X(_1463_));
 sg13g2_buf_1 _3126_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[7] ),
    .X(_1474_));
 sg13g2_o21ai_1 _3127_ (.B1(net240),
    .Y(_1485_),
    .A1(net220),
    .A2(_1463_));
 sg13g2_buf_2 _3128_ (.A(_1485_),
    .X(_1496_));
 sg13g2_buf_2 _3129_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ),
    .X(_1507_));
 sg13g2_inv_1 _3130_ (.Y(_1518_),
    .A(_1507_));
 sg13g2_nand2b_1 _3131_ (.Y(_1529_),
    .B(_1518_),
    .A_N(_1496_));
 sg13g2_buf_1 _3132_ (.A(net220),
    .X(_1540_));
 sg13g2_buf_1 _3133_ (.A(net189),
    .X(_1551_));
 sg13g2_buf_1 _3134_ (.A(net190),
    .X(_1562_));
 sg13g2_and2_1 _3135_ (.A(net191),
    .B(net167),
    .X(_1573_));
 sg13g2_buf_2 _3136_ (.A(_1573_),
    .X(_1584_));
 sg13g2_nand2_1 _3137_ (.Y(_1595_),
    .A(net168),
    .B(_1584_));
 sg13g2_nand2_1 _3138_ (.Y(_1606_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ),
    .B(_1595_));
 sg13g2_nor2_1 _3139_ (.A(_1529_),
    .B(_1606_),
    .Y(_0004_));
 sg13g2_buf_1 _3140_ (.A(\audio_engine_1.counter[10] ),
    .X(_1627_));
 sg13g2_buf_1 _3141_ (.A(\audio_engine_1.seq_time[3] ),
    .X(_1638_));
 sg13g2_buf_1 _3142_ (.A(_1638_),
    .X(_1649_));
 sg13g2_buf_1 _3143_ (.A(\audio_engine_1.seq_time[4] ),
    .X(_1660_));
 sg13g2_nand2_1 _3144_ (.Y(_1671_),
    .A(net217),
    .B(net239));
 sg13g2_buf_1 _3145_ (.A(\audio_engine_1.seq_time[1] ),
    .X(_1682_));
 sg13g2_buf_1 _3146_ (.A(_1682_),
    .X(_1693_));
 sg13g2_buf_2 _3147_ (.A(\audio_engine_1.seq_time[2] ),
    .X(_1704_));
 sg13g2_buf_1 _3148_ (.A(\audio_engine_1.seq_time[0] ),
    .X(_1715_));
 sg13g2_nor2b_1 _3149_ (.A(_1704_),
    .B_N(net237),
    .Y(_1726_));
 sg13g2_buf_2 _3150_ (.A(\audio_engine_1.seq_time[6] ),
    .X(_1737_));
 sg13g2_nand2b_1 _3151_ (.Y(_1748_),
    .B(_1704_),
    .A_N(net237));
 sg13g2_nor2_1 _3152_ (.A(_1737_),
    .B(_1748_),
    .Y(_1759_));
 sg13g2_or2_1 _3153_ (.X(_1770_),
    .B(_1759_),
    .A(_1726_));
 sg13g2_buf_1 _3154_ (.A(_1715_),
    .X(_1781_));
 sg13g2_buf_1 _3155_ (.A(_1704_),
    .X(_1792_));
 sg13g2_nor3_1 _3156_ (.A(net216),
    .B(net215),
    .C(net214),
    .Y(_1803_));
 sg13g2_a21oi_1 _3157_ (.A1(_1693_),
    .A2(_1770_),
    .Y(_1814_),
    .B1(_1803_));
 sg13g2_buf_1 _3158_ (.A(_1737_),
    .X(_1825_));
 sg13g2_inv_1 _3159_ (.Y(_1836_),
    .A(_1682_));
 sg13g2_nor2b_1 _3160_ (.A(_1649_),
    .B_N(net237),
    .Y(_1847_));
 sg13g2_inv_2 _3161_ (.Y(_1858_),
    .A(_1638_));
 sg13g2_nor2_2 _3162_ (.A(_1858_),
    .B(net239),
    .Y(_1869_));
 sg13g2_a22oi_1 _3163_ (.Y(_1880_),
    .B1(_1869_),
    .B2(_0034_),
    .A2(_1847_),
    .A1(_1836_));
 sg13g2_nand2_1 _3164_ (.Y(_1891_),
    .A(net237),
    .B(_1869_));
 sg13g2_o21ai_1 _3165_ (.B1(_1891_),
    .Y(_1902_),
    .A1(net237),
    .A2(net217));
 sg13g2_nor2_1 _3166_ (.A(net238),
    .B(net215),
    .Y(_1913_));
 sg13g2_a221oi_1 _3167_ (.B2(_1869_),
    .C1(net214),
    .B1(_1913_),
    .A1(net238),
    .Y(_1924_),
    .A2(_1902_));
 sg13g2_a21oi_1 _3168_ (.A1(net214),
    .A2(_1880_),
    .Y(_1935_),
    .B1(_1924_));
 sg13g2_a21oi_1 _3169_ (.A1(_1836_),
    .A2(_1748_),
    .Y(_1946_),
    .B1(_1726_));
 sg13g2_nand2_1 _3170_ (.Y(_1957_),
    .A(net213),
    .B(_1946_));
 sg13g2_o21ai_1 _3171_ (.B1(_1957_),
    .Y(_1968_),
    .A1(_1825_),
    .A2(_1935_));
 sg13g2_o21ai_1 _3172_ (.B1(_1968_),
    .Y(_1979_),
    .A1(_1671_),
    .A2(_1814_));
 sg13g2_xor2_1 _3173_ (.B(_1979_),
    .A(_0010_),
    .X(_1990_));
 sg13g2_nor2b_1 _3174_ (.A(net238),
    .B_N(_1704_),
    .Y(_2001_));
 sg13g2_buf_1 _3175_ (.A(_2001_),
    .X(_2012_));
 sg13g2_nor2_1 _3176_ (.A(_1704_),
    .B(_1858_),
    .Y(_2023_));
 sg13g2_nand2_1 _3177_ (.Y(_2034_),
    .A(_1836_),
    .B(_2023_));
 sg13g2_nor2_1 _3178_ (.A(_1704_),
    .B(_1649_),
    .Y(_2045_));
 sg13g2_and2_1 _3179_ (.A(_1704_),
    .B(_1638_),
    .X(_2056_));
 sg13g2_buf_1 _3180_ (.A(_2056_),
    .X(_2067_));
 sg13g2_o21ai_1 _3181_ (.B1(net216),
    .Y(_2078_),
    .A1(_2045_),
    .A2(_2067_));
 sg13g2_a21oi_1 _3182_ (.A1(_2034_),
    .A2(_2078_),
    .Y(_2089_),
    .B1(net215));
 sg13g2_a21oi_1 _3183_ (.A1(_1869_),
    .A2(_2012_),
    .Y(_2100_),
    .B1(_2089_));
 sg13g2_nand3_1 _3184_ (.B(net213),
    .C(_0007_),
    .A(net216),
    .Y(_2111_));
 sg13g2_o21ai_1 _3185_ (.B1(_2111_),
    .Y(_2122_),
    .A1(net213),
    .A2(_2100_));
 sg13g2_xor2_1 _3186_ (.B(_2122_),
    .A(_0012_),
    .X(_2133_));
 sg13g2_nand2_1 _3187_ (.Y(_2144_),
    .A(_1792_),
    .B(net213));
 sg13g2_and2_1 _3188_ (.A(net238),
    .B(_1715_),
    .X(_2155_));
 sg13g2_buf_1 _3189_ (.A(_2155_),
    .X(_2166_));
 sg13g2_mux2_1 _3190_ (.A0(_2166_),
    .A1(_1836_),
    .S(_1671_),
    .X(_2177_));
 sg13g2_nor2_2 _3191_ (.A(_1858_),
    .B(_1737_),
    .Y(_2188_));
 sg13g2_nor2_1 _3192_ (.A(net216),
    .B(_0007_),
    .Y(_2199_));
 sg13g2_nand4_1 _3193_ (.B(_0008_),
    .C(_2188_),
    .A(net215),
    .Y(_2210_),
    .D(_2199_));
 sg13g2_o21ai_1 _3194_ (.B1(_2210_),
    .Y(_2221_),
    .A1(_2144_),
    .A2(_2177_));
 sg13g2_xnor2_1 _3195_ (.Y(_2230_),
    .A(_0009_),
    .B(_2221_));
 sg13g2_nand2_1 _3196_ (.Y(_2241_),
    .A(net237),
    .B(net239));
 sg13g2_nor2_1 _3197_ (.A(net217),
    .B(_1737_),
    .Y(_2252_));
 sg13g2_a22oi_1 _3198_ (.Y(_2262_),
    .B1(_2252_),
    .B2(_2199_),
    .A2(_2023_),
    .A1(net216));
 sg13g2_nand2b_1 _3199_ (.Y(_2272_),
    .B(_1737_),
    .A_N(net214));
 sg13g2_xor2_1 _3200_ (.B(net217),
    .A(net237),
    .X(_2283_));
 sg13g2_a221oi_1 _3201_ (.B2(_2283_),
    .C1(net239),
    .B1(_2012_),
    .A1(net217),
    .Y(_2294_),
    .A2(_2166_));
 sg13g2_or2_1 _3202_ (.X(_2305_),
    .B(_2294_),
    .A(_1737_));
 sg13g2_o21ai_1 _3203_ (.B1(_2305_),
    .Y(_2316_),
    .A1(_2166_),
    .A2(_2272_));
 sg13g2_o21ai_1 _3204_ (.B1(_2316_),
    .Y(_2327_),
    .A1(_2241_),
    .A2(_2262_));
 sg13g2_xnor2_1 _3205_ (.Y(_2338_),
    .A(_0011_),
    .B(_2327_));
 sg13g2_buf_1 _3206_ (.A(\audio_engine_1.freq_synth1.hp_ctr[0] ),
    .X(_2349_));
 sg13g2_and3_1 _3207_ (.X(_2360_),
    .A(_1792_),
    .B(net217),
    .C(net239));
 sg13g2_nor2_1 _3208_ (.A(_1836_),
    .B(_2360_),
    .Y(_2371_));
 sg13g2_a21oi_1 _3209_ (.A1(_0034_),
    .A2(_2360_),
    .Y(_2382_),
    .B1(_2371_));
 sg13g2_nor2_1 _3210_ (.A(net238),
    .B(_1858_),
    .Y(_2393_));
 sg13g2_a21oi_1 _3211_ (.A1(net238),
    .A2(_2045_),
    .Y(_2404_),
    .B1(_2393_));
 sg13g2_nor2_1 _3212_ (.A(net215),
    .B(_2404_),
    .Y(_2415_));
 sg13g2_nor4_1 _3213_ (.A(net239),
    .B(_1737_),
    .C(_2415_),
    .D(_2067_),
    .Y(_2426_));
 sg13g2_a21oi_1 _3214_ (.A1(net213),
    .A2(_2382_),
    .Y(_2436_),
    .B1(_2426_));
 sg13g2_xor2_1 _3215_ (.B(_2436_),
    .A(_2349_),
    .X(_2444_));
 sg13g2_nand2_1 _3216_ (.Y(_2445_),
    .A(_0007_),
    .B(_2166_));
 sg13g2_nor2b_1 _3217_ (.A(net217),
    .B_N(_0007_),
    .Y(_2446_));
 sg13g2_o21ai_1 _3218_ (.B1(net238),
    .Y(_2447_),
    .A1(_2067_),
    .A2(_2446_));
 sg13g2_a21oi_1 _3219_ (.A1(_2034_),
    .A2(_2447_),
    .Y(_2448_),
    .B1(net215));
 sg13g2_a22oi_1 _3220_ (.Y(_2449_),
    .B1(_2012_),
    .B2(_1858_),
    .A2(_2023_),
    .A1(net238));
 sg13g2_nand2_1 _3221_ (.Y(_2450_),
    .A(_1869_),
    .B(_2012_));
 sg13g2_o21ai_1 _3222_ (.B1(_2450_),
    .Y(_2451_),
    .A1(_2241_),
    .A2(_2449_));
 sg13g2_nor3_1 _3223_ (.A(net213),
    .B(_2448_),
    .C(_2451_),
    .Y(_2452_));
 sg13g2_a21oi_1 _3224_ (.A1(net213),
    .A2(_2445_),
    .Y(_2453_),
    .B1(_2452_));
 sg13g2_xor2_1 _3225_ (.B(_2453_),
    .A(_0014_),
    .X(_2454_));
 sg13g2_nand4_1 _3226_ (.B(_2338_),
    .C(_2444_),
    .A(_2230_),
    .Y(_2455_),
    .D(_2454_));
 sg13g2_buf_1 _3227_ (.A(\audio_engine_1.freq_synth1.hp_ctr[1] ),
    .X(_2456_));
 sg13g2_a21oi_1 _3228_ (.A1(_1704_),
    .A2(_2188_),
    .Y(_2457_),
    .B1(_2045_));
 sg13g2_nor2_1 _3229_ (.A(_1781_),
    .B(_2457_),
    .Y(_2458_));
 sg13g2_a21oi_1 _3230_ (.A1(_1726_),
    .A2(_2188_),
    .Y(_2459_),
    .B1(_2458_));
 sg13g2_nor2_1 _3231_ (.A(net237),
    .B(net214),
    .Y(_2460_));
 sg13g2_a221oi_1 _3232_ (.B2(_2460_),
    .C1(net216),
    .B1(_2188_),
    .A1(net214),
    .Y(_2461_),
    .A2(_1847_));
 sg13g2_a21oi_1 _3233_ (.A1(net216),
    .A2(_2459_),
    .Y(_2462_),
    .B1(_2461_));
 sg13g2_nor2b_1 _3234_ (.A(_2462_),
    .B_N(net239),
    .Y(_2463_));
 sg13g2_mux2_1 _3235_ (.A0(_2188_),
    .A1(_1737_),
    .S(_1781_),
    .X(_2464_));
 sg13g2_a21oi_1 _3236_ (.A1(_2012_),
    .A2(_2464_),
    .Y(_2465_),
    .B1(_1660_));
 sg13g2_nand3_1 _3237_ (.B(net213),
    .C(_2460_),
    .A(_1693_),
    .Y(_2466_));
 sg13g2_o21ai_1 _3238_ (.B1(_2466_),
    .Y(_2467_),
    .A1(_2463_),
    .A2(_2465_));
 sg13g2_xnor2_1 _3239_ (.Y(_2468_),
    .A(_2456_),
    .B(_2467_));
 sg13g2_nor4_1 _3240_ (.A(_1990_),
    .B(_2133_),
    .C(_2455_),
    .D(_2468_),
    .Y(_2469_));
 sg13g2_buf_2 _3241_ (.A(_2469_),
    .X(_2470_));
 sg13g2_nand3_1 _3242_ (.B(_1627_),
    .C(_2470_),
    .A(\audio_engine_1.freq_synth1.en_synth_clk ),
    .Y(_2471_));
 sg13g2_mux2_1 _3243_ (.A0(_0002_),
    .A1(\audio_engine_1.freq_synth1.audio_reg ),
    .S(_2471_),
    .X(_0058_));
 sg13g2_nand2_2 _3244_ (.Y(_2472_),
    .A(\audio_engine_1.freq_synth1.en_synth_clk ),
    .B(_1627_));
 sg13g2_buf_1 _3245_ (.A(_2472_),
    .X(_2473_));
 sg13g2_nand2b_1 _3246_ (.Y(_2474_),
    .B(_2349_),
    .A_N(_2470_));
 sg13g2_nand2_1 _3247_ (.Y(_2475_),
    .A(_0036_),
    .B(net188));
 sg13g2_o21ai_1 _3248_ (.B1(_2475_),
    .Y(_0059_),
    .A1(net188),
    .A2(_2474_));
 sg13g2_or2_1 _3249_ (.X(_2476_),
    .B(_2472_),
    .A(_2456_));
 sg13g2_nor2_1 _3250_ (.A(_2349_),
    .B(_2470_),
    .Y(_2477_));
 sg13g2_o21ai_1 _3251_ (.B1(_2456_),
    .Y(_2478_),
    .A1(net188),
    .A2(_2477_));
 sg13g2_o21ai_1 _3252_ (.B1(_2478_),
    .Y(_0060_),
    .A1(_2474_),
    .A2(_2476_));
 sg13g2_nand2_1 _3253_ (.Y(_2479_),
    .A(_2349_),
    .B(_2456_));
 sg13g2_xnor2_1 _3254_ (.Y(_2480_),
    .A(_0009_),
    .B(_2479_));
 sg13g2_nor3_1 _3255_ (.A(_2470_),
    .B(_2473_),
    .C(_2480_),
    .Y(_2481_));
 sg13g2_a21o_1 _3256_ (.A2(_2473_),
    .A1(\audio_engine_1.freq_synth1.hp_ctr[2] ),
    .B1(_2481_),
    .X(_0061_));
 sg13g2_nand3_1 _3257_ (.B(_2456_),
    .C(\audio_engine_1.freq_synth1.hp_ctr[2] ),
    .A(_2349_),
    .Y(_2482_));
 sg13g2_xnor2_1 _3258_ (.Y(_2483_),
    .A(_0010_),
    .B(_2482_));
 sg13g2_nor3_1 _3259_ (.A(_2470_),
    .B(net188),
    .C(_2483_),
    .Y(_2484_));
 sg13g2_a21o_1 _3260_ (.A2(net188),
    .A1(\audio_engine_1.freq_synth1.hp_ctr[3] ),
    .B1(_2484_),
    .X(_0062_));
 sg13g2_inv_1 _3261_ (.Y(_2485_),
    .A(\audio_engine_1.freq_synth1.hp_ctr[3] ));
 sg13g2_nor2_1 _3262_ (.A(_2485_),
    .B(_2482_),
    .Y(_2486_));
 sg13g2_xor2_1 _3263_ (.B(_2486_),
    .A(_0011_),
    .X(_2487_));
 sg13g2_nor3_1 _3264_ (.A(_2470_),
    .B(_2472_),
    .C(_2487_),
    .Y(_2488_));
 sg13g2_a21o_1 _3265_ (.A2(net188),
    .A1(\audio_engine_1.freq_synth1.hp_ctr[4] ),
    .B1(_2488_),
    .X(_0063_));
 sg13g2_nand2_1 _3266_ (.Y(_2489_),
    .A(\audio_engine_1.freq_synth1.hp_ctr[4] ),
    .B(_2486_));
 sg13g2_xnor2_1 _3267_ (.Y(_2490_),
    .A(_0012_),
    .B(_2489_));
 sg13g2_nor3_1 _3268_ (.A(_2470_),
    .B(_2472_),
    .C(_2490_),
    .Y(_2491_));
 sg13g2_a21o_1 _3269_ (.A2(net188),
    .A1(\audio_engine_1.freq_synth1.hp_ctr[5] ),
    .B1(_2491_),
    .X(_0064_));
 sg13g2_nand3_1 _3270_ (.B(\audio_engine_1.freq_synth1.hp_ctr[5] ),
    .C(_2486_),
    .A(\audio_engine_1.freq_synth1.hp_ctr[4] ),
    .Y(_2492_));
 sg13g2_xnor2_1 _3271_ (.Y(_2493_),
    .A(_0014_),
    .B(_2492_));
 sg13g2_nor3_1 _3272_ (.A(_2470_),
    .B(_2472_),
    .C(_2493_),
    .Y(_2494_));
 sg13g2_a21o_1 _3273_ (.A2(net188),
    .A1(\audio_engine_1.freq_synth1.hp_ctr[6] ),
    .B1(_2494_),
    .X(_0065_));
 sg13g2_buf_2 _3274_ (.A(\audio_engine_1.seq_ctr[0] ),
    .X(_2495_));
 sg13g2_buf_1 _3275_ (.A(\audio_engine_1.counter[17] ),
    .X(_2496_));
 sg13g2_nand2_2 _3276_ (.Y(_2497_),
    .A(_2496_),
    .B(\audio_engine_1.en_seq_clk ));
 sg13g2_xnor2_1 _3277_ (.Y(_0066_),
    .A(_2495_),
    .B(_2497_));
 sg13g2_buf_1 _3278_ (.A(\audio_engine_1.seq_ctr[1] ),
    .X(_2498_));
 sg13g2_nand3_1 _3279_ (.B(\audio_engine_1.en_seq_clk ),
    .C(_2495_),
    .A(_2496_),
    .Y(_2499_));
 sg13g2_xnor2_1 _3280_ (.Y(_0067_),
    .A(_2498_),
    .B(_2499_));
 sg13g2_buf_2 _3281_ (.A(\audio_engine_1.seq_ctr[2] ),
    .X(_2500_));
 sg13g2_nand4_1 _3282_ (.B(\audio_engine_1.en_seq_clk ),
    .C(_2498_),
    .A(_2496_),
    .Y(_2501_),
    .D(_2495_));
 sg13g2_buf_2 _3283_ (.A(\audio_engine_1.seq_ctr[3] ),
    .X(_2502_));
 sg13g2_buf_1 _3284_ (.A(_0006_),
    .X(_2503_));
 sg13g2_nor2_1 _3285_ (.A(_2502_),
    .B(_2503_),
    .Y(_2504_));
 sg13g2_nor3_1 _3286_ (.A(_2500_),
    .B(_2501_),
    .C(_2504_),
    .Y(_2505_));
 sg13g2_a21o_1 _3287_ (.A2(_2501_),
    .A1(_2500_),
    .B1(_2505_),
    .X(_0068_));
 sg13g2_nand2_1 _3288_ (.Y(_2506_),
    .A(_2498_),
    .B(_2500_));
 sg13g2_nor3_1 _3289_ (.A(_0015_),
    .B(_2497_),
    .C(_2506_),
    .Y(_2507_));
 sg13g2_xor2_1 _3290_ (.B(_2507_),
    .A(_2502_),
    .X(_0069_));
 sg13g2_nand4_1 _3291_ (.B(_2495_),
    .C(_2500_),
    .A(_2498_),
    .Y(_2508_),
    .D(_2503_));
 sg13g2_o21ai_1 _3292_ (.B1(_2508_),
    .Y(_2509_),
    .A1(_2500_),
    .A2(_2503_));
 sg13g2_nand2b_1 _3293_ (.Y(_2510_),
    .B(_2500_),
    .A_N(_2502_));
 sg13g2_nand3_1 _3294_ (.B(_2495_),
    .C(_2510_),
    .A(_2498_),
    .Y(_2511_));
 sg13g2_inv_1 _3295_ (.Y(_2512_),
    .A(_2503_));
 sg13g2_a22oi_1 _3296_ (.Y(_2513_),
    .B1(_2511_),
    .B2(_2512_),
    .A2(_2509_),
    .A1(_2502_));
 sg13g2_nand2_1 _3297_ (.Y(_2514_),
    .A(\audio_engine_1.seq_ctr[4] ),
    .B(_2497_));
 sg13g2_o21ai_1 _3298_ (.B1(_2514_),
    .Y(_0070_),
    .A1(_2497_),
    .A2(_2513_));
 sg13g2_nor4_2 _3299_ (.A(_2502_),
    .B(_2500_),
    .C(_2503_),
    .Y(_2515_),
    .D(_2501_));
 sg13g2_mux2_1 _3300_ (.A0(net215),
    .A1(_0034_),
    .S(_2515_),
    .X(_0071_));
 sg13g2_nand2_1 _3301_ (.Y(_2516_),
    .A(net215),
    .B(_2515_));
 sg13g2_xnor2_1 _3302_ (.Y(_0072_),
    .A(net216),
    .B(_2516_));
 sg13g2_nand2_1 _3303_ (.Y(_2517_),
    .A(_2166_),
    .B(_2515_));
 sg13g2_xnor2_1 _3304_ (.Y(_0073_),
    .A(net214),
    .B(_2517_));
 sg13g2_nand3_1 _3305_ (.B(_2166_),
    .C(_2515_),
    .A(net214),
    .Y(_2518_));
 sg13g2_xnor2_1 _3306_ (.Y(_0074_),
    .A(net217),
    .B(_2518_));
 sg13g2_nor2_1 _3307_ (.A(_1858_),
    .B(_2518_),
    .Y(_2519_));
 sg13g2_xor2_1 _3308_ (.B(_2519_),
    .A(net239),
    .X(_0075_));
 sg13g2_nor2_1 _3309_ (.A(_1671_),
    .B(_2518_),
    .Y(_2520_));
 sg13g2_xor2_1 _3310_ (.B(_2520_),
    .A(\audio_engine_1.seq_time[5] ),
    .X(_0076_));
 sg13g2_nand2_1 _3311_ (.Y(_2521_),
    .A(\audio_engine_1.seq_time[5] ),
    .B(_2520_));
 sg13g2_xnor2_1 _3312_ (.Y(_0077_),
    .A(_1825_),
    .B(_2521_));
 sg13g2_buf_8 _3313_ (.A(\graphics_engine_1.ctr[0] ),
    .X(_2522_));
 sg13g2_inv_1 _3314_ (.Y(_2523_),
    .A(net7));
 sg13g2_nand3_1 _3315_ (.B(\graphics_engine_1.en_v_sync ),
    .C(\graphics_engine_1.v_sync ),
    .A(_2523_),
    .Y(_2524_));
 sg13g2_mux2_1 _3316_ (.A0(_0035_),
    .A1(_2522_),
    .S(_2524_),
    .X(_0078_));
 sg13g2_buf_8 _3317_ (.A(\graphics_engine_1.ctr[1] ),
    .X(_2525_));
 sg13g2_buf_1 _3318_ (.A(_2525_),
    .X(_2526_));
 sg13g2_inv_1 _3319_ (.Y(_2527_),
    .A(_2522_));
 sg13g2_nor2_1 _3320_ (.A(_2527_),
    .B(_2524_),
    .Y(_2528_));
 sg13g2_xor2_1 _3321_ (.B(_2528_),
    .A(net212),
    .X(_0079_));
 sg13g2_buf_2 _3322_ (.A(\graphics_engine_1.ctr[2] ),
    .X(_2529_));
 sg13g2_buf_1 _3323_ (.A(net235),
    .X(_2530_));
 sg13g2_and2_1 _3324_ (.A(net212),
    .B(_2528_),
    .X(_2531_));
 sg13g2_xor2_1 _3325_ (.B(_2531_),
    .A(net211),
    .X(_0080_));
 sg13g2_buf_1 _3326_ (.A(\graphics_engine_1.ctr[3] ),
    .X(_2532_));
 sg13g2_buf_1 _3327_ (.A(_2532_),
    .X(_2533_));
 sg13g2_buf_1 _3328_ (.A(net210),
    .X(_2534_));
 sg13g2_nand2_1 _3329_ (.Y(_2535_),
    .A(net211),
    .B(_2531_));
 sg13g2_xnor2_1 _3330_ (.Y(_0081_),
    .A(net187),
    .B(_2535_));
 sg13g2_buf_1 _3331_ (.A(\graphics_engine_1.ctr[4] ),
    .X(_2536_));
 sg13g2_inv_1 _3332_ (.Y(_2537_),
    .A(net234));
 sg13g2_inv_1 _3333_ (.Y(_2538_),
    .A(net210));
 sg13g2_buf_1 _3334_ (.A(_2538_),
    .X(_2539_));
 sg13g2_nor2_1 _3335_ (.A(net166),
    .B(_2535_),
    .Y(_2540_));
 sg13g2_xnor2_1 _3336_ (.Y(_0082_),
    .A(_2537_),
    .B(_2540_));
 sg13g2_buf_1 _3337_ (.A(\graphics_engine_1.ctr[5] ),
    .X(_2541_));
 sg13g2_buf_1 _3338_ (.A(_2541_),
    .X(_2542_));
 sg13g2_buf_1 _3339_ (.A(net234),
    .X(_2543_));
 sg13g2_nand2_1 _3340_ (.Y(_2544_),
    .A(net208),
    .B(_2540_));
 sg13g2_xnor2_1 _3341_ (.Y(_0083_),
    .A(net209),
    .B(_2544_));
 sg13g2_buf_1 _3342_ (.A(\graphics_engine_1.ctr[6] ),
    .X(_2545_));
 sg13g2_nand3_1 _3343_ (.B(_2542_),
    .C(_2540_),
    .A(net208),
    .Y(_2546_));
 sg13g2_xnor2_1 _3344_ (.Y(_0084_),
    .A(net232),
    .B(_2546_));
 sg13g2_buf_1 _3345_ (.A(\graphics_engine_1.ctr[7] ),
    .X(_2547_));
 sg13g2_inv_1 _3346_ (.Y(_2548_),
    .A(net209));
 sg13g2_inv_1 _3347_ (.Y(_2549_),
    .A(_2545_));
 sg13g2_nor3_1 _3348_ (.A(_2548_),
    .B(_2549_),
    .C(_2544_),
    .Y(_2550_));
 sg13g2_xor2_1 _3349_ (.B(_2550_),
    .A(_2547_),
    .X(_0085_));
 sg13g2_nand2_1 _3350_ (.Y(_2551_),
    .A(_2547_),
    .B(_2550_));
 sg13g2_xnor2_1 _3351_ (.Y(_0086_),
    .A(\graphics_engine_1.ctr[8] ),
    .B(_2551_));
 sg13g2_buf_2 _3352_ (.A(net247),
    .X(_2552_));
 sg13g2_inv_1 _3353_ (.Y(_2553_),
    .A(net244));
 sg13g2_buf_1 _3354_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ),
    .X(_2554_));
 sg13g2_buf_1 _3355_ (.A(net221),
    .X(_2555_));
 sg13g2_nand2_2 _3356_ (.Y(_2556_),
    .A(net186),
    .B(net169));
 sg13g2_or2_1 _3357_ (.X(_2557_),
    .B(net225),
    .A(net222));
 sg13g2_buf_1 _3358_ (.A(_2557_),
    .X(_2558_));
 sg13g2_nor4_1 _3359_ (.A(net242),
    .B(net231),
    .C(_2556_),
    .D(_2558_),
    .Y(_2559_));
 sg13g2_nor2_1 _3360_ (.A(net245),
    .B(_1134_),
    .Y(_2560_));
 sg13g2_nand4_1 _3361_ (.B(_1068_),
    .C(_2559_),
    .A(_2553_),
    .Y(_2561_),
    .D(_2560_));
 sg13g2_nand2_1 _3362_ (.Y(_2562_),
    .A(_2552_),
    .B(_2561_));
 sg13g2_buf_1 _3363_ (.A(_2562_),
    .X(_2563_));
 sg13g2_inv_2 _3364_ (.Y(_2564_),
    .A(_1430_));
 sg13g2_buf_1 _3365_ (.A(net185),
    .X(_2565_));
 sg13g2_buf_1 _3366_ (.A(net165),
    .X(_2566_));
 sg13g2_buf_2 _3367_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[2] ),
    .X(_2567_));
 sg13g2_buf_1 _3368_ (.A(_2567_),
    .X(_2568_));
 sg13g2_buf_1 _3369_ (.A(_2568_),
    .X(_2569_));
 sg13g2_buf_2 _3370_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_x[0] ),
    .X(_2570_));
 sg13g2_buf_1 _3371_ (.A(_2570_),
    .X(_2571_));
 sg13g2_buf_1 _3372_ (.A(net206),
    .X(_2572_));
 sg13g2_nand2_1 _3373_ (.Y(_2573_),
    .A(net184),
    .B(net183));
 sg13g2_buf_2 _3374_ (.A(_2573_),
    .X(_2574_));
 sg13g2_buf_1 _3375_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ),
    .X(_2575_));
 sg13g2_buf_8 _3376_ (.A(\graphics_engine_1.anim_2x[0] ),
    .X(_2576_));
 sg13g2_nand2_1 _3377_ (.Y(_2577_),
    .A(net230),
    .B(_2576_));
 sg13g2_nor3_2 _3378_ (.A(net144),
    .B(_2574_),
    .C(_2577_),
    .Y(_2578_));
 sg13g2_nor2_1 _3379_ (.A(_1408_),
    .B(net220),
    .Y(_2579_));
 sg13g2_buf_1 _3380_ (.A(net240),
    .X(_2580_));
 sg13g2_nor2b_1 _3381_ (.A(net205),
    .B_N(\graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ),
    .Y(_2581_));
 sg13g2_and4_1 _3382_ (.A(_1507_),
    .B(_2578_),
    .C(_2579_),
    .D(_2581_),
    .X(_2582_));
 sg13g2_buf_1 _3383_ (.A(_2582_),
    .X(_2583_));
 sg13g2_nand2_1 _3384_ (.Y(_2584_),
    .A(_0031_),
    .B(_2583_));
 sg13g2_nand3b_1 _3385_ (.B(net231),
    .C(_2552_),
    .Y(_2585_),
    .A_N(_2583_));
 sg13g2_o21ai_1 _3386_ (.B1(_2585_),
    .Y(_0098_),
    .A1(net67),
    .A2(_2584_));
 sg13g2_nand2_1 _3387_ (.Y(_2586_),
    .A(net231),
    .B(_2583_));
 sg13g2_xnor2_1 _3388_ (.Y(_2587_),
    .A(net242),
    .B(_2586_));
 sg13g2_and2_1 _3389_ (.A(_2552_),
    .B(_2587_),
    .X(_0099_));
 sg13g2_nor2b_1 _3390_ (.A(_2583_),
    .B_N(_2552_),
    .Y(_2588_));
 sg13g2_buf_1 _3391_ (.A(_2588_),
    .X(_2589_));
 sg13g2_nor2_1 _3392_ (.A(net67),
    .B(_2589_),
    .Y(_2590_));
 sg13g2_buf_2 _3393_ (.A(_2590_),
    .X(_2591_));
 sg13g2_nand4_1 _3394_ (.B(net231),
    .C(_1332_),
    .A(net242),
    .Y(_2592_),
    .D(_2591_));
 sg13g2_a21oi_1 _3395_ (.A1(net242),
    .A2(net231),
    .Y(_2593_),
    .B1(_2563_));
 sg13g2_o21ai_1 _3396_ (.B1(net186),
    .Y(_2594_),
    .A1(_2589_),
    .A2(_2593_));
 sg13g2_nand2_1 _3397_ (.Y(_0100_),
    .A(_2592_),
    .B(_2594_));
 sg13g2_buf_1 _3398_ (.A(net169),
    .X(_2595_));
 sg13g2_and3_1 _3399_ (.X(_2596_),
    .A(net242),
    .B(net231),
    .C(net186));
 sg13g2_buf_1 _3400_ (.A(_2596_),
    .X(_2597_));
 sg13g2_nand2_1 _3401_ (.Y(_2598_),
    .A(_2591_),
    .B(_2597_));
 sg13g2_nand2b_1 _3402_ (.Y(_2599_),
    .B(_2552_),
    .A_N(_2583_));
 sg13g2_buf_1 _3403_ (.A(_2599_),
    .X(_2600_));
 sg13g2_o21ai_1 _3404_ (.B1(net54),
    .Y(_2601_),
    .A1(_2563_),
    .A2(_2597_));
 sg13g2_nand2_1 _3405_ (.Y(_2602_),
    .A(net143),
    .B(_2601_));
 sg13g2_o21ai_1 _3406_ (.B1(_2602_),
    .Y(_0101_),
    .A1(net143),
    .A2(_2598_));
 sg13g2_a21oi_1 _3407_ (.A1(net143),
    .A2(_2597_),
    .Y(_2603_),
    .B1(net67));
 sg13g2_buf_1 _3408_ (.A(net192),
    .X(_2604_));
 sg13g2_buf_1 _3409_ (.A(net164),
    .X(_2605_));
 sg13g2_buf_1 _3410_ (.A(net142),
    .X(_2606_));
 sg13g2_o21ai_1 _3411_ (.B1(net120),
    .Y(_2607_),
    .A1(_2589_),
    .A2(_2603_));
 sg13g2_o21ai_1 _3412_ (.B1(_2607_),
    .Y(_0102_),
    .A1(_1288_),
    .A2(_2598_));
 sg13g2_buf_1 _3413_ (.A(net194),
    .X(_2608_));
 sg13g2_buf_1 _3414_ (.A(net163),
    .X(_2609_));
 sg13g2_buf_1 _3415_ (.A(net141),
    .X(_2610_));
 sg13g2_and2_1 _3416_ (.A(net193),
    .B(net164),
    .X(_2611_));
 sg13g2_buf_2 _3417_ (.A(_2611_),
    .X(_2612_));
 sg13g2_and2_1 _3418_ (.A(_2597_),
    .B(_2612_),
    .X(_2613_));
 sg13g2_buf_1 _3419_ (.A(_2613_),
    .X(_2614_));
 sg13g2_nand2_1 _3420_ (.Y(_2615_),
    .A(_2591_),
    .B(_2614_));
 sg13g2_o21ai_1 _3421_ (.B1(net54),
    .Y(_2616_),
    .A1(net67),
    .A2(_2614_));
 sg13g2_nand2_1 _3422_ (.Y(_2617_),
    .A(net119),
    .B(_2616_));
 sg13g2_o21ai_1 _3423_ (.B1(_2617_),
    .Y(_0103_),
    .A1(net119),
    .A2(_2615_));
 sg13g2_buf_1 _3424_ (.A(net224),
    .X(_2618_));
 sg13g2_buf_1 _3425_ (.A(net182),
    .X(_2619_));
 sg13g2_buf_1 _3426_ (.A(net162),
    .X(_2620_));
 sg13g2_buf_1 _3427_ (.A(net140),
    .X(_2621_));
 sg13g2_and2_1 _3428_ (.A(net119),
    .B(_2614_),
    .X(_2622_));
 sg13g2_buf_1 _3429_ (.A(_2622_),
    .X(_2623_));
 sg13g2_nand2_1 _3430_ (.Y(_2624_),
    .A(_2591_),
    .B(_2623_));
 sg13g2_o21ai_1 _3431_ (.B1(net54),
    .Y(_2625_),
    .A1(net67),
    .A2(_2623_));
 sg13g2_nand2_1 _3432_ (.Y(_2626_),
    .A(net118),
    .B(_2625_));
 sg13g2_o21ai_1 _3433_ (.B1(_2626_),
    .Y(_0104_),
    .A1(net118),
    .A2(_2624_));
 sg13g2_and2_1 _3434_ (.A(net118),
    .B(_2623_),
    .X(_2627_));
 sg13g2_buf_1 _3435_ (.A(_2627_),
    .X(_2628_));
 sg13g2_nand2_1 _3436_ (.Y(_2629_),
    .A(_2591_),
    .B(_2628_));
 sg13g2_o21ai_1 _3437_ (.B1(net54),
    .Y(_2630_),
    .A1(net67),
    .A2(_2628_));
 sg13g2_nand2_1 _3438_ (.Y(_2631_),
    .A(net245),
    .B(_2630_));
 sg13g2_o21ai_1 _3439_ (.B1(_2631_),
    .Y(_0105_),
    .A1(net245),
    .A2(_2629_));
 sg13g2_and2_1 _3440_ (.A(net245),
    .B(_2628_),
    .X(_2632_));
 sg13g2_buf_1 _3441_ (.A(_2632_),
    .X(_2633_));
 sg13g2_nand2_1 _3442_ (.Y(_2634_),
    .A(_2591_),
    .B(_2633_));
 sg13g2_o21ai_1 _3443_ (.B1(_2599_),
    .Y(_2635_),
    .A1(net67),
    .A2(_2633_));
 sg13g2_nand2_1 _3444_ (.Y(_2636_),
    .A(net244),
    .B(_2635_));
 sg13g2_o21ai_1 _3445_ (.B1(_2636_),
    .Y(_0106_),
    .A1(net244),
    .A2(_2634_));
 sg13g2_nand3_1 _3446_ (.B(_2591_),
    .C(_2633_),
    .A(net244),
    .Y(_2637_));
 sg13g2_a21oi_1 _3447_ (.A1(net244),
    .A2(_2633_),
    .Y(_2638_),
    .B1(net67));
 sg13g2_o21ai_1 _3448_ (.B1(_1068_),
    .Y(_2639_),
    .A1(_2589_),
    .A2(_2638_));
 sg13g2_o21ai_1 _3449_ (.B1(_2639_),
    .Y(_0107_),
    .A1(_1068_),
    .A2(_2637_));
 sg13g2_mux2_1 _3450_ (.A0(_0033_),
    .A1(\audio_engine_1.counter[0] ),
    .S(net8),
    .X(_0040_));
 sg13g2_inv_1 _3451_ (.Y(_2640_),
    .A(\audio_engine_1.counter[7] ));
 sg13g2_nor2b_1 _3452_ (.A(net8),
    .B_N(\audio_engine_1.counter[0] ),
    .Y(_2641_));
 sg13g2_and3_1 _3453_ (.X(_2642_),
    .A(\audio_engine_1.counter[1] ),
    .B(\audio_engine_1.counter[2] ),
    .C(_2641_));
 sg13g2_buf_1 _3454_ (.A(_2642_),
    .X(_2643_));
 sg13g2_and3_1 _3455_ (.X(_2644_),
    .A(\audio_engine_1.counter[3] ),
    .B(\audio_engine_1.counter[4] ),
    .C(_2643_));
 sg13g2_buf_1 _3456_ (.A(_2644_),
    .X(_2645_));
 sg13g2_nand3_1 _3457_ (.B(\audio_engine_1.counter[6] ),
    .C(_2645_),
    .A(\audio_engine_1.counter[5] ),
    .Y(_2646_));
 sg13g2_nor2_1 _3458_ (.A(_2640_),
    .B(_2646_),
    .Y(_2647_));
 sg13g2_nand3_1 _3459_ (.B(\audio_engine_1.counter[9] ),
    .C(_2647_),
    .A(\audio_engine_1.counter[8] ),
    .Y(_2648_));
 sg13g2_xnor2_1 _3460_ (.Y(_0041_),
    .A(_1627_),
    .B(_2648_));
 sg13g2_inv_1 _3461_ (.Y(_2649_),
    .A(_1627_));
 sg13g2_nor2_1 _3462_ (.A(_2649_),
    .B(_2648_),
    .Y(_2650_));
 sg13g2_xor2_1 _3463_ (.B(_2650_),
    .A(\audio_engine_1.counter[11] ),
    .X(_0042_));
 sg13g2_nand2_1 _3464_ (.Y(_2651_),
    .A(\audio_engine_1.counter[11] ),
    .B(_2650_));
 sg13g2_xnor2_1 _3465_ (.Y(_0043_),
    .A(\audio_engine_1.counter[12] ),
    .B(_2651_));
 sg13g2_nand3_1 _3466_ (.B(\audio_engine_1.counter[12] ),
    .C(_2650_),
    .A(\audio_engine_1.counter[11] ),
    .Y(_2652_));
 sg13g2_xnor2_1 _3467_ (.Y(_0044_),
    .A(\audio_engine_1.counter[13] ),
    .B(_2652_));
 sg13g2_buf_1 _3468_ (.A(\audio_engine_1.counter[14] ),
    .X(_2653_));
 sg13g2_inv_1 _3469_ (.Y(_2654_),
    .A(\audio_engine_1.counter[13] ));
 sg13g2_nor2_2 _3470_ (.A(_2654_),
    .B(_2652_),
    .Y(_2655_));
 sg13g2_xor2_1 _3471_ (.B(_2655_),
    .A(_2653_),
    .X(_0045_));
 sg13g2_nand2_1 _3472_ (.Y(_2656_),
    .A(_2653_),
    .B(_2655_));
 sg13g2_xnor2_1 _3473_ (.Y(_0046_),
    .A(\audio_engine_1.counter[15] ),
    .B(_2656_));
 sg13g2_nand3_1 _3474_ (.B(\audio_engine_1.counter[15] ),
    .C(_2655_),
    .A(_2653_),
    .Y(_2657_));
 sg13g2_xnor2_1 _3475_ (.Y(_0047_),
    .A(\audio_engine_1.counter[16] ),
    .B(_2657_));
 sg13g2_nand4_1 _3476_ (.B(\audio_engine_1.counter[15] ),
    .C(\audio_engine_1.counter[16] ),
    .A(_2653_),
    .Y(_2658_),
    .D(_2655_));
 sg13g2_xnor2_1 _3477_ (.Y(_0048_),
    .A(_2496_),
    .B(_2658_));
 sg13g2_xor2_1 _3478_ (.B(_2641_),
    .A(\audio_engine_1.counter[1] ),
    .X(_0049_));
 sg13g2_nand2_1 _3479_ (.Y(_2659_),
    .A(\audio_engine_1.counter[1] ),
    .B(_2641_));
 sg13g2_xnor2_1 _3480_ (.Y(_0050_),
    .A(\audio_engine_1.counter[2] ),
    .B(_2659_));
 sg13g2_xor2_1 _3481_ (.B(_2643_),
    .A(\audio_engine_1.counter[3] ),
    .X(_0051_));
 sg13g2_nand2_1 _3482_ (.Y(_2660_),
    .A(\audio_engine_1.counter[3] ),
    .B(_2643_));
 sg13g2_xnor2_1 _3483_ (.Y(_0052_),
    .A(\audio_engine_1.counter[4] ),
    .B(_2660_));
 sg13g2_xor2_1 _3484_ (.B(_2645_),
    .A(\audio_engine_1.counter[5] ),
    .X(_0053_));
 sg13g2_nand2_1 _3485_ (.Y(_2661_),
    .A(\audio_engine_1.counter[5] ),
    .B(_2645_));
 sg13g2_xnor2_1 _3486_ (.Y(_0054_),
    .A(\audio_engine_1.counter[6] ),
    .B(_2661_));
 sg13g2_xnor2_1 _3487_ (.Y(_0055_),
    .A(\audio_engine_1.counter[7] ),
    .B(_2646_));
 sg13g2_xor2_1 _3488_ (.B(_2647_),
    .A(\audio_engine_1.counter[8] ),
    .X(_0056_));
 sg13g2_nand2_1 _3489_ (.Y(_2662_),
    .A(\audio_engine_1.counter[8] ),
    .B(_2647_));
 sg13g2_xnor2_1 _3490_ (.Y(_0057_),
    .A(\audio_engine_1.counter[9] ),
    .B(_2662_));
 sg13g2_nor2_1 _3491_ (.A(_2523_),
    .B(_0037_),
    .Y(_2663_));
 sg13g2_a21oi_1 _3492_ (.A1(_2523_),
    .A2(_0003_),
    .Y(_0087_),
    .B1(_2663_));
 sg13g2_and2_1 _3493_ (.A(_0032_),
    .B(_2589_),
    .X(_0088_));
 sg13g2_xor2_1 _3494_ (.B(_2576_),
    .A(net230),
    .X(_2664_));
 sg13g2_and2_1 _3495_ (.A(_2552_),
    .B(_2664_),
    .X(_0089_));
 sg13g2_inv_2 _3496_ (.Y(_2665_),
    .A(net184));
 sg13g2_xnor2_1 _3497_ (.Y(_2666_),
    .A(_2665_),
    .B(_2577_));
 sg13g2_nor2_1 _3498_ (.A(net54),
    .B(_2666_),
    .Y(_0090_));
 sg13g2_inv_2 _3499_ (.Y(_2667_),
    .A(net206));
 sg13g2_buf_1 _3500_ (.A(_2667_),
    .X(_2668_));
 sg13g2_buf_1 _3501_ (.A(net161),
    .X(_2669_));
 sg13g2_buf_1 _3502_ (.A(_2569_),
    .X(_2670_));
 sg13g2_nand3_1 _3503_ (.B(_2576_),
    .C(net160),
    .A(net230),
    .Y(_2671_));
 sg13g2_xnor2_1 _3504_ (.Y(_2672_),
    .A(net139),
    .B(_2671_));
 sg13g2_nor2_1 _3505_ (.A(net54),
    .B(_2672_),
    .Y(_0091_));
 sg13g2_nor2_1 _3506_ (.A(_2574_),
    .B(_2577_),
    .Y(_2673_));
 sg13g2_xnor2_1 _3507_ (.Y(_2674_),
    .A(_2566_),
    .B(_2673_));
 sg13g2_and2_1 _3508_ (.A(_2552_),
    .B(_2674_),
    .X(_0092_));
 sg13g2_buf_1 _3509_ (.A(net191),
    .X(_2675_));
 sg13g2_buf_1 _3510_ (.A(net159),
    .X(_2676_));
 sg13g2_buf_1 _3511_ (.A(net138),
    .X(_2677_));
 sg13g2_xnor2_1 _3512_ (.Y(_2678_),
    .A(net117),
    .B(_2578_));
 sg13g2_nor2_1 _3513_ (.A(net54),
    .B(_2678_),
    .Y(_0093_));
 sg13g2_nand2_1 _3514_ (.Y(_2679_),
    .A(net117),
    .B(_2578_));
 sg13g2_xnor2_1 _3515_ (.Y(_2680_),
    .A(net168),
    .B(_2679_));
 sg13g2_and2_1 _3516_ (.A(_2552_),
    .B(_2680_),
    .X(_0094_));
 sg13g2_nand3_1 _3517_ (.B(_1551_),
    .C(_2578_),
    .A(net117),
    .Y(_2681_));
 sg13g2_xor2_1 _3518_ (.B(_2681_),
    .A(net205),
    .X(_2682_));
 sg13g2_nor2_1 _3519_ (.A(net54),
    .B(_2682_),
    .Y(_0095_));
 sg13g2_nand4_1 _3520_ (.B(_1551_),
    .C(_1584_),
    .A(_2580_),
    .Y(_2683_),
    .D(_2673_));
 sg13g2_xnor2_1 _3521_ (.Y(_2684_),
    .A(_1518_),
    .B(_2683_));
 sg13g2_nor2_1 _3522_ (.A(_2600_),
    .B(_2684_),
    .Y(_0096_));
 sg13g2_nand2_1 _3523_ (.Y(_2685_),
    .A(net205),
    .B(_1507_));
 sg13g2_or2_1 _3524_ (.X(_2686_),
    .B(_2685_),
    .A(_2681_));
 sg13g2_xor2_1 _3525_ (.B(_2686_),
    .A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ),
    .X(_2687_));
 sg13g2_nor2_1 _3526_ (.A(_2600_),
    .B(_2687_),
    .Y(_0097_));
 sg13g2_inv_1 _3527_ (.Y(_0038_),
    .A(_0000_));
 sg13g2_inv_1 _3528_ (.Y(_0039_),
    .A(_0001_));
 sg13g2_inv_1 _3529_ (.Y(_2688_),
    .A(\audio_engine_1.freq_synth1.audio_reg ));
 sg13g2_o21ai_1 _3530_ (.B1(_0015_),
    .Y(_2689_),
    .A1(_2495_),
    .A2(_2512_));
 sg13g2_a21oi_1 _3531_ (.A1(_2498_),
    .A2(_2689_),
    .Y(_2690_),
    .B1(_2500_));
 sg13g2_nor2b_1 _3532_ (.A(_2690_),
    .B_N(_2502_),
    .Y(_2691_));
 sg13g2_nor4_1 _3533_ (.A(\audio_engine_1.seq_ctr[4] ),
    .B(_2688_),
    .C(net8),
    .D(_2691_),
    .Y(audio));
 sg13g2_inv_1 _3534_ (.Y(_2692_),
    .A(_1068_));
 sg13g2_buf_1 _3535_ (.A(_0018_),
    .X(_2693_));
 sg13g2_inv_1 _3536_ (.Y(_2694_),
    .A(net229));
 sg13g2_buf_1 _3537_ (.A(_2694_),
    .X(_2695_));
 sg13g2_o21ai_1 _3538_ (.B1(\graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ),
    .Y(_2696_),
    .A1(_1507_),
    .A2(net181));
 sg13g2_and3_1 _3539_ (.X(_2697_),
    .A(_2692_),
    .B(_1178_),
    .C(_2696_));
 sg13g2_nor2b_1 _3540_ (.A(net2),
    .B_N(_2697_),
    .Y(_2698_));
 sg13g2_buf_2 _3541_ (.A(_2698_),
    .X(_2699_));
 sg13g2_and2_1 _3542_ (.A(net2),
    .B(_2697_),
    .X(_2700_));
 sg13g2_buf_2 _3543_ (.A(_2700_),
    .X(_2701_));
 sg13g2_buf_1 _3544_ (.A(_2693_),
    .X(_2702_));
 sg13g2_or2_1 _3545_ (.X(_2703_),
    .B(net206),
    .A(net207));
 sg13g2_buf_1 _3546_ (.A(_2703_),
    .X(_2704_));
 sg13g2_nor3_2 _3547_ (.A(_1375_),
    .B(_1463_),
    .C(net158),
    .Y(_2705_));
 sg13g2_xnor2_1 _3548_ (.Y(_2706_),
    .A(net204),
    .B(_2705_));
 sg13g2_buf_2 _3549_ (.A(_0020_),
    .X(_2707_));
 sg13g2_nor4_2 _3550_ (.A(net207),
    .B(net206),
    .C(net219),
    .Y(_2708_),
    .D(net190));
 sg13g2_xor2_1 _3551_ (.B(_2708_),
    .A(_2707_),
    .X(_2709_));
 sg13g2_buf_2 _3552_ (.A(_2709_),
    .X(_2710_));
 sg13g2_buf_1 _3553_ (.A(_0019_),
    .X(_2711_));
 sg13g2_inv_1 _3554_ (.Y(_2712_),
    .A(_2711_));
 sg13g2_and2_1 _3555_ (.A(_2567_),
    .B(_2570_),
    .X(_2713_));
 sg13g2_buf_2 _3556_ (.A(_2713_),
    .X(_2714_));
 sg13g2_nor2_1 _3557_ (.A(net184),
    .B(net183),
    .Y(_2715_));
 sg13g2_buf_2 _3558_ (.A(_2715_),
    .X(_2716_));
 sg13g2_nand2b_1 _3559_ (.Y(_2717_),
    .B(net167),
    .A_N(_2711_));
 sg13g2_buf_1 _3560_ (.A(_0024_),
    .X(_2718_));
 sg13g2_inv_1 _3561_ (.Y(_2719_),
    .A(net228));
 sg13g2_a221oi_1 _3562_ (.B2(_2717_),
    .C1(net203),
    .B1(_2716_),
    .A1(_2712_),
    .Y(_2720_),
    .A2(_2714_));
 sg13g2_buf_1 _3563_ (.A(net167),
    .X(_2721_));
 sg13g2_nor4_1 _3564_ (.A(_2721_),
    .B(_2711_),
    .C(net228),
    .D(net158),
    .Y(_2722_));
 sg13g2_nor3_2 _3565_ (.A(_2710_),
    .B(_2720_),
    .C(_2722_),
    .Y(_2723_));
 sg13g2_xnor2_1 _3566_ (.Y(_2724_),
    .A(_2706_),
    .B(_2723_));
 sg13g2_inv_2 _3567_ (.Y(_2725_),
    .A(net224));
 sg13g2_nor4_1 _3568_ (.A(_1310_),
    .B(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[0] ),
    .C(_1233_),
    .D(_1101_),
    .Y(_2726_));
 sg13g2_buf_2 _3569_ (.A(_2726_),
    .X(_2727_));
 sg13g2_buf_2 _3570_ (.A(_0013_),
    .X(_2728_));
 sg13g2_buf_2 _3571_ (.A(_0030_),
    .X(_2729_));
 sg13g2_nand2b_1 _3572_ (.Y(_2730_),
    .B(_2729_),
    .A_N(_2728_));
 sg13g2_a21o_1 _3573_ (.A2(_2727_),
    .A1(net180),
    .B1(_2730_),
    .X(_2731_));
 sg13g2_buf_1 _3574_ (.A(_2731_),
    .X(_2732_));
 sg13g2_or4_1 _3575_ (.A(_1310_),
    .B(net243),
    .C(_1233_),
    .D(net225),
    .X(_2733_));
 sg13g2_buf_1 _3576_ (.A(_2733_),
    .X(_2734_));
 sg13g2_xnor2_1 _3577_ (.Y(_2735_),
    .A(net245),
    .B(_2728_));
 sg13g2_or4_1 _3578_ (.A(_1145_),
    .B(_2729_),
    .C(_2734_),
    .D(_2735_),
    .X(_2736_));
 sg13g2_buf_1 _3579_ (.A(_2736_),
    .X(_2737_));
 sg13g2_nand2_1 _3580_ (.Y(_2738_),
    .A(net136),
    .B(net116));
 sg13g2_or3_1 _3581_ (.A(_1321_),
    .B(_1189_),
    .C(_1244_),
    .X(_2739_));
 sg13g2_buf_1 _3582_ (.A(_2739_),
    .X(_2740_));
 sg13g2_buf_1 _3583_ (.A(_0029_),
    .X(_2741_));
 sg13g2_buf_1 _3584_ (.A(_2741_),
    .X(_2742_));
 sg13g2_buf_1 _3585_ (.A(net202),
    .X(_2743_));
 sg13g2_buf_1 _3586_ (.A(_0023_),
    .X(_2744_));
 sg13g2_nor2_1 _3587_ (.A(net179),
    .B(net227),
    .Y(_2745_));
 sg13g2_nand2_2 _3588_ (.Y(_2746_),
    .A(_2740_),
    .B(_2745_));
 sg13g2_nor3_2 _3589_ (.A(net221),
    .B(net243),
    .C(net222),
    .Y(_2747_));
 sg13g2_xor2_1 _3590_ (.B(net202),
    .A(net225),
    .X(_2748_));
 sg13g2_nand3_1 _3591_ (.B(_2747_),
    .C(_2748_),
    .A(net227),
    .Y(_2749_));
 sg13g2_buf_2 _3592_ (.A(_2749_),
    .X(_2750_));
 sg13g2_nand2_2 _3593_ (.Y(_2751_),
    .A(_2746_),
    .B(_2750_));
 sg13g2_nand2_1 _3594_ (.Y(_2752_),
    .A(_2738_),
    .B(_2751_));
 sg13g2_or2_1 _3595_ (.X(_2753_),
    .B(net243),
    .A(net221));
 sg13g2_buf_1 _3596_ (.A(_2753_),
    .X(_2754_));
 sg13g2_nor2_1 _3597_ (.A(_1266_),
    .B(_2754_),
    .Y(_2755_));
 sg13g2_nor2b_2 _3598_ (.A(net202),
    .B_N(net227),
    .Y(_2756_));
 sg13g2_nor2b_1 _3599_ (.A(net227),
    .B_N(net202),
    .Y(_2757_));
 sg13g2_buf_1 _3600_ (.A(_0028_),
    .X(_2758_));
 sg13g2_mux2_1 _3601_ (.A0(_2756_),
    .A1(_2757_),
    .S(net226),
    .X(_2759_));
 sg13g2_nand2b_2 _3602_ (.Y(_2760_),
    .B(net194),
    .A_N(net192));
 sg13g2_nor2_1 _3603_ (.A(_2754_),
    .B(_2760_),
    .Y(_2761_));
 sg13g2_or2_1 _3604_ (.X(_2762_),
    .B(net227),
    .A(_2741_));
 sg13g2_buf_1 _3605_ (.A(_2762_),
    .X(_2763_));
 sg13g2_nand3_1 _3606_ (.B(_2742_),
    .C(net227),
    .A(net226),
    .Y(_2764_));
 sg13g2_o21ai_1 _3607_ (.B1(_2764_),
    .Y(_2765_),
    .A1(net226),
    .A2(_2763_));
 sg13g2_a22oi_1 _3608_ (.Y(_2766_),
    .B1(_2761_),
    .B2(_2765_),
    .A2(_2759_),
    .A1(_2755_));
 sg13g2_buf_1 _3609_ (.A(_2766_),
    .X(_2767_));
 sg13g2_nor2_2 _3610_ (.A(net192),
    .B(net194),
    .Y(_2768_));
 sg13g2_inv_2 _3611_ (.Y(_2769_),
    .A(net226));
 sg13g2_mux2_1 _3612_ (.A0(_2756_),
    .A1(_2757_),
    .S(_2769_),
    .X(_2770_));
 sg13g2_o21ai_1 _3613_ (.B1(_2770_),
    .Y(_2771_),
    .A1(_2768_),
    .A2(_2754_));
 sg13g2_buf_1 _3614_ (.A(_2771_),
    .X(_2772_));
 sg13g2_a221oi_1 _3615_ (.B2(_2772_),
    .C1(_2556_),
    .B1(_2767_),
    .A1(net136),
    .Y(_2773_),
    .A2(net116));
 sg13g2_buf_1 _3616_ (.A(net226),
    .X(_2774_));
 sg13g2_buf_1 _3617_ (.A(net201),
    .X(_2775_));
 sg13g2_a21oi_2 _3618_ (.B1(_2730_),
    .Y(_2776_),
    .A2(_2727_),
    .A1(net180));
 sg13g2_buf_1 _3619_ (.A(_2729_),
    .X(_2777_));
 sg13g2_nor4_2 _3620_ (.A(net224),
    .B(net200),
    .C(_2734_),
    .Y(_2778_),
    .D(_2735_));
 sg13g2_nor2_2 _3621_ (.A(_2776_),
    .B(_2778_),
    .Y(_2779_));
 sg13g2_nor2_1 _3622_ (.A(net221),
    .B(net243),
    .Y(_2780_));
 sg13g2_xnor2_1 _3623_ (.Y(_2781_),
    .A(net226),
    .B(net227));
 sg13g2_a21o_1 _3624_ (.A2(_2780_),
    .A1(_2604_),
    .B1(_2781_),
    .X(_2782_));
 sg13g2_buf_1 _3625_ (.A(_2780_),
    .X(_2783_));
 sg13g2_nand3_1 _3626_ (.B(net157),
    .C(_2781_),
    .A(_2604_),
    .Y(_2784_));
 sg13g2_inv_1 _3627_ (.Y(_2785_),
    .A(net202));
 sg13g2_xnor2_1 _3628_ (.Y(_2786_),
    .A(net177),
    .B(_2727_));
 sg13g2_a21o_1 _3629_ (.A2(_2784_),
    .A1(_2782_),
    .B1(_2786_),
    .X(_2787_));
 sg13g2_nor4_1 _3630_ (.A(_1332_),
    .B(net178),
    .C(_2779_),
    .D(_2787_),
    .Y(_2788_));
 sg13g2_o21ai_1 _3631_ (.B1(net157),
    .Y(_2789_),
    .A1(_2776_),
    .A2(_2778_));
 sg13g2_o21ai_1 _3632_ (.B1(net178),
    .Y(_2790_),
    .A1(_2776_),
    .A2(_2778_));
 sg13g2_a22oi_1 _3633_ (.Y(_2791_),
    .B1(_2789_),
    .B2(_2790_),
    .A2(_2772_),
    .A1(_2767_));
 sg13g2_nor2b_1 _3634_ (.A(_2758_),
    .B_N(net223),
    .Y(_2792_));
 sg13g2_buf_1 _3635_ (.A(_2792_),
    .X(_2793_));
 sg13g2_inv_1 _3636_ (.Y(_2794_),
    .A(_2793_));
 sg13g2_nand2_1 _3637_ (.Y(_2795_),
    .A(net201),
    .B(net157));
 sg13g2_a221oi_1 _3638_ (.B2(_2795_),
    .C1(_2787_),
    .B1(_2794_),
    .A1(net136),
    .Y(_2796_),
    .A2(net116));
 sg13g2_nor4_2 _3639_ (.A(_2773_),
    .B(_2788_),
    .C(_2791_),
    .Y(_2797_),
    .D(_2796_));
 sg13g2_buf_1 _3640_ (.A(net227),
    .X(_2798_));
 sg13g2_nor2b_1 _3641_ (.A(net199),
    .B_N(_1200_),
    .Y(_2799_));
 sg13g2_xnor2_1 _3642_ (.Y(_2800_),
    .A(_1200_),
    .B(net199));
 sg13g2_mux2_1 _3643_ (.A0(_2799_),
    .A1(_2800_),
    .S(_1321_),
    .X(_2801_));
 sg13g2_xor2_1 _3644_ (.B(net199),
    .A(net164),
    .X(_2802_));
 sg13g2_nor3_1 _3645_ (.A(net201),
    .B(_2754_),
    .C(_2802_),
    .Y(_2803_));
 sg13g2_a21o_1 _3646_ (.A2(_2801_),
    .A1(net178),
    .B1(_2803_),
    .X(_2804_));
 sg13g2_buf_1 _3647_ (.A(_2804_),
    .X(_2805_));
 sg13g2_a21oi_2 _3648_ (.B1(_2786_),
    .Y(_2806_),
    .A2(_2737_),
    .A1(_2732_));
 sg13g2_nand2_2 _3649_ (.Y(_2807_),
    .A(_2805_),
    .B(_2806_));
 sg13g2_or2_1 _3650_ (.X(_2808_),
    .B(_2722_),
    .A(_2720_));
 sg13g2_buf_2 _3651_ (.A(_2808_),
    .X(_2809_));
 sg13g2_buf_1 _3652_ (.A(_2711_),
    .X(_2810_));
 sg13g2_nor2_2 _3653_ (.A(net198),
    .B(_2574_),
    .Y(_2811_));
 sg13g2_nor3_2 _3654_ (.A(net207),
    .B(net183),
    .C(net190),
    .Y(_2812_));
 sg13g2_xnor2_1 _3655_ (.Y(_2813_),
    .A(net228),
    .B(_2812_));
 sg13g2_buf_2 _3656_ (.A(_2813_),
    .X(_2814_));
 sg13g2_buf_1 _3657_ (.A(_2712_),
    .X(_2815_));
 sg13g2_xnor2_1 _3658_ (.Y(_2816_),
    .A(net167),
    .B(net228));
 sg13g2_nor3_1 _3659_ (.A(net176),
    .B(net158),
    .C(_2816_),
    .Y(_2817_));
 sg13g2_a21o_1 _3660_ (.A2(_2814_),
    .A1(_2811_),
    .B1(_2817_),
    .X(_2818_));
 sg13g2_buf_2 _3661_ (.A(_2818_),
    .X(_2819_));
 sg13g2_xnor2_1 _3662_ (.Y(_2820_),
    .A(_2707_),
    .B(_2708_));
 sg13g2_mux2_1 _3663_ (.A0(_2809_),
    .A1(_2819_),
    .S(_2820_),
    .X(_2821_));
 sg13g2_nand2_1 _3664_ (.Y(_2822_),
    .A(_2574_),
    .B(net158));
 sg13g2_buf_1 _3665_ (.A(_2822_),
    .X(_2823_));
 sg13g2_buf_1 _3666_ (.A(net101),
    .X(_2824_));
 sg13g2_nand3_1 _3667_ (.B(_2821_),
    .C(_2824_),
    .A(_2807_),
    .Y(_2825_));
 sg13g2_a21oi_1 _3668_ (.A1(_2752_),
    .A2(_2797_),
    .Y(_2826_),
    .B1(_2825_));
 sg13g2_nand2_1 _3669_ (.Y(_2827_),
    .A(net176),
    .B(_2714_));
 sg13g2_nand2_1 _3670_ (.Y(_2828_),
    .A(net198),
    .B(_2716_));
 sg13g2_and2_1 _3671_ (.A(_2827_),
    .B(_2828_),
    .X(_2829_));
 sg13g2_xor2_1 _3672_ (.B(net243),
    .A(net221),
    .X(_2830_));
 sg13g2_buf_2 _3673_ (.A(_2830_),
    .X(_2831_));
 sg13g2_nand2_1 _3674_ (.Y(_2832_),
    .A(net201),
    .B(_2831_));
 sg13g2_buf_2 _3675_ (.A(_2832_),
    .X(_2833_));
 sg13g2_a21oi_2 _3676_ (.B1(_2833_),
    .Y(_2834_),
    .A2(_2750_),
    .A1(_2746_));
 sg13g2_nand2_1 _3677_ (.Y(_2835_),
    .A(_2767_),
    .B(_2772_));
 sg13g2_buf_1 _3678_ (.A(net198),
    .X(_2836_));
 sg13g2_and2_1 _3679_ (.A(net201),
    .B(_2831_),
    .X(_2837_));
 sg13g2_buf_1 _3680_ (.A(_2837_),
    .X(_2838_));
 sg13g2_nor2b_2 _3681_ (.A(net193),
    .B_N(_2758_),
    .Y(_2839_));
 sg13g2_mux2_1 _3682_ (.A0(_2793_),
    .A1(_2839_),
    .S(_1332_),
    .X(_2840_));
 sg13g2_buf_2 _3683_ (.A(_2840_),
    .X(_2841_));
 sg13g2_nor2_1 _3684_ (.A(_2838_),
    .B(_2841_),
    .Y(_2842_));
 sg13g2_nor4_1 _3685_ (.A(net175),
    .B(_2779_),
    .C(net101),
    .D(_2842_),
    .Y(_2843_));
 sg13g2_o21ai_1 _3686_ (.B1(_2843_),
    .Y(_2844_),
    .A1(_2834_),
    .A2(_2835_));
 sg13g2_nor2b_1 _3687_ (.A(_2787_),
    .B_N(_2841_),
    .Y(_2845_));
 sg13g2_nor2_1 _3688_ (.A(net176),
    .B(_2714_),
    .Y(_2846_));
 sg13g2_nor2_2 _3689_ (.A(_2811_),
    .B(_2846_),
    .Y(_2847_));
 sg13g2_inv_1 _3690_ (.Y(_2848_),
    .A(_2831_));
 sg13g2_nor2_1 _3691_ (.A(net201),
    .B(_2848_),
    .Y(_2849_));
 sg13g2_buf_2 _3692_ (.A(_2849_),
    .X(_2850_));
 sg13g2_nor3_1 _3693_ (.A(_2779_),
    .B(_2847_),
    .C(_2850_),
    .Y(_2851_));
 sg13g2_o21ai_1 _3694_ (.B1(_2851_),
    .Y(_2852_),
    .A1(_2835_),
    .A2(_2845_));
 sg13g2_and4_1 _3695_ (.A(_2821_),
    .B(_2829_),
    .C(_2844_),
    .D(_2852_),
    .X(_2853_));
 sg13g2_nor3_1 _3696_ (.A(_2724_),
    .B(_2826_),
    .C(_2853_),
    .Y(_2854_));
 sg13g2_buf_2 _3697_ (.A(_0017_),
    .X(_2855_));
 sg13g2_nor2b_2 _3698_ (.A(net240),
    .B_N(_2705_),
    .Y(_2856_));
 sg13g2_xnor2_1 _3699_ (.Y(_2857_),
    .A(_2855_),
    .B(_2856_));
 sg13g2_buf_2 _3700_ (.A(_2857_),
    .X(_2858_));
 sg13g2_nor2_1 _3701_ (.A(_2706_),
    .B(_2723_),
    .Y(_2859_));
 sg13g2_xnor2_1 _3702_ (.Y(_2860_),
    .A(_2858_),
    .B(_2859_));
 sg13g2_nand2b_1 _3703_ (.Y(_2861_),
    .B(_2860_),
    .A_N(_2854_));
 sg13g2_nor2_1 _3704_ (.A(_2714_),
    .B(_2716_),
    .Y(_2862_));
 sg13g2_buf_2 _3705_ (.A(_2862_),
    .X(_2863_));
 sg13g2_buf_1 _3706_ (.A(_2863_),
    .X(_2864_));
 sg13g2_buf_1 _3707_ (.A(net85),
    .X(_2865_));
 sg13g2_a221oi_1 _3708_ (.B2(_2784_),
    .C1(_2786_),
    .B1(_2782_),
    .A1(net136),
    .Y(_2866_),
    .A2(net116));
 sg13g2_buf_1 _3709_ (.A(_2866_),
    .X(_2867_));
 sg13g2_a21oi_1 _3710_ (.A1(_2767_),
    .A2(_2772_),
    .Y(_2868_),
    .B1(_2779_));
 sg13g2_o21ai_1 _3711_ (.B1(_2841_),
    .Y(_2869_),
    .A1(_2867_),
    .A2(_2868_));
 sg13g2_xnor2_1 _3712_ (.Y(_2870_),
    .A(_2769_),
    .B(net157));
 sg13g2_a221oi_1 _3713_ (.B2(_2870_),
    .C1(net85),
    .B1(_2868_),
    .A1(_2850_),
    .Y(_2871_),
    .A2(_2867_));
 sg13g2_a21oi_1 _3714_ (.A1(net66),
    .A2(_2869_),
    .Y(_2872_),
    .B1(_2871_));
 sg13g2_nor2_1 _3715_ (.A(_2847_),
    .B(_2872_),
    .Y(_2873_));
 sg13g2_nand2_1 _3716_ (.Y(_2874_),
    .A(net175),
    .B(_2574_));
 sg13g2_nand2_2 _3717_ (.Y(_2875_),
    .A(_2827_),
    .B(_2874_));
 sg13g2_and2_1 _3718_ (.A(_2752_),
    .B(_2797_),
    .X(_2876_));
 sg13g2_buf_1 _3719_ (.A(_2876_),
    .X(_2877_));
 sg13g2_o21ai_1 _3720_ (.B1(_2738_),
    .Y(_2878_),
    .A1(_2751_),
    .A2(_2835_));
 sg13g2_nand2_1 _3721_ (.Y(_2879_),
    .A(net85),
    .B(_2838_));
 sg13g2_nand3_1 _3722_ (.B(_2850_),
    .C(_2867_),
    .A(net85),
    .Y(_2880_));
 sg13g2_o21ai_1 _3723_ (.B1(_2880_),
    .Y(_2881_),
    .A1(_2878_),
    .A2(_2879_));
 sg13g2_nor2_1 _3724_ (.A(_2807_),
    .B(_2863_),
    .Y(_2882_));
 sg13g2_nor4_1 _3725_ (.A(_2875_),
    .B(_2877_),
    .C(_2881_),
    .D(_2882_),
    .Y(_2883_));
 sg13g2_nor4_1 _3726_ (.A(_2710_),
    .B(_2809_),
    .C(_2819_),
    .D(_2858_),
    .Y(_2884_));
 sg13g2_o21ai_1 _3727_ (.B1(_2884_),
    .Y(_2885_),
    .A1(_2873_),
    .A2(_2883_));
 sg13g2_nor4_1 _3728_ (.A(net221),
    .B(_1189_),
    .C(net192),
    .D(_2744_),
    .Y(_2886_));
 sg13g2_a22oi_1 _3729_ (.Y(_2887_),
    .B1(_2748_),
    .B2(_2886_),
    .A2(_2756_),
    .A1(_2740_));
 sg13g2_buf_1 _3730_ (.A(_2887_),
    .X(_2888_));
 sg13g2_or3_1 _3731_ (.A(_2779_),
    .B(_2870_),
    .C(_2888_),
    .X(_2889_));
 sg13g2_buf_1 _3732_ (.A(_2889_),
    .X(_2890_));
 sg13g2_nor2_1 _3733_ (.A(_2890_),
    .B(_2824_),
    .Y(_2891_));
 sg13g2_or3_1 _3734_ (.A(_2847_),
    .B(_2882_),
    .C(_2891_),
    .X(_2892_));
 sg13g2_nand2_1 _3735_ (.Y(_2893_),
    .A(_2740_),
    .B(_2756_));
 sg13g2_nand2_1 _3736_ (.Y(_2894_),
    .A(_2748_),
    .B(_2886_));
 sg13g2_a221oi_1 _3737_ (.B2(_2894_),
    .C1(_2870_),
    .B1(_2893_),
    .A1(_2732_),
    .Y(_2895_),
    .A2(_2737_));
 sg13g2_or2_1 _3738_ (.X(_2896_),
    .B(_2895_),
    .A(net175));
 sg13g2_buf_1 _3739_ (.A(net137),
    .X(_2897_));
 sg13g2_buf_1 _3740_ (.A(_2897_),
    .X(_2898_));
 sg13g2_nor2_1 _3741_ (.A(net160),
    .B(net100),
    .Y(_2899_));
 sg13g2_buf_1 _3742_ (.A(net175),
    .X(_2900_));
 sg13g2_a22oi_1 _3743_ (.Y(_2901_),
    .B1(_2899_),
    .B2(net156),
    .A2(net85),
    .A1(_2896_));
 sg13g2_buf_1 _3744_ (.A(net115),
    .X(_2902_));
 sg13g2_nand2_1 _3745_ (.Y(_2903_),
    .A(net99),
    .B(net175));
 sg13g2_nor2_1 _3746_ (.A(net158),
    .B(_2903_),
    .Y(_2904_));
 sg13g2_nor3_1 _3747_ (.A(net203),
    .B(_2811_),
    .C(_2904_),
    .Y(_2905_));
 sg13g2_a21oi_1 _3748_ (.A1(net203),
    .A2(_2901_),
    .Y(_2906_),
    .B1(_2905_));
 sg13g2_o21ai_1 _3749_ (.B1(_2906_),
    .Y(_2907_),
    .A1(_2877_),
    .A2(_2892_));
 sg13g2_nor2_1 _3750_ (.A(net161),
    .B(_2836_),
    .Y(_2908_));
 sg13g2_inv_1 _3751_ (.Y(_2909_),
    .A(_2908_));
 sg13g2_a221oi_1 _3752_ (.B2(_2750_),
    .C1(_2833_),
    .B1(_2746_),
    .A1(net136),
    .Y(_2910_),
    .A2(net116));
 sg13g2_buf_1 _3753_ (.A(_2910_),
    .X(_2911_));
 sg13g2_buf_1 _3754_ (.A(_2572_),
    .X(_2912_));
 sg13g2_buf_1 _3755_ (.A(net155),
    .X(_2913_));
 sg13g2_buf_1 _3756_ (.A(net135),
    .X(_2914_));
 sg13g2_nor2_1 _3757_ (.A(net114),
    .B(net176),
    .Y(_2915_));
 sg13g2_a21oi_1 _3758_ (.A1(_2909_),
    .A2(_2911_),
    .Y(_2916_),
    .B1(_2915_));
 sg13g2_nor3_1 _3759_ (.A(_2665_),
    .B(net203),
    .C(_2916_),
    .Y(_2917_));
 sg13g2_xnor2_1 _3760_ (.Y(_2918_),
    .A(net203),
    .B(_2812_));
 sg13g2_buf_1 _3761_ (.A(_2918_),
    .X(_2919_));
 sg13g2_nor2_1 _3762_ (.A(net184),
    .B(net161),
    .Y(_2920_));
 sg13g2_nand3_1 _3763_ (.B(net113),
    .C(_2920_),
    .A(net156),
    .Y(_2921_));
 sg13g2_buf_1 _3764_ (.A(_2814_),
    .X(_2922_));
 sg13g2_nand4_1 _3765_ (.B(_2806_),
    .C(_2811_),
    .A(_2805_),
    .Y(_2923_),
    .D(net98));
 sg13g2_nand3_1 _3766_ (.B(_2806_),
    .C(_2817_),
    .A(_2805_),
    .Y(_2924_));
 sg13g2_nand4_1 _3767_ (.B(net176),
    .C(net113),
    .A(_2665_),
    .Y(_2925_),
    .D(_2911_));
 sg13g2_nand4_1 _3768_ (.B(_2923_),
    .C(_2924_),
    .A(_2921_),
    .Y(_2926_),
    .D(_2925_));
 sg13g2_nor2_1 _3769_ (.A(_2888_),
    .B(_2838_),
    .Y(_2927_));
 sg13g2_or2_1 _3770_ (.X(_2928_),
    .B(_2834_),
    .A(_2927_));
 sg13g2_nand2_1 _3771_ (.Y(_2929_),
    .A(_2738_),
    .B(_2928_));
 sg13g2_o21ai_1 _3772_ (.B1(net66),
    .Y(_2930_),
    .A1(_2815_),
    .A2(_2929_));
 sg13g2_o21ai_1 _3773_ (.B1(_2930_),
    .Y(_2931_),
    .A1(_2917_),
    .A2(_2926_));
 sg13g2_a22oi_1 _3774_ (.Y(_2932_),
    .B1(_2746_),
    .B2(_2750_),
    .A2(net116),
    .A1(net136));
 sg13g2_buf_1 _3775_ (.A(_2932_),
    .X(_2933_));
 sg13g2_nand2_1 _3776_ (.Y(_2934_),
    .A(_2933_),
    .B(_2850_));
 sg13g2_a22oi_1 _3777_ (.Y(_2935_),
    .B1(_2934_),
    .B2(_2890_),
    .A2(_2929_),
    .A1(_2875_));
 sg13g2_nand4_1 _3778_ (.B(net158),
    .C(_2809_),
    .A(_2574_),
    .Y(_2936_),
    .D(_2935_));
 sg13g2_xnor2_1 _3779_ (.Y(_2937_),
    .A(_2710_),
    .B(_2809_));
 sg13g2_buf_1 _3780_ (.A(_2706_),
    .X(_2938_));
 sg13g2_xnor2_1 _3781_ (.Y(_2939_),
    .A(_2858_),
    .B(_2938_));
 sg13g2_nor2_1 _3782_ (.A(_2937_),
    .B(_2939_),
    .Y(_2940_));
 sg13g2_nand4_1 _3783_ (.B(_2931_),
    .C(_2936_),
    .A(_2907_),
    .Y(_2941_),
    .D(_2940_));
 sg13g2_nand3_1 _3784_ (.B(_2885_),
    .C(_2941_),
    .A(_2861_),
    .Y(_2942_));
 sg13g2_nor2_1 _3785_ (.A(net85),
    .B(_2841_),
    .Y(_2943_));
 sg13g2_a221oi_1 _3786_ (.B2(net201),
    .C1(_2888_),
    .B1(_2831_),
    .A1(net136),
    .Y(_2944_),
    .A2(net116));
 sg13g2_buf_1 _3787_ (.A(_2944_),
    .X(_2945_));
 sg13g2_nor2b_1 _3788_ (.A(_2945_),
    .B_N(_2841_),
    .Y(_2946_));
 sg13g2_a221oi_1 _3789_ (.B2(_2864_),
    .C1(_2752_),
    .B1(_2946_),
    .A1(_2807_),
    .Y(_2947_),
    .A2(_2943_));
 sg13g2_o21ai_1 _3790_ (.B1(_2906_),
    .Y(_2948_),
    .A1(_2847_),
    .A2(_2947_));
 sg13g2_a21o_1 _3791_ (.A2(_2945_),
    .A1(net66),
    .B1(_2882_),
    .X(_2949_));
 sg13g2_nand3b_1 _3792_ (.B(_2906_),
    .C(_2949_),
    .Y(_2950_),
    .A_N(_2797_));
 sg13g2_nand3_1 _3793_ (.B(_2948_),
    .C(_2950_),
    .A(_2931_),
    .Y(_2951_));
 sg13g2_and2_1 _3794_ (.A(_2937_),
    .B(_2724_),
    .X(_2952_));
 sg13g2_nor2_1 _3795_ (.A(net66),
    .B(_2797_),
    .Y(_2953_));
 sg13g2_a21oi_1 _3796_ (.A1(_2846_),
    .A2(_2877_),
    .Y(_2954_),
    .B1(_2953_));
 sg13g2_nand2_1 _3797_ (.Y(_2955_),
    .A(_2833_),
    .B(_2933_));
 sg13g2_nor2_1 _3798_ (.A(_2833_),
    .B(_2874_),
    .Y(_2956_));
 sg13g2_nor2_1 _3799_ (.A(_2809_),
    .B(_2819_),
    .Y(_2957_));
 sg13g2_a221oi_1 _3800_ (.B2(_2933_),
    .C1(_2957_),
    .B1(_2956_),
    .A1(_2811_),
    .Y(_2958_),
    .A2(_2955_));
 sg13g2_buf_1 _3801_ (.A(_2718_),
    .X(_2959_));
 sg13g2_nor2b_1 _3802_ (.A(net198),
    .B_N(net197),
    .Y(_2960_));
 sg13g2_nor2_1 _3803_ (.A(net160),
    .B(net197),
    .Y(_2961_));
 sg13g2_a21oi_1 _3804_ (.A1(net160),
    .A2(_2960_),
    .Y(_2962_),
    .B1(_2961_));
 sg13g2_nand2_1 _3805_ (.Y(_2963_),
    .A(_2769_),
    .B(net157));
 sg13g2_and2_1 _3806_ (.A(net223),
    .B(net226),
    .X(_2964_));
 sg13g2_buf_2 _3807_ (.A(_2964_),
    .X(_2965_));
 sg13g2_nand2_1 _3808_ (.Y(_2966_),
    .A(net186),
    .B(_2965_));
 sg13g2_a221oi_1 _3809_ (.B2(_2966_),
    .C1(_2888_),
    .B1(_2963_),
    .A1(net136),
    .Y(_2967_),
    .A2(net116));
 sg13g2_buf_1 _3810_ (.A(_2967_),
    .X(_2968_));
 sg13g2_nor3_1 _3811_ (.A(net156),
    .B(net113),
    .C(_2968_),
    .Y(_2969_));
 sg13g2_a21o_1 _3812_ (.A2(_2919_),
    .A1(_2915_),
    .B1(net160),
    .X(_2970_));
 sg13g2_nand2_1 _3813_ (.Y(_2971_),
    .A(net156),
    .B(net98));
 sg13g2_a21oi_1 _3814_ (.A1(net139),
    .A2(_2719_),
    .Y(_2972_),
    .B1(_2665_));
 sg13g2_o21ai_1 _3815_ (.B1(_2972_),
    .Y(_2973_),
    .A1(_2968_),
    .A2(_2971_));
 sg13g2_o21ai_1 _3816_ (.B1(_2973_),
    .Y(_2974_),
    .A1(_2969_),
    .A2(_2970_));
 sg13g2_o21ai_1 _3817_ (.B1(_2974_),
    .Y(_2975_),
    .A1(net139),
    .A2(_2962_));
 sg13g2_o21ai_1 _3818_ (.B1(_2880_),
    .Y(_2976_),
    .A1(_2865_),
    .A2(_2929_));
 sg13g2_nand2_1 _3819_ (.Y(_2977_),
    .A(_2875_),
    .B(_2976_));
 sg13g2_nand2b_1 _3820_ (.Y(_2978_),
    .B(_2724_),
    .A_N(_2937_));
 sg13g2_a221oi_1 _3821_ (.B2(_2977_),
    .C1(_2978_),
    .B1(_2975_),
    .A1(_2954_),
    .Y(_2979_),
    .A2(_2958_));
 sg13g2_a21oi_1 _3822_ (.A1(_2951_),
    .A2(_2952_),
    .Y(_2980_),
    .B1(_2979_));
 sg13g2_mux2_1 _3823_ (.A0(_2807_),
    .A1(_2890_),
    .S(net139),
    .X(_2981_));
 sg13g2_nand3_1 _3824_ (.B(_2900_),
    .C(_2981_),
    .A(_2665_),
    .Y(_2982_));
 sg13g2_a22oi_1 _3825_ (.Y(_2983_),
    .B1(_2915_),
    .B2(_2807_),
    .A2(_2908_),
    .A1(_2890_));
 sg13g2_nand2b_1 _3826_ (.Y(_2984_),
    .B(net160),
    .A_N(_2983_));
 sg13g2_nand2_1 _3827_ (.Y(_2985_),
    .A(_2823_),
    .B(_2945_));
 sg13g2_nand2_1 _3828_ (.Y(_2986_),
    .A(_2838_),
    .B(_2933_));
 sg13g2_nand3_1 _3829_ (.B(_2986_),
    .C(_2847_),
    .A(_2985_),
    .Y(_2987_));
 sg13g2_nand4_1 _3830_ (.B(_2984_),
    .C(_2821_),
    .A(_2982_),
    .Y(_2988_),
    .D(_2987_));
 sg13g2_buf_1 _3831_ (.A(_2707_),
    .X(_2989_));
 sg13g2_nor3_1 _3832_ (.A(_2665_),
    .B(_2989_),
    .C(net197),
    .Y(_2990_));
 sg13g2_a21oi_1 _3833_ (.A1(_2665_),
    .A2(net196),
    .Y(_2991_),
    .B1(_2990_));
 sg13g2_and2_1 _3834_ (.A(net184),
    .B(net196),
    .X(_2992_));
 sg13g2_o21ai_1 _3835_ (.B1(_2992_),
    .Y(_2993_),
    .A1(net139),
    .A2(_2959_));
 sg13g2_o21ai_1 _3836_ (.B1(_2993_),
    .Y(_2994_),
    .A1(net139),
    .A2(_2991_));
 sg13g2_buf_1 _3837_ (.A(_2820_),
    .X(_2995_));
 sg13g2_xnor2_1 _3838_ (.Y(_2996_),
    .A(net112),
    .B(_2922_));
 sg13g2_nor3_2 _3839_ (.A(net184),
    .B(net183),
    .C(_2711_),
    .Y(_2997_));
 sg13g2_a22oi_1 _3840_ (.Y(_2998_),
    .B1(_2996_),
    .B2(_2997_),
    .A2(_2994_),
    .A1(net156));
 sg13g2_nor2_1 _3841_ (.A(_2929_),
    .B(_2998_),
    .Y(_2999_));
 sg13g2_nand2_1 _3842_ (.Y(_3000_),
    .A(_2863_),
    .B(_2968_));
 sg13g2_nand3_1 _3843_ (.B(_2850_),
    .C(_2867_),
    .A(_2822_),
    .Y(_3001_));
 sg13g2_a21o_1 _3844_ (.A2(_3001_),
    .A1(_3000_),
    .B1(net112),
    .X(_3002_));
 sg13g2_or2_1 _3845_ (.X(_3003_),
    .B(_2968_),
    .A(_2823_));
 sg13g2_nand3_1 _3846_ (.B(_2833_),
    .C(_2933_),
    .A(net101),
    .Y(_3004_));
 sg13g2_nand4_1 _3847_ (.B(_3003_),
    .C(_3004_),
    .A(_2875_),
    .Y(_3005_),
    .D(_2937_));
 sg13g2_o21ai_1 _3848_ (.B1(_3005_),
    .Y(_3006_),
    .A1(_2875_),
    .A2(_3002_));
 sg13g2_o21ai_1 _3849_ (.B1(_2957_),
    .Y(_3007_),
    .A1(_2999_),
    .A2(_3006_));
 sg13g2_inv_1 _3850_ (.Y(_3008_),
    .A(_2860_));
 sg13g2_nand4_1 _3851_ (.B(_3007_),
    .C(_2724_),
    .A(_2988_),
    .Y(_3009_),
    .D(_3008_));
 sg13g2_xor2_1 _3852_ (.B(_2856_),
    .A(_2855_),
    .X(_3010_));
 sg13g2_buf_2 _3853_ (.A(_0016_),
    .X(_3011_));
 sg13g2_nand2_1 _3854_ (.Y(_3012_),
    .A(_1518_),
    .B(_2856_));
 sg13g2_xor2_1 _3855_ (.B(_3012_),
    .A(_3011_),
    .X(_3013_));
 sg13g2_nor2b_1 _3856_ (.A(_3013_),
    .B_N(_2859_),
    .Y(_3014_));
 sg13g2_xnor2_1 _3857_ (.Y(_3015_),
    .A(net181),
    .B(_2705_));
 sg13g2_nand2_1 _3858_ (.Y(_3016_),
    .A(_2710_),
    .B(_3015_));
 sg13g2_or3_1 _3859_ (.A(_2819_),
    .B(_2858_),
    .C(_3016_),
    .X(_3017_));
 sg13g2_a22oi_1 _3860_ (.Y(_3018_),
    .B1(_3017_),
    .B2(_3013_),
    .A2(_3014_),
    .A1(_3010_));
 sg13g2_a21oi_1 _3861_ (.A1(_2890_),
    .A2(_2878_),
    .Y(_3019_),
    .B1(net5));
 sg13g2_nand2_1 _3862_ (.Y(_3020_),
    .A(net156),
    .B(net66));
 sg13g2_a21oi_1 _3863_ (.A1(_2752_),
    .A2(_2797_),
    .Y(_3021_),
    .B1(_2968_));
 sg13g2_a21o_1 _3864_ (.A2(_2797_),
    .A1(_2986_),
    .B1(net66),
    .X(_3022_));
 sg13g2_o21ai_1 _3865_ (.B1(_3022_),
    .Y(_3023_),
    .A1(_3020_),
    .A2(_3021_));
 sg13g2_nor3_1 _3866_ (.A(net112),
    .B(_2809_),
    .C(_2819_),
    .Y(_3024_));
 sg13g2_nand2_1 _3867_ (.Y(_3025_),
    .A(_2716_),
    .B(_2945_));
 sg13g2_mux2_1 _3868_ (.A0(_2945_),
    .A1(_2911_),
    .S(_2668_),
    .X(_3026_));
 sg13g2_a22oi_1 _3869_ (.Y(_3027_),
    .B1(_3026_),
    .B2(net160),
    .A2(_2911_),
    .A1(_2920_));
 sg13g2_mux4_1 _3870_ (.S0(_2900_),
    .A0(_2574_),
    .A1(_2704_),
    .A2(_3025_),
    .A3(_3027_),
    .S1(_2919_),
    .X(_3028_));
 sg13g2_nor3_1 _3871_ (.A(_2995_),
    .B(_3010_),
    .C(_3015_),
    .Y(_3029_));
 sg13g2_nand2_1 _3872_ (.Y(_3030_),
    .A(_2957_),
    .B(_3001_));
 sg13g2_nand2_1 _3873_ (.Y(_3031_),
    .A(_2895_),
    .B(_2908_));
 sg13g2_o21ai_1 _3874_ (.B1(_3031_),
    .Y(_3032_),
    .A1(_2815_),
    .A2(_2807_));
 sg13g2_and2_1 _3875_ (.A(net155),
    .B(_2711_),
    .X(_3033_));
 sg13g2_buf_1 _3876_ (.A(_3033_),
    .X(_3034_));
 sg13g2_nand3_1 _3877_ (.B(_2806_),
    .C(_3034_),
    .A(_2805_),
    .Y(_3035_));
 sg13g2_nand3_1 _3878_ (.B(_2895_),
    .C(_2716_),
    .A(net175),
    .Y(_3036_));
 sg13g2_nand3_1 _3879_ (.B(_2806_),
    .C(_2997_),
    .A(_2805_),
    .Y(_3037_));
 sg13g2_nand3_1 _3880_ (.B(_3036_),
    .C(_3037_),
    .A(_3035_),
    .Y(_3038_));
 sg13g2_a221oi_1 _3881_ (.B2(net160),
    .C1(_3038_),
    .B1(_3032_),
    .A1(_2937_),
    .Y(_3039_),
    .A2(_3030_));
 sg13g2_buf_1 _3882_ (.A(_2855_),
    .X(_3040_));
 sg13g2_nand2_1 _3883_ (.Y(_3041_),
    .A(_2580_),
    .B(_2705_));
 sg13g2_xnor2_1 _3884_ (.Y(_3042_),
    .A(net181),
    .B(_2723_));
 sg13g2_mux2_1 _3885_ (.A0(_2705_),
    .A1(_3041_),
    .S(_3042_),
    .X(_3043_));
 sg13g2_nand3_1 _3886_ (.B(_2856_),
    .C(_3042_),
    .A(_3040_),
    .Y(_3044_));
 sg13g2_o21ai_1 _3887_ (.B1(_3044_),
    .Y(_3045_),
    .A1(_3040_),
    .A2(_3043_));
 sg13g2_nand3_1 _3888_ (.B(_2819_),
    .C(_2985_),
    .A(_2995_),
    .Y(_3046_));
 sg13g2_nor3_1 _3889_ (.A(_3010_),
    .B(_2938_),
    .C(_3046_),
    .Y(_3047_));
 sg13g2_a221oi_1 _3890_ (.B2(_3045_),
    .C1(_3047_),
    .B1(_3039_),
    .A1(_3028_),
    .Y(_3048_),
    .A2(_3029_));
 sg13g2_a21o_1 _3891_ (.A2(_3024_),
    .A1(_3023_),
    .B1(_3048_),
    .X(_3049_));
 sg13g2_nand4_1 _3892_ (.B(_3018_),
    .C(_3019_),
    .A(_3009_),
    .Y(_3050_),
    .D(_3049_));
 sg13g2_a21o_1 _3893_ (.A2(_2980_),
    .A1(_2942_),
    .B1(_3050_),
    .X(_0108_));
 sg13g2_xnor2_1 _3894_ (.Y(_0109_),
    .A(net198),
    .B(_2716_));
 sg13g2_nand2_1 _3895_ (.Y(_0110_),
    .A(_2814_),
    .B(_0109_));
 sg13g2_nor2_2 _3896_ (.A(_2710_),
    .B(_0110_),
    .Y(_0111_));
 sg13g2_nand2_1 _3897_ (.Y(_0112_),
    .A(net84),
    .B(_0111_));
 sg13g2_a21oi_1 _3898_ (.A1(net184),
    .A2(_3034_),
    .Y(_0113_),
    .B1(_2997_));
 sg13g2_inv_1 _3899_ (.Y(_0114_),
    .A(_0113_));
 sg13g2_nand2b_1 _3900_ (.Y(_0115_),
    .B(_2728_),
    .A_N(_2729_));
 sg13g2_buf_1 _3901_ (.A(net200),
    .X(_0116_));
 sg13g2_nand2_1 _3902_ (.Y(_0117_),
    .A(net174),
    .B(_2735_));
 sg13g2_or2_1 _3903_ (.X(_0118_),
    .B(_2735_),
    .A(net174));
 sg13g2_nor2_1 _3904_ (.A(net140),
    .B(_2734_),
    .Y(_0119_));
 sg13g2_buf_1 _3905_ (.A(_2743_),
    .X(_0120_));
 sg13g2_nand2b_1 _3906_ (.Y(_0121_),
    .B(_2774_),
    .A_N(_1211_));
 sg13g2_a22oi_1 _3907_ (.Y(_0122_),
    .B1(_0121_),
    .B2(net221),
    .A2(_2783_),
    .A1(_2558_));
 sg13g2_nor2_1 _3908_ (.A(net179),
    .B(_2793_),
    .Y(_0123_));
 sg13g2_a22oi_1 _3909_ (.Y(_0124_),
    .B1(_0122_),
    .B2(_0123_),
    .A2(_2734_),
    .A1(net154));
 sg13g2_nor2_1 _3910_ (.A(_2751_),
    .B(_0124_),
    .Y(_0125_));
 sg13g2_mux4_1 _3911_ (.S0(_0119_),
    .A0(_0115_),
    .A1(_0117_),
    .A2(_2730_),
    .A3(_0118_),
    .S1(_0125_),
    .X(_0126_));
 sg13g2_buf_1 _3912_ (.A(_0126_),
    .X(_0127_));
 sg13g2_nand2_1 _3913_ (.Y(_0128_),
    .A(_2963_),
    .B(_2966_));
 sg13g2_and2_1 _3914_ (.A(_2751_),
    .B(_0128_),
    .X(_0129_));
 sg13g2_buf_1 _3915_ (.A(_0129_),
    .X(_0130_));
 sg13g2_nor2_1 _3916_ (.A(_2834_),
    .B(_0130_),
    .Y(_0131_));
 sg13g2_nand4_1 _3917_ (.B(net200),
    .C(_2727_),
    .A(net180),
    .Y(_0132_),
    .D(_2735_));
 sg13g2_buf_1 _3918_ (.A(_0132_),
    .X(_0133_));
 sg13g2_a21o_1 _3919_ (.A2(_2727_),
    .A1(net180),
    .B1(_0115_),
    .X(_0134_));
 sg13g2_buf_1 _3920_ (.A(_0134_),
    .X(_0135_));
 sg13g2_nand2_2 _3921_ (.Y(_0136_),
    .A(_0133_),
    .B(_0135_));
 sg13g2_nand3_1 _3922_ (.B(_2850_),
    .C(_0136_),
    .A(_2751_),
    .Y(_0137_));
 sg13g2_buf_2 _3923_ (.A(_0137_),
    .X(_0138_));
 sg13g2_o21ai_1 _3924_ (.B1(_0138_),
    .Y(_0139_),
    .A1(net65),
    .A2(_0131_));
 sg13g2_xnor2_1 _3925_ (.Y(_0140_),
    .A(_2712_),
    .B(_2716_));
 sg13g2_nor2_1 _3926_ (.A(net113),
    .B(_0140_),
    .Y(_0141_));
 sg13g2_buf_1 _3927_ (.A(_0141_),
    .X(_0142_));
 sg13g2_or2_1 _3928_ (.X(_0143_),
    .B(net154),
    .A(net178));
 sg13g2_o21ai_1 _3929_ (.B1(net179),
    .Y(_0144_),
    .A1(_1244_),
    .A2(net225));
 sg13g2_buf_1 _3930_ (.A(_0144_),
    .X(_0145_));
 sg13g2_or3_1 _3931_ (.A(_2605_),
    .B(net163),
    .C(net179),
    .X(_0146_));
 sg13g2_nand4_1 _3932_ (.B(net157),
    .C(_0145_),
    .A(_2775_),
    .Y(_0147_),
    .D(_0146_));
 sg13g2_o21ai_1 _3933_ (.B1(_0147_),
    .Y(_0148_),
    .A1(_2556_),
    .A2(_0143_));
 sg13g2_a21oi_1 _3934_ (.A1(_2834_),
    .A2(net83),
    .Y(_0149_),
    .B1(_0148_));
 sg13g2_a21o_1 _3935_ (.A2(_0149_),
    .A1(_0138_),
    .B1(net113),
    .X(_0150_));
 sg13g2_nor2_1 _3936_ (.A(_2814_),
    .B(_0140_),
    .Y(_0151_));
 sg13g2_or3_1 _3937_ (.A(_2822_),
    .B(_2834_),
    .C(_0148_),
    .X(_0152_));
 sg13g2_a22oi_1 _3938_ (.Y(_0153_),
    .B1(_0151_),
    .B2(_0152_),
    .A2(net83),
    .A1(_0130_));
 sg13g2_buf_1 _3939_ (.A(net178),
    .X(_0154_));
 sg13g2_buf_1 _3940_ (.A(net199),
    .X(_0155_));
 sg13g2_a21o_1 _3941_ (.A2(net173),
    .A1(net153),
    .B1(_2556_),
    .X(_0156_));
 sg13g2_o21ai_1 _3942_ (.B1(net157),
    .Y(_0157_),
    .A1(net153),
    .A2(_2802_));
 sg13g2_a21oi_1 _3943_ (.A1(_0156_),
    .A2(_0157_),
    .Y(_0158_),
    .B1(_2786_));
 sg13g2_nand2_1 _3944_ (.Y(_0159_),
    .A(_0151_),
    .B(_0158_));
 sg13g2_a221oi_1 _3945_ (.B2(net86),
    .C1(net65),
    .B1(_0159_),
    .A1(_0150_),
    .Y(_0160_),
    .A2(_0153_));
 sg13g2_a21oi_1 _3946_ (.A1(_0114_),
    .A2(_0139_),
    .Y(_0161_),
    .B1(_0160_));
 sg13g2_nor2_1 _3947_ (.A(net112),
    .B(net83),
    .Y(_0162_));
 sg13g2_nor2_1 _3948_ (.A(net84),
    .B(_0111_),
    .Y(_0163_));
 sg13g2_o21ai_1 _3949_ (.B1(_0163_),
    .Y(_0164_),
    .A1(_0161_),
    .A2(_0162_));
 sg13g2_buf_1 _3950_ (.A(net153),
    .X(_0165_));
 sg13g2_nand2_1 _3951_ (.Y(_0166_),
    .A(net178),
    .B(net154));
 sg13g2_o21ai_1 _3952_ (.B1(_0166_),
    .Y(_0167_),
    .A1(_0165_),
    .A2(_2786_));
 sg13g2_nand3_1 _3953_ (.B(_2831_),
    .C(_0167_),
    .A(net173),
    .Y(_0168_));
 sg13g2_nand2_2 _3954_ (.Y(_0169_),
    .A(_2814_),
    .B(_0140_));
 sg13g2_nor2_1 _3955_ (.A(net85),
    .B(_0169_),
    .Y(_0170_));
 sg13g2_o21ai_1 _3956_ (.B1(_0170_),
    .Y(_0171_),
    .A1(net65),
    .A2(_0168_));
 sg13g2_o21ai_1 _3957_ (.B1(_0171_),
    .Y(_0172_),
    .A1(_0111_),
    .A2(_0162_));
 sg13g2_inv_1 _3958_ (.Y(_0173_),
    .A(_0158_));
 sg13g2_o21ai_1 _3959_ (.B1(_0138_),
    .Y(_0174_),
    .A1(net65),
    .A2(_0173_));
 sg13g2_nor2_1 _3960_ (.A(_2848_),
    .B(_2764_),
    .Y(_0175_));
 sg13g2_nor2_1 _3961_ (.A(_2870_),
    .B(_2888_),
    .Y(_0176_));
 sg13g2_nor2_1 _3962_ (.A(_0175_),
    .B(_0176_),
    .Y(_0177_));
 sg13g2_nor2_1 _3963_ (.A(net66),
    .B(_0177_),
    .Y(_0178_));
 sg13g2_a21oi_1 _3964_ (.A1(_0133_),
    .A2(_0135_),
    .Y(_0179_),
    .B1(_0125_));
 sg13g2_o21ai_1 _3965_ (.B1(_0125_),
    .Y(_0180_),
    .A1(_2776_),
    .A2(_2778_));
 sg13g2_nand2b_1 _3966_ (.Y(_0181_),
    .B(_0180_),
    .A_N(_0179_));
 sg13g2_a221oi_1 _3967_ (.B2(_0181_),
    .C1(_0162_),
    .B1(_0178_),
    .A1(net66),
    .Y(_0182_),
    .A2(_0174_));
 sg13g2_a21oi_1 _3968_ (.A1(net169),
    .A2(_2745_),
    .Y(_0183_),
    .B1(net186));
 sg13g2_o21ai_1 _3969_ (.B1(_0183_),
    .Y(_0184_),
    .A1(net143),
    .A2(_2888_));
 sg13g2_o21ai_1 _3970_ (.B1(net186),
    .Y(_0185_),
    .A1(net143),
    .A2(_2763_));
 sg13g2_and3_1 _3971_ (.X(_0186_),
    .A(net153),
    .B(_0184_),
    .C(_0185_));
 sg13g2_xnor2_1 _3972_ (.Y(_0187_),
    .A(net173),
    .B(_2747_));
 sg13g2_nor2_1 _3973_ (.A(_0154_),
    .B(_2754_),
    .Y(_0188_));
 sg13g2_a21oi_1 _3974_ (.A1(_0143_),
    .A2(_0166_),
    .Y(_0189_),
    .B1(_2556_));
 sg13g2_a21oi_1 _3975_ (.A1(_2786_),
    .A2(_0188_),
    .Y(_0190_),
    .B1(_0189_));
 sg13g2_o21ai_1 _3976_ (.B1(_0114_),
    .Y(_0191_),
    .A1(_0187_),
    .A2(_0190_));
 sg13g2_nor3_1 _3977_ (.A(_0130_),
    .B(_0186_),
    .C(_0191_),
    .Y(_0192_));
 sg13g2_nand2_2 _3978_ (.Y(_0193_),
    .A(_2827_),
    .B(_2828_));
 sg13g2_inv_1 _3979_ (.Y(_0194_),
    .A(net194));
 sg13g2_buf_1 _3980_ (.A(_0194_),
    .X(_0195_));
 sg13g2_nand2_1 _3981_ (.Y(_0196_),
    .A(net179),
    .B(net199));
 sg13g2_nand2_1 _3982_ (.Y(_0197_),
    .A(_2769_),
    .B(_2757_));
 sg13g2_nor2_1 _3983_ (.A(net133),
    .B(_2756_),
    .Y(_0198_));
 sg13g2_a221oi_1 _3984_ (.B2(_0198_),
    .C1(net120),
    .B1(_0197_),
    .A1(net133),
    .Y(_0199_),
    .A2(_0196_));
 sg13g2_o21ai_1 _3985_ (.B1(_2763_),
    .Y(_0200_),
    .A1(net178),
    .A2(_0196_));
 sg13g2_nor3_1 _3986_ (.A(_2609_),
    .B(net178),
    .C(_2763_),
    .Y(_0201_));
 sg13g2_a21o_1 _3987_ (.A2(_0200_),
    .A1(net120),
    .B1(_0201_),
    .X(_0202_));
 sg13g2_o21ai_1 _3988_ (.B1(net157),
    .Y(_0203_),
    .A1(_0199_),
    .A2(_0202_));
 sg13g2_and2_1 _3989_ (.A(net179),
    .B(net199),
    .X(_0204_));
 sg13g2_inv_2 _3990_ (.Y(_0205_),
    .A(net193));
 sg13g2_o21ai_1 _3991_ (.B1(_2764_),
    .Y(_0206_),
    .A1(_0205_),
    .A2(_2763_));
 sg13g2_a22oi_1 _3992_ (.Y(_0207_),
    .B1(_0206_),
    .B2(net186),
    .A2(_0204_),
    .A1(_2965_));
 sg13g2_nand3_1 _3993_ (.B(_0203_),
    .C(_0207_),
    .A(_0193_),
    .Y(_0208_));
 sg13g2_nor2b_1 _3994_ (.A(_0192_),
    .B_N(_0208_),
    .Y(_0209_));
 sg13g2_nand2_1 _3995_ (.Y(_0210_),
    .A(_0203_),
    .B(_0207_));
 sg13g2_nor3_1 _3996_ (.A(_2834_),
    .B(_0176_),
    .C(_0210_),
    .Y(_0211_));
 sg13g2_nor4_1 _3997_ (.A(net98),
    .B(net65),
    .C(_0209_),
    .D(_0211_),
    .Y(_0212_));
 sg13g2_nor3_1 _3998_ (.A(_0172_),
    .B(_0182_),
    .C(_0212_),
    .Y(_0213_));
 sg13g2_or2_1 _3999_ (.X(_0214_),
    .B(_0211_),
    .A(net65));
 sg13g2_xnor2_1 _4000_ (.Y(_0215_),
    .A(net154),
    .B(_2727_));
 sg13g2_xnor2_1 _4001_ (.Y(_0216_),
    .A(_0154_),
    .B(_0215_));
 sg13g2_a21oi_1 _4002_ (.A1(_2783_),
    .A2(_0216_),
    .Y(_0217_),
    .B1(_0189_));
 sg13g2_nor2_1 _4003_ (.A(_0187_),
    .B(_0217_),
    .Y(_0218_));
 sg13g2_and2_1 _4004_ (.A(net198),
    .B(net228),
    .X(_0219_));
 sg13g2_and2_1 _4005_ (.A(_2816_),
    .B(_2997_),
    .X(_0220_));
 sg13g2_a21o_1 _4006_ (.A2(_0219_),
    .A1(net158),
    .B1(_0220_),
    .X(_0221_));
 sg13g2_buf_1 _4007_ (.A(_0221_),
    .X(_0222_));
 sg13g2_nand2_1 _4008_ (.Y(_0223_),
    .A(_0222_),
    .B(_0187_));
 sg13g2_a22oi_1 _4009_ (.Y(_0224_),
    .B1(_0223_),
    .B2(_0130_),
    .A2(_0218_),
    .A1(net113));
 sg13g2_nor2_1 _4010_ (.A(net86),
    .B(net83),
    .Y(_0225_));
 sg13g2_o21ai_1 _4011_ (.B1(_0225_),
    .Y(_0226_),
    .A1(net65),
    .A2(_0224_));
 sg13g2_a21o_1 _4012_ (.A2(_0214_),
    .A1(_0138_),
    .B1(_0226_),
    .X(_0227_));
 sg13g2_a22oi_1 _4013_ (.Y(_0228_),
    .B1(_0213_),
    .B2(_0227_),
    .A2(_0164_),
    .A1(_0112_));
 sg13g2_nand2_1 _4014_ (.Y(_0229_),
    .A(net112),
    .B(net83));
 sg13g2_nand2_1 _4015_ (.Y(_0230_),
    .A(_2838_),
    .B(_2751_));
 sg13g2_nor2_1 _4016_ (.A(_0230_),
    .B(net65),
    .Y(_0231_));
 sg13g2_nand3_1 _4017_ (.B(_0193_),
    .C(_0138_),
    .A(net113),
    .Y(_0232_));
 sg13g2_nor2_1 _4018_ (.A(net112),
    .B(_2922_),
    .Y(_0233_));
 sg13g2_o21ai_1 _4019_ (.B1(_0233_),
    .Y(_0234_),
    .A1(_0231_),
    .A2(_0232_));
 sg13g2_nand3_1 _4020_ (.B(_0229_),
    .C(_0234_),
    .A(net84),
    .Y(_0235_));
 sg13g2_o21ai_1 _4021_ (.B1(_0181_),
    .Y(_0236_),
    .A1(_2928_),
    .A2(_0210_));
 sg13g2_o21ai_1 _4022_ (.B1(_2858_),
    .Y(_0237_),
    .A1(_0233_),
    .A2(_3015_));
 sg13g2_nand3_1 _4023_ (.B(net84),
    .C(_0111_),
    .A(_3010_),
    .Y(_0238_));
 sg13g2_a221oi_1 _4024_ (.B2(_0238_),
    .C1(net5),
    .B1(_0237_),
    .A1(_0138_),
    .Y(_0239_),
    .A2(_0236_));
 sg13g2_o21ai_1 _4025_ (.B1(_0138_),
    .Y(_0240_),
    .A1(_0230_),
    .A2(_0127_));
 sg13g2_a221oi_1 _4026_ (.B2(_0193_),
    .C1(net83),
    .B1(_0240_),
    .A1(_0181_),
    .Y(_0241_),
    .A2(_0158_));
 sg13g2_nand2_1 _4027_ (.Y(_0242_),
    .A(_2819_),
    .B(_0240_));
 sg13g2_nor2_1 _4028_ (.A(net84),
    .B(_0229_),
    .Y(_0243_));
 sg13g2_a22oi_1 _4029_ (.Y(_0244_),
    .B1(_0242_),
    .B2(_0243_),
    .A2(_0241_),
    .A1(net84));
 sg13g2_nand3_1 _4030_ (.B(_0239_),
    .C(_0244_),
    .A(_0235_),
    .Y(_0245_));
 sg13g2_or2_1 _4031_ (.X(_0246_),
    .B(_0245_),
    .A(_0228_));
 sg13g2_inv_1 _4032_ (.Y(_0247_),
    .A(net5));
 sg13g2_and2_1 _4033_ (.A(net222),
    .B(_1101_),
    .X(_0248_));
 sg13g2_buf_2 _4034_ (.A(_0248_),
    .X(_0249_));
 sg13g2_nor2_1 _4035_ (.A(net162),
    .B(_0249_),
    .Y(_0250_));
 sg13g2_nand2_1 _4036_ (.Y(_0251_),
    .A(net222),
    .B(net225));
 sg13g2_inv_1 _4037_ (.Y(_0252_),
    .A(_2728_));
 sg13g2_a21oi_1 _4038_ (.A1(_2560_),
    .A2(_0251_),
    .Y(_0253_),
    .B1(_0252_));
 sg13g2_nor4_1 _4039_ (.A(_1079_),
    .B(net224),
    .C(_2728_),
    .D(_0249_),
    .Y(_0254_));
 sg13g2_nor2b_1 _4040_ (.A(_2729_),
    .B_N(_2741_),
    .Y(_0255_));
 sg13g2_nand3b_1 _4041_ (.B(_1101_),
    .C(net222),
    .Y(_0256_),
    .A_N(_1134_));
 sg13g2_buf_1 _4042_ (.A(_0256_),
    .X(_0257_));
 sg13g2_nor2b_1 _4043_ (.A(_1134_),
    .B_N(_2729_),
    .Y(_0258_));
 sg13g2_nor2b_1 _4044_ (.A(net202),
    .B_N(_2729_),
    .Y(_0259_));
 sg13g2_a221oi_1 _4045_ (.B2(_0249_),
    .C1(_0259_),
    .B1(_0258_),
    .A1(_0255_),
    .Y(_0260_),
    .A2(_0257_));
 sg13g2_buf_1 _4046_ (.A(_0260_),
    .X(_0261_));
 sg13g2_or3_1 _4047_ (.A(_0253_),
    .B(_0254_),
    .C(_0261_),
    .X(_0262_));
 sg13g2_buf_1 _4048_ (.A(_0262_),
    .X(_0263_));
 sg13g2_nor2_1 _4049_ (.A(_0250_),
    .B(net82),
    .Y(_0264_));
 sg13g2_inv_2 _4050_ (.Y(_0265_),
    .A(net219));
 sg13g2_and2_1 _4051_ (.A(net183),
    .B(net167),
    .X(_0266_));
 sg13g2_buf_1 _4052_ (.A(_0266_),
    .X(_0267_));
 sg13g2_nand2_1 _4053_ (.Y(_0268_),
    .A(_0265_),
    .B(net111));
 sg13g2_buf_1 _4054_ (.A(_0268_),
    .X(_0269_));
 sg13g2_buf_1 _4055_ (.A(_0253_),
    .X(_0270_));
 sg13g2_buf_1 _4056_ (.A(_0254_),
    .X(_0271_));
 sg13g2_buf_1 _4057_ (.A(_0261_),
    .X(_0272_));
 sg13g2_nor2_2 _4058_ (.A(net191),
    .B(net137),
    .Y(_0273_));
 sg13g2_nor2_1 _4059_ (.A(net223),
    .B(net192),
    .Y(_0274_));
 sg13g2_buf_2 _4060_ (.A(_0274_),
    .X(_0275_));
 sg13g2_nand3_1 _4061_ (.B(_0273_),
    .C(_0275_),
    .A(_1167_),
    .Y(_0276_));
 sg13g2_or4_1 _4062_ (.A(net132),
    .B(net110),
    .C(net97),
    .D(_0276_),
    .X(_0277_));
 sg13g2_buf_1 _4063_ (.A(_2912_),
    .X(_0278_));
 sg13g2_xor2_1 _4064_ (.B(_2729_),
    .A(net179),
    .X(_0279_));
 sg13g2_buf_2 _4065_ (.A(_0279_),
    .X(_0280_));
 sg13g2_nor2b_1 _4066_ (.A(_2728_),
    .B_N(net224),
    .Y(_0281_));
 sg13g2_buf_1 _4067_ (.A(_0281_),
    .X(_0282_));
 sg13g2_and2_1 _4068_ (.A(_0280_),
    .B(_0282_),
    .X(_0283_));
 sg13g2_buf_1 _4069_ (.A(_0283_),
    .X(_0284_));
 sg13g2_and2_1 _4070_ (.A(net223),
    .B(net194),
    .X(_0285_));
 sg13g2_buf_1 _4071_ (.A(_0285_),
    .X(_0286_));
 sg13g2_nor4_1 _4072_ (.A(_1266_),
    .B(net155),
    .C(net159),
    .D(_0286_),
    .Y(_0287_));
 sg13g2_nor2_1 _4073_ (.A(net155),
    .B(_1463_),
    .Y(_0288_));
 sg13g2_a221oi_1 _4074_ (.B2(_0287_),
    .C1(_0288_),
    .B1(_0284_),
    .A1(net131),
    .Y(_0289_),
    .A2(_1584_));
 sg13g2_nor2_1 _4075_ (.A(net163),
    .B(net155),
    .Y(_0290_));
 sg13g2_xor2_1 _4076_ (.B(_2608_),
    .A(net193),
    .X(_0291_));
 sg13g2_mux2_1 _4077_ (.A0(_0290_),
    .A1(_0291_),
    .S(_1266_),
    .X(_0292_));
 sg13g2_xor2_1 _4078_ (.B(net167),
    .A(net183),
    .X(_0293_));
 sg13g2_a21oi_1 _4079_ (.A1(_0284_),
    .A2(_0292_),
    .Y(_0294_),
    .B1(_0293_));
 sg13g2_a21o_1 _4080_ (.A2(_0289_),
    .A1(_0277_),
    .B1(_0294_),
    .X(_0295_));
 sg13g2_nor2b_2 _4081_ (.A(net194),
    .B_N(_1255_),
    .Y(_0296_));
 sg13g2_nand3_1 _4082_ (.B(_0282_),
    .C(_0296_),
    .A(_0280_),
    .Y(_0297_));
 sg13g2_buf_1 _4083_ (.A(_0297_),
    .X(_0298_));
 sg13g2_a21o_1 _4084_ (.A2(_2612_),
    .A1(net141),
    .B1(_2620_),
    .X(_0299_));
 sg13g2_nand2_1 _4085_ (.Y(_0300_),
    .A(_0298_),
    .B(_0299_));
 sg13g2_nand2_2 _4086_ (.Y(_0301_),
    .A(_2667_),
    .B(net159));
 sg13g2_a21oi_1 _4087_ (.A1(net99),
    .A2(_0298_),
    .Y(_0302_),
    .B1(_0301_));
 sg13g2_o21ai_1 _4088_ (.B1(_0302_),
    .Y(_0303_),
    .A1(net82),
    .A2(_0300_));
 sg13g2_a22oi_1 _4089_ (.Y(_0304_),
    .B1(_0295_),
    .B2(_0303_),
    .A2(_0269_),
    .A1(net197));
 sg13g2_nor2_1 _4090_ (.A(net169),
    .B(net141),
    .Y(_0305_));
 sg13g2_o21ai_1 _4091_ (.B1(net140),
    .Y(_0306_),
    .A1(net142),
    .A2(_0305_));
 sg13g2_nor2_1 _4092_ (.A(net164),
    .B(net182),
    .Y(_0307_));
 sg13g2_nand2b_1 _4093_ (.Y(_0308_),
    .B(_0286_),
    .A_N(_0307_));
 sg13g2_a21oi_1 _4094_ (.A1(_0306_),
    .A2(_0308_),
    .Y(_0309_),
    .B1(net82));
 sg13g2_nor2_1 _4095_ (.A(_0269_),
    .B(_0309_),
    .Y(_0310_));
 sg13g2_inv_2 _4096_ (.Y(_0311_),
    .A(net241));
 sg13g2_o21ai_1 _4097_ (.B1(_0311_),
    .Y(_0312_),
    .A1(_0304_),
    .A2(_0310_));
 sg13g2_nand3_1 _4098_ (.B(_0280_),
    .C(_0251_),
    .A(_0252_),
    .Y(_0313_));
 sg13g2_a21oi_1 _4099_ (.A1(_2621_),
    .A2(_0313_),
    .Y(_0314_),
    .B1(net169));
 sg13g2_nor4_1 _4100_ (.A(net144),
    .B(_0250_),
    .C(net82),
    .D(_0314_),
    .Y(_0315_));
 sg13g2_nor2b_1 _4101_ (.A(net182),
    .B_N(_2608_),
    .Y(_0316_));
 sg13g2_nor2b_1 _4102_ (.A(net194),
    .B_N(net224),
    .Y(_0317_));
 sg13g2_buf_2 _4103_ (.A(_0317_),
    .X(_0318_));
 sg13g2_o21ai_1 _4104_ (.B1(_2612_),
    .Y(_0319_),
    .A1(_0316_),
    .A2(_0318_));
 sg13g2_o21ai_1 _4105_ (.B1(net144),
    .Y(_0320_),
    .A1(net82),
    .A2(_0319_));
 sg13g2_nor2b_1 _4106_ (.A(_0315_),
    .B_N(_0320_),
    .Y(_0321_));
 sg13g2_buf_1 _4107_ (.A(_0265_),
    .X(_0322_));
 sg13g2_a21oi_1 _4108_ (.A1(net165),
    .A2(_0319_),
    .Y(_0323_),
    .B1(net135));
 sg13g2_nor2_1 _4109_ (.A(net152),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_nor3_1 _4110_ (.A(net132),
    .B(net110),
    .C(_0272_),
    .Y(_0325_));
 sg13g2_buf_1 _4111_ (.A(_0205_),
    .X(_0326_));
 sg13g2_nor2_1 _4112_ (.A(net141),
    .B(net115),
    .Y(_0327_));
 sg13g2_a22oi_1 _4113_ (.Y(_0328_),
    .B1(_0327_),
    .B2(net140),
    .A2(_0316_),
    .A1(net142));
 sg13g2_nor2b_1 _4114_ (.A(net142),
    .B_N(net182),
    .Y(_0329_));
 sg13g2_nand2b_1 _4115_ (.Y(_0330_),
    .B(net141),
    .A_N(net137));
 sg13g2_nand3_1 _4116_ (.B(_0329_),
    .C(_0330_),
    .A(_0205_),
    .Y(_0331_));
 sg13g2_o21ai_1 _4117_ (.B1(_0331_),
    .Y(_0332_),
    .A1(net130),
    .A2(_0328_));
 sg13g2_nand3_1 _4118_ (.B(_0325_),
    .C(_0332_),
    .A(net139),
    .Y(_0333_));
 sg13g2_a21oi_1 _4119_ (.A1(net168),
    .A2(_0267_),
    .Y(_0334_),
    .B1(net138));
 sg13g2_nor2_1 _4120_ (.A(net141),
    .B(_2612_),
    .Y(_0335_));
 sg13g2_a21oi_1 _4121_ (.A1(_0284_),
    .A2(_0335_),
    .Y(_0336_),
    .B1(_0269_));
 sg13g2_and2_1 _4122_ (.A(net220),
    .B(net228),
    .X(_0337_));
 sg13g2_nor2_1 _4123_ (.A(net189),
    .B(net197),
    .Y(_0338_));
 sg13g2_a21oi_1 _4124_ (.A1(_0269_),
    .A2(_0337_),
    .Y(_0339_),
    .B1(_0338_));
 sg13g2_nand2b_1 _4125_ (.Y(_0340_),
    .B(_0339_),
    .A_N(_0336_));
 sg13g2_a221oi_1 _4126_ (.B2(_0334_),
    .C1(_0340_),
    .B1(_0333_),
    .A1(_0309_),
    .Y(_0341_),
    .A2(_0324_));
 sg13g2_o21ai_1 _4127_ (.B1(_0341_),
    .Y(_0342_),
    .A1(_0301_),
    .A2(_0321_));
 sg13g2_o21ai_1 _4128_ (.B1(net220),
    .Y(_0343_),
    .A1(net191),
    .A2(_0266_));
 sg13g2_buf_2 _4129_ (.A(_0343_),
    .X(_0344_));
 sg13g2_nand3b_1 _4130_ (.B(net204),
    .C(net205),
    .Y(_0345_),
    .A_N(net195));
 sg13g2_o21ai_1 _4131_ (.B1(net204),
    .Y(_0346_),
    .A1(net205),
    .A2(_0344_));
 sg13g2_nand2b_1 _4132_ (.Y(_0347_),
    .B(net181),
    .A_N(_0344_));
 sg13g2_nand3_1 _4133_ (.B(_0346_),
    .C(_0347_),
    .A(net195),
    .Y(_0348_));
 sg13g2_o21ai_1 _4134_ (.B1(_0348_),
    .Y(_0349_),
    .A1(_0344_),
    .A2(_0345_));
 sg13g2_nand2_1 _4135_ (.Y(_0350_),
    .A(_0269_),
    .B(_0337_));
 sg13g2_a21o_1 _4136_ (.A2(_0303_),
    .A1(_0295_),
    .B1(_0350_),
    .X(_0351_));
 sg13g2_nand4_1 _4137_ (.B(_0342_),
    .C(_0349_),
    .A(_0312_),
    .Y(_0352_),
    .D(_0351_));
 sg13g2_nand3b_1 _4138_ (.B(_1518_),
    .C(_0344_),
    .Y(_0353_),
    .A_N(net205));
 sg13g2_xnor2_1 _4139_ (.Y(_0354_),
    .A(_3011_),
    .B(_0353_));
 sg13g2_nor2_1 _4140_ (.A(net99),
    .B(_0301_),
    .Y(_0355_));
 sg13g2_nor2b_1 _4141_ (.A(net223),
    .B_N(net192),
    .Y(_0356_));
 sg13g2_buf_2 _4142_ (.A(_0356_),
    .X(_0357_));
 sg13g2_and4_1 _4143_ (.A(_0194_),
    .B(_0280_),
    .C(_0282_),
    .D(_0357_),
    .X(_0358_));
 sg13g2_buf_1 _4144_ (.A(_0358_),
    .X(_0359_));
 sg13g2_nand2_2 _4145_ (.Y(_0360_),
    .A(net183),
    .B(net137));
 sg13g2_mux2_1 _4146_ (.A0(_0311_),
    .A1(_0337_),
    .S(_0360_),
    .X(_0361_));
 sg13g2_nor2_1 _4147_ (.A(net159),
    .B(net181),
    .Y(_0362_));
 sg13g2_nand2_1 _4148_ (.Y(_0363_),
    .A(net191),
    .B(net220));
 sg13g2_nand2b_1 _4149_ (.Y(_0364_),
    .B(net228),
    .A_N(net229));
 sg13g2_nor2_1 _4150_ (.A(_0363_),
    .B(_0364_),
    .Y(_0365_));
 sg13g2_a221oi_1 _4151_ (.B2(_0362_),
    .C1(_0365_),
    .B1(_0361_),
    .A1(net204),
    .Y(_0366_),
    .A2(_0338_));
 sg13g2_a21oi_1 _4152_ (.A1(_0355_),
    .A2(_0359_),
    .Y(_0367_),
    .B1(_0366_));
 sg13g2_a21oi_1 _4153_ (.A1(net140),
    .A2(_2760_),
    .Y(_0368_),
    .B1(_1222_));
 sg13g2_or2_1 _4154_ (.X(_0369_),
    .B(_0368_),
    .A(_0250_));
 sg13g2_o21ai_1 _4155_ (.B1(_0288_),
    .Y(_0370_),
    .A1(_0263_),
    .A2(_0369_));
 sg13g2_buf_2 _4156_ (.A(_0021_),
    .X(_0371_));
 sg13g2_inv_2 _4157_ (.Y(_0372_),
    .A(_0371_));
 sg13g2_a21oi_1 _4158_ (.A1(_2612_),
    .A2(_0316_),
    .Y(_0373_),
    .B1(net111));
 sg13g2_nor2b_1 _4159_ (.A(_1255_),
    .B_N(net243),
    .Y(_0374_));
 sg13g2_buf_2 _4160_ (.A(_0374_),
    .X(_0375_));
 sg13g2_o21ai_1 _4161_ (.B1(_0318_),
    .Y(_0376_),
    .A1(_0265_),
    .A2(_0375_));
 sg13g2_o21ai_1 _4162_ (.B1(_0376_),
    .Y(_0377_),
    .A1(net138),
    .A2(_0373_));
 sg13g2_nand4_1 _4163_ (.B(_0293_),
    .C(_0325_),
    .A(_0372_),
    .Y(_0378_),
    .D(_0377_));
 sg13g2_nand2_1 _4164_ (.Y(_0379_),
    .A(_1167_),
    .B(_0275_));
 sg13g2_nor4_2 _4165_ (.A(net132),
    .B(net110),
    .C(net97),
    .Y(_0380_),
    .D(_0379_));
 sg13g2_and3_1 _4166_ (.X(_0381_),
    .A(_0252_),
    .B(_1167_),
    .C(_0280_));
 sg13g2_nand2_1 _4167_ (.Y(_0382_),
    .A(net138),
    .B(_0381_));
 sg13g2_o21ai_1 _4168_ (.B1(net163),
    .Y(_0383_),
    .A1(net223),
    .A2(net164));
 sg13g2_buf_1 _4169_ (.A(_0383_),
    .X(_0384_));
 sg13g2_or3_1 _4170_ (.A(net243),
    .B(net192),
    .C(_1112_),
    .X(_0385_));
 sg13g2_nand4_1 _4171_ (.B(_0282_),
    .C(_0384_),
    .A(_0280_),
    .Y(_0386_),
    .D(_0385_));
 sg13g2_a21oi_1 _4172_ (.A1(net152),
    .A2(_0386_),
    .Y(_0387_),
    .B1(_0360_));
 sg13g2_o21ai_1 _4173_ (.B1(_0387_),
    .Y(_0388_),
    .A1(_0380_),
    .A2(_0382_));
 sg13g2_nand4_1 _4174_ (.B(_0370_),
    .C(_0378_),
    .A(_0367_),
    .Y(_0389_),
    .D(_0388_));
 sg13g2_xnor2_1 _4175_ (.Y(_0390_),
    .A(net195),
    .B(_0346_));
 sg13g2_nand2_1 _4176_ (.Y(_0391_),
    .A(_0389_),
    .B(_0390_));
 sg13g2_nand2_1 _4177_ (.Y(_0392_),
    .A(_0375_),
    .B(_0318_));
 sg13g2_or4_1 _4178_ (.A(net132),
    .B(net110),
    .C(_0261_),
    .D(_0392_),
    .X(_0393_));
 sg13g2_buf_1 _4179_ (.A(_0393_),
    .X(_0394_));
 sg13g2_nor2b_1 _4180_ (.A(net155),
    .B_N(net142),
    .Y(_0395_));
 sg13g2_nor2b_1 _4181_ (.A(net164),
    .B_N(net183),
    .Y(_0396_));
 sg13g2_o21ai_1 _4182_ (.B1(net169),
    .Y(_0397_),
    .A1(_0395_),
    .A2(_0396_));
 sg13g2_nand2b_1 _4183_ (.Y(_0398_),
    .B(_0318_),
    .A_N(_0396_));
 sg13g2_nor4_1 _4184_ (.A(net132),
    .B(net110),
    .C(net97),
    .D(_0398_),
    .Y(_0399_));
 sg13g2_nand2_1 _4185_ (.Y(_0400_),
    .A(_0280_),
    .B(_0282_));
 sg13g2_nand2b_1 _4186_ (.Y(_0401_),
    .B(net142),
    .A_N(net169));
 sg13g2_a21oi_1 _4187_ (.A1(net141),
    .A2(_0401_),
    .Y(_0402_),
    .B1(_0395_));
 sg13g2_nor2_1 _4188_ (.A(_0400_),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_o21ai_1 _4189_ (.B1(_0403_),
    .Y(_0404_),
    .A1(_0397_),
    .A2(_0399_));
 sg13g2_a21oi_1 _4190_ (.A1(_0394_),
    .A2(_0404_),
    .Y(_0405_),
    .B1(_0269_));
 sg13g2_o21ai_1 _4191_ (.B1(net161),
    .Y(_0406_),
    .A1(net185),
    .A2(_0372_));
 sg13g2_o21ai_1 _4192_ (.B1(_0406_),
    .Y(_0407_),
    .A1(net99),
    .A2(_0371_));
 sg13g2_a22oi_1 _4193_ (.Y(_0408_),
    .B1(_0407_),
    .B2(net152),
    .A2(_1584_),
    .A1(_2913_));
 sg13g2_nand4_1 _4194_ (.B(net185),
    .C(_0375_),
    .A(_2667_),
    .Y(_0409_),
    .D(_0318_));
 sg13g2_nor4_1 _4195_ (.A(net132),
    .B(net110),
    .C(net97),
    .D(_0409_),
    .Y(_0410_));
 sg13g2_nand3_1 _4196_ (.B(net111),
    .C(_0318_),
    .A(_0375_),
    .Y(_0411_));
 sg13g2_nor4_1 _4197_ (.A(_0270_),
    .B(_0271_),
    .C(net97),
    .D(_0411_),
    .Y(_0412_));
 sg13g2_nor3_1 _4198_ (.A(net131),
    .B(net99),
    .C(_0298_),
    .Y(_0413_));
 sg13g2_nor4_1 _4199_ (.A(_0380_),
    .B(_0410_),
    .C(_0412_),
    .D(_0413_),
    .Y(_0414_));
 sg13g2_nand2b_1 _4200_ (.Y(_0415_),
    .B(net220),
    .A_N(net191));
 sg13g2_mux2_1 _4201_ (.A0(net189),
    .A1(_0415_),
    .S(net203),
    .X(_0416_));
 sg13g2_nand3_1 _4202_ (.B(_0311_),
    .C(net197),
    .A(net159),
    .Y(_0417_));
 sg13g2_o21ai_1 _4203_ (.B1(_0417_),
    .Y(_0418_),
    .A1(net111),
    .A2(_0416_));
 sg13g2_nand2_1 _4204_ (.Y(_0419_),
    .A(_2675_),
    .B(net203));
 sg13g2_nand2_1 _4205_ (.Y(_0420_),
    .A(_1540_),
    .B(net181));
 sg13g2_a21oi_1 _4206_ (.A1(_0269_),
    .A2(_0419_),
    .Y(_0421_),
    .B1(_0420_));
 sg13g2_a21o_1 _4207_ (.A2(_0418_),
    .A1(net204),
    .B1(_0421_),
    .X(_0422_));
 sg13g2_o21ai_1 _4208_ (.B1(_0422_),
    .Y(_0423_),
    .A1(_0408_),
    .A2(_0414_));
 sg13g2_buf_1 _4209_ (.A(net99),
    .X(_0424_));
 sg13g2_and2_1 _4210_ (.A(net165),
    .B(_0394_),
    .X(_0425_));
 sg13g2_a221oi_1 _4211_ (.B2(_0425_),
    .C1(_0301_),
    .B1(_0404_),
    .A1(net81),
    .Y(_0426_),
    .A2(_0298_));
 sg13g2_nor3_1 _4212_ (.A(_0405_),
    .B(_0423_),
    .C(_0426_),
    .Y(_0427_));
 sg13g2_nand2_1 _4213_ (.Y(_0428_),
    .A(net99),
    .B(_0381_));
 sg13g2_nand2_1 _4214_ (.Y(_0429_),
    .A(_0278_),
    .B(_0265_));
 sg13g2_a21oi_1 _4215_ (.A1(net165),
    .A2(_0298_),
    .Y(_0430_),
    .B1(_0429_));
 sg13g2_o21ai_1 _4216_ (.B1(_0430_),
    .Y(_0431_),
    .A1(_0380_),
    .A2(_0428_));
 sg13g2_nor2b_1 _4217_ (.A(net141),
    .B_N(_1211_),
    .Y(_0432_));
 sg13g2_nor2_1 _4218_ (.A(net133),
    .B(net111),
    .Y(_0433_));
 sg13g2_a22oi_1 _4219_ (.Y(_0434_),
    .B1(_0433_),
    .B2(net130),
    .A2(_0432_),
    .A1(net165));
 sg13g2_nand2_1 _4220_ (.Y(_0435_),
    .A(_1277_),
    .B(_0265_));
 sg13g2_or3_1 _4221_ (.A(_0400_),
    .B(_0434_),
    .C(_0435_),
    .X(_0436_));
 sg13g2_nand2_1 _4222_ (.Y(_0437_),
    .A(_0372_),
    .B(_0293_));
 sg13g2_nand4_1 _4223_ (.B(_0280_),
    .C(_0282_),
    .A(net111),
    .Y(_0438_),
    .D(_0296_));
 sg13g2_o21ai_1 _4224_ (.B1(_0438_),
    .Y(_0439_),
    .A1(_0437_),
    .A2(_0386_));
 sg13g2_o21ai_1 _4225_ (.B1(net117),
    .Y(_0440_),
    .A1(_0410_),
    .A2(_0439_));
 sg13g2_nand4_1 _4226_ (.B(_0422_),
    .C(_0436_),
    .A(_0431_),
    .Y(_0441_),
    .D(_0440_));
 sg13g2_and2_1 _4227_ (.A(net115),
    .B(_0298_),
    .X(_0442_));
 sg13g2_nand3_1 _4228_ (.B(_0360_),
    .C(_0318_),
    .A(_0375_),
    .Y(_0443_));
 sg13g2_or4_1 _4229_ (.A(_0270_),
    .B(_0271_),
    .C(_0272_),
    .D(_0443_),
    .X(_0444_));
 sg13g2_and2_1 _4230_ (.A(_0265_),
    .B(_0298_),
    .X(_0445_));
 sg13g2_nand2b_1 _4231_ (.Y(_0446_),
    .B(net191),
    .A_N(net190));
 sg13g2_buf_2 _4232_ (.A(_0446_),
    .X(_0447_));
 sg13g2_nand2b_1 _4233_ (.Y(_0448_),
    .B(net190),
    .A_N(net219));
 sg13g2_buf_1 _4234_ (.A(_0448_),
    .X(_0449_));
 sg13g2_nand2_1 _4235_ (.Y(_0450_),
    .A(net161),
    .B(_0449_));
 sg13g2_o21ai_1 _4236_ (.B1(_0450_),
    .Y(_0451_),
    .A1(_0359_),
    .A2(_0447_));
 sg13g2_a221oi_1 _4237_ (.B2(_0445_),
    .C1(_0451_),
    .B1(_0444_),
    .A1(_0442_),
    .Y(_0452_),
    .A2(_0394_));
 sg13g2_nand2_1 _4238_ (.Y(_0453_),
    .A(_0360_),
    .B(_0291_));
 sg13g2_nand3_1 _4239_ (.B(_0290_),
    .C(_0357_),
    .A(net115),
    .Y(_0454_));
 sg13g2_o21ai_1 _4240_ (.B1(_0454_),
    .Y(_0455_),
    .A1(net120),
    .A2(_0453_));
 sg13g2_nor2_1 _4241_ (.A(net152),
    .B(_0400_),
    .Y(_0456_));
 sg13g2_nor2_1 _4242_ (.A(net159),
    .B(_0311_),
    .Y(_0457_));
 sg13g2_nor2_1 _4243_ (.A(net229),
    .B(net228),
    .Y(_0458_));
 sg13g2_mux2_1 _4244_ (.A0(net229),
    .A1(_0458_),
    .S(_0360_),
    .X(_0459_));
 sg13g2_nand3b_1 _4245_ (.B(net229),
    .C(net220),
    .Y(_0460_),
    .A_N(net197));
 sg13g2_o21ai_1 _4246_ (.B1(_0460_),
    .Y(_0461_),
    .A1(net189),
    .A2(_0364_));
 sg13g2_nor3_1 _4247_ (.A(net189),
    .B(net111),
    .C(_0364_),
    .Y(_0462_));
 sg13g2_a221oi_1 _4248_ (.B2(net138),
    .C1(_0462_),
    .B1(_0461_),
    .A1(_0457_),
    .Y(_0463_),
    .A2(_0459_));
 sg13g2_a221oi_1 _4249_ (.B2(_0456_),
    .C1(_0463_),
    .B1(_0455_),
    .A1(_0380_),
    .Y(_0464_),
    .A2(_0288_));
 sg13g2_nand2b_1 _4250_ (.Y(_0465_),
    .B(_0464_),
    .A_N(_0452_));
 sg13g2_and2_1 _4251_ (.A(_0371_),
    .B(_0293_),
    .X(_0466_));
 sg13g2_nor2b_1 _4252_ (.A(_0466_),
    .B_N(net205),
    .Y(_0467_));
 sg13g2_o21ai_1 _4253_ (.B1(net204),
    .Y(_0468_),
    .A1(_0344_),
    .A2(_0467_));
 sg13g2_buf_1 _4254_ (.A(net180),
    .X(_0469_));
 sg13g2_o21ai_1 _4255_ (.B1(net145),
    .Y(_0470_),
    .A1(net151),
    .A2(_0432_));
 sg13g2_o21ai_1 _4256_ (.B1(_0470_),
    .Y(_0471_),
    .A1(net140),
    .A2(_0286_));
 sg13g2_o21ai_1 _4257_ (.B1(_0355_),
    .Y(_0472_),
    .A1(_0263_),
    .A2(_0471_));
 sg13g2_and2_1 _4258_ (.A(_0447_),
    .B(_0449_),
    .X(_0473_));
 sg13g2_buf_1 _4259_ (.A(_0473_),
    .X(_0474_));
 sg13g2_nand2_1 _4260_ (.Y(_0475_),
    .A(net162),
    .B(_0384_));
 sg13g2_nand2_1 _4261_ (.Y(_0476_),
    .A(_2612_),
    .B(_0316_));
 sg13g2_nor2_1 _4262_ (.A(net155),
    .B(_1584_),
    .Y(_0477_));
 sg13g2_a221oi_1 _4263_ (.B2(_0476_),
    .C1(_0477_),
    .B1(_0475_),
    .A1(net131),
    .Y(_0478_),
    .A2(_0474_));
 sg13g2_nand3_1 _4264_ (.B(_0267_),
    .C(_0296_),
    .A(net159),
    .Y(_0479_));
 sg13g2_o21ai_1 _4265_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0435_),
    .A2(_0453_));
 sg13g2_nor3_1 _4266_ (.A(_2694_),
    .B(net203),
    .C(_0363_),
    .Y(_0481_));
 sg13g2_nor3_1 _4267_ (.A(net111),
    .B(_0415_),
    .C(_0364_),
    .Y(_0482_));
 sg13g2_nor4_1 _4268_ (.A(_2675_),
    .B(net189),
    .C(net229),
    .D(_0360_),
    .Y(_0483_));
 sg13g2_nor3_1 _4269_ (.A(net189),
    .B(net229),
    .C(net197),
    .Y(_0484_));
 sg13g2_nor4_1 _4270_ (.A(_0481_),
    .B(_0482_),
    .C(_0483_),
    .D(_0484_),
    .Y(_0485_));
 sg13g2_a221oi_1 _4271_ (.B2(_0284_),
    .C1(_0485_),
    .B1(_0480_),
    .A1(_0325_),
    .Y(_0486_),
    .A2(_0478_));
 sg13g2_a21oi_1 _4272_ (.A1(_0344_),
    .A2(_0466_),
    .Y(_0487_),
    .B1(net204));
 sg13g2_nor3_1 _4273_ (.A(net205),
    .B(_0344_),
    .C(_0466_),
    .Y(_0488_));
 sg13g2_nor3_1 _4274_ (.A(_2855_),
    .B(_0487_),
    .C(_0488_),
    .Y(_0489_));
 sg13g2_a221oi_1 _4275_ (.B2(_0486_),
    .C1(_0489_),
    .B1(_0472_),
    .A1(net195),
    .Y(_0490_),
    .A2(_0468_));
 sg13g2_nor3_1 _4276_ (.A(net165),
    .B(_0301_),
    .C(_0394_),
    .Y(_0491_));
 sg13g2_nand2_1 _4277_ (.Y(_0492_),
    .A(net135),
    .B(_0359_));
 sg13g2_nand2b_1 _4278_ (.Y(_0493_),
    .B(net161),
    .A_N(_0386_));
 sg13g2_a21oi_1 _4279_ (.A1(_0492_),
    .A2(_0493_),
    .Y(_0494_),
    .B1(_0447_));
 sg13g2_or3_1 _4280_ (.A(_0366_),
    .B(_0491_),
    .C(_0494_),
    .X(_0495_));
 sg13g2_nand4_1 _4281_ (.B(_0465_),
    .C(_0490_),
    .A(_0441_),
    .Y(_0496_),
    .D(_0495_));
 sg13g2_o21ai_1 _4282_ (.B1(_0496_),
    .Y(_0497_),
    .A1(_0391_),
    .A2(_0427_));
 sg13g2_nand4_1 _4283_ (.B(_0352_),
    .C(_0354_),
    .A(_0264_),
    .Y(_0498_),
    .D(_0497_));
 sg13g2_xnor2_1 _4284_ (.Y(_0499_),
    .A(net245),
    .B(net244));
 sg13g2_nand3_1 _4285_ (.B(_1167_),
    .C(_0499_),
    .A(net174),
    .Y(_0500_));
 sg13g2_buf_1 _4286_ (.A(_0500_),
    .X(_0501_));
 sg13g2_nor3_2 _4287_ (.A(_2618_),
    .B(_1090_),
    .C(net200),
    .Y(_0502_));
 sg13g2_nand2_1 _4288_ (.Y(_0503_),
    .A(_0275_),
    .B(_0502_));
 sg13g2_buf_2 _4289_ (.A(_0503_),
    .X(_0504_));
 sg13g2_nor4_1 _4290_ (.A(net163),
    .B(_2618_),
    .C(_1090_),
    .D(net200),
    .Y(_0505_));
 sg13g2_buf_1 _4291_ (.A(_0505_),
    .X(_0506_));
 sg13g2_nand2_1 _4292_ (.Y(_0507_),
    .A(_0205_),
    .B(_1266_));
 sg13g2_and4_1 _4293_ (.A(_2619_),
    .B(net174),
    .C(_0249_),
    .D(_0499_),
    .X(_0508_));
 sg13g2_buf_1 _4294_ (.A(_0508_),
    .X(_0509_));
 sg13g2_a221oi_1 _4295_ (.B2(_0507_),
    .C1(_0509_),
    .B1(net109),
    .A1(_2668_),
    .Y(_0510_),
    .A2(_0504_));
 sg13g2_o21ai_1 _4296_ (.B1(_0510_),
    .Y(_0511_),
    .A1(_1288_),
    .A2(_0501_));
 sg13g2_nor3_1 _4297_ (.A(_2913_),
    .B(_1288_),
    .C(_0501_),
    .Y(_0512_));
 sg13g2_nor2_1 _4298_ (.A(_0449_),
    .B(_0512_),
    .Y(_0513_));
 sg13g2_nand2_1 _4299_ (.Y(_0514_),
    .A(_0384_),
    .B(_0502_));
 sg13g2_o21ai_1 _4300_ (.B1(_0514_),
    .Y(_0515_),
    .A1(_0275_),
    .A2(_0501_));
 sg13g2_and2_1 _4301_ (.A(_0275_),
    .B(_0502_),
    .X(_0516_));
 sg13g2_buf_1 _4302_ (.A(_0516_),
    .X(_0517_));
 sg13g2_nand2_1 _4303_ (.Y(_0518_),
    .A(net131),
    .B(_0357_));
 sg13g2_nand2_1 _4304_ (.Y(_0519_),
    .A(_0397_),
    .B(_0518_));
 sg13g2_a221oi_1 _4305_ (.B2(_0519_),
    .C1(_0447_),
    .B1(_0506_),
    .A1(_0290_),
    .Y(_0520_),
    .A2(_0517_));
 sg13g2_and2_1 _4306_ (.A(_2707_),
    .B(_0273_),
    .X(_0521_));
 sg13g2_nand3_1 _4307_ (.B(_0507_),
    .C(net109),
    .A(_2667_),
    .Y(_0522_));
 sg13g2_nand2_1 _4308_ (.Y(_0523_),
    .A(_0504_),
    .B(_0522_));
 sg13g2_o21ai_1 _4309_ (.B1(_1584_),
    .Y(_0524_),
    .A1(_0371_),
    .A2(_0504_));
 sg13g2_nor2_1 _4310_ (.A(net196),
    .B(_0273_),
    .Y(_0525_));
 sg13g2_a22oi_1 _4311_ (.Y(_0526_),
    .B1(_0524_),
    .B2(_0525_),
    .A2(_0523_),
    .A1(_0521_));
 sg13g2_a221oi_1 _4312_ (.B2(_0520_),
    .C1(_0526_),
    .B1(_0515_),
    .A1(_0511_),
    .Y(_0527_),
    .A2(_0513_));
 sg13g2_nand2_1 _4313_ (.Y(_0528_),
    .A(net196),
    .B(_1463_));
 sg13g2_nor2_1 _4314_ (.A(_0195_),
    .B(_0504_),
    .Y(_0529_));
 sg13g2_nor3_1 _4315_ (.A(_2707_),
    .B(_0371_),
    .C(_1463_),
    .Y(_0530_));
 sg13g2_o21ai_1 _4316_ (.B1(_0530_),
    .Y(_0531_),
    .A1(_0509_),
    .A2(_0529_));
 sg13g2_nand2_1 _4317_ (.Y(_0532_),
    .A(net100),
    .B(_0522_));
 sg13g2_nand3_1 _4318_ (.B(_0507_),
    .C(net109),
    .A(_1584_),
    .Y(_0533_));
 sg13g2_o21ai_1 _4319_ (.B1(_0533_),
    .Y(_0534_),
    .A1(net100),
    .A2(_0504_));
 sg13g2_nand3_1 _4320_ (.B(_0507_),
    .C(net109),
    .A(net165),
    .Y(_0535_));
 sg13g2_nand2_1 _4321_ (.Y(_0536_),
    .A(_2902_),
    .B(_0517_));
 sg13g2_a21oi_1 _4322_ (.A1(_0535_),
    .A2(_0536_),
    .Y(_0537_),
    .B1(net114));
 sg13g2_a221oi_1 _4323_ (.B2(net114),
    .C1(_0537_),
    .B1(_0534_),
    .A1(net152),
    .Y(_0538_),
    .A2(_0532_));
 sg13g2_a21oi_1 _4324_ (.A1(_0528_),
    .A2(_0531_),
    .Y(_0539_),
    .B1(_0538_));
 sg13g2_nand2_1 _4325_ (.Y(_0540_),
    .A(_2810_),
    .B(_2579_));
 sg13g2_xnor2_1 _4326_ (.Y(_0541_),
    .A(net229),
    .B(_0540_));
 sg13g2_o21ai_1 _4327_ (.B1(_0541_),
    .Y(_0542_),
    .A1(_0527_),
    .A2(_0539_));
 sg13g2_nand2_2 _4328_ (.Y(_0543_),
    .A(net138),
    .B(net115));
 sg13g2_a21oi_1 _4329_ (.A1(net145),
    .A2(_0501_),
    .Y(_0544_),
    .B1(net130));
 sg13g2_nor2_1 _4330_ (.A(net135),
    .B(_0544_),
    .Y(_0545_));
 sg13g2_nor2b_1 _4331_ (.A(net109),
    .B_N(_0395_),
    .Y(_0546_));
 sg13g2_inv_1 _4332_ (.Y(_0547_),
    .A(net200));
 sg13g2_nor2_1 _4333_ (.A(_1123_),
    .B(net224),
    .Y(_0548_));
 sg13g2_nand3_1 _4334_ (.B(_0547_),
    .C(_0548_),
    .A(_2553_),
    .Y(_0549_));
 sg13g2_nand2_1 _4335_ (.Y(_0550_),
    .A(net135),
    .B(_0549_));
 sg13g2_nand2_1 _4336_ (.Y(_0551_),
    .A(net131),
    .B(_2612_));
 sg13g2_a21oi_1 _4337_ (.A1(_0550_),
    .A2(_0551_),
    .Y(_0552_),
    .B1(_0509_));
 sg13g2_nor3_1 _4338_ (.A(_0545_),
    .B(_0546_),
    .C(_0552_),
    .Y(_0553_));
 sg13g2_o21ai_1 _4339_ (.B1(_0447_),
    .Y(_0554_),
    .A1(_0371_),
    .A2(_0449_));
 sg13g2_nor2b_1 _4340_ (.A(_0529_),
    .B_N(_0554_),
    .Y(_0555_));
 sg13g2_and2_1 _4341_ (.A(_0384_),
    .B(_0502_),
    .X(_0556_));
 sg13g2_nand2_1 _4342_ (.Y(_0557_),
    .A(_0556_),
    .B(_0530_));
 sg13g2_a22oi_1 _4343_ (.Y(_0558_),
    .B1(_0557_),
    .B2(_0528_),
    .A2(_0555_),
    .A1(_0515_));
 sg13g2_o21ai_1 _4344_ (.B1(_0558_),
    .Y(_0559_),
    .A1(_0543_),
    .A2(_0553_));
 sg13g2_nand2b_1 _4345_ (.Y(_0560_),
    .B(net115),
    .A_N(_2707_));
 sg13g2_nand4_1 _4346_ (.B(net165),
    .C(_0375_),
    .A(net131),
    .Y(_0561_),
    .D(net109));
 sg13g2_a21oi_1 _4347_ (.A1(_0560_),
    .A2(_0561_),
    .Y(_0562_),
    .B1(net138));
 sg13g2_nor3_1 _4348_ (.A(_1288_),
    .B(_0549_),
    .C(_0560_),
    .Y(_0563_));
 sg13g2_nand3_1 _4349_ (.B(_0357_),
    .C(net109),
    .A(_0273_),
    .Y(_0564_));
 sg13g2_a21oi_1 _4350_ (.A1(net196),
    .A2(_0564_),
    .Y(_0565_),
    .B1(net135));
 sg13g2_nor3_1 _4351_ (.A(_0562_),
    .B(_0563_),
    .C(_0565_),
    .Y(_0566_));
 sg13g2_nor2_1 _4352_ (.A(net99),
    .B(net196),
    .Y(_0567_));
 sg13g2_nand3_1 _4353_ (.B(_0251_),
    .C(_0502_),
    .A(_0205_),
    .Y(_0568_));
 sg13g2_or2_1 _4354_ (.X(_0569_),
    .B(_0568_),
    .A(_2565_));
 sg13g2_a21oi_1 _4355_ (.A1(_2565_),
    .A2(net196),
    .Y(_0570_),
    .B1(_2676_));
 sg13g2_nor3_1 _4356_ (.A(net144),
    .B(_0301_),
    .C(_0556_),
    .Y(_0571_));
 sg13g2_a221oi_1 _4357_ (.B2(_0570_),
    .C1(_0571_),
    .B1(_0569_),
    .A1(_0504_),
    .Y(_0572_),
    .A2(_0567_));
 sg13g2_nand2b_1 _4358_ (.Y(_0573_),
    .B(_0572_),
    .A_N(_0566_));
 sg13g2_a21o_1 _4359_ (.A2(_0573_),
    .A1(_0559_),
    .B1(_0541_),
    .X(_0574_));
 sg13g2_nand2_1 _4360_ (.Y(_0575_),
    .A(_0514_),
    .B(_0501_));
 sg13g2_xor2_1 _4361_ (.B(_3011_),
    .A(_1507_),
    .X(_0576_));
 sg13g2_nand2_1 _4362_ (.Y(_0577_),
    .A(net195),
    .B(_0576_));
 sg13g2_nand3b_1 _4363_ (.B(_3011_),
    .C(_1496_),
    .Y(_0578_),
    .A_N(net195));
 sg13g2_o21ai_1 _4364_ (.B1(_0578_),
    .Y(_0579_),
    .A1(_1496_),
    .A2(_0577_));
 sg13g2_nand2_1 _4365_ (.Y(_0580_),
    .A(_0575_),
    .B(_0579_));
 sg13g2_a21o_1 _4366_ (.A2(_0574_),
    .A1(_0542_),
    .B1(_0580_),
    .X(_0581_));
 sg13g2_nand3_1 _4367_ (.B(net176),
    .C(_2693_),
    .A(_1375_),
    .Y(_0582_));
 sg13g2_nand2_1 _4368_ (.Y(_0583_),
    .A(_2810_),
    .B(_2695_));
 sg13g2_a21oi_1 _4369_ (.A1(_0582_),
    .A2(_0583_),
    .Y(_0584_),
    .B1(net115));
 sg13g2_o21ai_1 _4370_ (.B1(net159),
    .Y(_0585_),
    .A1(_1540_),
    .A2(net204));
 sg13g2_nand2_1 _4371_ (.Y(_0586_),
    .A(net152),
    .B(_0420_));
 sg13g2_o21ai_1 _4372_ (.B1(_0586_),
    .Y(_0587_),
    .A1(_0584_),
    .A2(_0585_));
 sg13g2_nand3_1 _4373_ (.B(net189),
    .C(_1584_),
    .A(net240),
    .Y(_0588_));
 sg13g2_xnor2_1 _4374_ (.Y(_0589_),
    .A(_1507_),
    .B(_0588_));
 sg13g2_nand4_1 _4375_ (.B(net224),
    .C(_2553_),
    .A(_1079_),
    .Y(_0590_),
    .D(_0385_));
 sg13g2_nor2b_1 _4376_ (.A(net245),
    .B_N(net244),
    .Y(_0591_));
 sg13g2_o21ai_1 _4377_ (.B1(net162),
    .Y(_0592_),
    .A1(net193),
    .A2(net163));
 sg13g2_nand3_1 _4378_ (.B(_0591_),
    .C(_0592_),
    .A(_1266_),
    .Y(_0593_));
 sg13g2_nand2_1 _4379_ (.Y(_0594_),
    .A(net193),
    .B(net199));
 sg13g2_nor2b_1 _4380_ (.A(net194),
    .B_N(_0022_),
    .Y(_0595_));
 sg13g2_buf_2 _4381_ (.A(_0595_),
    .X(_0596_));
 sg13g2_nand2_1 _4382_ (.Y(_0597_),
    .A(_0329_),
    .B(_0596_));
 sg13g2_o21ai_1 _4383_ (.B1(_0597_),
    .Y(_0598_),
    .A1(_2620_),
    .A2(_0596_));
 sg13g2_a22oi_1 _4384_ (.Y(_0599_),
    .B1(_0594_),
    .B2(_0598_),
    .A2(_0593_),
    .A1(_0590_));
 sg13g2_nand3_1 _4385_ (.B(_0589_),
    .C(_0599_),
    .A(_0587_),
    .Y(_0600_));
 sg13g2_nor2_1 _4386_ (.A(net175),
    .B(_0363_),
    .Y(_0601_));
 sg13g2_xnor2_1 _4387_ (.Y(_0602_),
    .A(net181),
    .B(_0601_));
 sg13g2_nand2b_1 _4388_ (.Y(_0603_),
    .B(_0602_),
    .A_N(_0600_));
 sg13g2_nor3_1 _4389_ (.A(net223),
    .B(net164),
    .C(net163),
    .Y(_0604_));
 sg13g2_o21ai_1 _4390_ (.B1(_0591_),
    .Y(_0605_),
    .A1(_2725_),
    .A2(_0604_));
 sg13g2_and2_1 _4391_ (.A(_0590_),
    .B(_0605_),
    .X(_0606_));
 sg13g2_buf_2 _4392_ (.A(_0606_),
    .X(_0607_));
 sg13g2_nor2_1 _4393_ (.A(_1595_),
    .B(_0607_),
    .Y(_0608_));
 sg13g2_nand2_1 _4394_ (.Y(_0609_),
    .A(_0307_),
    .B(_0596_));
 sg13g2_o21ai_1 _4395_ (.B1(_0609_),
    .Y(_0610_),
    .A1(net151),
    .A2(_0596_));
 sg13g2_nand2_1 _4396_ (.Y(_0611_),
    .A(_2799_),
    .B(_0610_));
 sg13g2_nor2_1 _4397_ (.A(net151),
    .B(net173),
    .Y(_0612_));
 sg13g2_nor2_1 _4398_ (.A(net145),
    .B(_0469_),
    .Y(_0613_));
 sg13g2_a221oi_1 _4399_ (.B2(net143),
    .C1(net114),
    .B1(_0613_),
    .A1(_0357_),
    .Y(_0614_),
    .A2(_0612_));
 sg13g2_and2_1 _4400_ (.A(net130),
    .B(_0610_),
    .X(_0615_));
 sg13g2_o21ai_1 _4401_ (.B1(net173),
    .Y(_0616_),
    .A1(_0613_),
    .A2(_0615_));
 sg13g2_a22oi_1 _4402_ (.Y(_0617_),
    .B1(_0616_),
    .B2(net114),
    .A2(_0614_),
    .A1(_0611_));
 sg13g2_a22oi_1 _4403_ (.Y(_0618_),
    .B1(_0608_),
    .B2(_0617_),
    .A2(_0543_),
    .A1(_0311_));
 sg13g2_inv_1 _4404_ (.Y(_0619_),
    .A(_0022_));
 sg13g2_o21ai_1 _4405_ (.B1(net162),
    .Y(_0620_),
    .A1(_0619_),
    .A2(_2558_));
 sg13g2_nand2_1 _4406_ (.Y(_0621_),
    .A(_0609_),
    .B(_0620_));
 sg13g2_nor2b_1 _4407_ (.A(_0607_),
    .B_N(_0621_),
    .Y(_0622_));
 sg13g2_nand2_1 _4408_ (.Y(_0623_),
    .A(_2606_),
    .B(net173));
 sg13g2_xnor2_1 _4409_ (.Y(_0624_),
    .A(_2619_),
    .B(_0596_));
 sg13g2_nor2_1 _4410_ (.A(_2605_),
    .B(_2798_),
    .Y(_0625_));
 sg13g2_o21ai_1 _4411_ (.B1(_0625_),
    .Y(_0626_),
    .A1(net130),
    .A2(_0624_));
 sg13g2_a21oi_1 _4412_ (.A1(_0623_),
    .A2(_0626_),
    .Y(_0627_),
    .B1(_0449_));
 sg13g2_nand3_1 _4413_ (.B(net173),
    .C(_0622_),
    .A(net130),
    .Y(_0628_));
 sg13g2_inv_1 _4414_ (.Y(_0629_),
    .A(_0447_));
 sg13g2_nand2b_1 _4415_ (.Y(_0630_),
    .B(_0022_),
    .A_N(net163));
 sg13g2_a22oi_1 _4416_ (.Y(_0631_),
    .B1(_0630_),
    .B2(_0329_),
    .A2(_0357_),
    .A1(net162));
 sg13g2_a21oi_1 _4417_ (.A1(_0609_),
    .A2(_0631_),
    .Y(_0632_),
    .B1(_2798_));
 sg13g2_o21ai_1 _4418_ (.B1(net140),
    .Y(_0633_),
    .A1(net142),
    .A2(_0596_));
 sg13g2_nand3_1 _4419_ (.B(net180),
    .C(_0630_),
    .A(net145),
    .Y(_0634_));
 sg13g2_a21o_1 _4420_ (.A2(_0634_),
    .A1(_0633_),
    .B1(_0594_),
    .X(_0635_));
 sg13g2_nand2_1 _4421_ (.Y(_0636_),
    .A(_0273_),
    .B(_0635_));
 sg13g2_xnor2_1 _4422_ (.Y(_0637_),
    .A(_0205_),
    .B(_0596_));
 sg13g2_mux2_1 _4423_ (.A0(net140),
    .A1(_0307_),
    .S(_0637_),
    .X(_0638_));
 sg13g2_a21oi_1 _4424_ (.A1(net173),
    .A2(_0638_),
    .Y(_0639_),
    .B1(_0613_));
 sg13g2_nor4_1 _4425_ (.A(_0607_),
    .B(_0632_),
    .C(_0636_),
    .D(_0639_),
    .Y(_0640_));
 sg13g2_a221oi_1 _4426_ (.B2(_0629_),
    .C1(_0640_),
    .B1(_0628_),
    .A1(_0622_),
    .Y(_0641_),
    .A2(_0627_));
 sg13g2_nor2_1 _4427_ (.A(net139),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_nor3_1 _4428_ (.A(_0155_),
    .B(_1288_),
    .C(_0624_),
    .Y(_0643_));
 sg13g2_nand2_1 _4429_ (.Y(_0644_),
    .A(net117),
    .B(_0643_));
 sg13g2_o21ai_1 _4430_ (.B1(_0543_),
    .Y(_0645_),
    .A1(_0607_),
    .A2(_0644_));
 sg13g2_nor2_1 _4431_ (.A(_2676_),
    .B(_0635_),
    .Y(_0646_));
 sg13g2_a21oi_1 _4432_ (.A1(net81),
    .A2(_0643_),
    .Y(_0647_),
    .B1(_0646_));
 sg13g2_xnor2_1 _4433_ (.Y(_0648_),
    .A(_0630_),
    .B(_0594_));
 sg13g2_nor2_1 _4434_ (.A(net120),
    .B(_0648_),
    .Y(_0649_));
 sg13g2_xnor2_1 _4435_ (.Y(_0650_),
    .A(_2621_),
    .B(_0649_));
 sg13g2_nor3_1 _4436_ (.A(net114),
    .B(_0607_),
    .C(_0650_),
    .Y(_0651_));
 sg13g2_o21ai_1 _4437_ (.B1(_0651_),
    .Y(_0652_),
    .A1(_0607_),
    .A2(_0647_));
 sg13g2_nor2_1 _4438_ (.A(_0645_),
    .B(_0652_),
    .Y(_0653_));
 sg13g2_or4_1 _4439_ (.A(_0603_),
    .B(_0618_),
    .C(_0642_),
    .D(_0653_),
    .X(_0654_));
 sg13g2_nor2_1 _4440_ (.A(_0205_),
    .B(net131),
    .Y(_0655_));
 sg13g2_a22oi_1 _4441_ (.Y(_0656_),
    .B1(_0612_),
    .B2(net130),
    .A2(_0621_),
    .A1(_0655_));
 sg13g2_nand3_1 _4442_ (.B(_0625_),
    .C(_0621_),
    .A(net135),
    .Y(_0657_));
 sg13g2_o21ai_1 _4443_ (.B1(_0657_),
    .Y(_0658_),
    .A1(net145),
    .A2(_0656_));
 sg13g2_a21oi_1 _4444_ (.A1(_0372_),
    .A2(_0632_),
    .Y(_0659_),
    .B1(net117));
 sg13g2_nor2_1 _4445_ (.A(_0607_),
    .B(_0659_),
    .Y(_0660_));
 sg13g2_o21ai_1 _4446_ (.B1(_0660_),
    .Y(_0661_),
    .A1(net152),
    .A2(_0658_));
 sg13g2_a21oi_1 _4447_ (.A1(net143),
    .A2(_0613_),
    .Y(_0662_),
    .B1(_0632_));
 sg13g2_nor3_1 _4448_ (.A(net168),
    .B(_0543_),
    .C(_0662_),
    .Y(_0663_));
 sg13g2_inv_1 _4449_ (.Y(_0664_),
    .A(net199));
 sg13g2_a21o_1 _4450_ (.A2(_0275_),
    .A1(_0664_),
    .B1(_2612_),
    .X(_0665_));
 sg13g2_and4_1 _4451_ (.A(net168),
    .B(_0543_),
    .C(_0621_),
    .D(_0665_),
    .X(_0666_));
 sg13g2_o21ai_1 _4452_ (.B1(_0651_),
    .Y(_0667_),
    .A1(_0663_),
    .A2(_0666_));
 sg13g2_o21ai_1 _4453_ (.B1(net169),
    .Y(_0668_),
    .A1(net142),
    .A2(_0664_));
 sg13g2_a221oi_1 _4454_ (.B2(_0590_),
    .C1(_0668_),
    .B1(_0593_),
    .A1(net145),
    .Y(_0669_),
    .A2(_0624_));
 sg13g2_nand2b_1 _4455_ (.Y(_0670_),
    .B(_0669_),
    .A_N(_0429_));
 sg13g2_a21o_1 _4456_ (.A2(_0670_),
    .A1(net81),
    .B1(_0311_),
    .X(_0671_));
 sg13g2_a221oi_1 _4457_ (.B2(_0671_),
    .C1(_0603_),
    .B1(_0667_),
    .A1(net144),
    .Y(_0672_),
    .A2(_0661_));
 sg13g2_a21oi_1 _4458_ (.A1(_0504_),
    .A2(_0522_),
    .Y(_0673_),
    .B1(_2902_));
 sg13g2_nand3_1 _4459_ (.B(_0372_),
    .C(_0517_),
    .A(_0322_),
    .Y(_0674_));
 sg13g2_nand2b_1 _4460_ (.Y(_0675_),
    .B(_0674_),
    .A_N(_0673_));
 sg13g2_nand2_1 _4461_ (.Y(_0676_),
    .A(net161),
    .B(_0375_));
 sg13g2_and2_1 _4462_ (.A(_0518_),
    .B(_0676_),
    .X(_0677_));
 sg13g2_nor2_1 _4463_ (.A(net196),
    .B(_1463_),
    .Y(_0678_));
 sg13g2_o21ai_1 _4464_ (.B1(_0678_),
    .Y(_0679_),
    .A1(_0549_),
    .A2(_0677_));
 sg13g2_nor3_1 _4465_ (.A(_0371_),
    .B(_0543_),
    .C(_0514_),
    .Y(_0680_));
 sg13g2_a221oi_1 _4466_ (.B2(_0528_),
    .C1(_0680_),
    .B1(_0679_),
    .A1(_2989_),
    .Y(_0681_),
    .A2(_0675_));
 sg13g2_nand2_1 _4467_ (.Y(_0682_),
    .A(net115),
    .B(_0556_));
 sg13g2_mux2_1 _4468_ (.A0(_0535_),
    .A1(_0682_),
    .S(net152),
    .X(_0683_));
 sg13g2_nand4_1 _4469_ (.B(_0357_),
    .C(_0474_),
    .A(net176),
    .Y(_0684_),
    .D(net109));
 sg13g2_a21oi_1 _4470_ (.A1(_0683_),
    .A2(_0684_),
    .Y(_0685_),
    .B1(net114));
 sg13g2_and2_1 _4471_ (.A(net138),
    .B(_0568_),
    .X(_0686_));
 sg13g2_nor3_1 _4472_ (.A(net100),
    .B(_0521_),
    .C(_0686_),
    .Y(_0687_));
 sg13g2_nand2_1 _4473_ (.Y(_0688_),
    .A(net176),
    .B(_0474_));
 sg13g2_o21ai_1 _4474_ (.B1(_0528_),
    .Y(_0689_),
    .A1(_0504_),
    .A2(_0688_));
 sg13g2_nor3_1 _4475_ (.A(_0685_),
    .B(_0687_),
    .C(_0689_),
    .Y(_0690_));
 sg13g2_nand2_1 _4476_ (.Y(_0691_),
    .A(_2702_),
    .B(_0540_));
 sg13g2_nand3_1 _4477_ (.B(net181),
    .C(_2579_),
    .A(net198),
    .Y(_0692_));
 sg13g2_xnor2_1 _4478_ (.Y(_0693_),
    .A(_2855_),
    .B(_1496_));
 sg13g2_nand4_1 _4479_ (.B(_0691_),
    .C(_0692_),
    .A(_0575_),
    .Y(_0694_),
    .D(_0693_));
 sg13g2_nor2_1 _4480_ (.A(_2855_),
    .B(_1496_),
    .Y(_0695_));
 sg13g2_o21ai_1 _4481_ (.B1(_0521_),
    .Y(_0696_),
    .A1(net161),
    .A2(_0372_));
 sg13g2_nand2b_1 _4482_ (.Y(_0697_),
    .B(_0696_),
    .A_N(_0541_));
 sg13g2_a22oi_1 _4483_ (.Y(_0698_),
    .B1(_0695_),
    .B2(_0697_),
    .A2(_1529_),
    .A1(net195));
 sg13g2_nand4_1 _4484_ (.B(_0691_),
    .C(_0692_),
    .A(_1496_),
    .Y(_0699_),
    .D(_0696_));
 sg13g2_o21ai_1 _4485_ (.B1(_0699_),
    .Y(_0700_),
    .A1(_1518_),
    .A2(_1496_));
 sg13g2_nor2b_1 _4486_ (.A(_3011_),
    .B_N(net195),
    .Y(_0701_));
 sg13g2_a22oi_1 _4487_ (.Y(_0702_),
    .B1(_0700_),
    .B2(_0701_),
    .A2(_0698_),
    .A1(_3011_));
 sg13g2_nor4_1 _4488_ (.A(_0681_),
    .B(_0690_),
    .C(_0694_),
    .D(_0702_),
    .Y(_0703_));
 sg13g2_or2_1 _4489_ (.X(_0704_),
    .B(_0669_),
    .A(net100));
 sg13g2_nand3_1 _4490_ (.B(net168),
    .C(_0372_),
    .A(net100),
    .Y(_0705_));
 sg13g2_o21ai_1 _4491_ (.B1(_0705_),
    .Y(_0706_),
    .A1(net81),
    .A2(net168));
 sg13g2_a22oi_1 _4492_ (.Y(_0707_),
    .B1(_0706_),
    .B2(_2677_),
    .A2(_0704_),
    .A1(_2579_));
 sg13g2_nor3_1 _4493_ (.A(_2595_),
    .B(_0155_),
    .C(_0477_),
    .Y(_0708_));
 sg13g2_a221oi_1 _4494_ (.B2(_0622_),
    .C1(_0273_),
    .B1(_0708_),
    .A1(_0477_),
    .Y(_0709_),
    .A2(_0669_));
 sg13g2_nand2_1 _4495_ (.Y(_0710_),
    .A(_0322_),
    .B(_2903_));
 sg13g2_o21ai_1 _4496_ (.B1(_0710_),
    .Y(_0711_),
    .A1(net168),
    .A2(net175));
 sg13g2_o21ai_1 _4497_ (.B1(_0582_),
    .Y(_0712_),
    .A1(_2702_),
    .A2(_2903_));
 sg13g2_a22oi_1 _4498_ (.Y(_0713_),
    .B1(_0712_),
    .B2(_2677_),
    .A2(_0711_),
    .A1(_2695_));
 sg13g2_nor4_1 _4499_ (.A(_0600_),
    .B(_0707_),
    .C(_0709_),
    .D(_0713_),
    .Y(_0714_));
 sg13g2_nor3_1 _4500_ (.A(_0672_),
    .B(_0703_),
    .C(_0714_),
    .Y(_0715_));
 sg13g2_nand4_1 _4501_ (.B(_0581_),
    .C(_0654_),
    .A(_0498_),
    .Y(_0716_),
    .D(_0715_));
 sg13g2_nand2_1 _4502_ (.Y(_0717_),
    .A(_2740_),
    .B(_0204_));
 sg13g2_nand3b_1 _4503_ (.B(_0664_),
    .C(_2747_),
    .Y(_0718_),
    .A_N(_2748_));
 sg13g2_a22oi_1 _4504_ (.Y(_0719_),
    .B1(_0717_),
    .B2(_0718_),
    .A2(_0135_),
    .A1(_0133_));
 sg13g2_nand3_1 _4505_ (.B(_2833_),
    .C(_0719_),
    .A(_2863_),
    .Y(_0720_));
 sg13g2_nand3_1 _4506_ (.B(net154),
    .C(_2831_),
    .A(_2775_),
    .Y(_0721_));
 sg13g2_a21oi_2 _4507_ (.B1(_0721_),
    .Y(_0722_),
    .A2(_0135_),
    .A1(_0133_));
 sg13g2_nand2_1 _4508_ (.Y(_0723_),
    .A(net101),
    .B(_0722_));
 sg13g2_a21oi_1 _4509_ (.A1(_0720_),
    .A2(_0723_),
    .Y(_0724_),
    .B1(_0169_));
 sg13g2_nand2_1 _4510_ (.Y(_0725_),
    .A(net113),
    .B(_0109_));
 sg13g2_nor2_1 _4511_ (.A(_1332_),
    .B(_2839_),
    .Y(_0726_));
 sg13g2_nor3_1 _4512_ (.A(net186),
    .B(_2965_),
    .C(_0275_),
    .Y(_0727_));
 sg13g2_o21ai_1 _4513_ (.B1(_0664_),
    .Y(_0728_),
    .A1(_0726_),
    .A2(_0727_));
 sg13g2_a21oi_1 _4514_ (.A1(_2609_),
    .A2(_0664_),
    .Y(_0729_),
    .B1(_2740_));
 sg13g2_nand3_1 _4515_ (.B(_2747_),
    .C(_2745_),
    .A(net133),
    .Y(_0730_));
 sg13g2_o21ai_1 _4516_ (.B1(_0730_),
    .Y(_0731_),
    .A1(net177),
    .A2(_0729_));
 sg13g2_nand3_1 _4517_ (.B(_0728_),
    .C(_0731_),
    .A(_0136_),
    .Y(_0732_));
 sg13g2_buf_1 _4518_ (.A(_0732_),
    .X(_0733_));
 sg13g2_nor3_1 _4519_ (.A(net86),
    .B(_0725_),
    .C(_0733_),
    .Y(_0734_));
 sg13g2_nor3_1 _4520_ (.A(_0222_),
    .B(_0724_),
    .C(_0734_),
    .Y(_0735_));
 sg13g2_nor2_1 _4521_ (.A(_2836_),
    .B(_2822_),
    .Y(_0736_));
 sg13g2_nand2b_1 _4522_ (.Y(_0737_),
    .B(_0136_),
    .A_N(_0721_));
 sg13g2_buf_1 _4523_ (.A(_0737_),
    .X(_0738_));
 sg13g2_buf_1 _4524_ (.A(_0719_),
    .X(_0739_));
 sg13g2_nand2_1 _4525_ (.Y(_0740_),
    .A(_2833_),
    .B(net96));
 sg13g2_nor2_1 _4526_ (.A(_2814_),
    .B(_0113_),
    .Y(_0741_));
 sg13g2_a22oi_1 _4527_ (.Y(_0742_),
    .B1(_0219_),
    .B2(net158),
    .A2(_2997_),
    .A1(_2816_));
 sg13g2_xnor2_1 _4528_ (.Y(_0743_),
    .A(_2710_),
    .B(_0742_));
 sg13g2_o21ai_1 _4529_ (.B1(_0743_),
    .Y(_0744_),
    .A1(_0142_),
    .A2(_0741_));
 sg13g2_a221oi_1 _4530_ (.B2(_0193_),
    .C1(_0744_),
    .B1(_0740_),
    .A1(_0736_),
    .Y(_0745_),
    .A2(_0738_));
 sg13g2_and2_1 _4531_ (.A(net200),
    .B(_2728_),
    .X(_0746_));
 sg13g2_o21ai_1 _4532_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net162),
    .A2(_2734_));
 sg13g2_nand4_1 _4533_ (.B(_0547_),
    .C(_2727_),
    .A(_2725_),
    .Y(_0748_),
    .D(_2735_));
 sg13g2_a22oi_1 _4534_ (.Y(_0749_),
    .B1(_0747_),
    .B2(_0748_),
    .A2(_2750_),
    .A1(_2746_));
 sg13g2_buf_1 _4535_ (.A(_0749_),
    .X(_0750_));
 sg13g2_nand2b_1 _4536_ (.Y(_0751_),
    .B(_0750_),
    .A_N(_2870_));
 sg13g2_a21oi_1 _4537_ (.A1(_0187_),
    .A2(_0722_),
    .Y(_0752_),
    .B1(net98));
 sg13g2_nand2_1 _4538_ (.Y(_0753_),
    .A(_0751_),
    .B(_0752_));
 sg13g2_nor2_1 _4539_ (.A(_2820_),
    .B(_0742_),
    .Y(_0754_));
 sg13g2_nor2_2 _4540_ (.A(_3015_),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_a21oi_1 _4541_ (.A1(_0745_),
    .A2(_0753_),
    .Y(_0756_),
    .B1(_0755_));
 sg13g2_o21ai_1 _4542_ (.B1(_0756_),
    .Y(_0757_),
    .A1(_3016_),
    .A2(_0735_));
 sg13g2_nand2_1 _4543_ (.Y(_0758_),
    .A(_2833_),
    .B(_0750_));
 sg13g2_and2_1 _4544_ (.A(_0733_),
    .B(_0758_),
    .X(_0759_));
 sg13g2_nand2_1 _4545_ (.Y(_0760_),
    .A(_2842_),
    .B(net96));
 sg13g2_a221oi_1 _4546_ (.B2(_2841_),
    .C1(net101),
    .B1(net96),
    .A1(_0136_),
    .Y(_0761_),
    .A2(_0175_));
 sg13g2_a21oi_1 _4547_ (.A1(net86),
    .A2(_0760_),
    .Y(_0762_),
    .B1(_0761_));
 sg13g2_nor3_1 _4548_ (.A(_0169_),
    .B(_0759_),
    .C(_0762_),
    .Y(_0763_));
 sg13g2_nand3_1 _4549_ (.B(_0128_),
    .C(_0750_),
    .A(_2863_),
    .Y(_0764_));
 sg13g2_nand3_1 _4550_ (.B(_0738_),
    .C(_0764_),
    .A(_0151_),
    .Y(_0765_));
 sg13g2_a21oi_1 _4551_ (.A1(_0193_),
    .A2(_0759_),
    .Y(_0766_),
    .B1(_0765_));
 sg13g2_a21o_1 _4552_ (.A2(_0720_),
    .A1(_0738_),
    .B1(_0736_),
    .X(_0767_));
 sg13g2_and3_1 _4553_ (.X(_0768_),
    .A(_0169_),
    .B(_0725_),
    .C(_0767_));
 sg13g2_nor4_1 _4554_ (.A(_0743_),
    .B(_0763_),
    .C(_0766_),
    .D(_0768_),
    .Y(_0769_));
 sg13g2_a21oi_1 _4555_ (.A1(_2963_),
    .A2(_2966_),
    .Y(_0770_),
    .B1(net85));
 sg13g2_nand3_1 _4556_ (.B(_2850_),
    .C(_0739_),
    .A(net156),
    .Y(_0771_));
 sg13g2_o21ai_1 _4557_ (.B1(_0771_),
    .Y(_0772_),
    .A1(net156),
    .A2(_0733_));
 sg13g2_a22oi_1 _4558_ (.Y(_0773_),
    .B1(_0772_),
    .B2(_2865_),
    .A2(_0770_),
    .A1(net96));
 sg13g2_nor2_1 _4559_ (.A(_0111_),
    .B(_0754_),
    .Y(_0774_));
 sg13g2_nand4_1 _4560_ (.B(_2863_),
    .C(_0140_),
    .A(net98),
    .Y(_0775_),
    .D(_0722_));
 sg13g2_nor2_1 _4561_ (.A(net112),
    .B(_0222_),
    .Y(_0776_));
 sg13g2_a21oi_1 _4562_ (.A1(net112),
    .A2(_0775_),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_nand2_1 _4563_ (.Y(_0778_),
    .A(_2850_),
    .B(net96));
 sg13g2_nand2_1 _4564_ (.Y(_0779_),
    .A(_0738_),
    .B(_0778_));
 sg13g2_nor3_1 _4565_ (.A(net98),
    .B(_0140_),
    .C(_0743_),
    .Y(_0780_));
 sg13g2_nor2_1 _4566_ (.A(_2706_),
    .B(_0754_),
    .Y(_0781_));
 sg13g2_a221oi_1 _4567_ (.B2(_0780_),
    .C1(_0781_),
    .B1(_0779_),
    .A1(net84),
    .Y(_0782_),
    .A2(_0777_));
 sg13g2_o21ai_1 _4568_ (.B1(_0782_),
    .Y(_0783_),
    .A1(_0773_),
    .A2(_0774_));
 sg13g2_o21ai_1 _4569_ (.B1(_0783_),
    .Y(_0784_),
    .A1(_0757_),
    .A2(_0769_));
 sg13g2_nor2_1 _4570_ (.A(_2814_),
    .B(_2828_),
    .Y(_0785_));
 sg13g2_and2_1 _4571_ (.A(_2814_),
    .B(_2997_),
    .X(_0786_));
 sg13g2_nand2_1 _4572_ (.Y(_0787_),
    .A(net184),
    .B(net198));
 sg13g2_a22oi_1 _4573_ (.Y(_0788_),
    .B1(_2960_),
    .B2(_2714_),
    .A2(_3034_),
    .A1(_2719_));
 sg13g2_o21ai_1 _4574_ (.B1(_0788_),
    .Y(_0789_),
    .A1(_2959_),
    .A2(_0787_));
 sg13g2_nor3_1 _4575_ (.A(_0785_),
    .B(_0786_),
    .C(_0789_),
    .Y(_0790_));
 sg13g2_a221oi_1 _4576_ (.B2(_0758_),
    .C1(_0790_),
    .B1(_0733_),
    .A1(_0187_),
    .Y(_0791_),
    .A2(_0722_));
 sg13g2_nor2b_1 _4577_ (.A(_0791_),
    .B_N(_0776_),
    .Y(_0792_));
 sg13g2_nor4_1 _4578_ (.A(_2710_),
    .B(net98),
    .C(_0113_),
    .D(_0733_),
    .Y(_0793_));
 sg13g2_a221oi_1 _4579_ (.B2(_0128_),
    .C1(net86),
    .B1(_0750_),
    .A1(_2841_),
    .Y(_0794_),
    .A2(net96));
 sg13g2_nand2_1 _4580_ (.Y(_0795_),
    .A(_0136_),
    .B(_0175_));
 sg13g2_and4_1 _4581_ (.A(net101),
    .B(_0751_),
    .C(_0760_),
    .D(_0795_),
    .X(_0796_));
 sg13g2_o21ai_1 _4582_ (.B1(net83),
    .Y(_0797_),
    .A1(_0794_),
    .A2(_0796_));
 sg13g2_o21ai_1 _4583_ (.B1(_0797_),
    .Y(_0798_),
    .A1(_0792_),
    .A2(_0793_));
 sg13g2_and2_1 _4584_ (.A(_3010_),
    .B(_0755_),
    .X(_0799_));
 sg13g2_nor2_1 _4585_ (.A(_3010_),
    .B(_0755_),
    .Y(_0800_));
 sg13g2_a21o_1 _4586_ (.A2(_0799_),
    .A1(_0798_),
    .B1(_0800_),
    .X(_0801_));
 sg13g2_o21ai_1 _4587_ (.B1(_0738_),
    .Y(_0802_),
    .A1(net86),
    .A2(_0778_));
 sg13g2_nand2_1 _4588_ (.Y(_0803_),
    .A(net83),
    .B(_0802_));
 sg13g2_nand2_1 _4589_ (.Y(_0804_),
    .A(_2858_),
    .B(_0755_));
 sg13g2_nand3_1 _4590_ (.B(_2829_),
    .C(_0779_),
    .A(net98),
    .Y(_0805_));
 sg13g2_nand2_1 _4591_ (.Y(_0806_),
    .A(_0169_),
    .B(_0725_));
 sg13g2_nand4_1 _4592_ (.B(_2848_),
    .C(_0739_),
    .A(_2864_),
    .Y(_0807_),
    .D(_0806_));
 sg13g2_a21oi_1 _4593_ (.A1(_0805_),
    .A2(_0807_),
    .Y(_0808_),
    .B1(_0109_));
 sg13g2_nor2_1 _4594_ (.A(_2831_),
    .B(_0169_),
    .Y(_0809_));
 sg13g2_a21oi_1 _4595_ (.A1(net96),
    .A2(_0809_),
    .Y(_0810_),
    .B1(_0151_));
 sg13g2_nor3_1 _4596_ (.A(net86),
    .B(_0733_),
    .C(_0810_),
    .Y(_0811_));
 sg13g2_nor4_1 _4597_ (.A(_0743_),
    .B(_0804_),
    .C(_0808_),
    .D(_0811_),
    .Y(_0812_));
 sg13g2_nand2_1 _4598_ (.Y(_0813_),
    .A(_2863_),
    .B(_2965_));
 sg13g2_nor2_1 _4599_ (.A(net193),
    .B(_2774_),
    .Y(_0814_));
 sg13g2_nand2_1 _4600_ (.Y(_0815_),
    .A(_0814_),
    .B(net101));
 sg13g2_a21oi_1 _4601_ (.A1(_0813_),
    .A2(_0815_),
    .Y(_0816_),
    .B1(_1332_));
 sg13g2_xnor2_1 _4602_ (.Y(_0817_),
    .A(net130),
    .B(net101));
 sg13g2_nor3_1 _4603_ (.A(_2555_),
    .B(_0165_),
    .C(_0817_),
    .Y(_0818_));
 sg13g2_o21ai_1 _4604_ (.B1(net96),
    .Y(_0819_),
    .A1(_0816_),
    .A2(_0818_));
 sg13g2_and3_1 _4605_ (.X(_0820_),
    .A(_0136_),
    .B(_0728_),
    .C(_0731_));
 sg13g2_a21oi_1 _4606_ (.A1(net86),
    .A2(_0820_),
    .Y(_0821_),
    .B1(_0110_));
 sg13g2_a221oi_1 _4607_ (.B2(_0222_),
    .C1(_0821_),
    .B1(_0819_),
    .A1(_0767_),
    .Y(_0822_),
    .A2(_0806_));
 sg13g2_nand3_1 _4608_ (.B(net84),
    .C(_0743_),
    .A(_2858_),
    .Y(_0823_));
 sg13g2_nor2_1 _4609_ (.A(_0820_),
    .B(_0750_),
    .Y(_0824_));
 sg13g2_nor2_1 _4610_ (.A(_2858_),
    .B(_0755_),
    .Y(_0825_));
 sg13g2_nor4_1 _4611_ (.A(net5),
    .B(_3013_),
    .C(_0824_),
    .D(_0825_),
    .Y(_0826_));
 sg13g2_o21ai_1 _4612_ (.B1(_0826_),
    .Y(_0827_),
    .A1(_0822_),
    .A2(_0823_));
 sg13g2_a221oi_1 _4613_ (.B2(_0812_),
    .C1(_0827_),
    .B1(_0803_),
    .A1(_0784_),
    .Y(_0828_),
    .A2(_0801_));
 sg13g2_a21oi_1 _4614_ (.A1(_0247_),
    .A2(_0716_),
    .Y(_0829_),
    .B1(_0828_));
 sg13g2_nand3_1 _4615_ (.B(_0246_),
    .C(_0829_),
    .A(_0108_),
    .Y(_0830_));
 sg13g2_buf_2 _4616_ (.A(_0830_),
    .X(_0831_));
 sg13g2_nor2_1 _4617_ (.A(net240),
    .B(_2547_),
    .Y(_0832_));
 sg13g2_nand2_1 _4618_ (.Y(_0833_),
    .A(_1386_),
    .B(net233));
 sg13g2_nand3_1 _4619_ (.B(net234),
    .C(net233),
    .A(net218),
    .Y(_0834_));
 sg13g2_nand3_1 _4620_ (.B(net218),
    .C(net234),
    .A(_1386_),
    .Y(_0835_));
 sg13g2_nand4_1 _4621_ (.B(_0833_),
    .C(_0834_),
    .A(_0311_),
    .Y(_0836_),
    .D(_0835_));
 sg13g2_nand3_1 _4622_ (.B(_0834_),
    .C(_0835_),
    .A(_0833_),
    .Y(_0837_));
 sg13g2_and2_1 _4623_ (.A(net240),
    .B(_2547_),
    .X(_0838_));
 sg13g2_a221oi_1 _4624_ (.B2(net241),
    .C1(_0838_),
    .B1(_0837_),
    .A1(net232),
    .Y(_0839_),
    .A2(_0836_));
 sg13g2_or2_1 _4625_ (.X(_0840_),
    .B(_0839_),
    .A(_0832_));
 sg13g2_buf_2 _4626_ (.A(_0840_),
    .X(_0841_));
 sg13g2_nand2_1 _4627_ (.Y(_0842_),
    .A(_2567_),
    .B(net235));
 sg13g2_a21oi_1 _4628_ (.A1(_2576_),
    .A2(net236),
    .Y(_0843_),
    .B1(_2525_));
 sg13g2_a21oi_1 _4629_ (.A1(_2567_),
    .A2(net235),
    .Y(_0844_),
    .B1(\graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ));
 sg13g2_nand3_1 _4630_ (.B(_2525_),
    .C(net236),
    .A(_2576_),
    .Y(_0845_));
 sg13g2_nor2_1 _4631_ (.A(_2567_),
    .B(net235),
    .Y(_0846_));
 sg13g2_a221oi_1 _4632_ (.B2(_0845_),
    .C1(_0846_),
    .B1(_0844_),
    .A1(_0842_),
    .Y(_0847_),
    .A2(_0843_));
 sg13g2_buf_2 _4633_ (.A(_0847_),
    .X(_0848_));
 sg13g2_and2_1 _4634_ (.A(_2570_),
    .B(_2532_),
    .X(_0849_));
 sg13g2_buf_1 _4635_ (.A(_0849_),
    .X(_0850_));
 sg13g2_or2_1 _4636_ (.X(_0851_),
    .B(_2532_),
    .A(_2570_));
 sg13g2_buf_1 _4637_ (.A(_0851_),
    .X(_0852_));
 sg13g2_o21ai_1 _4638_ (.B1(_0852_),
    .Y(_0853_),
    .A1(_0848_),
    .A2(_0850_));
 sg13g2_buf_1 _4639_ (.A(_0853_),
    .X(_0854_));
 sg13g2_xnor2_1 _4640_ (.Y(_0855_),
    .A(_1386_),
    .B(net233));
 sg13g2_xnor2_1 _4641_ (.Y(_0856_),
    .A(net218),
    .B(net234));
 sg13g2_buf_2 _4642_ (.A(_0856_),
    .X(_0857_));
 sg13g2_xnor2_1 _4643_ (.Y(_0858_),
    .A(_1364_),
    .B(net232));
 sg13g2_buf_1 _4644_ (.A(_0858_),
    .X(_0859_));
 sg13g2_nor4_2 _4645_ (.A(_0832_),
    .B(_0855_),
    .C(_0857_),
    .Y(_0860_),
    .D(net172));
 sg13g2_nand2b_1 _4646_ (.Y(_0861_),
    .B(_0860_),
    .A_N(net108));
 sg13g2_buf_2 _4647_ (.A(_0861_),
    .X(_0862_));
 sg13g2_xor2_1 _4648_ (.B(\graphics_engine_1.ctr[8] ),
    .A(_1507_),
    .X(_0863_));
 sg13g2_a21oi_2 _4649_ (.B1(_0863_),
    .Y(_0864_),
    .A2(_0862_),
    .A1(_0841_));
 sg13g2_buf_8 _4650_ (.A(_0864_),
    .X(_0865_));
 sg13g2_xnor2_1 _4651_ (.Y(_0866_),
    .A(_1507_),
    .B(\graphics_engine_1.ctr[8] ));
 sg13g2_buf_2 _4652_ (.A(_0866_),
    .X(_0867_));
 sg13g2_nor2_1 _4653_ (.A(_0832_),
    .B(_0839_),
    .Y(_0868_));
 sg13g2_buf_1 _4654_ (.A(_0868_),
    .X(_0869_));
 sg13g2_nor2b_1 _4655_ (.A(net108),
    .B_N(_0860_),
    .Y(_0870_));
 sg13g2_buf_2 _4656_ (.A(_0870_),
    .X(_0871_));
 sg13g2_nor3_1 _4657_ (.A(_0867_),
    .B(net95),
    .C(_0871_),
    .Y(_0872_));
 sg13g2_buf_1 _4658_ (.A(_0872_),
    .X(_0873_));
 sg13g2_nor2_2 _4659_ (.A(net53),
    .B(net52),
    .Y(_0874_));
 sg13g2_nand2_1 _4660_ (.Y(_0875_),
    .A(net119),
    .B(net134));
 sg13g2_buf_1 _4661_ (.A(_2769_),
    .X(_0876_));
 sg13g2_nand3_1 _4662_ (.B(net171),
    .C(_0874_),
    .A(net133),
    .Y(_0877_));
 sg13g2_o21ai_1 _4663_ (.B1(_0877_),
    .Y(_0878_),
    .A1(_0874_),
    .A2(_0875_));
 sg13g2_nor2_1 _4664_ (.A(net132),
    .B(net110),
    .Y(_0879_));
 sg13g2_buf_2 _4665_ (.A(_0879_),
    .X(_0880_));
 sg13g2_o21ai_1 _4666_ (.B1(_0867_),
    .Y(_0881_),
    .A1(net95),
    .A2(_0871_));
 sg13g2_buf_2 _4667_ (.A(_0881_),
    .X(_0882_));
 sg13g2_nand3_1 _4668_ (.B(_0841_),
    .C(_0862_),
    .A(_0863_),
    .Y(_0883_));
 sg13g2_buf_2 _4669_ (.A(_0883_),
    .X(_0884_));
 sg13g2_nand2_1 _4670_ (.Y(_0885_),
    .A(net164),
    .B(_0194_));
 sg13g2_nand2_1 _4671_ (.Y(_0886_),
    .A(_2760_),
    .B(_0885_));
 sg13g2_buf_1 _4672_ (.A(_0886_),
    .X(_0887_));
 sg13g2_buf_1 _4673_ (.A(net97),
    .X(_0888_));
 sg13g2_a221oi_1 _4674_ (.B2(net151),
    .C1(net80),
    .B1(net94),
    .A1(_0882_),
    .Y(_0889_),
    .A2(_0884_));
 sg13g2_xnor2_1 _4675_ (.Y(_0890_),
    .A(_0880_),
    .B(_0889_));
 sg13g2_nand2_2 _4676_ (.Y(_0891_),
    .A(_0882_),
    .B(_0884_));
 sg13g2_xnor2_1 _4677_ (.Y(_0892_),
    .A(_2769_),
    .B(_0867_));
 sg13g2_o21ai_1 _4678_ (.B1(_0892_),
    .Y(_0893_),
    .A1(net95),
    .A2(_0871_));
 sg13g2_buf_1 _4679_ (.A(_0893_),
    .X(_0894_));
 sg13g2_nand3b_1 _4680_ (.B(_0862_),
    .C(_0841_),
    .Y(_0895_),
    .A_N(_0892_));
 sg13g2_buf_1 _4681_ (.A(_0895_),
    .X(_0896_));
 sg13g2_nand2_1 _4682_ (.Y(_0897_),
    .A(_0894_),
    .B(_0896_));
 sg13g2_buf_2 _4683_ (.A(_0897_),
    .X(_0898_));
 sg13g2_nor3_1 _4684_ (.A(net118),
    .B(net53),
    .C(net52),
    .Y(_0899_));
 sg13g2_a221oi_1 _4685_ (.B2(net119),
    .C1(_0899_),
    .B1(_0898_),
    .A1(_0318_),
    .Y(_0900_),
    .A2(_0891_));
 sg13g2_nand2b_1 _4686_ (.Y(_0901_),
    .B(_0900_),
    .A_N(_0890_));
 sg13g2_nand2_1 _4687_ (.Y(_0902_),
    .A(net151),
    .B(net171));
 sg13g2_nor3_1 _4688_ (.A(net53),
    .B(net52),
    .C(_0902_),
    .Y(_0903_));
 sg13g2_nand2_1 _4689_ (.Y(_0904_),
    .A(net118),
    .B(net134));
 sg13g2_a21oi_1 _4690_ (.A1(_0902_),
    .A2(_0904_),
    .Y(_0905_),
    .B1(net119));
 sg13g2_nor2_1 _4691_ (.A(_0903_),
    .B(_0905_),
    .Y(_0906_));
 sg13g2_a21oi_1 _4692_ (.A1(_0890_),
    .A2(_0906_),
    .Y(_0907_),
    .B1(net120));
 sg13g2_a22oi_1 _4693_ (.Y(_0908_),
    .B1(_0901_),
    .B2(_0907_),
    .A2(_0878_),
    .A1(net151));
 sg13g2_nand2_1 _4694_ (.Y(_0909_),
    .A(net133),
    .B(_0898_));
 sg13g2_nand2_1 _4695_ (.Y(_0910_),
    .A(net119),
    .B(net118));
 sg13g2_mux2_1 _4696_ (.A0(net118),
    .A1(_0910_),
    .S(_0874_),
    .X(_0911_));
 sg13g2_a21o_1 _4697_ (.A2(_0911_),
    .A1(_0909_),
    .B1(_0890_),
    .X(_0912_));
 sg13g2_nor2b_1 _4698_ (.A(_1134_),
    .B_N(_0028_),
    .Y(_0913_));
 sg13g2_and3_1 _4699_ (.X(_0914_),
    .A(net119),
    .B(_0902_),
    .C(_0904_));
 sg13g2_a22oi_1 _4700_ (.Y(_0915_),
    .B1(_0914_),
    .B2(_0890_),
    .A2(_0913_),
    .A1(_0891_));
 sg13g2_a21o_1 _4701_ (.A2(_0915_),
    .A1(_0912_),
    .B1(net145),
    .X(_0916_));
 sg13g2_xnor2_1 _4702_ (.Y(_0917_),
    .A(net222),
    .B(net225));
 sg13g2_buf_1 _4703_ (.A(_0917_),
    .X(_0918_));
 sg13g2_nor3_1 _4704_ (.A(net182),
    .B(_0867_),
    .C(net150),
    .Y(_0919_));
 sg13g2_nand2b_1 _4705_ (.Y(_0920_),
    .B(_0919_),
    .A_N(_0860_));
 sg13g2_nand2_1 _4706_ (.Y(_0921_),
    .A(net108),
    .B(_0919_));
 sg13g2_a21o_1 _4707_ (.A2(_0921_),
    .A1(_0920_),
    .B1(net95),
    .X(_0922_));
 sg13g2_nor3_1 _4708_ (.A(net182),
    .B(_0863_),
    .C(net150),
    .Y(_0923_));
 sg13g2_nand2_1 _4709_ (.Y(_0924_),
    .A(_0860_),
    .B(_0923_));
 sg13g2_o21ai_1 _4710_ (.B1(net97),
    .Y(_0925_),
    .A1(net108),
    .A2(_0924_));
 sg13g2_a21oi_1 _4711_ (.A1(net95),
    .A2(_0923_),
    .Y(_0926_),
    .B1(_0925_));
 sg13g2_nor2b_1 _4712_ (.A(net97),
    .B_N(_0919_),
    .Y(_0927_));
 sg13g2_nor2_1 _4713_ (.A(net95),
    .B(_0871_),
    .Y(_0928_));
 sg13g2_a21oi_1 _4714_ (.A1(net179),
    .A2(_0257_),
    .Y(_0929_),
    .B1(_0547_));
 sg13g2_a21o_1 _4715_ (.A2(_0257_),
    .A1(_0255_),
    .B1(_0929_),
    .X(_0930_));
 sg13g2_buf_1 _4716_ (.A(_0930_),
    .X(_0931_));
 sg13g2_nand2_1 _4717_ (.Y(_0932_),
    .A(_0931_),
    .B(_0923_));
 sg13g2_a21oi_1 _4718_ (.A1(_0841_),
    .A2(_0862_),
    .Y(_0933_),
    .B1(_0932_));
 sg13g2_a221oi_1 _4719_ (.B2(_0928_),
    .C1(_0933_),
    .B1(_0927_),
    .A1(_0922_),
    .Y(_0934_),
    .A2(_0926_));
 sg13g2_buf_2 _4720_ (.A(_0934_),
    .X(_0935_));
 sg13g2_buf_1 _4721_ (.A(net150),
    .X(_0936_));
 sg13g2_xnor2_1 _4722_ (.Y(_0937_),
    .A(net182),
    .B(_2768_));
 sg13g2_nor2_1 _4723_ (.A(net93),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_o21ai_1 _4724_ (.B1(_0938_),
    .Y(_0939_),
    .A1(_0864_),
    .A2(_0872_));
 sg13g2_buf_1 _4725_ (.A(_0939_),
    .X(_0940_));
 sg13g2_nand3_1 _4726_ (.B(_0882_),
    .C(_0884_),
    .A(net93),
    .Y(_0941_));
 sg13g2_nand3_1 _4727_ (.B(_0940_),
    .C(_0941_),
    .A(net171),
    .Y(_0942_));
 sg13g2_xnor2_1 _4728_ (.Y(_0943_),
    .A(net180),
    .B(_0249_));
 sg13g2_nand4_1 _4729_ (.B(_0882_),
    .C(_0884_),
    .A(net80),
    .Y(_0944_),
    .D(_0943_));
 sg13g2_buf_1 _4730_ (.A(_0944_),
    .X(_0945_));
 sg13g2_o21ai_1 _4731_ (.B1(net93),
    .Y(_0946_),
    .A1(net53),
    .A2(net52));
 sg13g2_nand3_1 _4732_ (.B(_0945_),
    .C(_0946_),
    .A(net134),
    .Y(_0947_));
 sg13g2_nand4_1 _4733_ (.B(_0890_),
    .C(_0942_),
    .A(net129),
    .Y(_0948_),
    .D(_0947_));
 sg13g2_nand3_1 _4734_ (.B(_0888_),
    .C(net94),
    .A(net134),
    .Y(_0949_));
 sg13g2_nand4_1 _4735_ (.B(net93),
    .C(_0882_),
    .A(net171),
    .Y(_0950_),
    .D(_0884_));
 sg13g2_o21ai_1 _4736_ (.B1(_0950_),
    .Y(_0951_),
    .A1(_0874_),
    .A2(_0949_));
 sg13g2_nand3_1 _4737_ (.B(_0890_),
    .C(_0951_),
    .A(net151),
    .Y(_0952_));
 sg13g2_nor2_1 _4738_ (.A(_0880_),
    .B(_0935_),
    .Y(_0953_));
 sg13g2_nand2_1 _4739_ (.Y(_0954_),
    .A(_0867_),
    .B(_0937_));
 sg13g2_a21oi_1 _4740_ (.A1(_0841_),
    .A2(_0862_),
    .Y(_0955_),
    .B1(_0954_));
 sg13g2_xnor2_1 _4741_ (.Y(_0956_),
    .A(net180),
    .B(_2768_));
 sg13g2_nor4_1 _4742_ (.A(_0867_),
    .B(net95),
    .C(_0871_),
    .D(_0956_),
    .Y(_0957_));
 sg13g2_xnor2_1 _4743_ (.Y(_0958_),
    .A(net182),
    .B(_0249_));
 sg13g2_nand2_1 _4744_ (.Y(_0959_),
    .A(_0863_),
    .B(_0958_));
 sg13g2_a21oi_1 _4745_ (.A1(_0841_),
    .A2(_0862_),
    .Y(_0960_),
    .B1(_0959_));
 sg13g2_nor4_1 _4746_ (.A(_0863_),
    .B(net95),
    .C(_0871_),
    .D(_0943_),
    .Y(_0961_));
 sg13g2_nor4_1 _4747_ (.A(_0955_),
    .B(_0957_),
    .C(_0960_),
    .D(_0961_),
    .Y(_0962_));
 sg13g2_buf_2 _4748_ (.A(_0962_),
    .X(_0963_));
 sg13g2_o21ai_1 _4749_ (.B1(_0963_),
    .Y(_0964_),
    .A1(net94),
    .A2(_0898_));
 sg13g2_nor2_1 _4750_ (.A(net162),
    .B(net150),
    .Y(_0965_));
 sg13g2_o21ai_1 _4751_ (.B1(_0965_),
    .Y(_0966_),
    .A1(_0864_),
    .A2(_0872_));
 sg13g2_buf_1 _4752_ (.A(_0966_),
    .X(_0967_));
 sg13g2_or2_1 _4753_ (.X(_0968_),
    .B(_0254_),
    .A(_0253_));
 sg13g2_buf_1 _4754_ (.A(_0968_),
    .X(_0969_));
 sg13g2_nor2_1 _4755_ (.A(_2769_),
    .B(_0958_),
    .Y(_0970_));
 sg13g2_nand4_1 _4756_ (.B(_0882_),
    .C(_0884_),
    .A(net92),
    .Y(_0971_),
    .D(_0970_));
 sg13g2_o21ai_1 _4757_ (.B1(_0261_),
    .Y(_0972_),
    .A1(net132),
    .A2(net110));
 sg13g2_buf_1 _4758_ (.A(_0972_),
    .X(_0973_));
 sg13g2_nand2_1 _4759_ (.Y(_0974_),
    .A(_2769_),
    .B(_0956_));
 sg13g2_a21oi_1 _4760_ (.A1(net82),
    .A2(_0973_),
    .Y(_0975_),
    .B1(_0974_));
 sg13g2_o21ai_1 _4761_ (.B1(_0975_),
    .Y(_0976_),
    .A1(net53),
    .A2(net52));
 sg13g2_a22oi_1 _4762_ (.Y(_0977_),
    .B1(_0971_),
    .B2(_0976_),
    .A2(_0967_),
    .A1(net80));
 sg13g2_nand2_1 _4763_ (.Y(_0978_),
    .A(net92),
    .B(net94));
 sg13g2_a21o_1 _4764_ (.A2(_0896_),
    .A1(_0894_),
    .B1(_0978_),
    .X(_0979_));
 sg13g2_buf_1 _4765_ (.A(_0979_),
    .X(_0980_));
 sg13g2_a21oi_2 _4766_ (.B1(_0980_),
    .Y(_0981_),
    .A2(_0945_),
    .A1(_0940_));
 sg13g2_a221oi_1 _4767_ (.B2(net129),
    .C1(_0981_),
    .B1(_0977_),
    .A1(_0953_),
    .Y(_0982_),
    .A2(_0964_));
 sg13g2_nand4_1 _4768_ (.B(_0948_),
    .C(_0952_),
    .A(_0935_),
    .Y(_0983_),
    .D(_0982_));
 sg13g2_a21oi_2 _4769_ (.B1(_0983_),
    .Y(_0984_),
    .A2(_0916_),
    .A1(_0908_));
 sg13g2_or2_1 _4770_ (.X(_0985_),
    .B(_2576_),
    .A(net231));
 sg13g2_nor3_1 _4771_ (.A(net153),
    .B(_0252_),
    .C(net150),
    .Y(_0986_));
 sg13g2_nand4_1 _4772_ (.B(_0884_),
    .C(_0943_),
    .A(_0882_),
    .Y(_0987_),
    .D(_0986_));
 sg13g2_buf_1 _4773_ (.A(_0987_),
    .X(_0988_));
 sg13g2_nand3_1 _4774_ (.B(net153),
    .C(net94),
    .A(net118),
    .Y(_0989_));
 sg13g2_a21oi_1 _4775_ (.A1(net82),
    .A2(_0973_),
    .Y(_0990_),
    .B1(_0989_));
 sg13g2_o21ai_1 _4776_ (.B1(_0990_),
    .Y(_0991_),
    .A1(net53),
    .A2(net52));
 sg13g2_buf_1 _4777_ (.A(_0991_),
    .X(_0992_));
 sg13g2_nand2_2 _4778_ (.Y(_0993_),
    .A(_0988_),
    .B(_0992_));
 sg13g2_nor2_1 _4779_ (.A(_0935_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_nand4_1 _4780_ (.B(_0952_),
    .C(_0982_),
    .A(_0948_),
    .Y(_0995_),
    .D(_0994_));
 sg13g2_nand3b_1 _4781_ (.B(_0985_),
    .C(_0995_),
    .Y(_0996_),
    .A_N(net4));
 sg13g2_or2_1 _4782_ (.X(_0997_),
    .B(_0996_),
    .A(_0984_));
 sg13g2_buf_1 _4783_ (.A(_0997_),
    .X(_0998_));
 sg13g2_nor2_1 _4784_ (.A(_0831_),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_nand2_2 _4785_ (.Y(_1000_),
    .A(net93),
    .B(net150));
 sg13g2_nor4_1 _4786_ (.A(net134),
    .B(_0880_),
    .C(_0958_),
    .D(_1000_),
    .Y(_1001_));
 sg13g2_nor4_1 _4787_ (.A(net171),
    .B(net92),
    .C(_0937_),
    .D(_1000_),
    .Y(_1002_));
 sg13g2_mux2_1 _4788_ (.A0(_1001_),
    .A1(_1002_),
    .S(_0891_),
    .X(_1003_));
 sg13g2_buf_2 _4789_ (.A(_1003_),
    .X(_1004_));
 sg13g2_xnor2_1 _4790_ (.Y(_1005_),
    .A(net240),
    .B(_2547_));
 sg13g2_and2_1 _4791_ (.A(net219),
    .B(_2542_),
    .X(_1006_));
 sg13g2_a221oi_1 _4792_ (.B2(net241),
    .C1(_1006_),
    .B1(net232),
    .A1(net167),
    .Y(_1007_),
    .A2(net208));
 sg13g2_nor3_1 _4793_ (.A(_1441_),
    .B(net208),
    .C(net209),
    .Y(_1008_));
 sg13g2_o21ai_1 _4794_ (.B1(net209),
    .Y(_1009_),
    .A1(_1441_),
    .A2(net208));
 sg13g2_o21ai_1 _4795_ (.B1(_1009_),
    .Y(_1010_),
    .A1(_0265_),
    .A2(_1008_));
 sg13g2_a21oi_1 _4796_ (.A1(net241),
    .A2(net232),
    .Y(_1011_),
    .B1(_1010_));
 sg13g2_a221oi_1 _4797_ (.B2(_1007_),
    .C1(_1011_),
    .B1(net108),
    .A1(_0311_),
    .Y(_1012_),
    .A2(_2549_));
 sg13g2_xor2_1 _4798_ (.B(_1012_),
    .A(_1005_),
    .X(_1013_));
 sg13g2_buf_8 _4799_ (.A(_1013_),
    .X(_1014_));
 sg13g2_buf_1 _4800_ (.A(_1014_),
    .X(_1015_));
 sg13g2_xor2_1 _4801_ (.B(net232),
    .A(_1364_),
    .X(_1016_));
 sg13g2_buf_1 _4802_ (.A(_1016_),
    .X(_1017_));
 sg13g2_nand2_1 _4803_ (.Y(_1018_),
    .A(net170),
    .B(_1010_));
 sg13g2_nand2b_1 _4804_ (.Y(_1019_),
    .B(net172),
    .A_N(_0837_));
 sg13g2_and2_1 _4805_ (.A(_1018_),
    .B(_1019_),
    .X(_1020_));
 sg13g2_buf_1 _4806_ (.A(_1020_),
    .X(_1021_));
 sg13g2_nor2_1 _4807_ (.A(net218),
    .B(net234),
    .Y(_1022_));
 sg13g2_nor2_2 _4808_ (.A(net191),
    .B(net209),
    .Y(_1023_));
 sg13g2_nor3_1 _4809_ (.A(net170),
    .B(_1022_),
    .C(_1023_),
    .Y(_1024_));
 sg13g2_nor2_1 _4810_ (.A(net185),
    .B(_2537_),
    .Y(_1025_));
 sg13g2_nor3_1 _4811_ (.A(_1006_),
    .B(_1025_),
    .C(net172),
    .Y(_1026_));
 sg13g2_mux2_1 _4812_ (.A0(_1024_),
    .A1(_1026_),
    .S(net108),
    .X(_1027_));
 sg13g2_nor2_1 _4813_ (.A(_1021_),
    .B(_1027_),
    .Y(_1028_));
 sg13g2_buf_1 _4814_ (.A(_1028_),
    .X(_1029_));
 sg13g2_nor2_1 _4815_ (.A(_2667_),
    .B(_1022_),
    .Y(_1030_));
 sg13g2_o21ai_1 _4816_ (.B1(_1030_),
    .Y(_1031_),
    .A1(net210),
    .A2(_0848_));
 sg13g2_o21ai_1 _4817_ (.B1(net210),
    .Y(_1032_),
    .A1(net207),
    .A2(net235));
 sg13g2_a221oi_1 _4818_ (.B2(_0845_),
    .C1(_1032_),
    .B1(_0844_),
    .A1(_0842_),
    .Y(_1033_),
    .A2(_0843_));
 sg13g2_nand2_1 _4819_ (.Y(_1034_),
    .A(_2564_),
    .B(_2537_));
 sg13g2_o21ai_1 _4820_ (.B1(_1034_),
    .Y(_1035_),
    .A1(_1025_),
    .A2(_1033_));
 sg13g2_nor2_1 _4821_ (.A(_0265_),
    .B(net233),
    .Y(_1036_));
 sg13g2_nor2b_1 _4822_ (.A(net219),
    .B_N(net233),
    .Y(_1037_));
 sg13g2_or2_1 _4823_ (.X(_1038_),
    .B(_1037_),
    .A(_1036_));
 sg13g2_buf_1 _4824_ (.A(_1038_),
    .X(_1039_));
 sg13g2_a21o_1 _4825_ (.A2(_1035_),
    .A1(_1031_),
    .B1(_1039_),
    .X(_1040_));
 sg13g2_buf_2 _4826_ (.A(_1040_),
    .X(_1041_));
 sg13g2_buf_1 _4827_ (.A(_1031_),
    .X(_1042_));
 sg13g2_buf_1 _4828_ (.A(_1035_),
    .X(_1043_));
 sg13g2_nand3_1 _4829_ (.B(net107),
    .C(net106),
    .A(_1039_),
    .Y(_1044_));
 sg13g2_buf_2 _4830_ (.A(_1044_),
    .X(_1045_));
 sg13g2_nand2_1 _4831_ (.Y(_1046_),
    .A(_1041_),
    .B(_1045_));
 sg13g2_buf_1 _4832_ (.A(_1046_),
    .X(_1047_));
 sg13g2_buf_1 _4833_ (.A(_1047_),
    .X(_1048_));
 sg13g2_xnor2_1 _4834_ (.Y(_1049_),
    .A(net108),
    .B(_0857_));
 sg13g2_buf_8 _4835_ (.A(_0848_),
    .X(_1050_));
 sg13g2_xnor2_1 _4836_ (.Y(_1051_),
    .A(net187),
    .B(net128));
 sg13g2_xnor2_1 _4837_ (.Y(_1052_),
    .A(_2667_),
    .B(_1051_));
 sg13g2_buf_8 _4838_ (.A(_1052_),
    .X(_1053_));
 sg13g2_nand2_2 _4839_ (.Y(_1054_),
    .A(_1049_),
    .B(_1053_));
 sg13g2_nand2_1 _4840_ (.Y(_1055_),
    .A(net34),
    .B(_1054_));
 sg13g2_nor2_1 _4841_ (.A(net49),
    .B(_1054_),
    .Y(_1056_));
 sg13g2_a21oi_1 _4842_ (.A1(_1029_),
    .A2(_1055_),
    .Y(_1057_),
    .B1(_1056_));
 sg13g2_nand2_1 _4843_ (.Y(_1058_),
    .A(_1018_),
    .B(_1019_));
 sg13g2_or3_1 _4844_ (.A(net170),
    .B(_1022_),
    .C(_1023_),
    .X(_1059_));
 sg13g2_nand2_1 _4845_ (.Y(_1060_),
    .A(net167),
    .B(net208));
 sg13g2_nand3_1 _4846_ (.B(_1060_),
    .C(net170),
    .A(_0833_),
    .Y(_1061_));
 sg13g2_mux2_1 _4847_ (.A0(_1059_),
    .A1(_1061_),
    .S(_0854_),
    .X(_1062_));
 sg13g2_nand2_1 _4848_ (.Y(_1063_),
    .A(_1058_),
    .B(_1062_));
 sg13g2_buf_1 _4849_ (.A(_1063_),
    .X(_1064_));
 sg13g2_xor2_1 _4850_ (.B(net208),
    .A(net218),
    .X(_1065_));
 sg13g2_xnor2_1 _4851_ (.Y(_1066_),
    .A(net108),
    .B(_1065_));
 sg13g2_buf_2 _4852_ (.A(_1066_),
    .X(_1067_));
 sg13g2_buf_1 _4853_ (.A(_1067_),
    .X(_1069_));
 sg13g2_nand4_1 _4854_ (.B(_1048_),
    .C(net62),
    .A(_1064_),
    .Y(_1070_),
    .D(net64));
 sg13g2_o21ai_1 _4855_ (.B1(_1070_),
    .Y(_1071_),
    .A1(_1015_),
    .A2(_1057_));
 sg13g2_xnor2_1 _4856_ (.Y(_1072_),
    .A(net166),
    .B(net128));
 sg13g2_nor2_1 _4857_ (.A(net155),
    .B(_0857_),
    .Y(_1073_));
 sg13g2_and2_1 _4858_ (.A(_0850_),
    .B(_0857_),
    .X(_1074_));
 sg13g2_nand3_1 _4859_ (.B(net166),
    .C(_1065_),
    .A(_2572_),
    .Y(_1075_));
 sg13g2_nor2_1 _4860_ (.A(net128),
    .B(_1075_),
    .Y(_1076_));
 sg13g2_a221oi_1 _4861_ (.B2(net128),
    .C1(_1076_),
    .B1(_1074_),
    .A1(_1072_),
    .Y(_1077_),
    .A2(_1073_));
 sg13g2_buf_2 _4862_ (.A(_1077_),
    .X(_1078_));
 sg13g2_buf_1 _4863_ (.A(_1078_),
    .X(_1080_));
 sg13g2_xnor2_1 _4864_ (.Y(_1081_),
    .A(_1005_),
    .B(_1012_));
 sg13g2_buf_1 _4865_ (.A(_1081_),
    .X(_1082_));
 sg13g2_nand2_1 _4866_ (.Y(_1083_),
    .A(net170),
    .B(_1023_));
 sg13g2_a21o_1 _4867_ (.A2(net106),
    .A1(net107),
    .B1(_1083_),
    .X(_1084_));
 sg13g2_nand4_1 _4868_ (.B(net170),
    .C(net107),
    .A(_1037_),
    .Y(_1085_),
    .D(net106));
 sg13g2_nand4_1 _4869_ (.B(_1017_),
    .C(net107),
    .A(_1036_),
    .Y(_1086_),
    .D(net106));
 sg13g2_nand2_1 _4870_ (.Y(_1087_),
    .A(_1006_),
    .B(_0859_));
 sg13g2_a21o_1 _4871_ (.A2(_1043_),
    .A1(_1042_),
    .B1(_1087_),
    .X(_1088_));
 sg13g2_nand4_1 _4872_ (.B(_1085_),
    .C(_1086_),
    .A(_1084_),
    .Y(_1089_),
    .D(_1088_));
 sg13g2_buf_2 _4873_ (.A(_1089_),
    .X(_1091_));
 sg13g2_nand2_2 _4874_ (.Y(_1092_),
    .A(net60),
    .B(_1091_));
 sg13g2_nor2_1 _4875_ (.A(net61),
    .B(_1092_),
    .Y(_1093_));
 sg13g2_nand2_1 _4876_ (.Y(_1094_),
    .A(_1028_),
    .B(net64));
 sg13g2_buf_1 _4877_ (.A(_1094_),
    .X(_1095_));
 sg13g2_inv_1 _4878_ (.Y(_1096_),
    .A(_1073_));
 sg13g2_nand2_1 _4879_ (.Y(_1097_),
    .A(_0850_),
    .B(_0857_));
 sg13g2_mux2_1 _4880_ (.A0(_1075_),
    .A1(_1097_),
    .S(net128),
    .X(_1098_));
 sg13g2_o21ai_1 _4881_ (.B1(_1098_),
    .Y(_1099_),
    .A1(_1051_),
    .A2(_1096_));
 sg13g2_buf_1 _4882_ (.A(_1099_),
    .X(_1100_));
 sg13g2_buf_1 _4883_ (.A(_1100_),
    .X(_1102_));
 sg13g2_a21oi_2 _4884_ (.B1(net59),
    .Y(_1103_),
    .A2(_1045_),
    .A1(_1041_));
 sg13g2_nor2_1 _4885_ (.A(net33),
    .B(_1103_),
    .Y(_1104_));
 sg13g2_or2_1 _4886_ (.X(_1105_),
    .B(_1104_),
    .A(_1093_));
 sg13g2_a21oi_2 _4887_ (.B1(net93),
    .Y(_1106_),
    .A2(_0992_),
    .A1(_0988_));
 sg13g2_nand2_1 _4888_ (.Y(_1107_),
    .A(_0922_),
    .B(_0926_));
 sg13g2_nand2_1 _4889_ (.Y(_1108_),
    .A(_1107_),
    .B(_0993_));
 sg13g2_buf_1 _4890_ (.A(net63),
    .X(_1109_));
 sg13g2_buf_1 _4891_ (.A(_1109_),
    .X(_1110_));
 sg13g2_buf_1 _4892_ (.A(net60),
    .X(_1111_));
 sg13g2_buf_1 _4893_ (.A(net47),
    .X(_1113_));
 sg13g2_xnor2_1 _4894_ (.Y(_1114_),
    .A(net49),
    .B(_1067_));
 sg13g2_nor2_1 _4895_ (.A(net49),
    .B(_1067_),
    .Y(_1115_));
 sg13g2_nor2_1 _4896_ (.A(_1067_),
    .B(_1053_),
    .Y(_1116_));
 sg13g2_a21oi_1 _4897_ (.A1(_1113_),
    .A2(_1115_),
    .Y(_1117_),
    .B1(_1116_));
 sg13g2_o21ai_1 _4898_ (.B1(_1117_),
    .Y(_1118_),
    .A1(_1113_),
    .A2(_1114_));
 sg13g2_buf_1 _4899_ (.A(net64),
    .X(_1119_));
 sg13g2_nor3_1 _4900_ (.A(net48),
    .B(net46),
    .C(_1055_),
    .Y(_1120_));
 sg13g2_a21oi_1 _4901_ (.A1(net32),
    .A2(_1118_),
    .Y(_1121_),
    .B1(_1120_));
 sg13g2_nand2_1 _4902_ (.Y(_1122_),
    .A(_1036_),
    .B(net172));
 sg13g2_nand2_1 _4903_ (.Y(_1124_),
    .A(_1037_),
    .B(net172));
 sg13g2_a22oi_1 _4904_ (.Y(_1125_),
    .B1(_1122_),
    .B2(_1124_),
    .A2(_1043_),
    .A1(_1042_));
 sg13g2_nand4_1 _4905_ (.B(net107),
    .C(net106),
    .A(net170),
    .Y(_1126_),
    .D(_1023_));
 sg13g2_nor2_1 _4906_ (.A(_0833_),
    .B(net170),
    .Y(_1127_));
 sg13g2_nand3_1 _4907_ (.B(net106),
    .C(_1127_),
    .A(net107),
    .Y(_1128_));
 sg13g2_nand3b_1 _4908_ (.B(_1126_),
    .C(_1128_),
    .Y(_1129_),
    .A_N(_1125_));
 sg13g2_buf_1 _4909_ (.A(_1129_),
    .X(_1130_));
 sg13g2_buf_1 _4910_ (.A(_1130_),
    .X(_1131_));
 sg13g2_and2_1 _4911_ (.A(_1041_),
    .B(_1045_),
    .X(_1132_));
 sg13g2_buf_1 _4912_ (.A(_1132_),
    .X(_1133_));
 sg13g2_buf_1 _4913_ (.A(_1133_),
    .X(_1135_));
 sg13g2_nor2_1 _4914_ (.A(net30),
    .B(_1078_),
    .Y(_1136_));
 sg13g2_a221oi_1 _4915_ (.B2(_0976_),
    .C1(net129),
    .B1(_0971_),
    .A1(net80),
    .Y(_1137_),
    .A2(_0967_));
 sg13g2_buf_1 _4916_ (.A(_1137_),
    .X(_1138_));
 sg13g2_o21ai_1 _4917_ (.B1(_1138_),
    .Y(_1139_),
    .A1(net45),
    .A2(_1136_));
 sg13g2_o21ai_1 _4918_ (.B1(_1139_),
    .Y(_1140_),
    .A1(_1108_),
    .A2(_1121_));
 sg13g2_a221oi_1 _4919_ (.B2(_1106_),
    .C1(_1140_),
    .B1(_1105_),
    .A1(_1004_),
    .Y(_1141_),
    .A2(_1071_));
 sg13g2_nand4_1 _4920_ (.B(_0931_),
    .C(_0863_),
    .A(net92),
    .Y(_1142_),
    .D(_0958_));
 sg13g2_a21oi_1 _4921_ (.A1(_0841_),
    .A2(_0862_),
    .Y(_1143_),
    .B1(_1142_));
 sg13g2_nand4_1 _4922_ (.B(net93),
    .C(_0867_),
    .A(net92),
    .Y(_1144_),
    .D(_0958_));
 sg13g2_nor3_1 _4923_ (.A(_0869_),
    .B(_0871_),
    .C(_1144_),
    .Y(_1146_));
 sg13g2_o21ai_1 _4924_ (.B1(net171),
    .Y(_1147_),
    .A1(_1143_),
    .A2(_1146_));
 sg13g2_mux2_1 _4925_ (.A0(net82),
    .A1(_0973_),
    .S(_0965_),
    .X(_1148_));
 sg13g2_nor3_1 _4926_ (.A(net171),
    .B(_0956_),
    .C(_1148_),
    .Y(_1149_));
 sg13g2_o21ai_1 _4927_ (.B1(_1149_),
    .Y(_1150_),
    .A1(net53),
    .A2(net52));
 sg13g2_a21o_1 _4928_ (.A2(_1150_),
    .A1(_1147_),
    .B1(net150),
    .X(_1151_));
 sg13g2_buf_1 _4929_ (.A(_1151_),
    .X(_1152_));
 sg13g2_a21oi_2 _4930_ (.B1(_1000_),
    .Y(_1153_),
    .A2(_0976_),
    .A1(_0971_));
 sg13g2_nand2_1 _4931_ (.Y(_1154_),
    .A(_1153_),
    .B(net31));
 sg13g2_nand3_1 _4932_ (.B(_1045_),
    .C(_1100_),
    .A(_1041_),
    .Y(_1155_));
 sg13g2_buf_2 _4933_ (.A(_1155_),
    .X(_1157_));
 sg13g2_a221oi_1 _4934_ (.B2(_1154_),
    .C1(_1157_),
    .B1(_1152_),
    .A1(_1058_),
    .Y(_1158_),
    .A2(_1062_));
 sg13g2_nand4_1 _4935_ (.B(net129),
    .C(_0894_),
    .A(net92),
    .Y(_1159_),
    .D(_0896_));
 sg13g2_a21oi_2 _4936_ (.B1(_1159_),
    .Y(_1160_),
    .A2(_0945_),
    .A1(_0940_));
 sg13g2_nor2_1 _4937_ (.A(net32),
    .B(_1114_),
    .Y(_1161_));
 sg13g2_a21oi_1 _4938_ (.A1(net45),
    .A2(_1116_),
    .Y(_1162_),
    .B1(_1161_));
 sg13g2_buf_1 _4939_ (.A(net60),
    .X(_1163_));
 sg13g2_buf_8 _4940_ (.A(_1054_),
    .X(_1164_));
 sg13g2_nand3_1 _4941_ (.B(net43),
    .C(_1091_),
    .A(net44),
    .Y(_1165_));
 sg13g2_o21ai_1 _4942_ (.B1(_1165_),
    .Y(_1166_),
    .A1(net31),
    .A2(_1162_));
 sg13g2_and2_1 _4943_ (.A(_1160_),
    .B(_1166_),
    .X(_1168_));
 sg13g2_nor2_1 _4944_ (.A(net34),
    .B(net44),
    .Y(_1169_));
 sg13g2_nor2_1 _4945_ (.A(net131),
    .B(_1033_),
    .Y(_1170_));
 sg13g2_nor2_1 _4946_ (.A(_1170_),
    .B(_1065_),
    .Y(_1171_));
 sg13g2_nand2_1 _4947_ (.Y(_1172_),
    .A(net135),
    .B(_1051_));
 sg13g2_nor3_1 _4948_ (.A(net128),
    .B(_0852_),
    .C(_0857_),
    .Y(_1173_));
 sg13g2_a21oi_2 _4949_ (.B1(_1173_),
    .Y(_1174_),
    .A2(_1172_),
    .A1(_1171_));
 sg13g2_nand3_1 _4950_ (.B(_1062_),
    .C(_1100_),
    .A(_1058_),
    .Y(_1175_));
 sg13g2_buf_1 _4951_ (.A(_1175_),
    .X(_1176_));
 sg13g2_o21ai_1 _4952_ (.B1(_1176_),
    .Y(_1177_),
    .A1(net50),
    .A2(_1174_));
 sg13g2_nor3_1 _4953_ (.A(net63),
    .B(net59),
    .C(net60),
    .Y(_1179_));
 sg13g2_a21o_1 _4954_ (.A2(net31),
    .A1(net32),
    .B1(_1179_),
    .X(_1180_));
 sg13g2_buf_1 _4955_ (.A(net49),
    .X(_1181_));
 sg13g2_buf_1 _4956_ (.A(net29),
    .X(_1182_));
 sg13g2_a22oi_1 _4957_ (.Y(_1183_),
    .B1(_1180_),
    .B2(net24),
    .A2(_1177_),
    .A1(_1169_));
 sg13g2_o21ai_1 _4958_ (.B1(net134),
    .Y(_1184_),
    .A1(_1143_),
    .A2(_1146_));
 sg13g2_nor3_1 _4959_ (.A(net153),
    .B(_0956_),
    .C(_1148_),
    .Y(_1185_));
 sg13g2_o21ai_1 _4960_ (.B1(_1185_),
    .Y(_1186_),
    .A1(_0865_),
    .A2(_0873_));
 sg13g2_a21oi_2 _4961_ (.B1(_0936_),
    .Y(_1187_),
    .A2(_1186_),
    .A1(_1184_));
 sg13g2_nor2b_1 _4962_ (.A(_1183_),
    .B_N(_1187_),
    .Y(_1188_));
 sg13g2_nand2_1 _4963_ (.Y(_1190_),
    .A(_2912_),
    .B(_1065_));
 sg13g2_nand2b_1 _4964_ (.Y(_1191_),
    .B(_0857_),
    .A_N(_0852_));
 sg13g2_nand3_1 _4965_ (.B(net187),
    .C(_1065_),
    .A(_2667_),
    .Y(_1192_));
 sg13g2_mux2_1 _4966_ (.A0(_1191_),
    .A1(_1192_),
    .S(net128),
    .X(_1193_));
 sg13g2_o21ai_1 _4967_ (.B1(_1193_),
    .Y(_1194_),
    .A1(_1051_),
    .A2(_1190_));
 sg13g2_buf_1 _4968_ (.A(_1194_),
    .X(_1195_));
 sg13g2_buf_1 _4969_ (.A(net79),
    .X(_1196_));
 sg13g2_nor3_1 _4970_ (.A(net63),
    .B(net49),
    .C(net60),
    .Y(_1197_));
 sg13g2_buf_1 _4971_ (.A(_1197_),
    .X(_1198_));
 sg13g2_nand2_1 _4972_ (.Y(_1199_),
    .A(net58),
    .B(net23));
 sg13g2_o21ai_1 _4973_ (.B1(_0956_),
    .Y(_1201_),
    .A1(net53),
    .A2(net52));
 sg13g2_nand3_1 _4974_ (.B(_0884_),
    .C(_0943_),
    .A(_0882_),
    .Y(_1202_));
 sg13g2_mux2_1 _4975_ (.A0(_1201_),
    .A1(_1202_),
    .S(_0880_),
    .X(_1203_));
 sg13g2_nand3_1 _4976_ (.B(net129),
    .C(_0898_),
    .A(net93),
    .Y(_1204_));
 sg13g2_nor3_1 _4977_ (.A(_1199_),
    .B(_1203_),
    .C(_1204_),
    .Y(_1205_));
 sg13g2_nor4_1 _4978_ (.A(_1158_),
    .B(_1168_),
    .C(_1188_),
    .D(_1205_),
    .Y(_1206_));
 sg13g2_nand2_1 _4979_ (.Y(_1207_),
    .A(net63),
    .B(net49));
 sg13g2_a21oi_2 _4980_ (.B1(net94),
    .Y(_1208_),
    .A2(_1186_),
    .A1(_1184_));
 sg13g2_nor2_1 _4981_ (.A(net134),
    .B(_0880_),
    .Y(_1209_));
 sg13g2_o21ai_1 _4982_ (.B1(_1209_),
    .Y(_1210_),
    .A1(_0960_),
    .A2(_0961_));
 sg13g2_nor2_1 _4983_ (.A(net171),
    .B(net92),
    .Y(_1212_));
 sg13g2_o21ai_1 _4984_ (.B1(_1212_),
    .Y(_1213_),
    .A1(_0955_),
    .A2(_0957_));
 sg13g2_a21oi_2 _4985_ (.B1(_1000_),
    .Y(_1214_),
    .A2(_1213_),
    .A1(_1210_));
 sg13g2_xnor2_1 _4986_ (.Y(_1215_),
    .A(_0278_),
    .B(_1051_));
 sg13g2_buf_2 _4987_ (.A(_1215_),
    .X(_1216_));
 sg13g2_nand2_1 _4988_ (.Y(_1217_),
    .A(_1049_),
    .B(_1216_));
 sg13g2_buf_1 _4989_ (.A(_1217_),
    .X(_1218_));
 sg13g2_nor2_1 _4990_ (.A(net42),
    .B(net31),
    .Y(_1219_));
 sg13g2_a22oi_1 _4991_ (.Y(_1220_),
    .B1(_1214_),
    .B2(_1219_),
    .A2(_1208_),
    .A1(net58));
 sg13g2_nor2_1 _4992_ (.A(_1207_),
    .B(_1220_),
    .Y(_1221_));
 sg13g2_xnor2_1 _4993_ (.Y(_1223_),
    .A(net32),
    .B(net43));
 sg13g2_buf_1 _4994_ (.A(_1028_),
    .X(_1224_));
 sg13g2_nand3_1 _4995_ (.B(_1048_),
    .C(net79),
    .A(_1224_),
    .Y(_1225_));
 sg13g2_o21ai_1 _4996_ (.B1(_1225_),
    .Y(_1226_),
    .A1(net24),
    .A2(_1223_));
 sg13g2_buf_1 _4997_ (.A(_1049_),
    .X(_1227_));
 sg13g2_nor2_1 _4998_ (.A(net78),
    .B(_1092_),
    .Y(_1228_));
 sg13g2_a21oi_1 _4999_ (.A1(net51),
    .A2(_1226_),
    .Y(_1229_),
    .B1(_1228_));
 sg13g2_o21ai_1 _5000_ (.B1(_0257_),
    .Y(_1230_),
    .A1(_0469_),
    .A2(_2558_));
 sg13g2_nand4_1 _5001_ (.B(_2728_),
    .C(_0888_),
    .A(net134),
    .Y(_1231_),
    .D(_1230_));
 sg13g2_a22oi_1 _5002_ (.Y(_1232_),
    .B1(_2768_),
    .B2(net151),
    .A2(_1167_),
    .A1(net120));
 sg13g2_nor3_1 _5003_ (.A(net153),
    .B(_0973_),
    .C(_1232_),
    .Y(_1234_));
 sg13g2_o21ai_1 _5004_ (.B1(_1234_),
    .Y(_1235_),
    .A1(_0865_),
    .A2(_0873_));
 sg13g2_o21ai_1 _5005_ (.B1(_1235_),
    .Y(_1236_),
    .A1(_0891_),
    .A2(_1231_));
 sg13g2_buf_1 _5006_ (.A(_1236_),
    .X(_1237_));
 sg13g2_nor2b_1 _5007_ (.A(_1229_),
    .B_N(_1237_),
    .Y(_1238_));
 sg13g2_and2_1 _5008_ (.A(_0894_),
    .B(_0896_),
    .X(_1239_));
 sg13g2_buf_1 _5009_ (.A(_1239_),
    .X(_1240_));
 sg13g2_nor2_1 _5010_ (.A(_0880_),
    .B(net129),
    .Y(_1241_));
 sg13g2_nor2_1 _5011_ (.A(_0935_),
    .B(_0963_),
    .Y(_1242_));
 sg13g2_nand3_1 _5012_ (.B(_1241_),
    .C(_1242_),
    .A(_1240_),
    .Y(_1243_));
 sg13g2_nor3_1 _5013_ (.A(net33),
    .B(_1157_),
    .C(_1243_),
    .Y(_1245_));
 sg13g2_nand3_1 _5014_ (.B(_1240_),
    .C(net23),
    .A(net129),
    .Y(_1246_));
 sg13g2_or3_1 _5015_ (.A(net80),
    .B(_1203_),
    .C(_1246_),
    .X(_1247_));
 sg13g2_nor2_1 _5016_ (.A(net42),
    .B(_1247_),
    .Y(_1248_));
 sg13g2_nor4_1 _5017_ (.A(_1221_),
    .B(_1238_),
    .C(_1245_),
    .D(_1248_),
    .Y(_1249_));
 sg13g2_nand3_1 _5018_ (.B(net80),
    .C(net150),
    .A(_0969_),
    .Y(_1250_));
 sg13g2_nor3_2 _5019_ (.A(_0898_),
    .B(_0963_),
    .C(_1250_),
    .Y(_1251_));
 sg13g2_nand2_1 _5020_ (.Y(_1252_),
    .A(net24),
    .B(_1053_));
 sg13g2_nor3_2 _5021_ (.A(_1240_),
    .B(_0963_),
    .C(_1250_),
    .Y(_1253_));
 sg13g2_a22oi_1 _5022_ (.Y(_1254_),
    .B1(_1253_),
    .B2(_1053_),
    .A2(_1252_),
    .A1(_1251_));
 sg13g2_nor3_1 _5023_ (.A(net62),
    .B(net33),
    .C(_1254_),
    .Y(_1256_));
 sg13g2_nand2_1 _5024_ (.Y(_1257_),
    .A(net41),
    .B(_1082_));
 sg13g2_nor2_1 _5025_ (.A(_1115_),
    .B(_1257_),
    .Y(_1258_));
 sg13g2_nand2_2 _5026_ (.Y(_1259_),
    .A(net107),
    .B(net106));
 sg13g2_nand4_1 _5027_ (.B(net172),
    .C(_1259_),
    .A(net209),
    .Y(_1260_),
    .D(net59));
 sg13g2_nand4_1 _5028_ (.B(net172),
    .C(_1259_),
    .A(net117),
    .Y(_1261_),
    .D(_1102_));
 sg13g2_o21ai_1 _5029_ (.B1(_1127_),
    .Y(_1262_),
    .A1(_1259_),
    .A2(_1102_));
 sg13g2_and3_1 _5030_ (.X(_1263_),
    .A(_1260_),
    .B(_1261_),
    .C(_1262_));
 sg13g2_o21ai_1 _5031_ (.B1(net117),
    .Y(_1264_),
    .A1(net209),
    .A2(_1259_));
 sg13g2_nand4_1 _5032_ (.B(net106),
    .C(_1023_),
    .A(net107),
    .Y(_1265_),
    .D(_1078_));
 sg13g2_a21oi_1 _5033_ (.A1(net209),
    .A2(_1259_),
    .Y(_1267_),
    .B1(net172));
 sg13g2_nand3_1 _5034_ (.B(_1265_),
    .C(_1267_),
    .A(_1264_),
    .Y(_1268_));
 sg13g2_a21oi_1 _5035_ (.A1(_1263_),
    .A2(_1268_),
    .Y(_1269_),
    .B1(_1111_));
 sg13g2_o21ai_1 _5036_ (.B1(_1153_),
    .Y(_1270_),
    .A1(_1258_),
    .A2(_1269_));
 sg13g2_and2_1 _5037_ (.A(net60),
    .B(_1091_),
    .X(_1271_));
 sg13g2_buf_1 _5038_ (.A(_1271_),
    .X(_1272_));
 sg13g2_nor2_2 _5039_ (.A(net63),
    .B(_1082_),
    .Y(_1273_));
 sg13g2_nor4_1 _5040_ (.A(net41),
    .B(_1047_),
    .C(_1078_),
    .D(net64),
    .Y(_1274_));
 sg13g2_a221oi_1 _5041_ (.B2(net29),
    .C1(_1274_),
    .B1(_1273_),
    .A1(_1078_),
    .Y(_1275_),
    .A2(_1272_));
 sg13g2_or2_1 _5042_ (.X(_1276_),
    .B(_1275_),
    .A(_1152_));
 sg13g2_nand3_1 _5043_ (.B(net49),
    .C(_1067_),
    .A(net41),
    .Y(_1278_));
 sg13g2_nand3_1 _5044_ (.B(net30),
    .C(_1227_),
    .A(net63),
    .Y(_1279_));
 sg13g2_a21oi_1 _5045_ (.A1(_1278_),
    .A2(_1279_),
    .Y(_1280_),
    .B1(net47));
 sg13g2_nor2_1 _5046_ (.A(_1133_),
    .B(net79),
    .Y(_1281_));
 sg13g2_nor4_1 _5047_ (.A(net50),
    .B(net46),
    .C(_1281_),
    .D(_1056_),
    .Y(_1282_));
 sg13g2_o21ai_1 _5048_ (.B1(_1214_),
    .Y(_1283_),
    .A1(_1280_),
    .A2(_1282_));
 sg13g2_a221oi_1 _5049_ (.B2(net50),
    .C1(net44),
    .B1(_1281_),
    .A1(_1130_),
    .Y(_1284_),
    .A2(_1195_));
 sg13g2_o21ai_1 _5050_ (.B1(_1111_),
    .Y(_1285_),
    .A1(_1029_),
    .A2(_1114_));
 sg13g2_nand3b_1 _5051_ (.B(_1285_),
    .C(_1208_),
    .Y(_1286_),
    .A_N(_1284_));
 sg13g2_nand4_1 _5052_ (.B(_1276_),
    .C(_1283_),
    .A(_1270_),
    .Y(_1287_),
    .D(_1286_));
 sg13g2_nand2_1 _5053_ (.Y(_1289_),
    .A(_0940_),
    .B(_0945_));
 sg13g2_a21o_1 _5054_ (.A2(_1172_),
    .A1(_1171_),
    .B1(_1173_),
    .X(_1290_));
 sg13g2_buf_1 _5055_ (.A(_1290_),
    .X(_1291_));
 sg13g2_a22oi_1 _5056_ (.Y(_1292_),
    .B1(net57),
    .B2(_1242_),
    .A2(_1157_),
    .A1(_1289_));
 sg13g2_nand2_1 _5057_ (.Y(_1293_),
    .A(_1289_),
    .B(net57));
 sg13g2_o21ai_1 _5058_ (.B1(_1293_),
    .Y(_1294_),
    .A1(net24),
    .A2(_1292_));
 sg13g2_and4_1 _5059_ (.A(_0898_),
    .B(_1241_),
    .C(_1273_),
    .D(_1294_),
    .X(_1295_));
 sg13g2_nor3_1 _5060_ (.A(_1256_),
    .B(_1287_),
    .C(_1295_),
    .Y(_1296_));
 sg13g2_nand4_1 _5061_ (.B(_1206_),
    .C(_1249_),
    .A(_1141_),
    .Y(_1297_),
    .D(_1296_));
 sg13g2_inv_1 _5062_ (.Y(_1298_),
    .A(net230));
 sg13g2_a21oi_1 _5063_ (.A1(_1298_),
    .A2(_0845_),
    .Y(_1300_),
    .B1(_0843_));
 sg13g2_xor2_1 _5064_ (.B(net211),
    .A(_2569_),
    .X(_1301_));
 sg13g2_xnor2_1 _5065_ (.Y(_1302_),
    .A(_1300_),
    .B(_1301_));
 sg13g2_nand2b_2 _5066_ (.Y(_1303_),
    .B(net242),
    .A_N(_1302_));
 sg13g2_nor2_1 _5067_ (.A(_1053_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_a21oi_1 _5068_ (.A1(_1053_),
    .A2(_1303_),
    .Y(_1305_),
    .B1(_1332_));
 sg13g2_or2_1 _5069_ (.X(_1306_),
    .B(_1305_),
    .A(_1304_));
 sg13g2_xnor2_1 _5070_ (.Y(_1307_),
    .A(net143),
    .B(_1067_));
 sg13g2_inv_1 _5071_ (.Y(_1308_),
    .A(_1307_));
 sg13g2_a22oi_1 _5072_ (.Y(_1309_),
    .B1(_1306_),
    .B2(_1308_),
    .A2(_1067_),
    .A1(_0619_));
 sg13g2_xnor2_1 _5073_ (.Y(_1311_),
    .A(net120),
    .B(net30));
 sg13g2_xnor2_1 _5074_ (.Y(_1312_),
    .A(_1309_),
    .B(_1311_));
 sg13g2_buf_1 _5075_ (.A(_1312_),
    .X(_1313_));
 sg13g2_xnor2_1 _5076_ (.Y(_1314_),
    .A(_1306_),
    .B(_1308_));
 sg13g2_buf_2 _5077_ (.A(_1314_),
    .X(_1315_));
 sg13g2_xnor2_1 _5078_ (.Y(_1316_),
    .A(_2555_),
    .B(_1216_));
 sg13g2_buf_2 _5079_ (.A(_1316_),
    .X(_1317_));
 sg13g2_xnor2_1 _5080_ (.Y(_1318_),
    .A(_1303_),
    .B(_1317_));
 sg13g2_nor2_1 _5081_ (.A(_1315_),
    .B(_1318_),
    .Y(_1319_));
 sg13g2_xnor2_1 _5082_ (.Y(_1320_),
    .A(net18),
    .B(_1319_));
 sg13g2_xnor2_1 _5083_ (.Y(_1322_),
    .A(net240),
    .B(net232));
 sg13g2_xnor2_1 _5084_ (.Y(_1323_),
    .A(_1386_),
    .B(net234));
 sg13g2_buf_2 _5085_ (.A(_1323_),
    .X(_1324_));
 sg13g2_nor2_1 _5086_ (.A(\graphics_engine_1.overlay_creator1.text_demosiine1.x[6] ),
    .B(net233),
    .Y(_1325_));
 sg13g2_nor2_1 _5087_ (.A(_1419_),
    .B(_2532_),
    .Y(_1326_));
 sg13g2_buf_2 _5088_ (.A(_1326_),
    .X(_1327_));
 sg13g2_nor3_1 _5089_ (.A(_1324_),
    .B(_1325_),
    .C(_1327_),
    .Y(_1328_));
 sg13g2_nor2_2 _5090_ (.A(_2567_),
    .B(_2525_),
    .Y(_1329_));
 sg13g2_a22oi_1 _5091_ (.Y(_1330_),
    .B1(net236),
    .B2(net230),
    .A2(_2525_),
    .A1(_2567_));
 sg13g2_buf_2 _5092_ (.A(_1330_),
    .X(_1331_));
 sg13g2_a22oi_1 _5093_ (.Y(_1333_),
    .B1(net211),
    .B2(net206),
    .A2(_2532_),
    .A1(net218));
 sg13g2_o21ai_1 _5094_ (.B1(_1333_),
    .Y(_1334_),
    .A1(_1329_),
    .A2(_1331_));
 sg13g2_nand2_1 _5095_ (.Y(_1335_),
    .A(_1419_),
    .B(_2532_));
 sg13g2_buf_2 _5096_ (.A(_1335_),
    .X(_1336_));
 sg13g2_nor2_1 _5097_ (.A(_2570_),
    .B(net235),
    .Y(_1337_));
 sg13g2_buf_1 _5098_ (.A(_1337_),
    .X(_1338_));
 sg13g2_nand2_1 _5099_ (.Y(_1339_),
    .A(_1336_),
    .B(_1338_));
 sg13g2_nand4_1 _5100_ (.B(_1328_),
    .C(_1334_),
    .A(_1322_),
    .Y(_1340_),
    .D(_1339_));
 sg13g2_a22oi_1 _5101_ (.Y(_1341_),
    .B1(net233),
    .B2(net241),
    .A2(net234),
    .A1(_1386_));
 sg13g2_nor2_1 _5102_ (.A(_1325_),
    .B(_1341_),
    .Y(_1342_));
 sg13g2_nand2_1 _5103_ (.Y(_1344_),
    .A(_1322_),
    .B(_1342_));
 sg13g2_xor2_1 _5104_ (.B(net232),
    .A(_1474_),
    .X(_1345_));
 sg13g2_o21ai_1 _5105_ (.B1(_1345_),
    .Y(_1346_),
    .A1(_1325_),
    .A2(_1341_));
 sg13g2_or2_1 _5106_ (.X(_1347_),
    .B(_1346_),
    .A(_1334_));
 sg13g2_a21o_1 _5107_ (.A2(_1339_),
    .A1(_1328_),
    .B1(_1346_),
    .X(_1348_));
 sg13g2_nand4_1 _5108_ (.B(_1344_),
    .C(_1347_),
    .A(_1340_),
    .Y(_1349_),
    .D(_1348_));
 sg13g2_buf_1 _5109_ (.A(_1349_),
    .X(_1350_));
 sg13g2_buf_1 _5110_ (.A(_1350_),
    .X(_1351_));
 sg13g2_nor2_1 _5111_ (.A(net133),
    .B(net154),
    .Y(_1352_));
 sg13g2_o21ai_1 _5112_ (.B1(_1352_),
    .Y(_1353_),
    .A1(_1277_),
    .A2(net77));
 sg13g2_buf_2 _5113_ (.A(_1353_),
    .X(_1354_));
 sg13g2_and4_1 _5114_ (.A(_1340_),
    .B(_1344_),
    .C(_1347_),
    .D(_1348_),
    .X(_1355_));
 sg13g2_buf_2 _5115_ (.A(_1355_),
    .X(_1356_));
 sg13g2_buf_1 _5116_ (.A(_1356_),
    .X(_1357_));
 sg13g2_nor2_1 _5117_ (.A(net225),
    .B(net202),
    .Y(_1358_));
 sg13g2_nand3_1 _5118_ (.B(net76),
    .C(_1358_),
    .A(_2606_),
    .Y(_1359_));
 sg13g2_buf_2 _5119_ (.A(_1359_),
    .X(_1360_));
 sg13g2_and2_1 _5120_ (.A(_1354_),
    .B(_1360_),
    .X(_1361_));
 sg13g2_or2_1 _5121_ (.X(_1362_),
    .B(net235),
    .A(net206));
 sg13g2_buf_2 _5122_ (.A(_1362_),
    .X(_1363_));
 sg13g2_nand2_2 _5123_ (.Y(_1365_),
    .A(net210),
    .B(_1363_));
 sg13g2_nor4_1 _5124_ (.A(_1329_),
    .B(_1331_),
    .C(_1324_),
    .D(_1365_),
    .Y(_1366_));
 sg13g2_xor2_1 _5125_ (.B(net208),
    .A(net219),
    .X(_1367_));
 sg13g2_nand3_1 _5126_ (.B(_1363_),
    .C(_1367_),
    .A(_1562_),
    .Y(_1368_));
 sg13g2_nor3_1 _5127_ (.A(_1329_),
    .B(_1331_),
    .C(_1368_),
    .Y(_1369_));
 sg13g2_buf_1 _5128_ (.A(_1324_),
    .X(_1370_));
 sg13g2_nor2_1 _5129_ (.A(_1336_),
    .B(net149),
    .Y(_1371_));
 sg13g2_and2_1 _5130_ (.A(_2570_),
    .B(net235),
    .X(_1372_));
 sg13g2_buf_1 _5131_ (.A(_1372_),
    .X(_1373_));
 sg13g2_nand2_1 _5132_ (.Y(_1374_),
    .A(net187),
    .B(_1373_));
 sg13g2_nand2_1 _5133_ (.Y(_1376_),
    .A(_1562_),
    .B(_1373_));
 sg13g2_a21oi_1 _5134_ (.A1(_1374_),
    .A2(_1376_),
    .Y(_1377_),
    .B1(net149));
 sg13g2_nor4_1 _5135_ (.A(_1366_),
    .B(_1369_),
    .C(_1371_),
    .D(_1377_),
    .Y(_1378_));
 sg13g2_buf_2 _5136_ (.A(_1378_),
    .X(_1379_));
 sg13g2_nand2_1 _5137_ (.Y(_1380_),
    .A(net206),
    .B(net211));
 sg13g2_o21ai_1 _5138_ (.B1(_1380_),
    .Y(_1381_),
    .A1(_1329_),
    .A2(_1331_));
 sg13g2_a21oi_1 _5139_ (.A1(_1381_),
    .A2(_1363_),
    .Y(_1382_),
    .B1(net187));
 sg13g2_buf_2 _5140_ (.A(_1382_),
    .X(_1383_));
 sg13g2_buf_1 _5141_ (.A(_1381_),
    .X(_1384_));
 sg13g2_nor2_1 _5142_ (.A(_2538_),
    .B(_1338_),
    .Y(_1385_));
 sg13g2_a21oi_1 _5143_ (.A1(net127),
    .A2(_1385_),
    .Y(_1387_),
    .B1(net137));
 sg13g2_buf_1 _5144_ (.A(_1370_),
    .X(_1388_));
 sg13g2_o21ai_1 _5145_ (.B1(_1388_),
    .Y(_1389_),
    .A1(_1383_),
    .A2(_1387_));
 sg13g2_buf_2 _5146_ (.A(_1389_),
    .X(_1390_));
 sg13g2_xor2_1 _5147_ (.B(net210),
    .A(net218),
    .X(_1391_));
 sg13g2_buf_1 _5148_ (.A(_1391_),
    .X(_1392_));
 sg13g2_nor2_1 _5149_ (.A(_1338_),
    .B(_1392_),
    .Y(_1393_));
 sg13g2_and2_1 _5150_ (.A(_1384_),
    .B(_1393_),
    .X(_1394_));
 sg13g2_buf_1 _5151_ (.A(_1394_),
    .X(_1395_));
 sg13g2_xnor2_1 _5152_ (.Y(_1396_),
    .A(net190),
    .B(net210));
 sg13g2_a21oi_2 _5153_ (.B1(_1396_),
    .Y(_1398_),
    .A2(_1363_),
    .A1(net127));
 sg13g2_and2_1 _5154_ (.A(net230),
    .B(net236),
    .X(_1399_));
 sg13g2_buf_2 _5155_ (.A(_1399_),
    .X(_1400_));
 sg13g2_xnor2_1 _5156_ (.Y(_1401_),
    .A(net207),
    .B(net212));
 sg13g2_xnor2_1 _5157_ (.Y(_1402_),
    .A(_1400_),
    .B(_1401_));
 sg13g2_xnor2_1 _5158_ (.Y(_1403_),
    .A(_2570_),
    .B(_2529_));
 sg13g2_o21ai_1 _5159_ (.B1(_1403_),
    .Y(_1404_),
    .A1(_1329_),
    .A2(_1331_));
 sg13g2_buf_1 _5160_ (.A(_1404_),
    .X(_1405_));
 sg13g2_or3_1 _5161_ (.A(_1329_),
    .B(_1331_),
    .C(_1403_),
    .X(_1406_));
 sg13g2_buf_1 _5162_ (.A(_1406_),
    .X(_1407_));
 sg13g2_and3_1 _5163_ (.X(_1409_),
    .A(_1402_),
    .B(net125),
    .C(net124));
 sg13g2_buf_1 _5164_ (.A(_1409_),
    .X(_1410_));
 sg13g2_o21ai_1 _5165_ (.B1(_1410_),
    .Y(_1411_),
    .A1(_1395_),
    .A2(_1398_));
 sg13g2_buf_1 _5166_ (.A(_1411_),
    .X(_1412_));
 sg13g2_buf_1 _5167_ (.A(_1384_),
    .X(_1413_));
 sg13g2_nand2_2 _5168_ (.Y(_1414_),
    .A(net105),
    .B(_1393_));
 sg13g2_or2_1 _5169_ (.X(_1415_),
    .B(_2525_),
    .A(net207));
 sg13g2_and2_1 _5170_ (.A(net207),
    .B(_2525_),
    .X(_1416_));
 sg13g2_a221oi_1 _5171_ (.B2(_1400_),
    .C1(_1416_),
    .B1(_1415_),
    .A1(_2571_),
    .Y(_1417_),
    .A2(_2530_));
 sg13g2_buf_2 _5172_ (.A(_1417_),
    .X(_1418_));
 sg13g2_buf_1 _5173_ (.A(_1418_),
    .X(_1420_));
 sg13g2_buf_1 _5174_ (.A(_1338_),
    .X(_1421_));
 sg13g2_o21ai_1 _5175_ (.B1(net148),
    .Y(_1422_),
    .A1(net104),
    .A2(net147));
 sg13g2_buf_1 _5176_ (.A(_1422_),
    .X(_1423_));
 sg13g2_nand2_1 _5177_ (.Y(_1424_),
    .A(net230),
    .B(net236));
 sg13g2_xnor2_1 _5178_ (.Y(_1425_),
    .A(_1424_),
    .B(_1401_));
 sg13g2_buf_1 _5179_ (.A(_1425_),
    .X(_1426_));
 sg13g2_and3_1 _5180_ (.X(_1427_),
    .A(_1426_),
    .B(net125),
    .C(net124));
 sg13g2_buf_1 _5181_ (.A(_1427_),
    .X(_1428_));
 sg13g2_nand3_1 _5182_ (.B(_1423_),
    .C(_1428_),
    .A(_1414_),
    .Y(_1429_));
 sg13g2_a22oi_1 _5183_ (.Y(_1431_),
    .B1(_1412_),
    .B2(_1429_),
    .A2(_1390_),
    .A1(_1379_));
 sg13g2_nand4_1 _5184_ (.B(_2530_),
    .C(_2526_),
    .A(net230),
    .Y(_1432_),
    .D(net236));
 sg13g2_nand4_1 _5185_ (.B(net207),
    .C(net211),
    .A(_2575_),
    .Y(_1433_),
    .D(net236));
 sg13g2_nand3_1 _5186_ (.B(net211),
    .C(net212),
    .A(_2568_),
    .Y(_1434_));
 sg13g2_nand4_1 _5187_ (.B(net206),
    .C(net212),
    .A(_2575_),
    .Y(_1435_),
    .D(net236));
 sg13g2_and4_1 _5188_ (.A(_1432_),
    .B(_1433_),
    .C(_1434_),
    .D(_1435_),
    .X(_1436_));
 sg13g2_buf_1 _5189_ (.A(_1436_),
    .X(_1437_));
 sg13g2_a221oi_1 _5190_ (.B2(_2714_),
    .C1(_1373_),
    .B1(_1400_),
    .A1(_2571_),
    .Y(_1438_),
    .A2(_1416_));
 sg13g2_buf_1 _5191_ (.A(_1438_),
    .X(_1439_));
 sg13g2_and2_1 _5192_ (.A(net219),
    .B(_2543_),
    .X(_1440_));
 sg13g2_xor2_1 _5193_ (.B(_2541_),
    .A(net241),
    .X(_1442_));
 sg13g2_nor2_1 _5194_ (.A(_1440_),
    .B(_1442_),
    .Y(_1443_));
 sg13g2_nand4_1 _5195_ (.B(_1437_),
    .C(_1439_),
    .A(net166),
    .Y(_1444_),
    .D(_1443_));
 sg13g2_or2_1 _5196_ (.X(_1445_),
    .B(_2536_),
    .A(_1397_));
 sg13g2_buf_1 _5197_ (.A(_1445_),
    .X(_1446_));
 sg13g2_nor2_1 _5198_ (.A(_1442_),
    .B(_1446_),
    .Y(_1447_));
 sg13g2_inv_1 _5199_ (.Y(_1448_),
    .A(_1447_));
 sg13g2_xnor2_1 _5200_ (.Y(_1449_),
    .A(net241),
    .B(net233));
 sg13g2_a21oi_1 _5201_ (.A1(_1397_),
    .A2(_2543_),
    .Y(_1450_),
    .B1(net218));
 sg13g2_and2_1 _5202_ (.A(_1449_),
    .B(_1450_),
    .X(_1451_));
 sg13g2_o21ai_1 _5203_ (.B1(_1451_),
    .Y(_1453_),
    .A1(_1418_),
    .A2(_1365_));
 sg13g2_and3_1 _5204_ (.X(_1454_),
    .A(_1444_),
    .B(_1448_),
    .C(_1453_));
 sg13g2_buf_2 _5205_ (.A(_1454_),
    .X(_1455_));
 sg13g2_o21ai_1 _5206_ (.B1(_1450_),
    .Y(_1456_),
    .A1(_1418_),
    .A2(_1365_));
 sg13g2_nor2_1 _5207_ (.A(net210),
    .B(_1440_),
    .Y(_1457_));
 sg13g2_o21ai_1 _5208_ (.B1(_1457_),
    .Y(_1458_),
    .A1(_1418_),
    .A2(_1338_));
 sg13g2_nand4_1 _5209_ (.B(_1446_),
    .C(_1456_),
    .A(_1442_),
    .Y(_1459_),
    .D(_1458_));
 sg13g2_buf_2 _5210_ (.A(_1459_),
    .X(_1460_));
 sg13g2_nand2_1 _5211_ (.Y(_1461_),
    .A(_1455_),
    .B(_1460_));
 sg13g2_buf_2 _5212_ (.A(_1461_),
    .X(_1462_));
 sg13g2_buf_1 _5213_ (.A(_1462_),
    .X(_1464_));
 sg13g2_buf_1 _5214_ (.A(net28),
    .X(_1465_));
 sg13g2_and2_1 _5215_ (.A(net125),
    .B(net124),
    .X(_1466_));
 sg13g2_buf_1 _5216_ (.A(_1466_),
    .X(_1467_));
 sg13g2_o21ai_1 _5217_ (.B1(net166),
    .Y(_1468_),
    .A1(_1418_),
    .A2(_1338_));
 sg13g2_buf_1 _5218_ (.A(_1468_),
    .X(_1469_));
 sg13g2_nand2_1 _5219_ (.Y(_1470_),
    .A(net137),
    .B(_1324_));
 sg13g2_a21oi_1 _5220_ (.A1(net127),
    .A2(_1385_),
    .Y(_1471_),
    .B1(_1470_));
 sg13g2_buf_1 _5221_ (.A(_1367_),
    .X(_1472_));
 sg13g2_nor2_1 _5222_ (.A(net137),
    .B(net146),
    .Y(_1473_));
 sg13g2_nor2_2 _5223_ (.A(net104),
    .B(_1365_),
    .Y(_1475_));
 sg13g2_buf_1 _5224_ (.A(_1363_),
    .X(_1476_));
 sg13g2_nand2_1 _5225_ (.Y(_1477_),
    .A(net146),
    .B(_1327_));
 sg13g2_a21oi_1 _5226_ (.A1(net127),
    .A2(net123),
    .Y(_1478_),
    .B1(_1477_));
 sg13g2_a221oi_1 _5227_ (.B2(_1475_),
    .C1(_1478_),
    .B1(_1473_),
    .A1(_1469_),
    .Y(_1479_),
    .A2(_1471_));
 sg13g2_buf_2 _5228_ (.A(_1479_),
    .X(_1480_));
 sg13g2_or2_1 _5229_ (.X(_1481_),
    .B(_1480_),
    .A(net90));
 sg13g2_buf_1 _5230_ (.A(_1481_),
    .X(_1482_));
 sg13g2_nand3b_1 _5231_ (.B(net22),
    .C(_1482_),
    .Y(_1483_),
    .A_N(_1431_));
 sg13g2_nand3_1 _5232_ (.B(_1448_),
    .C(_1453_),
    .A(_1444_),
    .Y(_1484_));
 sg13g2_and4_1 _5233_ (.A(_1442_),
    .B(_1446_),
    .C(_1456_),
    .D(_1458_),
    .X(_1486_));
 sg13g2_buf_1 _5234_ (.A(_1486_),
    .X(_1487_));
 sg13g2_nor2_1 _5235_ (.A(_1484_),
    .B(_1487_),
    .Y(_1488_));
 sg13g2_buf_1 _5236_ (.A(_1488_),
    .X(_1489_));
 sg13g2_buf_1 _5237_ (.A(_1489_),
    .X(_1490_));
 sg13g2_a21oi_1 _5238_ (.A1(net125),
    .A2(net124),
    .Y(_1491_),
    .B1(_1426_));
 sg13g2_buf_1 _5239_ (.A(_1491_),
    .X(_1492_));
 sg13g2_nand4_1 _5240_ (.B(_1363_),
    .C(net146),
    .A(net127),
    .Y(_1493_),
    .D(_1327_));
 sg13g2_nand2b_1 _5241_ (.Y(_1494_),
    .B(_2533_),
    .A_N(net190));
 sg13g2_nor2_1 _5242_ (.A(_1324_),
    .B(_1494_),
    .Y(_1495_));
 sg13g2_o21ai_1 _5243_ (.B1(_1495_),
    .Y(_1497_),
    .A1(_1418_),
    .A2(net147));
 sg13g2_nor2_1 _5244_ (.A(net185),
    .B(_2533_),
    .Y(_1498_));
 sg13g2_nand4_1 _5245_ (.B(_1439_),
    .C(net146),
    .A(_1437_),
    .Y(_1499_),
    .D(_1498_));
 sg13g2_nor2_2 _5246_ (.A(net185),
    .B(net166),
    .Y(_1500_));
 sg13g2_nand4_1 _5247_ (.B(net127),
    .C(_1363_),
    .A(_1500_),
    .Y(_1501_),
    .D(_1370_));
 sg13g2_nand4_1 _5248_ (.B(_1497_),
    .C(_1499_),
    .A(_1493_),
    .Y(_1502_),
    .D(_1501_));
 sg13g2_buf_1 _5249_ (.A(_1502_),
    .X(_1503_));
 sg13g2_nand2_1 _5250_ (.Y(_1504_),
    .A(net89),
    .B(net75));
 sg13g2_nand2_1 _5251_ (.Y(_1505_),
    .A(net174),
    .B(_0814_));
 sg13g2_xnor2_1 _5252_ (.Y(_1506_),
    .A(_2777_),
    .B(_0145_));
 sg13g2_nand2_1 _5253_ (.Y(_1508_),
    .A(_2793_),
    .B(_1506_));
 sg13g2_mux2_1 _5254_ (.A0(_1505_),
    .A1(_1508_),
    .S(net77),
    .X(_1509_));
 sg13g2_buf_1 _5255_ (.A(_1509_),
    .X(_1510_));
 sg13g2_buf_1 _5256_ (.A(_1510_),
    .X(_1511_));
 sg13g2_a21oi_1 _5257_ (.A1(net27),
    .A2(_1504_),
    .Y(_1512_),
    .B1(net26));
 sg13g2_buf_1 _5258_ (.A(_1488_),
    .X(_1513_));
 sg13g2_a21o_1 _5259_ (.A2(net124),
    .A1(net125),
    .B1(_1402_),
    .X(_1514_));
 sg13g2_buf_2 _5260_ (.A(_1514_),
    .X(_1515_));
 sg13g2_nor2_1 _5261_ (.A(_1515_),
    .B(_1480_),
    .Y(_1516_));
 sg13g2_o21ai_1 _5262_ (.B1(net90),
    .Y(_1517_),
    .A1(_1395_),
    .A2(_1398_));
 sg13g2_nand3_1 _5263_ (.B(_1423_),
    .C(_1492_),
    .A(_1414_),
    .Y(_1519_));
 sg13g2_a22oi_1 _5264_ (.Y(_1520_),
    .B1(_1517_),
    .B2(_1519_),
    .A2(_1390_),
    .A1(_1379_));
 sg13g2_or3_1 _5265_ (.A(net39),
    .B(_1516_),
    .C(_1520_),
    .X(_1521_));
 sg13g2_nand2_1 _5266_ (.Y(_1522_),
    .A(net75),
    .B(net91));
 sg13g2_nand2_1 _5267_ (.Y(_1523_),
    .A(net174),
    .B(_2793_));
 sg13g2_nand2_1 _5268_ (.Y(_1524_),
    .A(_0814_),
    .B(_1506_));
 sg13g2_mux2_1 _5269_ (.A0(_1523_),
    .A1(_1524_),
    .S(_1350_),
    .X(_1525_));
 sg13g2_buf_2 _5270_ (.A(_1525_),
    .X(_1526_));
 sg13g2_a21oi_1 _5271_ (.A1(_1490_),
    .A2(_1522_),
    .Y(_1527_),
    .B1(_1526_));
 sg13g2_a22oi_1 _5272_ (.Y(_1528_),
    .B1(_1521_),
    .B2(_1527_),
    .A2(_1512_),
    .A1(_1483_));
 sg13g2_o21ai_1 _5273_ (.B1(net185),
    .Y(_1530_),
    .A1(net104),
    .A2(_1365_));
 sg13g2_nand3_1 _5274_ (.B(_1469_),
    .C(_1530_),
    .A(net126),
    .Y(_1531_));
 sg13g2_buf_2 _5275_ (.A(_1531_),
    .X(_1532_));
 sg13g2_o21ai_1 _5276_ (.B1(_1472_),
    .Y(_1533_),
    .A1(_1383_),
    .A2(_1387_));
 sg13g2_buf_1 _5277_ (.A(_1533_),
    .X(_1534_));
 sg13g2_nand2_1 _5278_ (.Y(_1535_),
    .A(_1532_),
    .B(_1534_));
 sg13g2_buf_1 _5279_ (.A(_1535_),
    .X(_1536_));
 sg13g2_buf_1 _5280_ (.A(_1402_),
    .X(_1537_));
 sg13g2_a21oi_1 _5281_ (.A1(_1405_),
    .A2(net124),
    .Y(_1538_),
    .B1(net122));
 sg13g2_buf_1 _5282_ (.A(_1538_),
    .X(_1539_));
 sg13g2_o21ai_1 _5283_ (.B1(net88),
    .Y(_1541_),
    .A1(_1395_),
    .A2(_1398_));
 sg13g2_buf_1 _5284_ (.A(_1541_),
    .X(_1542_));
 sg13g2_nor3_1 _5285_ (.A(net27),
    .B(net25),
    .C(_1542_),
    .Y(_1543_));
 sg13g2_nand3_1 _5286_ (.B(net125),
    .C(net124),
    .A(net122),
    .Y(_1544_));
 sg13g2_buf_1 _5287_ (.A(_1544_),
    .X(_1545_));
 sg13g2_buf_1 _5288_ (.A(_1545_),
    .X(_1546_));
 sg13g2_buf_1 _5289_ (.A(_1515_),
    .X(_1547_));
 sg13g2_o21ai_1 _5290_ (.B1(net73),
    .Y(_1548_),
    .A1(_1484_),
    .A2(_1487_));
 sg13g2_buf_1 _5291_ (.A(_1480_),
    .X(_1549_));
 sg13g2_a21oi_1 _5292_ (.A1(_1546_),
    .A2(_1548_),
    .Y(_1550_),
    .B1(_1549_));
 sg13g2_nand2_1 _5293_ (.Y(_1552_),
    .A(net133),
    .B(net154));
 sg13g2_inv_1 _5294_ (.Y(_1553_),
    .A(_1552_));
 sg13g2_and2_1 _5295_ (.A(net222),
    .B(net202),
    .X(_1554_));
 sg13g2_mux2_1 _5296_ (.A0(_1554_),
    .A1(_1358_),
    .S(_0913_),
    .X(_1555_));
 sg13g2_nand2b_1 _5297_ (.Y(_1556_),
    .B(net226),
    .A_N(_1134_));
 sg13g2_nand2_1 _5298_ (.Y(_1557_),
    .A(net225),
    .B(_2742_));
 sg13g2_o21ai_1 _5299_ (.B1(_1557_),
    .Y(_1558_),
    .A1(_2558_),
    .A2(_1556_));
 sg13g2_or3_1 _5300_ (.A(_2777_),
    .B(_1555_),
    .C(_1558_),
    .X(_1559_));
 sg13g2_buf_1 _5301_ (.A(_1559_),
    .X(_1560_));
 sg13g2_o21ai_1 _5302_ (.B1(net174),
    .Y(_1561_),
    .A1(_1555_),
    .A2(_1558_));
 sg13g2_buf_1 _5303_ (.A(_1561_),
    .X(_1563_));
 sg13g2_and4_1 _5304_ (.A(_1553_),
    .B(_2965_),
    .C(_1560_),
    .D(_1563_),
    .X(_1564_));
 sg13g2_xnor2_1 _5305_ (.Y(_1565_),
    .A(net200),
    .B(_0548_));
 sg13g2_nor2_1 _5306_ (.A(_0121_),
    .B(_1565_),
    .Y(_1566_));
 sg13g2_nand2_1 _5307_ (.Y(_1567_),
    .A(_0120_),
    .B(_0249_));
 sg13g2_nand2_1 _5308_ (.Y(_1568_),
    .A(_0146_),
    .B(_1567_));
 sg13g2_and2_1 _5309_ (.A(_1566_),
    .B(_1568_),
    .X(_1569_));
 sg13g2_mux2_1 _5310_ (.A0(_1564_),
    .A1(_1569_),
    .S(net76),
    .X(_1570_));
 sg13g2_buf_1 _5311_ (.A(_1570_),
    .X(_1571_));
 sg13g2_o21ai_1 _5312_ (.B1(_1571_),
    .Y(_1572_),
    .A1(_1543_),
    .A2(_1550_));
 sg13g2_o21ai_1 _5313_ (.B1(_1572_),
    .Y(_1574_),
    .A1(_1361_),
    .A2(_1528_));
 sg13g2_nand2_1 _5314_ (.Y(_1575_),
    .A(_1414_),
    .B(_1423_));
 sg13g2_buf_1 _5315_ (.A(_1575_),
    .X(_1576_));
 sg13g2_nand2_1 _5316_ (.Y(_1577_),
    .A(_1379_),
    .B(_1390_));
 sg13g2_buf_1 _5317_ (.A(_1577_),
    .X(_1578_));
 sg13g2_nor2_1 _5318_ (.A(net39),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_nor3_1 _5319_ (.A(net28),
    .B(net122),
    .C(net25),
    .Y(_1580_));
 sg13g2_nand2_1 _5320_ (.Y(_1581_),
    .A(net125),
    .B(_1407_));
 sg13g2_buf_1 _5321_ (.A(_1581_),
    .X(_1582_));
 sg13g2_buf_1 _5322_ (.A(_1582_),
    .X(_1583_));
 sg13g2_o21ai_1 _5323_ (.B1(_1583_),
    .Y(_1585_),
    .A1(_1579_),
    .A2(_1580_));
 sg13g2_buf_1 _5324_ (.A(_1426_),
    .X(_1586_));
 sg13g2_o21ai_1 _5325_ (.B1(_1583_),
    .Y(_1587_),
    .A1(net103),
    .A2(net36));
 sg13g2_nand2_1 _5326_ (.Y(_1588_),
    .A(net27),
    .B(_1587_));
 sg13g2_buf_1 _5327_ (.A(_1410_),
    .X(_1589_));
 sg13g2_a21oi_1 _5328_ (.A1(_1536_),
    .A2(net71),
    .Y(_1590_),
    .B1(net37));
 sg13g2_nand3_1 _5329_ (.B(_0296_),
    .C(_1345_),
    .A(_2743_),
    .Y(_1591_));
 sg13g2_inv_1 _5330_ (.Y(_1592_),
    .A(_1591_));
 sg13g2_nor3_1 _5331_ (.A(_1322_),
    .B(_1342_),
    .C(_1557_),
    .Y(_1593_));
 sg13g2_nand3_1 _5332_ (.B(_1334_),
    .C(_1339_),
    .A(_1328_),
    .Y(_1594_));
 sg13g2_mux2_1 _5333_ (.A0(_1592_),
    .A1(_1593_),
    .S(_1594_),
    .X(_1596_));
 sg13g2_nor2_1 _5334_ (.A(_1345_),
    .B(_1557_),
    .Y(_1597_));
 sg13g2_nor4_1 _5335_ (.A(net177),
    .B(_0885_),
    .C(_1345_),
    .D(_1342_),
    .Y(_1598_));
 sg13g2_mux2_1 _5336_ (.A0(_1597_),
    .A1(_1598_),
    .S(_1594_),
    .X(_1599_));
 sg13g2_or2_1 _5337_ (.X(_1600_),
    .B(_1557_),
    .A(_1345_));
 sg13g2_or2_1 _5338_ (.X(_1601_),
    .B(_1341_),
    .A(_1325_));
 sg13g2_a21o_1 _5339_ (.A2(_1600_),
    .A1(_1591_),
    .B1(_1601_),
    .X(_1602_));
 sg13g2_o21ai_1 _5340_ (.B1(_1602_),
    .Y(_1603_),
    .A1(net177),
    .A2(_2760_));
 sg13g2_or3_1 _5341_ (.A(_1596_),
    .B(_1599_),
    .C(_1603_),
    .X(_1604_));
 sg13g2_buf_1 _5342_ (.A(_1604_),
    .X(_1605_));
 sg13g2_nor2_1 _5343_ (.A(_0547_),
    .B(_2794_),
    .Y(_1607_));
 sg13g2_and2_1 _5344_ (.A(_0814_),
    .B(_1506_),
    .X(_1608_));
 sg13g2_mux2_1 _5345_ (.A0(_1607_),
    .A1(_1608_),
    .S(net77),
    .X(_1609_));
 sg13g2_nand2_1 _5346_ (.Y(_1610_),
    .A(_1605_),
    .B(_1609_));
 sg13g2_a221oi_1 _5347_ (.B2(_1590_),
    .C1(_1610_),
    .B1(_1588_),
    .A1(net37),
    .Y(_1611_),
    .A2(_1585_));
 sg13g2_nor2_1 _5348_ (.A(net87),
    .B(_1470_),
    .Y(_1612_));
 sg13g2_nand2_1 _5349_ (.Y(_1613_),
    .A(net126),
    .B(_1426_));
 sg13g2_buf_1 _5350_ (.A(net146),
    .X(_1614_));
 sg13g2_nand2_1 _5351_ (.Y(_1615_),
    .A(net121),
    .B(net122));
 sg13g2_and4_1 _5352_ (.A(net144),
    .B(net87),
    .C(_1613_),
    .D(_1615_),
    .X(_1616_));
 sg13g2_nor2_1 _5353_ (.A(_1475_),
    .B(_1383_),
    .Y(_1617_));
 sg13g2_o21ai_1 _5354_ (.B1(_1617_),
    .Y(_1618_),
    .A1(_1612_),
    .A2(_1616_));
 sg13g2_mux2_1 _5355_ (.A0(_1475_),
    .A1(_1383_),
    .S(net126),
    .X(_1619_));
 sg13g2_and2_1 _5356_ (.A(net100),
    .B(net89),
    .X(_1620_));
 sg13g2_mux2_1 _5357_ (.A0(net90),
    .A1(net88),
    .S(net100),
    .X(_1621_));
 sg13g2_mux2_1 _5358_ (.A0(_1475_),
    .A1(_1383_),
    .S(_1472_),
    .X(_1622_));
 sg13g2_a22oi_1 _5359_ (.Y(_1623_),
    .B1(_1621_),
    .B2(_1622_),
    .A2(_1620_),
    .A1(_1619_));
 sg13g2_a21o_1 _5360_ (.A2(_1623_),
    .A1(_1618_),
    .B1(net39),
    .X(_1624_));
 sg13g2_o21ai_1 _5361_ (.B1(_1537_),
    .Y(_1625_),
    .A1(net104),
    .A2(net147));
 sg13g2_nand4_1 _5362_ (.B(net123),
    .C(net126),
    .A(net105),
    .Y(_1626_),
    .D(net103));
 sg13g2_o21ai_1 _5363_ (.B1(_1626_),
    .Y(_1628_),
    .A1(net126),
    .A2(_1625_));
 sg13g2_nor3_1 _5364_ (.A(_1420_),
    .B(_1421_),
    .C(_1426_),
    .Y(_1629_));
 sg13g2_a21oi_1 _5365_ (.A1(net105),
    .A2(net123),
    .Y(_1630_),
    .B1(_1537_));
 sg13g2_or2_1 _5366_ (.X(_1631_),
    .B(_1630_),
    .A(_1629_));
 sg13g2_o21ai_1 _5367_ (.B1(_1477_),
    .Y(_1632_),
    .A1(_1336_),
    .A2(net121));
 sg13g2_a22oi_1 _5368_ (.Y(_1633_),
    .B1(_1631_),
    .B2(_1632_),
    .A2(_1628_),
    .A1(net148));
 sg13g2_or3_1 _5369_ (.A(net28),
    .B(net87),
    .C(_1633_),
    .X(_1634_));
 sg13g2_nand2b_1 _5370_ (.Y(_1635_),
    .B(_1356_),
    .A_N(_0146_));
 sg13g2_buf_1 _5371_ (.A(_1635_),
    .X(_1636_));
 sg13g2_mux2_1 _5372_ (.A0(_1552_),
    .A1(_1567_),
    .S(_1356_),
    .X(_1637_));
 sg13g2_buf_1 _5373_ (.A(_1637_),
    .X(_1639_));
 sg13g2_a21o_1 _5374_ (.A2(_1639_),
    .A1(_1636_),
    .B1(_1526_),
    .X(_1640_));
 sg13g2_buf_1 _5375_ (.A(_1640_),
    .X(_1641_));
 sg13g2_a21oi_1 _5376_ (.A1(_1624_),
    .A2(_1634_),
    .Y(_1642_),
    .B1(_1641_));
 sg13g2_nand2_1 _5377_ (.Y(_1643_),
    .A(net71),
    .B(net75));
 sg13g2_nand2b_1 _5378_ (.Y(_1644_),
    .B(_1490_),
    .A_N(_1643_));
 sg13g2_nor2_1 _5379_ (.A(_1418_),
    .B(net147),
    .Y(_1645_));
 sg13g2_buf_2 _5380_ (.A(_1645_),
    .X(_1646_));
 sg13g2_nand2_1 _5381_ (.Y(_1647_),
    .A(net185),
    .B(net149));
 sg13g2_a21oi_1 _5382_ (.A1(net127),
    .A2(_1385_),
    .Y(_1648_),
    .B1(_1647_));
 sg13g2_and4_1 _5383_ (.A(_1437_),
    .B(_1439_),
    .C(net149),
    .D(_1498_),
    .X(_1650_));
 sg13g2_a221oi_1 _5384_ (.B2(_1469_),
    .C1(_1650_),
    .B1(_1648_),
    .A1(_1646_),
    .Y(_1651_),
    .A2(_1371_));
 sg13g2_buf_1 _5385_ (.A(_1651_),
    .X(_1652_));
 sg13g2_nand2_1 _5386_ (.Y(_1653_),
    .A(_1515_),
    .B(net56));
 sg13g2_nand2_1 _5387_ (.Y(_1654_),
    .A(_2721_),
    .B(net146));
 sg13g2_a21oi_1 _5388_ (.A1(net127),
    .A2(_1385_),
    .Y(_1655_),
    .B1(_1654_));
 sg13g2_nor2_1 _5389_ (.A(net137),
    .B(net149),
    .Y(_1656_));
 sg13g2_nand2_1 _5390_ (.Y(_1657_),
    .A(net149),
    .B(_1327_));
 sg13g2_a21oi_1 _5391_ (.A1(net105),
    .A2(net123),
    .Y(_1658_),
    .B1(_1657_));
 sg13g2_a221oi_1 _5392_ (.B2(_1475_),
    .C1(_1658_),
    .B1(_1656_),
    .A1(_1469_),
    .Y(_1659_),
    .A2(_1655_));
 sg13g2_buf_1 _5393_ (.A(_1659_),
    .X(_1661_));
 sg13g2_buf_1 _5394_ (.A(net88),
    .X(_1662_));
 sg13g2_nand2_1 _5395_ (.Y(_1663_),
    .A(net55),
    .B(net70));
 sg13g2_nand3_1 _5396_ (.B(_1653_),
    .C(_1663_),
    .A(_1464_),
    .Y(_1664_));
 sg13g2_nor2_1 _5397_ (.A(net154),
    .B(_0918_),
    .Y(_1665_));
 sg13g2_nand2_1 _5398_ (.Y(_1666_),
    .A(_1566_),
    .B(_1665_));
 sg13g2_and2_1 _5399_ (.A(net201),
    .B(_0286_),
    .X(_1667_));
 sg13g2_nand4_1 _5400_ (.B(_1560_),
    .C(_1563_),
    .A(net177),
    .Y(_1668_),
    .D(_1667_));
 sg13g2_mux2_1 _5401_ (.A0(_1666_),
    .A1(_1668_),
    .S(net77),
    .X(_1669_));
 sg13g2_buf_1 _5402_ (.A(_1669_),
    .X(_1670_));
 sg13g2_a21oi_1 _5403_ (.A1(_1644_),
    .A2(_1664_),
    .Y(_1672_),
    .B1(_1670_));
 sg13g2_nand2b_1 _5404_ (.Y(_1673_),
    .B(_1605_),
    .A_N(_1510_));
 sg13g2_buf_2 _5405_ (.A(_1673_),
    .X(_1674_));
 sg13g2_nor2_2 _5406_ (.A(_1395_),
    .B(_1398_),
    .Y(_1675_));
 sg13g2_o21ai_1 _5407_ (.B1(_1581_),
    .Y(_1676_),
    .A1(_1395_),
    .A2(_1398_));
 sg13g2_buf_1 _5408_ (.A(_1676_),
    .X(_1677_));
 sg13g2_nand3_1 _5409_ (.B(_1414_),
    .C(_1423_),
    .A(_1467_),
    .Y(_1678_));
 sg13g2_and2_1 _5410_ (.A(_1677_),
    .B(_1678_),
    .X(_1679_));
 sg13g2_a221oi_1 _5411_ (.B2(net36),
    .C1(net28),
    .B1(_1679_),
    .A1(_1675_),
    .Y(_1680_),
    .A2(net70));
 sg13g2_and4_1 _5412_ (.A(_1493_),
    .B(_1497_),
    .C(_1499_),
    .D(_1501_),
    .X(_1681_));
 sg13g2_buf_1 _5413_ (.A(_1681_),
    .X(_1683_));
 sg13g2_nor2_2 _5414_ (.A(net87),
    .B(_1683_),
    .Y(_1684_));
 sg13g2_nor2_1 _5415_ (.A(_1489_),
    .B(_1684_),
    .Y(_1685_));
 sg13g2_nor3_1 _5416_ (.A(_1674_),
    .B(_1680_),
    .C(_1685_),
    .Y(_1686_));
 sg13g2_or3_1 _5417_ (.A(_1642_),
    .B(_1672_),
    .C(_1686_),
    .X(_1687_));
 sg13g2_nor2b_1 _5418_ (.A(_1565_),
    .B_N(_2965_),
    .Y(_1688_));
 sg13g2_nand2_1 _5419_ (.Y(_1689_),
    .A(_1688_),
    .B(_1665_));
 sg13g2_nand4_1 _5420_ (.B(net177),
    .C(_0116_),
    .A(_2610_),
    .Y(_1690_),
    .D(_2839_));
 sg13g2_mux2_1 _5421_ (.A0(_1689_),
    .A1(_1690_),
    .S(net77),
    .X(_1691_));
 sg13g2_or2_1 _5422_ (.X(_1692_),
    .B(_1691_),
    .A(net71));
 sg13g2_buf_1 _5423_ (.A(_1692_),
    .X(_1694_));
 sg13g2_nor2_1 _5424_ (.A(net40),
    .B(net56),
    .Y(_1695_));
 sg13g2_nor2b_1 _5425_ (.A(_1694_),
    .B_N(_1695_),
    .Y(_1696_));
 sg13g2_nand2_1 _5426_ (.Y(_1697_),
    .A(_0195_),
    .B(net177));
 sg13g2_nand2_1 _5427_ (.Y(_1698_),
    .A(net177),
    .B(_0249_));
 sg13g2_mux2_1 _5428_ (.A0(_1697_),
    .A1(_1698_),
    .S(_1356_),
    .X(_1699_));
 sg13g2_buf_1 _5429_ (.A(_1699_),
    .X(_1700_));
 sg13g2_nand3_1 _5430_ (.B(_2768_),
    .C(net76),
    .A(_0120_),
    .Y(_1701_));
 sg13g2_buf_2 _5431_ (.A(_1701_),
    .X(_1702_));
 sg13g2_a22oi_1 _5432_ (.Y(_1703_),
    .B1(_1542_),
    .B2(_1678_),
    .A2(_1390_),
    .A1(_1379_));
 sg13g2_nand3_1 _5433_ (.B(_1609_),
    .C(_1703_),
    .A(net22),
    .Y(_1705_));
 sg13g2_nand2b_1 _5434_ (.Y(_1706_),
    .B(_2965_),
    .A_N(_1565_));
 sg13g2_nand3_1 _5435_ (.B(_1560_),
    .C(_1563_),
    .A(_2839_),
    .Y(_1707_));
 sg13g2_mux2_1 _5436_ (.A0(_1706_),
    .A1(_1707_),
    .S(net77),
    .X(_1708_));
 sg13g2_buf_1 _5437_ (.A(_1708_),
    .X(_1709_));
 sg13g2_and3_1 _5438_ (.X(_1710_),
    .A(_1437_),
    .B(_1439_),
    .C(_1327_));
 sg13g2_buf_1 _5439_ (.A(_1710_),
    .X(_1711_));
 sg13g2_nor4_1 _5440_ (.A(_2534_),
    .B(_2537_),
    .C(_0447_),
    .D(_1449_),
    .Y(_1712_));
 sg13g2_o21ai_1 _5441_ (.B1(_1712_),
    .Y(_1713_),
    .A1(net104),
    .A2(net147));
 sg13g2_nor2_1 _5442_ (.A(net149),
    .B(_1449_),
    .Y(_1714_));
 sg13g2_nand4_1 _5443_ (.B(net123),
    .C(_1498_),
    .A(net105),
    .Y(_1716_),
    .D(_1714_));
 sg13g2_nor3_1 _5444_ (.A(net149),
    .B(_1449_),
    .C(_1494_),
    .Y(_1717_));
 sg13g2_nand3_1 _5445_ (.B(net123),
    .C(_1717_),
    .A(net105),
    .Y(_1718_));
 sg13g2_nand4_1 _5446_ (.B(_1437_),
    .C(_1439_),
    .A(_1500_),
    .Y(_1719_),
    .D(_1714_));
 sg13g2_nand4_1 _5447_ (.B(_1716_),
    .C(_1718_),
    .A(_1713_),
    .Y(_1720_),
    .D(_1719_));
 sg13g2_a21oi_1 _5448_ (.A1(_1447_),
    .A2(_1711_),
    .Y(_1721_),
    .B1(_1720_));
 sg13g2_buf_2 _5449_ (.A(_1721_),
    .X(_1722_));
 sg13g2_or3_1 _5450_ (.A(net35),
    .B(net71),
    .C(_1722_),
    .X(_1723_));
 sg13g2_a22oi_1 _5451_ (.Y(_1724_),
    .B1(_1705_),
    .B2(_1723_),
    .A2(_1702_),
    .A1(_1700_));
 sg13g2_inv_1 _5452_ (.Y(_1725_),
    .A(_0145_));
 sg13g2_nand3_1 _5453_ (.B(_1725_),
    .C(net77),
    .A(_0547_),
    .Y(_1727_));
 sg13g2_o21ai_1 _5454_ (.B1(net174),
    .Y(_1728_),
    .A1(_0145_),
    .A2(net76));
 sg13g2_nand4_1 _5455_ (.B(_1605_),
    .C(_1727_),
    .A(_0876_),
    .Y(_1729_),
    .D(_1728_));
 sg13g2_xnor2_1 _5456_ (.Y(_1730_),
    .A(_0326_),
    .B(net76));
 sg13g2_o21ai_1 _5457_ (.B1(net72),
    .Y(_1731_),
    .A1(net103),
    .A2(_1730_));
 sg13g2_nor3_1 _5458_ (.A(_1729_),
    .B(_1722_),
    .C(_1731_),
    .Y(_1732_));
 sg13g2_or3_1 _5459_ (.A(_1696_),
    .B(_1724_),
    .C(_1732_),
    .X(_1733_));
 sg13g2_nor4_1 _5460_ (.A(_1574_),
    .B(_1611_),
    .C(_1687_),
    .D(_1733_),
    .Y(_1734_));
 sg13g2_nand2_1 _5461_ (.Y(_1735_),
    .A(net105),
    .B(net123));
 sg13g2_buf_1 _5462_ (.A(_1735_),
    .X(_1736_));
 sg13g2_xnor2_1 _5463_ (.Y(_1738_),
    .A(net69),
    .B(net88));
 sg13g2_nand2_1 _5464_ (.Y(_1739_),
    .A(_1632_),
    .B(_1738_));
 sg13g2_buf_1 _5465_ (.A(net126),
    .X(_1740_));
 sg13g2_nand4_1 _5466_ (.B(net102),
    .C(net148),
    .A(_1646_),
    .Y(_1741_),
    .D(net70));
 sg13g2_nand4_1 _5467_ (.B(net121),
    .C(net148),
    .A(net69),
    .Y(_1742_),
    .D(net73));
 sg13g2_nand4_1 _5468_ (.B(_1739_),
    .C(_1741_),
    .A(_1412_),
    .Y(_1743_),
    .D(_1742_));
 sg13g2_nor2b_1 _5469_ (.A(net35),
    .B_N(_1743_),
    .Y(_1744_));
 sg13g2_o21ai_1 _5470_ (.B1(_1412_),
    .Y(_1745_),
    .A1(_1484_),
    .A2(_1487_));
 sg13g2_nand3_1 _5471_ (.B(_1423_),
    .C(net71),
    .A(_1414_),
    .Y(_1746_));
 sg13g2_nand4_1 _5472_ (.B(_1460_),
    .C(_1677_),
    .A(_1455_),
    .Y(_1747_),
    .D(_1746_));
 sg13g2_nand3_1 _5473_ (.B(_1745_),
    .C(_1747_),
    .A(_1536_),
    .Y(_1749_));
 sg13g2_nor2_1 _5474_ (.A(_1410_),
    .B(net88),
    .Y(_1750_));
 sg13g2_nand2b_1 _5475_ (.Y(_1751_),
    .B(_1750_),
    .A_N(_1651_));
 sg13g2_nand2b_1 _5476_ (.Y(_1752_),
    .B(_1750_),
    .A_N(net38));
 sg13g2_mux2_1 _5477_ (.A0(_1751_),
    .A1(_1752_),
    .S(net22),
    .X(_1753_));
 sg13g2_and3_1 _5478_ (.X(_1754_),
    .A(_2965_),
    .B(_1560_),
    .C(_1563_));
 sg13g2_mux2_1 _5479_ (.A0(_1566_),
    .A1(_1754_),
    .S(_1351_),
    .X(_1755_));
 sg13g2_buf_1 _5480_ (.A(_1755_),
    .X(_1756_));
 sg13g2_inv_1 _5481_ (.Y(_1757_),
    .A(_1756_));
 sg13g2_a21oi_1 _5482_ (.A1(_1749_),
    .A2(_1753_),
    .Y(_1758_),
    .B1(_1757_));
 sg13g2_o21ai_1 _5483_ (.B1(_1605_),
    .Y(_1760_),
    .A1(_1744_),
    .A2(_1758_));
 sg13g2_nand2_1 _5484_ (.Y(_1761_),
    .A(net121),
    .B(net103));
 sg13g2_o21ai_1 _5485_ (.B1(_1761_),
    .Y(_1762_),
    .A1(net121),
    .A2(net74));
 sg13g2_nand2_1 _5486_ (.Y(_1763_),
    .A(_1711_),
    .B(_1762_));
 sg13g2_o21ai_1 _5487_ (.B1(net81),
    .Y(_1764_),
    .A1(_1475_),
    .A2(_1383_));
 sg13g2_o21ai_1 _5488_ (.B1(_1613_),
    .Y(_1765_),
    .A1(net102),
    .A2(net74));
 sg13g2_nand3_1 _5489_ (.B(_1764_),
    .C(_1765_),
    .A(_1530_),
    .Y(_1766_));
 sg13g2_nand3_1 _5490_ (.B(_1763_),
    .C(_1766_),
    .A(_1482_),
    .Y(_1767_));
 sg13g2_nor2_1 _5491_ (.A(net27),
    .B(net35),
    .Y(_1768_));
 sg13g2_nand3_1 _5492_ (.B(_1460_),
    .C(_1503_),
    .A(_1455_),
    .Y(_1769_));
 sg13g2_buf_1 _5493_ (.A(_1769_),
    .X(_1771_));
 sg13g2_nor3_1 _5494_ (.A(_1709_),
    .B(net73),
    .C(_1771_),
    .Y(_1772_));
 sg13g2_a21o_1 _5495_ (.A2(_1768_),
    .A1(_1767_),
    .B1(_1772_),
    .X(_1773_));
 sg13g2_nand2_2 _5496_ (.Y(_1774_),
    .A(_1426_),
    .B(_1467_));
 sg13g2_nor2_1 _5497_ (.A(_1774_),
    .B(net56),
    .Y(_1775_));
 sg13g2_nor2_1 _5498_ (.A(_1545_),
    .B(_1480_),
    .Y(_1776_));
 sg13g2_buf_1 _5499_ (.A(net90),
    .X(_1777_));
 sg13g2_nor2_1 _5500_ (.A(net68),
    .B(_1683_),
    .Y(_1778_));
 sg13g2_nor4_1 _5501_ (.A(net27),
    .B(_1775_),
    .C(_1776_),
    .D(_1778_),
    .Y(_1779_));
 sg13g2_nand2_2 _5502_ (.Y(_1780_),
    .A(net122),
    .B(net87));
 sg13g2_nor2_1 _5503_ (.A(_1780_),
    .B(net38),
    .Y(_1782_));
 sg13g2_nor3_1 _5504_ (.A(net22),
    .B(_1684_),
    .C(_1782_),
    .Y(_1783_));
 sg13g2_nor3_1 _5505_ (.A(net26),
    .B(_1779_),
    .C(_1783_),
    .Y(_1784_));
 sg13g2_nand2_1 _5506_ (.Y(_1785_),
    .A(_1636_),
    .B(_1639_));
 sg13g2_o21ai_1 _5507_ (.B1(_1785_),
    .Y(_1786_),
    .A1(_1773_),
    .A2(_1784_));
 sg13g2_nor3_1 _5508_ (.A(net68),
    .B(net26),
    .C(net56),
    .Y(_1787_));
 sg13g2_o21ai_1 _5509_ (.B1(_1756_),
    .Y(_1788_),
    .A1(net122),
    .A2(net68));
 sg13g2_nand2b_1 _5510_ (.Y(_1789_),
    .B(net71),
    .A_N(net26));
 sg13g2_a21oi_1 _5511_ (.A1(_1788_),
    .A2(_1789_),
    .Y(_1790_),
    .B1(net55));
 sg13g2_buf_1 _5512_ (.A(net27),
    .X(_1791_));
 sg13g2_a21oi_1 _5513_ (.A1(_1700_),
    .A2(_1702_),
    .Y(_1793_),
    .B1(net21));
 sg13g2_o21ai_1 _5514_ (.B1(_1793_),
    .Y(_1794_),
    .A1(_1787_),
    .A2(_1790_));
 sg13g2_and3_1 _5515_ (.X(_1795_),
    .A(_1760_),
    .B(_1786_),
    .C(_1794_));
 sg13g2_and2_1 _5516_ (.A(_1734_),
    .B(_1795_),
    .X(_1796_));
 sg13g2_nand3_1 _5517_ (.B(_2576_),
    .C(net6),
    .A(net231),
    .Y(_1797_));
 sg13g2_buf_1 _5518_ (.A(_1797_),
    .X(_1798_));
 sg13g2_nand2b_1 _5519_ (.Y(_1799_),
    .B(_1785_),
    .A_N(_1511_));
 sg13g2_nor2_1 _5520_ (.A(net103),
    .B(net37),
    .Y(_1800_));
 sg13g2_o21ai_1 _5521_ (.B1(net148),
    .Y(_1801_),
    .A1(_1646_),
    .A2(net91));
 sg13g2_nor3_1 _5522_ (.A(_2898_),
    .B(net104),
    .C(net147),
    .Y(_1802_));
 sg13g2_a221oi_1 _5523_ (.B2(_1802_),
    .C1(net121),
    .B1(net91),
    .A1(_1500_),
    .Y(_1804_),
    .A2(net69));
 sg13g2_nor3_1 _5524_ (.A(_1336_),
    .B(net104),
    .C(net147),
    .Y(_1805_));
 sg13g2_a221oi_1 _5525_ (.B2(_1805_),
    .C1(_1740_),
    .B1(net91),
    .A1(net144),
    .Y(_1806_),
    .A2(_1383_));
 sg13g2_a21oi_1 _5526_ (.A1(_1801_),
    .A2(_1804_),
    .Y(_1807_),
    .B1(_1806_));
 sg13g2_o21ai_1 _5527_ (.B1(_1807_),
    .Y(_1808_),
    .A1(_1465_),
    .A2(_1800_));
 sg13g2_nand2_1 _5528_ (.Y(_1809_),
    .A(net103),
    .B(net37));
 sg13g2_nand4_1 _5529_ (.B(_1460_),
    .C(_1379_),
    .A(_1455_),
    .Y(_1810_),
    .D(_1390_));
 sg13g2_a21o_1 _5530_ (.A2(_1809_),
    .A1(_1780_),
    .B1(_1810_),
    .X(_1811_));
 sg13g2_and2_1 _5531_ (.A(_1808_),
    .B(_1811_),
    .X(_1812_));
 sg13g2_nor2_1 _5532_ (.A(_1799_),
    .B(_1812_),
    .Y(_1813_));
 sg13g2_a21oi_2 _5533_ (.B1(_1722_),
    .Y(_1815_),
    .A2(_1702_),
    .A1(_1700_));
 sg13g2_nand2_1 _5534_ (.Y(_1816_),
    .A(net28),
    .B(_1684_));
 sg13g2_nand4_1 _5535_ (.B(net36),
    .C(_1412_),
    .A(net39),
    .Y(_1817_),
    .D(_1429_));
 sg13g2_nor3_2 _5536_ (.A(_1596_),
    .B(_1599_),
    .C(_1603_),
    .Y(_1818_));
 sg13g2_a21oi_1 _5537_ (.A1(_1816_),
    .A2(_1817_),
    .Y(_1819_),
    .B1(_1818_));
 sg13g2_a21o_1 _5538_ (.A2(_1702_),
    .A1(_1700_),
    .B1(_1722_),
    .X(_1820_));
 sg13g2_nand2_1 _5539_ (.Y(_1821_),
    .A(_1756_),
    .B(net72));
 sg13g2_o21ai_1 _5540_ (.B1(net26),
    .Y(_1822_),
    .A1(_1820_),
    .A2(_1821_));
 sg13g2_o21ai_1 _5541_ (.B1(_1822_),
    .Y(_1823_),
    .A1(_1815_),
    .A2(_1819_));
 sg13g2_a21oi_2 _5542_ (.B1(_1526_),
    .Y(_1824_),
    .A2(_1360_),
    .A1(_1354_));
 sg13g2_nand2_1 _5543_ (.Y(_1826_),
    .A(_1462_),
    .B(_1577_));
 sg13g2_a21oi_1 _5544_ (.A1(net37),
    .A2(net74),
    .Y(_1827_),
    .B1(_1800_));
 sg13g2_nand2b_1 _5545_ (.Y(_1828_),
    .B(_1428_),
    .A_N(_1771_));
 sg13g2_o21ai_1 _5546_ (.B1(_1828_),
    .Y(_1829_),
    .A1(_1826_),
    .A2(_1827_));
 sg13g2_a21oi_1 _5547_ (.A1(_1636_),
    .A2(_1639_),
    .Y(_1830_),
    .B1(net35));
 sg13g2_o21ai_1 _5548_ (.B1(net40),
    .Y(_1831_),
    .A1(net89),
    .A2(_1683_));
 sg13g2_and2_1 _5549_ (.A(_1830_),
    .B(_1831_),
    .X(_1832_));
 sg13g2_mux2_1 _5550_ (.A0(_1383_),
    .A1(_1617_),
    .S(_2566_),
    .X(_1833_));
 sg13g2_a221oi_1 _5551_ (.B2(_1833_),
    .C1(_1614_),
    .B1(_1515_),
    .A1(_1327_),
    .Y(_1834_),
    .A2(_1589_));
 sg13g2_a21oi_1 _5552_ (.A1(_1646_),
    .A2(_1515_),
    .Y(_1835_),
    .B1(_1410_));
 sg13g2_nand2_1 _5553_ (.Y(_1837_),
    .A(_1646_),
    .B(_1410_));
 sg13g2_o21ai_1 _5554_ (.B1(_1837_),
    .Y(_1838_),
    .A1(net166),
    .A2(_1835_));
 sg13g2_a221oi_1 _5555_ (.B2(net81),
    .C1(_1740_),
    .B1(_1838_),
    .A1(_1475_),
    .Y(_1839_),
    .A2(_1589_));
 sg13g2_nor2_1 _5556_ (.A(net39),
    .B(_1516_),
    .Y(_1840_));
 sg13g2_o21ai_1 _5557_ (.B1(_1840_),
    .Y(_1841_),
    .A1(_1834_),
    .A2(_1839_));
 sg13g2_inv_1 _5558_ (.Y(_1842_),
    .A(_1571_));
 sg13g2_nor2_1 _5559_ (.A(net88),
    .B(_1683_),
    .Y(_1843_));
 sg13g2_nor3_1 _5560_ (.A(net28),
    .B(_1843_),
    .C(_1776_),
    .Y(_1844_));
 sg13g2_nor2_1 _5561_ (.A(_1777_),
    .B(_1480_),
    .Y(_1845_));
 sg13g2_nor2_1 _5562_ (.A(net89),
    .B(net56),
    .Y(_1846_));
 sg13g2_nor3_1 _5563_ (.A(net39),
    .B(_1845_),
    .C(_1846_),
    .Y(_1848_));
 sg13g2_nor3_1 _5564_ (.A(_1842_),
    .B(_1844_),
    .C(_1848_),
    .Y(_1849_));
 sg13g2_a221oi_1 _5565_ (.B2(_1841_),
    .C1(_1849_),
    .B1(_1832_),
    .A1(_1824_),
    .Y(_1850_),
    .A2(_1829_));
 sg13g2_a221oi_1 _5566_ (.B2(_1500_),
    .C1(net126),
    .B1(_1629_),
    .A1(net87),
    .Y(_1851_),
    .A2(_1711_));
 sg13g2_and4_1 _5567_ (.A(_1413_),
    .B(_1476_),
    .C(net125),
    .D(net124),
    .X(_1852_));
 sg13g2_nor3_1 _5568_ (.A(_1396_),
    .B(_1852_),
    .C(_1630_),
    .Y(_1853_));
 sg13g2_a21oi_1 _5569_ (.A1(_1413_),
    .A2(_1476_),
    .Y(_1854_),
    .B1(_1336_));
 sg13g2_a22oi_1 _5570_ (.Y(_1855_),
    .B1(_1629_),
    .B2(_1327_),
    .A2(_1854_),
    .A1(net87));
 sg13g2_nand3b_1 _5571_ (.B(_1855_),
    .C(net126),
    .Y(_1856_),
    .A_N(_1853_));
 sg13g2_nand3b_1 _5572_ (.B(_1462_),
    .C(_1856_),
    .Y(_1857_),
    .A_N(_1851_));
 sg13g2_nor2_1 _5573_ (.A(_1480_),
    .B(_1774_),
    .Y(_1859_));
 sg13g2_a21oi_1 _5574_ (.A1(net40),
    .A2(net75),
    .Y(_1860_),
    .B1(_1859_));
 sg13g2_a21o_1 _5575_ (.A2(_1860_),
    .A1(_1857_),
    .B1(_1641_),
    .X(_1861_));
 sg13g2_nor2_1 _5576_ (.A(_1586_),
    .B(_1771_),
    .Y(_1862_));
 sg13g2_o21ai_1 _5577_ (.B1(_1652_),
    .Y(_1863_),
    .A1(_1661_),
    .A2(_1774_));
 sg13g2_and2_1 _5578_ (.A(_1462_),
    .B(_1863_),
    .X(_1864_));
 sg13g2_a21oi_2 _5579_ (.B1(_1510_),
    .Y(_1865_),
    .A2(_1360_),
    .A1(_1354_));
 sg13g2_o21ai_1 _5580_ (.B1(_1865_),
    .Y(_1866_),
    .A1(_1862_),
    .A2(_1864_));
 sg13g2_nor2_1 _5581_ (.A(_1818_),
    .B(net35),
    .Y(_1867_));
 sg13g2_nand3_1 _5582_ (.B(net90),
    .C(_1622_),
    .A(net81),
    .Y(_1868_));
 sg13g2_nand2_1 _5583_ (.Y(_1870_),
    .A(net144),
    .B(net89));
 sg13g2_a22oi_1 _5584_ (.Y(_1871_),
    .B1(_1492_),
    .B2(_2898_),
    .A2(_1656_),
    .A1(net90));
 sg13g2_mux2_1 _5585_ (.A0(_1870_),
    .A1(_1871_),
    .S(_1617_),
    .X(_1872_));
 sg13g2_nand3_1 _5586_ (.B(_1534_),
    .C(_1412_),
    .A(_1532_),
    .Y(_1873_));
 sg13g2_and3_1 _5587_ (.X(_1874_),
    .A(_1868_),
    .B(_1872_),
    .C(_1873_));
 sg13g2_nand3_1 _5588_ (.B(_1423_),
    .C(_1515_),
    .A(_1414_),
    .Y(_1875_));
 sg13g2_buf_1 _5589_ (.A(_1875_),
    .X(_1876_));
 sg13g2_and2_1 _5590_ (.A(_1542_),
    .B(_1876_),
    .X(_1877_));
 sg13g2_nor4_1 _5591_ (.A(net40),
    .B(_1535_),
    .C(_1691_),
    .D(_1877_),
    .Y(_1878_));
 sg13g2_a21oi_1 _5592_ (.A1(_1867_),
    .A2(_1874_),
    .Y(_1879_),
    .B1(_1878_));
 sg13g2_a21oi_1 _5593_ (.A1(net40),
    .A2(_1643_),
    .Y(_1881_),
    .B1(_1670_));
 sg13g2_a22oi_1 _5594_ (.Y(_1882_),
    .B1(_1677_),
    .B2(_1678_),
    .A2(_1390_),
    .A1(_1379_));
 sg13g2_nor2_1 _5595_ (.A(_1661_),
    .B(_1515_),
    .Y(_1883_));
 sg13g2_or3_1 _5596_ (.A(_1488_),
    .B(_1882_),
    .C(_1883_),
    .X(_1884_));
 sg13g2_a22oi_1 _5597_ (.Y(_1885_),
    .B1(_1607_),
    .B2(_1545_),
    .A2(net88),
    .A1(_1688_));
 sg13g2_and3_1 _5598_ (.X(_1886_),
    .A(_2839_),
    .B(_1560_),
    .C(_1563_));
 sg13g2_a221oi_1 _5599_ (.B2(_1545_),
    .C1(net76),
    .B1(_1608_),
    .A1(_1886_),
    .Y(_1887_),
    .A2(net88));
 sg13g2_a21oi_1 _5600_ (.A1(net76),
    .A2(_1885_),
    .Y(_1888_),
    .B1(_1887_));
 sg13g2_a22oi_1 _5601_ (.Y(_1889_),
    .B1(_1888_),
    .B2(_1815_),
    .A2(_1884_),
    .A1(_1881_));
 sg13g2_and4_1 _5602_ (.A(_1861_),
    .B(_1866_),
    .C(_1879_),
    .D(_1889_),
    .X(_1890_));
 sg13g2_nand4_1 _5603_ (.B(_1560_),
    .C(_1563_),
    .A(net77),
    .Y(_1892_),
    .D(_1667_));
 sg13g2_nand3_1 _5604_ (.B(net76),
    .C(_1566_),
    .A(_0887_),
    .Y(_1893_));
 sg13g2_a21oi_2 _5605_ (.B1(_2785_),
    .Y(_1894_),
    .A2(_1893_),
    .A1(_1892_));
 sg13g2_a21oi_1 _5606_ (.A1(_1455_),
    .A2(_1460_),
    .Y(_1895_),
    .B1(_1503_));
 sg13g2_and3_1 _5607_ (.X(_1896_),
    .A(net40),
    .B(net38),
    .C(_1751_));
 sg13g2_o21ai_1 _5608_ (.B1(_1752_),
    .Y(_1897_),
    .A1(_1895_),
    .A2(_1896_));
 sg13g2_a221oi_1 _5609_ (.B2(_1500_),
    .C1(_1388_),
    .B1(_1852_),
    .A1(_1581_),
    .Y(_1898_),
    .A2(_1711_));
 sg13g2_nor4_1 _5610_ (.A(_1736_),
    .B(_1614_),
    .C(net90),
    .D(net148),
    .Y(_1899_));
 sg13g2_nor4_1 _5611_ (.A(_1646_),
    .B(net121),
    .C(net87),
    .D(_1392_),
    .Y(_1900_));
 sg13g2_a221oi_1 _5612_ (.B2(net123),
    .C1(net146),
    .B1(net105),
    .A1(_2897_),
    .Y(_1901_),
    .A2(net187));
 sg13g2_nor4_1 _5613_ (.A(_1420_),
    .B(_1421_),
    .C(net146),
    .D(_1327_),
    .Y(_1903_));
 sg13g2_mux2_1 _5614_ (.A0(_1901_),
    .A1(_1903_),
    .S(net90),
    .X(_1904_));
 sg13g2_nor4_1 _5615_ (.A(_1898_),
    .B(_1899_),
    .C(_1900_),
    .D(_1904_),
    .Y(_1905_));
 sg13g2_o21ai_1 _5616_ (.B1(_1513_),
    .Y(_1906_),
    .A1(_1905_),
    .A2(_1703_));
 sg13g2_nand2_1 _5617_ (.Y(_1907_),
    .A(_1677_),
    .B(_1546_));
 sg13g2_nand3_1 _5618_ (.B(net25),
    .C(_1907_),
    .A(net28),
    .Y(_1908_));
 sg13g2_a21oi_1 _5619_ (.A1(_1906_),
    .A2(_1908_),
    .Y(_1909_),
    .B1(_1610_));
 sg13g2_a21oi_1 _5620_ (.A1(_1894_),
    .A2(_1897_),
    .Y(_1910_),
    .B1(_1909_));
 sg13g2_nand4_1 _5621_ (.B(_1850_),
    .C(_1890_),
    .A(_1823_),
    .Y(_1911_),
    .D(_1910_));
 sg13g2_buf_1 _5622_ (.A(_1911_),
    .X(_1912_));
 sg13g2_or3_1 _5623_ (.A(_1462_),
    .B(net36),
    .C(_1679_),
    .X(_1914_));
 sg13g2_nand2_1 _5624_ (.Y(_1915_),
    .A(_1539_),
    .B(_1480_));
 sg13g2_nand3_1 _5625_ (.B(_1653_),
    .C(_1915_),
    .A(_1464_),
    .Y(_1916_));
 sg13g2_a21o_1 _5626_ (.A2(_1916_),
    .A1(_1914_),
    .B1(_1641_),
    .X(_1917_));
 sg13g2_xnor2_1 _5627_ (.Y(_1918_),
    .A(_1675_),
    .B(_1410_));
 sg13g2_and3_1 _5628_ (.X(_1919_),
    .A(net40),
    .B(_1535_),
    .C(_1918_));
 sg13g2_o21ai_1 _5629_ (.B1(_1571_),
    .Y(_1920_),
    .A1(_1695_),
    .A2(_1919_));
 sg13g2_a22oi_1 _5630_ (.Y(_1921_),
    .B1(_1675_),
    .B2(_1586_),
    .A2(_1534_),
    .A1(_1532_));
 sg13g2_mux2_1 _5631_ (.A0(_1578_),
    .A1(_1921_),
    .S(_1462_),
    .X(_1922_));
 sg13g2_nor2_1 _5632_ (.A(_1777_),
    .B(net37),
    .Y(_1923_));
 sg13g2_nor3_1 _5633_ (.A(_1818_),
    .B(_1526_),
    .C(_1923_),
    .Y(_1925_));
 sg13g2_a21oi_1 _5634_ (.A1(_1636_),
    .A2(_1639_),
    .Y(_1926_),
    .B1(_1510_));
 sg13g2_a22oi_1 _5635_ (.Y(_1927_),
    .B1(_1542_),
    .B2(_1876_),
    .A2(_1534_),
    .A1(_1532_));
 sg13g2_mux2_1 _5636_ (.A0(_1927_),
    .A1(_1905_),
    .S(net28),
    .X(_1928_));
 sg13g2_a22oi_1 _5637_ (.Y(_1929_),
    .B1(_1926_),
    .B2(_1928_),
    .A2(_1925_),
    .A1(_1922_));
 sg13g2_a22oi_1 _5638_ (.Y(_1930_),
    .B1(_1542_),
    .B2(_1876_),
    .A2(_1390_),
    .A1(_1379_));
 sg13g2_mux2_1 _5639_ (.A0(_1684_),
    .A1(_1930_),
    .S(_1462_),
    .X(_1931_));
 sg13g2_mux2_1 _5640_ (.A0(_1882_),
    .A1(_1843_),
    .S(net40),
    .X(_1932_));
 sg13g2_a22oi_1 _5641_ (.Y(_1933_),
    .B1(_1932_),
    .B2(_1865_),
    .A2(_1931_),
    .A1(_1824_));
 sg13g2_nand4_1 _5642_ (.B(_1920_),
    .C(_1929_),
    .A(_1917_),
    .Y(_1934_),
    .D(_1933_));
 sg13g2_and3_1 _5643_ (.X(_1936_),
    .A(_1455_),
    .B(_1460_),
    .C(_1480_));
 sg13g2_o21ai_1 _5644_ (.B1(_1662_),
    .Y(_1937_),
    .A1(_1895_),
    .A2(_1936_));
 sg13g2_nand2_1 _5645_ (.Y(_1938_),
    .A(net68),
    .B(net38));
 sg13g2_nand3_1 _5646_ (.B(_1532_),
    .C(_1534_),
    .A(_1582_),
    .Y(_1939_));
 sg13g2_a21o_1 _5647_ (.A2(_1939_),
    .A1(_1938_),
    .B1(net39),
    .X(_1940_));
 sg13g2_nand3_1 _5648_ (.B(_1482_),
    .C(_1652_),
    .A(net39),
    .Y(_1941_));
 sg13g2_nand4_1 _5649_ (.B(_1937_),
    .C(_1940_),
    .A(_1894_),
    .Y(_1942_),
    .D(_1941_));
 sg13g2_o21ai_1 _5650_ (.B1(net36),
    .Y(_1943_),
    .A1(_1675_),
    .A2(_1662_));
 sg13g2_or3_1 _5651_ (.A(_1674_),
    .B(_1685_),
    .C(_1943_),
    .X(_1944_));
 sg13g2_o21ai_1 _5652_ (.B1(_1549_),
    .Y(_1945_),
    .A1(net25),
    .A2(_1412_));
 sg13g2_nand2_1 _5653_ (.Y(_1947_),
    .A(_1867_),
    .B(_1945_));
 sg13g2_nor2_1 _5654_ (.A(net68),
    .B(_1510_),
    .Y(_1948_));
 sg13g2_nor2_1 _5655_ (.A(net73),
    .B(_1526_),
    .Y(_1949_));
 sg13g2_o21ai_1 _5656_ (.B1(_1815_),
    .Y(_1950_),
    .A1(_1948_),
    .A2(_1949_));
 sg13g2_nand4_1 _5657_ (.B(_1944_),
    .C(_1947_),
    .A(_1942_),
    .Y(_1951_),
    .D(_1950_));
 sg13g2_nor2_1 _5658_ (.A(_1816_),
    .B(_1674_),
    .Y(_1952_));
 sg13g2_a22oi_1 _5659_ (.Y(_1953_),
    .B1(_1379_),
    .B2(_1390_),
    .A2(_1460_),
    .A1(_1455_));
 sg13g2_buf_1 _5660_ (.A(_1953_),
    .X(_1954_));
 sg13g2_a22oi_1 _5661_ (.Y(_1955_),
    .B1(_1918_),
    .B2(_1954_),
    .A2(net75),
    .A1(_1513_));
 sg13g2_nor2b_1 _5662_ (.A(_1955_),
    .B_N(_1830_),
    .Y(_1956_));
 sg13g2_a21oi_1 _5663_ (.A1(_1694_),
    .A2(_1670_),
    .Y(_1958_),
    .B1(_1722_));
 sg13g2_nor3_1 _5664_ (.A(net74),
    .B(_1771_),
    .C(_1670_),
    .Y(_1959_));
 sg13g2_or4_1 _5665_ (.A(_1952_),
    .B(_1956_),
    .C(_1958_),
    .D(_1959_),
    .X(_1960_));
 sg13g2_or3_1 _5666_ (.A(_1934_),
    .B(_1951_),
    .C(_1960_),
    .X(_1961_));
 sg13g2_nor4_1 _5667_ (.A(_1798_),
    .B(_1813_),
    .C(_1912_),
    .D(_1961_),
    .Y(_1962_));
 sg13g2_nor2_1 _5668_ (.A(_2610_),
    .B(_1556_),
    .Y(_1963_));
 sg13g2_xnor2_1 _5669_ (.Y(_1964_),
    .A(_0116_),
    .B(_1963_));
 sg13g2_a22oi_1 _5670_ (.Y(_1965_),
    .B1(_1605_),
    .B2(_2595_),
    .A2(_1964_),
    .A1(_1725_));
 sg13g2_or2_1 _5671_ (.X(_1966_),
    .B(_1965_),
    .A(_1357_));
 sg13g2_a21oi_1 _5672_ (.A1(_1725_),
    .A2(_1351_),
    .Y(_1967_),
    .B1(_1964_));
 sg13g2_a21oi_1 _5673_ (.A1(_0326_),
    .A2(_1357_),
    .Y(_1969_),
    .B1(_0876_));
 sg13g2_nor2_1 _5674_ (.A(_1818_),
    .B(_1969_),
    .Y(_1970_));
 sg13g2_nor2_1 _5675_ (.A(_1967_),
    .B(_1970_),
    .Y(_1971_));
 sg13g2_nand3b_1 _5676_ (.B(_2576_),
    .C(_2554_),
    .Y(_1972_),
    .A_N(net3));
 sg13g2_a21oi_2 _5677_ (.B1(_1972_),
    .Y(_1973_),
    .A2(_1971_),
    .A1(_1966_));
 sg13g2_nor2_1 _5678_ (.A(_1973_),
    .B(_1798_),
    .Y(_1974_));
 sg13g2_a21oi_1 _5679_ (.A1(_1796_),
    .A2(_1962_),
    .Y(_1975_),
    .B1(_1974_));
 sg13g2_nand2_1 _5680_ (.Y(_1976_),
    .A(_1700_),
    .B(_1702_));
 sg13g2_nand2_1 _5681_ (.Y(_1977_),
    .A(_1976_),
    .B(_1948_));
 sg13g2_a22oi_1 _5682_ (.Y(_1978_),
    .B1(_1694_),
    .B2(_1977_),
    .A2(net37),
    .A1(net72));
 sg13g2_nor2_1 _5683_ (.A(net122),
    .B(net35),
    .Y(_1980_));
 sg13g2_a21oi_1 _5684_ (.A1(net122),
    .A2(_1756_),
    .Y(_1981_),
    .B1(_1980_));
 sg13g2_nor2_1 _5685_ (.A(net72),
    .B(net55),
    .Y(_1982_));
 sg13g2_nand2_1 _5686_ (.Y(_1983_),
    .A(_1976_),
    .B(_1982_));
 sg13g2_nor2_1 _5687_ (.A(net26),
    .B(_1780_),
    .Y(_1984_));
 sg13g2_o21ai_1 _5688_ (.B1(_1976_),
    .Y(_1985_),
    .A1(_1949_),
    .A2(_1984_));
 sg13g2_o21ai_1 _5689_ (.B1(_1985_),
    .Y(_1986_),
    .A1(_1981_),
    .A2(_1983_));
 sg13g2_o21ai_1 _5690_ (.B1(_1954_),
    .Y(_1987_),
    .A1(_1978_),
    .A2(_1986_));
 sg13g2_nor2_1 _5691_ (.A(net38),
    .B(_1842_),
    .Y(_1988_));
 sg13g2_a21oi_1 _5692_ (.A1(net55),
    .A2(_1867_),
    .Y(_1989_),
    .B1(_1988_));
 sg13g2_nand2b_1 _5693_ (.Y(_1991_),
    .B(net71),
    .A_N(_1989_));
 sg13g2_nor2_1 _5694_ (.A(_1791_),
    .B(net38),
    .Y(_1992_));
 sg13g2_nor2_1 _5695_ (.A(net22),
    .B(_1683_),
    .Y(_1993_));
 sg13g2_a221oi_1 _5696_ (.B2(_1992_),
    .C1(_1993_),
    .B1(net91),
    .A1(_1954_),
    .Y(_1994_),
    .A2(_1918_));
 sg13g2_nor2b_1 _5697_ (.A(_1994_),
    .B_N(_1830_),
    .Y(_1995_));
 sg13g2_buf_1 _5698_ (.A(net22),
    .X(_1996_));
 sg13g2_nand3_1 _5699_ (.B(net89),
    .C(_1730_),
    .A(net19),
    .Y(_1997_));
 sg13g2_nor3_1 _5700_ (.A(net55),
    .B(_1729_),
    .C(_1997_),
    .Y(_1998_));
 sg13g2_a21oi_1 _5701_ (.A1(net55),
    .A2(net73),
    .Y(_1999_),
    .B1(net75));
 sg13g2_nand2_1 _5702_ (.Y(_2000_),
    .A(net21),
    .B(_1999_));
 sg13g2_a21oi_1 _5703_ (.A1(_1816_),
    .A2(_2000_),
    .Y(_2002_),
    .B1(_1674_));
 sg13g2_or2_1 _5704_ (.X(_2003_),
    .B(_1927_),
    .A(net22));
 sg13g2_a221oi_1 _5705_ (.B2(_1360_),
    .C1(net38),
    .B1(_1354_),
    .A1(net103),
    .Y(_2004_),
    .A2(net72));
 sg13g2_a21oi_1 _5706_ (.A1(_1785_),
    .A2(_2003_),
    .Y(_2005_),
    .B1(_2004_));
 sg13g2_nor3_1 _5707_ (.A(net26),
    .B(_1504_),
    .C(_2005_),
    .Y(_2006_));
 sg13g2_nor4_1 _5708_ (.A(_1995_),
    .B(_1998_),
    .C(_2002_),
    .D(_2006_),
    .Y(_2007_));
 sg13g2_or2_1 _5709_ (.X(_2008_),
    .B(_1684_),
    .A(net22));
 sg13g2_nand3_1 _5710_ (.B(_1824_),
    .C(_2008_),
    .A(_1516_),
    .Y(_2009_));
 sg13g2_nand3_1 _5711_ (.B(_1992_),
    .C(_1865_),
    .A(net89),
    .Y(_2010_));
 sg13g2_o21ai_1 _5712_ (.B1(net21),
    .Y(_2011_),
    .A1(net36),
    .A2(_1679_));
 sg13g2_nand4_1 _5713_ (.B(_1785_),
    .C(net75),
    .A(_1949_),
    .Y(_2013_),
    .D(_2011_));
 sg13g2_nand3_1 _5714_ (.B(_2010_),
    .C(_2013_),
    .A(_2009_),
    .Y(_2014_));
 sg13g2_nor2b_1 _5715_ (.A(net35),
    .B_N(net55),
    .Y(_2015_));
 sg13g2_nor3_1 _5716_ (.A(net19),
    .B(net74),
    .C(_1526_),
    .Y(_2016_));
 sg13g2_nor2_1 _5717_ (.A(_1818_),
    .B(net37),
    .Y(_2017_));
 sg13g2_o21ai_1 _5718_ (.B1(_2017_),
    .Y(_2018_),
    .A1(_2015_),
    .A2(_2016_));
 sg13g2_or2_1 _5719_ (.X(_2019_),
    .B(net56),
    .A(net70));
 sg13g2_and4_1 _5720_ (.A(net27),
    .B(_1504_),
    .C(_1482_),
    .D(_2019_),
    .X(_2020_));
 sg13g2_and2_1 _5721_ (.A(_1677_),
    .B(_1876_),
    .X(_2021_));
 sg13g2_o21ai_1 _5722_ (.B1(net19),
    .Y(_2022_),
    .A1(net36),
    .A2(_2021_));
 sg13g2_nand3b_1 _5723_ (.B(_1894_),
    .C(_2022_),
    .Y(_2024_),
    .A_N(_2020_));
 sg13g2_nor2_1 _5724_ (.A(net74),
    .B(_1670_),
    .Y(_2025_));
 sg13g2_nand2b_1 _5725_ (.Y(_2026_),
    .B(_1771_),
    .A_N(_1954_));
 sg13g2_nor2_1 _5726_ (.A(_1670_),
    .B(_1722_),
    .Y(_2027_));
 sg13g2_a21oi_1 _5727_ (.A1(_2025_),
    .A2(_2026_),
    .Y(_2028_),
    .B1(_2027_));
 sg13g2_nand3_1 _5728_ (.B(_2024_),
    .C(_2028_),
    .A(_2018_),
    .Y(_2029_));
 sg13g2_nor4_1 _5729_ (.A(net73),
    .B(_1729_),
    .C(_1730_),
    .D(_1722_),
    .Y(_2030_));
 sg13g2_nor4_1 _5730_ (.A(_2014_),
    .B(_2029_),
    .C(_1934_),
    .D(_2030_),
    .Y(_2031_));
 sg13g2_nand4_1 _5731_ (.B(_1991_),
    .C(_2007_),
    .A(_1987_),
    .Y(_2032_),
    .D(_2031_));
 sg13g2_nand2_1 _5732_ (.Y(_2033_),
    .A(_1973_),
    .B(_2032_));
 sg13g2_o21ai_1 _5733_ (.B1(_2033_),
    .Y(_2035_),
    .A1(_1320_),
    .A2(_1975_));
 sg13g2_nor2_1 _5734_ (.A(_0984_),
    .B(_0996_),
    .Y(_2036_));
 sg13g2_o21ai_1 _5735_ (.B1(_1176_),
    .Y(_2037_),
    .A1(net41),
    .A2(net58));
 sg13g2_a22oi_1 _5736_ (.Y(_2038_),
    .B1(_2037_),
    .B2(_1181_),
    .A2(net58),
    .A1(net45));
 sg13g2_nand2b_1 _5737_ (.Y(_2039_),
    .B(_1138_),
    .A_N(_2038_));
 sg13g2_nor2_2 _5738_ (.A(net30),
    .B(_1227_),
    .Y(_2040_));
 sg13g2_nor2_1 _5739_ (.A(net41),
    .B(net60),
    .Y(_2041_));
 sg13g2_and2_1 _5740_ (.A(_2040_),
    .B(_2041_),
    .X(_2042_));
 sg13g2_nor3_2 _5741_ (.A(_1021_),
    .B(_1024_),
    .C(_1067_),
    .Y(_2043_));
 sg13g2_o21ai_1 _5742_ (.B1(net30),
    .Y(_2044_),
    .A1(net79),
    .A2(_2043_));
 sg13g2_a21oi_1 _5743_ (.A1(_1278_),
    .A2(_2044_),
    .Y(_2046_),
    .B1(net51));
 sg13g2_o21ai_1 _5744_ (.B1(_1004_),
    .Y(_2047_),
    .A1(_2042_),
    .A2(_2046_));
 sg13g2_a22oi_1 _5745_ (.Y(_2048_),
    .B1(_0988_),
    .B2(_0992_),
    .A2(_0967_),
    .A1(net80));
 sg13g2_nor2_1 _5746_ (.A(net49),
    .B(net59),
    .Y(_2049_));
 sg13g2_o21ai_1 _5747_ (.B1(net47),
    .Y(_2050_),
    .A1(_2040_),
    .A2(_2049_));
 sg13g2_nand3_1 _5748_ (.B(_1045_),
    .C(_1078_),
    .A(_1041_),
    .Y(_2051_));
 sg13g2_nor2_1 _5749_ (.A(net79),
    .B(_2051_),
    .Y(_2052_));
 sg13g2_or3_1 _5750_ (.A(_1136_),
    .B(_1163_),
    .C(_2052_),
    .X(_2053_));
 sg13g2_nand4_1 _5751_ (.B(_2048_),
    .C(_2050_),
    .A(_1109_),
    .Y(_2054_),
    .D(_2053_));
 sg13g2_mux2_1 _5752_ (.A0(_1116_),
    .A1(net79),
    .S(net63),
    .X(_2055_));
 sg13g2_buf_1 _5753_ (.A(net30),
    .X(_2057_));
 sg13g2_a221oi_1 _5754_ (.B2(net20),
    .C1(net47),
    .B1(_2055_),
    .A1(net50),
    .Y(_2058_),
    .A2(_2040_));
 sg13g2_o21ai_1 _5755_ (.B1(net44),
    .Y(_2059_),
    .A1(_1207_),
    .A2(_1174_));
 sg13g2_nand3b_1 _5756_ (.B(_1237_),
    .C(_2059_),
    .Y(_2060_),
    .A_N(_2058_));
 sg13g2_nand4_1 _5757_ (.B(_2047_),
    .C(_2054_),
    .A(_2039_),
    .Y(_2061_),
    .D(_2060_));
 sg13g2_nor2_2 _5758_ (.A(_2057_),
    .B(_1094_),
    .Y(_2062_));
 sg13g2_nand2_1 _5759_ (.Y(_2063_),
    .A(net64),
    .B(_1054_));
 sg13g2_o21ai_1 _5760_ (.B1(_2063_),
    .Y(_2064_),
    .A1(net61),
    .A2(net51));
 sg13g2_a22oi_1 _5761_ (.Y(_2065_),
    .B1(_2064_),
    .B2(net45),
    .A2(_2062_),
    .A1(net58));
 sg13g2_xnor2_1 _5762_ (.Y(_2066_),
    .A(_0963_),
    .B(net29));
 sg13g2_nor3_1 _5763_ (.A(_0935_),
    .B(_0980_),
    .C(net33),
    .Y(_2068_));
 sg13g2_nand3_1 _5764_ (.B(_2066_),
    .C(_2068_),
    .A(net61),
    .Y(_2069_));
 sg13g2_o21ai_1 _5765_ (.B1(_2069_),
    .Y(_2070_),
    .A1(_1152_),
    .A2(_2065_));
 sg13g2_and3_1 _5766_ (.X(_2071_),
    .A(_1196_),
    .B(_1253_),
    .C(_2062_));
 sg13g2_nand2_1 _5767_ (.Y(_2072_),
    .A(net59),
    .B(net46));
 sg13g2_o21ai_1 _5768_ (.B1(_2072_),
    .Y(_2073_),
    .A1(net42),
    .A2(net51));
 sg13g2_xnor2_1 _5769_ (.Y(_2074_),
    .A(net78),
    .B(net46));
 sg13g2_a22oi_1 _5770_ (.Y(_2075_),
    .B1(_2074_),
    .B2(_1091_),
    .A2(_2073_),
    .A1(net45));
 sg13g2_nand4_1 _5771_ (.B(net34),
    .C(net64),
    .A(net41),
    .Y(_2076_),
    .D(net57));
 sg13g2_a221oi_1 _5772_ (.B2(_2076_),
    .C1(_1000_),
    .B1(_2075_),
    .A1(_1210_),
    .Y(_2077_),
    .A2(_1213_));
 sg13g2_nor4_1 _5773_ (.A(_2061_),
    .B(_2070_),
    .C(_2071_),
    .D(_2077_),
    .Y(_2079_));
 sg13g2_o21ai_1 _5774_ (.B1(net63),
    .Y(_2080_),
    .A1(net30),
    .A2(net78));
 sg13g2_o21ai_1 _5775_ (.B1(net51),
    .Y(_2081_),
    .A1(_2049_),
    .A2(_2080_));
 sg13g2_nand3b_1 _5776_ (.B(net43),
    .C(_2057_),
    .Y(_2082_),
    .A_N(_2043_));
 sg13g2_nand3_1 _5777_ (.B(_1225_),
    .C(_2082_),
    .A(net47),
    .Y(_2083_));
 sg13g2_nand3_1 _5778_ (.B(_2081_),
    .C(_2083_),
    .A(_1153_),
    .Y(_2084_));
 sg13g2_o21ai_1 _5779_ (.B1(_2084_),
    .Y(_2085_),
    .A1(net62),
    .A2(_1247_));
 sg13g2_nand3_1 _5780_ (.B(_0898_),
    .C(net62),
    .A(net129),
    .Y(_2086_));
 sg13g2_nand3_1 _5781_ (.B(_1240_),
    .C(net43),
    .A(net94),
    .Y(_2087_));
 sg13g2_nand2_1 _5782_ (.Y(_2088_),
    .A(net92),
    .B(net23));
 sg13g2_a21oi_1 _5783_ (.A1(_2086_),
    .A2(_2087_),
    .Y(_2090_),
    .B1(_2088_));
 sg13g2_nor2_1 _5784_ (.A(net46),
    .B(net43),
    .Y(_2091_));
 sg13g2_xnor2_1 _5785_ (.Y(_2092_),
    .A(net48),
    .B(net61));
 sg13g2_a22oi_1 _5786_ (.Y(_2093_),
    .B1(_2092_),
    .B2(_1169_),
    .A2(_2091_),
    .A1(_1091_));
 sg13g2_nor2b_1 _5787_ (.A(_2093_),
    .B_N(_1187_),
    .Y(_2094_));
 sg13g2_a21o_1 _5788_ (.A2(_2090_),
    .A1(_1242_),
    .B1(_2094_),
    .X(_2095_));
 sg13g2_mux2_1 _5789_ (.A0(net62),
    .A1(_1174_),
    .S(net41),
    .X(_2096_));
 sg13g2_a21o_1 _5790_ (.A2(_1176_),
    .A1(net34),
    .B1(net44),
    .X(_2097_));
 sg13g2_a21oi_1 _5791_ (.A1(net20),
    .A2(_2096_),
    .Y(_2098_),
    .B1(_2097_));
 sg13g2_nor2_1 _5792_ (.A(net42),
    .B(_1092_),
    .Y(_2099_));
 sg13g2_o21ai_1 _5793_ (.B1(_1160_),
    .Y(_2101_),
    .A1(_2098_),
    .A2(_2099_));
 sg13g2_nor3_1 _5794_ (.A(net20),
    .B(net42),
    .C(net33),
    .Y(_2102_));
 sg13g2_nor2_1 _5795_ (.A(net34),
    .B(net57),
    .Y(_2103_));
 sg13g2_nand2_1 _5796_ (.Y(_2104_),
    .A(net62),
    .B(net46));
 sg13g2_mux2_1 _5797_ (.A0(_1078_),
    .A1(_1054_),
    .S(net64),
    .X(_2105_));
 sg13g2_a221oi_1 _5798_ (.B2(net29),
    .C1(net50),
    .B1(_2105_),
    .A1(_2103_),
    .Y(_2106_),
    .A2(_2104_));
 sg13g2_o21ai_1 _5799_ (.B1(_1208_),
    .Y(_2107_),
    .A1(_2102_),
    .A2(_2106_));
 sg13g2_nand3b_1 _5800_ (.B(_2101_),
    .C(_2107_),
    .Y(_2108_),
    .A_N(_1205_));
 sg13g2_nand3_1 _5801_ (.B(net59),
    .C(net44),
    .A(net48),
    .Y(_2109_));
 sg13g2_o21ai_1 _5802_ (.B1(_2109_),
    .Y(_2110_),
    .A1(net48),
    .A2(_2063_));
 sg13g2_a221oi_1 _5803_ (.B2(_1182_),
    .C1(_0935_),
    .B1(_2110_),
    .A1(net58),
    .Y(_2112_),
    .A2(net23));
 sg13g2_nor2_2 _5804_ (.A(_1100_),
    .B(net79),
    .Y(_2113_));
 sg13g2_nand4_1 _5805_ (.B(net34),
    .C(net60),
    .A(net41),
    .Y(_2114_),
    .D(_2113_));
 sg13g2_nand2_1 _5806_ (.Y(_2115_),
    .A(_0935_),
    .B(_2114_));
 sg13g2_nand2_1 _5807_ (.Y(_2116_),
    .A(_0993_),
    .B(_2115_));
 sg13g2_nand2_1 _5808_ (.Y(_2117_),
    .A(_1182_),
    .B(_1069_));
 sg13g2_nand4_1 _5809_ (.B(_1273_),
    .C(_1251_),
    .A(_2117_),
    .Y(_2118_),
    .D(_2051_));
 sg13g2_o21ai_1 _5810_ (.B1(_2118_),
    .Y(_2119_),
    .A1(_2112_),
    .A2(_2116_));
 sg13g2_nor4_2 _5811_ (.A(_2085_),
    .B(_2095_),
    .C(_2108_),
    .Y(_2120_),
    .D(_2119_));
 sg13g2_nand3_1 _5812_ (.B(net44),
    .C(_1091_),
    .A(net61),
    .Y(_2121_));
 sg13g2_o21ai_1 _5813_ (.B1(net45),
    .Y(_2123_),
    .A1(_1216_),
    .A2(net46));
 sg13g2_nand3_1 _5814_ (.B(_2076_),
    .C(_2123_),
    .A(_2121_),
    .Y(_2124_));
 sg13g2_nand2b_1 _5815_ (.Y(_2125_),
    .B(net29),
    .A_N(_1176_));
 sg13g2_nor2_1 _5816_ (.A(net29),
    .B(net42),
    .Y(_2126_));
 sg13g2_a21oi_1 _5817_ (.A1(_2080_),
    .A2(_2125_),
    .Y(_2127_),
    .B1(_2126_));
 sg13g2_a22oi_1 _5818_ (.Y(_2128_),
    .B1(_2127_),
    .B2(_1138_),
    .A2(_2124_),
    .A1(_1214_));
 sg13g2_and2_1 _5819_ (.A(net61),
    .B(_1198_),
    .X(_2129_));
 sg13g2_nand2_1 _5820_ (.Y(_2130_),
    .A(_1253_),
    .B(_2129_));
 sg13g2_nor3_1 _5821_ (.A(_1281_),
    .B(_1056_),
    .C(_1094_),
    .Y(_2131_));
 sg13g2_nand2_1 _5822_ (.Y(_2132_),
    .A(_0981_),
    .B(_2131_));
 sg13g2_nor2_1 _5823_ (.A(net33),
    .B(_2103_),
    .Y(_2134_));
 sg13g2_nor2_1 _5824_ (.A(_1053_),
    .B(_1092_),
    .Y(_2135_));
 sg13g2_o21ai_1 _5825_ (.B1(_1160_),
    .Y(_2136_),
    .A1(_2134_),
    .A2(_2135_));
 sg13g2_nand4_1 _5826_ (.B(_2130_),
    .C(_2132_),
    .A(_2128_),
    .Y(_2137_),
    .D(_2136_));
 sg13g2_nand3_1 _5827_ (.B(net44),
    .C(net57),
    .A(net48),
    .Y(_2138_));
 sg13g2_nand3_1 _5828_ (.B(_1080_),
    .C(_1119_),
    .A(_1130_),
    .Y(_2139_));
 sg13g2_nand4_1 _5829_ (.B(net34),
    .C(_1216_),
    .A(_1224_),
    .Y(_2140_),
    .D(net46));
 sg13g2_nand4_1 _5830_ (.B(_2138_),
    .C(_2139_),
    .A(_1092_),
    .Y(_2141_),
    .D(_2140_));
 sg13g2_nor3_1 _5831_ (.A(_1021_),
    .B(_1027_),
    .C(net79),
    .Y(_2142_));
 sg13g2_a22oi_1 _5832_ (.Y(_2143_),
    .B1(_2142_),
    .B2(_2051_),
    .A2(_1196_),
    .A1(_1131_));
 sg13g2_nand3_1 _5833_ (.B(net47),
    .C(_1091_),
    .A(net42),
    .Y(_2145_));
 sg13g2_o21ai_1 _5834_ (.B1(_2145_),
    .Y(_2146_),
    .A1(net47),
    .A2(_2143_));
 sg13g2_a22oi_1 _5835_ (.Y(_2147_),
    .B1(_2146_),
    .B2(_1187_),
    .A2(_2141_),
    .A1(_1208_));
 sg13g2_nor2_1 _5836_ (.A(_1069_),
    .B(_1014_),
    .Y(_2148_));
 sg13g2_o21ai_1 _5837_ (.B1(_1157_),
    .Y(_2149_),
    .A1(_1135_),
    .A2(net57));
 sg13g2_nor2_1 _5838_ (.A(net166),
    .B(_0855_),
    .Y(_2150_));
 sg13g2_nor2_1 _5839_ (.A(_2669_),
    .B(_0855_),
    .Y(_2151_));
 sg13g2_o21ai_1 _5840_ (.B1(_1050_),
    .Y(_2152_),
    .A1(_2150_),
    .A2(_2151_));
 sg13g2_o21ai_1 _5841_ (.B1(_0850_),
    .Y(_2153_),
    .A1(_1050_),
    .A2(_1039_));
 sg13g2_a21oi_1 _5842_ (.A1(_2152_),
    .A2(_2153_),
    .Y(_2154_),
    .B1(_0857_));
 sg13g2_o21ai_1 _5843_ (.B1(net114),
    .Y(_2156_),
    .A1(net187),
    .A2(net128));
 sg13g2_o21ai_1 _5844_ (.B1(_2156_),
    .Y(_2157_),
    .A1(_2914_),
    .A2(_1072_));
 sg13g2_nand2_1 _5845_ (.Y(_2158_),
    .A(_0855_),
    .B(_1022_));
 sg13g2_o21ai_1 _5846_ (.B1(_2158_),
    .Y(_2159_),
    .A1(_1060_),
    .A2(_0855_));
 sg13g2_nand2b_1 _5847_ (.Y(_2160_),
    .B(_2159_),
    .A_N(_0852_));
 sg13g2_o21ai_1 _5848_ (.B1(_2160_),
    .Y(_2161_),
    .A1(_1065_),
    .A2(_2157_));
 sg13g2_nor4_1 _5849_ (.A(net48),
    .B(_1119_),
    .C(_2154_),
    .D(_2161_),
    .Y(_2162_));
 sg13g2_a221oi_1 _5850_ (.B2(_2041_),
    .C1(_2162_),
    .B1(_2149_),
    .A1(_1131_),
    .Y(_2163_),
    .A2(_2148_));
 sg13g2_nand2b_1 _5851_ (.Y(_2164_),
    .B(_1153_),
    .A_N(_2163_));
 sg13g2_nor3_1 _5852_ (.A(net34),
    .B(_1163_),
    .C(_2113_),
    .Y(_2165_));
 sg13g2_o21ai_1 _5853_ (.B1(net48),
    .Y(_2167_),
    .A1(_1135_),
    .A2(net64));
 sg13g2_o21ai_1 _5854_ (.B1(_2114_),
    .Y(_2168_),
    .A1(_2165_),
    .A2(_2167_));
 sg13g2_nand3_1 _5855_ (.B(_0993_),
    .C(_2168_),
    .A(_1107_),
    .Y(_2169_));
 sg13g2_a21oi_1 _5856_ (.A1(net20),
    .A2(_1174_),
    .Y(_2170_),
    .B1(_1103_));
 sg13g2_o21ai_1 _5857_ (.B1(_1070_),
    .Y(_2171_),
    .A1(_1257_),
    .A2(_2170_));
 sg13g2_nand2_1 _5858_ (.Y(_2172_),
    .A(_1004_),
    .B(_2171_));
 sg13g2_nand4_1 _5859_ (.B(_2164_),
    .C(_2169_),
    .A(_2147_),
    .Y(_2173_),
    .D(_2172_));
 sg13g2_nand2_1 _5860_ (.Y(_2174_),
    .A(_1218_),
    .B(_2062_));
 sg13g2_nand2_1 _5861_ (.Y(_2175_),
    .A(net30),
    .B(net78));
 sg13g2_nor2_1 _5862_ (.A(net47),
    .B(_2175_),
    .Y(_2176_));
 sg13g2_a21oi_1 _5863_ (.A1(_1055_),
    .A2(_1157_),
    .Y(_2178_),
    .B1(_1015_));
 sg13g2_o21ai_1 _5864_ (.B1(net48),
    .Y(_2179_),
    .A1(_2176_),
    .A2(_2178_));
 sg13g2_a21oi_1 _5865_ (.A1(_2174_),
    .A2(_2179_),
    .Y(_2180_),
    .B1(_1152_));
 sg13g2_a21oi_1 _5866_ (.A1(net94),
    .A2(net62),
    .Y(_2181_),
    .B1(_0880_));
 sg13g2_nand3_1 _5867_ (.B(_0896_),
    .C(_2181_),
    .A(_0894_),
    .Y(_2182_));
 sg13g2_o21ai_1 _5868_ (.B1(_2182_),
    .Y(_2183_),
    .A1(_0980_),
    .A2(net43));
 sg13g2_nand3_1 _5869_ (.B(_1242_),
    .C(_2183_),
    .A(net23),
    .Y(_2184_));
 sg13g2_a21o_1 _5870_ (.A2(_1216_),
    .A1(net20),
    .B1(_1103_),
    .X(_2185_));
 sg13g2_a22oi_1 _5871_ (.Y(_2186_),
    .B1(_2185_),
    .B2(_1273_),
    .A2(_1291_),
    .A1(_1272_));
 sg13g2_nand2b_1 _5872_ (.Y(_2187_),
    .B(_1237_),
    .A_N(_2186_));
 sg13g2_nor3_1 _5873_ (.A(_2040_),
    .B(_1095_),
    .C(_2126_),
    .Y(_2189_));
 sg13g2_o21ai_1 _5874_ (.B1(_1106_),
    .Y(_2190_),
    .A1(_1093_),
    .A2(_2189_));
 sg13g2_nand3_1 _5875_ (.B(_2187_),
    .C(_2190_),
    .A(_2184_),
    .Y(_2191_));
 sg13g2_nor4_2 _5876_ (.A(_2137_),
    .B(_2173_),
    .C(_2180_),
    .Y(_2192_),
    .D(_2191_));
 sg13g2_o21ai_1 _5877_ (.B1(_1070_),
    .Y(_2193_),
    .A1(_1281_),
    .A2(_1257_));
 sg13g2_a22oi_1 _5878_ (.Y(_2194_),
    .B1(_2193_),
    .B2(_1004_),
    .A2(_2129_),
    .A1(_0981_));
 sg13g2_o21ai_1 _5879_ (.B1(_1237_),
    .Y(_2195_),
    .A1(_1228_),
    .A2(_2131_));
 sg13g2_a22oi_1 _5880_ (.Y(_2196_),
    .B1(_1093_),
    .B2(_1106_),
    .A2(net45),
    .A1(_1138_));
 sg13g2_nor2_1 _5881_ (.A(_2175_),
    .B(net33),
    .Y(_2197_));
 sg13g2_o21ai_1 _5882_ (.B1(_1165_),
    .Y(_2198_),
    .A1(_1114_),
    .A2(net33));
 sg13g2_a22oi_1 _5883_ (.Y(_2200_),
    .B1(_2198_),
    .B2(_1160_),
    .A2(_2197_),
    .A1(_1251_));
 sg13g2_nand4_1 _5884_ (.B(_2195_),
    .C(_2196_),
    .A(_2194_),
    .Y(_2201_),
    .D(_2200_));
 sg13g2_nor3_1 _5885_ (.A(_0936_),
    .B(net20),
    .C(net61),
    .Y(_2202_));
 sg13g2_a22oi_1 _5886_ (.Y(_2203_),
    .B1(_2202_),
    .B2(_0977_),
    .A2(_1169_),
    .A1(_1106_));
 sg13g2_and2_1 _5887_ (.A(net58),
    .B(net23),
    .X(_2204_));
 sg13g2_nand2_1 _5888_ (.Y(_2205_),
    .A(_2204_),
    .B(_1253_));
 sg13g2_o21ai_1 _5889_ (.B1(_2205_),
    .Y(_2206_),
    .A1(net32),
    .A2(_2203_));
 sg13g2_nand2_1 _5890_ (.Y(_2207_),
    .A(net29),
    .B(net78));
 sg13g2_o21ai_1 _5891_ (.B1(_2207_),
    .Y(_2208_),
    .A1(net29),
    .A2(net58));
 sg13g2_a221oi_1 _5892_ (.B2(_2041_),
    .C1(_1120_),
    .B1(_2208_),
    .A1(net45),
    .Y(_2209_),
    .A2(_2148_));
 sg13g2_a221oi_1 _5893_ (.B2(net59),
    .C1(_1272_),
    .B1(net23),
    .A1(_1181_),
    .Y(_2211_),
    .A2(_1179_));
 sg13g2_nand2b_1 _5894_ (.Y(_2212_),
    .B(_1187_),
    .A_N(_2211_));
 sg13g2_o21ai_1 _5895_ (.B1(_2212_),
    .Y(_2213_),
    .A1(_1108_),
    .A2(_2209_));
 sg13g2_nor4_2 _5896_ (.A(_1287_),
    .B(_2201_),
    .C(_2206_),
    .Y(_2214_),
    .D(_2213_));
 sg13g2_nand4_1 _5897_ (.B(_2120_),
    .C(_2192_),
    .A(_2079_),
    .Y(_2215_),
    .D(_2214_));
 sg13g2_a21oi_1 _5898_ (.A1(_2036_),
    .A2(_2215_),
    .Y(_2216_),
    .B1(_0831_));
 sg13g2_and2_1 _5899_ (.A(_0247_),
    .B(_0716_),
    .X(_2217_));
 sg13g2_buf_2 _5900_ (.A(ui_in[4]),
    .X(_2218_));
 sg13g2_nand2_1 _5901_ (.Y(_2219_),
    .A(_2218_),
    .B(_1320_));
 sg13g2_nand2_1 _5902_ (.Y(_2220_),
    .A(_2217_),
    .B(_2219_));
 sg13g2_inv_1 _5903_ (.Y(_2222_),
    .A(_2220_));
 sg13g2_a221oi_1 _5904_ (.B2(_2216_),
    .C1(_2222_),
    .B1(_2035_),
    .A1(_0999_),
    .Y(_2223_),
    .A2(_1297_));
 sg13g2_mux2_1 _5905_ (.A0(_2699_),
    .A1(_2701_),
    .S(_2223_),
    .X(net10));
 sg13g2_nand2_1 _5906_ (.Y(_2224_),
    .A(_2218_),
    .B(_1313_));
 sg13g2_o21ai_1 _5907_ (.B1(_1973_),
    .Y(_2225_),
    .A1(_1813_),
    .A2(_1912_));
 sg13g2_o21ai_1 _5908_ (.B1(_2225_),
    .Y(_2226_),
    .A1(net18),
    .A2(_1975_));
 sg13g2_nor3_1 _5909_ (.A(_0831_),
    .B(_0998_),
    .C(_2192_),
    .Y(_2227_));
 sg13g2_a221oi_1 _5910_ (.B2(_2216_),
    .C1(_2227_),
    .B1(_2226_),
    .A1(_2217_),
    .Y(_2228_),
    .A2(_2224_));
 sg13g2_mux2_1 _5911_ (.A0(_2699_),
    .A1(_2701_),
    .S(_2228_),
    .X(net11));
 sg13g2_and3_1 _5912_ (.X(_2229_),
    .A(_0108_),
    .B(_0246_),
    .C(_0829_));
 sg13g2_buf_1 _5913_ (.A(_2229_),
    .X(_2231_));
 sg13g2_or4_1 _5914_ (.A(_2061_),
    .B(_2070_),
    .C(_2071_),
    .D(_2077_),
    .X(_2232_));
 sg13g2_or4_1 _5915_ (.A(_2085_),
    .B(_2095_),
    .C(_2108_),
    .D(_2119_),
    .X(_2233_));
 sg13g2_nor2_1 _5916_ (.A(_2232_),
    .B(_2233_),
    .Y(_2234_));
 sg13g2_nand2_1 _5917_ (.Y(_2235_),
    .A(_2192_),
    .B(_2214_));
 sg13g2_nand4_1 _5918_ (.B(_2036_),
    .C(_2234_),
    .A(_2231_),
    .Y(_2236_),
    .D(_2235_));
 sg13g2_inv_1 _5919_ (.Y(_2237_),
    .A(_2218_));
 sg13g2_nand2_1 _5920_ (.Y(_2238_),
    .A(_1315_),
    .B(_1318_));
 sg13g2_xnor2_1 _5921_ (.Y(_2239_),
    .A(net18),
    .B(_2238_));
 sg13g2_or2_1 _5922_ (.X(_2240_),
    .B(_2239_),
    .A(_2237_));
 sg13g2_and2_1 _5923_ (.A(_0716_),
    .B(_2240_),
    .X(_2242_));
 sg13g2_buf_1 _5924_ (.A(_2242_),
    .X(_2243_));
 sg13g2_or2_1 _5925_ (.X(_2244_),
    .B(_2243_),
    .A(_2231_));
 sg13g2_inv_1 _5926_ (.Y(_2245_),
    .A(_2701_));
 sg13g2_a21oi_1 _5927_ (.A1(_2236_),
    .A2(_2244_),
    .Y(_2246_),
    .B1(_2245_));
 sg13g2_a21o_1 _5928_ (.A2(_1971_),
    .A1(_1966_),
    .B1(_1972_),
    .X(_2247_));
 sg13g2_a21oi_1 _5929_ (.A1(_1734_),
    .A2(_1795_),
    .Y(_2248_),
    .B1(_2247_));
 sg13g2_a21oi_1 _5930_ (.A1(_2036_),
    .A2(_2215_),
    .Y(_2249_),
    .B1(_2248_));
 sg13g2_a21o_1 _5931_ (.A2(_1962_),
    .A1(_1796_),
    .B1(_1974_),
    .X(_2250_));
 sg13g2_a22oi_1 _5932_ (.Y(_2251_),
    .B1(_2243_),
    .B2(_0831_),
    .A2(_2239_),
    .A1(_2250_));
 sg13g2_and3_1 _5933_ (.X(_2253_),
    .A(_2701_),
    .B(_2249_),
    .C(_2251_));
 sg13g2_and2_1 _5934_ (.A(_2234_),
    .B(_2235_),
    .X(_2254_));
 sg13g2_o21ai_1 _5935_ (.B1(_2699_),
    .Y(_2255_),
    .A1(_2231_),
    .A2(_2243_));
 sg13g2_a221oi_1 _5936_ (.B2(_0999_),
    .C1(_2255_),
    .B1(_2254_),
    .A1(_2249_),
    .Y(_2256_),
    .A2(_2251_));
 sg13g2_or3_1 _5937_ (.A(_2246_),
    .B(_2253_),
    .C(_2256_),
    .X(net12));
 sg13g2_xor2_1 _5938_ (.B(_1302_),
    .A(net242),
    .X(_2257_));
 sg13g2_or2_1 _5939_ (.X(_2258_),
    .B(_2257_),
    .A(_1315_));
 sg13g2_nor3_1 _5940_ (.A(net18),
    .B(_1317_),
    .C(_2258_),
    .Y(_2259_));
 sg13g2_a21o_1 _5941_ (.A2(_2258_),
    .A1(net18),
    .B1(_2259_),
    .X(_2260_));
 sg13g2_nand2_1 _5942_ (.Y(_2261_),
    .A(_2218_),
    .B(_2260_));
 sg13g2_o21ai_1 _5943_ (.B1(_2261_),
    .Y(_2263_),
    .A1(_2218_),
    .A2(_0027_));
 sg13g2_and2_1 _5944_ (.A(_1973_),
    .B(_1961_),
    .X(_2264_));
 sg13g2_a21o_1 _5945_ (.A2(_2260_),
    .A1(_2250_),
    .B1(_2264_),
    .X(_2265_));
 sg13g2_nor3_1 _5946_ (.A(_0831_),
    .B(_0998_),
    .C(_2214_),
    .Y(_2266_));
 sg13g2_a221oi_1 _5947_ (.B2(_2216_),
    .C1(_2266_),
    .B1(_2265_),
    .A1(_0831_),
    .Y(_2267_),
    .A2(_2263_));
 sg13g2_mux2_1 _5948_ (.A0(_2699_),
    .A1(_2701_),
    .S(_2267_),
    .X(net14));
 sg13g2_nand3_1 _5949_ (.B(net50),
    .C(_2113_),
    .A(_0935_),
    .Y(_2268_));
 sg13g2_xnor2_1 _5950_ (.Y(_2269_),
    .A(net80),
    .B(_0967_));
 sg13g2_nand3_1 _5951_ (.B(_1110_),
    .C(net59),
    .A(_2269_),
    .Y(_2270_));
 sg13g2_a221oi_1 _5952_ (.B2(_2270_),
    .C1(net51),
    .B1(_2268_),
    .A1(_1041_),
    .Y(_2271_),
    .A2(_1045_));
 sg13g2_a21oi_1 _5953_ (.A1(_1164_),
    .A2(_1157_),
    .Y(_2273_),
    .B1(_1095_));
 sg13g2_nand2_1 _5954_ (.Y(_2274_),
    .A(net61),
    .B(_1164_));
 sg13g2_nor3_1 _5955_ (.A(_2269_),
    .B(_2274_),
    .C(_2167_),
    .Y(_2275_));
 sg13g2_a21o_1 _5956_ (.A2(_2273_),
    .A1(_2269_),
    .B1(_2275_),
    .X(_2276_));
 sg13g2_o21ai_1 _5957_ (.B1(_0993_),
    .Y(_2277_),
    .A1(_2271_),
    .A2(_2276_));
 sg13g2_or2_1 _5958_ (.X(_2278_),
    .B(_1243_),
    .A(_1199_));
 sg13g2_nand2_1 _5959_ (.Y(_2279_),
    .A(net24),
    .B(_2113_));
 sg13g2_o21ai_1 _5960_ (.B1(_2279_),
    .Y(_2280_),
    .A1(net24),
    .A2(_1174_));
 sg13g2_and2_1 _5961_ (.A(_1273_),
    .B(_2280_),
    .X(_2281_));
 sg13g2_o21ai_1 _5962_ (.B1(_1160_),
    .Y(_2282_),
    .A1(_2099_),
    .A2(_2281_));
 sg13g2_nor2_1 _5963_ (.A(net20),
    .B(_1176_),
    .Y(_2284_));
 sg13g2_a21oi_1 _5964_ (.A1(net43),
    .A2(_1157_),
    .Y(_2285_),
    .B1(net50));
 sg13g2_o21ai_1 _5965_ (.B1(_1138_),
    .Y(_2286_),
    .A1(_2284_),
    .A2(_2285_));
 sg13g2_nand3_1 _5966_ (.B(_2282_),
    .C(_2286_),
    .A(_2278_),
    .Y(_2287_));
 sg13g2_a21o_1 _5967_ (.A2(_2280_),
    .A1(net31),
    .B1(_2176_),
    .X(_2288_));
 sg13g2_a21oi_1 _5968_ (.A1(net32),
    .A2(_2288_),
    .Y(_2289_),
    .B1(_2102_));
 sg13g2_nor2b_1 _5969_ (.A(_2289_),
    .B_N(_1208_),
    .Y(_2290_));
 sg13g2_a22oi_1 _5970_ (.Y(_2291_),
    .B1(_2059_),
    .B2(_1237_),
    .A2(_2043_),
    .A1(_1004_));
 sg13g2_nor2_1 _5971_ (.A(net51),
    .B(_2291_),
    .Y(_2292_));
 sg13g2_nand2_1 _5972_ (.Y(_2293_),
    .A(net42),
    .B(_2049_));
 sg13g2_nand4_1 _5973_ (.B(_2043_),
    .C(_2059_),
    .A(_1237_),
    .Y(_2295_),
    .D(_2293_));
 sg13g2_nand2_1 _5974_ (.Y(_2296_),
    .A(_1004_),
    .B(_2042_));
 sg13g2_a221oi_1 _5975_ (.B2(net57),
    .C1(net24),
    .B1(net51),
    .A1(net78),
    .Y(_2297_),
    .A2(_1216_));
 sg13g2_a21oi_1 _5976_ (.A1(net78),
    .A2(net31),
    .Y(_2298_),
    .B1(net20));
 sg13g2_nor2_1 _5977_ (.A(_2297_),
    .B(_2298_),
    .Y(_2299_));
 sg13g2_a22oi_1 _5978_ (.Y(_2300_),
    .B1(_2299_),
    .B2(net32),
    .A2(_2062_),
    .A1(net57));
 sg13g2_nand2b_1 _5979_ (.Y(_2301_),
    .B(_1214_),
    .A_N(_2300_));
 sg13g2_nand3_1 _5980_ (.B(net62),
    .C(_1198_),
    .A(_0981_),
    .Y(_2302_));
 sg13g2_nand4_1 _5981_ (.B(_2296_),
    .C(_2301_),
    .A(_2295_),
    .Y(_2303_),
    .D(_2302_));
 sg13g2_nor4_1 _5982_ (.A(_2287_),
    .B(_2290_),
    .C(_2292_),
    .D(_2303_),
    .Y(_2304_));
 sg13g2_nand2_1 _5983_ (.Y(_2306_),
    .A(_2117_),
    .B(_1157_));
 sg13g2_a22oi_1 _5984_ (.Y(_2307_),
    .B1(_2306_),
    .B2(_1273_),
    .A2(_2274_),
    .A1(_1272_));
 sg13g2_nor2b_1 _5985_ (.A(_2307_),
    .B_N(_1187_),
    .Y(_2308_));
 sg13g2_nand2_1 _5986_ (.Y(_2309_),
    .A(net31),
    .B(_2040_));
 sg13g2_o21ai_1 _5987_ (.B1(_2309_),
    .Y(_2310_),
    .A1(net24),
    .A2(_2105_));
 sg13g2_a22oi_1 _5988_ (.Y(_2311_),
    .B1(_2310_),
    .B2(net32),
    .A2(_2274_),
    .A1(_2062_));
 sg13g2_nor2_1 _5989_ (.A(_1152_),
    .B(_2311_),
    .Y(_2312_));
 sg13g2_nand3_1 _5990_ (.B(_1080_),
    .C(_1115_),
    .A(net50),
    .Y(_2313_));
 sg13g2_o21ai_1 _5991_ (.B1(net43),
    .Y(_2314_),
    .A1(_1110_),
    .A2(_1103_));
 sg13g2_nand3_1 _5992_ (.B(_2313_),
    .C(_2314_),
    .A(_1207_),
    .Y(_2315_));
 sg13g2_nand2_1 _5993_ (.Y(_2317_),
    .A(_1153_),
    .B(_2081_));
 sg13g2_a21oi_1 _5994_ (.A1(net31),
    .A2(_2315_),
    .Y(_2318_),
    .B1(_2317_));
 sg13g2_a22oi_1 _5995_ (.Y(_2319_),
    .B1(_2113_),
    .B2(_1251_),
    .A2(_1253_),
    .A1(net78));
 sg13g2_nor2b_1 _5996_ (.A(_2319_),
    .B_N(net23),
    .Y(_2320_));
 sg13g2_nor4_1 _5997_ (.A(_2308_),
    .B(_2312_),
    .C(_2318_),
    .D(_2320_),
    .Y(_2321_));
 sg13g2_nand3_1 _5998_ (.B(_2304_),
    .C(_2321_),
    .A(_2277_),
    .Y(_2322_));
 sg13g2_nor2_1 _5999_ (.A(_1315_),
    .B(_1317_),
    .Y(_2323_));
 sg13g2_nor2_1 _6000_ (.A(net18),
    .B(_2323_),
    .Y(_2324_));
 sg13g2_nand3b_1 _6001_ (.B(_1302_),
    .C(_1317_),
    .Y(_2325_),
    .A_N(_1299_));
 sg13g2_o21ai_1 _6002_ (.B1(_2325_),
    .Y(_2326_),
    .A1(_1303_),
    .A2(_1317_));
 sg13g2_nand2_1 _6003_ (.Y(_2328_),
    .A(_1315_),
    .B(_2326_));
 sg13g2_xor2_1 _6004_ (.B(_1317_),
    .A(_1299_),
    .X(_2329_));
 sg13g2_and2_1 _6005_ (.A(_1315_),
    .B(_2329_),
    .X(_2330_));
 sg13g2_mux2_1 _6006_ (.A0(_2328_),
    .A1(_2330_),
    .S(net18),
    .X(_2331_));
 sg13g2_o21ai_1 _6007_ (.B1(_2331_),
    .Y(_2332_),
    .A1(_2257_),
    .A2(_2324_));
 sg13g2_nor2_1 _6008_ (.A(_1798_),
    .B(_2332_),
    .Y(_2333_));
 sg13g2_and2_1 _6009_ (.A(_1547_),
    .B(_1746_),
    .X(_2334_));
 sg13g2_nand2_1 _6010_ (.Y(_2335_),
    .A(_1867_),
    .B(_1873_));
 sg13g2_a21oi_1 _6011_ (.A1(net25),
    .A2(_2334_),
    .Y(_2336_),
    .B1(_2335_));
 sg13g2_nand2b_1 _6012_ (.Y(_2337_),
    .B(net68),
    .A_N(_1691_));
 sg13g2_nand3_1 _6013_ (.B(net72),
    .C(_1609_),
    .A(_1976_),
    .Y(_2339_));
 sg13g2_a21oi_1 _6014_ (.A1(_2337_),
    .A2(_2339_),
    .Y(_2340_),
    .B1(_1722_));
 sg13g2_nand2_1 _6015_ (.Y(_2341_),
    .A(net74),
    .B(net73));
 sg13g2_nand3_1 _6016_ (.B(net75),
    .C(_2341_),
    .A(net21),
    .Y(_2342_));
 sg13g2_o21ai_1 _6017_ (.B1(net56),
    .Y(_2343_),
    .A1(net103),
    .A2(net55));
 sg13g2_nand3_1 _6018_ (.B(net68),
    .C(_2343_),
    .A(net19),
    .Y(_2344_));
 sg13g2_a221oi_1 _6019_ (.B2(_2344_),
    .C1(net35),
    .B1(_2342_),
    .A1(_1636_),
    .Y(_2345_),
    .A2(_1639_));
 sg13g2_nor2_1 _6020_ (.A(_1774_),
    .B(_1810_),
    .Y(_2346_));
 sg13g2_a21oi_1 _6021_ (.A1(net19),
    .A2(_1845_),
    .Y(_2347_),
    .B1(_2346_));
 sg13g2_o21ai_1 _6022_ (.B1(net89),
    .Y(_2348_),
    .A1(_1993_),
    .A2(_1695_));
 sg13g2_a21oi_1 _6023_ (.A1(_2347_),
    .A2(_2348_),
    .Y(_2350_),
    .B1(_1641_));
 sg13g2_nor3_1 _6024_ (.A(net104),
    .B(net102),
    .C(_1365_),
    .Y(_2351_));
 sg13g2_a21oi_1 _6025_ (.A1(net69),
    .A2(net71),
    .Y(_2352_),
    .B1(net70));
 sg13g2_nand2_1 _6026_ (.Y(_2353_),
    .A(net69),
    .B(net70));
 sg13g2_o21ai_1 _6027_ (.B1(_2353_),
    .Y(_2354_),
    .A1(net187),
    .A2(_2352_));
 sg13g2_a22oi_1 _6028_ (.Y(_2355_),
    .B1(_2354_),
    .B2(net102),
    .A2(_2341_),
    .A1(_2351_));
 sg13g2_nor2_1 _6029_ (.A(net102),
    .B(_1469_),
    .Y(_2356_));
 sg13g2_o21ai_1 _6030_ (.B1(net73),
    .Y(_2357_),
    .A1(_2534_),
    .A2(net74));
 sg13g2_nand2_1 _6031_ (.Y(_2358_),
    .A(_1646_),
    .B(_2357_));
 sg13g2_o21ai_1 _6032_ (.B1(_2358_),
    .Y(_2359_),
    .A1(_2539_),
    .A2(_2352_));
 sg13g2_a221oi_1 _6033_ (.B2(net102),
    .C1(net81),
    .B1(_2359_),
    .A1(net70),
    .Y(_2361_),
    .A2(_2356_));
 sg13g2_a21o_1 _6034_ (.A2(_2355_),
    .A1(_0424_),
    .B1(_2361_),
    .X(_2362_));
 sg13g2_o21ai_1 _6035_ (.B1(_1571_),
    .Y(_2363_),
    .A1(_2008_),
    .A2(_1776_));
 sg13g2_a21oi_1 _6036_ (.A1(net19),
    .A2(_2362_),
    .Y(_2364_),
    .B1(_2363_));
 sg13g2_a21oi_1 _6037_ (.A1(_1791_),
    .A2(_1778_),
    .Y(_2365_),
    .B1(_1782_));
 sg13g2_nand2_1 _6038_ (.Y(_2366_),
    .A(net38),
    .B(net56));
 sg13g2_nand3_1 _6039_ (.B(net91),
    .C(_2366_),
    .A(_1996_),
    .Y(_2367_));
 sg13g2_a21oi_1 _6040_ (.A1(_2365_),
    .A2(_2367_),
    .Y(_2368_),
    .B1(_1799_));
 sg13g2_or4_1 _6041_ (.A(_2345_),
    .B(_2350_),
    .C(_2364_),
    .D(_2368_),
    .X(_2369_));
 sg13g2_nand3_1 _6042_ (.B(net72),
    .C(net36),
    .A(net21),
    .Y(_2370_));
 sg13g2_a21oi_1 _6043_ (.A1(_1816_),
    .A2(_2370_),
    .Y(_2372_),
    .B1(_1674_));
 sg13g2_nand2_1 _6044_ (.Y(_2373_),
    .A(net212),
    .B(_1400_));
 sg13g2_o21ai_1 _6045_ (.B1(_2353_),
    .Y(_2374_),
    .A1(_1380_),
    .A2(_2373_));
 sg13g2_nor2_1 _6046_ (.A(_1403_),
    .B(net148),
    .Y(_2375_));
 sg13g2_nand2b_1 _6047_ (.Y(_2376_),
    .B(_1424_),
    .A_N(net212));
 sg13g2_nand2_1 _6048_ (.Y(_2377_),
    .A(net147),
    .B(_1396_));
 sg13g2_o21ai_1 _6049_ (.B1(_2377_),
    .Y(_2378_),
    .A1(_1380_),
    .A2(_1396_));
 sg13g2_nand3_1 _6050_ (.B(_1400_),
    .C(_1403_),
    .A(net212),
    .Y(_2379_));
 sg13g2_o21ai_1 _6051_ (.B1(_2379_),
    .Y(_2380_),
    .A1(_1403_),
    .A2(_2376_));
 sg13g2_a21oi_1 _6052_ (.A1(_2376_),
    .A2(_2378_),
    .Y(_2381_),
    .B1(_2380_));
 sg13g2_a22oi_1 _6053_ (.Y(_2383_),
    .B1(_2373_),
    .B2(_2669_),
    .A2(_2376_),
    .A1(_1373_));
 sg13g2_xnor2_1 _6054_ (.Y(_2384_),
    .A(_2526_),
    .B(_1424_));
 sg13g2_xor2_1 _6055_ (.B(net211),
    .A(_2914_),
    .X(_2385_));
 sg13g2_a221oi_1 _6056_ (.B2(_2385_),
    .C1(_2670_),
    .B1(_2384_),
    .A1(_1396_),
    .Y(_2386_),
    .A2(_2383_));
 sg13g2_a21oi_1 _6057_ (.A1(_2670_),
    .A2(_2381_),
    .Y(_2387_),
    .B1(_2386_));
 sg13g2_a221oi_1 _6058_ (.B2(_2373_),
    .C1(_2387_),
    .B1(_2375_),
    .A1(net148),
    .Y(_2388_),
    .A2(_2374_));
 sg13g2_or3_1 _6059_ (.A(_1996_),
    .B(net25),
    .C(_2388_),
    .X(_2389_));
 sg13g2_o21ai_1 _6060_ (.B1(net27),
    .Y(_2390_),
    .A1(_1576_),
    .A2(_1547_));
 sg13g2_nand3_1 _6061_ (.B(_1677_),
    .C(_1746_),
    .A(_1465_),
    .Y(_2391_));
 sg13g2_nand3_1 _6062_ (.B(_2390_),
    .C(_2391_),
    .A(net25),
    .Y(_2392_));
 sg13g2_a21oi_1 _6063_ (.A1(_2389_),
    .A2(_2392_),
    .Y(_2394_),
    .B1(_1610_));
 sg13g2_nor2_1 _6064_ (.A(_2372_),
    .B(_2394_),
    .Y(_2395_));
 sg13g2_nor2_1 _6065_ (.A(net21),
    .B(net68),
    .Y(_2396_));
 sg13g2_a22oi_1 _6066_ (.Y(_2397_),
    .B1(_2343_),
    .B2(_2396_),
    .A2(net91),
    .A1(_1993_));
 sg13g2_nand2b_1 _6067_ (.Y(_2398_),
    .B(_1824_),
    .A_N(_2397_));
 sg13g2_o21ai_1 _6068_ (.B1(net19),
    .Y(_2399_),
    .A1(net25),
    .A2(_2334_));
 sg13g2_nand2b_1 _6069_ (.Y(_2400_),
    .B(net21),
    .A_N(_2366_));
 sg13g2_and3_1 _6070_ (.X(_2401_),
    .A(_1826_),
    .B(_1894_),
    .C(_2400_));
 sg13g2_a22oi_1 _6071_ (.Y(_2402_),
    .B1(_2401_),
    .B2(_1750_),
    .A2(_2399_),
    .A1(_1881_));
 sg13g2_o21ai_1 _6072_ (.B1(_1774_),
    .Y(_2403_),
    .A1(net69),
    .A2(_1780_));
 sg13g2_o21ai_1 _6073_ (.B1(_1657_),
    .Y(_2405_),
    .A1(_1336_),
    .A2(net102));
 sg13g2_a22oi_1 _6074_ (.Y(_2406_),
    .B1(_2403_),
    .B2(_2405_),
    .A2(_2351_),
    .A1(net91));
 sg13g2_o21ai_1 _6075_ (.B1(_1774_),
    .Y(_2407_),
    .A1(_2539_),
    .A2(_1780_));
 sg13g2_nand4_1 _6076_ (.B(net69),
    .C(net102),
    .A(_1336_),
    .Y(_2408_),
    .D(_2407_));
 sg13g2_nor3_1 _6077_ (.A(net69),
    .B(net72),
    .C(_1761_),
    .Y(_2409_));
 sg13g2_nor3_1 _6078_ (.A(net121),
    .B(_1469_),
    .C(_1780_),
    .Y(_2410_));
 sg13g2_o21ai_1 _6079_ (.B1(_0424_),
    .Y(_2411_),
    .A1(_2409_),
    .A2(_2410_));
 sg13g2_nand4_1 _6080_ (.B(_2406_),
    .C(_2408_),
    .A(net19),
    .Y(_2412_),
    .D(_2411_));
 sg13g2_a221oi_1 _6081_ (.B2(_1360_),
    .C1(_1511_),
    .B1(_1354_),
    .A1(net21),
    .Y(_2413_),
    .A2(_1504_));
 sg13g2_nand2_1 _6082_ (.Y(_2414_),
    .A(_1756_),
    .B(net70));
 sg13g2_o21ai_1 _6083_ (.B1(_2414_),
    .Y(_2416_),
    .A1(net26),
    .A2(_2341_));
 sg13g2_a22oi_1 _6084_ (.Y(_2417_),
    .B1(_2416_),
    .B2(_1815_),
    .A2(_2413_),
    .A1(_2412_));
 sg13g2_nand4_1 _6085_ (.B(_2398_),
    .C(_2402_),
    .A(_2395_),
    .Y(_2418_),
    .D(_2417_));
 sg13g2_or4_1 _6086_ (.A(_2336_),
    .B(_2340_),
    .C(_2369_),
    .D(_2418_),
    .X(_2419_));
 sg13g2_nand3_1 _6087_ (.B(_1920_),
    .C(_1929_),
    .A(_1917_),
    .Y(_2420_));
 sg13g2_o21ai_1 _6088_ (.B1(_1933_),
    .Y(_2421_),
    .A1(_1799_),
    .A2(_1812_));
 sg13g2_or4_1 _6089_ (.A(_2420_),
    .B(_1951_),
    .C(_1960_),
    .D(_2421_),
    .X(_2422_));
 sg13g2_nor2_1 _6090_ (.A(_1912_),
    .B(_2422_),
    .Y(_2423_));
 sg13g2_a21oi_1 _6091_ (.A1(_1796_),
    .A2(_2423_),
    .Y(_2424_),
    .B1(_2247_));
 sg13g2_mux2_1 _6092_ (.A0(_2333_),
    .A1(_2419_),
    .S(_2424_),
    .X(_2425_));
 sg13g2_mux2_1 _6093_ (.A0(_0026_),
    .A1(_2332_),
    .S(_2218_),
    .X(_2427_));
 sg13g2_nor2_1 _6094_ (.A(_2231_),
    .B(_2427_),
    .Y(_2428_));
 sg13g2_a221oi_1 _6095_ (.B2(_2216_),
    .C1(_2428_),
    .B1(_2425_),
    .A1(_0999_),
    .Y(_2429_),
    .A2(_2322_));
 sg13g2_mux2_1 _6096_ (.A0(_2699_),
    .A1(_2701_),
    .S(_2429_),
    .X(net15));
 sg13g2_and2_1 _6097_ (.A(_1315_),
    .B(_2257_),
    .X(_2430_));
 sg13g2_o21ai_1 _6098_ (.B1(_1315_),
    .Y(_2431_),
    .A1(_1317_),
    .A2(_2257_));
 sg13g2_mux2_1 _6099_ (.A0(_2430_),
    .A1(_2431_),
    .S(net18),
    .X(_2432_));
 sg13g2_nand2_1 _6100_ (.Y(_2433_),
    .A(_2218_),
    .B(_2432_));
 sg13g2_o21ai_1 _6101_ (.B1(_2433_),
    .Y(_2434_),
    .A1(_0025_),
    .A2(_2218_));
 sg13g2_and4_1 _6102_ (.A(_2079_),
    .B(_2120_),
    .C(_2192_),
    .D(_2214_),
    .X(_2435_));
 sg13g2_o21ai_1 _6103_ (.B1(_1973_),
    .Y(_2437_),
    .A1(_1912_),
    .A2(_2422_));
 sg13g2_nor2b_1 _6104_ (.A(_1798_),
    .B_N(_2432_),
    .Y(_2438_));
 sg13g2_a21oi_1 _6105_ (.A1(_2437_),
    .A2(_2438_),
    .Y(_2439_),
    .B1(_2248_));
 sg13g2_o21ai_1 _6106_ (.B1(_2439_),
    .Y(_2440_),
    .A1(_0998_),
    .A2(_2435_));
 sg13g2_nor4_1 _6107_ (.A(_0984_),
    .B(_0996_),
    .C(_2232_),
    .D(_2233_),
    .Y(_2441_));
 sg13g2_a21oi_1 _6108_ (.A1(_2235_),
    .A2(_2441_),
    .Y(_2442_),
    .B1(_0831_));
 sg13g2_a22oi_1 _6109_ (.Y(_2443_),
    .B1(_2440_),
    .B2(_2442_),
    .A2(_2434_),
    .A1(_0831_));
 sg13g2_mux2_1 _6110_ (.A0(_2699_),
    .A1(_2701_),
    .S(_2443_),
    .X(net16));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _6120__268 (.L_HI(net268));
 sg13g2_buf_1 _6113_ (.A(net254),
    .X(uio_oe[0]));
 sg13g2_buf_1 _6114_ (.A(net255),
    .X(uio_oe[1]));
 sg13g2_buf_1 _6115_ (.A(net256),
    .X(uio_oe[2]));
 sg13g2_buf_1 _6116_ (.A(net257),
    .X(uio_oe[3]));
 sg13g2_buf_1 _6117_ (.A(net258),
    .X(uio_oe[4]));
 sg13g2_buf_1 _6118_ (.A(net259),
    .X(uio_oe[5]));
 sg13g2_buf_1 _6119_ (.A(net260),
    .X(uio_oe[6]));
 sg13g2_buf_1 _6120_ (.A(net268),
    .X(uio_oe[7]));
 sg13g2_buf_1 _6121_ (.A(net261),
    .X(uio_out[0]));
 sg13g2_buf_1 _6122_ (.A(net262),
    .X(uio_out[1]));
 sg13g2_buf_1 _6123_ (.A(net263),
    .X(uio_out[2]));
 sg13g2_buf_1 _6124_ (.A(net264),
    .X(uio_out[3]));
 sg13g2_buf_1 _6125_ (.A(net265),
    .X(uio_out[4]));
 sg13g2_buf_1 _6126_ (.A(net266),
    .X(uio_out[5]));
 sg13g2_buf_1 _6127_ (.A(net267),
    .X(uio_out[6]));
 sg13g2_buf_1 _6128_ (.A(audio),
    .X(net9));
 sg13g2_buf_1 _6129_ (.A(\graphics_engine_1.v_sync ),
    .X(net13));
 sg13g2_buf_1 _6130_ (.A(h_sync),
    .X(net17));
 sg13g2_dfrbp_1 \audio_engine_1.counter[0]$_DFFE_PN0N_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net252),
    .D(_0040_),
    .Q_N(_0033_),
    .Q(\audio_engine_1.counter[0] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[10]$_DFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net250),
    .D(_0041_),
    .Q_N(_0001_),
    .Q(\audio_engine_1.counter[10] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[11]$_DFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net248),
    .D(_0042_),
    .Q_N(_3083_),
    .Q(\audio_engine_1.counter[11] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[12]$_DFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net248),
    .D(_0043_),
    .Q_N(_3082_),
    .Q(\audio_engine_1.counter[12] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[13]$_DFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net248),
    .D(_0044_),
    .Q_N(_3081_),
    .Q(\audio_engine_1.counter[13] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[14]$_DFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net248),
    .D(_0045_),
    .Q_N(_3080_),
    .Q(\audio_engine_1.counter[14] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[15]$_DFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net248),
    .D(_0046_),
    .Q_N(_3079_),
    .Q(\audio_engine_1.counter[15] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[16]$_DFFE_PN0N_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net248),
    .D(_0047_),
    .Q_N(_3078_),
    .Q(\audio_engine_1.counter[16] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[17]$_DFFE_PN0N_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net249),
    .D(_0048_),
    .Q_N(_0000_),
    .Q(\audio_engine_1.counter[17] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[1]$_DFFE_PN0N_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net252),
    .D(_0049_),
    .Q_N(_3077_),
    .Q(\audio_engine_1.counter[1] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[2]$_DFFE_PN0N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net252),
    .D(_0050_),
    .Q_N(_3076_),
    .Q(\audio_engine_1.counter[2] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[3]$_DFFE_PN0N_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net251),
    .D(_0051_),
    .Q_N(_3075_),
    .Q(\audio_engine_1.counter[3] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[4]$_DFFE_PN0N_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net251),
    .D(_0052_),
    .Q_N(_3074_),
    .Q(\audio_engine_1.counter[4] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[5]$_DFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net250),
    .D(_0053_),
    .Q_N(_3073_),
    .Q(\audio_engine_1.counter[5] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[6]$_DFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net250),
    .D(_0054_),
    .Q_N(_3072_),
    .Q(\audio_engine_1.counter[6] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[7]$_DFFE_PN0N_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net250),
    .D(_0055_),
    .Q_N(_3071_),
    .Q(\audio_engine_1.counter[7] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[8]$_DFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net248),
    .D(_0056_),
    .Q_N(_3070_),
    .Q(\audio_engine_1.counter[8] ));
 sg13g2_dfrbp_1 \audio_engine_1.counter[9]$_DFFE_PN0N_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net248),
    .D(_0057_),
    .Q_N(_3069_),
    .Q(\audio_engine_1.counter[9] ));
 sg13g2_dfrbp_1 \audio_engine_1.en_seq_clk$_DFF_PN1_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net249),
    .D(_0038_),
    .Q_N(\audio_engine_1.en_seq_clk ),
    .Q(_3085_));
 sg13g2_dfrbp_1 \audio_engine_1.freq_synth1.audio_reg$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net249),
    .D(_0058_),
    .Q_N(_0002_),
    .Q(\audio_engine_1.freq_synth1.audio_reg ));
 sg13g2_dfrbp_1 \audio_engine_1.freq_synth1.en_synth_clk$_DFF_PN1_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net250),
    .D(_0039_),
    .Q_N(\audio_engine_1.freq_synth1.en_synth_clk ),
    .Q(_3086_));
 sg13g2_dfrbp_1 \audio_engine_1.freq_synth1.hp_ctr[0]$_DFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net250),
    .D(_0059_),
    .Q_N(\audio_engine_1.freq_synth1.hp_ctr[0] ),
    .Q(_0036_));
 sg13g2_dfrbp_1 \audio_engine_1.freq_synth1.hp_ctr[1]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net250),
    .D(_0060_),
    .Q_N(_3068_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[1] ));
 sg13g2_dfrbp_1 \audio_engine_1.freq_synth1.hp_ctr[2]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net247),
    .D(_0061_),
    .Q_N(_0009_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[2] ));
 sg13g2_dfrbp_1 \audio_engine_1.freq_synth1.hp_ctr[3]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net247),
    .D(_0062_),
    .Q_N(_0010_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[3] ));
 sg13g2_dfrbp_1 \audio_engine_1.freq_synth1.hp_ctr[4]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net246),
    .D(_0063_),
    .Q_N(_0011_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[4] ));
 sg13g2_dfrbp_1 \audio_engine_1.freq_synth1.hp_ctr[5]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net246),
    .D(_0064_),
    .Q_N(_0012_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[5] ));
 sg13g2_dfrbp_1 \audio_engine_1.freq_synth1.hp_ctr[6]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net246),
    .D(_0065_),
    .Q_N(_0014_),
    .Q(\audio_engine_1.freq_synth1.hp_ctr[6] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_ctr[0]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net249),
    .D(_0066_),
    .Q_N(_0015_),
    .Q(\audio_engine_1.seq_ctr[0] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_ctr[1]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net249),
    .D(_0067_),
    .Q_N(_3067_),
    .Q(\audio_engine_1.seq_ctr[1] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_ctr[2]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net251),
    .D(_0068_),
    .Q_N(_3066_),
    .Q(\audio_engine_1.seq_ctr[2] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_ctr[3]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net252),
    .D(_0069_),
    .Q_N(_3065_),
    .Q(\audio_engine_1.seq_ctr[3] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_ctr[4]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net252),
    .D(_0070_),
    .Q_N(_0006_),
    .Q(\audio_engine_1.seq_ctr[4] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_time[0]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net251),
    .D(_0071_),
    .Q_N(_0034_),
    .Q(\audio_engine_1.seq_time[0] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_time[1]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net247),
    .D(_0072_),
    .Q_N(_3064_),
    .Q(\audio_engine_1.seq_time[1] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_time[2]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net246),
    .D(_0073_),
    .Q_N(_0007_),
    .Q(\audio_engine_1.seq_time[2] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_time[3]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net246),
    .D(_0074_),
    .Q_N(_3063_),
    .Q(\audio_engine_1.seq_time[3] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_time[4]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net246),
    .D(_0075_),
    .Q_N(_0008_),
    .Q(\audio_engine_1.seq_time[4] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_time[5]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net246),
    .D(_0076_),
    .Q_N(_3062_),
    .Q(\audio_engine_1.seq_time[5] ));
 sg13g2_dfrbp_1 \audio_engine_1.seq_time[6]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net246),
    .D(_0077_),
    .Q_N(_3061_),
    .Q(\audio_engine_1.seq_time[6] ));
 sg13g2_dfrbp_1 \graphics_engine_1.ctr[0]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net252),
    .D(_0078_),
    .Q_N(_0035_),
    .Q(\graphics_engine_1.ctr[0] ));
 sg13g2_dfrbp_1 \graphics_engine_1.ctr[1]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net251),
    .D(_0079_),
    .Q_N(_3060_),
    .Q(\graphics_engine_1.ctr[1] ));
 sg13g2_dfrbp_1 \graphics_engine_1.ctr[2]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net247),
    .D(_0080_),
    .Q_N(_3059_),
    .Q(\graphics_engine_1.ctr[2] ));
 sg13g2_dfrbp_1 \graphics_engine_1.ctr[3]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net247),
    .D(_0081_),
    .Q_N(_3058_),
    .Q(\graphics_engine_1.ctr[3] ));
 sg13g2_dfrbp_1 \graphics_engine_1.ctr[4]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net251),
    .D(_0082_),
    .Q_N(_3057_),
    .Q(\graphics_engine_1.ctr[4] ));
 sg13g2_dfrbp_1 \graphics_engine_1.ctr[5]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net251),
    .D(_0083_),
    .Q_N(_0025_),
    .Q(\graphics_engine_1.ctr[5] ));
 sg13g2_dfrbp_1 \graphics_engine_1.ctr[6]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net252),
    .D(_0084_),
    .Q_N(_0026_),
    .Q(\graphics_engine_1.ctr[6] ));
 sg13g2_dfrbp_1 \graphics_engine_1.ctr[7]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net251),
    .D(_0085_),
    .Q_N(_0027_),
    .Q(\graphics_engine_1.ctr[7] ));
 sg13g2_dfrbp_1 \graphics_engine_1.ctr[8]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net247),
    .D(_0086_),
    .Q_N(_3056_),
    .Q(\graphics_engine_1.ctr[8] ));
 sg13g2_dfrbp_1 \graphics_engine_1.en_v_sync$_DFFE_PN1N_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net253),
    .D(_0087_),
    .Q_N(\graphics_engine_1.en_v_sync ),
    .Q(_0037_));
 sg13g2_dfrbp_1 \vga_controller_1.h_sync$_DFF_P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net269),
    .D(_0004_),
    .Q_N(_3084_),
    .Q(h_sync));
 sg13g2_dfrbp_1 \vga_controller_1.v_sync$_DFF_P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net270),
    .D(_0005_),
    .Q_N(_0003_),
    .Q(\graphics_engine_1.v_sync ));
 sg13g2_dfrbp_1 \vga_controller_1.x[0]$_SDFF_PP0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net271),
    .D(_0088_),
    .Q_N(_0032_),
    .Q(\graphics_engine_1.anim_2x[0] ));
 sg13g2_dfrbp_1 \vga_controller_1.x[1]$_SDFF_PP0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net272),
    .D(_0089_),
    .Q_N(_3055_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[1] ));
 sg13g2_dfrbp_1 \vga_controller_1.x[2]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net273),
    .D(_0090_),
    .Q_N(_3054_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[2] ));
 sg13g2_dfrbp_1 \vga_controller_1.x[3]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net274),
    .D(_0091_),
    .Q_N(_0021_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_x[0] ));
 sg13g2_dfrbp_1 \vga_controller_1.x[4]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net275),
    .D(_0092_),
    .Q_N(_0019_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[4] ));
 sg13g2_dfrbp_1 \vga_controller_1.x[5]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net276),
    .D(_0093_),
    .Q_N(_0024_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[5] ));
 sg13g2_dfrbp_1 \vga_controller_1.x[6]$_SDFF_PP0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net277),
    .D(_0094_),
    .Q_N(_0020_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[6] ));
 sg13g2_dfrbp_1 \vga_controller_1.x[7]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net278),
    .D(_0095_),
    .Q_N(_0018_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[7] ));
 sg13g2_dfrbp_1 \vga_controller_1.x[8]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net279),
    .D(_0096_),
    .Q_N(_0017_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[8] ));
 sg13g2_dfrbp_1 \vga_controller_1.x[9]$_SDFF_PP0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net280),
    .D(_0097_),
    .Q_N(_0016_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.x[9] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[0]$_SDFFCE_PP0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net281),
    .D(_0098_),
    .Q_N(_0031_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[0] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[1]$_SDFFCE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net282),
    .D(_0099_),
    .Q_N(_3053_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[1] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[2]$_SDFFCE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net283),
    .D(_0100_),
    .Q_N(_3052_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[2] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[3]$_SDFFCE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net284),
    .D(_0101_),
    .Q_N(_0022_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[0] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[4]$_SDFFCE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net285),
    .D(_0102_),
    .Q_N(_0028_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.demosiine_off_y[1] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[5]$_SDFFCE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net286),
    .D(_0103_),
    .Q_N(_0023_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[5] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[6]$_SDFFCE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net287),
    .D(_0104_),
    .Q_N(_0029_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[6] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[7]$_SDFFCE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net288),
    .D(_0105_),
    .Q_N(_0030_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[7] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[8]$_SDFFCE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net289),
    .D(_0106_),
    .Q_N(_0013_),
    .Q(\graphics_engine_1.overlay_creator1.text_demosiine1.y[8] ));
 sg13g2_dfrbp_1 \vga_controller_1.y[9]$_SDFFCE_PP0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net290),
    .D(_0107_),
    .Q_N(_3051_),
    .Q(\vga_controller_1.y[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[7]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[0]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[1]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[2]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[3]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[6]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout18 (.A(_1313_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_1996_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_2057_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1791_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1465_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_1198_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1182_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1536_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_1511_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1490_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1464_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1181_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1135_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1113_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1110_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1095_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1048_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1709_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1578_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1576_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1549_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1513_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1489_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1224_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1218_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1164_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1163_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1131_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1119_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1111_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1109_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1047_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1029_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1015_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0873_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0865_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2600_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1661_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1652_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1291_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1196_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1102_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1082_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1080_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1069_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1064_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1014_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0127_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_2865_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_2563_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1777_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1736_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1662_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1589_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_1583_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1547_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1546_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1503_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1357_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1351_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1227_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1195_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0888_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0424_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0263_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0142_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_2938_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_2864_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_2824_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1582_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1539_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1492_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1467_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1428_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0969_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0931_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0887_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0869_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0739_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0272_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_2922_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_2902_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_2898_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_2823_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_1740_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_1586_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_1420_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_1413_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_1043_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_1042_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0854_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0506_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_0271_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0267_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_2995_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_2919_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_2914_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_2897_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_2737_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_2677_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_2621_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_2610_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_2606_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_1614_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_1537_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_1476_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_1407_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_1405_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_1388_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_1384_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_1050_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_0936_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0326_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_0278_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_0270_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_0195_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_0165_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_2913_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_2732_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_2721_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_2676_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_2669_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_2620_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_2609_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_2605_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_2595_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_2566_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_1277_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_1472_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_1421_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_1392_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_1370_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_0918_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_0469_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_0322_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_0154_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_0120_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_2912_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_2900_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_2783_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_2704_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_2675_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_2670_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_2668_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_2619_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_2608_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_2604_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_2565_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_2539_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_1562_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_1551_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_1222_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_1017_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_0876_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0859_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_0155_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_0116_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_2836_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_2815_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_2785_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_2775_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_2743_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_2725_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_2695_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_2618_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_2572_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_2569_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_2564_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_2555_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_2534_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_2473_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_1540_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_1441_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_1408_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_1255_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_1211_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_1123_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_3040_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_2989_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_2959_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_2810_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_2798_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_2777_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_2774_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_2742_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_2719_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_2702_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_2580_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_2571_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_2568_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_2543_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_2542_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_2533_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_2530_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_2526_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_1825_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_1792_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_1781_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_1693_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_1649_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_1430_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_1397_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_1375_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_1321_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_1244_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_1200_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_1145_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_1112_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_2758_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_2744_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_2718_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_2693_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_2575_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_2554_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_2545_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_2541_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_2536_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_2529_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_2522_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_1715_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_1682_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_1660_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_1474_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_1364_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_1299_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_1189_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_1090_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_1079_),
    .X(net245));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(net247));
 sg13g2_buf_4 fanout247 (.X(net247),
    .A(net1));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(net253));
 sg13g2_buf_2 fanout249 (.A(net250),
    .X(net249));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(net253));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(net252));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(net253));
 sg13g2_buf_1 fanout253 (.A(net1),
    .X(net253));
 sg13g2_tielo _6113__254 (.L_LO(net254));
 sg13g2_tielo _6114__255 (.L_LO(net255));
 sg13g2_tielo _6115__256 (.L_LO(net256));
 sg13g2_tielo _6116__257 (.L_LO(net257));
 sg13g2_tielo _6117__258 (.L_LO(net258));
 sg13g2_tielo _6118__259 (.L_LO(net259));
 sg13g2_tielo _6119__260 (.L_LO(net260));
 sg13g2_tielo _6121__261 (.L_LO(net261));
 sg13g2_tielo _6122__262 (.L_LO(net262));
 sg13g2_tielo _6123__263 (.L_LO(net263));
 sg13g2_tielo _6124__264 (.L_LO(net264));
 sg13g2_tielo _6125__265 (.L_LO(net265));
 sg13g2_tielo _6126__266 (.L_LO(net266));
 sg13g2_tielo _6127__267 (.L_LO(net267));
 sg13g2_tiehi \vga_controller_1.h_sync$_DFF_P__269  (.L_HI(net269));
 sg13g2_tiehi \vga_controller_1.v_sync$_DFF_P__270  (.L_HI(net270));
 sg13g2_tiehi \vga_controller_1.x[0]$_SDFF_PP0__271  (.L_HI(net271));
 sg13g2_tiehi \vga_controller_1.x[1]$_SDFF_PP0__272  (.L_HI(net272));
 sg13g2_tiehi \vga_controller_1.x[2]$_SDFF_PP0__273  (.L_HI(net273));
 sg13g2_tiehi \vga_controller_1.x[3]$_SDFF_PP0__274  (.L_HI(net274));
 sg13g2_tiehi \vga_controller_1.x[4]$_SDFF_PP0__275  (.L_HI(net275));
 sg13g2_tiehi \vga_controller_1.x[5]$_SDFF_PP0__276  (.L_HI(net276));
 sg13g2_tiehi \vga_controller_1.x[6]$_SDFF_PP0__277  (.L_HI(net277));
 sg13g2_tiehi \vga_controller_1.x[7]$_SDFF_PP0__278  (.L_HI(net278));
 sg13g2_tiehi \vga_controller_1.x[8]$_SDFF_PP0__279  (.L_HI(net279));
 sg13g2_tiehi \vga_controller_1.x[9]$_SDFF_PP0__280  (.L_HI(net280));
 sg13g2_tiehi \vga_controller_1.y[0]$_SDFFCE_PP0P__281  (.L_HI(net281));
 sg13g2_tiehi \vga_controller_1.y[1]$_SDFFCE_PP0P__282  (.L_HI(net282));
 sg13g2_tiehi \vga_controller_1.y[2]$_SDFFCE_PP0P__283  (.L_HI(net283));
 sg13g2_tiehi \vga_controller_1.y[3]$_SDFFCE_PP0P__284  (.L_HI(net284));
 sg13g2_tiehi \vga_controller_1.y[4]$_SDFFCE_PP0P__285  (.L_HI(net285));
 sg13g2_tiehi \vga_controller_1.y[5]$_SDFFCE_PP0P__286  (.L_HI(net286));
 sg13g2_tiehi \vga_controller_1.y[6]$_SDFFCE_PP0P__287  (.L_HI(net287));
 sg13g2_tiehi \vga_controller_1.y[7]$_SDFFCE_PP0P__288  (.L_HI(net288));
 sg13g2_tiehi \vga_controller_1.y[8]$_SDFFCE_PP0P__289  (.L_HI(net289));
 sg13g2_tiehi \vga_controller_1.y[9]$_SDFFCE_PP0P__290  (.L_HI(net290));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_15_0_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0004_));
 sg13g2_antennanp ANTENNA_2 (.A(_0005_));
 sg13g2_antennanp ANTENNA_3 (.A(_0995_));
 sg13g2_antennanp ANTENNA_4 (.A(_1297_));
 sg13g2_antennanp ANTENNA_5 (.A(_0004_));
 sg13g2_antennanp ANTENNA_6 (.A(_0005_));
 sg13g2_antennanp ANTENNA_7 (.A(_0995_));
 sg13g2_antennanp ANTENNA_8 (.A(_0004_));
 sg13g2_antennanp ANTENNA_9 (.A(_0005_));
 sg13g2_antennanp ANTENNA_10 (.A(_0995_));
 sg13g2_antennanp ANTENNA_11 (.A(_0004_));
 sg13g2_antennanp ANTENNA_12 (.A(_0005_));
 sg13g2_antennanp ANTENNA_13 (.A(_0995_));
 sg13g2_antennanp ANTENNA_14 (.A(_0004_));
 sg13g2_antennanp ANTENNA_15 (.A(_0005_));
 sg13g2_antennanp ANTENNA_16 (.A(_0995_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_204 ();
 sg13g2_fill_1 FILLER_0_211 ();
 sg13g2_decap_4 FILLER_0_216 ();
 sg13g2_fill_1 FILLER_0_220 ();
 sg13g2_decap_8 FILLER_0_229 ();
 sg13g2_decap_8 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_243 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_4 FILLER_0_425 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_fill_2 FILLER_1_154 ();
 sg13g2_fill_1 FILLER_1_156 ();
 sg13g2_fill_1 FILLER_1_161 ();
 sg13g2_fill_1 FILLER_1_188 ();
 sg13g2_fill_1 FILLER_1_194 ();
 sg13g2_decap_4 FILLER_1_200 ();
 sg13g2_fill_1 FILLER_1_204 ();
 sg13g2_fill_2 FILLER_1_210 ();
 sg13g2_fill_2 FILLER_1_239 ();
 sg13g2_decap_4 FILLER_1_245 ();
 sg13g2_fill_1 FILLER_1_253 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_4 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_191 ();
 sg13g2_fill_1 FILLER_2_201 ();
 sg13g2_fill_1 FILLER_2_227 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_4 FILLER_3_176 ();
 sg13g2_fill_1 FILLER_3_185 ();
 sg13g2_fill_1 FILLER_3_195 ();
 sg13g2_decap_4 FILLER_3_201 ();
 sg13g2_fill_1 FILLER_3_205 ();
 sg13g2_fill_2 FILLER_3_223 ();
 sg13g2_fill_1 FILLER_3_225 ();
 sg13g2_fill_2 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_237 ();
 sg13g2_decap_8 FILLER_3_244 ();
 sg13g2_fill_2 FILLER_3_251 ();
 sg13g2_fill_1 FILLER_3_258 ();
 sg13g2_decap_8 FILLER_3_267 ();
 sg13g2_decap_4 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_282 ();
 sg13g2_fill_1 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_299 ();
 sg13g2_decap_8 FILLER_3_306 ();
 sg13g2_decap_8 FILLER_3_313 ();
 sg13g2_decap_8 FILLER_3_320 ();
 sg13g2_decap_8 FILLER_3_327 ();
 sg13g2_decap_8 FILLER_3_334 ();
 sg13g2_fill_2 FILLER_3_341 ();
 sg13g2_fill_1 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_353 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_367 ();
 sg13g2_decap_8 FILLER_3_374 ();
 sg13g2_decap_8 FILLER_3_381 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_4 FILLER_4_215 ();
 sg13g2_fill_1 FILLER_4_219 ();
 sg13g2_fill_2 FILLER_4_224 ();
 sg13g2_fill_1 FILLER_4_226 ();
 sg13g2_decap_8 FILLER_4_258 ();
 sg13g2_decap_4 FILLER_4_265 ();
 sg13g2_fill_1 FILLER_4_269 ();
 sg13g2_decap_4 FILLER_4_286 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_4 FILLER_4_305 ();
 sg13g2_fill_1 FILLER_4_309 ();
 sg13g2_decap_8 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_330 ();
 sg13g2_fill_2 FILLER_4_341 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_fill_2 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_174 ();
 sg13g2_decap_8 FILLER_5_181 ();
 sg13g2_decap_8 FILLER_5_192 ();
 sg13g2_decap_8 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_5_206 ();
 sg13g2_decap_4 FILLER_5_213 ();
 sg13g2_fill_1 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_fill_2 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_274 ();
 sg13g2_fill_1 FILLER_5_280 ();
 sg13g2_fill_1 FILLER_5_286 ();
 sg13g2_fill_1 FILLER_5_306 ();
 sg13g2_fill_1 FILLER_5_312 ();
 sg13g2_decap_4 FILLER_5_317 ();
 sg13g2_fill_2 FILLER_5_333 ();
 sg13g2_fill_1 FILLER_5_335 ();
 sg13g2_decap_4 FILLER_5_341 ();
 sg13g2_fill_1 FILLER_5_345 ();
 sg13g2_decap_4 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_4 FILLER_5_424 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_140 ();
 sg13g2_decap_4 FILLER_6_162 ();
 sg13g2_decap_8 FILLER_6_176 ();
 sg13g2_fill_1 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_201 ();
 sg13g2_fill_2 FILLER_6_211 ();
 sg13g2_fill_2 FILLER_6_228 ();
 sg13g2_fill_1 FILLER_6_230 ();
 sg13g2_fill_2 FILLER_6_287 ();
 sg13g2_fill_1 FILLER_6_302 ();
 sg13g2_fill_1 FILLER_6_340 ();
 sg13g2_fill_1 FILLER_6_345 ();
 sg13g2_fill_2 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_4 FILLER_7_133 ();
 sg13g2_fill_1 FILLER_7_142 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_160 ();
 sg13g2_decap_4 FILLER_7_178 ();
 sg13g2_fill_1 FILLER_7_182 ();
 sg13g2_fill_2 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_189 ();
 sg13g2_fill_1 FILLER_7_195 ();
 sg13g2_fill_2 FILLER_7_208 ();
 sg13g2_fill_2 FILLER_7_237 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_decap_8 FILLER_7_250 ();
 sg13g2_fill_2 FILLER_7_257 ();
 sg13g2_fill_2 FILLER_7_264 ();
 sg13g2_fill_1 FILLER_7_266 ();
 sg13g2_fill_2 FILLER_7_272 ();
 sg13g2_fill_1 FILLER_7_274 ();
 sg13g2_fill_2 FILLER_7_289 ();
 sg13g2_fill_1 FILLER_7_295 ();
 sg13g2_decap_4 FILLER_7_305 ();
 sg13g2_fill_1 FILLER_7_324 ();
 sg13g2_fill_2 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_fill_1 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_decap_8 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_7_414 ();
 sg13g2_decap_8 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_4 FILLER_8_112 ();
 sg13g2_fill_1 FILLER_8_143 ();
 sg13g2_fill_1 FILLER_8_153 ();
 sg13g2_fill_1 FILLER_8_158 ();
 sg13g2_fill_1 FILLER_8_164 ();
 sg13g2_fill_2 FILLER_8_177 ();
 sg13g2_fill_1 FILLER_8_184 ();
 sg13g2_fill_2 FILLER_8_215 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_decap_4 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_241 ();
 sg13g2_decap_4 FILLER_8_267 ();
 sg13g2_fill_2 FILLER_8_271 ();
 sg13g2_fill_1 FILLER_8_278 ();
 sg13g2_decap_8 FILLER_8_283 ();
 sg13g2_fill_1 FILLER_8_295 ();
 sg13g2_fill_1 FILLER_8_301 ();
 sg13g2_decap_4 FILLER_8_343 ();
 sg13g2_fill_1 FILLER_8_351 ();
 sg13g2_decap_4 FILLER_8_357 ();
 sg13g2_fill_2 FILLER_8_361 ();
 sg13g2_fill_1 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_380 ();
 sg13g2_decap_8 FILLER_8_387 ();
 sg13g2_decap_8 FILLER_8_394 ();
 sg13g2_decap_8 FILLER_8_401 ();
 sg13g2_decap_8 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_8_415 ();
 sg13g2_decap_8 FILLER_8_422 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_4 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_123 ();
 sg13g2_fill_2 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_184 ();
 sg13g2_decap_8 FILLER_9_204 ();
 sg13g2_decap_4 FILLER_9_211 ();
 sg13g2_fill_1 FILLER_9_215 ();
 sg13g2_fill_2 FILLER_9_220 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_decap_4 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_fill_1 FILLER_9_281 ();
 sg13g2_fill_1 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_298 ();
 sg13g2_fill_1 FILLER_9_314 ();
 sg13g2_fill_2 FILLER_9_324 ();
 sg13g2_fill_1 FILLER_9_336 ();
 sg13g2_fill_2 FILLER_9_346 ();
 sg13g2_decap_4 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_381 ();
 sg13g2_decap_8 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_395 ();
 sg13g2_decap_8 FILLER_9_402 ();
 sg13g2_decap_8 FILLER_9_409 ();
 sg13g2_decap_8 FILLER_9_416 ();
 sg13g2_decap_8 FILLER_9_423 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_4 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_100 ();
 sg13g2_decap_4 FILLER_10_151 ();
 sg13g2_fill_1 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_184 ();
 sg13g2_fill_2 FILLER_10_191 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_decap_4 FILLER_10_203 ();
 sg13g2_fill_1 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_213 ();
 sg13g2_decap_8 FILLER_10_220 ();
 sg13g2_decap_4 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_235 ();
 sg13g2_fill_1 FILLER_10_237 ();
 sg13g2_decap_8 FILLER_10_258 ();
 sg13g2_decap_8 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_fill_2 FILLER_10_293 ();
 sg13g2_fill_1 FILLER_10_305 ();
 sg13g2_fill_1 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_fill_2 FILLER_10_334 ();
 sg13g2_fill_1 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_fill_1 FILLER_10_360 ();
 sg13g2_decap_4 FILLER_10_366 ();
 sg13g2_fill_1 FILLER_10_370 ();
 sg13g2_decap_4 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_8 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_10_412 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_decap_4 FILLER_10_426 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_91 ();
 sg13g2_fill_2 FILLER_11_106 ();
 sg13g2_fill_1 FILLER_11_108 ();
 sg13g2_fill_1 FILLER_11_113 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_fill_1 FILLER_11_140 ();
 sg13g2_decap_4 FILLER_11_146 ();
 sg13g2_decap_4 FILLER_11_159 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_4 FILLER_11_196 ();
 sg13g2_fill_2 FILLER_11_200 ();
 sg13g2_fill_1 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_213 ();
 sg13g2_decap_8 FILLER_11_220 ();
 sg13g2_decap_4 FILLER_11_258 ();
 sg13g2_fill_1 FILLER_11_266 ();
 sg13g2_fill_2 FILLER_11_272 ();
 sg13g2_fill_1 FILLER_11_274 ();
 sg13g2_fill_2 FILLER_11_279 ();
 sg13g2_fill_1 FILLER_11_281 ();
 sg13g2_fill_2 FILLER_11_295 ();
 sg13g2_fill_1 FILLER_11_301 ();
 sg13g2_fill_1 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_fill_2 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_fill_1 FILLER_12_95 ();
 sg13g2_fill_1 FILLER_12_108 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_fill_1 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_decap_8 FILLER_12_152 ();
 sg13g2_decap_8 FILLER_12_159 ();
 sg13g2_decap_8 FILLER_12_166 ();
 sg13g2_decap_8 FILLER_12_173 ();
 sg13g2_decap_8 FILLER_12_180 ();
 sg13g2_decap_8 FILLER_12_187 ();
 sg13g2_decap_8 FILLER_12_194 ();
 sg13g2_fill_1 FILLER_12_206 ();
 sg13g2_fill_2 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_255 ();
 sg13g2_decap_8 FILLER_12_288 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_fill_2 FILLER_12_312 ();
 sg13g2_decap_4 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_fill_2 FILLER_12_347 ();
 sg13g2_fill_1 FILLER_12_354 ();
 sg13g2_fill_2 FILLER_12_363 ();
 sg13g2_fill_1 FILLER_12_365 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_4 FILLER_12_377 ();
 sg13g2_fill_1 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_decap_8 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_12_414 ();
 sg13g2_decap_8 FILLER_12_421 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_4 FILLER_13_91 ();
 sg13g2_fill_2 FILLER_13_105 ();
 sg13g2_fill_2 FILLER_13_113 ();
 sg13g2_decap_4 FILLER_13_143 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_159 ();
 sg13g2_decap_4 FILLER_13_169 ();
 sg13g2_fill_1 FILLER_13_173 ();
 sg13g2_fill_2 FILLER_13_187 ();
 sg13g2_fill_1 FILLER_13_204 ();
 sg13g2_decap_4 FILLER_13_221 ();
 sg13g2_decap_4 FILLER_13_230 ();
 sg13g2_decap_4 FILLER_13_264 ();
 sg13g2_fill_2 FILLER_13_268 ();
 sg13g2_fill_2 FILLER_13_282 ();
 sg13g2_fill_1 FILLER_13_284 ();
 sg13g2_fill_2 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_fill_2 FILLER_13_296 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_fill_1 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_fill_2 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_8 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_13_412 ();
 sg13g2_decap_8 FILLER_13_419 ();
 sg13g2_decap_4 FILLER_13_426 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_fill_2 FILLER_14_91 ();
 sg13g2_fill_1 FILLER_14_93 ();
 sg13g2_fill_1 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_167 ();
 sg13g2_fill_2 FILLER_14_174 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_decap_4 FILLER_14_205 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_2 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_244 ();
 sg13g2_fill_2 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_258 ();
 sg13g2_decap_4 FILLER_14_264 ();
 sg13g2_fill_1 FILLER_14_268 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_decap_4 FILLER_14_303 ();
 sg13g2_fill_1 FILLER_14_307 ();
 sg13g2_fill_1 FILLER_14_317 ();
 sg13g2_decap_4 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_fill_1 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_363 ();
 sg13g2_fill_2 FILLER_14_370 ();
 sg13g2_fill_2 FILLER_14_383 ();
 sg13g2_fill_1 FILLER_14_385 ();
 sg13g2_fill_1 FILLER_14_392 ();
 sg13g2_fill_1 FILLER_14_401 ();
 sg13g2_decap_8 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_14_414 ();
 sg13g2_decap_8 FILLER_14_421 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_4 FILLER_15_77 ();
 sg13g2_fill_2 FILLER_15_85 ();
 sg13g2_fill_1 FILLER_15_97 ();
 sg13g2_fill_2 FILLER_15_103 ();
 sg13g2_fill_2 FILLER_15_117 ();
 sg13g2_fill_1 FILLER_15_119 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_fill_2 FILLER_15_200 ();
 sg13g2_fill_1 FILLER_15_202 ();
 sg13g2_fill_2 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_4 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_fill_2 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_311 ();
 sg13g2_decap_4 FILLER_15_318 ();
 sg13g2_fill_2 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_337 ();
 sg13g2_fill_2 FILLER_15_369 ();
 sg13g2_decap_4 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_418 ();
 sg13g2_decap_4 FILLER_15_425 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_4 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_81 ();
 sg13g2_fill_1 FILLER_16_99 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_107 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_decap_4 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_147 ();
 sg13g2_fill_1 FILLER_16_153 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_fill_2 FILLER_16_174 ();
 sg13g2_decap_4 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_192 ();
 sg13g2_decap_8 FILLER_16_204 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_fill_1 FILLER_16_222 ();
 sg13g2_fill_2 FILLER_16_228 ();
 sg13g2_fill_1 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_244 ();
 sg13g2_fill_2 FILLER_16_253 ();
 sg13g2_fill_1 FILLER_16_255 ();
 sg13g2_decap_4 FILLER_16_261 ();
 sg13g2_fill_1 FILLER_16_265 ();
 sg13g2_fill_1 FILLER_16_282 ();
 sg13g2_fill_1 FILLER_16_288 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_1 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_314 ();
 sg13g2_fill_2 FILLER_16_321 ();
 sg13g2_fill_2 FILLER_16_327 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_fill_2 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_358 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_fill_2 FILLER_16_366 ();
 sg13g2_fill_1 FILLER_16_381 ();
 sg13g2_fill_1 FILLER_16_403 ();
 sg13g2_decap_4 FILLER_16_414 ();
 sg13g2_fill_2 FILLER_16_418 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_4 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_97 ();
 sg13g2_decap_4 FILLER_17_125 ();
 sg13g2_fill_1 FILLER_17_129 ();
 sg13g2_decap_8 FILLER_17_143 ();
 sg13g2_decap_8 FILLER_17_150 ();
 sg13g2_decap_8 FILLER_17_157 ();
 sg13g2_decap_8 FILLER_17_164 ();
 sg13g2_fill_1 FILLER_17_176 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_4 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_decap_4 FILLER_17_203 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_220 ();
 sg13g2_decap_4 FILLER_17_244 ();
 sg13g2_fill_2 FILLER_17_248 ();
 sg13g2_decap_8 FILLER_17_255 ();
 sg13g2_fill_2 FILLER_17_262 ();
 sg13g2_fill_2 FILLER_17_269 ();
 sg13g2_decap_4 FILLER_17_278 ();
 sg13g2_fill_1 FILLER_17_296 ();
 sg13g2_fill_2 FILLER_17_310 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_fill_2 FILLER_17_337 ();
 sg13g2_fill_1 FILLER_17_339 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_fill_1 FILLER_17_357 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_fill_2 FILLER_17_377 ();
 sg13g2_decap_4 FILLER_17_401 ();
 sg13g2_fill_2 FILLER_17_405 ();
 sg13g2_decap_4 FILLER_17_425 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_fill_2 FILLER_18_77 ();
 sg13g2_fill_1 FILLER_18_102 ();
 sg13g2_fill_2 FILLER_18_122 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_fill_1 FILLER_18_158 ();
 sg13g2_fill_1 FILLER_18_164 ();
 sg13g2_decap_4 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_188 ();
 sg13g2_fill_2 FILLER_18_222 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_253 ();
 sg13g2_fill_2 FILLER_18_260 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_4 FILLER_18_284 ();
 sg13g2_fill_1 FILLER_18_288 ();
 sg13g2_fill_1 FILLER_18_299 ();
 sg13g2_decap_4 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_314 ();
 sg13g2_fill_2 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_334 ();
 sg13g2_decap_4 FILLER_18_344 ();
 sg13g2_decap_4 FILLER_18_356 ();
 sg13g2_fill_1 FILLER_18_360 ();
 sg13g2_decap_4 FILLER_18_366 ();
 sg13g2_decap_4 FILLER_18_374 ();
 sg13g2_fill_2 FILLER_18_387 ();
 sg13g2_decap_4 FILLER_18_393 ();
 sg13g2_decap_4 FILLER_18_407 ();
 sg13g2_fill_2 FILLER_18_411 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_4 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_2 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_88 ();
 sg13g2_fill_2 FILLER_19_99 ();
 sg13g2_fill_1 FILLER_19_101 ();
 sg13g2_decap_4 FILLER_19_121 ();
 sg13g2_fill_2 FILLER_19_125 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_149 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_179 ();
 sg13g2_fill_2 FILLER_19_184 ();
 sg13g2_fill_1 FILLER_19_186 ();
 sg13g2_fill_1 FILLER_19_192 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_4 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_fill_2 FILLER_19_238 ();
 sg13g2_decap_4 FILLER_19_257 ();
 sg13g2_fill_2 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_300 ();
 sg13g2_decap_8 FILLER_19_307 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_fill_2 FILLER_19_356 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_decap_4 FILLER_19_373 ();
 sg13g2_fill_1 FILLER_19_377 ();
 sg13g2_fill_2 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_4 FILLER_19_395 ();
 sg13g2_fill_1 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_405 ();
 sg13g2_decap_4 FILLER_19_412 ();
 sg13g2_fill_2 FILLER_19_416 ();
 sg13g2_decap_4 FILLER_19_425 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_93 ();
 sg13g2_decap_8 FILLER_20_100 ();
 sg13g2_decap_4 FILLER_20_115 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_decap_4 FILLER_20_131 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_decap_8 FILLER_20_153 ();
 sg13g2_decap_4 FILLER_20_160 ();
 sg13g2_fill_1 FILLER_20_164 ();
 sg13g2_decap_4 FILLER_20_170 ();
 sg13g2_fill_2 FILLER_20_174 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_223 ();
 sg13g2_fill_2 FILLER_20_238 ();
 sg13g2_fill_1 FILLER_20_240 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_271 ();
 sg13g2_decap_4 FILLER_20_289 ();
 sg13g2_fill_2 FILLER_20_293 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_decap_4 FILLER_20_306 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_4 FILLER_20_353 ();
 sg13g2_fill_2 FILLER_20_361 ();
 sg13g2_fill_2 FILLER_20_369 ();
 sg13g2_decap_4 FILLER_20_388 ();
 sg13g2_fill_2 FILLER_20_392 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_64 ();
 sg13g2_fill_1 FILLER_21_71 ();
 sg13g2_decap_8 FILLER_21_76 ();
 sg13g2_fill_2 FILLER_21_98 ();
 sg13g2_decap_4 FILLER_21_105 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_122 ();
 sg13g2_fill_2 FILLER_21_129 ();
 sg13g2_decap_8 FILLER_21_156 ();
 sg13g2_decap_8 FILLER_21_163 ();
 sg13g2_decap_8 FILLER_21_170 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_fill_1 FILLER_21_179 ();
 sg13g2_fill_2 FILLER_21_188 ();
 sg13g2_fill_2 FILLER_21_194 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_decap_4 FILLER_21_225 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_decap_4 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_fill_2 FILLER_21_272 ();
 sg13g2_fill_1 FILLER_21_274 ();
 sg13g2_decap_4 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_296 ();
 sg13g2_decap_8 FILLER_21_303 ();
 sg13g2_decap_4 FILLER_21_310 ();
 sg13g2_fill_2 FILLER_21_314 ();
 sg13g2_fill_2 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_341 ();
 sg13g2_fill_2 FILLER_21_351 ();
 sg13g2_fill_1 FILLER_21_361 ();
 sg13g2_fill_1 FILLER_21_366 ();
 sg13g2_fill_1 FILLER_21_372 ();
 sg13g2_fill_1 FILLER_21_381 ();
 sg13g2_fill_1 FILLER_21_387 ();
 sg13g2_fill_1 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_413 ();
 sg13g2_fill_2 FILLER_21_419 ();
 sg13g2_decap_4 FILLER_21_426 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_49 ();
 sg13g2_fill_1 FILLER_22_59 ();
 sg13g2_fill_2 FILLER_22_80 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_fill_1 FILLER_22_88 ();
 sg13g2_fill_1 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_107 ();
 sg13g2_decap_4 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_123 ();
 sg13g2_decap_8 FILLER_22_142 ();
 sg13g2_decap_8 FILLER_22_149 ();
 sg13g2_decap_8 FILLER_22_156 ();
 sg13g2_decap_4 FILLER_22_163 ();
 sg13g2_fill_2 FILLER_22_167 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_255 ();
 sg13g2_fill_1 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_289 ();
 sg13g2_decap_4 FILLER_22_296 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_decap_8 FILLER_22_307 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_324 ();
 sg13g2_fill_2 FILLER_22_330 ();
 sg13g2_fill_2 FILLER_22_339 ();
 sg13g2_fill_2 FILLER_22_349 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_fill_1 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_388 ();
 sg13g2_fill_2 FILLER_22_394 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_fill_2 FILLER_22_416 ();
 sg13g2_decap_4 FILLER_22_426 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_49 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_fill_1 FILLER_23_80 ();
 sg13g2_decap_4 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_92 ();
 sg13g2_fill_2 FILLER_23_113 ();
 sg13g2_fill_1 FILLER_23_115 ();
 sg13g2_decap_4 FILLER_23_121 ();
 sg13g2_fill_2 FILLER_23_133 ();
 sg13g2_fill_2 FILLER_23_141 ();
 sg13g2_fill_1 FILLER_23_143 ();
 sg13g2_fill_1 FILLER_23_180 ();
 sg13g2_decap_4 FILLER_23_186 ();
 sg13g2_fill_2 FILLER_23_190 ();
 sg13g2_fill_2 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_207 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_278 ();
 sg13g2_fill_2 FILLER_23_285 ();
 sg13g2_fill_1 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_292 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_315 ();
 sg13g2_fill_2 FILLER_23_320 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_327 ();
 sg13g2_decap_4 FILLER_23_341 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_decap_4 FILLER_23_352 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_fill_2 FILLER_23_375 ();
 sg13g2_fill_1 FILLER_23_382 ();
 sg13g2_fill_2 FILLER_23_387 ();
 sg13g2_fill_2 FILLER_23_393 ();
 sg13g2_fill_2 FILLER_23_408 ();
 sg13g2_fill_1 FILLER_23_410 ();
 sg13g2_decap_4 FILLER_23_415 ();
 sg13g2_decap_8 FILLER_23_423 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_49 ();
 sg13g2_fill_2 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_fill_2 FILLER_24_106 ();
 sg13g2_fill_1 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_fill_2 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_150 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_163 ();
 sg13g2_fill_2 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_fill_2 FILLER_24_184 ();
 sg13g2_fill_2 FILLER_24_195 ();
 sg13g2_fill_2 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_204 ();
 sg13g2_decap_8 FILLER_24_220 ();
 sg13g2_fill_2 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_fill_1 FILLER_24_250 ();
 sg13g2_fill_2 FILLER_24_256 ();
 sg13g2_fill_1 FILLER_24_258 ();
 sg13g2_fill_2 FILLER_24_265 ();
 sg13g2_fill_1 FILLER_24_267 ();
 sg13g2_decap_4 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_325 ();
 sg13g2_fill_1 FILLER_24_332 ();
 sg13g2_decap_4 FILLER_24_338 ();
 sg13g2_fill_2 FILLER_24_342 ();
 sg13g2_decap_4 FILLER_24_349 ();
 sg13g2_fill_1 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_24_379 ();
 sg13g2_decap_4 FILLER_24_387 ();
 sg13g2_fill_2 FILLER_24_391 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_24_414 ();
 sg13g2_decap_8 FILLER_24_421 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_4 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_93 ();
 sg13g2_decap_8 FILLER_25_100 ();
 sg13g2_decap_8 FILLER_25_115 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_decap_4 FILLER_25_138 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_decap_4 FILLER_25_222 ();
 sg13g2_fill_2 FILLER_25_226 ();
 sg13g2_decap_4 FILLER_25_233 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_decap_8 FILLER_25_248 ();
 sg13g2_fill_2 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_309 ();
 sg13g2_fill_1 FILLER_25_321 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_fill_1 FILLER_25_334 ();
 sg13g2_fill_1 FILLER_25_339 ();
 sg13g2_fill_1 FILLER_25_356 ();
 sg13g2_fill_1 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_decap_4 FILLER_25_377 ();
 sg13g2_fill_2 FILLER_25_381 ();
 sg13g2_fill_2 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_fill_2 FILLER_25_427 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_66 ();
 sg13g2_fill_1 FILLER_26_68 ();
 sg13g2_decap_4 FILLER_26_78 ();
 sg13g2_fill_2 FILLER_26_82 ();
 sg13g2_decap_4 FILLER_26_93 ();
 sg13g2_fill_1 FILLER_26_97 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_fill_1 FILLER_26_109 ();
 sg13g2_decap_8 FILLER_26_120 ();
 sg13g2_decap_8 FILLER_26_135 ();
 sg13g2_decap_8 FILLER_26_142 ();
 sg13g2_decap_8 FILLER_26_149 ();
 sg13g2_decap_8 FILLER_26_156 ();
 sg13g2_decap_4 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_174 ();
 sg13g2_fill_1 FILLER_26_181 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_fill_2 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_230 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_fill_2 FILLER_26_346 ();
 sg13g2_fill_1 FILLER_26_348 ();
 sg13g2_fill_2 FILLER_26_353 ();
 sg13g2_fill_1 FILLER_26_381 ();
 sg13g2_fill_1 FILLER_26_390 ();
 sg13g2_fill_1 FILLER_26_395 ();
 sg13g2_fill_2 FILLER_26_401 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_4 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_46 ();
 sg13g2_decap_4 FILLER_27_94 ();
 sg13g2_fill_2 FILLER_27_98 ();
 sg13g2_fill_1 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_134 ();
 sg13g2_fill_2 FILLER_27_139 ();
 sg13g2_decap_4 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_179 ();
 sg13g2_decap_4 FILLER_27_195 ();
 sg13g2_decap_4 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_decap_4 FILLER_27_230 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_decap_4 FILLER_27_254 ();
 sg13g2_fill_1 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_268 ();
 sg13g2_decap_8 FILLER_27_274 ();
 sg13g2_fill_2 FILLER_27_281 ();
 sg13g2_decap_4 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_300 ();
 sg13g2_decap_8 FILLER_27_307 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_4 FILLER_27_330 ();
 sg13g2_decap_4 FILLER_27_338 ();
 sg13g2_fill_2 FILLER_27_342 ();
 sg13g2_fill_2 FILLER_27_369 ();
 sg13g2_fill_1 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_fill_2 FILLER_27_400 ();
 sg13g2_fill_1 FILLER_27_402 ();
 sg13g2_decap_4 FILLER_27_425 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_49 ();
 sg13g2_fill_2 FILLER_28_72 ();
 sg13g2_fill_1 FILLER_28_74 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_decap_4 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_fill_1 FILLER_28_113 ();
 sg13g2_decap_4 FILLER_28_130 ();
 sg13g2_fill_2 FILLER_28_134 ();
 sg13g2_decap_4 FILLER_28_160 ();
 sg13g2_fill_1 FILLER_28_164 ();
 sg13g2_decap_8 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_232 ();
 sg13g2_fill_1 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_decap_8 FILLER_28_254 ();
 sg13g2_fill_1 FILLER_28_261 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_decap_4 FILLER_28_275 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_decap_4 FILLER_28_284 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_327 ();
 sg13g2_fill_2 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_341 ();
 sg13g2_decap_4 FILLER_28_348 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_fill_2 FILLER_28_386 ();
 sg13g2_decap_4 FILLER_28_393 ();
 sg13g2_fill_2 FILLER_28_397 ();
 sg13g2_decap_8 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_411 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_4 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_46 ();
 sg13g2_decap_4 FILLER_29_72 ();
 sg13g2_fill_1 FILLER_29_80 ();
 sg13g2_decap_8 FILLER_29_86 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_fill_2 FILLER_29_133 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_decap_8 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_166 ();
 sg13g2_fill_2 FILLER_29_173 ();
 sg13g2_fill_1 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_193 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_decap_4 FILLER_29_216 ();
 sg13g2_fill_1 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_231 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_247 ();
 sg13g2_decap_8 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_261 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_decap_4 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_278 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_4 FILLER_29_315 ();
 sg13g2_fill_2 FILLER_29_323 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_fill_2 FILLER_29_357 ();
 sg13g2_fill_2 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_369 ();
 sg13g2_fill_1 FILLER_29_375 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_fill_1 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_413 ();
 sg13g2_decap_4 FILLER_29_424 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_58 ();
 sg13g2_fill_1 FILLER_30_65 ();
 sg13g2_decap_4 FILLER_30_96 ();
 sg13g2_fill_1 FILLER_30_100 ();
 sg13g2_fill_2 FILLER_30_105 ();
 sg13g2_fill_1 FILLER_30_107 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_decap_8 FILLER_30_122 ();
 sg13g2_decap_8 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_1 FILLER_30_157 ();
 sg13g2_decap_8 FILLER_30_163 ();
 sg13g2_decap_4 FILLER_30_170 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_216 ();
 sg13g2_decap_8 FILLER_30_223 ();
 sg13g2_fill_2 FILLER_30_230 ();
 sg13g2_fill_1 FILLER_30_235 ();
 sg13g2_decap_4 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_decap_4 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_267 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_decap_4 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_316 ();
 sg13g2_fill_2 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_fill_1 FILLER_30_335 ();
 sg13g2_fill_2 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_364 ();
 sg13g2_fill_2 FILLER_30_379 ();
 sg13g2_fill_2 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_4 FILLER_30_405 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_decap_4 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_74 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_decap_4 FILLER_31_89 ();
 sg13g2_fill_2 FILLER_31_120 ();
 sg13g2_fill_1 FILLER_31_127 ();
 sg13g2_decap_8 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_143 ();
 sg13g2_decap_8 FILLER_31_153 ();
 sg13g2_decap_8 FILLER_31_160 ();
 sg13g2_decap_4 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_240 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_fill_1 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_302 ();
 sg13g2_decap_8 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_fill_2 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_325 ();
 sg13g2_decap_4 FILLER_31_340 ();
 sg13g2_fill_1 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_349 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_fill_1 FILLER_31_369 ();
 sg13g2_decap_4 FILLER_31_389 ();
 sg13g2_fill_1 FILLER_31_393 ();
 sg13g2_fill_2 FILLER_31_409 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_fill_2 FILLER_31_427 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_59 ();
 sg13g2_fill_2 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_108 ();
 sg13g2_fill_2 FILLER_32_113 ();
 sg13g2_decap_4 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_138 ();
 sg13g2_decap_8 FILLER_32_149 ();
 sg13g2_decap_8 FILLER_32_156 ();
 sg13g2_decap_4 FILLER_32_163 ();
 sg13g2_decap_4 FILLER_32_171 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_fill_2 FILLER_32_192 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_265 ();
 sg13g2_fill_1 FILLER_32_274 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_fill_2 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_326 ();
 sg13g2_fill_1 FILLER_32_331 ();
 sg13g2_decap_8 FILLER_32_338 ();
 sg13g2_decap_8 FILLER_32_345 ();
 sg13g2_fill_2 FILLER_32_352 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_363 ();
 sg13g2_decap_4 FILLER_32_370 ();
 sg13g2_fill_2 FILLER_32_379 ();
 sg13g2_fill_1 FILLER_32_381 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_fill_1 FILLER_32_393 ();
 sg13g2_fill_2 FILLER_32_402 ();
 sg13g2_fill_1 FILLER_32_412 ();
 sg13g2_decap_8 FILLER_32_418 ();
 sg13g2_decap_4 FILLER_32_425 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_44 ();
 sg13g2_fill_2 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_71 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_79 ();
 sg13g2_fill_2 FILLER_33_85 ();
 sg13g2_fill_2 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_108 ();
 sg13g2_fill_2 FILLER_33_114 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_125 ();
 sg13g2_decap_8 FILLER_33_132 ();
 sg13g2_fill_2 FILLER_33_139 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_decap_8 FILLER_33_152 ();
 sg13g2_fill_2 FILLER_33_159 ();
 sg13g2_decap_4 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_181 ();
 sg13g2_fill_2 FILLER_33_193 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_232 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_fill_2 FILLER_33_281 ();
 sg13g2_decap_4 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_295 ();
 sg13g2_decap_8 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_309 ();
 sg13g2_decap_8 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_328 ();
 sg13g2_fill_1 FILLER_33_335 ();
 sg13g2_decap_8 FILLER_33_361 ();
 sg13g2_decap_8 FILLER_33_368 ();
 sg13g2_fill_2 FILLER_33_375 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_33_389 ();
 sg13g2_fill_1 FILLER_33_394 ();
 sg13g2_fill_2 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_47 ();
 sg13g2_fill_1 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_75 ();
 sg13g2_decap_8 FILLER_34_122 ();
 sg13g2_decap_4 FILLER_34_133 ();
 sg13g2_fill_1 FILLER_34_137 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_fill_1 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_4 FILLER_34_182 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_decap_4 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_decap_8 FILLER_34_221 ();
 sg13g2_decap_4 FILLER_34_228 ();
 sg13g2_fill_2 FILLER_34_232 ();
 sg13g2_fill_2 FILLER_34_255 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_269 ();
 sg13g2_fill_1 FILLER_34_271 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_fill_1 FILLER_34_307 ();
 sg13g2_fill_2 FILLER_34_330 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_decap_4 FILLER_34_377 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_decap_8 FILLER_34_415 ();
 sg13g2_decap_8 FILLER_34_422 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_4 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_46 ();
 sg13g2_fill_2 FILLER_35_59 ();
 sg13g2_fill_1 FILLER_35_61 ();
 sg13g2_decap_4 FILLER_35_88 ();
 sg13g2_fill_2 FILLER_35_92 ();
 sg13g2_decap_4 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_124 ();
 sg13g2_decap_8 FILLER_35_137 ();
 sg13g2_fill_2 FILLER_35_144 ();
 sg13g2_decap_4 FILLER_35_166 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_4 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_211 ();
 sg13g2_fill_1 FILLER_35_213 ();
 sg13g2_decap_8 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_225 ();
 sg13g2_decap_4 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_236 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_decap_4 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_decap_4 FILLER_35_316 ();
 sg13g2_fill_1 FILLER_35_320 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_decap_4 FILLER_35_335 ();
 sg13g2_fill_2 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_fill_2 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_368 ();
 sg13g2_fill_1 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_384 ();
 sg13g2_fill_1 FILLER_35_390 ();
 sg13g2_fill_1 FILLER_35_397 ();
 sg13g2_fill_1 FILLER_35_406 ();
 sg13g2_decap_4 FILLER_35_424 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_73 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_fill_2 FILLER_36_80 ();
 sg13g2_fill_1 FILLER_36_82 ();
 sg13g2_decap_8 FILLER_36_96 ();
 sg13g2_decap_4 FILLER_36_116 ();
 sg13g2_fill_2 FILLER_36_120 ();
 sg13g2_fill_2 FILLER_36_129 ();
 sg13g2_decap_8 FILLER_36_139 ();
 sg13g2_decap_8 FILLER_36_146 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_fill_2 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_181 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_decap_4 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_decap_4 FILLER_36_252 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_decap_4 FILLER_36_290 ();
 sg13g2_fill_2 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_307 ();
 sg13g2_fill_2 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_decap_4 FILLER_36_347 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_373 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_decap_4 FILLER_36_402 ();
 sg13g2_fill_1 FILLER_36_406 ();
 sg13g2_fill_2 FILLER_36_412 ();
 sg13g2_decap_4 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_81 ();
 sg13g2_decap_8 FILLER_37_88 ();
 sg13g2_fill_1 FILLER_37_95 ();
 sg13g2_decap_4 FILLER_37_100 ();
 sg13g2_decap_8 FILLER_37_114 ();
 sg13g2_decap_8 FILLER_37_121 ();
 sg13g2_decap_8 FILLER_37_128 ();
 sg13g2_decap_4 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_139 ();
 sg13g2_fill_1 FILLER_37_167 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_fill_1 FILLER_37_181 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_205 ();
 sg13g2_fill_1 FILLER_37_212 ();
 sg13g2_fill_2 FILLER_37_217 ();
 sg13g2_fill_1 FILLER_37_219 ();
 sg13g2_fill_2 FILLER_37_230 ();
 sg13g2_decap_4 FILLER_37_237 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_decap_8 FILLER_37_274 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_decap_8 FILLER_37_296 ();
 sg13g2_decap_4 FILLER_37_303 ();
 sg13g2_decap_8 FILLER_37_311 ();
 sg13g2_decap_4 FILLER_37_318 ();
 sg13g2_fill_2 FILLER_37_330 ();
 sg13g2_fill_2 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_339 ();
 sg13g2_decap_8 FILLER_37_349 ();
 sg13g2_fill_2 FILLER_37_356 ();
 sg13g2_decap_4 FILLER_37_374 ();
 sg13g2_decap_4 FILLER_37_382 ();
 sg13g2_fill_2 FILLER_37_391 ();
 sg13g2_fill_1 FILLER_37_393 ();
 sg13g2_fill_1 FILLER_37_400 ();
 sg13g2_fill_1 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_412 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_4 FILLER_38_49 ();
 sg13g2_fill_2 FILLER_38_57 ();
 sg13g2_fill_1 FILLER_38_59 ();
 sg13g2_fill_2 FILLER_38_74 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_99 ();
 sg13g2_fill_2 FILLER_38_103 ();
 sg13g2_fill_1 FILLER_38_114 ();
 sg13g2_decap_4 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_134 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_210 ();
 sg13g2_fill_2 FILLER_38_223 ();
 sg13g2_fill_2 FILLER_38_230 ();
 sg13g2_fill_1 FILLER_38_232 ();
 sg13g2_fill_2 FILLER_38_237 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_272 ();
 sg13g2_decap_8 FILLER_38_282 ();
 sg13g2_fill_2 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_300 ();
 sg13g2_fill_1 FILLER_38_307 ();
 sg13g2_fill_2 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_323 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_336 ();
 sg13g2_fill_2 FILLER_38_343 ();
 sg13g2_fill_2 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_fill_2 FILLER_38_371 ();
 sg13g2_fill_2 FILLER_38_379 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_4 FILLER_38_405 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_4 FILLER_39_49 ();
 sg13g2_fill_2 FILLER_39_53 ();
 sg13g2_fill_1 FILLER_39_85 ();
 sg13g2_fill_2 FILLER_39_117 ();
 sg13g2_decap_4 FILLER_39_127 ();
 sg13g2_fill_2 FILLER_39_131 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_fill_1 FILLER_39_147 ();
 sg13g2_decap_4 FILLER_39_153 ();
 sg13g2_fill_2 FILLER_39_157 ();
 sg13g2_decap_4 FILLER_39_164 ();
 sg13g2_fill_1 FILLER_39_178 ();
 sg13g2_fill_1 FILLER_39_189 ();
 sg13g2_fill_1 FILLER_39_195 ();
 sg13g2_fill_1 FILLER_39_201 ();
 sg13g2_fill_1 FILLER_39_206 ();
 sg13g2_fill_2 FILLER_39_216 ();
 sg13g2_fill_1 FILLER_39_218 ();
 sg13g2_fill_1 FILLER_39_232 ();
 sg13g2_decap_4 FILLER_39_241 ();
 sg13g2_fill_1 FILLER_39_245 ();
 sg13g2_fill_1 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_278 ();
 sg13g2_decap_8 FILLER_39_285 ();
 sg13g2_fill_1 FILLER_39_292 ();
 sg13g2_decap_8 FILLER_39_297 ();
 sg13g2_fill_1 FILLER_39_304 ();
 sg13g2_decap_4 FILLER_39_330 ();
 sg13g2_fill_1 FILLER_39_334 ();
 sg13g2_fill_2 FILLER_39_361 ();
 sg13g2_fill_1 FILLER_39_363 ();
 sg13g2_fill_1 FILLER_39_374 ();
 sg13g2_decap_8 FILLER_39_380 ();
 sg13g2_fill_1 FILLER_39_400 ();
 sg13g2_fill_1 FILLER_39_407 ();
 sg13g2_fill_1 FILLER_39_417 ();
 sg13g2_decap_4 FILLER_39_424 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_fill_2 FILLER_40_49 ();
 sg13g2_fill_1 FILLER_40_51 ();
 sg13g2_fill_1 FILLER_40_85 ();
 sg13g2_fill_1 FILLER_40_102 ();
 sg13g2_fill_1 FILLER_40_108 ();
 sg13g2_fill_1 FILLER_40_115 ();
 sg13g2_decap_8 FILLER_40_130 ();
 sg13g2_decap_8 FILLER_40_137 ();
 sg13g2_decap_4 FILLER_40_144 ();
 sg13g2_fill_2 FILLER_40_148 ();
 sg13g2_decap_8 FILLER_40_158 ();
 sg13g2_decap_8 FILLER_40_165 ();
 sg13g2_fill_2 FILLER_40_172 ();
 sg13g2_fill_2 FILLER_40_182 ();
 sg13g2_fill_2 FILLER_40_187 ();
 sg13g2_decap_8 FILLER_40_193 ();
 sg13g2_decap_4 FILLER_40_200 ();
 sg13g2_fill_2 FILLER_40_204 ();
 sg13g2_decap_4 FILLER_40_219 ();
 sg13g2_decap_8 FILLER_40_228 ();
 sg13g2_fill_1 FILLER_40_235 ();
 sg13g2_decap_8 FILLER_40_240 ();
 sg13g2_decap_8 FILLER_40_247 ();
 sg13g2_decap_8 FILLER_40_254 ();
 sg13g2_decap_8 FILLER_40_276 ();
 sg13g2_fill_1 FILLER_40_283 ();
 sg13g2_decap_8 FILLER_40_289 ();
 sg13g2_decap_8 FILLER_40_296 ();
 sg13g2_fill_2 FILLER_40_303 ();
 sg13g2_fill_1 FILLER_40_305 ();
 sg13g2_decap_8 FILLER_40_319 ();
 sg13g2_decap_8 FILLER_40_326 ();
 sg13g2_decap_4 FILLER_40_333 ();
 sg13g2_fill_1 FILLER_40_337 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_fill_2 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_362 ();
 sg13g2_fill_2 FILLER_40_369 ();
 sg13g2_fill_1 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_383 ();
 sg13g2_fill_1 FILLER_40_398 ();
 sg13g2_fill_1 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_409 ();
 sg13g2_fill_2 FILLER_40_415 ();
 sg13g2_fill_1 FILLER_40_417 ();
 sg13g2_decap_8 FILLER_40_423 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_4 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_46 ();
 sg13g2_fill_1 FILLER_41_53 ();
 sg13g2_fill_1 FILLER_41_63 ();
 sg13g2_fill_2 FILLER_41_94 ();
 sg13g2_fill_1 FILLER_41_96 ();
 sg13g2_fill_2 FILLER_41_123 ();
 sg13g2_decap_8 FILLER_41_139 ();
 sg13g2_fill_2 FILLER_41_146 ();
 sg13g2_fill_1 FILLER_41_148 ();
 sg13g2_decap_8 FILLER_41_162 ();
 sg13g2_decap_8 FILLER_41_169 ();
 sg13g2_fill_2 FILLER_41_190 ();
 sg13g2_decap_8 FILLER_41_200 ();
 sg13g2_fill_2 FILLER_41_207 ();
 sg13g2_fill_1 FILLER_41_209 ();
 sg13g2_decap_4 FILLER_41_220 ();
 sg13g2_fill_1 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_234 ();
 sg13g2_decap_4 FILLER_41_241 ();
 sg13g2_fill_2 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_251 ();
 sg13g2_fill_1 FILLER_41_258 ();
 sg13g2_decap_4 FILLER_41_267 ();
 sg13g2_fill_2 FILLER_41_271 ();
 sg13g2_decap_4 FILLER_41_306 ();
 sg13g2_decap_4 FILLER_41_323 ();
 sg13g2_fill_1 FILLER_41_327 ();
 sg13g2_decap_8 FILLER_41_338 ();
 sg13g2_fill_2 FILLER_41_366 ();
 sg13g2_fill_1 FILLER_41_368 ();
 sg13g2_fill_2 FILLER_41_387 ();
 sg13g2_fill_1 FILLER_41_394 ();
 sg13g2_fill_1 FILLER_41_407 ();
 sg13g2_decap_8 FILLER_41_423 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_4 FILLER_42_49 ();
 sg13g2_decap_4 FILLER_42_58 ();
 sg13g2_fill_2 FILLER_42_62 ();
 sg13g2_fill_1 FILLER_42_68 ();
 sg13g2_fill_2 FILLER_42_88 ();
 sg13g2_fill_1 FILLER_42_90 ();
 sg13g2_fill_2 FILLER_42_96 ();
 sg13g2_fill_1 FILLER_42_98 ();
 sg13g2_fill_1 FILLER_42_108 ();
 sg13g2_decap_8 FILLER_42_113 ();
 sg13g2_decap_8 FILLER_42_120 ();
 sg13g2_decap_4 FILLER_42_127 ();
 sg13g2_decap_8 FILLER_42_139 ();
 sg13g2_decap_4 FILLER_42_146 ();
 sg13g2_fill_2 FILLER_42_150 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_fill_2 FILLER_42_175 ();
 sg13g2_fill_1 FILLER_42_177 ();
 sg13g2_fill_1 FILLER_42_203 ();
 sg13g2_fill_1 FILLER_42_209 ();
 sg13g2_fill_1 FILLER_42_215 ();
 sg13g2_fill_1 FILLER_42_221 ();
 sg13g2_decap_4 FILLER_42_247 ();
 sg13g2_fill_2 FILLER_42_263 ();
 sg13g2_fill_2 FILLER_42_270 ();
 sg13g2_decap_4 FILLER_42_335 ();
 sg13g2_fill_2 FILLER_42_339 ();
 sg13g2_decap_8 FILLER_42_349 ();
 sg13g2_fill_2 FILLER_42_356 ();
 sg13g2_fill_2 FILLER_42_363 ();
 sg13g2_fill_1 FILLER_42_365 ();
 sg13g2_fill_1 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_411 ();
 sg13g2_decap_8 FILLER_42_418 ();
 sg13g2_decap_4 FILLER_42_425 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_4 FILLER_43_49 ();
 sg13g2_fill_1 FILLER_43_53 ();
 sg13g2_fill_1 FILLER_43_58 ();
 sg13g2_fill_2 FILLER_43_73 ();
 sg13g2_decap_4 FILLER_43_84 ();
 sg13g2_fill_1 FILLER_43_97 ();
 sg13g2_fill_1 FILLER_43_106 ();
 sg13g2_fill_1 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_117 ();
 sg13g2_decap_4 FILLER_43_124 ();
 sg13g2_decap_8 FILLER_43_132 ();
 sg13g2_decap_4 FILLER_43_171 ();
 sg13g2_fill_2 FILLER_43_184 ();
 sg13g2_fill_1 FILLER_43_186 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_fill_1 FILLER_43_209 ();
 sg13g2_fill_1 FILLER_43_215 ();
 sg13g2_decap_4 FILLER_43_223 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_decap_4 FILLER_43_233 ();
 sg13g2_fill_1 FILLER_43_237 ();
 sg13g2_decap_4 FILLER_43_242 ();
 sg13g2_fill_1 FILLER_43_254 ();
 sg13g2_fill_2 FILLER_43_259 ();
 sg13g2_fill_1 FILLER_43_261 ();
 sg13g2_fill_2 FILLER_43_267 ();
 sg13g2_decap_4 FILLER_43_275 ();
 sg13g2_decap_4 FILLER_43_302 ();
 sg13g2_fill_1 FILLER_43_306 ();
 sg13g2_decap_4 FILLER_43_318 ();
 sg13g2_fill_1 FILLER_43_337 ();
 sg13g2_decap_8 FILLER_43_348 ();
 sg13g2_decap_8 FILLER_43_355 ();
 sg13g2_fill_2 FILLER_43_362 ();
 sg13g2_fill_1 FILLER_43_364 ();
 sg13g2_decap_4 FILLER_43_369 ();
 sg13g2_fill_2 FILLER_43_373 ();
 sg13g2_decap_8 FILLER_43_416 ();
 sg13g2_decap_8 FILLER_43_423 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_fill_1 FILLER_44_71 ();
 sg13g2_fill_2 FILLER_44_95 ();
 sg13g2_fill_2 FILLER_44_101 ();
 sg13g2_decap_8 FILLER_44_124 ();
 sg13g2_decap_8 FILLER_44_135 ();
 sg13g2_fill_2 FILLER_44_142 ();
 sg13g2_fill_1 FILLER_44_152 ();
 sg13g2_decap_8 FILLER_44_167 ();
 sg13g2_decap_8 FILLER_44_174 ();
 sg13g2_decap_8 FILLER_44_181 ();
 sg13g2_decap_8 FILLER_44_188 ();
 sg13g2_decap_4 FILLER_44_195 ();
 sg13g2_fill_1 FILLER_44_199 ();
 sg13g2_fill_1 FILLER_44_204 ();
 sg13g2_decap_8 FILLER_44_209 ();
 sg13g2_fill_2 FILLER_44_224 ();
 sg13g2_fill_1 FILLER_44_226 ();
 sg13g2_decap_4 FILLER_44_232 ();
 sg13g2_fill_1 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_241 ();
 sg13g2_fill_1 FILLER_44_252 ();
 sg13g2_decap_4 FILLER_44_258 ();
 sg13g2_fill_1 FILLER_44_266 ();
 sg13g2_decap_4 FILLER_44_298 ();
 sg13g2_decap_8 FILLER_44_310 ();
 sg13g2_fill_2 FILLER_44_317 ();
 sg13g2_fill_1 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_358 ();
 sg13g2_decap_8 FILLER_44_365 ();
 sg13g2_decap_4 FILLER_44_372 ();
 sg13g2_fill_2 FILLER_44_376 ();
 sg13g2_fill_2 FILLER_44_382 ();
 sg13g2_decap_4 FILLER_44_389 ();
 sg13g2_fill_1 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_44_402 ();
 sg13g2_decap_8 FILLER_44_409 ();
 sg13g2_decap_8 FILLER_44_416 ();
 sg13g2_decap_8 FILLER_44_423 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_fill_2 FILLER_45_56 ();
 sg13g2_fill_1 FILLER_45_58 ();
 sg13g2_fill_2 FILLER_45_72 ();
 sg13g2_fill_1 FILLER_45_98 ();
 sg13g2_fill_2 FILLER_45_107 ();
 sg13g2_fill_1 FILLER_45_109 ();
 sg13g2_fill_2 FILLER_45_123 ();
 sg13g2_fill_1 FILLER_45_125 ();
 sg13g2_fill_1 FILLER_45_135 ();
 sg13g2_decap_8 FILLER_45_163 ();
 sg13g2_decap_8 FILLER_45_170 ();
 sg13g2_fill_2 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_decap_4 FILLER_45_186 ();
 sg13g2_decap_4 FILLER_45_198 ();
 sg13g2_fill_1 FILLER_45_202 ();
 sg13g2_fill_2 FILLER_45_212 ();
 sg13g2_fill_1 FILLER_45_214 ();
 sg13g2_fill_1 FILLER_45_223 ();
 sg13g2_fill_2 FILLER_45_230 ();
 sg13g2_fill_1 FILLER_45_232 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_4 FILLER_45_266 ();
 sg13g2_fill_1 FILLER_45_270 ();
 sg13g2_decap_8 FILLER_45_275 ();
 sg13g2_fill_1 FILLER_45_282 ();
 sg13g2_decap_4 FILLER_45_287 ();
 sg13g2_fill_1 FILLER_45_291 ();
 sg13g2_fill_2 FILLER_45_300 ();
 sg13g2_fill_1 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_306 ();
 sg13g2_fill_1 FILLER_45_312 ();
 sg13g2_decap_4 FILLER_45_318 ();
 sg13g2_fill_2 FILLER_45_322 ();
 sg13g2_decap_4 FILLER_45_337 ();
 sg13g2_decap_8 FILLER_45_360 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_fill_2 FILLER_45_427 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_fill_2 FILLER_46_49 ();
 sg13g2_fill_2 FILLER_46_61 ();
 sg13g2_fill_1 FILLER_46_77 ();
 sg13g2_fill_1 FILLER_46_84 ();
 sg13g2_fill_1 FILLER_46_93 ();
 sg13g2_fill_1 FILLER_46_99 ();
 sg13g2_decap_8 FILLER_46_104 ();
 sg13g2_decap_4 FILLER_46_111 ();
 sg13g2_fill_1 FILLER_46_115 ();
 sg13g2_fill_1 FILLER_46_121 ();
 sg13g2_fill_2 FILLER_46_128 ();
 sg13g2_fill_2 FILLER_46_135 ();
 sg13g2_fill_1 FILLER_46_137 ();
 sg13g2_fill_1 FILLER_46_142 ();
 sg13g2_fill_2 FILLER_46_161 ();
 sg13g2_fill_2 FILLER_46_189 ();
 sg13g2_fill_1 FILLER_46_191 ();
 sg13g2_decap_4 FILLER_46_199 ();
 sg13g2_fill_1 FILLER_46_203 ();
 sg13g2_fill_1 FILLER_46_212 ();
 sg13g2_decap_8 FILLER_46_257 ();
 sg13g2_decap_8 FILLER_46_264 ();
 sg13g2_decap_4 FILLER_46_271 ();
 sg13g2_fill_2 FILLER_46_275 ();
 sg13g2_decap_8 FILLER_46_282 ();
 sg13g2_decap_8 FILLER_46_319 ();
 sg13g2_fill_1 FILLER_46_326 ();
 sg13g2_fill_2 FILLER_46_332 ();
 sg13g2_decap_8 FILLER_46_341 ();
 sg13g2_decap_4 FILLER_46_361 ();
 sg13g2_decap_8 FILLER_46_382 ();
 sg13g2_decap_8 FILLER_46_389 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_decap_8 FILLER_46_403 ();
 sg13g2_decap_8 FILLER_46_410 ();
 sg13g2_decap_8 FILLER_46_417 ();
 sg13g2_decap_4 FILLER_46_424 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_63 ();
 sg13g2_fill_2 FILLER_47_69 ();
 sg13g2_fill_1 FILLER_47_71 ();
 sg13g2_fill_1 FILLER_47_80 ();
 sg13g2_fill_2 FILLER_47_90 ();
 sg13g2_fill_1 FILLER_47_110 ();
 sg13g2_fill_1 FILLER_47_115 ();
 sg13g2_decap_8 FILLER_47_120 ();
 sg13g2_fill_1 FILLER_47_127 ();
 sg13g2_fill_1 FILLER_47_132 ();
 sg13g2_decap_8 FILLER_47_148 ();
 sg13g2_fill_2 FILLER_47_155 ();
 sg13g2_fill_1 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_163 ();
 sg13g2_decap_4 FILLER_47_176 ();
 sg13g2_fill_2 FILLER_47_188 ();
 sg13g2_decap_4 FILLER_47_213 ();
 sg13g2_fill_1 FILLER_47_217 ();
 sg13g2_decap_4 FILLER_47_223 ();
 sg13g2_fill_2 FILLER_47_227 ();
 sg13g2_decap_4 FILLER_47_234 ();
 sg13g2_fill_1 FILLER_47_238 ();
 sg13g2_fill_2 FILLER_47_243 ();
 sg13g2_fill_1 FILLER_47_245 ();
 sg13g2_fill_1 FILLER_47_251 ();
 sg13g2_decap_8 FILLER_47_256 ();
 sg13g2_fill_1 FILLER_47_268 ();
 sg13g2_fill_2 FILLER_47_278 ();
 sg13g2_decap_8 FILLER_47_285 ();
 sg13g2_decap_8 FILLER_47_292 ();
 sg13g2_decap_8 FILLER_47_299 ();
 sg13g2_fill_2 FILLER_47_306 ();
 sg13g2_fill_1 FILLER_47_308 ();
 sg13g2_fill_1 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_320 ();
 sg13g2_fill_1 FILLER_47_325 ();
 sg13g2_decap_8 FILLER_47_335 ();
 sg13g2_decap_8 FILLER_47_347 ();
 sg13g2_decap_4 FILLER_47_354 ();
 sg13g2_fill_1 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_368 ();
 sg13g2_decap_8 FILLER_47_375 ();
 sg13g2_decap_8 FILLER_47_382 ();
 sg13g2_decap_8 FILLER_47_389 ();
 sg13g2_decap_8 FILLER_47_396 ();
 sg13g2_decap_8 FILLER_47_403 ();
 sg13g2_decap_8 FILLER_47_410 ();
 sg13g2_decap_8 FILLER_47_417 ();
 sg13g2_decap_4 FILLER_47_424 ();
 sg13g2_fill_2 FILLER_47_428 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_4 FILLER_48_70 ();
 sg13g2_fill_2 FILLER_48_82 ();
 sg13g2_fill_1 FILLER_48_84 ();
 sg13g2_fill_1 FILLER_48_89 ();
 sg13g2_decap_8 FILLER_48_99 ();
 sg13g2_decap_8 FILLER_48_106 ();
 sg13g2_decap_8 FILLER_48_113 ();
 sg13g2_fill_2 FILLER_48_120 ();
 sg13g2_decap_4 FILLER_48_131 ();
 sg13g2_fill_2 FILLER_48_135 ();
 sg13g2_decap_8 FILLER_48_142 ();
 sg13g2_fill_2 FILLER_48_149 ();
 sg13g2_fill_1 FILLER_48_151 ();
 sg13g2_decap_8 FILLER_48_157 ();
 sg13g2_fill_2 FILLER_48_164 ();
 sg13g2_fill_2 FILLER_48_171 ();
 sg13g2_fill_1 FILLER_48_173 ();
 sg13g2_fill_1 FILLER_48_187 ();
 sg13g2_fill_2 FILLER_48_192 ();
 sg13g2_fill_2 FILLER_48_202 ();
 sg13g2_fill_1 FILLER_48_204 ();
 sg13g2_fill_1 FILLER_48_209 ();
 sg13g2_decap_8 FILLER_48_236 ();
 sg13g2_decap_4 FILLER_48_243 ();
 sg13g2_fill_2 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_258 ();
 sg13g2_decap_8 FILLER_48_290 ();
 sg13g2_decap_8 FILLER_48_297 ();
 sg13g2_fill_1 FILLER_48_304 ();
 sg13g2_decap_8 FILLER_48_309 ();
 sg13g2_fill_2 FILLER_48_316 ();
 sg13g2_fill_1 FILLER_48_322 ();
 sg13g2_fill_2 FILLER_48_326 ();
 sg13g2_fill_1 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_354 ();
 sg13g2_fill_2 FILLER_48_361 ();
 sg13g2_fill_2 FILLER_48_368 ();
 sg13g2_decap_4 FILLER_48_375 ();
 sg13g2_fill_1 FILLER_48_379 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_fill_2 FILLER_48_392 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_decap_8 FILLER_48_400 ();
 sg13g2_decap_8 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_48_414 ();
 sg13g2_decap_8 FILLER_48_421 ();
 sg13g2_fill_2 FILLER_48_428 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_4 FILLER_49_70 ();
 sg13g2_fill_2 FILLER_49_74 ();
 sg13g2_fill_2 FILLER_49_80 ();
 sg13g2_decap_8 FILLER_49_87 ();
 sg13g2_fill_2 FILLER_49_94 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_4 FILLER_49_131 ();
 sg13g2_fill_1 FILLER_49_135 ();
 sg13g2_fill_1 FILLER_49_153 ();
 sg13g2_decap_8 FILLER_49_167 ();
 sg13g2_decap_8 FILLER_49_174 ();
 sg13g2_decap_8 FILLER_49_181 ();
 sg13g2_decap_8 FILLER_49_192 ();
 sg13g2_decap_4 FILLER_49_199 ();
 sg13g2_fill_1 FILLER_49_208 ();
 sg13g2_fill_1 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_fill_1 FILLER_49_256 ();
 sg13g2_fill_1 FILLER_49_261 ();
 sg13g2_decap_8 FILLER_49_267 ();
 sg13g2_fill_2 FILLER_49_274 ();
 sg13g2_fill_2 FILLER_49_296 ();
 sg13g2_decap_4 FILLER_49_302 ();
 sg13g2_decap_4 FILLER_49_310 ();
 sg13g2_fill_2 FILLER_49_314 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_fill_2 FILLER_49_364 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_decap_4 FILLER_49_371 ();
 sg13g2_fill_2 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_381 ();
 sg13g2_decap_4 FILLER_49_388 ();
 sg13g2_fill_1 FILLER_49_392 ();
 sg13g2_fill_2 FILLER_49_397 ();
 sg13g2_decap_8 FILLER_49_411 ();
 sg13g2_decap_8 FILLER_49_418 ();
 sg13g2_decap_4 FILLER_49_425 ();
 sg13g2_fill_1 FILLER_49_429 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_11 ();
 sg13g2_decap_8 FILLER_50_51 ();
 sg13g2_decap_8 FILLER_50_58 ();
 sg13g2_decap_8 FILLER_50_65 ();
 sg13g2_decap_8 FILLER_50_72 ();
 sg13g2_decap_8 FILLER_50_79 ();
 sg13g2_fill_2 FILLER_50_86 ();
 sg13g2_fill_1 FILLER_50_88 ();
 sg13g2_decap_4 FILLER_50_121 ();
 sg13g2_decap_4 FILLER_50_133 ();
 sg13g2_fill_1 FILLER_50_137 ();
 sg13g2_fill_1 FILLER_50_156 ();
 sg13g2_decap_8 FILLER_50_170 ();
 sg13g2_decap_8 FILLER_50_177 ();
 sg13g2_decap_8 FILLER_50_188 ();
 sg13g2_fill_2 FILLER_50_195 ();
 sg13g2_fill_1 FILLER_50_197 ();
 sg13g2_fill_2 FILLER_50_206 ();
 sg13g2_fill_1 FILLER_50_208 ();
 sg13g2_fill_1 FILLER_50_213 ();
 sg13g2_fill_1 FILLER_50_230 ();
 sg13g2_decap_8 FILLER_50_270 ();
 sg13g2_fill_1 FILLER_50_308 ();
 sg13g2_decap_4 FILLER_50_318 ();
 sg13g2_fill_1 FILLER_50_332 ();
 sg13g2_fill_2 FILLER_50_358 ();
 sg13g2_decap_8 FILLER_50_364 ();
 sg13g2_fill_2 FILLER_50_371 ();
 sg13g2_fill_1 FILLER_50_373 ();
 sg13g2_fill_1 FILLER_50_387 ();
 sg13g2_fill_1 FILLER_50_398 ();
 sg13g2_decap_8 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_50_415 ();
 sg13g2_decap_8 FILLER_50_422 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_fill_2 FILLER_51_42 ();
 sg13g2_fill_1 FILLER_51_44 ();
 sg13g2_fill_2 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_81 ();
 sg13g2_fill_2 FILLER_51_90 ();
 sg13g2_fill_1 FILLER_51_92 ();
 sg13g2_fill_2 FILLER_51_106 ();
 sg13g2_fill_1 FILLER_51_128 ();
 sg13g2_fill_1 FILLER_51_162 ();
 sg13g2_decap_4 FILLER_51_171 ();
 sg13g2_fill_1 FILLER_51_175 ();
 sg13g2_fill_1 FILLER_51_181 ();
 sg13g2_fill_2 FILLER_51_186 ();
 sg13g2_fill_2 FILLER_51_219 ();
 sg13g2_fill_1 FILLER_51_221 ();
 sg13g2_decap_4 FILLER_51_235 ();
 sg13g2_fill_2 FILLER_51_239 ();
 sg13g2_fill_2 FILLER_51_249 ();
 sg13g2_fill_1 FILLER_51_257 ();
 sg13g2_fill_2 FILLER_51_262 ();
 sg13g2_decap_4 FILLER_51_272 ();
 sg13g2_fill_1 FILLER_51_286 ();
 sg13g2_decap_4 FILLER_51_291 ();
 sg13g2_fill_2 FILLER_51_299 ();
 sg13g2_fill_1 FILLER_51_301 ();
 sg13g2_fill_1 FILLER_51_312 ();
 sg13g2_decap_8 FILLER_51_317 ();
 sg13g2_decap_8 FILLER_51_324 ();
 sg13g2_decap_8 FILLER_51_331 ();
 sg13g2_fill_1 FILLER_51_338 ();
 sg13g2_fill_1 FILLER_51_352 ();
 sg13g2_decap_8 FILLER_51_357 ();
 sg13g2_fill_1 FILLER_51_364 ();
 sg13g2_decap_4 FILLER_51_376 ();
 sg13g2_fill_1 FILLER_51_380 ();
 sg13g2_fill_1 FILLER_51_414 ();
 sg13g2_decap_4 FILLER_51_426 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_14 ();
 sg13g2_fill_1 FILLER_52_16 ();
 sg13g2_decap_8 FILLER_52_43 ();
 sg13g2_fill_1 FILLER_52_50 ();
 sg13g2_decap_8 FILLER_52_55 ();
 sg13g2_decap_4 FILLER_52_62 ();
 sg13g2_fill_2 FILLER_52_66 ();
 sg13g2_decap_8 FILLER_52_73 ();
 sg13g2_decap_8 FILLER_52_80 ();
 sg13g2_decap_8 FILLER_52_87 ();
 sg13g2_decap_4 FILLER_52_94 ();
 sg13g2_fill_2 FILLER_52_98 ();
 sg13g2_fill_1 FILLER_52_105 ();
 sg13g2_fill_1 FILLER_52_112 ();
 sg13g2_fill_1 FILLER_52_119 ();
 sg13g2_decap_4 FILLER_52_125 ();
 sg13g2_fill_2 FILLER_52_149 ();
 sg13g2_fill_1 FILLER_52_160 ();
 sg13g2_decap_4 FILLER_52_166 ();
 sg13g2_fill_2 FILLER_52_170 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_1 FILLER_52_187 ();
 sg13g2_decap_4 FILLER_52_193 ();
 sg13g2_decap_8 FILLER_52_201 ();
 sg13g2_decap_8 FILLER_52_208 ();
 sg13g2_decap_8 FILLER_52_215 ();
 sg13g2_decap_4 FILLER_52_237 ();
 sg13g2_decap_4 FILLER_52_245 ();
 sg13g2_fill_1 FILLER_52_249 ();
 sg13g2_decap_8 FILLER_52_258 ();
 sg13g2_decap_8 FILLER_52_265 ();
 sg13g2_fill_2 FILLER_52_272 ();
 sg13g2_decap_8 FILLER_52_295 ();
 sg13g2_decap_8 FILLER_52_302 ();
 sg13g2_decap_8 FILLER_52_313 ();
 sg13g2_decap_8 FILLER_52_320 ();
 sg13g2_decap_8 FILLER_52_327 ();
 sg13g2_decap_4 FILLER_52_334 ();
 sg13g2_fill_2 FILLER_52_338 ();
 sg13g2_decap_8 FILLER_52_348 ();
 sg13g2_decap_8 FILLER_52_355 ();
 sg13g2_fill_1 FILLER_52_362 ();
 sg13g2_decap_4 FILLER_52_367 ();
 sg13g2_fill_2 FILLER_52_371 ();
 sg13g2_decap_4 FILLER_52_378 ();
 sg13g2_fill_2 FILLER_52_387 ();
 sg13g2_fill_2 FILLER_52_399 ();
 sg13g2_decap_4 FILLER_52_424 ();
 sg13g2_fill_2 FILLER_52_428 ();
 sg13g2_fill_1 FILLER_53_26 ();
 sg13g2_decap_8 FILLER_53_34 ();
 sg13g2_decap_4 FILLER_53_41 ();
 sg13g2_fill_2 FILLER_53_45 ();
 sg13g2_fill_1 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_4 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_118 ();
 sg13g2_fill_2 FILLER_53_143 ();
 sg13g2_fill_1 FILLER_53_145 ();
 sg13g2_fill_2 FILLER_53_157 ();
 sg13g2_decap_8 FILLER_53_163 ();
 sg13g2_fill_2 FILLER_53_170 ();
 sg13g2_decap_8 FILLER_53_198 ();
 sg13g2_fill_2 FILLER_53_205 ();
 sg13g2_decap_8 FILLER_53_212 ();
 sg13g2_fill_2 FILLER_53_219 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_decap_4 FILLER_53_260 ();
 sg13g2_fill_1 FILLER_53_264 ();
 sg13g2_decap_4 FILLER_53_270 ();
 sg13g2_fill_1 FILLER_53_274 ();
 sg13g2_fill_1 FILLER_53_287 ();
 sg13g2_decap_8 FILLER_53_296 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_decap_8 FILLER_53_315 ();
 sg13g2_decap_8 FILLER_53_322 ();
 sg13g2_decap_8 FILLER_53_329 ();
 sg13g2_decap_8 FILLER_53_336 ();
 sg13g2_decap_8 FILLER_53_343 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_383 ();
 sg13g2_fill_2 FILLER_53_390 ();
 sg13g2_fill_1 FILLER_53_392 ();
 sg13g2_decap_4 FILLER_53_398 ();
 sg13g2_decap_8 FILLER_53_411 ();
 sg13g2_decap_8 FILLER_53_418 ();
 sg13g2_decap_4 FILLER_53_425 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_7 ();
 sg13g2_fill_1 FILLER_54_11 ();
 sg13g2_fill_2 FILLER_54_19 ();
 sg13g2_fill_1 FILLER_54_21 ();
 sg13g2_fill_2 FILLER_54_27 ();
 sg13g2_decap_8 FILLER_54_72 ();
 sg13g2_fill_2 FILLER_54_79 ();
 sg13g2_fill_1 FILLER_54_81 ();
 sg13g2_decap_4 FILLER_54_86 ();
 sg13g2_fill_2 FILLER_54_90 ();
 sg13g2_decap_8 FILLER_54_96 ();
 sg13g2_decap_8 FILLER_54_103 ();
 sg13g2_fill_2 FILLER_54_110 ();
 sg13g2_decap_8 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_132 ();
 sg13g2_decap_4 FILLER_54_143 ();
 sg13g2_fill_1 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_156 ();
 sg13g2_decap_8 FILLER_54_163 ();
 sg13g2_decap_8 FILLER_54_170 ();
 sg13g2_fill_1 FILLER_54_177 ();
 sg13g2_decap_8 FILLER_54_182 ();
 sg13g2_decap_4 FILLER_54_210 ();
 sg13g2_fill_2 FILLER_54_214 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_decap_8 FILLER_54_226 ();
 sg13g2_decap_8 FILLER_54_233 ();
 sg13g2_decap_8 FILLER_54_240 ();
 sg13g2_decap_8 FILLER_54_247 ();
 sg13g2_decap_8 FILLER_54_259 ();
 sg13g2_decap_8 FILLER_54_266 ();
 sg13g2_decap_8 FILLER_54_273 ();
 sg13g2_fill_2 FILLER_54_280 ();
 sg13g2_decap_8 FILLER_54_287 ();
 sg13g2_decap_4 FILLER_54_294 ();
 sg13g2_fill_1 FILLER_54_298 ();
 sg13g2_decap_8 FILLER_54_303 ();
 sg13g2_decap_4 FILLER_54_310 ();
 sg13g2_fill_2 FILLER_54_323 ();
 sg13g2_fill_1 FILLER_54_325 ();
 sg13g2_decap_8 FILLER_54_335 ();
 sg13g2_fill_2 FILLER_54_342 ();
 sg13g2_fill_1 FILLER_54_354 ();
 sg13g2_fill_2 FILLER_54_359 ();
 sg13g2_fill_1 FILLER_54_361 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_fill_2 FILLER_54_400 ();
 sg13g2_fill_1 FILLER_54_402 ();
 sg13g2_fill_1 FILLER_54_412 ();
 sg13g2_decap_8 FILLER_54_418 ();
 sg13g2_decap_4 FILLER_54_425 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_18 ();
 sg13g2_fill_1 FILLER_55_24 ();
 sg13g2_fill_1 FILLER_55_34 ();
 sg13g2_decap_8 FILLER_55_43 ();
 sg13g2_fill_2 FILLER_55_50 ();
 sg13g2_fill_1 FILLER_55_52 ();
 sg13g2_fill_1 FILLER_55_58 ();
 sg13g2_fill_1 FILLER_55_63 ();
 sg13g2_fill_1 FILLER_55_72 ();
 sg13g2_fill_1 FILLER_55_78 ();
 sg13g2_fill_2 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_97 ();
 sg13g2_fill_2 FILLER_55_104 ();
 sg13g2_fill_1 FILLER_55_106 ();
 sg13g2_fill_2 FILLER_55_112 ();
 sg13g2_fill_1 FILLER_55_114 ();
 sg13g2_decap_4 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_127 ();
 sg13g2_fill_2 FILLER_55_137 ();
 sg13g2_fill_1 FILLER_55_139 ();
 sg13g2_decap_8 FILLER_55_168 ();
 sg13g2_fill_2 FILLER_55_175 ();
 sg13g2_decap_4 FILLER_55_182 ();
 sg13g2_fill_1 FILLER_55_186 ();
 sg13g2_decap_8 FILLER_55_243 ();
 sg13g2_decap_8 FILLER_55_250 ();
 sg13g2_decap_8 FILLER_55_257 ();
 sg13g2_fill_2 FILLER_55_264 ();
 sg13g2_fill_1 FILLER_55_266 ();
 sg13g2_fill_1 FILLER_55_271 ();
 sg13g2_decap_4 FILLER_55_277 ();
 sg13g2_fill_1 FILLER_55_281 ();
 sg13g2_decap_8 FILLER_55_286 ();
 sg13g2_decap_8 FILLER_55_293 ();
 sg13g2_decap_8 FILLER_55_300 ();
 sg13g2_fill_2 FILLER_55_307 ();
 sg13g2_fill_1 FILLER_55_333 ();
 sg13g2_fill_1 FILLER_55_341 ();
 sg13g2_decap_4 FILLER_55_387 ();
 sg13g2_fill_1 FILLER_55_391 ();
 sg13g2_decap_4 FILLER_55_402 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_1 FILLER_55_414 ();
 sg13g2_decap_4 FILLER_55_426 ();
 sg13g2_decap_8 FILLER_56_31 ();
 sg13g2_decap_8 FILLER_56_38 ();
 sg13g2_decap_8 FILLER_56_45 ();
 sg13g2_decap_4 FILLER_56_52 ();
 sg13g2_fill_2 FILLER_56_82 ();
 sg13g2_fill_2 FILLER_56_133 ();
 sg13g2_fill_1 FILLER_56_135 ();
 sg13g2_fill_1 FILLER_56_149 ();
 sg13g2_fill_2 FILLER_56_163 ();
 sg13g2_decap_4 FILLER_56_169 ();
 sg13g2_fill_2 FILLER_56_173 ();
 sg13g2_fill_1 FILLER_56_185 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_fill_1 FILLER_56_201 ();
 sg13g2_decap_4 FILLER_56_220 ();
 sg13g2_fill_2 FILLER_56_228 ();
 sg13g2_fill_2 FILLER_56_257 ();
 sg13g2_fill_1 FILLER_56_259 ();
 sg13g2_decap_8 FILLER_56_269 ();
 sg13g2_decap_4 FILLER_56_276 ();
 sg13g2_fill_1 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_285 ();
 sg13g2_decap_8 FILLER_56_292 ();
 sg13g2_decap_8 FILLER_56_299 ();
 sg13g2_fill_2 FILLER_56_332 ();
 sg13g2_decap_8 FILLER_56_340 ();
 sg13g2_decap_8 FILLER_56_347 ();
 sg13g2_decap_4 FILLER_56_354 ();
 sg13g2_fill_1 FILLER_56_362 ();
 sg13g2_fill_1 FILLER_56_398 ();
 sg13g2_decap_4 FILLER_56_404 ();
 sg13g2_fill_2 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_56_421 ();
 sg13g2_fill_2 FILLER_56_428 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_18 ();
 sg13g2_decap_8 FILLER_57_27 ();
 sg13g2_decap_8 FILLER_57_34 ();
 sg13g2_fill_2 FILLER_57_41 ();
 sg13g2_decap_4 FILLER_57_51 ();
 sg13g2_fill_2 FILLER_57_55 ();
 sg13g2_fill_1 FILLER_57_66 ();
 sg13g2_fill_1 FILLER_57_75 ();
 sg13g2_decap_4 FILLER_57_81 ();
 sg13g2_fill_2 FILLER_57_90 ();
 sg13g2_fill_1 FILLER_57_92 ();
 sg13g2_fill_2 FILLER_57_98 ();
 sg13g2_fill_1 FILLER_57_100 ();
 sg13g2_fill_2 FILLER_57_106 ();
 sg13g2_fill_1 FILLER_57_135 ();
 sg13g2_fill_1 FILLER_57_141 ();
 sg13g2_decap_4 FILLER_57_150 ();
 sg13g2_fill_2 FILLER_57_158 ();
 sg13g2_fill_1 FILLER_57_170 ();
 sg13g2_decap_8 FILLER_57_202 ();
 sg13g2_decap_8 FILLER_57_209 ();
 sg13g2_decap_8 FILLER_57_216 ();
 sg13g2_decap_8 FILLER_57_223 ();
 sg13g2_decap_8 FILLER_57_230 ();
 sg13g2_fill_1 FILLER_57_237 ();
 sg13g2_fill_2 FILLER_57_243 ();
 sg13g2_decap_4 FILLER_57_250 ();
 sg13g2_fill_2 FILLER_57_258 ();
 sg13g2_decap_4 FILLER_57_268 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_fill_1 FILLER_57_280 ();
 sg13g2_fill_1 FILLER_57_285 ();
 sg13g2_fill_2 FILLER_57_299 ();
 sg13g2_fill_1 FILLER_57_314 ();
 sg13g2_fill_1 FILLER_57_324 ();
 sg13g2_decap_8 FILLER_57_335 ();
 sg13g2_fill_2 FILLER_57_342 ();
 sg13g2_fill_1 FILLER_57_363 ();
 sg13g2_fill_2 FILLER_57_369 ();
 sg13g2_fill_1 FILLER_57_371 ();
 sg13g2_fill_2 FILLER_57_392 ();
 sg13g2_fill_1 FILLER_57_410 ();
 sg13g2_decap_8 FILLER_57_421 ();
 sg13g2_fill_2 FILLER_57_428 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_15 ();
 sg13g2_fill_2 FILLER_58_19 ();
 sg13g2_fill_2 FILLER_58_25 ();
 sg13g2_fill_2 FILLER_58_35 ();
 sg13g2_fill_1 FILLER_58_45 ();
 sg13g2_fill_2 FILLER_58_66 ();
 sg13g2_decap_8 FILLER_58_94 ();
 sg13g2_decap_8 FILLER_58_101 ();
 sg13g2_fill_2 FILLER_58_108 ();
 sg13g2_fill_2 FILLER_58_126 ();
 sg13g2_fill_1 FILLER_58_128 ();
 sg13g2_decap_4 FILLER_58_134 ();
 sg13g2_fill_2 FILLER_58_142 ();
 sg13g2_decap_8 FILLER_58_149 ();
 sg13g2_decap_8 FILLER_58_156 ();
 sg13g2_decap_4 FILLER_58_163 ();
 sg13g2_fill_2 FILLER_58_167 ();
 sg13g2_fill_1 FILLER_58_174 ();
 sg13g2_fill_2 FILLER_58_189 ();
 sg13g2_fill_1 FILLER_58_191 ();
 sg13g2_fill_2 FILLER_58_209 ();
 sg13g2_fill_1 FILLER_58_211 ();
 sg13g2_fill_2 FILLER_58_217 ();
 sg13g2_fill_1 FILLER_58_219 ();
 sg13g2_fill_1 FILLER_58_228 ();
 sg13g2_decap_4 FILLER_58_242 ();
 sg13g2_fill_1 FILLER_58_255 ();
 sg13g2_fill_1 FILLER_58_261 ();
 sg13g2_fill_1 FILLER_58_278 ();
 sg13g2_fill_1 FILLER_58_291 ();
 sg13g2_fill_1 FILLER_58_297 ();
 sg13g2_fill_1 FILLER_58_303 ();
 sg13g2_fill_1 FILLER_58_327 ();
 sg13g2_fill_1 FILLER_58_333 ();
 sg13g2_decap_4 FILLER_58_343 ();
 sg13g2_fill_1 FILLER_58_347 ();
 sg13g2_fill_1 FILLER_58_352 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_2 FILLER_58_389 ();
 sg13g2_fill_2 FILLER_58_396 ();
 sg13g2_fill_1 FILLER_58_398 ();
 sg13g2_fill_2 FILLER_58_404 ();
 sg13g2_fill_1 FILLER_58_406 ();
 sg13g2_decap_8 FILLER_58_418 ();
 sg13g2_decap_4 FILLER_58_425 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_2 FILLER_59_31 ();
 sg13g2_fill_1 FILLER_59_33 ();
 sg13g2_fill_2 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_97 ();
 sg13g2_decap_8 FILLER_59_104 ();
 sg13g2_decap_4 FILLER_59_111 ();
 sg13g2_fill_1 FILLER_59_115 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_fill_2 FILLER_59_146 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_fill_2 FILLER_59_179 ();
 sg13g2_fill_1 FILLER_59_181 ();
 sg13g2_fill_2 FILLER_59_198 ();
 sg13g2_decap_8 FILLER_59_209 ();
 sg13g2_fill_2 FILLER_59_216 ();
 sg13g2_fill_2 FILLER_59_226 ();
 sg13g2_decap_8 FILLER_59_232 ();
 sg13g2_fill_2 FILLER_59_248 ();
 sg13g2_fill_2 FILLER_59_256 ();
 sg13g2_fill_2 FILLER_59_263 ();
 sg13g2_fill_1 FILLER_59_265 ();
 sg13g2_fill_1 FILLER_59_277 ();
 sg13g2_fill_2 FILLER_59_282 ();
 sg13g2_fill_2 FILLER_59_289 ();
 sg13g2_fill_2 FILLER_59_299 ();
 sg13g2_fill_1 FILLER_59_306 ();
 sg13g2_decap_4 FILLER_59_320 ();
 sg13g2_fill_2 FILLER_59_324 ();
 sg13g2_decap_8 FILLER_59_331 ();
 sg13g2_fill_2 FILLER_59_338 ();
 sg13g2_fill_1 FILLER_59_364 ();
 sg13g2_fill_1 FILLER_59_379 ();
 sg13g2_fill_1 FILLER_59_385 ();
 sg13g2_fill_1 FILLER_59_399 ();
 sg13g2_fill_2 FILLER_59_406 ();
 sg13g2_fill_1 FILLER_59_413 ();
 sg13g2_decap_8 FILLER_59_423 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_fill_1 FILLER_60_50 ();
 sg13g2_fill_2 FILLER_60_76 ();
 sg13g2_fill_2 FILLER_60_96 ();
 sg13g2_fill_1 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_104 ();
 sg13g2_decap_8 FILLER_60_111 ();
 sg13g2_decap_8 FILLER_60_118 ();
 sg13g2_decap_8 FILLER_60_125 ();
 sg13g2_fill_1 FILLER_60_152 ();
 sg13g2_decap_8 FILLER_60_162 ();
 sg13g2_decap_8 FILLER_60_169 ();
 sg13g2_decap_4 FILLER_60_180 ();
 sg13g2_fill_1 FILLER_60_184 ();
 sg13g2_decap_8 FILLER_60_208 ();
 sg13g2_decap_4 FILLER_60_215 ();
 sg13g2_fill_1 FILLER_60_219 ();
 sg13g2_fill_2 FILLER_60_225 ();
 sg13g2_fill_1 FILLER_60_227 ();
 sg13g2_decap_4 FILLER_60_234 ();
 sg13g2_fill_1 FILLER_60_238 ();
 sg13g2_fill_2 FILLER_60_245 ();
 sg13g2_fill_1 FILLER_60_247 ();
 sg13g2_fill_2 FILLER_60_253 ();
 sg13g2_fill_1 FILLER_60_255 ();
 sg13g2_fill_2 FILLER_60_261 ();
 sg13g2_fill_1 FILLER_60_263 ();
 sg13g2_decap_8 FILLER_60_270 ();
 sg13g2_fill_2 FILLER_60_277 ();
 sg13g2_fill_1 FILLER_60_279 ();
 sg13g2_fill_1 FILLER_60_285 ();
 sg13g2_decap_4 FILLER_60_290 ();
 sg13g2_fill_1 FILLER_60_298 ();
 sg13g2_decap_8 FILLER_60_313 ();
 sg13g2_decap_8 FILLER_60_320 ();
 sg13g2_fill_1 FILLER_60_327 ();
 sg13g2_fill_2 FILLER_60_341 ();
 sg13g2_fill_1 FILLER_60_343 ();
 sg13g2_decap_8 FILLER_60_356 ();
 sg13g2_decap_8 FILLER_60_363 ();
 sg13g2_decap_4 FILLER_60_370 ();
 sg13g2_fill_1 FILLER_60_383 ();
 sg13g2_fill_2 FILLER_60_404 ();
 sg13g2_fill_1 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_413 ();
 sg13g2_decap_4 FILLER_60_424 ();
 sg13g2_fill_2 FILLER_60_428 ();
 sg13g2_fill_2 FILLER_61_31 ();
 sg13g2_fill_1 FILLER_61_33 ();
 sg13g2_fill_1 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_53 ();
 sg13g2_decap_4 FILLER_61_60 ();
 sg13g2_decap_4 FILLER_61_75 ();
 sg13g2_fill_2 FILLER_61_88 ();
 sg13g2_decap_4 FILLER_61_94 ();
 sg13g2_fill_2 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_fill_1 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_178 ();
 sg13g2_fill_1 FILLER_61_199 ();
 sg13g2_fill_2 FILLER_61_205 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_fill_2 FILLER_61_233 ();
 sg13g2_decap_4 FILLER_61_256 ();
 sg13g2_fill_2 FILLER_61_265 ();
 sg13g2_fill_2 FILLER_61_280 ();
 sg13g2_decap_4 FILLER_61_296 ();
 sg13g2_fill_1 FILLER_61_300 ();
 sg13g2_decap_4 FILLER_61_319 ();
 sg13g2_fill_1 FILLER_61_323 ();
 sg13g2_decap_8 FILLER_61_338 ();
 sg13g2_decap_8 FILLER_61_345 ();
 sg13g2_decap_8 FILLER_61_352 ();
 sg13g2_decap_8 FILLER_61_363 ();
 sg13g2_fill_1 FILLER_61_370 ();
 sg13g2_decap_4 FILLER_61_374 ();
 sg13g2_fill_1 FILLER_61_392 ();
 sg13g2_fill_2 FILLER_61_407 ();
 sg13g2_decap_4 FILLER_61_426 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_16 ();
 sg13g2_fill_1 FILLER_62_18 ();
 sg13g2_decap_8 FILLER_62_31 ();
 sg13g2_decap_8 FILLER_62_38 ();
 sg13g2_decap_4 FILLER_62_45 ();
 sg13g2_fill_1 FILLER_62_49 ();
 sg13g2_fill_2 FILLER_62_55 ();
 sg13g2_fill_1 FILLER_62_57 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_fill_1 FILLER_62_79 ();
 sg13g2_decap_8 FILLER_62_122 ();
 sg13g2_fill_1 FILLER_62_129 ();
 sg13g2_decap_4 FILLER_62_190 ();
 sg13g2_decap_8 FILLER_62_206 ();
 sg13g2_decap_4 FILLER_62_213 ();
 sg13g2_fill_1 FILLER_62_217 ();
 sg13g2_decap_8 FILLER_62_226 ();
 sg13g2_decap_8 FILLER_62_233 ();
 sg13g2_fill_1 FILLER_62_240 ();
 sg13g2_decap_4 FILLER_62_246 ();
 sg13g2_fill_1 FILLER_62_250 ();
 sg13g2_decap_8 FILLER_62_267 ();
 sg13g2_fill_1 FILLER_62_282 ();
 sg13g2_fill_1 FILLER_62_288 ();
 sg13g2_fill_2 FILLER_62_295 ();
 sg13g2_fill_2 FILLER_62_303 ();
 sg13g2_fill_2 FILLER_62_309 ();
 sg13g2_decap_4 FILLER_62_334 ();
 sg13g2_fill_2 FILLER_62_338 ();
 sg13g2_decap_8 FILLER_62_346 ();
 sg13g2_fill_2 FILLER_62_353 ();
 sg13g2_fill_2 FILLER_62_372 ();
 sg13g2_decap_4 FILLER_62_390 ();
 sg13g2_decap_8 FILLER_62_403 ();
 sg13g2_fill_2 FILLER_62_410 ();
 sg13g2_decap_8 FILLER_62_417 ();
 sg13g2_decap_4 FILLER_62_424 ();
 sg13g2_fill_2 FILLER_62_428 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_9 ();
 sg13g2_fill_2 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_34 ();
 sg13g2_fill_1 FILLER_63_41 ();
 sg13g2_decap_4 FILLER_63_50 ();
 sg13g2_fill_1 FILLER_63_54 ();
 sg13g2_decap_4 FILLER_63_65 ();
 sg13g2_fill_1 FILLER_63_81 ();
 sg13g2_fill_1 FILLER_63_95 ();
 sg13g2_decap_8 FILLER_63_100 ();
 sg13g2_decap_8 FILLER_63_107 ();
 sg13g2_decap_8 FILLER_63_114 ();
 sg13g2_decap_8 FILLER_63_121 ();
 sg13g2_decap_8 FILLER_63_128 ();
 sg13g2_decap_8 FILLER_63_135 ();
 sg13g2_decap_8 FILLER_63_142 ();
 sg13g2_fill_2 FILLER_63_149 ();
 sg13g2_fill_1 FILLER_63_151 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_63_194 ();
 sg13g2_fill_2 FILLER_63_201 ();
 sg13g2_fill_1 FILLER_63_203 ();
 sg13g2_fill_2 FILLER_63_222 ();
 sg13g2_decap_8 FILLER_63_228 ();
 sg13g2_fill_1 FILLER_63_276 ();
 sg13g2_fill_1 FILLER_63_281 ();
 sg13g2_decap_4 FILLER_63_294 ();
 sg13g2_fill_1 FILLER_63_298 ();
 sg13g2_decap_4 FILLER_63_303 ();
 sg13g2_fill_1 FILLER_63_307 ();
 sg13g2_decap_4 FILLER_63_324 ();
 sg13g2_fill_1 FILLER_63_328 ();
 sg13g2_decap_8 FILLER_63_334 ();
 sg13g2_fill_2 FILLER_63_341 ();
 sg13g2_decap_8 FILLER_63_349 ();
 sg13g2_fill_2 FILLER_63_361 ();
 sg13g2_fill_2 FILLER_63_416 ();
 sg13g2_decap_8 FILLER_63_423 ();
 sg13g2_decap_8 FILLER_64_39 ();
 sg13g2_fill_2 FILLER_64_46 ();
 sg13g2_fill_1 FILLER_64_48 ();
 sg13g2_fill_2 FILLER_64_90 ();
 sg13g2_fill_1 FILLER_64_92 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_4 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_120 ();
 sg13g2_decap_4 FILLER_64_127 ();
 sg13g2_decap_8 FILLER_64_135 ();
 sg13g2_fill_1 FILLER_64_151 ();
 sg13g2_fill_2 FILLER_64_156 ();
 sg13g2_fill_1 FILLER_64_158 ();
 sg13g2_decap_4 FILLER_64_163 ();
 sg13g2_fill_1 FILLER_64_167 ();
 sg13g2_decap_8 FILLER_64_181 ();
 sg13g2_decap_4 FILLER_64_188 ();
 sg13g2_fill_1 FILLER_64_192 ();
 sg13g2_fill_2 FILLER_64_206 ();
 sg13g2_fill_1 FILLER_64_239 ();
 sg13g2_decap_4 FILLER_64_257 ();
 sg13g2_fill_2 FILLER_64_271 ();
 sg13g2_fill_1 FILLER_64_300 ();
 sg13g2_fill_2 FILLER_64_311 ();
 sg13g2_fill_2 FILLER_64_318 ();
 sg13g2_fill_1 FILLER_64_320 ();
 sg13g2_fill_1 FILLER_64_331 ();
 sg13g2_decap_4 FILLER_64_342 ();
 sg13g2_fill_1 FILLER_64_346 ();
 sg13g2_fill_1 FILLER_64_362 ();
 sg13g2_fill_2 FILLER_64_367 ();
 sg13g2_fill_1 FILLER_64_369 ();
 sg13g2_fill_2 FILLER_64_385 ();
 sg13g2_fill_2 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_415 ();
 sg13g2_decap_8 FILLER_64_422 ();
 sg13g2_fill_1 FILLER_64_429 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_11 ();
 sg13g2_fill_1 FILLER_65_42 ();
 sg13g2_fill_1 FILLER_65_47 ();
 sg13g2_fill_1 FILLER_65_88 ();
 sg13g2_decap_8 FILLER_65_125 ();
 sg13g2_decap_8 FILLER_65_132 ();
 sg13g2_decap_4 FILLER_65_158 ();
 sg13g2_fill_2 FILLER_65_162 ();
 sg13g2_decap_8 FILLER_65_201 ();
 sg13g2_decap_8 FILLER_65_208 ();
 sg13g2_decap_4 FILLER_65_215 ();
 sg13g2_fill_2 FILLER_65_219 ();
 sg13g2_fill_2 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_250 ();
 sg13g2_decap_4 FILLER_65_257 ();
 sg13g2_fill_2 FILLER_65_261 ();
 sg13g2_fill_2 FILLER_65_268 ();
 sg13g2_fill_1 FILLER_65_270 ();
 sg13g2_decap_8 FILLER_65_295 ();
 sg13g2_decap_4 FILLER_65_302 ();
 sg13g2_fill_1 FILLER_65_312 ();
 sg13g2_fill_1 FILLER_65_318 ();
 sg13g2_decap_4 FILLER_65_329 ();
 sg13g2_decap_4 FILLER_65_344 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_fill_2 FILLER_65_376 ();
 sg13g2_fill_1 FILLER_65_391 ();
 sg13g2_fill_1 FILLER_65_398 ();
 sg13g2_fill_1 FILLER_65_404 ();
 sg13g2_decap_8 FILLER_65_421 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_4 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_18 ();
 sg13g2_fill_1 FILLER_66_51 ();
 sg13g2_fill_2 FILLER_66_56 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_decap_8 FILLER_66_94 ();
 sg13g2_decap_4 FILLER_66_101 ();
 sg13g2_fill_1 FILLER_66_105 ();
 sg13g2_fill_2 FILLER_66_114 ();
 sg13g2_fill_1 FILLER_66_147 ();
 sg13g2_fill_2 FILLER_66_156 ();
 sg13g2_decap_8 FILLER_66_162 ();
 sg13g2_fill_1 FILLER_66_169 ();
 sg13g2_fill_1 FILLER_66_174 ();
 sg13g2_fill_2 FILLER_66_180 ();
 sg13g2_fill_1 FILLER_66_187 ();
 sg13g2_fill_2 FILLER_66_193 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_fill_1 FILLER_66_217 ();
 sg13g2_decap_4 FILLER_66_232 ();
 sg13g2_fill_2 FILLER_66_236 ();
 sg13g2_decap_8 FILLER_66_254 ();
 sg13g2_decap_8 FILLER_66_270 ();
 sg13g2_decap_8 FILLER_66_277 ();
 sg13g2_fill_2 FILLER_66_284 ();
 sg13g2_fill_1 FILLER_66_286 ();
 sg13g2_decap_4 FILLER_66_292 ();
 sg13g2_fill_1 FILLER_66_296 ();
 sg13g2_fill_1 FILLER_66_311 ();
 sg13g2_fill_1 FILLER_66_320 ();
 sg13g2_decap_8 FILLER_66_341 ();
 sg13g2_decap_4 FILLER_66_348 ();
 sg13g2_fill_1 FILLER_66_352 ();
 sg13g2_decap_8 FILLER_66_362 ();
 sg13g2_decap_4 FILLER_66_369 ();
 sg13g2_fill_2 FILLER_66_373 ();
 sg13g2_fill_1 FILLER_66_379 ();
 sg13g2_fill_1 FILLER_66_384 ();
 sg13g2_decap_4 FILLER_66_389 ();
 sg13g2_fill_2 FILLER_66_393 ();
 sg13g2_fill_2 FILLER_66_400 ();
 sg13g2_fill_1 FILLER_66_402 ();
 sg13g2_fill_2 FILLER_66_408 ();
 sg13g2_fill_1 FILLER_66_410 ();
 sg13g2_decap_8 FILLER_66_416 ();
 sg13g2_decap_8 FILLER_66_423 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_4 FILLER_67_63 ();
 sg13g2_fill_2 FILLER_67_72 ();
 sg13g2_decap_8 FILLER_67_78 ();
 sg13g2_decap_8 FILLER_67_85 ();
 sg13g2_decap_8 FILLER_67_92 ();
 sg13g2_decap_4 FILLER_67_99 ();
 sg13g2_fill_2 FILLER_67_103 ();
 sg13g2_decap_8 FILLER_67_139 ();
 sg13g2_decap_4 FILLER_67_146 ();
 sg13g2_fill_1 FILLER_67_150 ();
 sg13g2_fill_2 FILLER_67_181 ();
 sg13g2_fill_2 FILLER_67_203 ();
 sg13g2_fill_1 FILLER_67_205 ();
 sg13g2_decap_4 FILLER_67_214 ();
 sg13g2_decap_4 FILLER_67_223 ();
 sg13g2_fill_2 FILLER_67_227 ();
 sg13g2_decap_4 FILLER_67_234 ();
 sg13g2_fill_1 FILLER_67_238 ();
 sg13g2_fill_2 FILLER_67_244 ();
 sg13g2_fill_1 FILLER_67_246 ();
 sg13g2_fill_2 FILLER_67_267 ();
 sg13g2_decap_8 FILLER_67_290 ();
 sg13g2_fill_2 FILLER_67_297 ();
 sg13g2_fill_1 FILLER_67_299 ();
 sg13g2_decap_4 FILLER_67_328 ();
 sg13g2_fill_2 FILLER_67_352 ();
 sg13g2_decap_4 FILLER_67_358 ();
 sg13g2_fill_2 FILLER_67_362 ();
 sg13g2_fill_1 FILLER_67_377 ();
 sg13g2_fill_2 FILLER_67_393 ();
 sg13g2_fill_1 FILLER_67_404 ();
 sg13g2_decap_8 FILLER_67_410 ();
 sg13g2_decap_8 FILLER_67_417 ();
 sg13g2_decap_4 FILLER_67_424 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_fill_2 FILLER_68_21 ();
 sg13g2_decap_4 FILLER_68_60 ();
 sg13g2_decap_8 FILLER_68_69 ();
 sg13g2_decap_8 FILLER_68_76 ();
 sg13g2_fill_2 FILLER_68_83 ();
 sg13g2_fill_2 FILLER_68_97 ();
 sg13g2_fill_2 FILLER_68_102 ();
 sg13g2_fill_1 FILLER_68_111 ();
 sg13g2_decap_8 FILLER_68_116 ();
 sg13g2_decap_4 FILLER_68_123 ();
 sg13g2_fill_1 FILLER_68_127 ();
 sg13g2_decap_8 FILLER_68_132 ();
 sg13g2_fill_1 FILLER_68_139 ();
 sg13g2_decap_4 FILLER_68_148 ();
 sg13g2_fill_2 FILLER_68_152 ();
 sg13g2_decap_8 FILLER_68_159 ();
 sg13g2_decap_8 FILLER_68_166 ();
 sg13g2_decap_4 FILLER_68_177 ();
 sg13g2_fill_1 FILLER_68_181 ();
 sg13g2_decap_4 FILLER_68_187 ();
 sg13g2_decap_8 FILLER_68_204 ();
 sg13g2_decap_8 FILLER_68_211 ();
 sg13g2_decap_8 FILLER_68_218 ();
 sg13g2_decap_8 FILLER_68_225 ();
 sg13g2_decap_8 FILLER_68_232 ();
 sg13g2_decap_8 FILLER_68_239 ();
 sg13g2_fill_2 FILLER_68_246 ();
 sg13g2_fill_2 FILLER_68_260 ();
 sg13g2_fill_1 FILLER_68_262 ();
 sg13g2_decap_4 FILLER_68_291 ();
 sg13g2_decap_8 FILLER_68_326 ();
 sg13g2_decap_8 FILLER_68_333 ();
 sg13g2_decap_4 FILLER_68_340 ();
 sg13g2_decap_4 FILLER_68_358 ();
 sg13g2_fill_2 FILLER_68_362 ();
 sg13g2_fill_1 FILLER_68_380 ();
 sg13g2_decap_4 FILLER_68_385 ();
 sg13g2_fill_1 FILLER_68_404 ();
 sg13g2_decap_8 FILLER_68_410 ();
 sg13g2_decap_8 FILLER_68_417 ();
 sg13g2_decap_4 FILLER_68_424 ();
 sg13g2_fill_2 FILLER_68_428 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_38 ();
 sg13g2_decap_8 FILLER_69_45 ();
 sg13g2_decap_8 FILLER_69_52 ();
 sg13g2_decap_8 FILLER_69_67 ();
 sg13g2_decap_8 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_81 ();
 sg13g2_decap_8 FILLER_69_113 ();
 sg13g2_decap_8 FILLER_69_120 ();
 sg13g2_fill_1 FILLER_69_127 ();
 sg13g2_decap_4 FILLER_69_136 ();
 sg13g2_fill_1 FILLER_69_140 ();
 sg13g2_decap_4 FILLER_69_153 ();
 sg13g2_fill_1 FILLER_69_157 ();
 sg13g2_decap_8 FILLER_69_162 ();
 sg13g2_decap_8 FILLER_69_169 ();
 sg13g2_fill_2 FILLER_69_176 ();
 sg13g2_fill_1 FILLER_69_178 ();
 sg13g2_decap_8 FILLER_69_183 ();
 sg13g2_fill_2 FILLER_69_190 ();
 sg13g2_fill_2 FILLER_69_197 ();
 sg13g2_fill_2 FILLER_69_203 ();
 sg13g2_fill_1 FILLER_69_205 ();
 sg13g2_decap_8 FILLER_69_214 ();
 sg13g2_decap_8 FILLER_69_221 ();
 sg13g2_decap_8 FILLER_69_228 ();
 sg13g2_decap_8 FILLER_69_235 ();
 sg13g2_decap_8 FILLER_69_242 ();
 sg13g2_decap_8 FILLER_69_249 ();
 sg13g2_decap_4 FILLER_69_256 ();
 sg13g2_fill_2 FILLER_69_260 ();
 sg13g2_decap_4 FILLER_69_275 ();
 sg13g2_fill_1 FILLER_69_279 ();
 sg13g2_decap_8 FILLER_69_289 ();
 sg13g2_decap_8 FILLER_69_296 ();
 sg13g2_decap_4 FILLER_69_313 ();
 sg13g2_fill_2 FILLER_69_317 ();
 sg13g2_decap_8 FILLER_69_324 ();
 sg13g2_fill_1 FILLER_69_331 ();
 sg13g2_fill_2 FILLER_69_341 ();
 sg13g2_fill_2 FILLER_69_383 ();
 sg13g2_decap_4 FILLER_69_403 ();
 sg13g2_decap_8 FILLER_69_412 ();
 sg13g2_decap_8 FILLER_69_419 ();
 sg13g2_decap_4 FILLER_69_426 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_4 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_40 ();
 sg13g2_decap_8 FILLER_70_47 ();
 sg13g2_decap_8 FILLER_70_54 ();
 sg13g2_fill_2 FILLER_70_61 ();
 sg13g2_decap_8 FILLER_70_92 ();
 sg13g2_decap_4 FILLER_70_125 ();
 sg13g2_decap_4 FILLER_70_181 ();
 sg13g2_fill_2 FILLER_70_185 ();
 sg13g2_decap_8 FILLER_70_202 ();
 sg13g2_fill_1 FILLER_70_209 ();
 sg13g2_decap_8 FILLER_70_218 ();
 sg13g2_decap_4 FILLER_70_233 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_decap_8 FILLER_70_243 ();
 sg13g2_decap_8 FILLER_70_250 ();
 sg13g2_decap_8 FILLER_70_257 ();
 sg13g2_decap_4 FILLER_70_264 ();
 sg13g2_fill_2 FILLER_70_268 ();
 sg13g2_fill_2 FILLER_70_297 ();
 sg13g2_fill_1 FILLER_70_304 ();
 sg13g2_fill_2 FILLER_70_320 ();
 sg13g2_decap_4 FILLER_70_328 ();
 sg13g2_fill_1 FILLER_70_332 ();
 sg13g2_fill_1 FILLER_70_347 ();
 sg13g2_fill_1 FILLER_70_364 ();
 sg13g2_fill_1 FILLER_70_371 ();
 sg13g2_fill_1 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_404 ();
 sg13g2_decap_4 FILLER_70_424 ();
 sg13g2_fill_2 FILLER_70_428 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_4 FILLER_71_21 ();
 sg13g2_fill_2 FILLER_71_25 ();
 sg13g2_fill_2 FILLER_71_31 ();
 sg13g2_fill_2 FILLER_71_79 ();
 sg13g2_decap_4 FILLER_71_98 ();
 sg13g2_fill_2 FILLER_71_121 ();
 sg13g2_fill_1 FILLER_71_133 ();
 sg13g2_fill_2 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_4 FILLER_71_182 ();
 sg13g2_fill_1 FILLER_71_186 ();
 sg13g2_decap_8 FILLER_71_220 ();
 sg13g2_decap_8 FILLER_71_227 ();
 sg13g2_fill_2 FILLER_71_234 ();
 sg13g2_fill_2 FILLER_71_245 ();
 sg13g2_fill_1 FILLER_71_247 ();
 sg13g2_decap_8 FILLER_71_253 ();
 sg13g2_decap_8 FILLER_71_260 ();
 sg13g2_decap_8 FILLER_71_267 ();
 sg13g2_fill_2 FILLER_71_274 ();
 sg13g2_fill_1 FILLER_71_276 ();
 sg13g2_fill_2 FILLER_71_317 ();
 sg13g2_fill_1 FILLER_71_319 ();
 sg13g2_fill_2 FILLER_71_337 ();
 sg13g2_fill_1 FILLER_71_339 ();
 sg13g2_fill_1 FILLER_71_344 ();
 sg13g2_fill_1 FILLER_71_352 ();
 sg13g2_fill_1 FILLER_71_358 ();
 sg13g2_fill_2 FILLER_71_364 ();
 sg13g2_fill_2 FILLER_71_370 ();
 sg13g2_fill_1 FILLER_71_372 ();
 sg13g2_fill_1 FILLER_71_392 ();
 sg13g2_fill_1 FILLER_71_398 ();
 sg13g2_fill_1 FILLER_71_403 ();
 sg13g2_fill_1 FILLER_71_423 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_fill_2 FILLER_72_30 ();
 sg13g2_fill_1 FILLER_72_32 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_fill_1 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_83 ();
 sg13g2_decap_8 FILLER_72_90 ();
 sg13g2_fill_2 FILLER_72_97 ();
 sg13g2_fill_1 FILLER_72_99 ();
 sg13g2_decap_4 FILLER_72_109 ();
 sg13g2_decap_8 FILLER_72_139 ();
 sg13g2_fill_2 FILLER_72_146 ();
 sg13g2_fill_1 FILLER_72_148 ();
 sg13g2_decap_4 FILLER_72_155 ();
 sg13g2_decap_8 FILLER_72_167 ();
 sg13g2_fill_2 FILLER_72_174 ();
 sg13g2_decap_8 FILLER_72_183 ();
 sg13g2_decap_4 FILLER_72_190 ();
 sg13g2_fill_2 FILLER_72_194 ();
 sg13g2_fill_1 FILLER_72_236 ();
 sg13g2_fill_1 FILLER_72_248 ();
 sg13g2_fill_2 FILLER_72_252 ();
 sg13g2_fill_1 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_264 ();
 sg13g2_decap_8 FILLER_72_271 ();
 sg13g2_decap_8 FILLER_72_278 ();
 sg13g2_decap_8 FILLER_72_285 ();
 sg13g2_decap_8 FILLER_72_296 ();
 sg13g2_decap_8 FILLER_72_303 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_4 FILLER_72_322 ();
 sg13g2_fill_2 FILLER_72_330 ();
 sg13g2_fill_1 FILLER_72_332 ();
 sg13g2_fill_1 FILLER_72_341 ();
 sg13g2_fill_1 FILLER_72_347 ();
 sg13g2_fill_1 FILLER_72_353 ();
 sg13g2_fill_1 FILLER_72_358 ();
 sg13g2_fill_1 FILLER_72_364 ();
 sg13g2_fill_2 FILLER_72_381 ();
 sg13g2_fill_1 FILLER_72_383 ();
 sg13g2_fill_2 FILLER_72_389 ();
 sg13g2_decap_4 FILLER_72_412 ();
 sg13g2_decap_8 FILLER_72_422 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_41 ();
 sg13g2_decap_8 FILLER_73_69 ();
 sg13g2_decap_8 FILLER_73_76 ();
 sg13g2_decap_8 FILLER_73_83 ();
 sg13g2_decap_8 FILLER_73_90 ();
 sg13g2_decap_8 FILLER_73_97 ();
 sg13g2_decap_4 FILLER_73_104 ();
 sg13g2_decap_8 FILLER_73_116 ();
 sg13g2_decap_8 FILLER_73_123 ();
 sg13g2_decap_8 FILLER_73_130 ();
 sg13g2_decap_8 FILLER_73_137 ();
 sg13g2_decap_8 FILLER_73_144 ();
 sg13g2_decap_8 FILLER_73_151 ();
 sg13g2_decap_8 FILLER_73_158 ();
 sg13g2_decap_8 FILLER_73_165 ();
 sg13g2_decap_8 FILLER_73_172 ();
 sg13g2_decap_4 FILLER_73_179 ();
 sg13g2_fill_1 FILLER_73_183 ();
 sg13g2_decap_8 FILLER_73_197 ();
 sg13g2_decap_8 FILLER_73_284 ();
 sg13g2_decap_8 FILLER_73_291 ();
 sg13g2_decap_8 FILLER_73_298 ();
 sg13g2_decap_8 FILLER_73_313 ();
 sg13g2_decap_8 FILLER_73_320 ();
 sg13g2_decap_4 FILLER_73_327 ();
 sg13g2_decap_8 FILLER_73_335 ();
 sg13g2_fill_2 FILLER_73_342 ();
 sg13g2_fill_1 FILLER_73_344 ();
 sg13g2_decap_8 FILLER_73_349 ();
 sg13g2_decap_8 FILLER_73_356 ();
 sg13g2_fill_1 FILLER_73_363 ();
 sg13g2_fill_2 FILLER_73_374 ();
 sg13g2_fill_1 FILLER_73_376 ();
 sg13g2_fill_1 FILLER_73_381 ();
 sg13g2_fill_1 FILLER_73_394 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_73_421 ();
 sg13g2_fill_2 FILLER_73_428 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_4 FILLER_74_42 ();
 sg13g2_fill_1 FILLER_74_108 ();
 sg13g2_decap_8 FILLER_74_121 ();
 sg13g2_fill_1 FILLER_74_128 ();
 sg13g2_fill_1 FILLER_74_163 ();
 sg13g2_decap_8 FILLER_74_190 ();
 sg13g2_fill_2 FILLER_74_197 ();
 sg13g2_fill_1 FILLER_74_213 ();
 sg13g2_decap_4 FILLER_74_226 ();
 sg13g2_fill_2 FILLER_74_230 ();
 sg13g2_fill_2 FILLER_74_238 ();
 sg13g2_decap_4 FILLER_74_257 ();
 sg13g2_fill_2 FILLER_74_276 ();
 sg13g2_decap_8 FILLER_74_283 ();
 sg13g2_fill_1 FILLER_74_290 ();
 sg13g2_decap_4 FILLER_74_323 ();
 sg13g2_fill_2 FILLER_74_327 ();
 sg13g2_decap_8 FILLER_74_334 ();
 sg13g2_decap_4 FILLER_74_341 ();
 sg13g2_fill_2 FILLER_74_345 ();
 sg13g2_fill_1 FILLER_74_356 ();
 sg13g2_fill_2 FILLER_74_362 ();
 sg13g2_decap_4 FILLER_74_376 ();
 sg13g2_fill_2 FILLER_74_391 ();
 sg13g2_fill_1 FILLER_74_398 ();
 sg13g2_fill_1 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_74_412 ();
 sg13g2_decap_8 FILLER_74_419 ();
 sg13g2_decap_4 FILLER_74_426 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_4 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_44 ();
 sg13g2_decap_8 FILLER_75_51 ();
 sg13g2_decap_8 FILLER_75_58 ();
 sg13g2_decap_8 FILLER_75_65 ();
 sg13g2_decap_8 FILLER_75_72 ();
 sg13g2_decap_8 FILLER_75_79 ();
 sg13g2_decap_4 FILLER_75_94 ();
 sg13g2_fill_2 FILLER_75_98 ();
 sg13g2_fill_1 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_164 ();
 sg13g2_decap_4 FILLER_75_171 ();
 sg13g2_fill_1 FILLER_75_175 ();
 sg13g2_fill_1 FILLER_75_199 ();
 sg13g2_fill_1 FILLER_75_216 ();
 sg13g2_fill_1 FILLER_75_222 ();
 sg13g2_fill_1 FILLER_75_231 ();
 sg13g2_fill_1 FILLER_75_237 ();
 sg13g2_fill_1 FILLER_75_243 ();
 sg13g2_fill_2 FILLER_75_280 ();
 sg13g2_fill_1 FILLER_75_290 ();
 sg13g2_fill_2 FILLER_75_307 ();
 sg13g2_fill_1 FILLER_75_309 ();
 sg13g2_fill_2 FILLER_75_321 ();
 sg13g2_fill_1 FILLER_75_334 ();
 sg13g2_decap_4 FILLER_75_339 ();
 sg13g2_fill_1 FILLER_75_350 ();
 sg13g2_fill_1 FILLER_75_355 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_fill_1 FILLER_75_366 ();
 sg13g2_fill_1 FILLER_75_372 ();
 sg13g2_fill_2 FILLER_75_379 ();
 sg13g2_decap_4 FILLER_75_397 ();
 sg13g2_fill_1 FILLER_75_401 ();
 sg13g2_decap_8 FILLER_75_422 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_4 FILLER_76_21 ();
 sg13g2_fill_1 FILLER_76_25 ();
 sg13g2_fill_2 FILLER_76_32 ();
 sg13g2_decap_4 FILLER_76_48 ();
 sg13g2_fill_2 FILLER_76_52 ();
 sg13g2_decap_8 FILLER_76_62 ();
 sg13g2_decap_8 FILLER_76_69 ();
 sg13g2_fill_2 FILLER_76_76 ();
 sg13g2_fill_1 FILLER_76_78 ();
 sg13g2_fill_1 FILLER_76_92 ();
 sg13g2_fill_2 FILLER_76_104 ();
 sg13g2_fill_2 FILLER_76_127 ();
 sg13g2_decap_8 FILLER_76_137 ();
 sg13g2_decap_8 FILLER_76_144 ();
 sg13g2_decap_8 FILLER_76_151 ();
 sg13g2_fill_2 FILLER_76_158 ();
 sg13g2_fill_1 FILLER_76_160 ();
 sg13g2_decap_8 FILLER_76_176 ();
 sg13g2_fill_2 FILLER_76_183 ();
 sg13g2_fill_1 FILLER_76_185 ();
 sg13g2_decap_4 FILLER_76_192 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_fill_1 FILLER_76_217 ();
 sg13g2_fill_2 FILLER_76_229 ();
 sg13g2_fill_1 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_237 ();
 sg13g2_decap_8 FILLER_76_249 ();
 sg13g2_decap_8 FILLER_76_256 ();
 sg13g2_decap_4 FILLER_76_263 ();
 sg13g2_fill_2 FILLER_76_267 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_4 FILLER_76_280 ();
 sg13g2_fill_2 FILLER_76_317 ();
 sg13g2_fill_1 FILLER_76_319 ();
 sg13g2_fill_1 FILLER_76_326 ();
 sg13g2_decap_4 FILLER_76_331 ();
 sg13g2_fill_1 FILLER_76_352 ();
 sg13g2_decap_4 FILLER_76_370 ();
 sg13g2_fill_1 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_383 ();
 sg13g2_decap_8 FILLER_76_395 ();
 sg13g2_decap_4 FILLER_76_402 ();
 sg13g2_fill_1 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_decap_4 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_30 ();
 sg13g2_decap_8 FILLER_77_44 ();
 sg13g2_decap_4 FILLER_77_51 ();
 sg13g2_fill_2 FILLER_77_55 ();
 sg13g2_decap_8 FILLER_77_83 ();
 sg13g2_decap_8 FILLER_77_90 ();
 sg13g2_decap_4 FILLER_77_97 ();
 sg13g2_decap_8 FILLER_77_136 ();
 sg13g2_decap_8 FILLER_77_143 ();
 sg13g2_decap_8 FILLER_77_150 ();
 sg13g2_decap_8 FILLER_77_157 ();
 sg13g2_fill_1 FILLER_77_208 ();
 sg13g2_decap_4 FILLER_77_213 ();
 sg13g2_fill_1 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_248 ();
 sg13g2_decap_4 FILLER_77_255 ();
 sg13g2_decap_8 FILLER_77_263 ();
 sg13g2_fill_1 FILLER_77_274 ();
 sg13g2_fill_2 FILLER_77_280 ();
 sg13g2_fill_2 FILLER_77_287 ();
 sg13g2_fill_2 FILLER_77_293 ();
 sg13g2_fill_1 FILLER_77_303 ();
 sg13g2_fill_1 FILLER_77_309 ();
 sg13g2_fill_1 FILLER_77_316 ();
 sg13g2_fill_2 FILLER_77_327 ();
 sg13g2_fill_1 FILLER_77_329 ();
 sg13g2_fill_2 FILLER_77_340 ();
 sg13g2_fill_1 FILLER_77_342 ();
 sg13g2_fill_2 FILLER_77_347 ();
 sg13g2_fill_1 FILLER_77_369 ();
 sg13g2_fill_2 FILLER_77_375 ();
 sg13g2_fill_1 FILLER_77_382 ();
 sg13g2_fill_2 FILLER_77_393 ();
 sg13g2_decap_4 FILLER_77_425 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_4 FILLER_78_7 ();
 sg13g2_fill_2 FILLER_78_11 ();
 sg13g2_decap_4 FILLER_78_51 ();
 sg13g2_fill_1 FILLER_78_55 ();
 sg13g2_decap_8 FILLER_78_109 ();
 sg13g2_decap_4 FILLER_78_116 ();
 sg13g2_fill_1 FILLER_78_120 ();
 sg13g2_fill_2 FILLER_78_127 ();
 sg13g2_decap_8 FILLER_78_152 ();
 sg13g2_fill_2 FILLER_78_159 ();
 sg13g2_fill_1 FILLER_78_161 ();
 sg13g2_fill_1 FILLER_78_226 ();
 sg13g2_decap_4 FILLER_78_247 ();
 sg13g2_fill_2 FILLER_78_266 ();
 sg13g2_decap_4 FILLER_78_275 ();
 sg13g2_fill_2 FILLER_78_279 ();
 sg13g2_fill_2 FILLER_78_301 ();
 sg13g2_fill_1 FILLER_78_303 ();
 sg13g2_fill_2 FILLER_78_313 ();
 sg13g2_fill_1 FILLER_78_358 ();
 sg13g2_fill_1 FILLER_78_369 ();
 sg13g2_fill_2 FILLER_78_382 ();
 sg13g2_fill_2 FILLER_78_396 ();
 sg13g2_fill_2 FILLER_78_427 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_4 FILLER_79_21 ();
 sg13g2_fill_2 FILLER_79_25 ();
 sg13g2_decap_4 FILLER_79_30 ();
 sg13g2_fill_1 FILLER_79_34 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_fill_1 FILLER_79_77 ();
 sg13g2_decap_4 FILLER_79_116 ();
 sg13g2_decap_4 FILLER_79_178 ();
 sg13g2_decap_4 FILLER_79_191 ();
 sg13g2_fill_2 FILLER_79_195 ();
 sg13g2_fill_1 FILLER_79_200 ();
 sg13g2_decap_4 FILLER_79_205 ();
 sg13g2_fill_2 FILLER_79_209 ();
 sg13g2_decap_8 FILLER_79_215 ();
 sg13g2_decap_8 FILLER_79_232 ();
 sg13g2_decap_8 FILLER_79_239 ();
 sg13g2_fill_1 FILLER_79_256 ();
 sg13g2_decap_8 FILLER_79_267 ();
 sg13g2_fill_1 FILLER_79_274 ();
 sg13g2_fill_2 FILLER_79_280 ();
 sg13g2_fill_2 FILLER_79_287 ();
 sg13g2_fill_2 FILLER_79_316 ();
 sg13g2_fill_1 FILLER_79_318 ();
 sg13g2_fill_2 FILLER_79_323 ();
 sg13g2_decap_4 FILLER_79_335 ();
 sg13g2_fill_1 FILLER_79_339 ();
 sg13g2_decap_8 FILLER_79_344 ();
 sg13g2_fill_2 FILLER_79_351 ();
 sg13g2_fill_2 FILLER_79_358 ();
 sg13g2_decap_8 FILLER_79_365 ();
 sg13g2_decap_4 FILLER_79_372 ();
 sg13g2_decap_4 FILLER_79_393 ();
 sg13g2_fill_2 FILLER_79_397 ();
 sg13g2_fill_1 FILLER_79_404 ();
 sg13g2_fill_1 FILLER_79_416 ();
 sg13g2_decap_8 FILLER_79_422 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_4 FILLER_80_28 ();
 sg13g2_fill_2 FILLER_80_32 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_77 ();
 sg13g2_decap_4 FILLER_80_86 ();
 sg13g2_fill_2 FILLER_80_90 ();
 sg13g2_fill_2 FILLER_80_100 ();
 sg13g2_fill_1 FILLER_80_102 ();
 sg13g2_fill_2 FILLER_80_107 ();
 sg13g2_fill_1 FILLER_80_109 ();
 sg13g2_fill_1 FILLER_80_118 ();
 sg13g2_fill_2 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_125 ();
 sg13g2_fill_2 FILLER_80_134 ();
 sg13g2_fill_1 FILLER_80_140 ();
 sg13g2_fill_1 FILLER_80_149 ();
 sg13g2_fill_2 FILLER_80_154 ();
 sg13g2_fill_1 FILLER_80_156 ();
 sg13g2_fill_2 FILLER_80_165 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_fill_2 FILLER_80_184 ();
 sg13g2_fill_1 FILLER_80_186 ();
 sg13g2_fill_1 FILLER_80_191 ();
 sg13g2_fill_1 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_201 ();
 sg13g2_decap_4 FILLER_80_209 ();
 sg13g2_decap_4 FILLER_80_221 ();
 sg13g2_fill_2 FILLER_80_225 ();
 sg13g2_decap_8 FILLER_80_235 ();
 sg13g2_fill_1 FILLER_80_242 ();
 sg13g2_decap_4 FILLER_80_247 ();
 sg13g2_decap_8 FILLER_80_269 ();
 sg13g2_decap_8 FILLER_80_276 ();
 sg13g2_fill_2 FILLER_80_283 ();
 sg13g2_decap_8 FILLER_80_290 ();
 sg13g2_decap_8 FILLER_80_297 ();
 sg13g2_decap_8 FILLER_80_304 ();
 sg13g2_decap_8 FILLER_80_311 ();
 sg13g2_decap_4 FILLER_80_318 ();
 sg13g2_decap_8 FILLER_80_333 ();
 sg13g2_fill_1 FILLER_80_340 ();
 sg13g2_decap_8 FILLER_80_345 ();
 sg13g2_fill_2 FILLER_80_352 ();
 sg13g2_fill_1 FILLER_80_354 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_decap_4 FILLER_80_378 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_decap_8 FILLER_80_407 ();
 sg13g2_decap_8 FILLER_80_414 ();
 sg13g2_decap_8 FILLER_80_421 ();
 sg13g2_fill_2 FILLER_80_428 ();
endmodule
