module tt_um_phansel_laplace_lut (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire clknet_0_clk;
 wire net243;
 wire \chars_remaining[0] ;
 wire \chars_remaining[1] ;
 wire \chars_remaining[2] ;
 wire \chars_remaining[3] ;
 wire \chars_remaining[4] ;
 wire \chars_remaining[5] ;
 wire \chars_remaining[6] ;
 wire \chars_remaining[7] ;
 wire \chars_remaining[8] ;
 wire \chars_remaining[9] ;
 wire clk_buffered;
 wire \clk_picker.clk_slow ;
 wire \clk_picker.counter[0] ;
 wire \clk_picker.counter[10] ;
 wire \clk_picker.counter[11] ;
 wire \clk_picker.counter[12] ;
 wire \clk_picker.counter[13] ;
 wire \clk_picker.counter[14] ;
 wire \clk_picker.counter[15] ;
 wire \clk_picker.counter[16] ;
 wire \clk_picker.counter[17] ;
 wire \clk_picker.counter[18] ;
 wire \clk_picker.counter[19] ;
 wire \clk_picker.counter[1] ;
 wire \clk_picker.counter[20] ;
 wire \clk_picker.counter[21] ;
 wire \clk_picker.counter[22] ;
 wire \clk_picker.counter[23] ;
 wire \clk_picker.counter[24] ;
 wire \clk_picker.counter[25] ;
 wire \clk_picker.counter[2] ;
 wire \clk_picker.counter[3] ;
 wire \clk_picker.counter[4] ;
 wire \clk_picker.counter[5] ;
 wire \clk_picker.counter[6] ;
 wire \clk_picker.counter[7] ;
 wire \clk_picker.counter[8] ;
 wire \clk_picker.counter[9] ;
 wire \line_mapper_1.pointer_addr[0] ;
 wire \line_mapper_1.pointer_addr[10] ;
 wire \line_mapper_1.pointer_addr[11] ;
 wire \line_mapper_1.pointer_addr[12] ;
 wire \line_mapper_1.pointer_addr[13] ;
 wire \line_mapper_1.pointer_addr[14] ;
 wire \line_mapper_1.pointer_addr[15] ;
 wire \line_mapper_1.pointer_addr[1] ;
 wire \line_mapper_1.pointer_addr[2] ;
 wire \line_mapper_1.pointer_addr[3] ;
 wire \line_mapper_1.pointer_addr[4] ;
 wire \line_mapper_1.pointer_addr[5] ;
 wire \line_mapper_1.pointer_addr[6] ;
 wire \line_mapper_1.pointer_addr[7] ;
 wire \line_mapper_1.pointer_addr[8] ;
 wire \line_mapper_1.pointer_addr[9] ;
 wire \mem_addr[0] ;
 wire \mem_addr[1] ;
 wire \mem_addr[2] ;
 wire \mem_addr[3] ;
 wire \mem_addr[4] ;
 wire \mem_addr[5] ;
 wire \mem_addr[6] ;
 wire \mem_addr[7] ;
 wire \mem_addr[8] ;
 wire \memory_1.mem_addr[9] ;
 wire \transformer_1.started ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_0_clk_buffered;
 wire clknet_3_0__leaf_clk_buffered;
 wire clknet_3_1__leaf_clk_buffered;
 wire clknet_3_2__leaf_clk_buffered;
 wire clknet_3_3__leaf_clk_buffered;
 wire clknet_3_4__leaf_clk_buffered;
 wire clknet_3_5__leaf_clk_buffered;
 wire clknet_3_6__leaf_clk_buffered;
 wire clknet_3_7__leaf_clk_buffered;

 sg13g2_buf_1 _3126_ (.A(\mem_addr[0] ),
    .X(_0725_));
 sg13g2_buf_1 _3127_ (.A(\mem_addr[1] ),
    .X(_0736_));
 sg13g2_nand2_1 _3128_ (.Y(_0747_),
    .A(net229),
    .B(net228));
 sg13g2_buf_2 _3129_ (.A(_0747_),
    .X(_0758_));
 sg13g2_buf_8 _3130_ (.A(\mem_addr[2] ),
    .X(_0769_));
 sg13g2_inv_2 _3131_ (.Y(_0780_),
    .A(_0769_));
 sg13g2_buf_8 _3132_ (.A(\mem_addr[3] ),
    .X(_0791_));
 sg13g2_inv_2 _3133_ (.Y(_0802_),
    .A(_0791_));
 sg13g2_nand3_1 _3134_ (.B(_0780_),
    .C(_0802_),
    .A(_0758_),
    .Y(_0813_));
 sg13g2_inv_4 _3135_ (.A(net229),
    .Y(_0823_));
 sg13g2_inv_4 _3136_ (.A(net228),
    .Y(_0834_));
 sg13g2_nand2_2 _3137_ (.Y(_0845_),
    .A(_0823_),
    .B(_0834_));
 sg13g2_nor2b_1 _3138_ (.A(_0813_),
    .B_N(_0845_),
    .Y(_0856_));
 sg13g2_buf_2 _3139_ (.A(_0856_),
    .X(_0867_));
 sg13g2_buf_8 _3140_ (.A(_0791_),
    .X(_0878_));
 sg13g2_nand2_1 _3141_ (.Y(_0889_),
    .A(net228),
    .B(_0769_));
 sg13g2_buf_2 _3142_ (.A(_0889_),
    .X(_0900_));
 sg13g2_nor2_2 _3143_ (.A(_0878_),
    .B(_0900_),
    .Y(_0911_));
 sg13g2_inv_1 _3144_ (.Y(_0922_),
    .A(_0911_));
 sg13g2_nor2b_1 _3145_ (.A(_0867_),
    .B_N(_0922_),
    .Y(_0933_));
 sg13g2_buf_2 _3146_ (.A(_0933_),
    .X(_0944_));
 sg13g2_buf_8 _3147_ (.A(net228),
    .X(_0955_));
 sg13g2_buf_8 _3148_ (.A(_0823_),
    .X(_0966_));
 sg13g2_nor2_2 _3149_ (.A(_0955_),
    .B(net210),
    .Y(_0976_));
 sg13g2_buf_8 _3150_ (.A(_0769_),
    .X(_0987_));
 sg13g2_buf_8 _3151_ (.A(net223),
    .X(_0998_));
 sg13g2_nand2_1 _3152_ (.Y(_1009_),
    .A(_0976_),
    .B(net209));
 sg13g2_buf_1 _3153_ (.A(_1009_),
    .X(_1020_));
 sg13g2_buf_8 _3154_ (.A(_0834_),
    .X(_1031_));
 sg13g2_nor2_2 _3155_ (.A(net223),
    .B(net208),
    .Y(_1042_));
 sg13g2_nand2_1 _3156_ (.Y(_1053_),
    .A(_1042_),
    .B(net210));
 sg13g2_buf_1 _3157_ (.A(_1053_),
    .X(_1064_));
 sg13g2_nand2_1 _3158_ (.Y(_1075_),
    .A(net83),
    .B(net82));
 sg13g2_buf_1 _3159_ (.A(net225),
    .X(_1086_));
 sg13g2_buf_8 _3160_ (.A(net207),
    .X(_1097_));
 sg13g2_buf_8 _3161_ (.A(net180),
    .X(_1108_));
 sg13g2_nand2_2 _3162_ (.Y(_1119_),
    .A(_1075_),
    .B(net132));
 sg13g2_buf_2 _3163_ (.A(\mem_addr[4] ),
    .X(_1130_));
 sg13g2_buf_1 _3164_ (.A(\mem_addr[5] ),
    .X(_1140_));
 sg13g2_nand2_1 _3165_ (.Y(_1151_),
    .A(_1130_),
    .B(net227));
 sg13g2_buf_2 _3166_ (.A(_1151_),
    .X(_1162_));
 sg13g2_buf_1 _3167_ (.A(_1162_),
    .X(_1173_));
 sg13g2_a21oi_1 _3168_ (.A1(_0944_),
    .A2(_1119_),
    .Y(_1184_),
    .B1(net179));
 sg13g2_nor2_1 _3169_ (.A(net229),
    .B(net228),
    .Y(_1195_));
 sg13g2_buf_2 _3170_ (.A(_1195_),
    .X(_1206_));
 sg13g2_nand2_1 _3171_ (.Y(_1217_),
    .A(_1206_),
    .B(net223));
 sg13g2_buf_1 _3172_ (.A(_1217_),
    .X(_1228_));
 sg13g2_buf_8 _3173_ (.A(net229),
    .X(_1239_));
 sg13g2_nand3_1 _3174_ (.B(net224),
    .C(_0987_),
    .A(net222),
    .Y(_1250_));
 sg13g2_buf_2 _3175_ (.A(_1250_),
    .X(_1261_));
 sg13g2_nand2_1 _3176_ (.Y(_1272_),
    .A(_0780_),
    .B(net229));
 sg13g2_buf_4 _3177_ (.X(_1283_),
    .A(_1272_));
 sg13g2_nand3_1 _3178_ (.B(_1261_),
    .C(_1283_),
    .A(net131),
    .Y(_1293_));
 sg13g2_buf_1 _3179_ (.A(net180),
    .X(_1304_));
 sg13g2_nand2_1 _3180_ (.Y(_1315_),
    .A(_1293_),
    .B(net130));
 sg13g2_nand2_1 _3181_ (.Y(_1326_),
    .A(_0802_),
    .B(net224));
 sg13g2_buf_2 _3182_ (.A(_1326_),
    .X(_1337_));
 sg13g2_buf_1 _3183_ (.A(_1337_),
    .X(_1348_));
 sg13g2_nand2_1 _3184_ (.Y(_1359_),
    .A(net210),
    .B(net223));
 sg13g2_buf_2 _3185_ (.A(_1359_),
    .X(_1370_));
 sg13g2_buf_8 _3186_ (.A(_1370_),
    .X(_1381_));
 sg13g2_inv_1 _3187_ (.Y(_1392_),
    .A(_1381_));
 sg13g2_nor2_1 _3188_ (.A(_1348_),
    .B(_1392_),
    .Y(_1403_));
 sg13g2_inv_2 _3189_ (.Y(_1413_),
    .A(_1403_));
 sg13g2_nor2_1 _3190_ (.A(_1130_),
    .B(net227),
    .Y(_1424_));
 sg13g2_buf_2 _3191_ (.A(_1424_),
    .X(_1435_));
 sg13g2_inv_1 _3192_ (.Y(_1446_),
    .A(_1435_));
 sg13g2_buf_1 _3193_ (.A(_1446_),
    .X(_1457_));
 sg13g2_buf_1 _3194_ (.A(net128),
    .X(_1468_));
 sg13g2_a21oi_1 _3195_ (.A1(_1315_),
    .A2(_1413_),
    .Y(_1479_),
    .B1(net80));
 sg13g2_nor2_1 _3196_ (.A(_1184_),
    .B(_1479_),
    .Y(_1490_));
 sg13g2_nand2_1 _3197_ (.Y(_1501_),
    .A(_0845_),
    .B(_0758_));
 sg13g2_buf_2 _3198_ (.A(_1501_),
    .X(_1512_));
 sg13g2_buf_8 _3199_ (.A(_1512_),
    .X(_1523_));
 sg13g2_buf_1 _3200_ (.A(_0780_),
    .X(_1534_));
 sg13g2_nand3_1 _3201_ (.B(net206),
    .C(net180),
    .A(net79),
    .Y(_1544_));
 sg13g2_buf_1 _3202_ (.A(_1544_),
    .X(_1555_));
 sg13g2_nand2_1 _3203_ (.Y(_1566_),
    .A(_0834_),
    .B(net229));
 sg13g2_buf_2 _3204_ (.A(_1566_),
    .X(_1577_));
 sg13g2_nand2_1 _3205_ (.Y(_1588_),
    .A(_0823_),
    .B(net228));
 sg13g2_buf_1 _3206_ (.A(_1588_),
    .X(_1599_));
 sg13g2_nand2_1 _3207_ (.Y(_1610_),
    .A(_1577_),
    .B(net178));
 sg13g2_buf_8 _3208_ (.A(_1610_),
    .X(_1621_));
 sg13g2_nor2_1 _3209_ (.A(net229),
    .B(_0769_),
    .Y(_1632_));
 sg13g2_buf_2 _3210_ (.A(_1632_),
    .X(_1643_));
 sg13g2_buf_1 _3211_ (.A(_1643_),
    .X(_1654_));
 sg13g2_nor2_1 _3212_ (.A(_1086_),
    .B(_1654_),
    .Y(_1664_));
 sg13g2_buf_2 _3213_ (.A(_1664_),
    .X(_1675_));
 sg13g2_nand2_1 _3214_ (.Y(_1686_),
    .A(net78),
    .B(_1675_));
 sg13g2_buf_8 _3215_ (.A(_0802_),
    .X(_1697_));
 sg13g2_buf_8 _3216_ (.A(net205),
    .X(_1708_));
 sg13g2_buf_1 _3217_ (.A(_0900_),
    .X(_1719_));
 sg13g2_nor2_2 _3218_ (.A(net176),
    .B(net175),
    .Y(_1730_));
 sg13g2_inv_2 _3219_ (.Y(_1741_),
    .A(_1730_));
 sg13g2_nand3_1 _3220_ (.B(_1686_),
    .C(_1741_),
    .A(_1555_),
    .Y(_1752_));
 sg13g2_inv_4 _3221_ (.A(_1130_),
    .Y(_1763_));
 sg13g2_nor2_1 _3222_ (.A(net227),
    .B(_1763_),
    .Y(_1774_));
 sg13g2_buf_2 _3223_ (.A(_1774_),
    .X(_1785_));
 sg13g2_buf_1 _3224_ (.A(_1785_),
    .X(_1796_));
 sg13g2_nand2_1 _3225_ (.Y(_1806_),
    .A(net228),
    .B(_0791_));
 sg13g2_buf_1 _3226_ (.A(_1806_),
    .X(_1817_));
 sg13g2_nand2_2 _3227_ (.Y(_1828_),
    .A(_0769_),
    .B(_0791_));
 sg13g2_nand2_1 _3228_ (.Y(_1839_),
    .A(net204),
    .B(_1828_));
 sg13g2_buf_8 _3229_ (.A(_1283_),
    .X(_1850_));
 sg13g2_nand3_1 _3230_ (.B(_1577_),
    .C(net126),
    .A(_1839_),
    .Y(_1861_));
 sg13g2_nand2_1 _3231_ (.Y(_1872_),
    .A(_1763_),
    .B(net227));
 sg13g2_nor2_2 _3232_ (.A(net207),
    .B(_1370_),
    .Y(_1882_));
 sg13g2_nor2_1 _3233_ (.A(_1872_),
    .B(_1882_),
    .Y(_1893_));
 sg13g2_nand2_1 _3234_ (.Y(_1904_),
    .A(_1861_),
    .B(_1893_));
 sg13g2_nor2_1 _3235_ (.A(_0867_),
    .B(_1904_),
    .Y(_1915_));
 sg13g2_a21oi_1 _3236_ (.A1(_1752_),
    .A2(net127),
    .Y(_1926_),
    .B1(_1915_));
 sg13g2_nand2_1 _3237_ (.Y(_1937_),
    .A(_1490_),
    .B(_1926_));
 sg13g2_buf_2 _3238_ (.A(\mem_addr[6] ),
    .X(_1948_));
 sg13g2_inv_1 _3239_ (.Y(_1959_),
    .A(_1948_));
 sg13g2_buf_1 _3240_ (.A(_1959_),
    .X(_1970_));
 sg13g2_buf_2 _3241_ (.A(net203),
    .X(_1981_));
 sg13g2_buf_1 _3242_ (.A(net174),
    .X(_1991_));
 sg13g2_nand2_1 _3243_ (.Y(_2002_),
    .A(_1937_),
    .B(net125));
 sg13g2_nand2_1 _3244_ (.Y(_2013_),
    .A(net222),
    .B(net223));
 sg13g2_buf_1 _3245_ (.A(_2013_),
    .X(_2024_));
 sg13g2_inv_1 _3246_ (.Y(_2035_),
    .A(net173));
 sg13g2_nand2_1 _3247_ (.Y(_2045_),
    .A(_1643_),
    .B(net208));
 sg13g2_buf_1 _3248_ (.A(_2045_),
    .X(_2056_));
 sg13g2_buf_8 _3249_ (.A(net176),
    .X(_2066_));
 sg13g2_nand2_2 _3250_ (.Y(_2077_),
    .A(_2056_),
    .B(net123));
 sg13g2_nor2_1 _3251_ (.A(_2035_),
    .B(_2077_),
    .Y(_2087_));
 sg13g2_nor2_2 _3252_ (.A(net222),
    .B(net208),
    .Y(_2097_));
 sg13g2_nor2_1 _3253_ (.A(_0769_),
    .B(_0966_),
    .Y(_2107_));
 sg13g2_buf_2 _3254_ (.A(_2107_),
    .X(_2117_));
 sg13g2_nand2_1 _3255_ (.Y(_2127_),
    .A(_2117_),
    .B(net208));
 sg13g2_buf_2 _3256_ (.A(_2127_),
    .X(_2137_));
 sg13g2_nand2_1 _3257_ (.Y(_2145_),
    .A(_2137_),
    .B(_1108_));
 sg13g2_nor2_1 _3258_ (.A(_2097_),
    .B(_2145_),
    .Y(_2155_));
 sg13g2_buf_1 _3259_ (.A(_1763_),
    .X(_2165_));
 sg13g2_buf_1 _3260_ (.A(net202),
    .X(_2175_));
 sg13g2_buf_1 _3261_ (.A(net172),
    .X(_2184_));
 sg13g2_o21ai_1 _3262_ (.B1(net122),
    .Y(_2195_),
    .A1(_2087_),
    .A2(_2155_));
 sg13g2_nand2_2 _3263_ (.Y(_2206_),
    .A(net173),
    .B(net224));
 sg13g2_inv_2 _3264_ (.Y(_2215_),
    .A(_1643_));
 sg13g2_buf_1 _3265_ (.A(_2215_),
    .X(_2225_));
 sg13g2_nand2_1 _3266_ (.Y(_2234_),
    .A(_2206_),
    .B(_2225_));
 sg13g2_nand2_1 _3267_ (.Y(_2242_),
    .A(net205),
    .B(_1130_));
 sg13g2_buf_2 _3268_ (.A(_2242_),
    .X(_2250_));
 sg13g2_inv_2 _3269_ (.Y(_2259_),
    .A(_2250_));
 sg13g2_nand2_2 _3270_ (.Y(_2267_),
    .A(net225),
    .B(_1130_));
 sg13g2_inv_1 _3271_ (.Y(_2273_),
    .A(_2267_));
 sg13g2_buf_1 _3272_ (.A(_2273_),
    .X(_2280_));
 sg13g2_nand2_1 _3273_ (.Y(_2289_),
    .A(net178),
    .B(_1534_));
 sg13g2_buf_2 _3274_ (.A(_0032_),
    .X(_2300_));
 sg13g2_nand2_1 _3275_ (.Y(_2309_),
    .A(_2300_),
    .B(net223));
 sg13g2_buf_2 _3276_ (.A(_2309_),
    .X(_2318_));
 sg13g2_nand2_1 _3277_ (.Y(_2327_),
    .A(_2289_),
    .B(_2318_));
 sg13g2_a22oi_1 _3278_ (.Y(_2335_),
    .B1(net120),
    .B2(_2327_),
    .A2(_2259_),
    .A1(_2234_));
 sg13g2_nand2_1 _3279_ (.Y(_2343_),
    .A(_2195_),
    .B(_2335_));
 sg13g2_nor2_1 _3280_ (.A(net227),
    .B(_1959_),
    .Y(_2352_));
 sg13g2_buf_1 _3281_ (.A(_2352_),
    .X(_2361_));
 sg13g2_buf_1 _3282_ (.A(net172),
    .X(_2370_));
 sg13g2_buf_1 _3283_ (.A(net119),
    .X(_2378_));
 sg13g2_buf_8 _3284_ (.A(net209),
    .X(_2379_));
 sg13g2_nand2_2 _3285_ (.Y(_2380_),
    .A(net208),
    .B(net225));
 sg13g2_nor2_2 _3286_ (.A(net170),
    .B(_2380_),
    .Y(_2381_));
 sg13g2_nand2_1 _3287_ (.Y(_2382_),
    .A(net229),
    .B(_0791_));
 sg13g2_buf_1 _3288_ (.A(_2382_),
    .X(_2383_));
 sg13g2_inv_2 _3289_ (.Y(_2384_),
    .A(net201));
 sg13g2_nand2_1 _3290_ (.Y(_2385_),
    .A(net208),
    .B(_2300_));
 sg13g2_buf_1 _3291_ (.A(net224),
    .X(_2386_));
 sg13g2_buf_2 _3292_ (.A(_0037_),
    .X(_2387_));
 sg13g2_buf_1 _3293_ (.A(_2387_),
    .X(_2388_));
 sg13g2_nand2_1 _3294_ (.Y(_2389_),
    .A(net200),
    .B(net221));
 sg13g2_buf_1 _3295_ (.A(_1086_),
    .X(_2390_));
 sg13g2_buf_1 _3296_ (.A(net169),
    .X(_2391_));
 sg13g2_a21oi_1 _3297_ (.A1(_2385_),
    .A2(_2389_),
    .Y(_2392_),
    .B1(_2391_));
 sg13g2_nor3_1 _3298_ (.A(_2381_),
    .B(_2384_),
    .C(_2392_),
    .Y(_2393_));
 sg13g2_nor2_1 _3299_ (.A(_0736_),
    .B(_0802_),
    .Y(_2394_));
 sg13g2_buf_1 _3300_ (.A(_2394_),
    .X(_2395_));
 sg13g2_nand2_1 _3301_ (.Y(_2396_),
    .A(net168),
    .B(_1643_));
 sg13g2_buf_2 _3302_ (.A(_2396_),
    .X(_2397_));
 sg13g2_buf_2 _3303_ (.A(_1130_),
    .X(_2398_));
 sg13g2_nand2_2 _3304_ (.Y(_2399_),
    .A(_2397_),
    .B(net220));
 sg13g2_nand2_1 _3305_ (.Y(_2400_),
    .A(_1283_),
    .B(_1370_));
 sg13g2_inv_2 _3306_ (.Y(_2401_),
    .A(_1337_));
 sg13g2_nand2_1 _3307_ (.Y(_2402_),
    .A(_2400_),
    .B(net117));
 sg13g2_inv_1 _3308_ (.Y(_2403_),
    .A(_2402_));
 sg13g2_nand2_1 _3309_ (.Y(_2404_),
    .A(net227),
    .B(_1948_));
 sg13g2_buf_2 _3310_ (.A(_2404_),
    .X(_2405_));
 sg13g2_inv_1 _3311_ (.Y(_2406_),
    .A(_2405_));
 sg13g2_o21ai_1 _3312_ (.B1(net167),
    .Y(_2407_),
    .A1(_2399_),
    .A2(_2403_));
 sg13g2_a21oi_1 _3313_ (.A1(net76),
    .A2(_2393_),
    .Y(_2408_),
    .B1(_2407_));
 sg13g2_a21oi_1 _3314_ (.A1(_2343_),
    .A2(net171),
    .Y(_2409_),
    .B1(_2408_));
 sg13g2_nand2_1 _3315_ (.Y(_2410_),
    .A(_2002_),
    .B(_2409_));
 sg13g2_buf_1 _3316_ (.A(\mem_addr[7] ),
    .X(_2411_));
 sg13g2_inv_2 _3317_ (.Y(_2412_),
    .A(_2411_));
 sg13g2_buf_1 _3318_ (.A(_2412_),
    .X(_2413_));
 sg13g2_buf_1 _3319_ (.A(net199),
    .X(_2414_));
 sg13g2_nand2_1 _3320_ (.Y(_2415_),
    .A(_2410_),
    .B(net166));
 sg13g2_nand2_1 _3321_ (.Y(_2416_),
    .A(_1948_),
    .B(_2411_));
 sg13g2_buf_2 _3322_ (.A(_2416_),
    .X(_2417_));
 sg13g2_buf_1 _3323_ (.A(_2417_),
    .X(_2418_));
 sg13g2_inv_1 _3324_ (.Y(_2419_),
    .A(net227));
 sg13g2_buf_1 _3325_ (.A(_2419_),
    .X(_2420_));
 sg13g2_buf_1 _3326_ (.A(net198),
    .X(_2421_));
 sg13g2_buf_1 _3327_ (.A(net164),
    .X(_2422_));
 sg13g2_buf_1 _3328_ (.A(_2422_),
    .X(_2423_));
 sg13g2_buf_1 _3329_ (.A(_2400_),
    .X(_2424_));
 sg13g2_buf_8 _3330_ (.A(net123),
    .X(_2425_));
 sg13g2_buf_1 _3331_ (.A(net74),
    .X(_2426_));
 sg13g2_nand2_1 _3332_ (.Y(_2427_),
    .A(net46),
    .B(net45));
 sg13g2_nand2_1 _3333_ (.Y(_2428_),
    .A(_0834_),
    .B(_0769_));
 sg13g2_buf_2 _3334_ (.A(_2428_),
    .X(_2429_));
 sg13g2_buf_1 _3335_ (.A(net220),
    .X(_2430_));
 sg13g2_buf_2 _3336_ (.A(net197),
    .X(_2431_));
 sg13g2_nand2_1 _3337_ (.Y(_2432_),
    .A(_2429_),
    .B(net163));
 sg13g2_nor2_2 _3338_ (.A(_1239_),
    .B(_2387_),
    .Y(_2433_));
 sg13g2_inv_2 _3339_ (.Y(_2434_),
    .A(_2433_));
 sg13g2_nor2_2 _3340_ (.A(net204),
    .B(_2434_),
    .Y(_2435_));
 sg13g2_nor2_1 _3341_ (.A(net220),
    .B(_2435_),
    .Y(_2436_));
 sg13g2_nor2_1 _3342_ (.A(_2387_),
    .B(net210),
    .Y(_2437_));
 sg13g2_nor2_1 _3343_ (.A(net224),
    .B(_0791_),
    .Y(_2438_));
 sg13g2_buf_4 _3344_ (.X(_2439_),
    .A(_2438_));
 sg13g2_nand2_1 _3345_ (.Y(_2440_),
    .A(_2437_),
    .B(_2439_));
 sg13g2_buf_1 _3346_ (.A(_2440_),
    .X(_2441_));
 sg13g2_nand2_1 _3347_ (.Y(_2442_),
    .A(_2436_),
    .B(net73));
 sg13g2_o21ai_1 _3348_ (.B1(_2442_),
    .Y(_2443_),
    .A1(_2427_),
    .A2(_2432_));
 sg13g2_nand2_1 _3349_ (.Y(_2444_),
    .A(_2384_),
    .B(_2429_));
 sg13g2_nand2_1 _3350_ (.Y(_2445_),
    .A(_1042_),
    .B(net207));
 sg13g2_nand2_1 _3351_ (.Y(_2446_),
    .A(_2444_),
    .B(_2445_));
 sg13g2_inv_2 _3352_ (.Y(_2447_),
    .A(_1872_));
 sg13g2_o21ai_1 _3353_ (.B1(_2447_),
    .Y(_2448_),
    .A1(_2446_),
    .A2(_2403_));
 sg13g2_nor2_1 _3354_ (.A(net169),
    .B(_2429_),
    .Y(_2449_));
 sg13g2_buf_8 _3355_ (.A(net205),
    .X(_2450_));
 sg13g2_inv_1 _3356_ (.Y(_2451_),
    .A(_0038_));
 sg13g2_nand2_1 _3357_ (.Y(_2452_),
    .A(net210),
    .B(_2451_));
 sg13g2_inv_2 _3358_ (.Y(_2453_),
    .A(_2387_));
 sg13g2_nand2_1 _3359_ (.Y(_2454_),
    .A(_2453_),
    .B(_0725_));
 sg13g2_buf_2 _3360_ (.A(_2454_),
    .X(_2455_));
 sg13g2_nand2_1 _3361_ (.Y(_2456_),
    .A(_2452_),
    .B(_2455_));
 sg13g2_nor2_1 _3362_ (.A(net162),
    .B(_2456_),
    .Y(_2457_));
 sg13g2_inv_1 _3363_ (.Y(_2458_),
    .A(_1162_));
 sg13g2_buf_1 _3364_ (.A(_2458_),
    .X(_2459_));
 sg13g2_o21ai_1 _3365_ (.B1(net115),
    .Y(_2460_),
    .A1(_2449_),
    .A2(_2457_));
 sg13g2_nor2_2 _3366_ (.A(_0998_),
    .B(_1206_),
    .Y(_2461_));
 sg13g2_buf_2 _3367_ (.A(net130),
    .X(_2462_));
 sg13g2_buf_1 _3368_ (.A(_1785_),
    .X(_2463_));
 sg13g2_nand3_1 _3369_ (.B(net72),
    .C(net114),
    .A(_2461_),
    .Y(_2464_));
 sg13g2_nand3_1 _3370_ (.B(_2460_),
    .C(_2464_),
    .A(_2448_),
    .Y(_2465_));
 sg13g2_a21oi_1 _3371_ (.A1(net75),
    .A2(_2443_),
    .Y(_2466_),
    .B1(_2465_));
 sg13g2_nor2_1 _3372_ (.A(net165),
    .B(_2466_),
    .Y(_2467_));
 sg13g2_nor2_1 _3373_ (.A(_1948_),
    .B(_2412_),
    .Y(_2468_));
 sg13g2_inv_1 _3374_ (.Y(_2469_),
    .A(_2468_));
 sg13g2_nand2_1 _3375_ (.Y(_2470_),
    .A(net131),
    .B(_1261_));
 sg13g2_nor2_1 _3376_ (.A(_2461_),
    .B(_2470_),
    .Y(_2471_));
 sg13g2_buf_8 _3377_ (.A(_2450_),
    .X(_2472_));
 sg13g2_nand2_1 _3378_ (.Y(_2473_),
    .A(_2471_),
    .B(net113));
 sg13g2_buf_1 _3379_ (.A(net210),
    .X(_2474_));
 sg13g2_nor2_1 _3380_ (.A(_0038_),
    .B(net160),
    .Y(_2475_));
 sg13g2_nor2_1 _3381_ (.A(net177),
    .B(_2475_),
    .Y(_2476_));
 sg13g2_nand2_1 _3382_ (.Y(_2477_),
    .A(_2476_),
    .B(net118));
 sg13g2_buf_1 _3383_ (.A(_1872_),
    .X(_2478_));
 sg13g2_buf_1 _3384_ (.A(net159),
    .X(_2479_));
 sg13g2_a21oi_1 _3385_ (.A1(_2473_),
    .A2(_2477_),
    .Y(_2480_),
    .B1(net112));
 sg13g2_nand2_1 _3386_ (.Y(_2481_),
    .A(_1512_),
    .B(net209));
 sg13g2_buf_2 _3387_ (.A(_2481_),
    .X(_2482_));
 sg13g2_nand2_1 _3388_ (.Y(_2483_),
    .A(_1610_),
    .B(net206));
 sg13g2_buf_1 _3389_ (.A(_2483_),
    .X(_2484_));
 sg13g2_nand2_1 _3390_ (.Y(_2485_),
    .A(_2482_),
    .B(net44));
 sg13g2_buf_2 _3391_ (.A(net118),
    .X(_2486_));
 sg13g2_buf_2 _3392_ (.A(net202),
    .X(_2487_));
 sg13g2_inv_4 _3393_ (.A(_2439_),
    .Y(_2488_));
 sg13g2_nor2_2 _3394_ (.A(_2455_),
    .B(_2488_),
    .Y(_2489_));
 sg13g2_nor2_2 _3395_ (.A(_2487_),
    .B(_2489_),
    .Y(_2490_));
 sg13g2_buf_1 _3396_ (.A(net227),
    .X(_2491_));
 sg13g2_buf_1 _3397_ (.A(net219),
    .X(_2492_));
 sg13g2_nand2_1 _3398_ (.Y(_2493_),
    .A(_2490_),
    .B(net196));
 sg13g2_a21oi_1 _3399_ (.A1(_2485_),
    .A2(net71),
    .Y(_2494_),
    .B1(_2493_));
 sg13g2_nand2_2 _3400_ (.Y(_2495_),
    .A(net178),
    .B(net209));
 sg13g2_nor2_1 _3401_ (.A(net223),
    .B(_2451_),
    .Y(_2496_));
 sg13g2_inv_1 _3402_ (.Y(_2497_),
    .A(_2496_));
 sg13g2_a21oi_2 _3403_ (.B1(net123),
    .Y(_2498_),
    .A2(_2497_),
    .A1(_2495_));
 sg13g2_nand2_2 _3404_ (.Y(_2499_),
    .A(_2498_),
    .B(net83));
 sg13g2_buf_1 _3405_ (.A(net220),
    .X(_2500_));
 sg13g2_buf_1 _3406_ (.A(net195),
    .X(_2501_));
 sg13g2_nor2_2 _3407_ (.A(net225),
    .B(_2387_),
    .Y(_2502_));
 sg13g2_nand2_1 _3408_ (.Y(_2503_),
    .A(net78),
    .B(_2502_));
 sg13g2_inv_1 _3409_ (.Y(_2504_),
    .A(_2503_));
 sg13g2_nor2_1 _3410_ (.A(net157),
    .B(_2504_),
    .Y(_2505_));
 sg13g2_nand2_2 _3411_ (.Y(_2506_),
    .A(_1381_),
    .B(net208));
 sg13g2_nand2_2 _3412_ (.Y(_2507_),
    .A(_2215_),
    .B(net173));
 sg13g2_a21oi_1 _3413_ (.A1(_2507_),
    .A2(_2280_),
    .Y(_2508_),
    .B1(net219));
 sg13g2_o21ai_1 _3414_ (.B1(_2508_),
    .Y(_2509_),
    .A1(_2506_),
    .A2(_2250_));
 sg13g2_a21oi_1 _3415_ (.A1(_2499_),
    .A2(_2505_),
    .Y(_2510_),
    .B1(_2509_));
 sg13g2_nor3_1 _3416_ (.A(_2480_),
    .B(_2494_),
    .C(_2510_),
    .Y(_2511_));
 sg13g2_nor2_1 _3417_ (.A(net161),
    .B(_2511_),
    .Y(_2512_));
 sg13g2_nor2_1 _3418_ (.A(_2467_),
    .B(_2512_),
    .Y(_2513_));
 sg13g2_nand2_1 _3419_ (.Y(_2514_),
    .A(_2415_),
    .B(_2513_));
 sg13g2_buf_1 _3420_ (.A(\mem_addr[8] ),
    .X(_2515_));
 sg13g2_inv_1 _3421_ (.Y(_2516_),
    .A(_2515_));
 sg13g2_buf_1 _3422_ (.A(net218),
    .X(_2517_));
 sg13g2_nand2_1 _3423_ (.Y(_2518_),
    .A(_2514_),
    .B(net194));
 sg13g2_nand2_2 _3424_ (.Y(_2519_),
    .A(net208),
    .B(net206));
 sg13g2_nand2_1 _3425_ (.Y(_2520_),
    .A(_2519_),
    .B(_0900_));
 sg13g2_buf_1 _3426_ (.A(_2520_),
    .X(_2521_));
 sg13g2_nand2_1 _3427_ (.Y(_2522_),
    .A(net70),
    .B(net160));
 sg13g2_buf_1 _3428_ (.A(_2472_),
    .X(_2523_));
 sg13g2_nand2_1 _3429_ (.Y(_2524_),
    .A(_2522_),
    .B(net69));
 sg13g2_inv_2 _3430_ (.Y(_2525_),
    .A(_1785_));
 sg13g2_buf_1 _3431_ (.A(_2525_),
    .X(_2526_));
 sg13g2_buf_1 _3432_ (.A(net68),
    .X(_2527_));
 sg13g2_a21oi_1 _3433_ (.A1(_2499_),
    .A2(_2524_),
    .Y(_2528_),
    .B1(net43));
 sg13g2_buf_1 _3434_ (.A(net128),
    .X(_2529_));
 sg13g2_a21o_1 _3435_ (.A2(_1119_),
    .A1(_0944_),
    .B1(net67),
    .X(_2530_));
 sg13g2_buf_1 _3436_ (.A(_2478_),
    .X(_2531_));
 sg13g2_nand2_1 _3437_ (.Y(_2532_),
    .A(_1577_),
    .B(_1534_));
 sg13g2_buf_2 _3438_ (.A(_2532_),
    .X(_2533_));
 sg13g2_nor2_1 _3439_ (.A(net162),
    .B(_2533_),
    .Y(_2534_));
 sg13g2_nor2_1 _3440_ (.A(net111),
    .B(_2534_),
    .Y(_2535_));
 sg13g2_nand2_1 _3441_ (.Y(_2536_),
    .A(net82),
    .B(net113));
 sg13g2_buf_1 _3442_ (.A(_2459_),
    .X(_2537_));
 sg13g2_nor2_2 _3443_ (.A(net224),
    .B(net206),
    .Y(_2538_));
 sg13g2_nor2_1 _3444_ (.A(net205),
    .B(_2538_),
    .Y(_2539_));
 sg13g2_buf_1 _3445_ (.A(_2539_),
    .X(_2540_));
 sg13g2_nand2_1 _3446_ (.Y(_2541_),
    .A(net65),
    .B(net121));
 sg13g2_nand3_1 _3447_ (.B(net126),
    .C(net69),
    .A(_2452_),
    .Y(_2542_));
 sg13g2_nand2_1 _3448_ (.Y(_2543_),
    .A(_2541_),
    .B(_2542_));
 sg13g2_a22oi_1 _3449_ (.Y(_2544_),
    .B1(net66),
    .B2(_2543_),
    .A2(_2536_),
    .A1(_2535_));
 sg13g2_nand3b_1 _3450_ (.B(_2530_),
    .C(_2544_),
    .Y(_2545_),
    .A_N(_2528_));
 sg13g2_buf_1 _3451_ (.A(_1948_),
    .X(_2546_));
 sg13g2_buf_1 _3452_ (.A(net217),
    .X(_2547_));
 sg13g2_buf_1 _3453_ (.A(net193),
    .X(_2548_));
 sg13g2_nand2_1 _3454_ (.Y(_2549_),
    .A(_2545_),
    .B(net156));
 sg13g2_buf_1 _3455_ (.A(net198),
    .X(_2550_));
 sg13g2_buf_1 _3456_ (.A(net155),
    .X(_2551_));
 sg13g2_nand2_1 _3457_ (.Y(_2552_),
    .A(_0780_),
    .B(net228));
 sg13g2_buf_1 _3458_ (.A(_2552_),
    .X(_2553_));
 sg13g2_nand2_1 _3459_ (.Y(_2554_),
    .A(net154),
    .B(_2429_));
 sg13g2_buf_1 _3460_ (.A(_2554_),
    .X(_2555_));
 sg13g2_nor2_2 _3461_ (.A(net207),
    .B(net64),
    .Y(_2556_));
 sg13g2_nand2_2 _3462_ (.Y(_2557_),
    .A(_1370_),
    .B(net225));
 sg13g2_nor2_2 _3463_ (.A(_2557_),
    .B(net70),
    .Y(_2558_));
 sg13g2_nor3_1 _3464_ (.A(net110),
    .B(_2556_),
    .C(_2558_),
    .Y(_2559_));
 sg13g2_buf_1 _3465_ (.A(net202),
    .X(_2560_));
 sg13g2_nor2_1 _3466_ (.A(net217),
    .B(net153),
    .Y(_2561_));
 sg13g2_inv_1 _3467_ (.Y(_2562_),
    .A(_2561_));
 sg13g2_nand2_1 _3468_ (.Y(_2563_),
    .A(_2506_),
    .B(net178));
 sg13g2_buf_1 _3469_ (.A(net74),
    .X(_2564_));
 sg13g2_nand2_1 _3470_ (.Y(_2565_),
    .A(_2563_),
    .B(net42));
 sg13g2_buf_1 _3471_ (.A(net164),
    .X(_2566_));
 sg13g2_nand2_1 _3472_ (.Y(_2567_),
    .A(_2565_),
    .B(net109));
 sg13g2_buf_2 _3473_ (.A(_2450_),
    .X(_2568_));
 sg13g2_nand2_1 _3474_ (.Y(_2569_),
    .A(_0845_),
    .B(net170));
 sg13g2_inv_1 _3475_ (.Y(_2570_),
    .A(_2569_));
 sg13g2_nor2_2 _3476_ (.A(_2097_),
    .B(_2533_),
    .Y(_2571_));
 sg13g2_nor3_2 _3477_ (.A(net108),
    .B(_2570_),
    .C(_2571_),
    .Y(_2572_));
 sg13g2_nor2_1 _3478_ (.A(_2567_),
    .B(_2572_),
    .Y(_2573_));
 sg13g2_nor3_1 _3479_ (.A(_2559_),
    .B(_2562_),
    .C(_2573_),
    .Y(_2574_));
 sg13g2_buf_1 _3480_ (.A(net196),
    .X(_2575_));
 sg13g2_nor2_1 _3481_ (.A(net205),
    .B(_2117_),
    .Y(_2576_));
 sg13g2_buf_2 _3482_ (.A(_2576_),
    .X(_2577_));
 sg13g2_nand2_1 _3483_ (.Y(_2578_),
    .A(_2577_),
    .B(net78));
 sg13g2_nor2_1 _3484_ (.A(net152),
    .B(_2578_),
    .Y(_2579_));
 sg13g2_nand2_1 _3485_ (.Y(_2580_),
    .A(_2300_),
    .B(net200));
 sg13g2_inv_1 _3486_ (.Y(_2581_),
    .A(_2580_));
 sg13g2_nor2_2 _3487_ (.A(net200),
    .B(_1828_),
    .Y(_2582_));
 sg13g2_a21oi_2 _3488_ (.B1(_2582_),
    .Y(_2583_),
    .A2(_2581_),
    .A1(net169));
 sg13g2_buf_1 _3489_ (.A(net79),
    .X(_2584_));
 sg13g2_nor2_2 _3490_ (.A(net180),
    .B(_1283_),
    .Y(_2585_));
 sg13g2_a21oi_1 _3491_ (.A1(net41),
    .A2(_2564_),
    .Y(_2586_),
    .B1(_2585_));
 sg13g2_o21ai_1 _3492_ (.B1(_2586_),
    .Y(_2587_),
    .A1(net109),
    .A2(_2583_));
 sg13g2_nor2_2 _3493_ (.A(_2500_),
    .B(_1948_),
    .Y(_2588_));
 sg13g2_o21ai_1 _3494_ (.B1(_2588_),
    .Y(_2589_),
    .A1(_2579_),
    .A2(_2587_));
 sg13g2_nor2b_1 _3495_ (.A(_2574_),
    .B_N(_2589_),
    .Y(_2590_));
 sg13g2_nand2_1 _3496_ (.Y(_2591_),
    .A(_2549_),
    .B(_2590_));
 sg13g2_buf_1 _3497_ (.A(_2411_),
    .X(_2592_));
 sg13g2_nor2_1 _3498_ (.A(net216),
    .B(net218),
    .Y(_2593_));
 sg13g2_buf_1 _3499_ (.A(_2593_),
    .X(_2594_));
 sg13g2_buf_1 _3500_ (.A(net111),
    .X(_2595_));
 sg13g2_nand2_1 _3501_ (.Y(_2596_),
    .A(net206),
    .B(_2300_));
 sg13g2_buf_2 _3502_ (.A(_2596_),
    .X(_2597_));
 sg13g2_nand2_1 _3503_ (.Y(_2598_),
    .A(_2495_),
    .B(net107));
 sg13g2_nand2_2 _3504_ (.Y(_2599_),
    .A(_2117_),
    .B(_2439_));
 sg13g2_inv_2 _3505_ (.Y(_2600_),
    .A(_2599_));
 sg13g2_a21oi_1 _3506_ (.A1(_2598_),
    .A2(net71),
    .Y(_2601_),
    .B1(_2600_));
 sg13g2_nand2_1 _3507_ (.Y(_2602_),
    .A(net154),
    .B(net173));
 sg13g2_a21oi_1 _3508_ (.A1(_2602_),
    .A2(net42),
    .Y(_2603_),
    .B1(net179));
 sg13g2_inv_1 _3509_ (.Y(_2604_),
    .A(_2318_));
 sg13g2_nor2_1 _3510_ (.A(net209),
    .B(_0758_),
    .Y(_2605_));
 sg13g2_buf_1 _3511_ (.A(_2605_),
    .X(_2606_));
 sg13g2_nor2_1 _3512_ (.A(_2604_),
    .B(net106),
    .Y(_2607_));
 sg13g2_nand2_1 _3513_ (.Y(_2608_),
    .A(_2607_),
    .B(net72));
 sg13g2_nand2_1 _3514_ (.Y(_2609_),
    .A(_2603_),
    .B(_2608_));
 sg13g2_o21ai_1 _3515_ (.B1(_2609_),
    .Y(_2610_),
    .A1(net63),
    .A2(_2601_));
 sg13g2_nor2_1 _3516_ (.A(_0955_),
    .B(_0987_),
    .Y(_2611_));
 sg13g2_buf_2 _3517_ (.A(_2611_),
    .X(_2612_));
 sg13g2_nor2_2 _3518_ (.A(_0966_),
    .B(_2612_),
    .Y(_2613_));
 sg13g2_nand2_1 _3519_ (.Y(_2614_),
    .A(_2613_),
    .B(net175));
 sg13g2_nand2_1 _3520_ (.Y(_2615_),
    .A(_2429_),
    .B(net210));
 sg13g2_nand2_1 _3521_ (.Y(_2616_),
    .A(_2614_),
    .B(_2615_));
 sg13g2_nand2_1 _3522_ (.Y(_2617_),
    .A(_2616_),
    .B(net42));
 sg13g2_nand2_2 _3523_ (.Y(_2618_),
    .A(net65),
    .B(_2533_));
 sg13g2_a21o_1 _3524_ (.A2(_2618_),
    .A1(_2617_),
    .B1(net67),
    .X(_2619_));
 sg13g2_nand2_1 _3525_ (.Y(_2620_),
    .A(_2519_),
    .B(_1283_));
 sg13g2_nor2_2 _3526_ (.A(net221),
    .B(_2097_),
    .Y(_2621_));
 sg13g2_nor2_1 _3527_ (.A(_2620_),
    .B(_2621_),
    .Y(_2622_));
 sg13g2_nand2_1 _3528_ (.Y(_2623_),
    .A(_2622_),
    .B(net132));
 sg13g2_buf_1 _3529_ (.A(net127),
    .X(_2624_));
 sg13g2_nand2_2 _3530_ (.Y(_2625_),
    .A(net81),
    .B(net205));
 sg13g2_nand3_1 _3531_ (.B(net62),
    .C(_2625_),
    .A(_2623_),
    .Y(_2626_));
 sg13g2_nand3b_1 _3532_ (.B(_2619_),
    .C(_2626_),
    .Y(_2627_),
    .A_N(_2610_));
 sg13g2_buf_1 _3533_ (.A(net217),
    .X(_2628_));
 sg13g2_buf_1 _3534_ (.A(net192),
    .X(_2629_));
 sg13g2_buf_1 _3535_ (.A(_2515_),
    .X(_2630_));
 sg13g2_nand2_1 _3536_ (.Y(_2631_),
    .A(net216),
    .B(net215));
 sg13g2_nor2_1 _3537_ (.A(net150),
    .B(_2631_),
    .Y(_2632_));
 sg13g2_nand2_1 _3538_ (.Y(_2633_),
    .A(_2627_),
    .B(_2632_));
 sg13g2_buf_1 _3539_ (.A(net157),
    .X(_2634_));
 sg13g2_inv_1 _3540_ (.Y(_2635_),
    .A(_0034_));
 sg13g2_nor4_1 _3541_ (.A(net105),
    .B(net218),
    .C(_2635_),
    .D(net165),
    .Y(_2636_));
 sg13g2_buf_1 _3542_ (.A(_2497_),
    .X(_2637_));
 sg13g2_nand2_1 _3543_ (.Y(_2638_),
    .A(net131),
    .B(_2637_));
 sg13g2_buf_2 _3544_ (.A(\memory_1.mem_addr[9] ),
    .X(_2639_));
 sg13g2_inv_1 _3545_ (.Y(_2640_),
    .A(_2639_));
 sg13g2_a21oi_1 _3546_ (.A1(_2636_),
    .A2(_2638_),
    .Y(_2641_),
    .B1(_2640_));
 sg13g2_nand2_1 _3547_ (.Y(_2642_),
    .A(_2633_),
    .B(_2641_));
 sg13g2_a21oi_1 _3548_ (.A1(_2591_),
    .A2(net151),
    .Y(_2643_),
    .B1(_2642_));
 sg13g2_inv_1 _3549_ (.Y(_2644_),
    .A(_2445_));
 sg13g2_a21oi_1 _3550_ (.A1(_2215_),
    .A2(_2318_),
    .Y(_2645_),
    .B1(net162));
 sg13g2_nor2_1 _3551_ (.A(_2644_),
    .B(_2645_),
    .Y(_2646_));
 sg13g2_nor2_1 _3552_ (.A(net225),
    .B(net210),
    .Y(_2647_));
 sg13g2_buf_1 _3553_ (.A(_2647_),
    .X(_2648_));
 sg13g2_nand2_1 _3554_ (.Y(_2649_),
    .A(net103),
    .B(net154));
 sg13g2_nand2_1 _3555_ (.Y(_2650_),
    .A(_2646_),
    .B(_2649_));
 sg13g2_nand2_1 _3556_ (.Y(_2651_),
    .A(_2650_),
    .B(net127));
 sg13g2_nand2_1 _3557_ (.Y(_2652_),
    .A(net177),
    .B(net176));
 sg13g2_inv_1 _3558_ (.Y(_2653_),
    .A(_2652_));
 sg13g2_a21oi_1 _3559_ (.A1(net79),
    .A2(net113),
    .Y(_2654_),
    .B1(_2653_));
 sg13g2_nand2_1 _3560_ (.Y(_2655_),
    .A(_0976_),
    .B(_2453_));
 sg13g2_nand2_2 _3561_ (.Y(_2656_),
    .A(_2655_),
    .B(_2390_));
 sg13g2_nand2_1 _3562_ (.Y(_2657_),
    .A(_2654_),
    .B(_2656_));
 sg13g2_buf_2 _3563_ (.A(_1435_),
    .X(_2658_));
 sg13g2_buf_1 _3564_ (.A(net149),
    .X(_2659_));
 sg13g2_nand2_1 _3565_ (.Y(_2660_),
    .A(_2657_),
    .B(net102));
 sg13g2_nand2_1 _3566_ (.Y(_2661_),
    .A(_2651_),
    .B(_2660_));
 sg13g2_nor2_2 _3567_ (.A(net224),
    .B(_1283_),
    .Y(_2662_));
 sg13g2_nor2_2 _3568_ (.A(_2625_),
    .B(_2662_),
    .Y(_2663_));
 sg13g2_inv_1 _3569_ (.Y(_2664_),
    .A(_2663_));
 sg13g2_buf_1 _3570_ (.A(net202),
    .X(_2665_));
 sg13g2_inv_2 _3571_ (.Y(_2666_),
    .A(net204));
 sg13g2_nor2_2 _3572_ (.A(net222),
    .B(_1828_),
    .Y(_2667_));
 sg13g2_nor3_1 _3573_ (.A(net148),
    .B(_2666_),
    .C(_2667_),
    .Y(_2668_));
 sg13g2_nand2_2 _3574_ (.Y(_2669_),
    .A(_2577_),
    .B(_2452_));
 sg13g2_nor2_2 _3575_ (.A(net225),
    .B(_1206_),
    .Y(_2670_));
 sg13g2_nand2_1 _3576_ (.Y(_2671_),
    .A(_2670_),
    .B(_1261_));
 sg13g2_nand3_1 _3577_ (.B(_2671_),
    .C(net153),
    .A(_2669_),
    .Y(_2672_));
 sg13g2_buf_1 _3578_ (.A(net219),
    .X(_2673_));
 sg13g2_nand2_1 _3579_ (.Y(_2674_),
    .A(_2672_),
    .B(net191));
 sg13g2_a21oi_1 _3580_ (.A1(_2664_),
    .A2(_2668_),
    .Y(_2675_),
    .B1(_2674_));
 sg13g2_nor2_1 _3581_ (.A(_2661_),
    .B(_2675_),
    .Y(_2676_));
 sg13g2_nor2_1 _3582_ (.A(net161),
    .B(_2676_),
    .Y(_2677_));
 sg13g2_nand2_1 _3583_ (.Y(_2678_),
    .A(_2234_),
    .B(net118));
 sg13g2_nand2_1 _3584_ (.Y(_2679_),
    .A(_2670_),
    .B(net154));
 sg13g2_a21oi_1 _3585_ (.A1(_2678_),
    .A2(_2679_),
    .Y(_2680_),
    .B1(_1468_));
 sg13g2_inv_1 _3586_ (.Y(_2681_),
    .A(_1828_));
 sg13g2_a21oi_1 _3587_ (.A1(net131),
    .A2(net104),
    .Y(_2682_),
    .B1(net118));
 sg13g2_o21ai_1 _3588_ (.B1(net115),
    .Y(_2683_),
    .A1(_2681_),
    .A2(_2682_));
 sg13g2_nand2b_1 _3589_ (.Y(_2684_),
    .B(_2683_),
    .A_N(_2680_));
 sg13g2_nand2_1 _3590_ (.Y(_2685_),
    .A(_1785_),
    .B(net162));
 sg13g2_buf_2 _3591_ (.A(_2685_),
    .X(_2686_));
 sg13g2_nand2_1 _3592_ (.Y(_2687_),
    .A(_2519_),
    .B(net178));
 sg13g2_nor2_1 _3593_ (.A(_2686_),
    .B(_2687_),
    .Y(_2688_));
 sg13g2_buf_1 _3594_ (.A(net204),
    .X(_2689_));
 sg13g2_nor2_1 _3595_ (.A(net147),
    .B(net46),
    .Y(_2690_));
 sg13g2_nand2_1 _3596_ (.Y(_2691_),
    .A(_1577_),
    .B(_2453_));
 sg13g2_nor2_1 _3597_ (.A(_2097_),
    .B(_2691_),
    .Y(_2692_));
 sg13g2_nor2_2 _3598_ (.A(net132),
    .B(_2692_),
    .Y(_2693_));
 sg13g2_o21ai_1 _3599_ (.B1(_2447_),
    .Y(_2694_),
    .A1(_2690_),
    .A2(_2693_));
 sg13g2_nand2b_1 _3600_ (.Y(_2695_),
    .B(_2694_),
    .A_N(_2688_));
 sg13g2_nor2_1 _3601_ (.A(_2684_),
    .B(_2695_),
    .Y(_2696_));
 sg13g2_nor2_1 _3602_ (.A(net165),
    .B(_2696_),
    .Y(_2697_));
 sg13g2_nor2_1 _3603_ (.A(_2677_),
    .B(_2697_),
    .Y(_2698_));
 sg13g2_nor2_1 _3604_ (.A(net225),
    .B(_2612_),
    .Y(_2699_));
 sg13g2_buf_1 _3605_ (.A(_2699_),
    .X(_2700_));
 sg13g2_buf_1 _3606_ (.A(_2525_),
    .X(_2701_));
 sg13g2_a21oi_1 _3607_ (.A1(net61),
    .A2(net126),
    .Y(_2702_),
    .B1(net60));
 sg13g2_nor2_2 _3608_ (.A(net205),
    .B(_1643_),
    .Y(_2703_));
 sg13g2_nand2_1 _3609_ (.Y(_2704_),
    .A(_2614_),
    .B(_2703_));
 sg13g2_buf_1 _3610_ (.A(_1162_),
    .X(_2705_));
 sg13g2_nor2_1 _3611_ (.A(net146),
    .B(_2556_),
    .Y(_2706_));
 sg13g2_a22oi_1 _3612_ (.Y(_2707_),
    .B1(_1555_),
    .B2(_2706_),
    .A2(_2704_),
    .A1(_2702_));
 sg13g2_inv_1 _3613_ (.Y(_2708_),
    .A(_2691_));
 sg13g2_nor2_1 _3614_ (.A(net207),
    .B(_2708_),
    .Y(_2709_));
 sg13g2_nor2_1 _3615_ (.A(net111),
    .B(_2709_),
    .Y(_2710_));
 sg13g2_buf_1 _3616_ (.A(net203),
    .X(_2711_));
 sg13g2_a21oi_1 _3617_ (.A1(_2710_),
    .A2(_1119_),
    .Y(_2712_),
    .B1(net145));
 sg13g2_inv_2 _3618_ (.Y(_2713_),
    .A(net106));
 sg13g2_buf_1 _3619_ (.A(net123),
    .X(_2714_));
 sg13g2_nand2_1 _3620_ (.Y(_2715_),
    .A(_2713_),
    .B(net59));
 sg13g2_a21o_1 _3621_ (.A2(_2715_),
    .A1(_2678_),
    .B1(net67),
    .X(_2716_));
 sg13g2_nand3_1 _3622_ (.B(_2712_),
    .C(_2716_),
    .A(_2707_),
    .Y(_2717_));
 sg13g2_inv_1 _3623_ (.Y(_2718_),
    .A(_2498_));
 sg13g2_nand2_1 _3624_ (.Y(_2719_),
    .A(_2429_),
    .B(net176));
 sg13g2_inv_2 _3625_ (.Y(_2720_),
    .A(_2719_));
 sg13g2_nor2_1 _3626_ (.A(net119),
    .B(_2720_),
    .Y(_2721_));
 sg13g2_nand2_1 _3627_ (.Y(_2722_),
    .A(_2718_),
    .B(_2721_));
 sg13g2_nand2_2 _3628_ (.Y(_2723_),
    .A(_1643_),
    .B(_2439_));
 sg13g2_nand2_2 _3629_ (.Y(_2724_),
    .A(_2723_),
    .B(_1763_));
 sg13g2_inv_2 _3630_ (.Y(_2725_),
    .A(_2724_));
 sg13g2_inv_1 _3631_ (.Y(_2726_),
    .A(_2435_));
 sg13g2_buf_1 _3632_ (.A(net196),
    .X(_2727_));
 sg13g2_a21oi_1 _3633_ (.A1(_2725_),
    .A2(_2726_),
    .Y(_2728_),
    .B1(net144));
 sg13g2_nand2_1 _3634_ (.Y(_2729_),
    .A(_2722_),
    .B(_2728_));
 sg13g2_nor2_1 _3635_ (.A(net111),
    .B(_2618_),
    .Y(_2730_));
 sg13g2_nand2_1 _3636_ (.Y(_2731_),
    .A(_1053_),
    .B(_1228_));
 sg13g2_nor2_1 _3637_ (.A(_0791_),
    .B(_1130_),
    .Y(_2732_));
 sg13g2_buf_2 _3638_ (.A(_2732_),
    .X(_2733_));
 sg13g2_inv_2 _3639_ (.Y(_2734_),
    .A(_2733_));
 sg13g2_nor2_2 _3640_ (.A(net198),
    .B(_2734_),
    .Y(_2735_));
 sg13g2_nand2_2 _3641_ (.Y(_2736_),
    .A(net154),
    .B(net222));
 sg13g2_nand2_1 _3642_ (.Y(_2737_),
    .A(_2735_),
    .B(_2736_));
 sg13g2_nor2_1 _3643_ (.A(_2731_),
    .B(_2737_),
    .Y(_2738_));
 sg13g2_nor3_1 _3644_ (.A(net193),
    .B(_2730_),
    .C(_2738_),
    .Y(_2739_));
 sg13g2_inv_1 _3645_ (.Y(_2740_),
    .A(_1882_));
 sg13g2_nand2_1 _3646_ (.Y(_2741_),
    .A(_2740_),
    .B(net129));
 sg13g2_nor2_1 _3647_ (.A(net177),
    .B(_2206_),
    .Y(_2742_));
 sg13g2_inv_1 _3648_ (.Y(_2743_),
    .A(_2742_));
 sg13g2_nand2_1 _3649_ (.Y(_2744_),
    .A(_2741_),
    .B(_2743_));
 sg13g2_nand3_1 _3650_ (.B(net154),
    .C(net131),
    .A(_2577_),
    .Y(_2745_));
 sg13g2_nand2_1 _3651_ (.Y(_2746_),
    .A(_2744_),
    .B(_2745_));
 sg13g2_nand2_1 _3652_ (.Y(_2747_),
    .A(_2746_),
    .B(net66));
 sg13g2_nand3_1 _3653_ (.B(_2739_),
    .C(_2747_),
    .A(_2729_),
    .Y(_2748_));
 sg13g2_buf_1 _3654_ (.A(net199),
    .X(_2749_));
 sg13g2_nand3_1 _3655_ (.B(_2748_),
    .C(net143),
    .A(_2717_),
    .Y(_2750_));
 sg13g2_buf_1 _3656_ (.A(net215),
    .X(_2751_));
 sg13g2_a21oi_1 _3657_ (.A1(_2698_),
    .A2(_2750_),
    .Y(_2752_),
    .B1(net190));
 sg13g2_nor2_1 _3658_ (.A(_2267_),
    .B(_2289_),
    .Y(_2753_));
 sg13g2_nor2_1 _3659_ (.A(_2753_),
    .B(_2663_),
    .Y(_2754_));
 sg13g2_nor2_1 _3660_ (.A(_1654_),
    .B(_2433_),
    .Y(_2755_));
 sg13g2_inv_2 _3661_ (.Y(_2756_),
    .A(_2755_));
 sg13g2_nand3_1 _3662_ (.B(_2175_),
    .C(net168),
    .A(_2756_),
    .Y(_2757_));
 sg13g2_nand2_1 _3663_ (.Y(_2758_),
    .A(_2754_),
    .B(_2757_));
 sg13g2_nand2_1 _3664_ (.Y(_2759_),
    .A(_2758_),
    .B(net116));
 sg13g2_nand2_1 _3665_ (.Y(_2760_),
    .A(_2485_),
    .B(net118));
 sg13g2_nand2_1 _3666_ (.Y(_2761_),
    .A(_0900_),
    .B(_0802_));
 sg13g2_buf_2 _3667_ (.A(_2761_),
    .X(_2762_));
 sg13g2_nand2_1 _3668_ (.Y(_2763_),
    .A(_2762_),
    .B(net158));
 sg13g2_nor2_1 _3669_ (.A(net155),
    .B(_2763_),
    .Y(_2764_));
 sg13g2_nand2_1 _3670_ (.Y(_2765_),
    .A(_2760_),
    .B(_2764_));
 sg13g2_inv_1 _3671_ (.Y(_2766_),
    .A(_2667_));
 sg13g2_nand2_1 _3672_ (.Y(_2767_),
    .A(_2766_),
    .B(net147));
 sg13g2_nand2_2 _3673_ (.Y(_2768_),
    .A(_0758_),
    .B(net206));
 sg13g2_buf_1 _3674_ (.A(_2390_),
    .X(_2769_));
 sg13g2_a21oi_1 _3675_ (.A1(_2768_),
    .A2(_2318_),
    .Y(_2770_),
    .B1(net101));
 sg13g2_buf_1 _3676_ (.A(_2459_),
    .X(_2771_));
 sg13g2_o21ai_1 _3677_ (.B1(net58),
    .Y(_2772_),
    .A1(_2767_),
    .A2(_2770_));
 sg13g2_nand3_1 _3678_ (.B(_2765_),
    .C(_2772_),
    .A(_2759_),
    .Y(_2773_));
 sg13g2_nand2_1 _3679_ (.Y(_2774_),
    .A(_2773_),
    .B(net125));
 sg13g2_nand2_2 _3680_ (.Y(_2775_),
    .A(net176),
    .B(net209));
 sg13g2_inv_1 _3681_ (.Y(_2776_),
    .A(_2775_));
 sg13g2_a21oi_2 _3682_ (.B1(_2585_),
    .Y(_2777_),
    .A2(_2776_),
    .A1(_1621_));
 sg13g2_nand2_1 _3683_ (.Y(_2778_),
    .A(_2777_),
    .B(_2444_));
 sg13g2_buf_1 _3684_ (.A(_1948_),
    .X(_2779_));
 sg13g2_nand3_1 _3685_ (.B(_2779_),
    .C(net102),
    .A(_2778_),
    .Y(_2780_));
 sg13g2_nand2_1 _3686_ (.Y(_2781_),
    .A(net81),
    .B(_0758_));
 sg13g2_nor2_2 _3687_ (.A(_2267_),
    .B(_2405_),
    .Y(_2782_));
 sg13g2_nand2_1 _3688_ (.Y(_2783_),
    .A(_1577_),
    .B(net223));
 sg13g2_buf_2 _3689_ (.A(_2783_),
    .X(_2784_));
 sg13g2_nand3_1 _3690_ (.B(net130),
    .C(net104),
    .A(_2784_),
    .Y(_2785_));
 sg13g2_nor2_1 _3691_ (.A(net177),
    .B(_2719_),
    .Y(_2786_));
 sg13g2_nor2_1 _3692_ (.A(net203),
    .B(_2525_),
    .Y(_2787_));
 sg13g2_nor2b_1 _3693_ (.A(_2786_),
    .B_N(_2787_),
    .Y(_2788_));
 sg13g2_a22oi_1 _3694_ (.Y(_2789_),
    .B1(_2785_),
    .B2(_2788_),
    .A2(_2782_),
    .A1(_2781_));
 sg13g2_nand2_1 _3695_ (.Y(_2790_),
    .A(_2780_),
    .B(_2789_));
 sg13g2_nand2_1 _3696_ (.Y(_2791_),
    .A(net154),
    .B(net81));
 sg13g2_nand2_1 _3697_ (.Y(_2792_),
    .A(_2791_),
    .B(net108));
 sg13g2_buf_1 _3698_ (.A(net195),
    .X(_2793_));
 sg13g2_a21o_1 _3699_ (.A2(_2792_),
    .A1(_2669_),
    .B1(net142),
    .X(_2794_));
 sg13g2_nand2_1 _3700_ (.Y(_2795_),
    .A(_2234_),
    .B(_2259_));
 sg13g2_a21oi_1 _3701_ (.A1(_2794_),
    .A2(_2795_),
    .Y(_2796_),
    .B1(_2405_));
 sg13g2_nor2_1 _3702_ (.A(_2790_),
    .B(_2796_),
    .Y(_2797_));
 sg13g2_nand2_1 _3703_ (.Y(_2798_),
    .A(_2774_),
    .B(_2797_));
 sg13g2_nand2_1 _3704_ (.Y(_2799_),
    .A(_2798_),
    .B(net151));
 sg13g2_nand2_1 _3705_ (.Y(_2800_),
    .A(net82),
    .B(_1261_));
 sg13g2_inv_1 _3706_ (.Y(_2801_),
    .A(_2800_));
 sg13g2_nand2_1 _3707_ (.Y(_2802_),
    .A(_2801_),
    .B(_2720_));
 sg13g2_a21oi_1 _3708_ (.A1(_2499_),
    .A2(_2802_),
    .Y(_2803_),
    .B1(net63));
 sg13g2_nand2_1 _3709_ (.Y(_2804_),
    .A(net44),
    .B(_2784_));
 sg13g2_buf_1 _3710_ (.A(net132),
    .X(_2805_));
 sg13g2_nand2_1 _3711_ (.Y(_2806_),
    .A(_2804_),
    .B(net57));
 sg13g2_nand2_1 _3712_ (.Y(_2807_),
    .A(_2756_),
    .B(_2439_));
 sg13g2_buf_1 _3713_ (.A(net179),
    .X(_2808_));
 sg13g2_a21oi_1 _3714_ (.A1(_2806_),
    .A2(_2807_),
    .Y(_2809_),
    .B1(net100));
 sg13g2_nor2_1 _3715_ (.A(_2803_),
    .B(_2809_),
    .Y(_2810_));
 sg13g2_nand2_2 _3716_ (.Y(_2811_),
    .A(_1283_),
    .B(net176));
 sg13g2_inv_1 _3717_ (.Y(_2812_),
    .A(_2811_));
 sg13g2_nand2_1 _3718_ (.Y(_2813_),
    .A(_2482_),
    .B(_2812_));
 sg13g2_nand2_1 _3719_ (.Y(_2814_),
    .A(_2731_),
    .B(net169));
 sg13g2_a21oi_1 _3720_ (.A1(_2813_),
    .A2(_2814_),
    .Y(_2815_),
    .B1(_2527_));
 sg13g2_nand2_1 _3721_ (.Y(_2816_),
    .A(net44),
    .B(_2720_));
 sg13g2_nand2_1 _3722_ (.Y(_2817_),
    .A(_2577_),
    .B(net83));
 sg13g2_nand2_1 _3723_ (.Y(_2818_),
    .A(_2816_),
    .B(_2817_));
 sg13g2_buf_2 _3724_ (.A(net149),
    .X(_2819_));
 sg13g2_nand2_1 _3725_ (.Y(_2820_),
    .A(_2818_),
    .B(net99));
 sg13g2_nand2_1 _3726_ (.Y(_2821_),
    .A(_2820_),
    .B(net193));
 sg13g2_nor2_1 _3727_ (.A(_2815_),
    .B(_2821_),
    .Y(_2822_));
 sg13g2_nand2_1 _3728_ (.Y(_2823_),
    .A(_2810_),
    .B(_2822_));
 sg13g2_a21oi_1 _3729_ (.A1(_1675_),
    .A2(net175),
    .Y(_2824_),
    .B1(net148));
 sg13g2_inv_2 _3730_ (.Y(_2825_),
    .A(net65));
 sg13g2_nand2_1 _3731_ (.Y(_2826_),
    .A(_2824_),
    .B(_2825_));
 sg13g2_nand2_1 _3732_ (.Y(_2827_),
    .A(_0758_),
    .B(net209));
 sg13g2_buf_2 _3733_ (.A(_2827_),
    .X(_2828_));
 sg13g2_nand2_2 _3734_ (.Y(_2829_),
    .A(_2828_),
    .B(net104));
 sg13g2_nor2_2 _3735_ (.A(_2398_),
    .B(net113),
    .Y(_2830_));
 sg13g2_nor2_1 _3736_ (.A(_2734_),
    .B(_2206_),
    .Y(_2831_));
 sg13g2_a21oi_1 _3737_ (.A1(_2829_),
    .A2(_2830_),
    .Y(_2832_),
    .B1(_2831_));
 sg13g2_nand2_1 _3738_ (.Y(_2833_),
    .A(_2826_),
    .B(_2832_));
 sg13g2_nand2_1 _3739_ (.Y(_2834_),
    .A(_2833_),
    .B(net75));
 sg13g2_nand2_1 _3740_ (.Y(_2835_),
    .A(_2829_),
    .B(net42));
 sg13g2_nand2_1 _3741_ (.Y(_2836_),
    .A(_2828_),
    .B(net107));
 sg13g2_nand2_1 _3742_ (.Y(_2837_),
    .A(_2836_),
    .B(net57));
 sg13g2_nand2_1 _3743_ (.Y(_2838_),
    .A(_2835_),
    .B(_2837_));
 sg13g2_buf_1 _3744_ (.A(_2447_),
    .X(_2839_));
 sg13g2_buf_1 _3745_ (.A(net192),
    .X(_2840_));
 sg13g2_a21oi_1 _3746_ (.A1(_2838_),
    .A2(net98),
    .Y(_2841_),
    .B1(net141));
 sg13g2_nor2_1 _3747_ (.A(net129),
    .B(_2117_),
    .Y(_2842_));
 sg13g2_inv_1 _3748_ (.Y(_2843_),
    .A(_2842_));
 sg13g2_nand2_1 _3749_ (.Y(_2844_),
    .A(_1315_),
    .B(_2843_));
 sg13g2_buf_2 _3750_ (.A(net58),
    .X(_2845_));
 sg13g2_nand2_1 _3751_ (.Y(_2846_),
    .A(_2844_),
    .B(net40));
 sg13g2_nand3_1 _3752_ (.B(_2841_),
    .C(_2846_),
    .A(_2834_),
    .Y(_2847_));
 sg13g2_inv_2 _3753_ (.Y(_2848_),
    .A(_2631_));
 sg13g2_nand3_1 _3754_ (.B(_2847_),
    .C(_2848_),
    .A(_2823_),
    .Y(_2849_));
 sg13g2_nand3_1 _3755_ (.B(_2849_),
    .C(_2640_),
    .A(_2799_),
    .Y(_2850_));
 sg13g2_nor2_1 _3756_ (.A(_2752_),
    .B(_2850_),
    .Y(_2851_));
 sg13g2_a21oi_1 _3757_ (.A1(_2518_),
    .A2(_2643_),
    .Y(_0016_),
    .B1(_2851_));
 sg13g2_nand2_1 _3758_ (.Y(_2852_),
    .A(_0758_),
    .B(_2453_));
 sg13g2_nor2_2 _3759_ (.A(_0802_),
    .B(_2852_),
    .Y(_2853_));
 sg13g2_inv_1 _3760_ (.Y(_2854_),
    .A(_2853_));
 sg13g2_nor2_1 _3761_ (.A(_1206_),
    .B(_2854_),
    .Y(_2855_));
 sg13g2_nand2_2 _3762_ (.Y(_2856_),
    .A(_2612_),
    .B(net205));
 sg13g2_nand2_1 _3763_ (.Y(_2857_),
    .A(_2856_),
    .B(net197));
 sg13g2_nor2_2 _3764_ (.A(net204),
    .B(_2455_),
    .Y(_2858_));
 sg13g2_nor2_1 _3765_ (.A(net197),
    .B(_2858_),
    .Y(_2859_));
 sg13g2_buf_1 _3766_ (.A(net164),
    .X(_2860_));
 sg13g2_a21oi_1 _3767_ (.A1(_2859_),
    .A2(_2649_),
    .Y(_2861_),
    .B1(net97));
 sg13g2_o21ai_1 _3768_ (.B1(_2861_),
    .Y(_2862_),
    .A1(_2855_),
    .A2(_2857_));
 sg13g2_buf_1 _3769_ (.A(_1839_),
    .X(_2863_));
 sg13g2_nand2_1 _3770_ (.Y(_2864_),
    .A(net96),
    .B(net160));
 sg13g2_o21ai_1 _3771_ (.B1(_2864_),
    .Y(_2865_),
    .A1(_2811_),
    .A2(net64));
 sg13g2_a21oi_1 _3772_ (.A1(_2865_),
    .A2(net99),
    .Y(_2866_),
    .B1(_2688_));
 sg13g2_a21oi_1 _3773_ (.A1(_2862_),
    .A2(_2866_),
    .Y(_2867_),
    .B1(_2417_));
 sg13g2_nand2_1 _3774_ (.Y(_2868_),
    .A(net207),
    .B(_1140_));
 sg13g2_nor2_1 _3775_ (.A(net175),
    .B(_2868_),
    .Y(_2869_));
 sg13g2_nor2_1 _3776_ (.A(_1337_),
    .B(_2455_),
    .Y(_2870_));
 sg13g2_buf_1 _3777_ (.A(_2870_),
    .X(_2871_));
 sg13g2_nor2_2 _3778_ (.A(_1283_),
    .B(_1337_),
    .Y(_2872_));
 sg13g2_nor2_1 _3779_ (.A(net56),
    .B(_2872_),
    .Y(_2873_));
 sg13g2_a21oi_1 _3780_ (.A1(_2873_),
    .A2(net172),
    .Y(_2874_),
    .B1(net164));
 sg13g2_inv_1 _3781_ (.Y(_2875_),
    .A(_2399_));
 sg13g2_nand2_1 _3782_ (.Y(_2876_),
    .A(_2708_),
    .B(net113));
 sg13g2_nand2_1 _3783_ (.Y(_2877_),
    .A(net168),
    .B(_2433_));
 sg13g2_buf_2 _3784_ (.A(_2877_),
    .X(_2878_));
 sg13g2_nand3_1 _3785_ (.B(_2876_),
    .C(_2878_),
    .A(_2875_),
    .Y(_2879_));
 sg13g2_o21ai_1 _3786_ (.B1(_2879_),
    .Y(_2880_),
    .A1(_2869_),
    .A2(_2874_));
 sg13g2_nand2_1 _3787_ (.Y(_2881_),
    .A(_2471_),
    .B(net130));
 sg13g2_buf_1 _3788_ (.A(net158),
    .X(_2882_));
 sg13g2_nand3_1 _3789_ (.B(net95),
    .C(_2843_),
    .A(_2881_),
    .Y(_2883_));
 sg13g2_nor2_1 _3790_ (.A(net221),
    .B(_1206_),
    .Y(_2884_));
 sg13g2_nand2_2 _3791_ (.Y(_2885_),
    .A(_2884_),
    .B(net180));
 sg13g2_nand3_1 _3792_ (.B(net197),
    .C(_0922_),
    .A(_2885_),
    .Y(_2886_));
 sg13g2_nor2b_1 _3793_ (.A(net196),
    .B_N(_2886_),
    .Y(_2887_));
 sg13g2_nand2_1 _3794_ (.Y(_2888_),
    .A(_2883_),
    .B(_2887_));
 sg13g2_nand2_1 _3795_ (.Y(_2889_),
    .A(_2880_),
    .B(_2888_));
 sg13g2_buf_1 _3796_ (.A(_2468_),
    .X(_2890_));
 sg13g2_nand2_1 _3797_ (.Y(_2891_),
    .A(_2889_),
    .B(net140));
 sg13g2_nand2b_1 _3798_ (.Y(_2892_),
    .B(_2891_),
    .A_N(_2867_));
 sg13g2_nor2_2 _3799_ (.A(net168),
    .B(_2703_),
    .Y(_2893_));
 sg13g2_nor2_1 _3800_ (.A(_2662_),
    .B(_2893_),
    .Y(_2894_));
 sg13g2_inv_1 _3801_ (.Y(_2895_),
    .A(_2894_));
 sg13g2_nand3_1 _3802_ (.B(net114),
    .C(_2077_),
    .A(_2895_),
    .Y(_2896_));
 sg13g2_inv_1 _3803_ (.Y(_2897_),
    .A(_2762_));
 sg13g2_nor2_1 _3804_ (.A(_1239_),
    .B(_2612_),
    .Y(_2898_));
 sg13g2_nand2_1 _3805_ (.Y(_2899_),
    .A(_2897_),
    .B(_2898_));
 sg13g2_inv_1 _3806_ (.Y(_2900_),
    .A(_2899_));
 sg13g2_o21ai_1 _3807_ (.B1(net102),
    .Y(_2901_),
    .A1(_2858_),
    .A2(_2900_));
 sg13g2_nand3_1 _3808_ (.B(net193),
    .C(_2901_),
    .A(_2896_),
    .Y(_2902_));
 sg13g2_nand2_1 _3809_ (.Y(_2903_),
    .A(net209),
    .B(_0038_));
 sg13g2_buf_1 _3810_ (.A(_2903_),
    .X(_2904_));
 sg13g2_nand2_2 _3811_ (.Y(_2905_),
    .A(_2713_),
    .B(net94));
 sg13g2_a22oi_1 _3812_ (.Y(_2906_),
    .B1(net45),
    .B2(_2905_),
    .A2(net81),
    .A1(_2666_));
 sg13g2_inv_1 _3813_ (.Y(_2907_),
    .A(_2814_));
 sg13g2_o21ai_1 _3814_ (.B1(net58),
    .Y(_2908_),
    .A1(_2600_),
    .A2(_2907_));
 sg13g2_o21ai_1 _3815_ (.B1(_2908_),
    .Y(_2909_),
    .A1(_2595_),
    .A2(_2906_));
 sg13g2_nor2_1 _3816_ (.A(_2902_),
    .B(_2909_),
    .Y(_2910_));
 sg13g2_a21oi_2 _3817_ (.B1(net101),
    .Y(_2911_),
    .A2(_2597_),
    .A1(net131));
 sg13g2_o21ai_1 _3818_ (.B1(net115),
    .Y(_2912_),
    .A1(_2582_),
    .A2(_2911_));
 sg13g2_nand2_2 _3819_ (.Y(_2913_),
    .A(net64),
    .B(net103));
 sg13g2_nor2_1 _3820_ (.A(net176),
    .B(net173),
    .Y(_2914_));
 sg13g2_inv_1 _3821_ (.Y(_2915_),
    .A(_2914_));
 sg13g2_nand2_1 _3822_ (.Y(_2916_),
    .A(_2913_),
    .B(_2915_));
 sg13g2_nand2_1 _3823_ (.Y(_2917_),
    .A(_2916_),
    .B(net127));
 sg13g2_nand3_1 _3824_ (.B(_2811_),
    .C(_2447_),
    .A(_2557_),
    .Y(_2918_));
 sg13g2_inv_1 _3825_ (.Y(_2919_),
    .A(_0036_));
 sg13g2_buf_1 _3826_ (.A(_2919_),
    .X(_2920_));
 sg13g2_nand2_1 _3827_ (.Y(_2921_),
    .A(_1435_),
    .B(net213));
 sg13g2_inv_1 _3828_ (.Y(_2922_),
    .A(_2921_));
 sg13g2_a21oi_1 _3829_ (.A1(_2922_),
    .A2(_2884_),
    .Y(_2923_),
    .B1(net214));
 sg13g2_nand4_1 _3830_ (.B(_2917_),
    .C(_2918_),
    .A(_2912_),
    .Y(_2924_),
    .D(_2923_));
 sg13g2_nand2_1 _3831_ (.Y(_2925_),
    .A(_2924_),
    .B(net199));
 sg13g2_nor2_1 _3832_ (.A(_2910_),
    .B(_2925_),
    .Y(_2926_));
 sg13g2_nor2_1 _3833_ (.A(_2892_),
    .B(_2926_),
    .Y(_2927_));
 sg13g2_nor2_1 _3834_ (.A(net190),
    .B(_2927_),
    .Y(_2928_));
 sg13g2_nor2_1 _3835_ (.A(_2380_),
    .B(_2507_),
    .Y(_2929_));
 sg13g2_nand2_1 _3836_ (.Y(_2930_),
    .A(_2929_),
    .B(net148));
 sg13g2_nand2_1 _3837_ (.Y(_2931_),
    .A(_2930_),
    .B(net155));
 sg13g2_nand2_1 _3838_ (.Y(_2932_),
    .A(net79),
    .B(net206));
 sg13g2_nand3_1 _3839_ (.B(net123),
    .C(_2828_),
    .A(_2932_),
    .Y(_2933_));
 sg13g2_inv_2 _3840_ (.Y(_2934_),
    .A(_2933_));
 sg13g2_nor3_1 _3841_ (.A(_2753_),
    .B(_2931_),
    .C(_2934_),
    .Y(_2935_));
 sg13g2_nor2_1 _3842_ (.A(_2066_),
    .B(_2768_),
    .Y(_2936_));
 sg13g2_inv_1 _3843_ (.Y(_2937_),
    .A(net56));
 sg13g2_nand2_2 _3844_ (.Y(_2938_),
    .A(_2937_),
    .B(net202));
 sg13g2_inv_1 _3845_ (.Y(_2939_),
    .A(_2938_));
 sg13g2_nand2_1 _3846_ (.Y(_2940_),
    .A(_2939_),
    .B(_2673_));
 sg13g2_nor2_1 _3847_ (.A(_2762_),
    .B(_2613_),
    .Y(_2941_));
 sg13g2_nand2_2 _3848_ (.Y(_2942_),
    .A(_2713_),
    .B(_2828_));
 sg13g2_nand2_1 _3849_ (.Y(_2943_),
    .A(_2942_),
    .B(_2462_));
 sg13g2_nand3b_1 _3850_ (.B(_2943_),
    .C(net58),
    .Y(_2944_),
    .A_N(_2941_));
 sg13g2_o21ai_1 _3851_ (.B1(_2944_),
    .Y(_2945_),
    .A1(_2936_),
    .A2(_2940_));
 sg13g2_buf_1 _3852_ (.A(net174),
    .X(_2946_));
 sg13g2_buf_1 _3853_ (.A(net93),
    .X(_2947_));
 sg13g2_o21ai_1 _3854_ (.B1(_2947_),
    .Y(_2948_),
    .A1(_2935_),
    .A2(_2945_));
 sg13g2_inv_1 _3855_ (.Y(_2949_),
    .A(_2594_));
 sg13g2_nand2_1 _3856_ (.Y(_2950_),
    .A(net121),
    .B(_2318_));
 sg13g2_nand2_2 _3857_ (.Y(_2951_),
    .A(_2950_),
    .B(net61));
 sg13g2_a21oi_1 _3858_ (.A1(_2951_),
    .A2(_2854_),
    .Y(_2952_),
    .B1(net179));
 sg13g2_nand3_1 _3859_ (.B(net101),
    .C(net107),
    .A(_2482_),
    .Y(_2953_));
 sg13g2_nand2_1 _3860_ (.Y(_2954_),
    .A(_2670_),
    .B(_2453_));
 sg13g2_nand3_1 _3861_ (.B(net127),
    .C(_2954_),
    .A(_2953_),
    .Y(_2955_));
 sg13g2_nand2b_1 _3862_ (.Y(_2956_),
    .B(_2955_),
    .A_N(_2952_));
 sg13g2_nor3_1 _3863_ (.A(_2681_),
    .B(net128),
    .C(_2736_),
    .Y(_2957_));
 sg13g2_a21oi_1 _3864_ (.A1(_2792_),
    .A2(_2885_),
    .Y(_2958_),
    .B1(net111));
 sg13g2_nor3_1 _3865_ (.A(net174),
    .B(_2957_),
    .C(_2958_),
    .Y(_2959_));
 sg13g2_nor2b_1 _3866_ (.A(_2956_),
    .B_N(_2959_),
    .Y(_2960_));
 sg13g2_nor2_1 _3867_ (.A(_2949_),
    .B(_2960_),
    .Y(_2961_));
 sg13g2_a21oi_1 _3868_ (.A1(_2948_),
    .A2(_2961_),
    .Y(_2962_),
    .B1(_2639_));
 sg13g2_nand2_2 _3869_ (.Y(_2963_),
    .A(_1850_),
    .B(net180));
 sg13g2_nor2_1 _3870_ (.A(net206),
    .B(_1512_),
    .Y(_2964_));
 sg13g2_nor2_1 _3871_ (.A(_2963_),
    .B(_2964_),
    .Y(_2965_));
 sg13g2_inv_1 _3872_ (.Y(_2966_),
    .A(_2965_));
 sg13g2_buf_1 _3873_ (.A(net153),
    .X(_2967_));
 sg13g2_inv_2 _3874_ (.Y(_2968_),
    .A(net94));
 sg13g2_o21ai_1 _3875_ (.B1(net59),
    .Y(_2969_),
    .A1(_2968_),
    .A2(_2461_));
 sg13g2_nand3_1 _3876_ (.B(net92),
    .C(_2969_),
    .A(_2966_),
    .Y(_2970_));
 sg13g2_buf_1 _3877_ (.A(net158),
    .X(_2971_));
 sg13g2_inv_1 _3878_ (.Y(_2972_),
    .A(_1261_));
 sg13g2_inv_2 _3879_ (.Y(_2973_),
    .A(_1839_));
 sg13g2_nor2_1 _3880_ (.A(_2972_),
    .B(_2973_),
    .Y(_2974_));
 sg13g2_nor2_1 _3881_ (.A(net91),
    .B(_2974_),
    .Y(_2975_));
 sg13g2_nand2_2 _3882_ (.Y(_2976_),
    .A(_2424_),
    .B(_2439_));
 sg13g2_a21oi_1 _3883_ (.A1(_2975_),
    .A2(_2976_),
    .Y(_2977_),
    .B1(net109));
 sg13g2_nand2_1 _3884_ (.Y(_2978_),
    .A(_2970_),
    .B(_2977_));
 sg13g2_nand2_1 _3885_ (.Y(_2979_),
    .A(_2507_),
    .B(net108));
 sg13g2_nor2_1 _3886_ (.A(net204),
    .B(_2215_),
    .Y(_2980_));
 sg13g2_inv_1 _3887_ (.Y(_2981_),
    .A(_2980_));
 sg13g2_nand2_1 _3888_ (.Y(_2982_),
    .A(_2979_),
    .B(_2981_));
 sg13g2_buf_1 _3889_ (.A(net114),
    .X(_2983_));
 sg13g2_buf_2 _3890_ (.A(net102),
    .X(_2984_));
 sg13g2_inv_1 _3891_ (.Y(_2985_),
    .A(_2786_));
 sg13g2_nand2_1 _3892_ (.Y(_2986_),
    .A(net107),
    .B(net175));
 sg13g2_nand2_1 _3893_ (.Y(_2987_),
    .A(_2986_),
    .B(net57));
 sg13g2_nand2_1 _3894_ (.Y(_2988_),
    .A(_2985_),
    .B(_2987_));
 sg13g2_a22oi_1 _3895_ (.Y(_2989_),
    .B1(net53),
    .B2(_2988_),
    .A2(net54),
    .A1(_2982_));
 sg13g2_a21oi_1 _3896_ (.A1(_2978_),
    .A2(_2989_),
    .Y(_2990_),
    .B1(net165));
 sg13g2_nand2_1 _3897_ (.Y(_2991_),
    .A(_2829_),
    .B(net72));
 sg13g2_a21oi_1 _3898_ (.A1(_2991_),
    .A2(_2951_),
    .Y(_2992_),
    .B1(net67));
 sg13g2_nor2_1 _3899_ (.A(net170),
    .B(_2383_),
    .Y(_2993_));
 sg13g2_nor2_1 _3900_ (.A(_2666_),
    .B(_2993_),
    .Y(_2994_));
 sg13g2_nand2_2 _3901_ (.Y(_2995_),
    .A(_2056_),
    .B(_1261_));
 sg13g2_nand2_1 _3902_ (.Y(_2996_),
    .A(_2995_),
    .B(net108));
 sg13g2_o21ai_1 _3903_ (.B1(_2996_),
    .Y(_2997_),
    .A1(_2492_),
    .A2(_2994_));
 sg13g2_buf_1 _3904_ (.A(net220),
    .X(_2998_));
 sg13g2_buf_1 _3905_ (.A(net189),
    .X(_2999_));
 sg13g2_nand2_1 _3906_ (.Y(_3000_),
    .A(_2997_),
    .B(_2999_));
 sg13g2_inv_1 _3907_ (.Y(_3001_),
    .A(_2852_));
 sg13g2_buf_1 _3908_ (.A(_0036_),
    .X(_3002_));
 sg13g2_nand2_1 _3909_ (.Y(_3003_),
    .A(_1097_),
    .B(net226));
 sg13g2_inv_1 _3910_ (.Y(_3004_),
    .A(_3003_));
 sg13g2_nor2_1 _3911_ (.A(net159),
    .B(_3004_),
    .Y(_3005_));
 sg13g2_a22oi_1 _3912_ (.Y(_3006_),
    .B1(net115),
    .B2(_2446_),
    .A2(_3005_),
    .A1(_3001_));
 sg13g2_nand2_1 _3913_ (.Y(_3007_),
    .A(_3000_),
    .B(_3006_));
 sg13g2_nor2_1 _3914_ (.A(_2992_),
    .B(_3007_),
    .Y(_3008_));
 sg13g2_nor2_1 _3915_ (.A(net161),
    .B(_3008_),
    .Y(_3009_));
 sg13g2_buf_1 _3916_ (.A(net215),
    .X(_3010_));
 sg13g2_o21ai_1 _3917_ (.B1(net188),
    .Y(_3011_),
    .A1(_2990_),
    .A2(_3009_));
 sg13g2_nand2_1 _3918_ (.Y(_3012_),
    .A(_2962_),
    .B(_3011_));
 sg13g2_nor2_1 _3919_ (.A(_2928_),
    .B(_3012_),
    .Y(_3013_));
 sg13g2_inv_2 _3920_ (.Y(_3014_),
    .A(_1719_));
 sg13g2_nand2_1 _3921_ (.Y(_3015_),
    .A(_1763_),
    .B(_2919_));
 sg13g2_nor2_2 _3922_ (.A(net198),
    .B(_3015_),
    .Y(_3016_));
 sg13g2_nand2_1 _3923_ (.Y(_3017_),
    .A(net79),
    .B(net96));
 sg13g2_nor2_1 _3924_ (.A(net80),
    .B(net117),
    .Y(_3018_));
 sg13g2_inv_1 _3925_ (.Y(_3019_),
    .A(_2381_));
 sg13g2_a21oi_1 _3926_ (.A1(_2951_),
    .A2(_3019_),
    .Y(_3020_),
    .B1(net146));
 sg13g2_a221oi_1 _3927_ (.B2(_3018_),
    .C1(_3020_),
    .B1(_3017_),
    .A1(_3014_),
    .Y(_3021_),
    .A2(_3016_));
 sg13g2_nand2_1 _3928_ (.Y(_3022_),
    .A(_3021_),
    .B(net156));
 sg13g2_a21oi_1 _3929_ (.A1(net131),
    .A2(_2597_),
    .Y(_3023_),
    .B1(net69));
 sg13g2_nor2_2 _3930_ (.A(net129),
    .B(_2434_),
    .Y(_3024_));
 sg13g2_nor2_1 _3931_ (.A(net195),
    .B(_3024_),
    .Y(_3025_));
 sg13g2_nand2b_1 _3932_ (.Y(_3026_),
    .B(_3025_),
    .A_N(_3023_));
 sg13g2_nor2_1 _3933_ (.A(net202),
    .B(_2504_),
    .Y(_3027_));
 sg13g2_inv_1 _3934_ (.Y(_3028_),
    .A(_2582_));
 sg13g2_nand2_1 _3935_ (.Y(_3029_),
    .A(_3027_),
    .B(_3028_));
 sg13g2_nand3_1 _3936_ (.B(_3029_),
    .C(net75),
    .A(_3026_),
    .Y(_3030_));
 sg13g2_nand2_2 _3937_ (.Y(_3031_),
    .A(_2097_),
    .B(_0998_));
 sg13g2_nand2_2 _3938_ (.Y(_3032_),
    .A(_2137_),
    .B(_3031_));
 sg13g2_nand2_1 _3939_ (.Y(_3033_),
    .A(_3032_),
    .B(net101));
 sg13g2_nor2_2 _3940_ (.A(net207),
    .B(net173),
    .Y(_3034_));
 sg13g2_inv_1 _3941_ (.Y(_3035_),
    .A(_3034_));
 sg13g2_nand2_1 _3942_ (.Y(_3036_),
    .A(_3033_),
    .B(_3035_));
 sg13g2_a21oi_1 _3943_ (.A1(_3036_),
    .A2(net98),
    .Y(_3037_),
    .B1(net141));
 sg13g2_nand2_1 _3944_ (.Y(_3038_),
    .A(_2556_),
    .B(net160));
 sg13g2_a21o_1 _3945_ (.A2(_3017_),
    .A1(_3038_),
    .B1(net100),
    .X(_3039_));
 sg13g2_nand3_1 _3946_ (.B(_3037_),
    .C(_3039_),
    .A(_3030_),
    .Y(_3040_));
 sg13g2_buf_1 _3947_ (.A(net216),
    .X(_3041_));
 sg13g2_buf_1 _3948_ (.A(net187),
    .X(_3042_));
 sg13g2_nand3_1 _3949_ (.B(_3040_),
    .C(net138),
    .A(_3022_),
    .Y(_3043_));
 sg13g2_buf_1 _3950_ (.A(net216),
    .X(_3044_));
 sg13g2_inv_2 _3951_ (.Y(_3045_),
    .A(_2352_));
 sg13g2_nand2_1 _3952_ (.Y(_3046_),
    .A(_2045_),
    .B(net94));
 sg13g2_nand2_1 _3953_ (.Y(_3047_),
    .A(_3046_),
    .B(net72));
 sg13g2_nor2_2 _3954_ (.A(net95),
    .B(net56),
    .Y(_3048_));
 sg13g2_nand2_2 _3955_ (.Y(_3049_),
    .A(_1261_),
    .B(_2497_));
 sg13g2_nand2_1 _3956_ (.Y(_3050_),
    .A(_3049_),
    .B(net74));
 sg13g2_nor2_2 _3957_ (.A(net123),
    .B(_2555_),
    .Y(_3051_));
 sg13g2_nor2_1 _3958_ (.A(net157),
    .B(_3051_),
    .Y(_3052_));
 sg13g2_a22oi_1 _3959_ (.Y(_3053_),
    .B1(_3050_),
    .B2(_3052_),
    .A2(_3048_),
    .A1(_3047_));
 sg13g2_nand2_1 _3960_ (.Y(_3054_),
    .A(_2578_),
    .B(_2665_));
 sg13g2_a21oi_1 _3961_ (.A1(_1042_),
    .A2(net113),
    .Y(_3055_),
    .B1(_2165_));
 sg13g2_inv_1 _3962_ (.Y(_0088_),
    .A(_3055_));
 sg13g2_o21ai_1 _3963_ (.B1(_0088_),
    .Y(_0089_),
    .A1(_2682_),
    .A2(_3054_));
 sg13g2_nand2_1 _3964_ (.Y(_0090_),
    .A(_0089_),
    .B(net167));
 sg13g2_o21ai_1 _3965_ (.B1(_0090_),
    .Y(_0091_),
    .A1(_3045_),
    .A2(_3053_));
 sg13g2_nor2_1 _3966_ (.A(net186),
    .B(_0091_),
    .Y(_0092_));
 sg13g2_nand2_2 _3967_ (.Y(_0093_),
    .A(net177),
    .B(net207));
 sg13g2_inv_1 _3968_ (.Y(_0094_),
    .A(_0093_));
 sg13g2_nor2_1 _3969_ (.A(net95),
    .B(_0094_),
    .Y(_0095_));
 sg13g2_nor2_1 _3970_ (.A(net189),
    .B(_2381_),
    .Y(_0096_));
 sg13g2_a21oi_1 _3971_ (.A1(_2720_),
    .A2(net79),
    .Y(_0097_),
    .B1(_2993_));
 sg13g2_a22oi_1 _3972_ (.Y(_0098_),
    .B1(_0096_),
    .B2(_0097_),
    .A2(_0095_),
    .A1(_2951_));
 sg13g2_nor2_1 _3973_ (.A(net201),
    .B(_2612_),
    .Y(_0099_));
 sg13g2_nor2_1 _3974_ (.A(net80),
    .B(_0099_),
    .Y(_0100_));
 sg13g2_nor3_1 _3975_ (.A(net68),
    .B(_3014_),
    .C(_2936_),
    .Y(_0101_));
 sg13g2_a21oi_1 _3976_ (.A1(_2744_),
    .A2(_0100_),
    .Y(_0102_),
    .B1(_0101_));
 sg13g2_o21ai_1 _3977_ (.B1(_0102_),
    .Y(_0103_),
    .A1(net75),
    .A2(_0098_));
 sg13g2_nand2_1 _3978_ (.Y(_0104_),
    .A(_0103_),
    .B(net55));
 sg13g2_nand2_1 _3979_ (.Y(_0105_),
    .A(_0092_),
    .B(_0104_));
 sg13g2_nand2_1 _3980_ (.Y(_0106_),
    .A(_3043_),
    .B(_0105_));
 sg13g2_nand2_2 _3981_ (.Y(_0107_),
    .A(net73),
    .B(net220));
 sg13g2_a21oi_2 _3982_ (.B1(net162),
    .Y(_0108_),
    .A2(net222),
    .A1(_2553_));
 sg13g2_nand2_1 _3983_ (.Y(_0109_),
    .A(_0108_),
    .B(net64));
 sg13g2_inv_1 _3984_ (.Y(_0110_),
    .A(_0109_));
 sg13g2_nor2_1 _3985_ (.A(net189),
    .B(_2489_),
    .Y(_0111_));
 sg13g2_a21oi_1 _3986_ (.A1(_0111_),
    .A2(_2878_),
    .Y(_0112_),
    .B1(net110));
 sg13g2_o21ai_1 _3987_ (.B1(_0112_),
    .Y(_0113_),
    .A1(_0107_),
    .A2(_0110_));
 sg13g2_buf_1 _3988_ (.A(net99),
    .X(_0114_));
 sg13g2_o21ai_1 _3989_ (.B1(net52),
    .Y(_0115_),
    .A1(_0094_),
    .A2(_0867_));
 sg13g2_nand2_1 _3990_ (.Y(_0116_),
    .A(net64),
    .B(net108));
 sg13g2_nand3_1 _3991_ (.B(net62),
    .C(_0116_),
    .A(_2745_),
    .Y(_0117_));
 sg13g2_buf_1 _3992_ (.A(net149),
    .X(_0118_));
 sg13g2_a21oi_1 _3993_ (.A1(_1882_),
    .A2(net90),
    .Y(_0119_),
    .B1(net145));
 sg13g2_nand4_1 _3994_ (.B(_0115_),
    .C(_0117_),
    .A(_0113_),
    .Y(_0120_),
    .D(_0119_));
 sg13g2_inv_1 _3995_ (.Y(_0121_),
    .A(_2625_));
 sg13g2_nor2_1 _3996_ (.A(net162),
    .B(_2483_),
    .Y(_0122_));
 sg13g2_buf_2 _3997_ (.A(_0122_),
    .X(_0123_));
 sg13g2_nor3_1 _3998_ (.A(net43),
    .B(_0121_),
    .C(_0123_),
    .Y(_0124_));
 sg13g2_inv_1 _3999_ (.Y(_0125_),
    .A(_2534_));
 sg13g2_nand2_1 _4000_ (.Y(_0126_),
    .A(_2756_),
    .B(net45));
 sg13g2_nand3_1 _4001_ (.B(_0126_),
    .C(net66),
    .A(_0125_),
    .Y(_0127_));
 sg13g2_nor2_1 _4002_ (.A(net163),
    .B(net103),
    .Y(_0128_));
 sg13g2_o21ai_1 _4003_ (.B1(_0128_),
    .Y(_0129_),
    .A1(net109),
    .A2(_2878_));
 sg13g2_nand2_1 _4004_ (.Y(_0130_),
    .A(_0127_),
    .B(_0129_));
 sg13g2_o21ai_1 _4005_ (.B1(net55),
    .Y(_0131_),
    .A1(_0124_),
    .A2(_0130_));
 sg13g2_nand3_1 _4006_ (.B(_0131_),
    .C(net151),
    .A(_0120_),
    .Y(_0132_));
 sg13g2_inv_1 _4007_ (.Y(_0133_),
    .A(_2995_));
 sg13g2_buf_1 _4008_ (.A(net132),
    .X(_0134_));
 sg13g2_nand2_1 _4009_ (.Y(_0135_),
    .A(_0133_),
    .B(net51));
 sg13g2_buf_2 _4010_ (.A(net197),
    .X(_0136_));
 sg13g2_nor2_2 _4011_ (.A(net221),
    .B(_0758_),
    .Y(_0137_));
 sg13g2_nor2_1 _4012_ (.A(net132),
    .B(_0137_),
    .Y(_0138_));
 sg13g2_nor2_2 _4013_ (.A(net137),
    .B(_0138_),
    .Y(_0139_));
 sg13g2_buf_1 _4014_ (.A(net219),
    .X(_0140_));
 sg13g2_buf_1 _4015_ (.A(net185),
    .X(_0141_));
 sg13g2_nand3_1 _4016_ (.B(_0139_),
    .C(net136),
    .A(_0135_),
    .Y(_0142_));
 sg13g2_nor2_1 _4017_ (.A(_1206_),
    .B(_2963_),
    .Y(_0143_));
 sg13g2_o21ai_1 _4018_ (.B1(net52),
    .Y(_0144_),
    .A1(_0143_),
    .A2(_0867_));
 sg13g2_nand2_1 _4019_ (.Y(_0145_),
    .A(_2878_),
    .B(_2856_));
 sg13g2_nor2_1 _4020_ (.A(net60),
    .B(_2687_),
    .Y(_0146_));
 sg13g2_a22oi_1 _4021_ (.Y(_0147_),
    .B1(_3035_),
    .B2(_0146_),
    .A2(net66),
    .A1(_0145_));
 sg13g2_nand3_1 _4022_ (.B(_0144_),
    .C(_0147_),
    .A(_0142_),
    .Y(_0148_));
 sg13g2_buf_2 _4023_ (.A(_0035_),
    .X(_0149_));
 sg13g2_nand2_1 _4024_ (.Y(_0150_),
    .A(_0034_),
    .B(_0149_));
 sg13g2_nor2_1 _4025_ (.A(_2417_),
    .B(_0150_),
    .Y(_0151_));
 sg13g2_nand2_1 _4026_ (.Y(_0152_),
    .A(_0151_),
    .B(net215));
 sg13g2_inv_2 _4027_ (.Y(_0153_),
    .A(_2397_));
 sg13g2_nor2_1 _4028_ (.A(_0153_),
    .B(_2911_),
    .Y(_0154_));
 sg13g2_o21ai_1 _4029_ (.B1(_2639_),
    .Y(_0155_),
    .A1(_0152_),
    .A2(_0154_));
 sg13g2_a21oi_1 _4030_ (.A1(_0148_),
    .A2(_2632_),
    .Y(_0156_),
    .B1(_0155_));
 sg13g2_nand2_1 _4031_ (.Y(_0157_),
    .A(_0132_),
    .B(_0156_));
 sg13g2_a21oi_1 _4032_ (.A1(_0106_),
    .A2(net194),
    .Y(_0158_),
    .B1(_0157_));
 sg13g2_nor2_1 _4033_ (.A(_3013_),
    .B(_0158_),
    .Y(_0021_));
 sg13g2_nand2_1 _4034_ (.Y(_0159_),
    .A(_2584_),
    .B(_2776_));
 sg13g2_nand3_1 _4035_ (.B(net126),
    .C(_2787_),
    .A(_0159_),
    .Y(_0160_));
 sg13g2_nand2_1 _4036_ (.Y(_0161_),
    .A(_2736_),
    .B(_1599_));
 sg13g2_nand2_1 _4037_ (.Y(_0162_),
    .A(_0161_),
    .B(_2782_));
 sg13g2_nand2_1 _4038_ (.Y(_0163_),
    .A(_0160_),
    .B(_0162_));
 sg13g2_nand2_1 _4039_ (.Y(_0164_),
    .A(_2784_),
    .B(_2289_));
 sg13g2_nor2_1 _4040_ (.A(net180),
    .B(_0164_),
    .Y(_0165_));
 sg13g2_nor2b_1 _4041_ (.A(_0165_),
    .B_N(_2444_),
    .Y(_0166_));
 sg13g2_nor3_1 _4042_ (.A(_1981_),
    .B(net67),
    .C(_0166_),
    .Y(_0167_));
 sg13g2_nand2_1 _4043_ (.Y(_0168_),
    .A(_3031_),
    .B(net61));
 sg13g2_nand2_1 _4044_ (.Y(_0169_),
    .A(net83),
    .B(_2703_));
 sg13g2_and3_1 _4045_ (.X(_0170_),
    .A(_0168_),
    .B(_0169_),
    .C(net91));
 sg13g2_nor3_1 _4046_ (.A(_2405_),
    .B(_3027_),
    .C(_0170_),
    .Y(_0171_));
 sg13g2_nor3_1 _4047_ (.A(_0163_),
    .B(_0167_),
    .C(_0171_),
    .Y(_0172_));
 sg13g2_inv_1 _4048_ (.Y(_0173_),
    .A(_2669_));
 sg13g2_nand2_1 _4049_ (.Y(_0174_),
    .A(_0900_),
    .B(_0878_));
 sg13g2_buf_2 _4050_ (.A(_0174_),
    .X(_0175_));
 sg13g2_nor2_1 _4051_ (.A(_0175_),
    .B(net78),
    .Y(_0176_));
 sg13g2_inv_1 _4052_ (.Y(_0177_),
    .A(_0176_));
 sg13g2_nand2_1 _4053_ (.Y(_0178_),
    .A(_0177_),
    .B(_2976_));
 sg13g2_a22oi_1 _4054_ (.Y(_0179_),
    .B1(net127),
    .B2(_0178_),
    .A2(net102),
    .A1(_0173_));
 sg13g2_a21oi_2 _4055_ (.B1(_2066_),
    .Y(_0180_),
    .A2(net94),
    .A1(_2137_));
 sg13g2_o21ai_1 _4056_ (.B1(_2771_),
    .Y(_0181_),
    .A1(_0180_),
    .A2(_0165_));
 sg13g2_inv_1 _4057_ (.Y(_0182_),
    .A(_2868_));
 sg13g2_nand3_1 _4058_ (.B(_2206_),
    .C(_0182_),
    .A(_2507_),
    .Y(_0183_));
 sg13g2_nand2_1 _4059_ (.Y(_0184_),
    .A(_2720_),
    .B(net78));
 sg13g2_nand2_1 _4060_ (.Y(_0185_),
    .A(_0183_),
    .B(_0184_));
 sg13g2_nand2_1 _4061_ (.Y(_0186_),
    .A(_0185_),
    .B(net122));
 sg13g2_nand3_1 _4062_ (.B(_0181_),
    .C(_0186_),
    .A(_0179_),
    .Y(_0187_));
 sg13g2_nand2_1 _4063_ (.Y(_0188_),
    .A(_0187_),
    .B(net125));
 sg13g2_nand2_1 _4064_ (.Y(_0189_),
    .A(_0172_),
    .B(_0188_));
 sg13g2_nand2_1 _4065_ (.Y(_0190_),
    .A(_0189_),
    .B(net151));
 sg13g2_buf_1 _4066_ (.A(net69),
    .X(_0191_));
 sg13g2_nor2_1 _4067_ (.A(_2496_),
    .B(_2964_),
    .Y(_0192_));
 sg13g2_o21ai_1 _4068_ (.B1(_2725_),
    .Y(_0193_),
    .A1(net39),
    .A2(_0192_));
 sg13g2_buf_1 _4069_ (.A(net191),
    .X(_0194_));
 sg13g2_nor2_1 _4070_ (.A(_2488_),
    .B(_2400_),
    .Y(_0195_));
 sg13g2_inv_1 _4071_ (.Y(_0196_),
    .A(_0195_));
 sg13g2_buf_2 _4072_ (.A(net163),
    .X(_0197_));
 sg13g2_nand2_1 _4073_ (.Y(_0198_),
    .A(_2621_),
    .B(net169));
 sg13g2_nand3_1 _4074_ (.B(net89),
    .C(_0198_),
    .A(_0196_),
    .Y(_0199_));
 sg13g2_nand3_1 _4075_ (.B(net135),
    .C(_0199_),
    .A(_0193_),
    .Y(_0200_));
 sg13g2_nand2_1 _4076_ (.Y(_0201_),
    .A(_2577_),
    .B(_2602_));
 sg13g2_nand2_1 _4077_ (.Y(_0202_),
    .A(_0201_),
    .B(_2488_));
 sg13g2_nor2_1 _4078_ (.A(_2525_),
    .B(_2720_),
    .Y(_0203_));
 sg13g2_inv_1 _4079_ (.Y(_0204_),
    .A(_2485_));
 sg13g2_nand2_1 _4080_ (.Y(_0205_),
    .A(_0204_),
    .B(net71));
 sg13g2_a22oi_1 _4081_ (.Y(_0206_),
    .B1(_0203_),
    .B2(_0205_),
    .A2(_0202_),
    .A1(net53));
 sg13g2_nand2_1 _4082_ (.Y(_0207_),
    .A(_0200_),
    .B(_0206_));
 sg13g2_inv_1 _4083_ (.Y(_0208_),
    .A(_1064_));
 sg13g2_o21ai_1 _4084_ (.B1(net74),
    .Y(_0209_),
    .A1(_2968_),
    .A2(_0208_));
 sg13g2_nand2_1 _4085_ (.Y(_0210_),
    .A(_2666_),
    .B(_2117_));
 sg13g2_buf_2 _4086_ (.A(_0210_),
    .X(_0211_));
 sg13g2_a21oi_1 _4087_ (.A1(_0209_),
    .A2(_0211_),
    .Y(_0212_),
    .B1(_0152_));
 sg13g2_nand2b_1 _4088_ (.Y(_0213_),
    .B(_2639_),
    .A_N(_0212_));
 sg13g2_a21oi_1 _4089_ (.A1(_0207_),
    .A2(_2632_),
    .Y(_0214_),
    .B1(_0213_));
 sg13g2_nand2_1 _4090_ (.Y(_0215_),
    .A(_0190_),
    .B(_0214_));
 sg13g2_inv_2 _4091_ (.Y(_0216_),
    .A(_2557_));
 sg13g2_nand3_1 _4092_ (.B(net122),
    .C(_0216_),
    .A(net44),
    .Y(_0217_));
 sg13g2_nor2_1 _4093_ (.A(net129),
    .B(_2755_),
    .Y(_0218_));
 sg13g2_nand2_1 _4094_ (.Y(_0219_),
    .A(_0218_),
    .B(net157));
 sg13g2_nand2_1 _4095_ (.Y(_0220_),
    .A(_2381_),
    .B(net142));
 sg13g2_a21oi_1 _4096_ (.A1(_2898_),
    .A2(_2733_),
    .Y(_0221_),
    .B1(_1970_));
 sg13g2_nand4_1 _4097_ (.B(_0219_),
    .C(_0220_),
    .A(_0217_),
    .Y(_0222_),
    .D(_0221_));
 sg13g2_nand2_1 _4098_ (.Y(_0223_),
    .A(_0222_),
    .B(_2405_));
 sg13g2_nand2_1 _4099_ (.Y(_0224_),
    .A(_3049_),
    .B(_2462_));
 sg13g2_nand3_1 _4100_ (.B(net92),
    .C(_0224_),
    .A(_2969_),
    .Y(_0225_));
 sg13g2_nand3_1 _4101_ (.B(net89),
    .C(_2445_),
    .A(_2873_),
    .Y(_0226_));
 sg13g2_nand3_1 _4102_ (.B(_0141_),
    .C(_0226_),
    .A(_0225_),
    .Y(_0227_));
 sg13g2_nand2_1 _4103_ (.Y(_0228_),
    .A(_0223_),
    .B(_0227_));
 sg13g2_nor2_1 _4104_ (.A(_0175_),
    .B(_2507_),
    .Y(_0229_));
 sg13g2_nor2_1 _4105_ (.A(net112),
    .B(_0229_),
    .Y(_0230_));
 sg13g2_nor2_1 _4106_ (.A(net221),
    .B(_0845_),
    .Y(_0231_));
 sg13g2_inv_1 _4107_ (.Y(_0232_),
    .A(_0231_));
 sg13g2_nand2_2 _4108_ (.Y(_0233_),
    .A(_0232_),
    .B(net42));
 sg13g2_inv_1 _4109_ (.Y(_0234_),
    .A(_2533_));
 sg13g2_nand2_2 _4110_ (.Y(_0235_),
    .A(_0234_),
    .B(net108));
 sg13g2_o21ai_1 _4111_ (.B1(_0235_),
    .Y(_0236_),
    .A1(net147),
    .A2(_1392_));
 sg13g2_a22oi_1 _4112_ (.Y(_0237_),
    .B1(net40),
    .B2(_0236_),
    .A2(_0233_),
    .A1(_0230_));
 sg13g2_nand2_1 _4113_ (.Y(_0238_),
    .A(net44),
    .B(net94));
 sg13g2_nand2_1 _4114_ (.Y(_0239_),
    .A(_0238_),
    .B(net69));
 sg13g2_a21oi_1 _4115_ (.A1(_3049_),
    .A2(net57),
    .Y(_0240_),
    .B1(net119));
 sg13g2_nand2_1 _4116_ (.Y(_0241_),
    .A(_0239_),
    .B(_0240_));
 sg13g2_nand2_1 _4117_ (.Y(_0242_),
    .A(_2555_),
    .B(_2384_));
 sg13g2_nor2_1 _4118_ (.A(_0136_),
    .B(_0911_),
    .Y(_0243_));
 sg13g2_a21oi_1 _4119_ (.A1(_0242_),
    .A2(_0243_),
    .Y(_0244_),
    .B1(net144));
 sg13g2_nand2_1 _4120_ (.Y(_0245_),
    .A(_0241_),
    .B(_0244_));
 sg13g2_nand3_1 _4121_ (.B(net125),
    .C(_0245_),
    .A(_0237_),
    .Y(_0246_));
 sg13g2_nand3_1 _4122_ (.B(_0246_),
    .C(net138),
    .A(_0228_),
    .Y(_0247_));
 sg13g2_nand2_2 _4123_ (.Y(_0248_),
    .A(_0900_),
    .B(net160));
 sg13g2_inv_1 _4124_ (.Y(_0249_),
    .A(_0248_));
 sg13g2_nand2_1 _4125_ (.Y(_0250_),
    .A(_0249_),
    .B(_2733_));
 sg13g2_nand2_1 _4126_ (.Y(_0251_),
    .A(_0250_),
    .B(net217));
 sg13g2_nor2_1 _4127_ (.A(net91),
    .B(_2873_),
    .Y(_0252_));
 sg13g2_nor2_1 _4128_ (.A(_0251_),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_nand2_1 _4129_ (.Y(_0254_),
    .A(_0180_),
    .B(net91));
 sg13g2_a21oi_1 _4130_ (.A1(_0253_),
    .A2(_0254_),
    .Y(_0255_),
    .B1(net171));
 sg13g2_inv_1 _4131_ (.Y(_0256_),
    .A(_0944_));
 sg13g2_o21ai_1 _4132_ (.B1(net139),
    .Y(_0257_),
    .A1(net201),
    .A2(net64));
 sg13g2_nor2_1 _4133_ (.A(net142),
    .B(_2974_),
    .Y(_0258_));
 sg13g2_nand2_1 _4134_ (.Y(_0259_),
    .A(_2986_),
    .B(net59));
 sg13g2_buf_1 _4135_ (.A(net196),
    .X(_0260_));
 sg13g2_a21oi_1 _4136_ (.A1(_0258_),
    .A2(_0259_),
    .Y(_0261_),
    .B1(net134));
 sg13g2_o21ai_1 _4137_ (.B1(_0261_),
    .Y(_0262_),
    .A1(_0256_),
    .A2(_0257_));
 sg13g2_nand2b_1 _4138_ (.Y(_0263_),
    .B(_0262_),
    .A_N(_0255_));
 sg13g2_nand2_1 _4139_ (.Y(_0264_),
    .A(_2756_),
    .B(_2395_));
 sg13g2_nand2_1 _4140_ (.Y(_0265_),
    .A(_3001_),
    .B(_2472_));
 sg13g2_nand2_1 _4141_ (.Y(_0266_),
    .A(_0264_),
    .B(_0265_));
 sg13g2_nand2_1 _4142_ (.Y(_0267_),
    .A(_2434_),
    .B(_2805_));
 sg13g2_o21ai_1 _4143_ (.B1(_2976_),
    .Y(_0268_),
    .A1(_2475_),
    .A2(_0267_));
 sg13g2_a22oi_1 _4144_ (.Y(_0269_),
    .B1(net53),
    .B2(_0268_),
    .A2(net98),
    .A1(_0266_));
 sg13g2_nand2b_1 _4145_ (.Y(_0270_),
    .B(net40),
    .A_N(_0166_));
 sg13g2_nor2_1 _4146_ (.A(net60),
    .B(_0108_),
    .Y(_0271_));
 sg13g2_buf_1 _4147_ (.A(net214),
    .X(_0272_));
 sg13g2_a21oi_1 _4148_ (.A1(_0271_),
    .A2(_2524_),
    .Y(_0273_),
    .B1(net184));
 sg13g2_nand3_1 _4149_ (.B(_0270_),
    .C(_0273_),
    .A(_0269_),
    .Y(_0274_));
 sg13g2_nand3_1 _4150_ (.B(_0274_),
    .C(net143),
    .A(_0263_),
    .Y(_0275_));
 sg13g2_a21oi_1 _4151_ (.A1(_0247_),
    .A2(_0275_),
    .Y(_0276_),
    .B1(_2751_));
 sg13g2_nor2_1 _4152_ (.A(_0215_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_nand2_1 _4153_ (.Y(_0278_),
    .A(_2482_),
    .B(_2137_));
 sg13g2_nand2_1 _4154_ (.Y(_0279_),
    .A(_0278_),
    .B(net59));
 sg13g2_nand2_1 _4155_ (.Y(_0280_),
    .A(net46),
    .B(_2666_));
 sg13g2_inv_1 _4156_ (.Y(_0281_),
    .A(_0280_));
 sg13g2_nor2_1 _4157_ (.A(net142),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_buf_2 _4158_ (.A(net97),
    .X(_0283_));
 sg13g2_a21oi_1 _4159_ (.A1(_0279_),
    .A2(_0282_),
    .Y(_0284_),
    .B1(net50));
 sg13g2_nor2_2 _4160_ (.A(net202),
    .B(_2855_),
    .Y(_0285_));
 sg13g2_nand2_1 _4161_ (.Y(_0286_),
    .A(_0285_),
    .B(_0196_));
 sg13g2_nand2_1 _4162_ (.Y(_0287_),
    .A(_0284_),
    .B(_0286_));
 sg13g2_nor2_1 _4163_ (.A(net43),
    .B(_2744_),
    .Y(_0288_));
 sg13g2_a21oi_1 _4164_ (.A1(_2704_),
    .A2(_0922_),
    .Y(_0289_),
    .B1(net67));
 sg13g2_nor2_1 _4165_ (.A(_0288_),
    .B(_0289_),
    .Y(_0290_));
 sg13g2_a21oi_1 _4166_ (.A1(_0287_),
    .A2(_0290_),
    .Y(_0291_),
    .B1(net165));
 sg13g2_nor2_1 _4167_ (.A(_2250_),
    .B(_0192_),
    .Y(_0292_));
 sg13g2_nand2_1 _4168_ (.Y(_0293_),
    .A(_2504_),
    .B(_2370_));
 sg13g2_o21ai_1 _4169_ (.B1(net120),
    .Y(_0294_),
    .A1(_2968_),
    .A2(_2461_));
 sg13g2_nand3_1 _4170_ (.B(_2830_),
    .C(net175),
    .A(net121),
    .Y(_0295_));
 sg13g2_nand3_1 _4171_ (.B(_0294_),
    .C(_0295_),
    .A(_0293_),
    .Y(_0296_));
 sg13g2_buf_1 _4172_ (.A(net109),
    .X(_0297_));
 sg13g2_o21ai_1 _4173_ (.B1(net49),
    .Y(_0298_),
    .A1(_0292_),
    .A2(_0296_));
 sg13g2_inv_1 _4174_ (.Y(_0299_),
    .A(_2856_));
 sg13g2_nor2_2 _4175_ (.A(net220),
    .B(_0299_),
    .Y(_0300_));
 sg13g2_inv_1 _4176_ (.Y(_0301_),
    .A(_0300_));
 sg13g2_nor3_1 _4177_ (.A(_2403_),
    .B(_0301_),
    .C(_2855_),
    .Y(_0302_));
 sg13g2_nor2_1 _4178_ (.A(net110),
    .B(_0302_),
    .Y(_0303_));
 sg13g2_buf_1 _4179_ (.A(net142),
    .X(_0304_));
 sg13g2_nand3_1 _4180_ (.B(net88),
    .C(_2671_),
    .A(_2760_),
    .Y(_0305_));
 sg13g2_nand2_1 _4181_ (.Y(_0306_),
    .A(_0303_),
    .B(_0305_));
 sg13g2_nand2_1 _4182_ (.Y(_0307_),
    .A(_0298_),
    .B(_0306_));
 sg13g2_buf_1 _4183_ (.A(net140),
    .X(_0308_));
 sg13g2_nand2_1 _4184_ (.Y(_0309_),
    .A(_0307_),
    .B(net87));
 sg13g2_nand2_2 _4185_ (.Y(_0310_),
    .A(_2615_),
    .B(_2736_));
 sg13g2_nand2_1 _4186_ (.Y(_0311_),
    .A(_0310_),
    .B(net72));
 sg13g2_nand2_1 _4187_ (.Y(_0312_),
    .A(_2482_),
    .B(net61));
 sg13g2_nand3_1 _4188_ (.B(_0312_),
    .C(net92),
    .A(_0311_),
    .Y(_0313_));
 sg13g2_inv_1 _4189_ (.Y(_0314_),
    .A(_0867_));
 sg13g2_a21oi_1 _4190_ (.A1(_0314_),
    .A2(_2668_),
    .Y(_0315_),
    .B1(net109));
 sg13g2_nand2_1 _4191_ (.Y(_0316_),
    .A(_0313_),
    .B(_0315_));
 sg13g2_a21oi_1 _4192_ (.A1(_1413_),
    .A2(_2380_),
    .Y(_0317_),
    .B1(_2701_));
 sg13g2_inv_1 _4193_ (.Y(_0318_),
    .A(_0175_));
 sg13g2_nor3_1 _4194_ (.A(net80),
    .B(_0318_),
    .C(_0195_),
    .Y(_0319_));
 sg13g2_nor3_1 _4195_ (.A(net145),
    .B(_0317_),
    .C(_0319_),
    .Y(_0320_));
 sg13g2_a21oi_1 _4196_ (.A1(_0316_),
    .A2(_0320_),
    .Y(_0321_),
    .B1(net187));
 sg13g2_nand2_1 _4197_ (.Y(_0322_),
    .A(_0285_),
    .B(_2617_));
 sg13g2_a21oi_1 _4198_ (.A1(_0111_),
    .A2(_0198_),
    .Y(_0323_),
    .B1(net144));
 sg13g2_a21oi_1 _4199_ (.A1(_0322_),
    .A2(_0323_),
    .Y(_0324_),
    .B1(net141));
 sg13g2_nor2_1 _4200_ (.A(net189),
    .B(_2900_),
    .Y(_0325_));
 sg13g2_nand2_1 _4201_ (.Y(_0326_),
    .A(net83),
    .B(net104));
 sg13g2_nand2_1 _4202_ (.Y(_0327_),
    .A(_0326_),
    .B(net72));
 sg13g2_a21oi_1 _4203_ (.A1(_0325_),
    .A2(_0327_),
    .Y(_0328_),
    .B1(net110));
 sg13g2_nand2_1 _4204_ (.Y(_0329_),
    .A(net79),
    .B(_2453_));
 sg13g2_nand2_1 _4205_ (.Y(_0330_),
    .A(_2932_),
    .B(_0329_));
 sg13g2_nand2_2 _4206_ (.Y(_0331_),
    .A(_0330_),
    .B(net118));
 sg13g2_nand2_1 _4207_ (.Y(_0332_),
    .A(_0331_),
    .B(_2824_));
 sg13g2_nand2_1 _4208_ (.Y(_0333_),
    .A(_0328_),
    .B(_0332_));
 sg13g2_nand2_1 _4209_ (.Y(_0334_),
    .A(_0324_),
    .B(_0333_));
 sg13g2_nand2_1 _4210_ (.Y(_0335_),
    .A(_0321_),
    .B(_0334_));
 sg13g2_nand3b_1 _4211_ (.B(_0309_),
    .C(_0335_),
    .Y(_0336_),
    .A_N(_0291_));
 sg13g2_nor2_1 _4212_ (.A(net101),
    .B(_2616_),
    .Y(_0337_));
 sg13g2_nand2_2 _4213_ (.Y(_0338_),
    .A(net73),
    .B(_2599_));
 sg13g2_nor2_1 _4214_ (.A(net148),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_a21oi_1 _4215_ (.A1(_0339_),
    .A2(_1119_),
    .Y(_0340_),
    .B1(net97));
 sg13g2_o21ai_1 _4216_ (.B1(_0340_),
    .Y(_0341_),
    .A1(_3054_),
    .A2(_0337_));
 sg13g2_nand2_1 _4217_ (.Y(_0342_),
    .A(net79),
    .B(_2700_));
 sg13g2_nand2_1 _4218_ (.Y(_0343_),
    .A(_0342_),
    .B(_0211_));
 sg13g2_inv_1 _4219_ (.Y(_0344_),
    .A(_2206_));
 sg13g2_nand2_2 _4220_ (.Y(_0345_),
    .A(_2215_),
    .B(net162));
 sg13g2_nand2_1 _4221_ (.Y(_0346_),
    .A(net96),
    .B(net178));
 sg13g2_o21ai_1 _4222_ (.B1(_0346_),
    .Y(_0347_),
    .A1(_0344_),
    .A2(_0345_));
 sg13g2_a22oi_1 _4223_ (.Y(_0348_),
    .B1(net90),
    .B2(_0347_),
    .A2(net54),
    .A1(_0343_));
 sg13g2_nand2_1 _4224_ (.Y(_0349_),
    .A(_0341_),
    .B(_0348_));
 sg13g2_inv_1 _4225_ (.Y(_0350_),
    .A(_2417_));
 sg13g2_buf_1 _4226_ (.A(_0350_),
    .X(_0351_));
 sg13g2_nand2_1 _4227_ (.Y(_0352_),
    .A(_0349_),
    .B(net86));
 sg13g2_nand2_2 _4228_ (.Y(_0353_),
    .A(net81),
    .B(net107));
 sg13g2_a22oi_1 _4229_ (.Y(_0354_),
    .B1(net65),
    .B2(_0353_),
    .A2(net103),
    .A1(net70));
 sg13g2_nand2_1 _4230_ (.Y(_0355_),
    .A(_2950_),
    .B(net96));
 sg13g2_nand3_1 _4231_ (.B(net137),
    .C(_0355_),
    .A(_3050_),
    .Y(_0356_));
 sg13g2_nand2_1 _4232_ (.Y(_0357_),
    .A(_0356_),
    .B(net146));
 sg13g2_o21ai_1 _4233_ (.B1(_0357_),
    .Y(_0358_),
    .A1(net110),
    .A2(_0354_));
 sg13g2_nand3_1 _4234_ (.B(net97),
    .C(_1675_),
    .A(_2614_),
    .Y(_0359_));
 sg13g2_nand3_1 _4235_ (.B(net185),
    .C(_2648_),
    .A(net64),
    .Y(_0360_));
 sg13g2_nand2_1 _4236_ (.Y(_0361_),
    .A(_1577_),
    .B(_2389_));
 sg13g2_a21oi_1 _4237_ (.A1(_0361_),
    .A2(net72),
    .Y(_0362_),
    .B1(_2501_));
 sg13g2_nand3_1 _4238_ (.B(_0360_),
    .C(_0362_),
    .A(_0359_),
    .Y(_0363_));
 sg13g2_nand3_1 _4239_ (.B(net140),
    .C(_0363_),
    .A(_0358_),
    .Y(_0364_));
 sg13g2_nand2_1 _4240_ (.Y(_0365_),
    .A(_0352_),
    .B(_0364_));
 sg13g2_nand2_1 _4241_ (.Y(_0366_),
    .A(_0365_),
    .B(net190));
 sg13g2_nand2_1 _4242_ (.Y(_0367_),
    .A(_2137_),
    .B(_1708_));
 sg13g2_inv_1 _4243_ (.Y(_0368_),
    .A(_0367_));
 sg13g2_a21oi_1 _4244_ (.A1(_0368_),
    .A2(_2784_),
    .Y(_0369_),
    .B1(net158));
 sg13g2_nor2_1 _4245_ (.A(net164),
    .B(_0216_),
    .Y(_0370_));
 sg13g2_nand2_1 _4246_ (.Y(_0371_),
    .A(_0369_),
    .B(_0370_));
 sg13g2_nor3_1 _4247_ (.A(_2525_),
    .B(_2612_),
    .C(_2963_),
    .Y(_0372_));
 sg13g2_nand2_1 _4248_ (.Y(_0373_),
    .A(_2434_),
    .B(_1697_));
 sg13g2_nor2_1 _4249_ (.A(_0976_),
    .B(_0373_),
    .Y(_0374_));
 sg13g2_nand2_1 _4250_ (.Y(_0375_),
    .A(_0374_),
    .B(_1785_));
 sg13g2_nand2_1 _4251_ (.Y(_0376_),
    .A(_0375_),
    .B(net217));
 sg13g2_nor2_1 _4252_ (.A(_0372_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_nand2_1 _4253_ (.Y(_0378_),
    .A(_0371_),
    .B(_0377_));
 sg13g2_nand3_1 _4254_ (.B(_2895_),
    .C(net102),
    .A(_2473_),
    .Y(_0379_));
 sg13g2_o21ai_1 _4255_ (.B1(_2915_),
    .Y(_0380_),
    .A1(_2538_),
    .A2(_2536_));
 sg13g2_buf_2 _4256_ (.A(_2447_),
    .X(_0381_));
 sg13g2_nand2_1 _4257_ (.Y(_0382_),
    .A(_0380_),
    .B(net85));
 sg13g2_nand2_1 _4258_ (.Y(_0383_),
    .A(_0379_),
    .B(_0382_));
 sg13g2_nor2_1 _4259_ (.A(_0378_),
    .B(_0383_),
    .Y(_0384_));
 sg13g2_nor2_1 _4260_ (.A(_2949_),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_nor2_1 _4261_ (.A(_3051_),
    .B(_2938_),
    .Y(_0386_));
 sg13g2_nor2_1 _4262_ (.A(_2267_),
    .B(_2905_),
    .Y(_0387_));
 sg13g2_nand2_1 _4263_ (.Y(_0388_),
    .A(_2137_),
    .B(net94));
 sg13g2_o21ai_1 _4264_ (.B1(net185),
    .Y(_0389_),
    .A1(_2250_),
    .A2(_0388_));
 sg13g2_nor3_1 _4265_ (.A(_0386_),
    .B(_0387_),
    .C(_0389_),
    .Y(_0390_));
 sg13g2_a22oi_1 _4266_ (.Y(_0391_),
    .B1(net157),
    .B2(_0176_),
    .A2(_2426_),
    .A1(_2829_));
 sg13g2_a21oi_1 _4267_ (.A1(_0391_),
    .A2(_0254_),
    .Y(_0392_),
    .B1(net152));
 sg13g2_nor2_1 _4268_ (.A(_0390_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_nand2_1 _4269_ (.Y(_0394_),
    .A(_0393_),
    .B(_2947_));
 sg13g2_a21oi_1 _4270_ (.A1(_0385_),
    .A2(_0394_),
    .Y(_0395_),
    .B1(_2639_));
 sg13g2_nand2_1 _4271_ (.Y(_0396_),
    .A(_0366_),
    .B(_0395_));
 sg13g2_a21oi_1 _4272_ (.A1(_0336_),
    .A2(net194),
    .Y(_0397_),
    .B1(_0396_));
 sg13g2_nor2_1 _4273_ (.A(_0277_),
    .B(_0397_),
    .Y(_0022_));
 sg13g2_a21oi_1 _4274_ (.A1(net41),
    .A2(net130),
    .Y(_0398_),
    .B1(_2117_));
 sg13g2_nand3_1 _4275_ (.B(_2658_),
    .C(_2766_),
    .A(_2913_),
    .Y(_0399_));
 sg13g2_o21ai_1 _4276_ (.B1(_0399_),
    .Y(_0400_),
    .A1(net179),
    .A2(_0398_));
 sg13g2_o21ai_1 _4277_ (.B1(net214),
    .Y(_0401_),
    .A1(_2525_),
    .A2(_0097_));
 sg13g2_nor2_1 _4278_ (.A(_0400_),
    .B(_0401_),
    .Y(_0402_));
 sg13g2_nand2_1 _4279_ (.Y(_0403_),
    .A(_0279_),
    .B(_2541_));
 sg13g2_nand2_1 _4280_ (.Y(_0404_),
    .A(_0403_),
    .B(net98));
 sg13g2_a21oi_1 _4281_ (.A1(_0402_),
    .A2(_0404_),
    .Y(_0405_),
    .B1(net199));
 sg13g2_nand2_1 _4282_ (.Y(_0406_),
    .A(net65),
    .B(net82));
 sg13g2_nor2_1 _4283_ (.A(net117),
    .B(_3034_),
    .Y(_0407_));
 sg13g2_a21oi_1 _4284_ (.A1(_0406_),
    .A2(_0407_),
    .Y(_0408_),
    .B1(net179));
 sg13g2_a21oi_1 _4285_ (.A1(_2876_),
    .A2(_0198_),
    .Y(_0409_),
    .B1(net128));
 sg13g2_nor3_1 _4286_ (.A(net192),
    .B(_0408_),
    .C(_0409_),
    .Y(_0410_));
 sg13g2_inv_1 _4287_ (.Y(_0411_),
    .A(_0312_));
 sg13g2_o21ai_1 _4288_ (.B1(_2983_),
    .Y(_0412_),
    .A1(_0411_),
    .A2(_2572_));
 sg13g2_nor2_1 _4289_ (.A(_0134_),
    .B(_0161_),
    .Y(_0413_));
 sg13g2_nor2_1 _4290_ (.A(net123),
    .B(_2571_),
    .Y(_0414_));
 sg13g2_o21ai_1 _4291_ (.B1(net85),
    .Y(_0415_),
    .A1(_0413_),
    .A2(_0414_));
 sg13g2_nand3_1 _4292_ (.B(_0412_),
    .C(_0415_),
    .A(_0410_),
    .Y(_0416_));
 sg13g2_nand2_1 _4293_ (.Y(_0417_),
    .A(_0405_),
    .B(_0416_));
 sg13g2_nand2_1 _4294_ (.Y(_0418_),
    .A(_2768_),
    .B(_2318_));
 sg13g2_nand2_1 _4295_ (.Y(_0419_),
    .A(_0418_),
    .B(net130));
 sg13g2_a21oi_1 _4296_ (.A1(_0419_),
    .A2(_1413_),
    .Y(_0420_),
    .B1(_2525_));
 sg13g2_a21oi_1 _4297_ (.A1(_0216_),
    .A2(_1621_),
    .Y(_0421_),
    .B1(_1446_));
 sg13g2_nand2_2 _4298_ (.Y(_0422_),
    .A(_3032_),
    .B(net123));
 sg13g2_nand2_1 _4299_ (.Y(_0423_),
    .A(_0421_),
    .B(_0422_));
 sg13g2_nand2_1 _4300_ (.Y(_0424_),
    .A(_0423_),
    .B(net214));
 sg13g2_nor2_1 _4301_ (.A(_0420_),
    .B(_0424_),
    .Y(_0425_));
 sg13g2_inv_1 _4302_ (.Y(_0426_),
    .A(_2670_));
 sg13g2_nor2_1 _4303_ (.A(net70),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_o21ai_1 _4304_ (.B1(net196),
    .Y(_0428_),
    .A1(_2399_),
    .A2(_0427_));
 sg13g2_nand2_2 _4305_ (.Y(_0429_),
    .A(_2533_),
    .B(_2691_));
 sg13g2_nand2_1 _4306_ (.Y(_0430_),
    .A(_0429_),
    .B(net108));
 sg13g2_nand3_1 _4307_ (.B(net95),
    .C(net201),
    .A(_0430_),
    .Y(_0431_));
 sg13g2_nand2b_1 _4308_ (.Y(_0432_),
    .B(_0431_),
    .A_N(_0428_));
 sg13g2_a21oi_1 _4309_ (.A1(_0425_),
    .A2(_0432_),
    .Y(_0433_),
    .B1(net187));
 sg13g2_nand2b_1 _4310_ (.Y(_0434_),
    .B(_0369_),
    .A_N(_2558_));
 sg13g2_a21oi_2 _4311_ (.B1(_1697_),
    .Y(_0435_),
    .A2(net224),
    .A1(_1643_));
 sg13g2_nand3_1 _4312_ (.B(_2137_),
    .C(_2784_),
    .A(_0435_),
    .Y(_0436_));
 sg13g2_buf_2 _4313_ (.A(_0436_),
    .X(_0437_));
 sg13g2_nand3_1 _4314_ (.B(net91),
    .C(_2777_),
    .A(_0437_),
    .Y(_0438_));
 sg13g2_nand3_1 _4315_ (.B(_0438_),
    .C(net144),
    .A(_0434_),
    .Y(_0439_));
 sg13g2_inv_1 _4316_ (.Y(_0440_),
    .A(_2731_));
 sg13g2_nand2_1 _4317_ (.Y(_0441_),
    .A(_0440_),
    .B(_0108_));
 sg13g2_nand2_1 _4318_ (.Y(_0442_),
    .A(_2622_),
    .B(net113));
 sg13g2_nand3_1 _4319_ (.B(_0442_),
    .C(net149),
    .A(_0441_),
    .Y(_0443_));
 sg13g2_nand2_1 _4320_ (.Y(_0444_),
    .A(_0443_),
    .B(net203));
 sg13g2_nand3_1 _4321_ (.B(net114),
    .C(_2664_),
    .A(_2623_),
    .Y(_0445_));
 sg13g2_nor2b_1 _4322_ (.A(_0444_),
    .B_N(_0445_),
    .Y(_0446_));
 sg13g2_nand2_1 _4323_ (.Y(_0447_),
    .A(_0439_),
    .B(_0446_));
 sg13g2_nand2_1 _4324_ (.Y(_0448_),
    .A(_0433_),
    .B(_0447_));
 sg13g2_nand2_1 _4325_ (.Y(_0449_),
    .A(_0417_),
    .B(_0448_));
 sg13g2_nand2_1 _4326_ (.Y(_0450_),
    .A(_0449_),
    .B(net194));
 sg13g2_nand2_1 _4327_ (.Y(_0451_),
    .A(_2720_),
    .B(_0353_));
 sg13g2_nand3_1 _4328_ (.B(_0451_),
    .C(net142),
    .A(_1861_),
    .Y(_0452_));
 sg13g2_nor2b_1 _4329_ (.A(net110),
    .B_N(_0452_),
    .Y(_0453_));
 sg13g2_nand2_1 _4330_ (.Y(_0454_),
    .A(_2616_),
    .B(net118));
 sg13g2_buf_1 _4331_ (.A(net95),
    .X(_0455_));
 sg13g2_nand3_1 _4332_ (.B(net48),
    .C(_0422_),
    .A(_0454_),
    .Y(_0456_));
 sg13g2_a21oi_1 _4333_ (.A1(_0453_),
    .A2(_0456_),
    .Y(_0457_),
    .B1(net150));
 sg13g2_nand2_1 _4334_ (.Y(_0458_),
    .A(_2812_),
    .B(_2506_));
 sg13g2_nand2_1 _4335_ (.Y(_0459_),
    .A(_0458_),
    .B(net189));
 sg13g2_a21oi_2 _4336_ (.B1(_1512_),
    .Y(_0460_),
    .A2(net221),
    .A1(net170));
 sg13g2_nand2_2 _4337_ (.Y(_0461_),
    .A(_0460_),
    .B(net74));
 sg13g2_a21oi_1 _4338_ (.A1(_0461_),
    .A2(_2436_),
    .Y(_0462_),
    .B1(net152));
 sg13g2_o21ai_1 _4339_ (.B1(_0462_),
    .Y(_0463_),
    .A1(_2572_),
    .A2(_0459_));
 sg13g2_nor2_1 _4340_ (.A(_0867_),
    .B(_2572_),
    .Y(_0464_));
 sg13g2_o21ai_1 _4341_ (.B1(net184),
    .Y(_0465_),
    .A1(_0150_),
    .A2(_0464_));
 sg13g2_nand2_1 _4342_ (.Y(_0466_),
    .A(_0465_),
    .B(_2848_));
 sg13g2_a21oi_1 _4343_ (.A1(_0457_),
    .A2(_0463_),
    .Y(_0467_),
    .B1(_0466_));
 sg13g2_a21oi_1 _4344_ (.A1(_2569_),
    .A2(net107),
    .Y(_0468_),
    .B1(net69));
 sg13g2_o21ai_1 _4345_ (.B1(_0118_),
    .Y(_0469_),
    .A1(_0468_),
    .A2(_2934_));
 sg13g2_o21ai_1 _4346_ (.B1(net85),
    .Y(_0470_),
    .A1(_2577_),
    .A2(_2934_));
 sg13g2_nand2_1 _4347_ (.Y(_0471_),
    .A(_0469_),
    .B(_0470_));
 sg13g2_a21oi_1 _4348_ (.A1(_2760_),
    .A2(_2976_),
    .Y(_0472_),
    .B1(net68));
 sg13g2_nor2_1 _4349_ (.A(net164),
    .B(_2250_),
    .Y(_0473_));
 sg13g2_a221oi_1 _4350_ (.B2(net115),
    .C1(net192),
    .B1(_2558_),
    .A1(_0361_),
    .Y(_0474_),
    .A2(_0473_));
 sg13g2_nand2b_1 _4351_ (.Y(_0475_),
    .B(_0474_),
    .A_N(_0472_));
 sg13g2_nor2_1 _4352_ (.A(_0471_),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_nand2_1 _4353_ (.Y(_0477_),
    .A(_2709_),
    .B(_2533_));
 sg13g2_nand2_1 _4354_ (.Y(_0478_),
    .A(_2974_),
    .B(_0248_));
 sg13g2_nand3_1 _4355_ (.B(_0478_),
    .C(net189),
    .A(_0477_),
    .Y(_0479_));
 sg13g2_o21ai_1 _4356_ (.B1(net172),
    .Y(_0480_),
    .A1(_2558_),
    .A2(_2709_));
 sg13g2_nand2_1 _4357_ (.Y(_0481_),
    .A(_0479_),
    .B(_0480_));
 sg13g2_buf_1 _4358_ (.A(net155),
    .X(_0482_));
 sg13g2_nand2_1 _4359_ (.Y(_0483_),
    .A(_0481_),
    .B(net84));
 sg13g2_nand2_1 _4360_ (.Y(_0484_),
    .A(_0093_),
    .B(net204));
 sg13g2_inv_1 _4361_ (.Y(_0485_),
    .A(_0484_));
 sg13g2_nand2_1 _4362_ (.Y(_0486_),
    .A(_2519_),
    .B(net103));
 sg13g2_a21oi_1 _4363_ (.A1(_0485_),
    .A2(_0486_),
    .Y(_0487_),
    .B1(net179));
 sg13g2_a21oi_1 _4364_ (.A1(_2541_),
    .A2(_0116_),
    .Y(_0488_),
    .B1(net111));
 sg13g2_nor3_1 _4365_ (.A(net174),
    .B(_0487_),
    .C(_0488_),
    .Y(_0489_));
 sg13g2_nand2_1 _4366_ (.Y(_0490_),
    .A(_0483_),
    .B(_0489_));
 sg13g2_nand2_1 _4367_ (.Y(_0491_),
    .A(_0490_),
    .B(net151));
 sg13g2_nor2_1 _4368_ (.A(_0476_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_nor2_1 _4369_ (.A(_0467_),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_nand2_1 _4370_ (.Y(_0494_),
    .A(_0450_),
    .B(_0493_));
 sg13g2_buf_1 _4371_ (.A(_2639_),
    .X(_0495_));
 sg13g2_nand2_1 _4372_ (.Y(_0496_),
    .A(_0494_),
    .B(net212));
 sg13g2_nor2_1 _4373_ (.A(net202),
    .B(_2941_),
    .Y(_0497_));
 sg13g2_a21oi_1 _4374_ (.A1(_2942_),
    .A2(net69),
    .Y(_0498_),
    .B1(net142));
 sg13g2_o21ai_1 _4375_ (.B1(_0485_),
    .Y(_0499_),
    .A1(_0497_),
    .A2(_0498_));
 sg13g2_nand2_1 _4376_ (.Y(_0500_),
    .A(_0499_),
    .B(net135));
 sg13g2_nor2_1 _4377_ (.A(net160),
    .B(_2538_),
    .Y(_0501_));
 sg13g2_inv_1 _4378_ (.Y(_0502_),
    .A(_0501_));
 sg13g2_nand2_1 _4379_ (.Y(_0503_),
    .A(_0502_),
    .B(net129));
 sg13g2_a21oi_1 _4380_ (.A1(_0503_),
    .A2(net52),
    .Y(_0504_),
    .B1(net93));
 sg13g2_nand2_2 _4381_ (.Y(_0505_),
    .A(_2571_),
    .B(net74));
 sg13g2_nand2_1 _4382_ (.Y(_0506_),
    .A(_0216_),
    .B(net78));
 sg13g2_a21o_1 _4383_ (.A2(_0506_),
    .A1(_0505_),
    .B1(net43),
    .X(_0507_));
 sg13g2_nand3_1 _4384_ (.B(_0504_),
    .C(_0507_),
    .A(_0500_),
    .Y(_0508_));
 sg13g2_nor2_1 _4385_ (.A(net129),
    .B(net46),
    .Y(_0509_));
 sg13g2_inv_1 _4386_ (.Y(_0510_),
    .A(_0509_));
 sg13g2_inv_1 _4387_ (.Y(_0511_),
    .A(_2449_));
 sg13g2_nand3_1 _4388_ (.B(_0511_),
    .C(_2669_),
    .A(_0510_),
    .Y(_0512_));
 sg13g2_nand2_1 _4389_ (.Y(_0513_),
    .A(_2533_),
    .B(_2828_));
 sg13g2_nand3_1 _4390_ (.B(net114),
    .C(_0513_),
    .A(_0109_),
    .Y(_0514_));
 sg13g2_nand2_1 _4391_ (.Y(_0515_),
    .A(_1850_),
    .B(_2455_));
 sg13g2_nand2_1 _4392_ (.Y(_0516_),
    .A(_0515_),
    .B(net168));
 sg13g2_nand2_1 _4393_ (.Y(_0517_),
    .A(net46),
    .B(net61));
 sg13g2_nand2_1 _4394_ (.Y(_0518_),
    .A(_0516_),
    .B(_0517_));
 sg13g2_nand2_1 _4395_ (.Y(_0519_),
    .A(_0518_),
    .B(_2447_));
 sg13g2_nand3_1 _4396_ (.B(_0519_),
    .C(_2923_),
    .A(_0514_),
    .Y(_0520_));
 sg13g2_a21oi_1 _4397_ (.A1(net40),
    .A2(_0512_),
    .Y(_0521_),
    .B1(_0520_));
 sg13g2_nor2_1 _4398_ (.A(net186),
    .B(_0521_),
    .Y(_0522_));
 sg13g2_nand2_1 _4399_ (.Y(_0523_),
    .A(_0508_),
    .B(_0522_));
 sg13g2_nand2_1 _4400_ (.Y(_0524_),
    .A(_3031_),
    .B(_2863_));
 sg13g2_nand2_1 _4401_ (.Y(_0525_),
    .A(_0524_),
    .B(_1348_));
 sg13g2_nand2_1 _4402_ (.Y(_0526_),
    .A(_2507_),
    .B(_1031_));
 sg13g2_nand2_2 _4403_ (.Y(_0527_),
    .A(_0526_),
    .B(_2564_));
 sg13g2_nand2_1 _4404_ (.Y(_0528_),
    .A(_2482_),
    .B(_0435_));
 sg13g2_nand2_1 _4405_ (.Y(_0529_),
    .A(_0527_),
    .B(_0528_));
 sg13g2_a22oi_1 _4406_ (.Y(_0530_),
    .B1(_2984_),
    .B2(_0529_),
    .A2(_0525_),
    .A1(_2537_));
 sg13g2_nand2_1 _4407_ (.Y(_0531_),
    .A(_1555_),
    .B(_1741_));
 sg13g2_buf_2 _4408_ (.A(net85),
    .X(_0532_));
 sg13g2_o21ai_1 _4409_ (.B1(net47),
    .Y(_0533_),
    .A1(_2087_),
    .A2(_0531_));
 sg13g2_inv_1 _4410_ (.Y(_0534_),
    .A(_2614_));
 sg13g2_nand2_1 _4411_ (.Y(_0535_),
    .A(_2482_),
    .B(_1839_));
 sg13g2_o21ai_1 _4412_ (.B1(_0535_),
    .Y(_0536_),
    .A1(_0345_),
    .A2(_0534_));
 sg13g2_nand2_1 _4413_ (.Y(_0537_),
    .A(_0536_),
    .B(_2624_));
 sg13g2_nand3_1 _4414_ (.B(_0533_),
    .C(_0537_),
    .A(_0530_),
    .Y(_0538_));
 sg13g2_nor2b_1 _4415_ (.A(_0345_),
    .B_N(net83),
    .Y(_0539_));
 sg13g2_a21oi_1 _4416_ (.A1(net160),
    .A2(_3051_),
    .Y(_0540_),
    .B1(_0539_));
 sg13g2_o21ai_1 _4417_ (.B1(net58),
    .Y(_0541_),
    .A1(_0099_),
    .A2(_2653_));
 sg13g2_o21ai_1 _4418_ (.B1(_0541_),
    .Y(_0542_),
    .A1(net63),
    .A2(_0540_));
 sg13g2_nand2_1 _4419_ (.Y(_0543_),
    .A(_0542_),
    .B(net86));
 sg13g2_nor2_1 _4420_ (.A(net177),
    .B(_2613_),
    .Y(_0544_));
 sg13g2_inv_1 _4421_ (.Y(_0545_),
    .A(_0544_));
 sg13g2_nor2_1 _4422_ (.A(_2430_),
    .B(_2457_),
    .Y(_0546_));
 sg13g2_o21ai_1 _4423_ (.B1(_0546_),
    .Y(_0547_),
    .A1(_2486_),
    .A2(_0545_));
 sg13g2_nor2_1 _4424_ (.A(net95),
    .B(_2858_),
    .Y(_0548_));
 sg13g2_nor2_1 _4425_ (.A(_2412_),
    .B(_3045_),
    .Y(_0549_));
 sg13g2_inv_1 _4426_ (.Y(_0550_),
    .A(_0549_));
 sg13g2_a21oi_1 _4427_ (.A1(_0548_),
    .A2(_2899_),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_a21oi_1 _4428_ (.A1(_0547_),
    .A2(_0551_),
    .Y(_0552_),
    .B1(net215));
 sg13g2_nand2_1 _4429_ (.Y(_0553_),
    .A(_0543_),
    .B(_0552_));
 sg13g2_a21oi_1 _4430_ (.A1(_0538_),
    .A2(net87),
    .Y(_0554_),
    .B1(_0553_));
 sg13g2_a21oi_1 _4431_ (.A1(_0523_),
    .A2(_0554_),
    .Y(_0555_),
    .B1(net212));
 sg13g2_buf_1 _4432_ (.A(net218),
    .X(_0556_));
 sg13g2_nor2_1 _4433_ (.A(net103),
    .B(_0299_),
    .Y(_0557_));
 sg13g2_inv_1 _4434_ (.Y(_0558_),
    .A(_0557_));
 sg13g2_a21oi_1 _4435_ (.A1(_2743_),
    .A2(net96),
    .Y(_0559_),
    .B1(_0558_));
 sg13g2_nand2_1 _4436_ (.Y(_0560_),
    .A(_0559_),
    .B(net48));
 sg13g2_nand2b_1 _4437_ (.Y(_0561_),
    .B(_2966_),
    .A_N(_0459_));
 sg13g2_nand3_1 _4438_ (.B(_0561_),
    .C(net75),
    .A(_0560_),
    .Y(_0562_));
 sg13g2_nand2_1 _4439_ (.Y(_0563_),
    .A(_2766_),
    .B(net153));
 sg13g2_nor3_1 _4440_ (.A(_0563_),
    .B(_0539_),
    .C(_0123_),
    .Y(_0564_));
 sg13g2_nand3_1 _4441_ (.B(net57),
    .C(net126),
    .A(_3031_),
    .Y(_0565_));
 sg13g2_a21oi_1 _4442_ (.A1(_0497_),
    .A2(_0565_),
    .Y(_0566_),
    .B1(net84));
 sg13g2_nand2b_1 _4443_ (.Y(_0567_),
    .B(_0566_),
    .A_N(_0564_));
 sg13g2_a21oi_1 _4444_ (.A1(_0562_),
    .A2(_0567_),
    .Y(_0568_),
    .B1(_2418_));
 sg13g2_nand2_1 _4445_ (.Y(_0569_),
    .A(_1523_),
    .B(net81));
 sg13g2_inv_1 _4446_ (.Y(_0570_),
    .A(_0569_));
 sg13g2_o21ai_1 _4447_ (.B1(_0480_),
    .Y(_0571_),
    .A1(_2267_),
    .A2(_0570_));
 sg13g2_nand2_1 _4448_ (.Y(_0572_),
    .A(_0571_),
    .B(net135));
 sg13g2_inv_1 _4449_ (.Y(_0573_),
    .A(_0437_));
 sg13g2_nand2_1 _4450_ (.Y(_0574_),
    .A(_2645_),
    .B(net114));
 sg13g2_nand2_1 _4451_ (.Y(_0575_),
    .A(net82),
    .B(net173));
 sg13g2_nand2_1 _4452_ (.Y(_0576_),
    .A(_0575_),
    .B(net77));
 sg13g2_inv_1 _4453_ (.Y(_0577_),
    .A(_2456_));
 sg13g2_nor2_2 _4454_ (.A(net219),
    .B(_2734_),
    .Y(_0578_));
 sg13g2_nand2_1 _4455_ (.Y(_0579_),
    .A(_0577_),
    .B(_0578_));
 sg13g2_nand3_1 _4456_ (.B(_0576_),
    .C(_0579_),
    .A(_0574_),
    .Y(_0580_));
 sg13g2_a21oi_1 _4457_ (.A1(net53),
    .A2(_0573_),
    .Y(_0581_),
    .B1(_0580_));
 sg13g2_a21oi_1 _4458_ (.A1(_0572_),
    .A2(_0581_),
    .Y(_0582_),
    .B1(net161));
 sg13g2_nor3_1 _4459_ (.A(net183),
    .B(_0568_),
    .C(_0582_),
    .Y(_0583_));
 sg13g2_o21ai_1 _4460_ (.B1(net92),
    .Y(_0584_),
    .A1(_2585_),
    .A2(_0573_));
 sg13g2_inv_1 _4461_ (.Y(_0585_),
    .A(_2506_));
 sg13g2_nor2_1 _4462_ (.A(_0585_),
    .B(_2742_),
    .Y(_0586_));
 sg13g2_a22oi_1 _4463_ (.Y(_0587_),
    .B1(net120),
    .B2(_0586_),
    .A2(_0577_),
    .A1(net77));
 sg13g2_nand2_1 _4464_ (.Y(_0588_),
    .A(_0584_),
    .B(_0587_));
 sg13g2_nand2_1 _4465_ (.Y(_0589_),
    .A(_0588_),
    .B(net167));
 sg13g2_nand2_1 _4466_ (.Y(_0590_),
    .A(_0422_),
    .B(net201));
 sg13g2_a21oi_1 _4467_ (.A1(_0169_),
    .A2(_3035_),
    .Y(_0591_),
    .B1(_2531_));
 sg13g2_a21oi_1 _4468_ (.A1(_0590_),
    .A2(net58),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_o21ai_1 _4469_ (.B1(_2399_),
    .Y(_0593_),
    .A1(net195),
    .A2(_2936_));
 sg13g2_nand2_1 _4470_ (.Y(_0594_),
    .A(_0593_),
    .B(_0461_));
 sg13g2_nand2_1 _4471_ (.Y(_0595_),
    .A(_0594_),
    .B(net116));
 sg13g2_nand2_1 _4472_ (.Y(_0596_),
    .A(_0592_),
    .B(_0595_));
 sg13g2_nand2_1 _4473_ (.Y(_0597_),
    .A(_0596_),
    .B(net93));
 sg13g2_a21oi_1 _4474_ (.A1(net41),
    .A2(net45),
    .Y(_0598_),
    .B1(_1882_));
 sg13g2_a21oi_1 _4475_ (.A1(net65),
    .A2(net78),
    .Y(_0599_),
    .B1(net122));
 sg13g2_nand3_1 _4476_ (.B(net45),
    .C(net131),
    .A(net44),
    .Y(_0600_));
 sg13g2_a22oi_1 _4477_ (.Y(_0601_),
    .B1(_0599_),
    .B2(_0600_),
    .A2(_0598_),
    .A1(_0282_));
 sg13g2_nand2_1 _4478_ (.Y(_0602_),
    .A(_0601_),
    .B(net171));
 sg13g2_nand3_1 _4479_ (.B(_0597_),
    .C(_0602_),
    .A(_0589_),
    .Y(_0603_));
 sg13g2_nand2_1 _4480_ (.Y(_0604_),
    .A(_0603_),
    .B(net166));
 sg13g2_nand2_1 _4481_ (.Y(_0605_),
    .A(_0583_),
    .B(_0604_));
 sg13g2_nand2_1 _4482_ (.Y(_0606_),
    .A(_0555_),
    .B(_0605_));
 sg13g2_nand2_1 _4483_ (.Y(_0023_),
    .A(_0496_),
    .B(_0606_));
 sg13g2_nand2_1 _4484_ (.Y(_0607_),
    .A(_0437_),
    .B(_0511_));
 sg13g2_a21oi_1 _4485_ (.A1(_3046_),
    .A2(net59),
    .Y(_0608_),
    .B1(_2606_));
 sg13g2_nor2_1 _4486_ (.A(_2526_),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_a21oi_1 _4487_ (.A1(_0607_),
    .A2(_2819_),
    .Y(_0610_),
    .B1(_0609_));
 sg13g2_nand2_1 _4488_ (.Y(_0611_),
    .A(_0248_),
    .B(net180));
 sg13g2_nor3_1 _4489_ (.A(net198),
    .B(_2972_),
    .C(_0611_),
    .Y(_0612_));
 sg13g2_nand2_1 _4490_ (.Y(_0613_),
    .A(_0107_),
    .B(net219));
 sg13g2_nand2b_1 _4491_ (.Y(_0614_),
    .B(_0613_),
    .A_N(_0612_));
 sg13g2_nand2_1 _4492_ (.Y(_0615_),
    .A(_2598_),
    .B(net59));
 sg13g2_nand3_1 _4493_ (.B(_2745_),
    .C(net91),
    .A(_0615_),
    .Y(_0616_));
 sg13g2_nand2_1 _4494_ (.Y(_0617_),
    .A(_0614_),
    .B(_0616_));
 sg13g2_nand2_1 _4495_ (.Y(_0618_),
    .A(_0610_),
    .B(_0617_));
 sg13g2_nand2_1 _4496_ (.Y(_0619_),
    .A(_0618_),
    .B(net86));
 sg13g2_nand2_1 _4497_ (.Y(_0620_),
    .A(_3031_),
    .B(_2637_));
 sg13g2_nand2_1 _4498_ (.Y(_0621_),
    .A(_0620_),
    .B(net74));
 sg13g2_nand3_1 _4499_ (.B(_0136_),
    .C(net147),
    .A(_0621_),
    .Y(_0622_));
 sg13g2_nor2_1 _4500_ (.A(_1206_),
    .B(_2437_),
    .Y(_0623_));
 sg13g2_a21oi_1 _4501_ (.A1(_0623_),
    .A2(_1304_),
    .Y(_0624_),
    .B1(net195));
 sg13g2_nand2_1 _4502_ (.Y(_0625_),
    .A(_0944_),
    .B(_0624_));
 sg13g2_nand3_1 _4503_ (.B(_0625_),
    .C(net116),
    .A(_0622_),
    .Y(_0626_));
 sg13g2_nor2_1 _4504_ (.A(net172),
    .B(_0484_),
    .Y(_0627_));
 sg13g2_nand2_1 _4505_ (.Y(_0628_),
    .A(_0422_),
    .B(_0627_));
 sg13g2_nand2_1 _4506_ (.Y(_0629_),
    .A(net65),
    .B(net46));
 sg13g2_nand3_1 _4507_ (.B(_2402_),
    .C(net95),
    .A(_0629_),
    .Y(_0630_));
 sg13g2_nand3_1 _4508_ (.B(_0630_),
    .C(net191),
    .A(_0628_),
    .Y(_0631_));
 sg13g2_nand2_1 _4509_ (.Y(_0632_),
    .A(_0626_),
    .B(_0631_));
 sg13g2_nand2_1 _4510_ (.Y(_0633_),
    .A(_0632_),
    .B(_2890_));
 sg13g2_nand2_1 _4511_ (.Y(_0634_),
    .A(_0619_),
    .B(_0633_));
 sg13g2_nand2_2 _4512_ (.Y(_0635_),
    .A(net78),
    .B(net170));
 sg13g2_nand3_1 _4513_ (.B(net45),
    .C(net124),
    .A(_0635_),
    .Y(_0636_));
 sg13g2_nand2_1 _4514_ (.Y(_0637_),
    .A(_0636_),
    .B(_2669_));
 sg13g2_nand3_1 _4515_ (.B(net88),
    .C(_0478_),
    .A(_0944_),
    .Y(_0638_));
 sg13g2_a21oi_1 _4516_ (.A1(_2784_),
    .A2(net104),
    .Y(_0639_),
    .B1(net51));
 sg13g2_nand2_1 _4517_ (.Y(_0640_),
    .A(_2708_),
    .B(net132));
 sg13g2_nand2_1 _4518_ (.Y(_0641_),
    .A(_0640_),
    .B(_2882_));
 sg13g2_nor2_1 _4519_ (.A(_0639_),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_nor2_1 _4520_ (.A(net50),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_a22oi_1 _4521_ (.Y(_0644_),
    .B1(_0638_),
    .B2(_0643_),
    .A2(_0637_),
    .A1(_2624_));
 sg13g2_nand2_1 _4522_ (.Y(_0645_),
    .A(_0414_),
    .B(_2828_));
 sg13g2_nand2_1 _4523_ (.Y(_0646_),
    .A(_0645_),
    .B(_0239_));
 sg13g2_a21oi_1 _4524_ (.A1(_0646_),
    .A2(_0114_),
    .Y(_0647_),
    .B1(_2946_));
 sg13g2_nand3_1 _4525_ (.B(_2793_),
    .C(_2583_),
    .A(_0209_),
    .Y(_0648_));
 sg13g2_nand2_1 _4526_ (.Y(_0649_),
    .A(_0216_),
    .B(_2713_));
 sg13g2_a21oi_1 _4527_ (.A1(_0649_),
    .A2(_3025_),
    .Y(_0650_),
    .B1(net97));
 sg13g2_nand2_1 _4528_ (.Y(_0651_),
    .A(_0648_),
    .B(_0650_));
 sg13g2_nand2_1 _4529_ (.Y(_0652_),
    .A(_2825_),
    .B(net149));
 sg13g2_o21ai_1 _4530_ (.B1(net203),
    .Y(_0653_),
    .A1(_2571_),
    .A2(_0652_));
 sg13g2_nand2_1 _4531_ (.Y(_0654_),
    .A(_0229_),
    .B(_1785_));
 sg13g2_o21ai_1 _4532_ (.B1(_0654_),
    .Y(_0655_),
    .A1(_2686_),
    .A2(_0570_));
 sg13g2_nor2_1 _4533_ (.A(_0653_),
    .B(_0655_),
    .Y(_0656_));
 sg13g2_nand2_1 _4534_ (.Y(_0657_),
    .A(_0651_),
    .B(_0656_));
 sg13g2_nand2_1 _4535_ (.Y(_0658_),
    .A(_0657_),
    .B(_2594_));
 sg13g2_a21oi_1 _4536_ (.A1(_0644_),
    .A2(_0647_),
    .Y(_0659_),
    .B1(_0658_));
 sg13g2_a21oi_1 _4537_ (.A1(_0634_),
    .A2(_3010_),
    .Y(_0660_),
    .B1(_0659_));
 sg13g2_nand2_1 _4538_ (.Y(_0661_),
    .A(_2620_),
    .B(net108));
 sg13g2_inv_1 _4539_ (.Y(_0662_),
    .A(_2858_));
 sg13g2_a21oi_1 _4540_ (.A1(_0661_),
    .A2(_0662_),
    .Y(_0663_),
    .B1(_1457_));
 sg13g2_nand2_1 _4541_ (.Y(_0664_),
    .A(_2280_),
    .B(net198));
 sg13g2_a21oi_1 _4542_ (.A1(net44),
    .A2(net94),
    .Y(_0665_),
    .B1(_0664_));
 sg13g2_nor3_1 _4543_ (.A(_0663_),
    .B(_0665_),
    .C(_0376_),
    .Y(_0666_));
 sg13g2_inv_1 _4544_ (.Y(_0667_),
    .A(_2699_));
 sg13g2_nor2_1 _4545_ (.A(_0667_),
    .B(_2964_),
    .Y(_0668_));
 sg13g2_nor2_1 _4546_ (.A(net195),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_nand2_1 _4547_ (.Y(_0670_),
    .A(_0669_),
    .B(_0454_));
 sg13g2_nor2_1 _4548_ (.A(_1763_),
    .B(_2872_),
    .Y(_0671_));
 sg13g2_inv_1 _4549_ (.Y(_0672_),
    .A(_2993_));
 sg13g2_a21oi_1 _4550_ (.A1(_0671_),
    .A2(_0672_),
    .Y(_0673_),
    .B1(net155));
 sg13g2_nand2_1 _4551_ (.Y(_0674_),
    .A(_0670_),
    .B(_0673_));
 sg13g2_a21oi_1 _4552_ (.A1(_0666_),
    .A2(_0674_),
    .Y(_0675_),
    .B1(net187));
 sg13g2_nand2_1 _4553_ (.Y(_0676_),
    .A(_0640_),
    .B(net137));
 sg13g2_nor2_1 _4554_ (.A(_2430_),
    .B(_2853_),
    .Y(_0677_));
 sg13g2_a21oi_1 _4555_ (.A1(_0677_),
    .A2(_0196_),
    .Y(_0678_),
    .B1(_2492_));
 sg13g2_o21ai_1 _4556_ (.B1(_0678_),
    .Y(_0679_),
    .A1(_0676_),
    .A2(_2934_));
 sg13g2_nor2_1 _4557_ (.A(net106),
    .B(_3046_),
    .Y(_0680_));
 sg13g2_nor2_1 _4558_ (.A(net59),
    .B(_0680_),
    .Y(_0681_));
 sg13g2_o21ai_1 _4559_ (.B1(_2771_),
    .Y(_0682_),
    .A1(_2693_),
    .A2(_0681_));
 sg13g2_nor3_1 _4560_ (.A(net159),
    .B(_0911_),
    .C(_2644_),
    .Y(_0683_));
 sg13g2_nor2_1 _4561_ (.A(net192),
    .B(_0683_),
    .Y(_0684_));
 sg13g2_nand3_1 _4562_ (.B(_0682_),
    .C(_0684_),
    .A(_0679_),
    .Y(_0685_));
 sg13g2_nand2_1 _4563_ (.Y(_0686_),
    .A(_0675_),
    .B(_0685_));
 sg13g2_nand2_1 _4564_ (.Y(_0687_),
    .A(_0460_),
    .B(net132));
 sg13g2_inv_1 _4565_ (.Y(_0688_),
    .A(_2556_));
 sg13g2_a21oi_1 _4566_ (.A1(_0687_),
    .A2(_0688_),
    .Y(_0689_),
    .B1(net68));
 sg13g2_nand2_1 _4567_ (.Y(_0690_),
    .A(_2484_),
    .B(_0922_));
 sg13g2_nor3_1 _4568_ (.A(net159),
    .B(net61),
    .C(_0318_),
    .Y(_0691_));
 sg13g2_a21oi_1 _4569_ (.A1(_0690_),
    .A2(_2458_),
    .Y(_0692_),
    .B1(_0691_));
 sg13g2_nand2_1 _4570_ (.Y(_0693_),
    .A(_0535_),
    .B(_2954_));
 sg13g2_nand2_1 _4571_ (.Y(_0694_),
    .A(_0693_),
    .B(net149));
 sg13g2_nand2_1 _4572_ (.Y(_0695_),
    .A(_0692_),
    .B(_0694_));
 sg13g2_nor2_1 _4573_ (.A(_0689_),
    .B(_0695_),
    .Y(_0696_));
 sg13g2_nor2_1 _4574_ (.A(net161),
    .B(_0696_),
    .Y(_0697_));
 sg13g2_a21oi_1 _4575_ (.A1(_1730_),
    .A2(net172),
    .Y(_0698_),
    .B1(net219));
 sg13g2_nand2_1 _4576_ (.Y(_0699_),
    .A(_0576_),
    .B(_0698_));
 sg13g2_o21ai_1 _4577_ (.B1(net148),
    .Y(_0700_),
    .A1(_3034_),
    .A2(_0123_));
 sg13g2_nor2b_1 _4578_ (.A(_0699_),
    .B_N(_0700_),
    .Y(_0701_));
 sg13g2_nand2_1 _4579_ (.Y(_0702_),
    .A(_3046_),
    .B(net113));
 sg13g2_a21oi_1 _4580_ (.A1(_0702_),
    .A2(_0280_),
    .Y(_0703_),
    .B1(net137));
 sg13g2_inv_1 _4581_ (.Y(_0704_),
    .A(_0338_));
 sg13g2_a21oi_1 _4582_ (.A1(_2273_),
    .A2(_2433_),
    .Y(_0705_),
    .B1(_2421_));
 sg13g2_o21ai_1 _4583_ (.B1(_0705_),
    .Y(_0706_),
    .A1(net153),
    .A2(_0704_));
 sg13g2_o21ai_1 _4584_ (.B1(_0350_),
    .Y(_0707_),
    .A1(_0703_),
    .A2(_0706_));
 sg13g2_nor2_1 _4585_ (.A(_0701_),
    .B(_0707_),
    .Y(_0708_));
 sg13g2_nor2_1 _4586_ (.A(_0697_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_nand2_1 _4587_ (.Y(_0710_),
    .A(_0686_),
    .B(_0709_));
 sg13g2_nand2_1 _4588_ (.Y(_0711_),
    .A(_0710_),
    .B(_0556_));
 sg13g2_nand2_1 _4589_ (.Y(_0712_),
    .A(_0660_),
    .B(_0711_));
 sg13g2_buf_1 _4590_ (.A(_2640_),
    .X(_0713_));
 sg13g2_nand2_1 _4591_ (.Y(_0714_),
    .A(_0712_),
    .B(net182));
 sg13g2_nand2_1 _4592_ (.Y(_0715_),
    .A(_0342_),
    .B(net137));
 sg13g2_a22oi_1 _4593_ (.Y(_0716_),
    .B1(_0563_),
    .B2(_0715_),
    .A2(_2733_),
    .A1(_0238_));
 sg13g2_o21ai_1 _4594_ (.B1(net199),
    .Y(_0717_),
    .A1(_2405_),
    .A2(_0716_));
 sg13g2_o21ai_1 _4595_ (.B1(_0485_),
    .Y(_0718_),
    .A1(_0134_),
    .A2(_2942_));
 sg13g2_nand2_2 _4596_ (.Y(_0719_),
    .A(_2995_),
    .B(net130));
 sg13g2_nand3_1 _4597_ (.B(_2793_),
    .C(_0719_),
    .A(_2933_),
    .Y(_0720_));
 sg13g2_o21ai_1 _4598_ (.B1(_0720_),
    .Y(_0721_),
    .A1(net139),
    .A2(_0718_));
 sg13g2_nor2_1 _4599_ (.A(_3045_),
    .B(_0721_),
    .Y(_0722_));
 sg13g2_nor2_1 _4600_ (.A(_0717_),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_inv_1 _4601_ (.Y(_0724_),
    .A(_2045_));
 sg13g2_o21ai_1 _4602_ (.B1(net176),
    .Y(_0726_),
    .A1(_2604_),
    .A2(_0724_));
 sg13g2_buf_1 _4603_ (.A(_0726_),
    .X(_0727_));
 sg13g2_nand2b_1 _4604_ (.Y(_0728_),
    .B(_0727_),
    .A_N(_2929_));
 sg13g2_nand2_1 _4605_ (.Y(_0729_),
    .A(_0728_),
    .B(net95));
 sg13g2_nand2_1 _4606_ (.Y(_0730_),
    .A(_0285_),
    .B(_0235_));
 sg13g2_nand2_1 _4607_ (.Y(_0731_),
    .A(_0729_),
    .B(_0730_));
 sg13g2_nand2_1 _4608_ (.Y(_0732_),
    .A(_0731_),
    .B(net134));
 sg13g2_inv_1 _4609_ (.Y(_0733_),
    .A(_2791_));
 sg13g2_nand2_1 _4610_ (.Y(_0734_),
    .A(_0733_),
    .B(_2812_));
 sg13g2_a21oi_1 _4611_ (.A1(_0734_),
    .A2(_0506_),
    .Y(_0735_),
    .B1(net68));
 sg13g2_a21oi_1 _4612_ (.A1(_0314_),
    .A2(_0125_),
    .Y(_0737_),
    .B1(net128));
 sg13g2_nor2_1 _4613_ (.A(_0735_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_nand2_1 _4614_ (.Y(_0739_),
    .A(_0732_),
    .B(_0738_));
 sg13g2_nand2_1 _4615_ (.Y(_0740_),
    .A(_0739_),
    .B(net125));
 sg13g2_nand2_1 _4616_ (.Y(_0741_),
    .A(_0723_),
    .B(_0740_));
 sg13g2_nand4_1 _4617_ (.B(net142),
    .C(_3019_),
    .A(_0461_),
    .Y(_0742_),
    .D(net201));
 sg13g2_inv_1 _4618_ (.Y(_0743_),
    .A(_0137_));
 sg13g2_nand2_2 _4619_ (.Y(_0744_),
    .A(_0743_),
    .B(net130));
 sg13g2_nor2_1 _4620_ (.A(net197),
    .B(_3034_),
    .Y(_0745_));
 sg13g2_a21oi_1 _4621_ (.A1(_0744_),
    .A2(_0745_),
    .Y(_0746_),
    .B1(net185));
 sg13g2_nand2_1 _4622_ (.Y(_0748_),
    .A(_0742_),
    .B(_0746_));
 sg13g2_nand2_1 _4623_ (.Y(_0749_),
    .A(_2557_),
    .B(_2775_));
 sg13g2_nand2_1 _4624_ (.Y(_0750_),
    .A(_2919_),
    .B(_1130_));
 sg13g2_nor2_1 _4625_ (.A(_2420_),
    .B(_0750_),
    .Y(_0751_));
 sg13g2_buf_2 _4626_ (.A(_0751_),
    .X(_0752_));
 sg13g2_a22oi_1 _4627_ (.Y(_0753_),
    .B1(_0752_),
    .B2(_0586_),
    .A2(_0749_),
    .A1(net85));
 sg13g2_nand2_1 _4628_ (.Y(_0754_),
    .A(_0748_),
    .B(_0753_));
 sg13g2_nand2_1 _4629_ (.Y(_0755_),
    .A(_0754_),
    .B(net125));
 sg13g2_nor2_1 _4630_ (.A(_2501_),
    .B(_2785_),
    .Y(_0756_));
 sg13g2_o21ai_1 _4631_ (.B1(_2361_),
    .Y(_0757_),
    .A1(_2399_),
    .A2(_0218_));
 sg13g2_nor2_1 _4632_ (.A(_2734_),
    .B(_0204_),
    .Y(_0759_));
 sg13g2_nor3_1 _4633_ (.A(_0756_),
    .B(_0757_),
    .C(_0759_),
    .Y(_0760_));
 sg13g2_nand2_1 _4634_ (.Y(_0761_),
    .A(_0719_),
    .B(_0704_));
 sg13g2_nand3_1 _4635_ (.B(_2628_),
    .C(_0381_),
    .A(_0761_),
    .Y(_0762_));
 sg13g2_nand2_1 _4636_ (.Y(_0763_),
    .A(_2379_),
    .B(net226));
 sg13g2_a21o_1 _4637_ (.A2(_0763_),
    .A1(_2533_),
    .B1(_2665_),
    .X(_0764_));
 sg13g2_nand2b_1 _4638_ (.Y(_0765_),
    .B(net167),
    .A_N(_0764_));
 sg13g2_nand3_1 _4639_ (.B(_0765_),
    .C(_2592_),
    .A(_0762_),
    .Y(_0766_));
 sg13g2_nor2_1 _4640_ (.A(_0760_),
    .B(_0766_),
    .Y(_0767_));
 sg13g2_nand2_1 _4641_ (.Y(_0768_),
    .A(_0755_),
    .B(_0767_));
 sg13g2_nand2_1 _4642_ (.Y(_0770_),
    .A(_0741_),
    .B(_0768_));
 sg13g2_nand2_1 _4643_ (.Y(_0771_),
    .A(_0770_),
    .B(net194));
 sg13g2_nor2_1 _4644_ (.A(net51),
    .B(_2461_),
    .Y(_0772_));
 sg13g2_nand2_1 _4645_ (.Y(_0773_),
    .A(_2768_),
    .B(_2904_));
 sg13g2_nand2_1 _4646_ (.Y(_0774_),
    .A(_0773_),
    .B(_1304_));
 sg13g2_nand3b_1 _4647_ (.B(_0774_),
    .C(net134),
    .Y(_0775_),
    .A_N(_0772_));
 sg13g2_inv_1 _4648_ (.Y(_0776_),
    .A(_2457_));
 sg13g2_nor2_1 _4649_ (.A(net196),
    .B(_2700_),
    .Y(_0777_));
 sg13g2_a21oi_1 _4650_ (.A1(_0776_),
    .A2(_0777_),
    .Y(_0778_),
    .B1(_2562_));
 sg13g2_nand2_1 _4651_ (.Y(_0779_),
    .A(_2740_),
    .B(net137));
 sg13g2_o21ai_1 _4652_ (.B1(_0779_),
    .Y(_0781_),
    .A1(net106),
    .A2(_2938_));
 sg13g2_nand3_1 _4653_ (.B(net157),
    .C(net96),
    .A(_2482_),
    .Y(_0782_));
 sg13g2_nand2_1 _4654_ (.Y(_0783_),
    .A(_0781_),
    .B(_0782_));
 sg13g2_a22oi_1 _4655_ (.Y(_0784_),
    .B1(net167),
    .B2(_0783_),
    .A2(_0778_),
    .A1(_0775_));
 sg13g2_a21oi_1 _4656_ (.A1(_0733_),
    .A2(_0182_),
    .Y(_0785_),
    .B1(_0368_));
 sg13g2_nand2_1 _4657_ (.Y(_0786_),
    .A(_2498_),
    .B(net97));
 sg13g2_nand2_1 _4658_ (.Y(_0787_),
    .A(_0785_),
    .B(_0786_));
 sg13g2_nor2_1 _4659_ (.A(_2842_),
    .B(_2857_),
    .Y(_0788_));
 sg13g2_nor2_1 _4660_ (.A(_2666_),
    .B(_2914_),
    .Y(_0789_));
 sg13g2_nor2_1 _4661_ (.A(_2431_),
    .B(_2776_),
    .Y(_0790_));
 sg13g2_nand2_1 _4662_ (.Y(_0792_),
    .A(_2433_),
    .B(_2386_));
 sg13g2_inv_1 _4663_ (.Y(_0793_),
    .A(_0792_));
 sg13g2_nor2_1 _4664_ (.A(_0793_),
    .B(_2656_),
    .Y(_0794_));
 sg13g2_inv_1 _4665_ (.Y(_0795_),
    .A(_0794_));
 sg13g2_a22oi_1 _4666_ (.Y(_0796_),
    .B1(_0790_),
    .B2(_0795_),
    .A2(_0789_),
    .A1(_0788_));
 sg13g2_a22oi_1 _4667_ (.Y(_0797_),
    .B1(net171),
    .B2(_0796_),
    .A2(_0787_),
    .A1(_2588_));
 sg13g2_nand2_1 _4668_ (.Y(_0798_),
    .A(_0784_),
    .B(_0797_));
 sg13g2_nand2_1 _4669_ (.Y(_0799_),
    .A(_0798_),
    .B(net166));
 sg13g2_nand2_1 _4670_ (.Y(_0800_),
    .A(_2137_),
    .B(_2318_));
 sg13g2_nand2_1 _4671_ (.Y(_0801_),
    .A(_0800_),
    .B(_2830_));
 sg13g2_nand2_1 _4672_ (.Y(_0803_),
    .A(_2995_),
    .B(_2733_));
 sg13g2_a21oi_1 _4673_ (.A1(_0801_),
    .A2(_0803_),
    .Y(_0804_),
    .B1(net84));
 sg13g2_nor3_1 _4674_ (.A(net139),
    .B(_2727_),
    .C(_0239_),
    .Y(_0805_));
 sg13g2_nor2_1 _4675_ (.A(_0804_),
    .B(_0805_),
    .Y(_0806_));
 sg13g2_inv_1 _4676_ (.Y(_0807_),
    .A(_0099_));
 sg13g2_nand2_1 _4677_ (.Y(_0808_),
    .A(_0704_),
    .B(_0807_));
 sg13g2_o21ai_1 _4678_ (.B1(_2913_),
    .Y(_0809_),
    .A1(net39),
    .A2(net46));
 sg13g2_a22oi_1 _4679_ (.Y(_0810_),
    .B1(net54),
    .B2(_0809_),
    .A2(net66),
    .A1(_0808_));
 sg13g2_a21oi_1 _4680_ (.A1(_0806_),
    .A2(_0810_),
    .Y(_0811_),
    .B1(net161));
 sg13g2_nand2_1 _4681_ (.Y(_0812_),
    .A(_1555_),
    .B(_0702_));
 sg13g2_a21oi_1 _4682_ (.A1(_0812_),
    .A2(_0151_),
    .Y(_0814_),
    .B1(net218));
 sg13g2_nor2b_1 _4683_ (.A(_0811_),
    .B_N(_0814_),
    .Y(_0815_));
 sg13g2_a21oi_1 _4684_ (.A1(_0799_),
    .A2(_0815_),
    .Y(_0816_),
    .B1(_2640_));
 sg13g2_nand2_1 _4685_ (.Y(_0817_),
    .A(_0771_),
    .B(_0816_));
 sg13g2_nand2_1 _4686_ (.Y(_0024_),
    .A(_0714_),
    .B(_0817_));
 sg13g2_nand2_1 _4687_ (.Y(_0818_),
    .A(_2801_),
    .B(net57));
 sg13g2_nand3_1 _4688_ (.B(net48),
    .C(_0233_),
    .A(_0818_),
    .Y(_0819_));
 sg13g2_nand3_1 _4689_ (.B(_2077_),
    .C(net89),
    .A(_0744_),
    .Y(_0820_));
 sg13g2_nand3_1 _4690_ (.B(net135),
    .C(_0820_),
    .A(_0819_),
    .Y(_0821_));
 sg13g2_inv_1 _4691_ (.Y(_0822_),
    .A(_0138_));
 sg13g2_a21o_1 _4692_ (.A2(_2656_),
    .A1(_0822_),
    .B1(net67),
    .X(_0824_));
 sg13g2_a21oi_1 _4693_ (.A1(net73),
    .A2(net62),
    .Y(_0825_),
    .B1(net150));
 sg13g2_nand3_1 _4694_ (.B(_0824_),
    .C(_0825_),
    .A(_0821_),
    .Y(_0826_));
 sg13g2_nand2_1 _4695_ (.Y(_0827_),
    .A(_0671_),
    .B(_2491_));
 sg13g2_nand2_1 _4696_ (.Y(_0828_),
    .A(_0827_),
    .B(_2547_));
 sg13g2_nor3_1 _4697_ (.A(_1730_),
    .B(_2479_),
    .C(_2600_),
    .Y(_0829_));
 sg13g2_nand2_1 _4698_ (.Y(_0830_),
    .A(net124),
    .B(net71));
 sg13g2_a21oi_1 _4699_ (.A1(_0139_),
    .A2(_0830_),
    .Y(_0831_),
    .B1(net152));
 sg13g2_nor3_1 _4700_ (.A(_0828_),
    .B(_0829_),
    .C(_0831_),
    .Y(_0832_));
 sg13g2_nor2_1 _4701_ (.A(net143),
    .B(_0832_),
    .Y(_0833_));
 sg13g2_inv_1 _4702_ (.Y(_0835_),
    .A(_0429_));
 sg13g2_inv_1 _4703_ (.Y(_0836_),
    .A(_0750_));
 sg13g2_a21oi_1 _4704_ (.A1(_0835_),
    .A2(_0836_),
    .Y(_0837_),
    .B1(net191));
 sg13g2_nand3_1 _4705_ (.B(_2893_),
    .C(_2184_),
    .A(_0367_),
    .Y(_0838_));
 sg13g2_nand2_1 _4706_ (.Y(_0839_),
    .A(_0837_),
    .B(_0838_));
 sg13g2_inv_1 _4707_ (.Y(_0840_),
    .A(_3024_));
 sg13g2_inv_1 _4708_ (.Y(_0841_),
    .A(_0211_));
 sg13g2_nor2_1 _4709_ (.A(_2489_),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_a22oi_1 _4710_ (.Y(_0843_),
    .B1(net66),
    .B2(_0842_),
    .A2(_0840_),
    .A1(net98));
 sg13g2_a21oi_1 _4711_ (.A1(_0839_),
    .A2(_0843_),
    .Y(_0844_),
    .B1(net150));
 sg13g2_nand2_1 _4712_ (.Y(_0846_),
    .A(_0792_),
    .B(_1097_));
 sg13g2_buf_2 _4713_ (.A(_0846_),
    .X(_0847_));
 sg13g2_nand2_1 _4714_ (.Y(_0848_),
    .A(_0847_),
    .B(net148));
 sg13g2_inv_1 _4715_ (.Y(_0849_),
    .A(_0848_));
 sg13g2_o21ai_1 _4716_ (.B1(_0849_),
    .Y(_0850_),
    .A1(net71),
    .A2(_2995_));
 sg13g2_a21oi_1 _4717_ (.A1(net56),
    .A2(_0197_),
    .Y(_0851_),
    .B1(_3045_));
 sg13g2_nor2_1 _4718_ (.A(net169),
    .B(_0310_),
    .Y(_0852_));
 sg13g2_o21ai_1 _4719_ (.B1(_0088_),
    .Y(_0853_),
    .A1(net88),
    .A2(_0852_));
 sg13g2_a22oi_1 _4720_ (.Y(_0854_),
    .B1(net167),
    .B2(_0853_),
    .A2(_0851_),
    .A1(_0850_));
 sg13g2_nand2b_1 _4721_ (.Y(_0855_),
    .B(_0854_),
    .A_N(_0844_));
 sg13g2_a22oi_1 _4722_ (.Y(_0857_),
    .B1(net166),
    .B2(_0855_),
    .A2(_0833_),
    .A1(_0826_));
 sg13g2_nand2_1 _4723_ (.Y(_0858_),
    .A(_0857_),
    .B(net194));
 sg13g2_nor3_1 _4724_ (.A(net189),
    .B(_3004_),
    .C(_2606_),
    .Y(_0859_));
 sg13g2_a21oi_1 _4725_ (.A1(_0208_),
    .A2(net213),
    .Y(_0860_),
    .B1(net153));
 sg13g2_nor2_1 _4726_ (.A(_0859_),
    .B(_0860_),
    .Y(_0861_));
 sg13g2_nand2_1 _4727_ (.Y(_0862_),
    .A(_0861_),
    .B(net152));
 sg13g2_nand3_1 _4728_ (.B(net54),
    .C(_2893_),
    .A(_2524_),
    .Y(_0863_));
 sg13g2_o21ai_1 _4729_ (.B1(net90),
    .Y(_0864_),
    .A1(_2489_),
    .A2(_0841_));
 sg13g2_nand4_1 _4730_ (.B(_0863_),
    .C(net141),
    .A(_0862_),
    .Y(_0865_),
    .D(_0864_));
 sg13g2_nor2_2 _4731_ (.A(_2488_),
    .B(_2434_),
    .Y(_0866_));
 sg13g2_nor2_1 _4732_ (.A(_1337_),
    .B(_2215_),
    .Y(_0868_));
 sg13g2_nor2_1 _4733_ (.A(_2500_),
    .B(_0868_),
    .Y(_0869_));
 sg13g2_a22oi_1 _4734_ (.Y(_0870_),
    .B1(_0869_),
    .B2(_0719_),
    .A2(net185),
    .A1(_2490_));
 sg13g2_o21ai_1 _4735_ (.B1(_0870_),
    .Y(_0871_),
    .A1(net43),
    .A2(_0866_));
 sg13g2_nand2_1 _4736_ (.Y(_0872_),
    .A(_0871_),
    .B(net93));
 sg13g2_nand2_1 _4737_ (.Y(_0873_),
    .A(_0865_),
    .B(_0872_));
 sg13g2_nand2_1 _4738_ (.Y(_0874_),
    .A(_0873_),
    .B(net166));
 sg13g2_nand2_1 _4739_ (.Y(_0875_),
    .A(_2662_),
    .B(net226));
 sg13g2_a21oi_1 _4740_ (.A1(net76),
    .A2(_0875_),
    .Y(_0876_),
    .B1(_0860_));
 sg13g2_nor2_1 _4741_ (.A(net226),
    .B(_0792_),
    .Y(_0877_));
 sg13g2_nor2_1 _4742_ (.A(net163),
    .B(_0877_),
    .Y(_0879_));
 sg13g2_nand2_2 _4743_ (.Y(_0880_),
    .A(_0137_),
    .B(net213));
 sg13g2_inv_1 _4744_ (.Y(_0881_),
    .A(_0880_));
 sg13g2_nor2_1 _4745_ (.A(net158),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_nor3_1 _4746_ (.A(net50),
    .B(_0879_),
    .C(_0882_),
    .Y(_0883_));
 sg13g2_a21oi_1 _4747_ (.A1(_0876_),
    .A2(_0297_),
    .Y(_0884_),
    .B1(_0883_));
 sg13g2_o21ai_1 _4748_ (.B1(_0351_),
    .Y(_0885_),
    .A1(net124),
    .A2(_2921_));
 sg13g2_nand2_1 _4749_ (.Y(_0886_),
    .A(_0885_),
    .B(_2630_));
 sg13g2_a21oi_1 _4750_ (.A1(_0884_),
    .A2(_2890_),
    .Y(_0887_),
    .B1(_0886_));
 sg13g2_a21oi_1 _4751_ (.A1(_0874_),
    .A2(_0887_),
    .Y(_0888_),
    .B1(_0713_));
 sg13g2_nand2_1 _4752_ (.Y(_0890_),
    .A(_0858_),
    .B(_0888_));
 sg13g2_nand2_1 _4753_ (.Y(_0891_),
    .A(_2662_),
    .B(net213));
 sg13g2_nand3_1 _4754_ (.B(_2893_),
    .C(net122),
    .A(_2715_),
    .Y(_0892_));
 sg13g2_inv_1 _4755_ (.Y(_0893_),
    .A(_0310_));
 sg13g2_a21oi_1 _4756_ (.A1(_0893_),
    .A2(_0836_),
    .Y(_0894_),
    .B1(_2860_));
 sg13g2_a22oi_1 _4757_ (.Y(_0895_),
    .B1(_0892_),
    .B2(_0894_),
    .A2(_0891_),
    .A1(net54));
 sg13g2_buf_1 _4758_ (.A(net193),
    .X(_0896_));
 sg13g2_nand2b_1 _4759_ (.Y(_0897_),
    .B(net133),
    .A_N(_0895_));
 sg13g2_nor2_1 _4760_ (.A(_2380_),
    .B(_2455_),
    .Y(_0898_));
 sg13g2_nor3_1 _4761_ (.A(net112),
    .B(_0898_),
    .C(_0866_),
    .Y(_0899_));
 sg13g2_nor2_1 _4762_ (.A(_2388_),
    .B(_1577_),
    .Y(_0901_));
 sg13g2_nand2_1 _4763_ (.Y(_0902_),
    .A(_0901_),
    .B(_2920_));
 sg13g2_inv_1 _4764_ (.Y(_0903_),
    .A(_0877_));
 sg13g2_a22oi_1 _4765_ (.Y(_0904_),
    .B1(net127),
    .B2(_0903_),
    .A2(_2658_),
    .A1(_0902_));
 sg13g2_nand3_1 _4766_ (.B(_2878_),
    .C(net115),
    .A(_2441_),
    .Y(_0905_));
 sg13g2_nand2_1 _4767_ (.Y(_0906_),
    .A(_0904_),
    .B(_0905_));
 sg13g2_o21ai_1 _4768_ (.B1(_1991_),
    .Y(_0907_),
    .A1(_0899_),
    .A2(_0906_));
 sg13g2_inv_1 _4769_ (.Y(_0908_),
    .A(_2859_));
 sg13g2_nor2_1 _4770_ (.A(_3045_),
    .B(_0908_),
    .Y(_0909_));
 sg13g2_inv_1 _4771_ (.Y(_0910_),
    .A(_0852_));
 sg13g2_a21oi_1 _4772_ (.A1(_0909_),
    .A2(_0910_),
    .Y(_0912_),
    .B1(net187));
 sg13g2_nand3_1 _4773_ (.B(_0907_),
    .C(_0912_),
    .A(_0897_),
    .Y(_0913_));
 sg13g2_nor2_2 _4774_ (.A(_2560_),
    .B(_3024_),
    .Y(_0914_));
 sg13g2_o21ai_1 _4775_ (.B1(net134),
    .Y(_0915_),
    .A1(_0914_),
    .A2(_0879_));
 sg13g2_nor2_1 _4776_ (.A(_1140_),
    .B(_0149_),
    .Y(_0916_));
 sg13g2_buf_2 _4777_ (.A(_0916_),
    .X(_0917_));
 sg13g2_nor2_1 _4778_ (.A(_0898_),
    .B(_3024_),
    .Y(_0918_));
 sg13g2_o21ai_1 _4779_ (.B1(_0918_),
    .Y(_0919_),
    .A1(net90),
    .A2(_0917_));
 sg13g2_a21oi_1 _4780_ (.A1(_0915_),
    .A2(_0919_),
    .Y(_0920_),
    .B1(net150));
 sg13g2_nand3_1 _4781_ (.B(net48),
    .C(_0847_),
    .A(_0233_),
    .Y(_0921_));
 sg13g2_a21oi_1 _4782_ (.A1(_2662_),
    .A2(net213),
    .Y(_0923_),
    .B1(_2998_));
 sg13g2_o21ai_1 _4783_ (.B1(net189),
    .Y(_0924_),
    .A1(net129),
    .A2(net121));
 sg13g2_nand2b_1 _4784_ (.Y(_0925_),
    .B(_0924_),
    .A_N(_0923_));
 sg13g2_a22oi_1 _4785_ (.Y(_0926_),
    .B1(_2361_),
    .B2(_0925_),
    .A2(net167),
    .A1(_0921_));
 sg13g2_nand3b_1 _4786_ (.B(net138),
    .C(_0926_),
    .Y(_0927_),
    .A_N(_0920_));
 sg13g2_nand2_1 _4787_ (.Y(_0928_),
    .A(_0913_),
    .B(_0927_));
 sg13g2_nand2_1 _4788_ (.Y(_0929_),
    .A(_0928_),
    .B(net194));
 sg13g2_nor2_1 _4789_ (.A(_2165_),
    .B(_0902_),
    .Y(_0930_));
 sg13g2_nor2_1 _4790_ (.A(_2421_),
    .B(_0930_),
    .Y(_0931_));
 sg13g2_o21ai_1 _4791_ (.B1(_0931_),
    .Y(_0932_),
    .A1(_3015_),
    .A2(_0513_));
 sg13g2_nand2_1 _4792_ (.Y(_0934_),
    .A(_3032_),
    .B(_3002_));
 sg13g2_inv_1 _4793_ (.Y(_0935_),
    .A(_0149_));
 sg13g2_nand2_1 _4794_ (.Y(_0936_),
    .A(_2175_),
    .B(_0935_));
 sg13g2_nand3_1 _4795_ (.B(net116),
    .C(_0936_),
    .A(_0934_),
    .Y(_0937_));
 sg13g2_nor2b_1 _4796_ (.A(net141),
    .B_N(_0937_),
    .Y(_0938_));
 sg13g2_nand2_1 _4797_ (.Y(_0939_),
    .A(_2768_),
    .B(_1708_));
 sg13g2_nor2_2 _4798_ (.A(_3001_),
    .B(_0939_),
    .Y(_0940_));
 sg13g2_nor2_1 _4799_ (.A(net60),
    .B(_0940_),
    .Y(_0941_));
 sg13g2_nand3_1 _4800_ (.B(net185),
    .C(_0936_),
    .A(_0875_),
    .Y(_0942_));
 sg13g2_inv_1 _4801_ (.Y(_0943_),
    .A(_0866_));
 sg13g2_a21oi_1 _4802_ (.A1(_0943_),
    .A2(net149),
    .Y(_0945_),
    .B1(net203));
 sg13g2_nand2_1 _4803_ (.Y(_0946_),
    .A(_0942_),
    .B(_0945_));
 sg13g2_o21ai_1 _4804_ (.B1(net199),
    .Y(_0947_),
    .A1(_0941_),
    .A2(_0946_));
 sg13g2_a21oi_1 _4805_ (.A1(_0932_),
    .A2(_0938_),
    .Y(_0948_),
    .B1(_0947_));
 sg13g2_nor3_1 _4806_ (.A(_2479_),
    .B(_3004_),
    .C(net106),
    .Y(_0949_));
 sg13g2_nand2_1 _4807_ (.Y(_0950_),
    .A(_2713_),
    .B(_1108_));
 sg13g2_a21oi_1 _4808_ (.A1(_0950_),
    .A2(_0367_),
    .Y(_0951_),
    .B1(net80));
 sg13g2_inv_1 _4809_ (.Y(_0952_),
    .A(_2622_));
 sg13g2_nand2_1 _4810_ (.Y(_0953_),
    .A(net220),
    .B(net226));
 sg13g2_inv_1 _4811_ (.Y(_0954_),
    .A(_0953_));
 sg13g2_a21oi_1 _4812_ (.A1(_0952_),
    .A2(net163),
    .Y(_0956_),
    .B1(_0954_));
 sg13g2_nand2b_1 _4813_ (.Y(_0957_),
    .B(_0956_),
    .A_N(_0951_));
 sg13g2_o21ai_1 _4814_ (.B1(net140),
    .Y(_0958_),
    .A1(_0949_),
    .A2(_0957_));
 sg13g2_o21ai_1 _4815_ (.B1(_0931_),
    .Y(_0959_),
    .A1(_2693_),
    .A2(_0848_));
 sg13g2_nor2_1 _4816_ (.A(_3004_),
    .B(_0901_),
    .Y(_0960_));
 sg13g2_a22oi_1 _4817_ (.Y(_0961_),
    .B1(net99),
    .B2(_0960_),
    .A2(net114),
    .A1(_0943_));
 sg13g2_nand2_1 _4818_ (.Y(_0962_),
    .A(_0959_),
    .B(_0961_));
 sg13g2_nand2_1 _4819_ (.Y(_0963_),
    .A(_0962_),
    .B(_0351_));
 sg13g2_nand2_1 _4820_ (.Y(_0964_),
    .A(_0958_),
    .B(_0963_));
 sg13g2_nor3_1 _4821_ (.A(net183),
    .B(_0948_),
    .C(_0964_),
    .Y(_0965_));
 sg13g2_nor2_1 _4822_ (.A(_2639_),
    .B(_0965_),
    .Y(_0967_));
 sg13g2_nand2_1 _4823_ (.Y(_0968_),
    .A(_0929_),
    .B(_0967_));
 sg13g2_nand2_1 _4824_ (.Y(_0025_),
    .A(_0890_),
    .B(_0968_));
 sg13g2_a21oi_1 _4825_ (.A1(_2932_),
    .A2(net39),
    .Y(_0969_),
    .B1(_3051_));
 sg13g2_a21oi_1 _4826_ (.A1(_0847_),
    .A2(_0790_),
    .Y(_0970_),
    .B1(_0482_));
 sg13g2_nor2_1 _4827_ (.A(_2391_),
    .B(_2437_),
    .Y(_0971_));
 sg13g2_inv_1 _4828_ (.Y(_0972_),
    .A(_0971_));
 sg13g2_nand3_1 _4829_ (.B(_0197_),
    .C(_0972_),
    .A(_0201_),
    .Y(_0973_));
 sg13g2_a22oi_1 _4830_ (.Y(_0974_),
    .B1(_0970_),
    .B2(_0973_),
    .A2(_0139_),
    .A1(_2423_));
 sg13g2_o21ai_1 _4831_ (.B1(_0974_),
    .Y(_0975_),
    .A1(net43),
    .A2(_0969_));
 sg13g2_nor2_1 _4832_ (.A(net197),
    .B(_2556_),
    .Y(_0977_));
 sg13g2_o21ai_1 _4833_ (.B1(_0977_),
    .Y(_0978_),
    .A1(net39),
    .A2(_2942_));
 sg13g2_a21oi_1 _4834_ (.A1(_0184_),
    .A2(_0095_),
    .Y(_0979_),
    .B1(_0550_));
 sg13g2_nand2_1 _4835_ (.Y(_0980_),
    .A(_0978_),
    .B(_0979_));
 sg13g2_a21oi_1 _4836_ (.A1(net101),
    .A2(net221),
    .Y(_0981_),
    .B1(net153));
 sg13g2_nand2_1 _4837_ (.Y(_0982_),
    .A(_0939_),
    .B(_0981_));
 sg13g2_nor2_1 _4838_ (.A(net116),
    .B(_2417_),
    .Y(_0983_));
 sg13g2_nand4_1 _4839_ (.B(_0982_),
    .C(_0295_),
    .A(_0803_),
    .Y(_0984_),
    .D(_0983_));
 sg13g2_nand3_1 _4840_ (.B(_0984_),
    .C(net218),
    .A(_0980_),
    .Y(_0985_));
 sg13g2_a21oi_1 _4841_ (.A1(_0975_),
    .A2(net87),
    .Y(_0986_),
    .B1(_0985_));
 sg13g2_a21oi_1 _4842_ (.A1(_2506_),
    .A2(_2897_),
    .Y(_0988_),
    .B1(_3023_));
 sg13g2_nand2_1 _4843_ (.Y(_0989_),
    .A(net117),
    .B(net66));
 sg13g2_o21ai_1 _4844_ (.B1(_0989_),
    .Y(_0990_),
    .A1(net63),
    .A2(_0988_));
 sg13g2_nand2_1 _4845_ (.Y(_0991_),
    .A(_0990_),
    .B(net133));
 sg13g2_nor2_2 _4846_ (.A(net170),
    .B(_1512_),
    .Y(_0992_));
 sg13g2_o21ai_1 _4847_ (.B1(_0788_),
    .Y(_0993_),
    .A1(_2557_),
    .A2(_0992_));
 sg13g2_nand2_1 _4848_ (.Y(_0994_),
    .A(_0232_),
    .B(net51));
 sg13g2_nand3_1 _4849_ (.B(net76),
    .C(_0259_),
    .A(_0994_),
    .Y(_0995_));
 sg13g2_nand3_1 _4850_ (.B(_0995_),
    .C(net171),
    .A(_0993_),
    .Y(_0996_));
 sg13g2_a21o_1 _4851_ (.A2(_0996_),
    .A1(_0991_),
    .B1(net138),
    .X(_0997_));
 sg13g2_a21oi_1 _4852_ (.A1(_2884_),
    .A2(net74),
    .Y(_0999_),
    .B1(net148));
 sg13g2_a21oi_1 _4853_ (.A1(_0999_),
    .A2(_0847_),
    .Y(_1000_),
    .B1(net50));
 sg13g2_nand2_1 _4854_ (.Y(_1001_),
    .A(_0164_),
    .B(_2714_));
 sg13g2_nand2_1 _4855_ (.Y(_1002_),
    .A(_0546_),
    .B(_1001_));
 sg13g2_nand2_1 _4856_ (.Y(_1003_),
    .A(_1000_),
    .B(_1002_));
 sg13g2_nand2_1 _4857_ (.Y(_1004_),
    .A(_2569_),
    .B(net104));
 sg13g2_nand2_1 _4858_ (.Y(_1005_),
    .A(_1004_),
    .B(_2805_));
 sg13g2_nand2_1 _4859_ (.Y(_1006_),
    .A(_1005_),
    .B(_2723_));
 sg13g2_nand3_1 _4860_ (.B(net105),
    .C(net75),
    .A(_1006_),
    .Y(_1007_));
 sg13g2_nand3_1 _4861_ (.B(_3033_),
    .C(net52),
    .A(_3038_),
    .Y(_1008_));
 sg13g2_nand3_1 _4862_ (.B(_1007_),
    .C(_1008_),
    .A(_1003_),
    .Y(_1010_));
 sg13g2_nor2_1 _4863_ (.A(net214),
    .B(net216),
    .Y(_1011_));
 sg13g2_nand2_1 _4864_ (.Y(_1012_),
    .A(_1010_),
    .B(_1011_));
 sg13g2_nand3_1 _4865_ (.B(_0997_),
    .C(_1012_),
    .A(_0986_),
    .Y(_1013_));
 sg13g2_nor2_1 _4866_ (.A(net60),
    .B(_2872_),
    .Y(_1014_));
 sg13g2_nor2_2 _4867_ (.A(_1162_),
    .B(_0866_),
    .Y(_1015_));
 sg13g2_nor2_1 _4868_ (.A(_0281_),
    .B(_0301_),
    .Y(_1016_));
 sg13g2_a221oi_1 _4869_ (.B2(_1741_),
    .C1(_1016_),
    .B1(_1015_),
    .A1(_1014_),
    .Y(_1017_),
    .A2(_2885_));
 sg13g2_a21oi_1 _4870_ (.A1(_1017_),
    .A2(net55),
    .Y(_1018_),
    .B1(net186));
 sg13g2_a21oi_1 _4871_ (.A1(_2569_),
    .A2(net121),
    .Y(_1019_),
    .B1(_2686_));
 sg13g2_a21oi_1 _4872_ (.A1(_2687_),
    .A2(_1828_),
    .Y(_1021_),
    .B1(net112));
 sg13g2_a21oi_1 _4873_ (.A1(_2679_),
    .A2(_0847_),
    .Y(_1022_),
    .B1(_1468_));
 sg13g2_nor4_1 _4874_ (.A(net145),
    .B(_1019_),
    .C(_1021_),
    .D(_1022_),
    .Y(_1023_));
 sg13g2_a21o_1 _4875_ (.A2(_3038_),
    .A1(_0135_),
    .B1(net100),
    .X(_1024_));
 sg13g2_o21ai_1 _4876_ (.B1(net62),
    .Y(_1025_),
    .A1(_1730_),
    .A2(_0123_));
 sg13g2_nand3_1 _4877_ (.B(_1024_),
    .C(_1025_),
    .A(_1023_),
    .Y(_1026_));
 sg13g2_nand2_1 _4878_ (.Y(_1027_),
    .A(_1018_),
    .B(_1026_));
 sg13g2_nand2_2 _4879_ (.Y(_1028_),
    .A(_0992_),
    .B(net169));
 sg13g2_nand2_1 _4880_ (.Y(_1029_),
    .A(_1028_),
    .B(_2915_));
 sg13g2_a21oi_1 _4881_ (.A1(_2490_),
    .A2(_0524_),
    .Y(_1030_),
    .B1(_0260_));
 sg13g2_o21ai_1 _4882_ (.B1(_1030_),
    .Y(_1032_),
    .A1(_2763_),
    .A2(_1029_));
 sg13g2_a21oi_1 _4883_ (.A1(_2725_),
    .A2(_2618_),
    .Y(_1033_),
    .B1(net84));
 sg13g2_nand2_2 _4884_ (.Y(_1034_),
    .A(_0773_),
    .B(_2568_));
 sg13g2_nor2_1 _4885_ (.A(net91),
    .B(_2914_),
    .Y(_1035_));
 sg13g2_nand2_1 _4886_ (.Y(_1036_),
    .A(_1034_),
    .B(_1035_));
 sg13g2_nand2_1 _4887_ (.Y(_1037_),
    .A(_1033_),
    .B(_1036_));
 sg13g2_a21oi_1 _4888_ (.A1(_1032_),
    .A2(_1037_),
    .Y(_1038_),
    .B1(net161));
 sg13g2_nor2_1 _4889_ (.A(_2425_),
    .B(_2289_),
    .Y(_1039_));
 sg13g2_inv_1 _4890_ (.Y(_1040_),
    .A(_1039_));
 sg13g2_nand2_1 _4891_ (.Y(_1041_),
    .A(_1034_),
    .B(_1040_));
 sg13g2_a21oi_1 _4892_ (.A1(_1041_),
    .A2(_0151_),
    .Y(_1043_),
    .B1(_2516_));
 sg13g2_nor2b_1 _4893_ (.A(_1038_),
    .B_N(_1043_),
    .Y(_1044_));
 sg13g2_a21oi_1 _4894_ (.A1(_1027_),
    .A2(_1044_),
    .Y(_1045_),
    .B1(net182));
 sg13g2_nand2_1 _4895_ (.Y(_1046_),
    .A(_1013_),
    .B(_1045_));
 sg13g2_a21oi_1 _4896_ (.A1(_0950_),
    .A2(_0342_),
    .Y(_1047_),
    .B1(net112));
 sg13g2_a21oi_1 _4897_ (.A1(_1034_),
    .A2(_3028_),
    .Y(_1048_),
    .B1(_2705_));
 sg13g2_inv_1 _4898_ (.Y(_1049_),
    .A(_0869_));
 sg13g2_a21oi_1 _4899_ (.A1(_0764_),
    .A2(_1049_),
    .Y(_1050_),
    .B1(_2931_));
 sg13g2_nor3_1 _4900_ (.A(_1047_),
    .B(_1048_),
    .C(_1050_),
    .Y(_1051_));
 sg13g2_a21oi_1 _4901_ (.A1(_1051_),
    .A2(net156),
    .Y(_1052_),
    .B1(net143));
 sg13g2_nor3_1 _4902_ (.A(_1730_),
    .B(_2857_),
    .C(_0123_),
    .Y(_1054_));
 sg13g2_a21oi_1 _4903_ (.A1(_0498_),
    .A2(_0818_),
    .Y(_1055_),
    .B1(_1054_));
 sg13g2_a21oi_1 _4904_ (.A1(_1055_),
    .A2(_0194_),
    .Y(_1056_),
    .B1(net133));
 sg13g2_a21oi_1 _4905_ (.A1(_0135_),
    .A2(_0527_),
    .Y(_1057_),
    .B1(net88));
 sg13g2_a21oi_1 _4906_ (.A1(_0687_),
    .A2(_2856_),
    .Y(_1058_),
    .B1(net48));
 sg13g2_o21ai_1 _4907_ (.B1(_0297_),
    .Y(_1059_),
    .A1(_1057_),
    .A2(_1058_));
 sg13g2_nand2_1 _4908_ (.Y(_1060_),
    .A(_1056_),
    .B(_1059_));
 sg13g2_nand2_1 _4909_ (.Y(_1061_),
    .A(_1052_),
    .B(_1060_));
 sg13g2_nand2_1 _4910_ (.Y(_1062_),
    .A(_0773_),
    .B(net91));
 sg13g2_nand2_1 _4911_ (.Y(_1063_),
    .A(_2566_),
    .B(_2920_));
 sg13g2_a21oi_1 _4912_ (.A1(_0577_),
    .A2(net88),
    .Y(_1065_),
    .B1(_1063_));
 sg13g2_inv_1 _4913_ (.Y(_1066_),
    .A(_3015_));
 sg13g2_a21oi_1 _4914_ (.A1(_3049_),
    .A2(_1066_),
    .Y(_1067_),
    .B1(net75));
 sg13g2_a21o_1 _4915_ (.A2(_3028_),
    .A1(_1034_),
    .B1(net76),
    .X(_1068_));
 sg13g2_a22oi_1 _4916_ (.Y(_1069_),
    .B1(_1067_),
    .B2(_1068_),
    .A2(_1065_),
    .A1(_1062_));
 sg13g2_nand2_1 _4917_ (.Y(_1070_),
    .A(_2743_),
    .B(net57));
 sg13g2_nand3_1 _4918_ (.B(net54),
    .C(_1413_),
    .A(_1070_),
    .Y(_1071_));
 sg13g2_nor2_1 _4919_ (.A(net111),
    .B(_0137_),
    .Y(_1072_));
 sg13g2_nand2_1 _4920_ (.Y(_1073_),
    .A(net149),
    .B(_0763_));
 sg13g2_inv_1 _4921_ (.Y(_1074_),
    .A(_1073_));
 sg13g2_a22oi_1 _4922_ (.Y(_1076_),
    .B1(_1074_),
    .B2(_2484_),
    .A2(_0972_),
    .A1(_1072_));
 sg13g2_nor3_1 _4923_ (.A(_2971_),
    .B(net155),
    .C(_2435_),
    .Y(_1077_));
 sg13g2_nand2_1 _4924_ (.Y(_1078_),
    .A(_1077_),
    .B(_0527_));
 sg13g2_nand3_1 _4925_ (.B(_1076_),
    .C(_1078_),
    .A(_1071_),
    .Y(_1079_));
 sg13g2_a21oi_1 _4926_ (.A1(_1079_),
    .A2(net156),
    .Y(_1080_),
    .B1(_3044_));
 sg13g2_o21ai_1 _4927_ (.B1(_1080_),
    .Y(_1081_),
    .A1(net156),
    .A2(_1069_));
 sg13g2_nand3_1 _4928_ (.B(_1081_),
    .C(net190),
    .A(_1061_),
    .Y(_1082_));
 sg13g2_a21oi_1 _4929_ (.A1(_1005_),
    .A2(_0822_),
    .Y(_1083_),
    .B1(net63));
 sg13g2_nand2_1 _4930_ (.Y(_1084_),
    .A(_0645_),
    .B(_1015_));
 sg13g2_nand3_1 _4931_ (.B(_2463_),
    .C(_0175_),
    .A(_1001_),
    .Y(_1085_));
 sg13g2_o21ai_1 _4932_ (.B1(_2659_),
    .Y(_1087_),
    .A1(_2681_),
    .A2(_2489_));
 sg13g2_nand4_1 _4933_ (.B(_1085_),
    .C(_2412_),
    .A(_1084_),
    .Y(_1088_),
    .D(_1087_));
 sg13g2_nor2_1 _4934_ (.A(_1083_),
    .B(_1088_),
    .Y(_1089_));
 sg13g2_nand2_1 _4935_ (.Y(_1090_),
    .A(_0211_),
    .B(net195));
 sg13g2_nor2_1 _4936_ (.A(net101),
    .B(_1004_),
    .Y(_1091_));
 sg13g2_nor3_1 _4937_ (.A(net185),
    .B(_1090_),
    .C(_1091_),
    .Y(_1092_));
 sg13g2_o21ai_1 _4938_ (.B1(_1893_),
    .Y(_1093_),
    .A1(net170),
    .A2(_2439_));
 sg13g2_nand2_1 _4939_ (.Y(_1094_),
    .A(_1093_),
    .B(net216));
 sg13g2_a21oi_1 _4940_ (.A1(_1031_),
    .A2(net221),
    .Y(_1095_),
    .B1(_2581_));
 sg13g2_a21oi_1 _4941_ (.A1(net51),
    .A2(_1095_),
    .Y(_1096_),
    .B1(_0827_));
 sg13g2_nor2_1 _4942_ (.A(_1094_),
    .B(_1096_),
    .Y(_1098_));
 sg13g2_nand2_1 _4943_ (.Y(_1099_),
    .A(_2897_),
    .B(net46));
 sg13g2_nand3_1 _4944_ (.B(net102),
    .C(_1099_),
    .A(_1028_),
    .Y(_1100_));
 sg13g2_nand3b_1 _4945_ (.B(_1098_),
    .C(_1100_),
    .Y(_1101_),
    .A_N(_1092_));
 sg13g2_nand2_1 _4946_ (.Y(_1102_),
    .A(_1101_),
    .B(_1991_));
 sg13g2_nor2_1 _4947_ (.A(_1089_),
    .B(_1102_),
    .Y(_1103_));
 sg13g2_o21ai_1 _4948_ (.B1(net216),
    .Y(_1104_),
    .A1(net68),
    .A2(_0168_));
 sg13g2_nand3_1 _4949_ (.B(net163),
    .C(_2726_),
    .A(_1034_),
    .Y(_1105_));
 sg13g2_nand2_1 _4950_ (.Y(_1106_),
    .A(net61),
    .B(net126));
 sg13g2_nand3_1 _4951_ (.B(_1106_),
    .C(net153),
    .A(_0485_),
    .Y(_1107_));
 sg13g2_nand3_1 _4952_ (.B(net191),
    .C(_1107_),
    .A(_1105_),
    .Y(_1109_));
 sg13g2_nand2_1 _4953_ (.Y(_1110_),
    .A(_1020_),
    .B(net124));
 sg13g2_o21ai_1 _4954_ (.B1(_2996_),
    .Y(_1111_),
    .A1(_2523_),
    .A2(_1110_));
 sg13g2_nand2_1 _4955_ (.Y(_1112_),
    .A(_1111_),
    .B(net99));
 sg13g2_nand3b_1 _4956_ (.B(_1109_),
    .C(_1112_),
    .Y(_1113_),
    .A_N(_1104_));
 sg13g2_nor2_1 _4957_ (.A(net177),
    .B(_2973_),
    .Y(_1114_));
 sg13g2_o21ai_1 _4958_ (.B1(net115),
    .Y(_1115_),
    .A1(_2600_),
    .A2(_1114_));
 sg13g2_nand3_1 _4959_ (.B(_2447_),
    .C(_0662_),
    .A(_0688_),
    .Y(_1116_));
 sg13g2_nand2_1 _4960_ (.Y(_1117_),
    .A(_1115_),
    .B(_1116_));
 sg13g2_nand3_1 _4961_ (.B(_1785_),
    .C(_1741_),
    .A(_0265_),
    .Y(_1118_));
 sg13g2_nand3_1 _4962_ (.B(net118),
    .C(_1435_),
    .A(_2986_),
    .Y(_1120_));
 sg13g2_a21oi_1 _4963_ (.A1(_1675_),
    .A2(_1435_),
    .Y(_1121_),
    .B1(_2411_));
 sg13g2_nand3_1 _4964_ (.B(_1120_),
    .C(_1121_),
    .A(_1118_),
    .Y(_1122_));
 sg13g2_nor2_1 _4965_ (.A(_1117_),
    .B(_1122_),
    .Y(_1123_));
 sg13g2_nor2_1 _4966_ (.A(net145),
    .B(_1123_),
    .Y(_1124_));
 sg13g2_nand2_1 _4967_ (.Y(_1125_),
    .A(_1113_),
    .B(_1124_));
 sg13g2_nand2_1 _4968_ (.Y(_1126_),
    .A(_1125_),
    .B(net183));
 sg13g2_nor2_1 _4969_ (.A(_1103_),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_nor2_1 _4970_ (.A(_2639_),
    .B(_1127_),
    .Y(_1128_));
 sg13g2_nand2_1 _4971_ (.Y(_1129_),
    .A(_1082_),
    .B(_1128_));
 sg13g2_nand2_1 _4972_ (.Y(_0026_),
    .A(_1046_),
    .B(_1129_));
 sg13g2_inv_1 _4973_ (.Y(_1131_),
    .A(_0180_));
 sg13g2_a21oi_1 _4974_ (.A1(_3027_),
    .A2(_1131_),
    .Y(_1132_),
    .B1(_0140_));
 sg13g2_a21oi_1 _4975_ (.A1(net41),
    .A2(_2502_),
    .Y(_1133_),
    .B1(net195));
 sg13g2_nand3_1 _4976_ (.B(_0505_),
    .C(_2981_),
    .A(_1133_),
    .Y(_1134_));
 sg13g2_nand2_1 _4977_ (.Y(_1135_),
    .A(_1132_),
    .B(_1134_));
 sg13g2_nand2_1 _4978_ (.Y(_1136_),
    .A(_0437_),
    .B(_2503_));
 sg13g2_nor3_1 _4979_ (.A(net159),
    .B(_0539_),
    .C(_2894_),
    .Y(_1137_));
 sg13g2_a21oi_1 _4980_ (.A1(_1136_),
    .A2(net58),
    .Y(_1138_),
    .B1(_1137_));
 sg13g2_nand2_1 _4981_ (.Y(_1139_),
    .A(_1135_),
    .B(_1138_));
 sg13g2_nand2_1 _4982_ (.Y(_1141_),
    .A(_1139_),
    .B(net140));
 sg13g2_nor2_1 _4983_ (.A(net219),
    .B(_2725_),
    .Y(_1142_));
 sg13g2_nand2b_1 _4984_ (.Y(_1143_),
    .B(_1142_),
    .A_N(_0882_));
 sg13g2_nand2_1 _4985_ (.Y(_1144_),
    .A(_2982_),
    .B(net85));
 sg13g2_nand3_1 _4986_ (.B(_0752_),
    .C(_2429_),
    .A(net82),
    .Y(_1145_));
 sg13g2_nand3_1 _4987_ (.B(_1144_),
    .C(_1145_),
    .A(_1143_),
    .Y(_1146_));
 sg13g2_nand2_1 _4988_ (.Y(_1147_),
    .A(_1146_),
    .B(net86));
 sg13g2_nand2_1 _4989_ (.Y(_1148_),
    .A(_1141_),
    .B(_1147_));
 sg13g2_nand2_1 _4990_ (.Y(_1149_),
    .A(_2117_),
    .B(net168));
 sg13g2_a21oi_1 _4991_ (.A1(_2565_),
    .A2(_1149_),
    .Y(_1150_),
    .B1(net80));
 sg13g2_a21oi_1 _4992_ (.A1(_2969_),
    .A2(_2825_),
    .Y(_1152_),
    .B1(net60));
 sg13g2_o21ai_1 _4993_ (.B1(_0502_),
    .Y(_1153_),
    .A1(net51),
    .A2(_0845_));
 sg13g2_o21ai_1 _4994_ (.B1(net174),
    .Y(_1154_),
    .A1(net112),
    .A2(_1153_));
 sg13g2_nor2_1 _4995_ (.A(net100),
    .B(_0464_),
    .Y(_1155_));
 sg13g2_nor4_1 _4996_ (.A(_1150_),
    .B(_1152_),
    .C(_1154_),
    .D(_1155_),
    .Y(_1156_));
 sg13g2_a21oi_1 _4997_ (.A1(_2577_),
    .A2(net70),
    .Y(_1157_),
    .B1(net197));
 sg13g2_nand2_2 _4998_ (.Y(_1158_),
    .A(_1523_),
    .B(_2502_));
 sg13g2_nand3_1 _4999_ (.B(_0505_),
    .C(_1158_),
    .A(_1157_),
    .Y(_1159_));
 sg13g2_nor2_1 _5000_ (.A(_0501_),
    .B(_0426_),
    .Y(_1160_));
 sg13g2_nor2_1 _5001_ (.A(net158),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_nand2b_1 _5002_ (.Y(_1163_),
    .B(_1161_),
    .A_N(_2929_));
 sg13g2_nand3_1 _5003_ (.B(net109),
    .C(_1163_),
    .A(_1159_),
    .Y(_1164_));
 sg13g2_o21ai_1 _5004_ (.B1(_1119_),
    .Y(_1165_),
    .A1(net41),
    .A2(_2762_));
 sg13g2_inv_1 _5005_ (.Y(_1166_),
    .A(_3016_));
 sg13g2_o21ai_1 _5006_ (.B1(net214),
    .Y(_1167_),
    .A1(_1166_),
    .A2(_2607_));
 sg13g2_a21oi_1 _5007_ (.A1(_1165_),
    .A2(net58),
    .Y(_1168_),
    .B1(_1167_));
 sg13g2_nand2_1 _5008_ (.Y(_1169_),
    .A(_1164_),
    .B(_1168_));
 sg13g2_nand2_1 _5009_ (.Y(_1170_),
    .A(_1169_),
    .B(net151));
 sg13g2_nor2_1 _5010_ (.A(_1156_),
    .B(_1170_),
    .Y(_1171_));
 sg13g2_a21oi_1 _5011_ (.A1(_1148_),
    .A2(net188),
    .Y(_1172_),
    .B1(_1171_));
 sg13g2_nand2_1 _5012_ (.Y(_1174_),
    .A(_2621_),
    .B(net162));
 sg13g2_o21ai_1 _5013_ (.B1(_1174_),
    .Y(_1175_),
    .A1(_2035_),
    .A2(net204));
 sg13g2_nand2_1 _5014_ (.Y(_1176_),
    .A(_1175_),
    .B(net164));
 sg13g2_nand2_1 _5015_ (.Y(_1177_),
    .A(_1176_),
    .B(_2526_));
 sg13g2_nor2_1 _5016_ (.A(net148),
    .B(_0427_),
    .Y(_1178_));
 sg13g2_nand2_1 _5017_ (.Y(_1179_),
    .A(_2499_),
    .B(_1178_));
 sg13g2_nand2_1 _5018_ (.Y(_1180_),
    .A(_1177_),
    .B(_1179_));
 sg13g2_nand2_1 _5019_ (.Y(_1181_),
    .A(_0388_),
    .B(_2425_));
 sg13g2_nand2_1 _5020_ (.Y(_1182_),
    .A(_0331_),
    .B(_1181_));
 sg13g2_nand2_1 _5021_ (.Y(_1183_),
    .A(_1182_),
    .B(net66));
 sg13g2_nand2_1 _5022_ (.Y(_1185_),
    .A(_0635_),
    .B(net107));
 sg13g2_o21ai_1 _5023_ (.B1(net214),
    .Y(_1186_),
    .A1(net159),
    .A2(_2618_));
 sg13g2_a21oi_1 _5024_ (.A1(_2735_),
    .A2(_1185_),
    .Y(_1187_),
    .B1(_1186_));
 sg13g2_nand3_1 _5025_ (.B(_1183_),
    .C(_1187_),
    .A(_1180_),
    .Y(_1188_));
 sg13g2_a21oi_1 _5026_ (.A1(_0300_),
    .A2(_3017_),
    .Y(_1189_),
    .B1(net155));
 sg13g2_o21ai_1 _5027_ (.B1(_2875_),
    .Y(_1190_),
    .A1(net51),
    .A2(_2742_));
 sg13g2_nand2_1 _5028_ (.Y(_1191_),
    .A(_1189_),
    .B(_1190_));
 sg13g2_nand2_1 _5029_ (.Y(_1192_),
    .A(_2692_),
    .B(_2769_));
 sg13g2_inv_1 _5030_ (.Y(_1193_),
    .A(_2723_));
 sg13g2_nand2_2 _5031_ (.Y(_1194_),
    .A(_1193_),
    .B(_1435_));
 sg13g2_nand2_2 _5032_ (.Y(_1196_),
    .A(_1194_),
    .B(net203));
 sg13g2_a21oi_1 _5033_ (.A1(_1192_),
    .A2(_0203_),
    .Y(_1197_),
    .B1(_1196_));
 sg13g2_a21oi_1 _5034_ (.A1(_1191_),
    .A2(_1197_),
    .Y(_1198_),
    .B1(_2413_));
 sg13g2_nand2_1 _5035_ (.Y(_1199_),
    .A(_1188_),
    .B(_1198_));
 sg13g2_o21ai_1 _5036_ (.B1(_0677_),
    .Y(_1200_),
    .A1(net51),
    .A2(_0680_));
 sg13g2_a21oi_1 _5037_ (.A1(_0497_),
    .A2(_0346_),
    .Y(_1201_),
    .B1(_2550_));
 sg13g2_nand2_1 _5038_ (.Y(_1202_),
    .A(_1200_),
    .B(_1201_));
 sg13g2_nor2_1 _5039_ (.A(_2568_),
    .B(_3001_),
    .Y(_1203_));
 sg13g2_nor3_1 _5040_ (.A(net128),
    .B(_1203_),
    .C(_0852_),
    .Y(_1204_));
 sg13g2_nor2_1 _5041_ (.A(_2491_),
    .B(_0750_),
    .Y(_1205_));
 sg13g2_a21oi_1 _5042_ (.A1(_2621_),
    .A2(_1205_),
    .Y(_1207_),
    .B1(net217));
 sg13g2_nor2b_1 _5043_ (.A(_1204_),
    .B_N(_1207_),
    .Y(_1208_));
 sg13g2_a21oi_1 _5044_ (.A1(_1202_),
    .A2(_1208_),
    .Y(_1209_),
    .B1(net216));
 sg13g2_nor2_1 _5045_ (.A(_1042_),
    .B(_2968_),
    .Y(_1210_));
 sg13g2_a21oi_1 _5046_ (.A1(_1210_),
    .A2(_2703_),
    .Y(_1211_),
    .B1(_2487_));
 sg13g2_nand2_1 _5047_ (.Y(_1212_),
    .A(_2473_),
    .B(_1211_));
 sg13g2_nand2_1 _5048_ (.Y(_1213_),
    .A(_1066_),
    .B(_3014_));
 sg13g2_nand2_1 _5049_ (.Y(_1214_),
    .A(_1212_),
    .B(_1213_));
 sg13g2_nand2_1 _5050_ (.Y(_1215_),
    .A(_1214_),
    .B(_2566_));
 sg13g2_a21oi_1 _5051_ (.A1(_0407_),
    .A2(_2397_),
    .Y(_1216_),
    .B1(net159));
 sg13g2_nor3_1 _5052_ (.A(net226),
    .B(_1162_),
    .C(_2800_),
    .Y(_1218_));
 sg13g2_nor3_1 _5053_ (.A(_1981_),
    .B(_1216_),
    .C(_1218_),
    .Y(_1219_));
 sg13g2_nand2_1 _5054_ (.Y(_1220_),
    .A(_1215_),
    .B(_1219_));
 sg13g2_nand2_1 _5055_ (.Y(_1221_),
    .A(_1209_),
    .B(_1220_));
 sg13g2_nand2_1 _5056_ (.Y(_1222_),
    .A(_1199_),
    .B(_1221_));
 sg13g2_nand2_1 _5057_ (.Y(_1223_),
    .A(_1222_),
    .B(net183));
 sg13g2_nand2_1 _5058_ (.Y(_1224_),
    .A(_1172_),
    .B(_1223_));
 sg13g2_nand2_1 _5059_ (.Y(_1225_),
    .A(_1224_),
    .B(net182));
 sg13g2_and3_1 _5060_ (.X(_1226_),
    .A(_0314_),
    .B(net76),
    .C(_2618_));
 sg13g2_a21o_1 _5061_ (.A2(net147),
    .A1(_3048_),
    .B1(net136),
    .X(_1227_));
 sg13g2_nand2_1 _5062_ (.Y(_1229_),
    .A(_0635_),
    .B(net61));
 sg13g2_nand2_1 _5063_ (.Y(_1230_),
    .A(_1229_),
    .B(_0807_));
 sg13g2_nor2_1 _5064_ (.A(net147),
    .B(net177),
    .Y(_1231_));
 sg13g2_nand2b_1 _5065_ (.Y(_1232_),
    .B(_0505_),
    .A_N(_1231_));
 sg13g2_a22oi_1 _5066_ (.Y(_1233_),
    .B1(net47),
    .B2(_1232_),
    .A2(net40),
    .A1(_1230_));
 sg13g2_o21ai_1 _5067_ (.B1(_1233_),
    .Y(_1234_),
    .A1(_1226_),
    .A2(_1227_));
 sg13g2_a22oi_1 _5068_ (.Y(_1235_),
    .B1(_0977_),
    .B2(_2881_),
    .A2(_0623_),
    .A1(net77));
 sg13g2_o21ai_1 _5069_ (.B1(net188),
    .Y(_1236_),
    .A1(_0550_),
    .A2(_1235_));
 sg13g2_a21oi_1 _5070_ (.A1(_1234_),
    .A2(net87),
    .Y(_1237_),
    .B1(_1236_));
 sg13g2_o21ai_1 _5071_ (.B1(_0430_),
    .Y(_1238_),
    .A1(net39),
    .A2(net70));
 sg13g2_a21oi_1 _5072_ (.A1(_1238_),
    .A2(net52),
    .Y(_1240_),
    .B1(net93));
 sg13g2_nand2_1 _5073_ (.Y(_1241_),
    .A(_2942_),
    .B(net45));
 sg13g2_nand3_1 _5074_ (.B(net48),
    .C(_0211_),
    .A(_1241_),
    .Y(_1242_));
 sg13g2_nand2_1 _5075_ (.Y(_1243_),
    .A(_0901_),
    .B(_0304_));
 sg13g2_nor2_1 _5076_ (.A(net164),
    .B(_0954_),
    .Y(_1244_));
 sg13g2_nand3_1 _5077_ (.B(_1243_),
    .C(_1244_),
    .A(_1242_),
    .Y(_1245_));
 sg13g2_nand2_1 _5078_ (.Y(_1246_),
    .A(_1240_),
    .B(_1245_));
 sg13g2_nand3_1 _5079_ (.B(_0455_),
    .C(_0994_),
    .A(_2586_),
    .Y(_1247_));
 sg13g2_nand2_1 _5080_ (.Y(_1248_),
    .A(_0548_),
    .B(_0813_));
 sg13g2_nand3_1 _5081_ (.B(net49),
    .C(_1248_),
    .A(_1247_),
    .Y(_1249_));
 sg13g2_nor3_2 _5082_ (.A(net198),
    .B(net213),
    .C(_0935_),
    .Y(_1251_));
 sg13g2_a21oi_1 _5083_ (.A1(_0952_),
    .A2(_1251_),
    .Y(_1252_),
    .B1(net150));
 sg13g2_nand2_1 _5084_ (.Y(_1253_),
    .A(_1249_),
    .B(_1252_));
 sg13g2_nand3_1 _5085_ (.B(_1253_),
    .C(net143),
    .A(_1246_),
    .Y(_1254_));
 sg13g2_nand2_1 _5086_ (.Y(_1255_),
    .A(_1237_),
    .B(_1254_));
 sg13g2_nor2b_1 _5087_ (.A(_1029_),
    .B_N(_0517_),
    .Y(_1256_));
 sg13g2_nor2_1 _5088_ (.A(_2853_),
    .B(_2936_),
    .Y(_1257_));
 sg13g2_o21ai_1 _5089_ (.B1(_1257_),
    .Y(_1258_),
    .A1(_0345_),
    .A2(_0344_));
 sg13g2_nor2_2 _5090_ (.A(net124),
    .B(_2686_),
    .Y(_1259_));
 sg13g2_a21oi_1 _5091_ (.A1(_1258_),
    .A2(_2984_),
    .Y(_1260_),
    .B1(_1259_));
 sg13g2_o21ai_1 _5092_ (.B1(_1260_),
    .Y(_1262_),
    .A1(net63),
    .A2(_1256_));
 sg13g2_nor2_1 _5093_ (.A(net112),
    .B(_2653_),
    .Y(_1263_));
 sg13g2_inv_1 _5094_ (.Y(_1264_),
    .A(_1114_));
 sg13g2_a22oi_1 _5095_ (.Y(_1265_),
    .B1(_1015_),
    .B2(_1264_),
    .A2(_0744_),
    .A1(_1263_));
 sg13g2_nand2_1 _5096_ (.Y(_1266_),
    .A(_0744_),
    .B(_0840_));
 sg13g2_inv_2 _5097_ (.Y(_1267_),
    .A(_0917_));
 sg13g2_nor2_1 _5098_ (.A(_2417_),
    .B(_1267_),
    .Y(_1268_));
 sg13g2_a21oi_1 _5099_ (.A1(_1266_),
    .A2(_1268_),
    .Y(_1269_),
    .B1(net215));
 sg13g2_o21ai_1 _5100_ (.B1(_1269_),
    .Y(_1270_),
    .A1(net165),
    .A2(_1265_));
 sg13g2_a21oi_1 _5101_ (.A1(_1262_),
    .A2(net87),
    .Y(_1271_),
    .B1(_1270_));
 sg13g2_a21oi_1 _5102_ (.A1(_1175_),
    .A2(net50),
    .Y(_1273_),
    .B1(net53));
 sg13g2_o21ai_1 _5103_ (.B1(_0774_),
    .Y(_1274_),
    .A1(_0426_),
    .A2(net106));
 sg13g2_nor2_2 _5104_ (.A(_0149_),
    .B(net198),
    .Y(_1275_));
 sg13g2_a21oi_1 _5105_ (.A1(_1274_),
    .A2(_1275_),
    .Y(_1276_),
    .B1(net150));
 sg13g2_o21ai_1 _5106_ (.B1(_1276_),
    .Y(_1277_),
    .A1(_0869_),
    .A2(_1273_));
 sg13g2_a21oi_1 _5107_ (.A1(net71),
    .A2(_0460_),
    .Y(_1278_),
    .B1(_0411_));
 sg13g2_nor3_1 _5108_ (.A(net109),
    .B(_3004_),
    .C(_1062_),
    .Y(_1279_));
 sg13g2_nand2_1 _5109_ (.Y(_1280_),
    .A(_2689_),
    .B(_1719_));
 sg13g2_a22oi_1 _5110_ (.Y(_1281_),
    .B1(_2659_),
    .B2(_2941_),
    .A2(_1280_),
    .A1(net114));
 sg13g2_nand2_1 _5111_ (.Y(_1282_),
    .A(_1281_),
    .B(net193));
 sg13g2_nor2_1 _5112_ (.A(_1279_),
    .B(_1282_),
    .Y(_1284_));
 sg13g2_o21ai_1 _5113_ (.B1(_1284_),
    .Y(_1285_),
    .A1(net100),
    .A2(_1278_));
 sg13g2_nand3_1 _5114_ (.B(_1285_),
    .C(net143),
    .A(_1277_),
    .Y(_1286_));
 sg13g2_nand2_1 _5115_ (.Y(_1287_),
    .A(_1271_),
    .B(_1286_));
 sg13g2_nand3_1 _5116_ (.B(_1287_),
    .C(net212),
    .A(_1255_),
    .Y(_1288_));
 sg13g2_nand2_1 _5117_ (.Y(_0027_),
    .A(_1225_),
    .B(_1288_));
 sg13g2_nand2_1 _5118_ (.Y(_1289_),
    .A(_0205_),
    .B(_2937_));
 sg13g2_nand2_1 _5119_ (.Y(_1290_),
    .A(_2495_),
    .B(net104));
 sg13g2_nand2b_1 _5120_ (.Y(_1291_),
    .B(_0220_),
    .A_N(_2831_));
 sg13g2_a21oi_1 _5121_ (.A1(net77),
    .A2(_1290_),
    .Y(_1292_),
    .B1(_1291_));
 sg13g2_a21oi_1 _5122_ (.A1(net41),
    .A2(net72),
    .Y(_1294_),
    .B1(_2667_));
 sg13g2_nand3_1 _5123_ (.B(net152),
    .C(_2876_),
    .A(_1294_),
    .Y(_1295_));
 sg13g2_nand3_1 _5124_ (.B(_0482_),
    .C(_2542_),
    .A(_1264_),
    .Y(_1296_));
 sg13g2_nand3_1 _5125_ (.B(_2588_),
    .C(_1296_),
    .A(_1295_),
    .Y(_1297_));
 sg13g2_o21ai_1 _5126_ (.B1(_1297_),
    .Y(_1298_),
    .A1(_2405_),
    .A2(_1292_));
 sg13g2_a22oi_1 _5127_ (.Y(_1299_),
    .B1(net138),
    .B2(_1298_),
    .A2(_1289_),
    .A1(_1268_));
 sg13g2_a21oi_1 _5128_ (.A1(_0177_),
    .A2(_1174_),
    .Y(_1300_),
    .B1(net43));
 sg13g2_inv_1 _5129_ (.Y(_1301_),
    .A(_1275_));
 sg13g2_a21oi_1 _5130_ (.A1(_2777_),
    .A2(_2766_),
    .Y(_1302_),
    .B1(_1301_));
 sg13g2_nor3_1 _5131_ (.A(_1196_),
    .B(_1300_),
    .C(_1302_),
    .Y(_1303_));
 sg13g2_a21oi_1 _5132_ (.A1(_0661_),
    .A2(_2967_),
    .Y(_1305_),
    .B1(net134));
 sg13g2_nand2_1 _5133_ (.Y(_1306_),
    .A(_1861_),
    .B(_3048_));
 sg13g2_nand2_1 _5134_ (.Y(_1307_),
    .A(_1305_),
    .B(_1306_));
 sg13g2_inv_1 _5135_ (.Y(_1308_),
    .A(_2613_));
 sg13g2_nand2_1 _5136_ (.Y(_1309_),
    .A(_1308_),
    .B(_0191_));
 sg13g2_nand3_1 _5137_ (.B(_2522_),
    .C(_2537_),
    .A(_1309_),
    .Y(_1310_));
 sg13g2_o21ai_1 _5138_ (.B1(net47),
    .Y(_1311_),
    .A1(_1882_),
    .A2(_1039_));
 sg13g2_nand4_1 _5139_ (.B(net133),
    .C(_1310_),
    .A(_1307_),
    .Y(_1312_),
    .D(_1311_));
 sg13g2_nand3b_1 _5140_ (.B(_1312_),
    .C(net166),
    .Y(_1313_),
    .A_N(_1303_));
 sg13g2_nand3_1 _5141_ (.B(_1313_),
    .C(_2517_),
    .A(_1299_),
    .Y(_1314_));
 sg13g2_a21oi_1 _5142_ (.A1(net124),
    .A2(_2318_),
    .Y(_1316_),
    .B1(net59));
 sg13g2_nand3_1 _5143_ (.B(_2719_),
    .C(net185),
    .A(_2963_),
    .Y(_1317_));
 sg13g2_nand2_1 _5144_ (.Y(_1318_),
    .A(_1317_),
    .B(net100));
 sg13g2_o21ai_1 _5145_ (.B1(_1318_),
    .Y(_1319_),
    .A1(_0107_),
    .A2(_1316_));
 sg13g2_nand2_1 _5146_ (.Y(_1320_),
    .A(_1319_),
    .B(_0119_));
 sg13g2_o21ai_1 _5147_ (.B1(net174),
    .Y(_1321_),
    .A1(_2519_),
    .A2(_2686_));
 sg13g2_a221oi_1 _5148_ (.B2(_1251_),
    .C1(_1321_),
    .B1(_0743_),
    .A1(net222),
    .Y(_1322_),
    .A2(_0578_));
 sg13g2_nand2_1 _5149_ (.Y(_1323_),
    .A(_0173_),
    .B(net52));
 sg13g2_a21oi_1 _5150_ (.A1(_1322_),
    .A2(_1323_),
    .Y(_1324_),
    .B1(net186));
 sg13g2_o21ai_1 _5151_ (.B1(_1324_),
    .Y(_1325_),
    .A1(_0737_),
    .A2(_1320_));
 sg13g2_nor2b_1 _5152_ (.A(_0681_),
    .B_N(_0813_),
    .Y(_1327_));
 sg13g2_nor2_1 _5153_ (.A(net146),
    .B(_2800_),
    .Y(_1328_));
 sg13g2_nand3_1 _5154_ (.B(net139),
    .C(_0847_),
    .A(_1158_),
    .Y(_1329_));
 sg13g2_nor2_1 _5155_ (.A(_2724_),
    .B(_0143_),
    .Y(_1330_));
 sg13g2_nor2_1 _5156_ (.A(net144),
    .B(_1330_),
    .Y(_1331_));
 sg13g2_a22oi_1 _5157_ (.Y(_1332_),
    .B1(_1329_),
    .B2(_1331_),
    .A2(_1328_),
    .A1(_2825_));
 sg13g2_o21ai_1 _5158_ (.B1(_1332_),
    .Y(_1333_),
    .A1(net63),
    .A2(_1327_));
 sg13g2_o21ai_1 _5159_ (.B1(_2967_),
    .Y(_1334_),
    .A1(_2644_),
    .A2(_2392_));
 sg13g2_nand2_1 _5160_ (.Y(_1335_),
    .A(_2495_),
    .B(_0954_));
 sg13g2_a21oi_1 _5161_ (.A1(_1334_),
    .A2(_1335_),
    .Y(_1336_),
    .B1(_0550_));
 sg13g2_nand2b_1 _5162_ (.Y(_1338_),
    .B(net215),
    .A_N(_1336_));
 sg13g2_a21oi_1 _5163_ (.A1(_1333_),
    .A2(net140),
    .Y(_1339_),
    .B1(_1338_));
 sg13g2_a21oi_1 _5164_ (.A1(_1325_),
    .A2(_1339_),
    .Y(_1340_),
    .B1(_2640_));
 sg13g2_nand2_1 _5165_ (.Y(_1341_),
    .A(_1314_),
    .B(_1340_));
 sg13g2_inv_1 _5166_ (.Y(_1342_),
    .A(_2461_));
 sg13g2_a22oi_1 _5167_ (.Y(_1343_),
    .B1(net105),
    .B2(_0338_),
    .A2(net120),
    .A1(_1342_));
 sg13g2_a21o_1 _5168_ (.A2(_2397_),
    .A1(_0939_),
    .B1(_0304_),
    .X(_1344_));
 sg13g2_a21oi_1 _5169_ (.A1(_1343_),
    .A2(_1344_),
    .Y(_1345_),
    .B1(net135));
 sg13g2_nand3_1 _5170_ (.B(_2378_),
    .C(_2145_),
    .A(_0621_),
    .Y(_1346_));
 sg13g2_nor2_1 _5171_ (.A(net172),
    .B(_1193_),
    .Y(_1347_));
 sg13g2_a21oi_1 _5172_ (.A1(_2583_),
    .A2(_1347_),
    .Y(_1349_),
    .B1(_0283_));
 sg13g2_a21o_1 _5173_ (.A2(_1349_),
    .A1(_1346_),
    .B1(net133),
    .X(_1350_));
 sg13g2_nor2b_1 _5174_ (.A(_1166_),
    .B_N(_2781_),
    .Y(_1351_));
 sg13g2_nor2_1 _5175_ (.A(_3051_),
    .B(_2493_),
    .Y(_1352_));
 sg13g2_nor3_1 _5176_ (.A(net145),
    .B(_1351_),
    .C(_1352_),
    .Y(_1353_));
 sg13g2_nor2_1 _5177_ (.A(net191),
    .B(_2938_),
    .Y(_1354_));
 sg13g2_a21oi_1 _5178_ (.A1(_0125_),
    .A2(_0667_),
    .Y(_1355_),
    .B1(net60));
 sg13g2_a21oi_1 _5179_ (.A1(_1354_),
    .A2(_0744_),
    .Y(_1356_),
    .B1(_1355_));
 sg13g2_a21oi_1 _5180_ (.A1(_1353_),
    .A2(_1356_),
    .Y(_1357_),
    .B1(_3044_));
 sg13g2_o21ai_1 _5181_ (.B1(_1357_),
    .Y(_1358_),
    .A1(_1345_),
    .A2(_1350_));
 sg13g2_nand2_2 _5182_ (.Y(_1360_),
    .A(_2703_),
    .B(net173));
 sg13g2_nand3_1 _5183_ (.B(_1360_),
    .C(net147),
    .A(_2503_),
    .Y(_1361_));
 sg13g2_nand2_1 _5184_ (.Y(_1362_),
    .A(_0528_),
    .B(_0914_));
 sg13g2_nor2_2 _5185_ (.A(_2398_),
    .B(_0153_),
    .Y(_1363_));
 sg13g2_a21oi_1 _5186_ (.A1(_1363_),
    .A2(_0667_),
    .Y(_1364_),
    .B1(net84));
 sg13g2_a22oi_1 _5187_ (.Y(_1365_),
    .B1(_1362_),
    .B2(_1364_),
    .A2(net54),
    .A1(_1361_));
 sg13g2_a21oi_1 _5188_ (.A1(_1354_),
    .A2(_2973_),
    .Y(_1366_),
    .B1(net141));
 sg13g2_nand2_1 _5189_ (.Y(_1367_),
    .A(_1365_),
    .B(_1366_));
 sg13g2_nor2_1 _5190_ (.A(_1267_),
    .B(_0880_),
    .Y(_1368_));
 sg13g2_a21oi_1 _5191_ (.A1(_1293_),
    .A2(_0752_),
    .Y(_1369_),
    .B1(_1368_));
 sg13g2_o21ai_1 _5192_ (.B1(net98),
    .Y(_1371_),
    .A1(_0153_),
    .A2(_2663_));
 sg13g2_nand3_1 _5193_ (.B(_1371_),
    .C(net133),
    .A(_1369_),
    .Y(_1372_));
 sg13g2_nand3_1 _5194_ (.B(net138),
    .C(_1372_),
    .A(_1367_),
    .Y(_1373_));
 sg13g2_nand3_1 _5195_ (.B(net190),
    .C(_1373_),
    .A(_1358_),
    .Y(_1374_));
 sg13g2_inv_1 _5196_ (.Y(_1375_),
    .A(_0752_));
 sg13g2_nor3_1 _5197_ (.A(net160),
    .B(_2538_),
    .C(_1375_),
    .Y(_1376_));
 sg13g2_a21oi_1 _5198_ (.A1(_1028_),
    .A2(_2913_),
    .Y(_1377_),
    .B1(net63));
 sg13g2_a21oi_1 _5199_ (.A1(_2540_),
    .A2(net126),
    .Y(_1378_),
    .B1(_2600_));
 sg13g2_nand2_1 _5200_ (.Y(_1379_),
    .A(_0880_),
    .B(net158));
 sg13g2_nand2_1 _5201_ (.Y(_1380_),
    .A(_1379_),
    .B(net155));
 sg13g2_a21oi_1 _5202_ (.A1(_1378_),
    .A2(net88),
    .Y(_1382_),
    .B1(_1380_));
 sg13g2_nor3_1 _5203_ (.A(_1376_),
    .B(_1377_),
    .C(_1382_),
    .Y(_1383_));
 sg13g2_nor2b_1 _5204_ (.A(net55),
    .B_N(_1383_),
    .Y(_1384_));
 sg13g2_nand3_1 _5205_ (.B(net76),
    .C(_1005_),
    .A(_0944_),
    .Y(_1385_));
 sg13g2_a21oi_1 _5206_ (.A1(_1035_),
    .A2(_2723_),
    .Y(_1386_),
    .B1(net152));
 sg13g2_nand2_1 _5207_ (.Y(_1387_),
    .A(_1385_),
    .B(_1386_));
 sg13g2_nor3_1 _5208_ (.A(net146),
    .B(_2502_),
    .C(_1203_),
    .Y(_1388_));
 sg13g2_a21oi_1 _5209_ (.A1(_1099_),
    .A2(_2885_),
    .Y(_1389_),
    .B1(_2595_));
 sg13g2_nor3_1 _5210_ (.A(net141),
    .B(_1388_),
    .C(_1389_),
    .Y(_1390_));
 sg13g2_a21o_1 _5211_ (.A2(_1390_),
    .A1(_1387_),
    .B1(net138),
    .X(_1391_));
 sg13g2_a22oi_1 _5212_ (.Y(_1393_),
    .B1(_0175_),
    .B2(_0745_),
    .A2(_0981_),
    .A1(_0407_));
 sg13g2_a21oi_1 _5213_ (.A1(_1393_),
    .A2(net75),
    .Y(_1394_),
    .B1(net93));
 sg13g2_a21oi_1 _5214_ (.A1(_1157_),
    .A2(_2654_),
    .Y(_1395_),
    .B1(net110));
 sg13g2_nor2_1 _5215_ (.A(net117),
    .B(_2585_),
    .Y(_1396_));
 sg13g2_nand3_1 _5216_ (.B(net89),
    .C(_1396_),
    .A(_1192_),
    .Y(_1397_));
 sg13g2_nand2_1 _5217_ (.Y(_1398_),
    .A(_1395_),
    .B(_1397_));
 sg13g2_nand2_1 _5218_ (.Y(_1399_),
    .A(_1394_),
    .B(_1398_));
 sg13g2_nand2_1 _5219_ (.Y(_1400_),
    .A(_0216_),
    .B(_1342_));
 sg13g2_inv_1 _5220_ (.Y(_1401_),
    .A(_1400_));
 sg13g2_o21ai_1 _5221_ (.B1(_1142_),
    .Y(_1402_),
    .A1(_0107_),
    .A2(_1401_));
 sg13g2_nor3_1 _5222_ (.A(net97),
    .B(net81),
    .C(_2250_),
    .Y(_1404_));
 sg13g2_nor2_1 _5223_ (.A(_1166_),
    .B(_2563_),
    .Y(_1405_));
 sg13g2_nor3_1 _5224_ (.A(net193),
    .B(_1404_),
    .C(_1405_),
    .Y(_1406_));
 sg13g2_a21oi_1 _5225_ (.A1(_1402_),
    .A2(_1406_),
    .Y(_1407_),
    .B1(net199));
 sg13g2_a21oi_1 _5226_ (.A1(_1399_),
    .A2(_1407_),
    .Y(_1408_),
    .B1(net188));
 sg13g2_o21ai_1 _5227_ (.B1(_1408_),
    .Y(_1409_),
    .A1(_1384_),
    .A2(_1391_));
 sg13g2_nand3_1 _5228_ (.B(_1409_),
    .C(net182),
    .A(_1374_),
    .Y(_1410_));
 sg13g2_nand2_1 _5229_ (.Y(_0028_),
    .A(_1341_),
    .B(_1410_));
 sg13g2_nand2_1 _5230_ (.Y(_1411_),
    .A(_0278_),
    .B(net57));
 sg13g2_nand2_1 _5231_ (.Y(_1412_),
    .A(_2905_),
    .B(net42));
 sg13g2_nand3_1 _5232_ (.B(net89),
    .C(_1412_),
    .A(_1411_),
    .Y(_1414_));
 sg13g2_a21oi_1 _5233_ (.A1(_0096_),
    .A2(_1158_),
    .Y(_1415_),
    .B1(net110));
 sg13g2_nand2_1 _5234_ (.Y(_1416_),
    .A(_1414_),
    .B(_1415_));
 sg13g2_nand3_1 _5235_ (.B(_2784_),
    .C(_2426_),
    .A(net82),
    .Y(_1417_));
 sg13g2_a21o_1 _5236_ (.A2(_1417_),
    .A1(_1131_),
    .B1(_2529_),
    .X(_1418_));
 sg13g2_nand3_1 _5237_ (.B(_2548_),
    .C(_1418_),
    .A(_1416_),
    .Y(_1419_));
 sg13g2_nor2_1 _5238_ (.A(net121),
    .B(_2686_),
    .Y(_1420_));
 sg13g2_nor3_1 _5239_ (.A(_2422_),
    .B(_0935_),
    .C(_2979_),
    .Y(_1421_));
 sg13g2_a21oi_1 _5240_ (.A1(_0184_),
    .A2(_1360_),
    .Y(_1422_),
    .B1(net80));
 sg13g2_nor3_1 _5241_ (.A(_1420_),
    .B(_1421_),
    .C(_1422_),
    .Y(_1423_));
 sg13g2_a21oi_1 _5242_ (.A1(_1423_),
    .A2(net125),
    .Y(_1425_),
    .B1(net187));
 sg13g2_nor2_1 _5243_ (.A(_2250_),
    .B(_0310_),
    .Y(_1426_));
 sg13g2_nor2_1 _5244_ (.A(_1817_),
    .B(_2755_),
    .Y(_1427_));
 sg13g2_inv_1 _5245_ (.Y(_1428_),
    .A(_1427_));
 sg13g2_a21oi_1 _5246_ (.A1(_1428_),
    .A2(_0235_),
    .Y(_1429_),
    .B1(net88));
 sg13g2_o21ai_1 _5247_ (.B1(_0549_),
    .Y(_1430_),
    .A1(_1426_),
    .A2(_1429_));
 sg13g2_nand2_1 _5248_ (.Y(_1431_),
    .A(_1430_),
    .B(_3010_));
 sg13g2_a21oi_1 _5249_ (.A1(_1419_),
    .A2(_1425_),
    .Y(_1432_),
    .B1(_1431_));
 sg13g2_o21ai_1 _5250_ (.B1(_0331_),
    .Y(_1433_),
    .A1(_0585_),
    .A2(_2762_));
 sg13g2_a22oi_1 _5251_ (.Y(_1434_),
    .B1(net62),
    .B2(_1433_),
    .A2(_0575_),
    .A1(_2922_));
 sg13g2_a21oi_1 _5252_ (.A1(_1675_),
    .A2(net70),
    .Y(_1436_),
    .B1(_1316_));
 sg13g2_nand2_1 _5253_ (.Y(_1437_),
    .A(_2932_),
    .B(net83));
 sg13g2_a22oi_1 _5254_ (.Y(_1438_),
    .B1(net77),
    .B2(_1437_),
    .A2(_1427_),
    .A1(net157));
 sg13g2_o21ai_1 _5255_ (.B1(_1438_),
    .Y(_1439_),
    .A1(net88),
    .A2(_1436_));
 sg13g2_nand2_1 _5256_ (.Y(_1440_),
    .A(_1439_),
    .B(net135));
 sg13g2_nand2_1 _5257_ (.Y(_1441_),
    .A(_1434_),
    .B(_1440_));
 sg13g2_nand2_1 _5258_ (.Y(_1442_),
    .A(_1441_),
    .B(_0308_));
 sg13g2_a21oi_1 _5259_ (.A1(_1432_),
    .A2(_1442_),
    .Y(_1443_),
    .B1(_0713_));
 sg13g2_o21ai_1 _5260_ (.B1(_0455_),
    .Y(_1444_),
    .A1(_0374_),
    .A2(_2907_));
 sg13g2_a21oi_1 _5261_ (.A1(net120),
    .A2(_0570_),
    .Y(_1445_),
    .B1(_1426_));
 sg13g2_a21o_1 _5262_ (.A2(_1445_),
    .A1(_1444_),
    .B1(_2405_),
    .X(_1447_));
 sg13g2_nor2_1 _5263_ (.A(net128),
    .B(_2856_),
    .Y(_1448_));
 sg13g2_inv_1 _5264_ (.Y(_1449_),
    .A(_2446_));
 sg13g2_nand2_1 _5265_ (.Y(_1450_),
    .A(_2812_),
    .B(net41));
 sg13g2_a21oi_1 _5266_ (.A1(_1449_),
    .A2(_1450_),
    .Y(_1451_),
    .B1(_1301_));
 sg13g2_a21oi_1 _5267_ (.A1(_0774_),
    .A2(net73),
    .Y(_1452_),
    .B1(net68));
 sg13g2_nor3_1 _5268_ (.A(_1448_),
    .B(_1451_),
    .C(_1452_),
    .Y(_1453_));
 sg13g2_nand2b_1 _5269_ (.Y(_1454_),
    .B(net125),
    .A_N(_1453_));
 sg13g2_a21oi_1 _5270_ (.A1(_3048_),
    .A2(_0516_),
    .Y(_1455_),
    .B1(_0325_));
 sg13g2_nand2_1 _5271_ (.Y(_1456_),
    .A(_1455_),
    .B(net171));
 sg13g2_nand3_1 _5272_ (.B(_1454_),
    .C(_1456_),
    .A(_1447_),
    .Y(_1458_));
 sg13g2_nand2_1 _5273_ (.Y(_1459_),
    .A(_1458_),
    .B(net166));
 sg13g2_inv_2 _5274_ (.Y(_1460_),
    .A(_2872_));
 sg13g2_nand3_1 _5275_ (.B(_0093_),
    .C(_1460_),
    .A(_0727_),
    .Y(_1461_));
 sg13g2_a22oi_1 _5276_ (.Y(_1462_),
    .B1(net40),
    .B2(_1461_),
    .A2(net136),
    .A1(_0759_));
 sg13g2_o21ai_1 _5277_ (.B1(_0917_),
    .Y(_1463_),
    .A1(_0911_),
    .A2(_0180_));
 sg13g2_a21oi_1 _5278_ (.A1(_1462_),
    .A2(_1463_),
    .Y(_1464_),
    .B1(net165));
 sg13g2_nand2_1 _5279_ (.Y(_1465_),
    .A(_2736_),
    .B(net169));
 sg13g2_nor2_1 _5280_ (.A(_1465_),
    .B(_2731_),
    .Y(_1466_));
 sg13g2_o21ai_1 _5281_ (.B1(net90),
    .Y(_1467_),
    .A1(_0338_),
    .A2(_1466_));
 sg13g2_nand2_1 _5282_ (.Y(_1469_),
    .A(_0629_),
    .B(_1158_));
 sg13g2_a21oi_1 _5283_ (.A1(_1469_),
    .A2(_2839_),
    .Y(_1470_),
    .B1(_1259_));
 sg13g2_nand2_1 _5284_ (.Y(_1471_),
    .A(_1467_),
    .B(_1470_));
 sg13g2_a21oi_1 _5285_ (.A1(_1471_),
    .A2(net140),
    .Y(_1472_),
    .B1(_2630_));
 sg13g2_nor2b_1 _5286_ (.A(_1464_),
    .B_N(_1472_),
    .Y(_1473_));
 sg13g2_nand2_1 _5287_ (.Y(_1474_),
    .A(_1459_),
    .B(_1473_));
 sg13g2_nand2_1 _5288_ (.Y(_1475_),
    .A(_1443_),
    .B(_1474_));
 sg13g2_a21oi_1 _5289_ (.A1(_1428_),
    .A2(_0914_),
    .Y(_1476_),
    .B1(net152));
 sg13g2_nand2_1 _5290_ (.Y(_1477_),
    .A(_1181_),
    .B(_1363_));
 sg13g2_nand2_1 _5291_ (.Y(_1478_),
    .A(_2806_),
    .B(_0914_));
 sg13g2_a22oi_1 _5292_ (.Y(_1480_),
    .B1(_2874_),
    .B2(_1478_),
    .A2(_1477_),
    .A1(_1476_));
 sg13g2_nor2_1 _5293_ (.A(_2469_),
    .B(_1480_),
    .Y(_1481_));
 sg13g2_nand3_1 _5294_ (.B(_3019_),
    .C(_1460_),
    .A(_0727_),
    .Y(_1482_));
 sg13g2_a22oi_1 _5295_ (.Y(_1483_),
    .B1(net76),
    .B2(_1482_),
    .A2(_0836_),
    .A1(_2476_));
 sg13g2_nor3_1 _5296_ (.A(_0034_),
    .B(net165),
    .C(_1483_),
    .Y(_1484_));
 sg13g2_nor2_1 _5297_ (.A(_1481_),
    .B(_1484_),
    .Y(_1485_));
 sg13g2_inv_1 _5298_ (.Y(_1486_),
    .A(_0165_));
 sg13g2_nand2_1 _5299_ (.Y(_1487_),
    .A(_1411_),
    .B(_1486_));
 sg13g2_nand2_1 _5300_ (.Y(_1488_),
    .A(_1487_),
    .B(net62));
 sg13g2_nand2b_1 _5301_ (.Y(_1489_),
    .B(_3038_),
    .A_N(_1231_));
 sg13g2_nand2_1 _5302_ (.Y(_1491_),
    .A(_1489_),
    .B(net47));
 sg13g2_nand3_1 _5303_ (.B(net53),
    .C(_2720_),
    .A(net44),
    .Y(_1492_));
 sg13g2_a21oi_1 _5304_ (.A1(_1075_),
    .A2(_0752_),
    .Y(_1493_),
    .B1(net184));
 sg13g2_nand4_1 _5305_ (.B(_1491_),
    .C(_1492_),
    .A(_1488_),
    .Y(_1494_),
    .D(_1493_));
 sg13g2_inv_1 _5306_ (.Y(_1495_),
    .A(_1181_));
 sg13g2_nor2_1 _5307_ (.A(net172),
    .B(_2980_),
    .Y(_1496_));
 sg13g2_nand2_1 _5308_ (.Y(_1497_),
    .A(net117),
    .B(net121));
 sg13g2_a21oi_1 _5309_ (.A1(_1496_),
    .A2(_1497_),
    .Y(_1498_),
    .B1(net144));
 sg13g2_o21ai_1 _5310_ (.B1(_1498_),
    .Y(_1499_),
    .A1(_0908_),
    .A2(_1495_));
 sg13g2_nand2_1 _5311_ (.Y(_1500_),
    .A(_2401_),
    .B(_2024_));
 sg13g2_a21oi_1 _5312_ (.A1(_0242_),
    .A2(_1500_),
    .Y(_1502_),
    .B1(net146));
 sg13g2_nand2_1 _5313_ (.Y(_1503_),
    .A(_3016_),
    .B(_2621_));
 sg13g2_o21ai_1 _5314_ (.B1(net192),
    .Y(_1504_),
    .A1(_0976_),
    .A2(_1503_));
 sg13g2_nor2_1 _5315_ (.A(_1502_),
    .B(_1504_),
    .Y(_1505_));
 sg13g2_a21oi_1 _5316_ (.A1(_1499_),
    .A2(_1505_),
    .Y(_1506_),
    .B1(net187));
 sg13g2_a21oi_1 _5317_ (.A1(_1494_),
    .A2(_1506_),
    .Y(_1507_),
    .B1(net183));
 sg13g2_nand2_1 _5318_ (.Y(_1508_),
    .A(_1485_),
    .B(_1507_));
 sg13g2_nand2_1 _5319_ (.Y(_1509_),
    .A(_1028_),
    .B(_2402_));
 sg13g2_nor2_1 _5320_ (.A(_0924_),
    .B(_1466_),
    .Y(_1510_));
 sg13g2_a21oi_1 _5321_ (.A1(_0278_),
    .A2(_0752_),
    .Y(_1511_),
    .B1(net174));
 sg13g2_o21ai_1 _5322_ (.B1(_1511_),
    .Y(_1513_),
    .A1(_1380_),
    .A2(_1510_));
 sg13g2_a21oi_1 _5323_ (.A1(net47),
    .A2(_1509_),
    .Y(_1514_),
    .B1(_1513_));
 sg13g2_nor2_1 _5324_ (.A(net186),
    .B(_1514_),
    .Y(_1515_));
 sg13g2_nand3_1 _5325_ (.B(net48),
    .C(_2915_),
    .A(_1486_),
    .Y(_1516_));
 sg13g2_nor2_1 _5326_ (.A(net158),
    .B(_2667_),
    .Y(_1517_));
 sg13g2_nand2_1 _5327_ (.Y(_1518_),
    .A(_2899_),
    .B(_1517_));
 sg13g2_nand3_1 _5328_ (.B(net135),
    .C(_1518_),
    .A(_1516_),
    .Y(_1519_));
 sg13g2_nand2_1 _5329_ (.Y(_1520_),
    .A(_0285_),
    .B(_2723_));
 sg13g2_nand3_1 _5330_ (.B(net122),
    .C(_1400_),
    .A(_0422_),
    .Y(_1521_));
 sg13g2_nand3_1 _5331_ (.B(net50),
    .C(_1521_),
    .A(_1520_),
    .Y(_1522_));
 sg13g2_nand3_1 _5332_ (.B(_1522_),
    .C(net55),
    .A(_1519_),
    .Y(_1524_));
 sg13g2_nand2_1 _5333_ (.Y(_1525_),
    .A(_1515_),
    .B(_1524_));
 sg13g2_a221oi_1 _5334_ (.B2(_0473_),
    .C1(net184),
    .B1(_1110_),
    .A1(_0231_),
    .Y(_1526_),
    .A2(_3016_));
 sg13g2_a21o_1 _5335_ (.A2(net73),
    .A1(_3033_),
    .B1(_1267_),
    .X(_1527_));
 sg13g2_a21oi_1 _5336_ (.A1(_1526_),
    .A2(_1527_),
    .Y(_1528_),
    .B1(net199));
 sg13g2_o21ai_1 _5337_ (.B1(_2859_),
    .Y(_1529_),
    .A1(_2625_),
    .A2(_0992_));
 sg13g2_nand3_1 _5338_ (.B(net139),
    .C(_2878_),
    .A(_2951_),
    .Y(_1530_));
 sg13g2_nand3_1 _5339_ (.B(_1530_),
    .C(net136),
    .A(_1529_),
    .Y(_1531_));
 sg13g2_nand2_1 _5340_ (.Y(_1532_),
    .A(_1509_),
    .B(net62));
 sg13g2_nand2_1 _5341_ (.Y(_1533_),
    .A(_0177_),
    .B(net73));
 sg13g2_a21oi_1 _5342_ (.A1(_1533_),
    .A2(net53),
    .Y(_1535_),
    .B1(net93));
 sg13g2_nand3_1 _5343_ (.B(_1532_),
    .C(_1535_),
    .A(_1531_),
    .Y(_1536_));
 sg13g2_a21oi_1 _5344_ (.A1(_1528_),
    .A2(_1536_),
    .Y(_1537_),
    .B1(net188));
 sg13g2_nand2_1 _5345_ (.Y(_1538_),
    .A(_1525_),
    .B(_1537_));
 sg13g2_nand3_1 _5346_ (.B(_1538_),
    .C(net182),
    .A(_1508_),
    .Y(_1539_));
 sg13g2_nand2_1 _5347_ (.Y(_0029_),
    .A(_1475_),
    .B(_1539_));
 sg13g2_o21ai_1 _5348_ (.B1(_0235_),
    .Y(_1540_),
    .A1(_3014_),
    .A2(_2963_));
 sg13g2_nand2_1 _5349_ (.Y(_1541_),
    .A(_2412_),
    .B(_2546_));
 sg13g2_a21oi_1 _5350_ (.A1(net115),
    .A2(_2384_),
    .Y(_1542_),
    .B1(_1541_));
 sg13g2_o21ai_1 _5351_ (.B1(_1542_),
    .Y(_1543_),
    .A1(_2705_),
    .A2(_0910_));
 sg13g2_a21oi_1 _5352_ (.A1(_0532_),
    .A2(_1540_),
    .Y(_1545_),
    .B1(_1543_));
 sg13g2_a22oi_1 _5353_ (.Y(_1546_),
    .B1(net120),
    .B2(_0620_),
    .A2(net56),
    .A1(net139));
 sg13g2_a21o_1 _5354_ (.A2(_0250_),
    .A1(_1546_),
    .B1(net136),
    .X(_1547_));
 sg13g2_a21oi_1 _5355_ (.A1(_2646_),
    .A2(_2503_),
    .Y(_1548_),
    .B1(_2527_));
 sg13g2_o21ai_1 _5356_ (.B1(_0734_),
    .Y(_1549_),
    .A1(net69),
    .A2(_1342_));
 sg13g2_nand2_1 _5357_ (.Y(_1550_),
    .A(_1549_),
    .B(_1275_));
 sg13g2_nand2_1 _5358_ (.Y(_1551_),
    .A(_2653_),
    .B(net99));
 sg13g2_nand3_1 _5359_ (.B(_1011_),
    .C(_1551_),
    .A(_1550_),
    .Y(_1552_));
 sg13g2_nor2_1 _5360_ (.A(_1548_),
    .B(_1552_),
    .Y(_1553_));
 sg13g2_a21oi_1 _5361_ (.A1(_1545_),
    .A2(_1547_),
    .Y(_1554_),
    .B1(_1553_));
 sg13g2_nand2_1 _5362_ (.Y(_1556_),
    .A(_1229_),
    .B(_2436_));
 sg13g2_nand2_1 _5363_ (.Y(_1557_),
    .A(_3014_),
    .B(_2384_));
 sg13g2_nand4_1 _5364_ (.B(_2998_),
    .C(net121),
    .A(_1557_),
    .Y(_1558_),
    .D(_2775_));
 sg13g2_nand3_1 _5365_ (.B(_1558_),
    .C(net191),
    .A(_1556_),
    .Y(_1559_));
 sg13g2_o21ai_1 _5366_ (.B1(_0917_),
    .Y(_1560_),
    .A1(net168),
    .A2(net56));
 sg13g2_nand3_1 _5367_ (.B(net184),
    .C(_1560_),
    .A(_1559_),
    .Y(_1561_));
 sg13g2_a21oi_1 _5368_ (.A1(_1174_),
    .A2(_0611_),
    .Y(_1562_),
    .B1(net159));
 sg13g2_a21oi_1 _5369_ (.A1(_1686_),
    .A2(_1465_),
    .Y(_1563_),
    .B1(net128));
 sg13g2_nor3_1 _5370_ (.A(_1259_),
    .B(_1562_),
    .C(_1563_),
    .Y(_1564_));
 sg13g2_nand2_1 _5371_ (.Y(_1565_),
    .A(_1564_),
    .B(_2711_));
 sg13g2_nand2_1 _5372_ (.Y(_1567_),
    .A(_1561_),
    .B(_1565_));
 sg13g2_nand2_1 _5373_ (.Y(_1568_),
    .A(_1567_),
    .B(_3042_));
 sg13g2_nand2_1 _5374_ (.Y(_1569_),
    .A(_1554_),
    .B(_1568_));
 sg13g2_nand2_1 _5375_ (.Y(_1570_),
    .A(_1569_),
    .B(_2517_));
 sg13g2_nor2_1 _5376_ (.A(_0414_),
    .B(_2934_),
    .Y(_1571_));
 sg13g2_nor2b_1 _5377_ (.A(_0544_),
    .B_N(_1251_),
    .Y(_1572_));
 sg13g2_nor3_1 _5378_ (.A(_0272_),
    .B(_1420_),
    .C(_1572_),
    .Y(_1573_));
 sg13g2_o21ai_1 _5379_ (.B1(_1573_),
    .Y(_1574_),
    .A1(net67),
    .A2(_1571_));
 sg13g2_nand2_1 _5380_ (.Y(_1575_),
    .A(_2615_),
    .B(_2488_));
 sg13g2_nand3_1 _5381_ (.B(_2999_),
    .C(_2775_),
    .A(_1575_),
    .Y(_1576_));
 sg13g2_nand2_1 _5382_ (.Y(_1578_),
    .A(_0458_),
    .B(_0096_));
 sg13g2_nand3_1 _5383_ (.B(_1578_),
    .C(_0141_),
    .A(_1576_),
    .Y(_1579_));
 sg13g2_o21ai_1 _5384_ (.B1(net94),
    .Y(_1580_),
    .A1(_0435_),
    .A2(_0772_));
 sg13g2_nand2_1 _5385_ (.Y(_1581_),
    .A(_1580_),
    .B(_0114_));
 sg13g2_nand3_1 _5386_ (.B(_1581_),
    .C(_0896_),
    .A(_1579_),
    .Y(_1582_));
 sg13g2_nand3_1 _5387_ (.B(net143),
    .C(_1582_),
    .A(_1574_),
    .Y(_1583_));
 sg13g2_a21oi_1 _5388_ (.A1(_2664_),
    .A2(_1496_),
    .Y(_1584_),
    .B1(_2551_));
 sg13g2_nand3_1 _5389_ (.B(_2985_),
    .C(net48),
    .A(_0419_),
    .Y(_1585_));
 sg13g2_nand2_1 _5390_ (.Y(_1586_),
    .A(_1584_),
    .B(_1585_));
 sg13g2_o21ai_1 _5391_ (.B1(net52),
    .Y(_1587_),
    .A1(_2435_),
    .A2(_0867_));
 sg13g2_a21oi_1 _5392_ (.A1(_0121_),
    .A2(net70),
    .Y(_1589_),
    .B1(net60));
 sg13g2_o21ai_1 _5393_ (.B1(_1589_),
    .Y(_1590_),
    .A1(_0353_),
    .A2(_0175_));
 sg13g2_nand3_1 _5394_ (.B(_1587_),
    .C(_1590_),
    .A(_1586_),
    .Y(_1591_));
 sg13g2_nand2_1 _5395_ (.Y(_1592_),
    .A(_1591_),
    .B(net87));
 sg13g2_a21oi_1 _5396_ (.A1(_2756_),
    .A2(_2486_),
    .Y(_1593_),
    .B1(_2634_));
 sg13g2_a221oi_1 _5397_ (.B2(_1417_),
    .C1(_0550_),
    .B1(_1593_),
    .A1(net105),
    .Y(_1594_),
    .A2(_1460_));
 sg13g2_nor2_1 _5398_ (.A(net183),
    .B(_1594_),
    .Y(_1595_));
 sg13g2_nand3_1 _5399_ (.B(_1592_),
    .C(_1595_),
    .A(_1583_),
    .Y(_1596_));
 sg13g2_nand3_1 _5400_ (.B(_1596_),
    .C(_0495_),
    .A(_1570_),
    .Y(_1597_));
 sg13g2_o21ai_1 _5401_ (.B1(_2634_),
    .Y(_1598_),
    .A1(_0911_),
    .A2(_0612_));
 sg13g2_nand2_1 _5402_ (.Y(_1600_),
    .A(_0557_),
    .B(net144));
 sg13g2_nor2_1 _5403_ (.A(net196),
    .B(net103),
    .Y(_1601_));
 sg13g2_a21oi_1 _5404_ (.A1(_1601_),
    .A2(_0093_),
    .Y(_1602_),
    .B1(net89));
 sg13g2_o21ai_1 _5405_ (.B1(_1602_),
    .Y(_1603_),
    .A1(_0123_),
    .A2(_1600_));
 sg13g2_nand3_1 _5406_ (.B(_0574_),
    .C(_1603_),
    .A(_1598_),
    .Y(_1604_));
 sg13g2_o21ai_1 _5407_ (.B1(net98),
    .Y(_1605_),
    .A1(_0094_),
    .A2(_0558_));
 sg13g2_a21oi_1 _5408_ (.A1(_1605_),
    .A2(_1194_),
    .Y(_1606_),
    .B1(_2417_));
 sg13g2_nor2_1 _5409_ (.A(_1375_),
    .B(_1437_),
    .Y(_1607_));
 sg13g2_a21oi_1 _5410_ (.A1(_1607_),
    .A2(net86),
    .Y(_1608_),
    .B1(net218));
 sg13g2_nand2b_1 _5411_ (.Y(_1609_),
    .B(_1608_),
    .A_N(_1606_));
 sg13g2_a21oi_1 _5412_ (.A1(_1604_),
    .A2(net87),
    .Y(_1611_),
    .B1(_1609_));
 sg13g2_nand2_1 _5413_ (.Y(_1612_),
    .A(_0557_),
    .B(net89));
 sg13g2_a21oi_1 _5414_ (.A1(_0719_),
    .A2(_0128_),
    .Y(_1613_),
    .B1(net134));
 sg13g2_o21ai_1 _5415_ (.B1(_1613_),
    .Y(_1614_),
    .A1(_2572_),
    .A2(_1612_));
 sg13g2_o21ai_1 _5416_ (.B1(_2777_),
    .Y(_1615_),
    .A1(_2973_),
    .A2(_0249_));
 sg13g2_nand2_1 _5417_ (.Y(_1616_),
    .A(_1615_),
    .B(net40));
 sg13g2_nand4_1 _5418_ (.B(net156),
    .C(_1503_),
    .A(_1614_),
    .Y(_1617_),
    .D(_1616_));
 sg13g2_inv_1 _5419_ (.Y(_1618_),
    .A(_0486_));
 sg13g2_nor2_1 _5420_ (.A(net103),
    .B(_2602_),
    .Y(_1619_));
 sg13g2_nor3_1 _5421_ (.A(net146),
    .B(_1618_),
    .C(_1619_),
    .Y(_1620_));
 sg13g2_a21oi_1 _5422_ (.A1(_0259_),
    .A2(net201),
    .Y(_1622_),
    .B1(net112));
 sg13g2_nor3_1 _5423_ (.A(net184),
    .B(_1620_),
    .C(_1622_),
    .Y(_1623_));
 sg13g2_nand3_1 _5424_ (.B(_1149_),
    .C(net92),
    .A(_2664_),
    .Y(_1624_));
 sg13g2_nand3_1 _5425_ (.B(net139),
    .C(_2811_),
    .A(_1360_),
    .Y(_1625_));
 sg13g2_nand3_1 _5426_ (.B(_1625_),
    .C(net50),
    .A(_1624_),
    .Y(_1626_));
 sg13g2_a21oi_1 _5427_ (.A1(_1623_),
    .A2(_1626_),
    .Y(_1627_),
    .B1(net186));
 sg13g2_nand2_1 _5428_ (.Y(_1628_),
    .A(_1617_),
    .B(_1627_));
 sg13g2_a21oi_1 _5429_ (.A1(_1611_),
    .A2(_1628_),
    .Y(_1629_),
    .B1(net212));
 sg13g2_a21oi_1 _5430_ (.A1(net81),
    .A2(net107),
    .Y(_1630_),
    .B1(net42));
 sg13g2_o21ai_1 _5431_ (.B1(net92),
    .Y(_1631_),
    .A1(_1630_),
    .A2(_2504_));
 sg13g2_o21ai_1 _5432_ (.B1(_0517_),
    .Y(_1633_),
    .A1(net42),
    .A2(_0248_));
 sg13g2_nand2_1 _5433_ (.Y(_1634_),
    .A(_1633_),
    .B(net89));
 sg13g2_a21o_1 _5434_ (.A2(_1634_),
    .A1(_1631_),
    .B1(net136),
    .X(_1635_));
 sg13g2_inv_1 _5435_ (.Y(_1636_),
    .A(_2300_));
 sg13g2_a21oi_1 _5436_ (.A1(_1636_),
    .A2(net39),
    .Y(_1637_),
    .B1(net146));
 sg13g2_o21ai_1 _5437_ (.B1(_0557_),
    .Y(_1638_),
    .A1(net201),
    .A2(net64));
 sg13g2_a22oi_1 _5438_ (.Y(_1639_),
    .B1(net47),
    .B2(_1638_),
    .A2(_1637_),
    .A1(_1449_));
 sg13g2_a21oi_1 _5439_ (.A1(_1635_),
    .A2(_1639_),
    .Y(_1640_),
    .B1(_2418_));
 sg13g2_a21oi_1 _5440_ (.A1(_0300_),
    .A2(_2854_),
    .Y(_1641_),
    .B1(net97));
 sg13g2_o21ai_1 _5441_ (.B1(_1641_),
    .Y(_1642_),
    .A1(_2399_),
    .A2(_2663_));
 sg13g2_nand2_1 _5442_ (.Y(_1644_),
    .A(_0999_),
    .B(_1360_));
 sg13g2_nand2_1 _5443_ (.Y(_1645_),
    .A(_1644_),
    .B(_1142_));
 sg13g2_a21oi_1 _5444_ (.A1(_1642_),
    .A2(_1645_),
    .Y(_1646_),
    .B1(net161));
 sg13g2_nor2_1 _5445_ (.A(net215),
    .B(_1646_),
    .Y(_1647_));
 sg13g2_nor2b_1 _5446_ (.A(_1640_),
    .B_N(_1647_),
    .Y(_1648_));
 sg13g2_nor2_1 _5447_ (.A(net43),
    .B(_0528_),
    .Y(_1649_));
 sg13g2_o21ai_1 _5448_ (.B1(net214),
    .Y(_1650_),
    .A1(_0248_),
    .A2(_2686_));
 sg13g2_a21oi_1 _5449_ (.A1(net90),
    .A2(_0881_),
    .Y(_1651_),
    .B1(_1650_));
 sg13g2_nand2_1 _5450_ (.Y(_1652_),
    .A(_2607_),
    .B(net45));
 sg13g2_nand3_1 _5451_ (.B(_1264_),
    .C(net98),
    .A(_1652_),
    .Y(_1653_));
 sg13g2_nand2_1 _5452_ (.Y(_1655_),
    .A(_1651_),
    .B(_1653_));
 sg13g2_nor3_1 _5453_ (.A(_1649_),
    .B(_1607_),
    .C(_1655_),
    .Y(_1656_));
 sg13g2_nor2b_1 _5454_ (.A(_2911_),
    .B_N(_1517_),
    .Y(_1657_));
 sg13g2_nor2_1 _5455_ (.A(net84),
    .B(_1657_),
    .Y(_1658_));
 sg13g2_o21ai_1 _5456_ (.B1(_1658_),
    .Y(_1659_),
    .A1(net105),
    .A2(_2916_));
 sg13g2_nand3_1 _5457_ (.B(net55),
    .C(_1659_),
    .A(_1522_),
    .Y(_1660_));
 sg13g2_nand3b_1 _5458_ (.B(_1660_),
    .C(net166),
    .Y(_1661_),
    .A_N(_1656_));
 sg13g2_nand2_1 _5459_ (.Y(_1662_),
    .A(_1648_),
    .B(_1661_));
 sg13g2_nand2_1 _5460_ (.Y(_1663_),
    .A(_1629_),
    .B(_1662_));
 sg13g2_nand2_1 _5461_ (.Y(_0017_),
    .A(_1597_),
    .B(_1663_));
 sg13g2_o21ai_1 _5462_ (.B1(_2769_),
    .Y(_1665_),
    .A1(_2968_),
    .A2(_2620_));
 sg13g2_nand3_1 _5463_ (.B(_2860_),
    .C(_1133_),
    .A(_1665_),
    .Y(_1666_));
 sg13g2_nand2_1 _5464_ (.Y(_1667_),
    .A(_2670_),
    .B(net126));
 sg13g2_nand3_1 _5465_ (.B(_2463_),
    .C(_1667_),
    .A(_1449_),
    .Y(_1668_));
 sg13g2_a21oi_1 _5466_ (.A1(_1666_),
    .A2(_1668_),
    .Y(_1669_),
    .B1(net145));
 sg13g2_nand3_1 _5467_ (.B(net200),
    .C(_1066_),
    .A(_0515_),
    .Y(_1670_));
 sg13g2_nor2_1 _5468_ (.A(_2550_),
    .B(_1670_),
    .Y(_1671_));
 sg13g2_nor2_1 _5469_ (.A(net200),
    .B(_1267_),
    .Y(_1672_));
 sg13g2_nand3_1 _5470_ (.B(_0373_),
    .C(_1672_),
    .A(_1360_),
    .Y(_1673_));
 sg13g2_nand2_1 _5471_ (.Y(_1674_),
    .A(_0866_),
    .B(_2458_));
 sg13g2_nand3_1 _5472_ (.B(_1970_),
    .C(_1674_),
    .A(_1673_),
    .Y(_1676_));
 sg13g2_nor2_1 _5473_ (.A(_1671_),
    .B(_1676_),
    .Y(_1677_));
 sg13g2_nor2_1 _5474_ (.A(_2412_),
    .B(_1677_),
    .Y(_1678_));
 sg13g2_nand2_1 _5475_ (.Y(_1679_),
    .A(_3051_),
    .B(_2474_));
 sg13g2_nand2_1 _5476_ (.Y(_1680_),
    .A(_0669_),
    .B(_1679_));
 sg13g2_nand4_1 _5477_ (.B(_0211_),
    .C(net163),
    .A(_1396_),
    .Y(_1681_),
    .D(_0662_));
 sg13g2_nand2_1 _5478_ (.Y(_1682_),
    .A(_1680_),
    .B(_1681_));
 sg13g2_nand2_1 _5479_ (.Y(_1683_),
    .A(_1682_),
    .B(_2406_));
 sg13g2_nand3b_1 _5480_ (.B(_1678_),
    .C(_1683_),
    .Y(_1684_),
    .A_N(_1669_));
 sg13g2_a21oi_1 _5481_ (.A1(_0640_),
    .A2(_2762_),
    .Y(_1685_),
    .B1(net137));
 sg13g2_nand2_1 _5482_ (.Y(_1687_),
    .A(_0577_),
    .B(_2714_));
 sg13g2_a21oi_1 _5483_ (.A1(_0478_),
    .A2(_1687_),
    .Y(_1688_),
    .B1(_2971_));
 sg13g2_o21ai_1 _5484_ (.B1(net134),
    .Y(_1689_),
    .A1(_1685_),
    .A2(_1688_));
 sg13g2_a21oi_1 _5485_ (.A1(_2424_),
    .A2(_2523_),
    .Y(_1690_),
    .B1(_1457_));
 sg13g2_a221oi_1 _5486_ (.B2(_2785_),
    .C1(net192),
    .B1(_1690_),
    .A1(_2708_),
    .Y(_1691_),
    .A2(_1205_));
 sg13g2_nand2_1 _5487_ (.Y(_1692_),
    .A(_1689_),
    .B(_1691_));
 sg13g2_a22oi_1 _5488_ (.Y(_1693_),
    .B1(net200),
    .B2(_2577_),
    .A2(_2648_),
    .A1(_2521_));
 sg13g2_nor2_1 _5489_ (.A(_2525_),
    .B(_1693_),
    .Y(_1694_));
 sg13g2_nor2_1 _5490_ (.A(_0792_),
    .B(_2921_),
    .Y(_1695_));
 sg13g2_nand3_1 _5491_ (.B(_0752_),
    .C(_2429_),
    .A(_2584_),
    .Y(_1696_));
 sg13g2_nand3b_1 _5492_ (.B(_1696_),
    .C(_2546_),
    .Y(_1698_),
    .A_N(_1695_));
 sg13g2_nor2_1 _5493_ (.A(_1694_),
    .B(_1698_),
    .Y(_1699_));
 sg13g2_nand2_1 _5494_ (.Y(_1700_),
    .A(_1486_),
    .B(_1149_));
 sg13g2_nand2_1 _5495_ (.Y(_1701_),
    .A(_1700_),
    .B(net85));
 sg13g2_a21oi_1 _5496_ (.A1(_1699_),
    .A2(_1701_),
    .Y(_1702_),
    .B1(net187));
 sg13g2_nand2_1 _5497_ (.Y(_1703_),
    .A(_1692_),
    .B(_1702_));
 sg13g2_nand2_1 _5498_ (.Y(_1704_),
    .A(_1684_),
    .B(_1703_));
 sg13g2_nand2_1 _5499_ (.Y(_1705_),
    .A(_1704_),
    .B(_0556_));
 sg13g2_nand2b_1 _5500_ (.Y(_1706_),
    .B(_0125_),
    .A_N(_2741_));
 sg13g2_nand2_1 _5501_ (.Y(_1707_),
    .A(_2225_),
    .B(net200));
 sg13g2_o21ai_1 _5502_ (.B1(net217),
    .Y(_1709_),
    .A1(_1707_),
    .A2(_1166_));
 sg13g2_a21oi_1 _5503_ (.A1(_1706_),
    .A2(_1796_),
    .Y(_1710_),
    .B1(_1709_));
 sg13g2_a21o_1 _5504_ (.A2(_0109_),
    .A1(_0430_),
    .B1(net179),
    .X(_1711_));
 sg13g2_inv_1 _5505_ (.Y(_1712_),
    .A(_0940_));
 sg13g2_nand3_1 _5506_ (.B(_2819_),
    .C(_0847_),
    .A(_1712_),
    .Y(_1713_));
 sg13g2_nand3_1 _5507_ (.B(_1711_),
    .C(_1713_),
    .A(_1710_),
    .Y(_1714_));
 sg13g2_nand2_1 _5508_ (.Y(_1715_),
    .A(_1714_),
    .B(net151));
 sg13g2_nor3_1 _5509_ (.A(net119),
    .B(_2600_),
    .C(_0173_),
    .Y(_1716_));
 sg13g2_inv_1 _5510_ (.Y(_1717_),
    .A(_1363_));
 sg13g2_a21oi_1 _5511_ (.A1(_1577_),
    .A2(_1675_),
    .Y(_1718_),
    .B1(_1717_));
 sg13g2_nor3_1 _5512_ (.A(net134),
    .B(_1716_),
    .C(_1718_),
    .Y(_1720_));
 sg13g2_a21o_1 _5513_ (.A2(_2723_),
    .A1(_2477_),
    .B1(net119),
    .X(_1721_));
 sg13g2_a22oi_1 _5514_ (.Y(_1722_),
    .B1(_2830_),
    .B2(_0429_),
    .A2(_2733_),
    .A1(_0326_));
 sg13g2_a21oi_1 _5515_ (.A1(_1721_),
    .A2(_1722_),
    .Y(_1723_),
    .B1(net50));
 sg13g2_nor3_1 _5516_ (.A(net150),
    .B(_1720_),
    .C(_1723_),
    .Y(_1724_));
 sg13g2_nor2_1 _5517_ (.A(_1715_),
    .B(_1724_),
    .Y(_1725_));
 sg13g2_nor2_1 _5518_ (.A(_1375_),
    .B(_0680_),
    .Y(_1726_));
 sg13g2_a21oi_1 _5519_ (.A1(_2792_),
    .A2(_3019_),
    .Y(_1727_),
    .B1(net111));
 sg13g2_nor4_1 _5520_ (.A(net174),
    .B(_1368_),
    .C(_1726_),
    .D(_1727_),
    .Y(_1728_));
 sg13g2_a21oi_1 _5521_ (.A1(_2994_),
    .A2(net73),
    .Y(_1729_),
    .B1(net68));
 sg13g2_nor3_1 _5522_ (.A(net96),
    .B(net80),
    .C(_0940_),
    .Y(_1731_));
 sg13g2_nor3_1 _5523_ (.A(_2547_),
    .B(_1729_),
    .C(_1731_),
    .Y(_1732_));
 sg13g2_o21ai_1 _5524_ (.B1(_0613_),
    .Y(_1733_),
    .A1(_2868_),
    .A2(_0534_));
 sg13g2_o21ai_1 _5525_ (.B1(_1733_),
    .Y(_1734_),
    .A1(_0668_),
    .A2(_1717_));
 sg13g2_nand2_1 _5526_ (.Y(_1735_),
    .A(_1732_),
    .B(_1734_));
 sg13g2_nand3b_1 _5527_ (.B(_1735_),
    .C(_2848_),
    .Y(_1736_),
    .A_N(_1728_));
 sg13g2_nor2b_1 _5528_ (.A(_1725_),
    .B_N(_1736_),
    .Y(_1737_));
 sg13g2_nand2_1 _5529_ (.Y(_1738_),
    .A(_1705_),
    .B(_1737_));
 sg13g2_nand2_1 _5530_ (.Y(_1739_),
    .A(_1738_),
    .B(net182));
 sg13g2_nand2_1 _5531_ (.Y(_1740_),
    .A(_0108_),
    .B(net82));
 sg13g2_a21o_1 _5532_ (.A2(_2937_),
    .A1(_1740_),
    .B1(_1267_),
    .X(_1742_));
 sg13g2_o21ai_1 _5533_ (.B1(net40),
    .Y(_1743_),
    .A1(_0123_),
    .A2(_1495_));
 sg13g2_o21ai_1 _5534_ (.B1(net47),
    .Y(_1744_),
    .A1(net117),
    .A2(_0137_));
 sg13g2_nand3_1 _5535_ (.B(_1743_),
    .C(_1744_),
    .A(_1742_),
    .Y(_1745_));
 sg13g2_a21oi_1 _5536_ (.A1(_1745_),
    .A2(net86),
    .Y(_1746_),
    .B1(net188));
 sg13g2_nand2_1 _5537_ (.Y(_1747_),
    .A(_1740_),
    .B(_1497_));
 sg13g2_nand3_1 _5538_ (.B(net83),
    .C(_2733_),
    .A(_1290_),
    .Y(_1748_));
 sg13g2_nand2_1 _5539_ (.Y(_1749_),
    .A(_0724_),
    .B(net77));
 sg13g2_nand3_1 _5540_ (.B(net122),
    .C(net178),
    .A(net96),
    .Y(_1750_));
 sg13g2_nand3_1 _5541_ (.B(_1749_),
    .C(_1750_),
    .A(_1748_),
    .Y(_1751_));
 sg13g2_a22oi_1 _5542_ (.Y(_1753_),
    .B1(net49),
    .B2(_1751_),
    .A2(_1747_),
    .A1(net47));
 sg13g2_nand2b_1 _5543_ (.Y(_1754_),
    .B(_0308_),
    .A_N(_1753_));
 sg13g2_nor2_1 _5544_ (.A(net39),
    .B(_2638_),
    .Y(_1755_));
 sg13g2_nor3_1 _5545_ (.A(_2551_),
    .B(_0301_),
    .C(_1755_),
    .Y(_1756_));
 sg13g2_a21oi_1 _5546_ (.A1(_0795_),
    .A2(_1106_),
    .Y(_1757_),
    .B1(net100));
 sg13g2_nand4_1 _5547_ (.B(_2397_),
    .C(_1796_),
    .A(_0373_),
    .Y(_1758_),
    .D(_2488_));
 sg13g2_nand2_1 _5548_ (.Y(_1759_),
    .A(_2638_),
    .B(_0578_));
 sg13g2_nand3_1 _5549_ (.B(net184),
    .C(_1759_),
    .A(_1758_),
    .Y(_1760_));
 sg13g2_nor3_1 _5550_ (.A(_1756_),
    .B(_1757_),
    .C(_1760_),
    .Y(_1761_));
 sg13g2_nor3_1 _5551_ (.A(_1301_),
    .B(_0094_),
    .C(net56),
    .Y(_1762_));
 sg13g2_nor3_1 _5552_ (.A(net184),
    .B(_1448_),
    .C(_1762_),
    .Y(_1764_));
 sg13g2_inv_1 _5553_ (.Y(_1765_),
    .A(_1158_));
 sg13g2_o21ai_1 _5554_ (.B1(net62),
    .Y(_1766_),
    .A1(net168),
    .A2(_1765_));
 sg13g2_a21oi_1 _5555_ (.A1(_1764_),
    .A2(_1766_),
    .Y(_1767_),
    .B1(net186));
 sg13g2_nand2b_1 _5556_ (.Y(_1768_),
    .B(_1767_),
    .A_N(_1761_));
 sg13g2_nand3_1 _5557_ (.B(_1754_),
    .C(_1768_),
    .A(_1746_),
    .Y(_1769_));
 sg13g2_a221oi_1 _5558_ (.B2(_0629_),
    .C1(_0550_),
    .B1(_0325_),
    .A1(_0727_),
    .Y(_1770_),
    .A2(net105));
 sg13g2_nor2_1 _5559_ (.A(net183),
    .B(_1770_),
    .Y(_1771_));
 sg13g2_nand2_1 _5560_ (.Y(_1772_),
    .A(_0992_),
    .B(net77));
 sg13g2_nand2_1 _5561_ (.Y(_1773_),
    .A(_0137_),
    .B(net120));
 sg13g2_nand3_1 _5562_ (.B(net119),
    .C(net147),
    .A(_2599_),
    .Y(_1775_));
 sg13g2_nand3_1 _5563_ (.B(_1773_),
    .C(_1775_),
    .A(_1772_),
    .Y(_1776_));
 sg13g2_a22oi_1 _5564_ (.Y(_1777_),
    .B1(net49),
    .B2(_1776_),
    .A2(_1251_),
    .A1(_0526_));
 sg13g2_nand2_1 _5565_ (.Y(_1778_),
    .A(_1777_),
    .B(net55));
 sg13g2_nand2_1 _5566_ (.Y(_1779_),
    .A(_1679_),
    .B(_0671_));
 sg13g2_nand3_1 _5567_ (.B(_0486_),
    .C(net92),
    .A(_0211_),
    .Y(_1780_));
 sg13g2_nand3_1 _5568_ (.B(net136),
    .C(_1780_),
    .A(_1779_),
    .Y(_1781_));
 sg13g2_o21ai_1 _5569_ (.B1(_0175_),
    .Y(_1782_),
    .A1(net106),
    .A2(_0426_));
 sg13g2_a21oi_1 _5570_ (.A1(_1782_),
    .A2(net53),
    .Y(_1783_),
    .B1(net93));
 sg13g2_a21oi_1 _5571_ (.A1(_1781_),
    .A2(_1783_),
    .Y(_1784_),
    .B1(net186));
 sg13g2_nand2_1 _5572_ (.Y(_1786_),
    .A(_1778_),
    .B(_1784_));
 sg13g2_a21oi_1 _5573_ (.A1(_1665_),
    .A2(_0510_),
    .Y(_1787_),
    .B1(_1267_));
 sg13g2_a21oi_1 _5574_ (.A1(_2835_),
    .A2(_0355_),
    .Y(_1788_),
    .B1(net100));
 sg13g2_inv_1 _5575_ (.Y(_1789_),
    .A(_2830_));
 sg13g2_nor2_1 _5576_ (.A(net116),
    .B(_1789_),
    .Y(_1790_));
 sg13g2_inv_1 _5577_ (.Y(_1791_),
    .A(_1095_));
 sg13g2_a22oi_1 _5578_ (.Y(_1792_),
    .B1(_2735_),
    .B2(_1791_),
    .A2(_1790_),
    .A1(_2905_));
 sg13g2_nand2b_1 _5579_ (.Y(_1793_),
    .B(_1792_),
    .A_N(_1788_));
 sg13g2_o21ai_1 _5580_ (.B1(net87),
    .Y(_1794_),
    .A1(_1787_),
    .A2(_1793_));
 sg13g2_nand3_1 _5581_ (.B(_1786_),
    .C(_1794_),
    .A(_1771_),
    .Y(_1795_));
 sg13g2_nand3_1 _5582_ (.B(_1795_),
    .C(net212),
    .A(_1769_),
    .Y(_1797_));
 sg13g2_nand2_1 _5583_ (.Y(_0018_),
    .A(_1739_),
    .B(_1797_));
 sg13g2_nor2_1 _5584_ (.A(_0923_),
    .B(_0882_),
    .Y(_1798_));
 sg13g2_a21oi_1 _5585_ (.A1(_1798_),
    .A2(_2575_),
    .Y(_1799_),
    .B1(_2711_));
 sg13g2_o21ai_1 _5586_ (.B1(_1799_),
    .Y(_1800_),
    .A1(_0903_),
    .A2(_1267_));
 sg13g2_o21ai_1 _5587_ (.B1(net99),
    .Y(_1801_),
    .A1(net226),
    .A2(_0133_));
 sg13g2_nand2_1 _5588_ (.Y(_1802_),
    .A(_0903_),
    .B(net139));
 sg13g2_nand2_1 _5589_ (.Y(_1803_),
    .A(_0880_),
    .B(_2447_));
 sg13g2_nand3_1 _5590_ (.B(_1802_),
    .C(_1803_),
    .A(_1801_),
    .Y(_1804_));
 sg13g2_nand2_1 _5591_ (.Y(_1805_),
    .A(_1804_),
    .B(_2946_));
 sg13g2_nand3_1 _5592_ (.B(net143),
    .C(_1805_),
    .A(_1800_),
    .Y(_1807_));
 sg13g2_nor2_1 _5593_ (.A(_2531_),
    .B(_0940_),
    .Y(_1808_));
 sg13g2_nor4_1 _5594_ (.A(_2184_),
    .B(_2673_),
    .C(_2980_),
    .D(_3024_),
    .Y(_1809_));
 sg13g2_nor4_1 _5595_ (.A(_2412_),
    .B(_0033_),
    .C(_1808_),
    .D(_1809_),
    .Y(_1810_));
 sg13g2_a21oi_1 _5596_ (.A1(net170),
    .A2(_2388_),
    .Y(_1811_),
    .B1(_1206_));
 sg13g2_nor2_1 _5597_ (.A(_3002_),
    .B(_1811_),
    .Y(_1812_));
 sg13g2_nor2_1 _5598_ (.A(_2529_),
    .B(_1812_),
    .Y(_1813_));
 sg13g2_a21oi_1 _5599_ (.A1(_0442_),
    .A2(_2845_),
    .Y(_1814_),
    .B1(_1813_));
 sg13g2_a21oi_1 _5600_ (.A1(_1810_),
    .A2(_1814_),
    .Y(_1815_),
    .B1(net188));
 sg13g2_nand2_1 _5601_ (.Y(_1816_),
    .A(_1807_),
    .B(_1815_));
 sg13g2_a21oi_1 _5602_ (.A1(_0231_),
    .A2(net213),
    .Y(_1818_),
    .B1(_2882_));
 sg13g2_a22oi_1 _5603_ (.Y(_1819_),
    .B1(net84),
    .B2(_1818_),
    .A2(_0118_),
    .A1(_1712_));
 sg13g2_nand3_1 _5604_ (.B(_2370_),
    .C(_2077_),
    .A(_1257_),
    .Y(_1820_));
 sg13g2_nand2_1 _5605_ (.Y(_1821_),
    .A(_1820_),
    .B(_0931_));
 sg13g2_a21oi_1 _5606_ (.A1(_1819_),
    .A2(_1821_),
    .Y(_1822_),
    .B1(_2629_));
 sg13g2_o21ai_1 _5607_ (.B1(_1379_),
    .Y(_1823_),
    .A1(_1090_),
    .A2(_2403_));
 sg13g2_inv_1 _5608_ (.Y(_1824_),
    .A(_1496_));
 sg13g2_nand2_1 _5609_ (.Y(_1825_),
    .A(_0477_),
    .B(net119));
 sg13g2_o21ai_1 _5610_ (.B1(_1825_),
    .Y(_1826_),
    .A1(_0940_),
    .A2(_1824_));
 sg13g2_a22oi_1 _5611_ (.Y(_1827_),
    .B1(net171),
    .B2(_1826_),
    .A2(_1823_),
    .A1(net167));
 sg13g2_nand2b_1 _5612_ (.Y(_1829_),
    .B(_1827_),
    .A_N(_1822_));
 sg13g2_nand2_1 _5613_ (.Y(_1830_),
    .A(_1829_),
    .B(net151));
 sg13g2_o21ai_1 _5614_ (.B1(_0956_),
    .Y(_1831_),
    .A1(_0153_),
    .A2(_1825_));
 sg13g2_nand2_1 _5615_ (.Y(_1832_),
    .A(_1831_),
    .B(net49));
 sg13g2_a21oi_1 _5616_ (.A1(_3032_),
    .A2(net213),
    .Y(_1833_),
    .B1(_2808_));
 sg13g2_nor3_1 _5617_ (.A(net141),
    .B(_1808_),
    .C(_1833_),
    .Y(_1834_));
 sg13g2_nand2_1 _5618_ (.Y(_1835_),
    .A(_1832_),
    .B(_1834_));
 sg13g2_a21oi_1 _5619_ (.A1(_1460_),
    .A2(_1363_),
    .Y(_1836_),
    .B1(_1818_));
 sg13g2_nand3_1 _5620_ (.B(net156),
    .C(_2635_),
    .A(_1836_),
    .Y(_1837_));
 sg13g2_nand3_1 _5621_ (.B(_2848_),
    .C(_1837_),
    .A(_1835_),
    .Y(_1838_));
 sg13g2_nand3_1 _5622_ (.B(_1830_),
    .C(_1838_),
    .A(_1816_),
    .Y(_1840_));
 sg13g2_nand2_1 _5623_ (.Y(_1841_),
    .A(_1840_),
    .B(net182));
 sg13g2_nand2_1 _5624_ (.Y(_1842_),
    .A(_0527_),
    .B(_2893_));
 sg13g2_a21oi_1 _5625_ (.A1(_1842_),
    .A2(_2845_),
    .Y(_1843_),
    .B1(_2840_));
 sg13g2_nor2_1 _5626_ (.A(_2701_),
    .B(_0868_),
    .Y(_1844_));
 sg13g2_o21ai_1 _5627_ (.B1(_1844_),
    .Y(_1845_),
    .A1(_0191_),
    .A2(_1811_));
 sg13g2_o21ai_1 _5628_ (.B1(net52),
    .Y(_1846_),
    .A1(net226),
    .A2(_2327_));
 sg13g2_nand3_1 _5629_ (.B(_0532_),
    .C(_2878_),
    .A(_0422_),
    .Y(_1847_));
 sg13g2_nand4_1 _5630_ (.B(_1845_),
    .C(_1846_),
    .A(_1843_),
    .Y(_1848_),
    .D(_1847_));
 sg13g2_a21oi_1 _5631_ (.A1(_1695_),
    .A2(_2548_),
    .Y(_1849_),
    .B1(_2413_));
 sg13g2_nand2_1 _5632_ (.Y(_1851_),
    .A(_1848_),
    .B(_1849_));
 sg13g2_nand3_1 _5633_ (.B(net90),
    .C(_2536_),
    .A(_0994_),
    .Y(_1852_));
 sg13g2_nand2_1 _5634_ (.Y(_1853_),
    .A(_0868_),
    .B(_2839_));
 sg13g2_a21o_1 _5635_ (.A2(_1853_),
    .A1(_1852_),
    .B1(net133),
    .X(_1854_));
 sg13g2_o21ai_1 _5636_ (.B1(_0283_),
    .Y(_1855_),
    .A1(_2734_),
    .A2(_0429_));
 sg13g2_nand4_1 _5637_ (.B(_2940_),
    .C(_0896_),
    .A(_1855_),
    .Y(_1856_),
    .D(_0827_));
 sg13g2_nand3_1 _5638_ (.B(_1856_),
    .C(_2749_),
    .A(_1854_),
    .Y(_1857_));
 sg13g2_nand3_1 _5639_ (.B(net190),
    .C(_1857_),
    .A(_1851_),
    .Y(_1858_));
 sg13g2_a21oi_1 _5640_ (.A1(_1257_),
    .A2(_0233_),
    .Y(_1859_),
    .B1(_2808_));
 sg13g2_o21ai_1 _5641_ (.B1(net116),
    .Y(_1860_),
    .A1(_0149_),
    .A2(_0891_));
 sg13g2_nand2_1 _5642_ (.Y(_1862_),
    .A(_1460_),
    .B(_0381_));
 sg13g2_nand2_1 _5643_ (.Y(_1863_),
    .A(_1860_),
    .B(_1862_));
 sg13g2_o21ai_1 _5644_ (.B1(net133),
    .Y(_1864_),
    .A1(_1859_),
    .A2(_1863_));
 sg13g2_a21oi_1 _5645_ (.A1(_1812_),
    .A2(_2983_),
    .Y(_1865_),
    .B1(_1196_));
 sg13g2_nand3_1 _5646_ (.B(_2077_),
    .C(_1275_),
    .A(_0950_),
    .Y(_1866_));
 sg13g2_a21oi_1 _5647_ (.A1(_1865_),
    .A2(_1866_),
    .Y(_1867_),
    .B1(_3041_));
 sg13g2_nand2_1 _5648_ (.Y(_1868_),
    .A(_1864_),
    .B(_1867_));
 sg13g2_nand3_1 _5649_ (.B(_0139_),
    .C(_2575_),
    .A(_1070_),
    .Y(_1869_));
 sg13g2_a21oi_1 _5650_ (.A1(_2922_),
    .A2(net106),
    .Y(_1870_),
    .B1(_0272_));
 sg13g2_nand2_1 _5651_ (.Y(_1871_),
    .A(_1869_),
    .B(_1870_));
 sg13g2_nand2_1 _5652_ (.Y(_1873_),
    .A(net56),
    .B(_0917_));
 sg13g2_nand4_1 _5653_ (.B(_1853_),
    .C(_1873_),
    .A(_1674_),
    .Y(_1874_),
    .D(_2840_));
 sg13g2_nand3_1 _5654_ (.B(_1874_),
    .C(_3042_),
    .A(_1871_),
    .Y(_1875_));
 sg13g2_a21o_1 _5655_ (.A2(_1875_),
    .A1(_1868_),
    .B1(_2751_),
    .X(_1876_));
 sg13g2_nand3_1 _5656_ (.B(_1876_),
    .C(_0495_),
    .A(_1858_),
    .Y(_1877_));
 sg13g2_nand2_1 _5657_ (.Y(_0019_),
    .A(_1841_),
    .B(_1877_));
 sg13g2_nand3_1 _5658_ (.B(_3055_),
    .C(_0159_),
    .A(_0177_),
    .Y(_1878_));
 sg13g2_o21ai_1 _5659_ (.B1(_1878_),
    .Y(_1879_),
    .A1(_2724_),
    .A2(_1029_));
 sg13g2_nand2_1 _5660_ (.Y(_1880_),
    .A(_0331_),
    .B(_0977_));
 sg13g2_nand3_1 _5661_ (.B(net137),
    .C(_2973_),
    .A(_0702_),
    .Y(_1881_));
 sg13g2_nand3_1 _5662_ (.B(net144),
    .C(_1881_),
    .A(_1880_),
    .Y(_1883_));
 sg13g2_o21ai_1 _5663_ (.B1(_1883_),
    .Y(_1884_),
    .A1(net136),
    .A2(_1879_));
 sg13g2_nand2_1 _5664_ (.Y(_1885_),
    .A(_1884_),
    .B(net140));
 sg13g2_o21ai_1 _5665_ (.B1(net92),
    .Y(_1886_),
    .A1(_1231_),
    .A2(_2911_));
 sg13g2_o21ai_1 _5666_ (.B1(_1886_),
    .Y(_1887_),
    .A1(_2035_),
    .A2(_0953_));
 sg13g2_nand2_1 _5667_ (.Y(_1888_),
    .A(_1887_),
    .B(_0549_));
 sg13g2_nand2_1 _5668_ (.Y(_1889_),
    .A(_1885_),
    .B(_1888_));
 sg13g2_nand2_1 _5669_ (.Y(_1890_),
    .A(_1889_),
    .B(net190));
 sg13g2_nand2_1 _5670_ (.Y(_1891_),
    .A(_2384_),
    .B(net154));
 sg13g2_nand3_1 _5671_ (.B(_2762_),
    .C(_0917_),
    .A(_1891_),
    .Y(_1892_));
 sg13g2_nand2_1 _5672_ (.Y(_1894_),
    .A(_1811_),
    .B(_2735_));
 sg13g2_nand3_1 _5673_ (.B(net217),
    .C(_1894_),
    .A(_1892_),
    .Y(_1895_));
 sg13g2_nand2_1 _5674_ (.Y(_1896_),
    .A(_1675_),
    .B(net178));
 sg13g2_a21oi_1 _5675_ (.A1(_1028_),
    .A2(_1896_),
    .Y(_1897_),
    .B1(_1173_));
 sg13g2_nor2_1 _5676_ (.A(_1895_),
    .B(_1897_),
    .Y(_1898_));
 sg13g2_nor2_1 _5677_ (.A(_2412_),
    .B(_1898_),
    .Y(_1899_));
 sg13g2_o21ai_1 _5678_ (.B1(net90),
    .Y(_1900_),
    .A1(_0229_),
    .A2(_0337_));
 sg13g2_a21oi_1 _5679_ (.A1(_2689_),
    .A2(net175),
    .Y(_1901_),
    .B1(_2478_));
 sg13g2_nor3_1 _5680_ (.A(_2779_),
    .B(_1901_),
    .C(_1259_),
    .Y(_1902_));
 sg13g2_nand2_1 _5681_ (.Y(_1903_),
    .A(_1900_),
    .B(_1902_));
 sg13g2_nand2_1 _5682_ (.Y(_1905_),
    .A(_1899_),
    .B(_1903_));
 sg13g2_nand2_1 _5683_ (.Y(_1906_),
    .A(_0546_),
    .B(_2077_));
 sg13g2_nand3_1 _5684_ (.B(_2431_),
    .C(_2775_),
    .A(_2825_),
    .Y(_1907_));
 sg13g2_nand3_1 _5685_ (.B(net191),
    .C(_1907_),
    .A(_1906_),
    .Y(_1908_));
 sg13g2_a221oi_1 _5686_ (.B2(_0578_),
    .C1(net203),
    .B1(_0577_),
    .A1(_1205_),
    .Y(_1909_),
    .A2(net124));
 sg13g2_nand2_1 _5687_ (.Y(_1910_),
    .A(_1908_),
    .B(_1909_));
 sg13g2_o21ai_1 _5688_ (.B1(net127),
    .Y(_1911_),
    .A1(_0176_),
    .A2(_1765_));
 sg13g2_nor3_1 _5689_ (.A(_1301_),
    .B(_2871_),
    .C(_2980_),
    .Y(_1912_));
 sg13g2_nor2_1 _5690_ (.A(_1196_),
    .B(_1912_),
    .Y(_1913_));
 sg13g2_a21oi_1 _5691_ (.A1(_1911_),
    .A2(_1913_),
    .Y(_1914_),
    .B1(_2592_));
 sg13g2_nand2_1 _5692_ (.Y(_1916_),
    .A(_1910_),
    .B(_1914_));
 sg13g2_nand2_1 _5693_ (.Y(_1917_),
    .A(_1905_),
    .B(_1916_));
 sg13g2_a21oi_1 _5694_ (.A1(_1040_),
    .A2(_0745_),
    .Y(_1918_),
    .B1(net84));
 sg13g2_a21oi_1 _5695_ (.A1(net65),
    .A2(_0353_),
    .Y(_1919_),
    .B1(net122));
 sg13g2_nand2_1 _5696_ (.Y(_1920_),
    .A(_1919_),
    .B(_1412_));
 sg13g2_nand3_1 _5697_ (.B(_1741_),
    .C(net102),
    .A(_1460_),
    .Y(_1921_));
 sg13g2_nand2_1 _5698_ (.Y(_1922_),
    .A(_1921_),
    .B(net193));
 sg13g2_a21oi_1 _5699_ (.A1(_1918_),
    .A2(_1920_),
    .Y(_1923_),
    .B1(_1922_));
 sg13g2_nand2_1 _5700_ (.Y(_1924_),
    .A(_2623_),
    .B(_0300_));
 sg13g2_nand2_1 _5701_ (.Y(_1925_),
    .A(_1924_),
    .B(_1772_));
 sg13g2_nand3_1 _5702_ (.B(net124),
    .C(_2828_),
    .A(_1251_),
    .Y(_1927_));
 sg13g2_nand2_1 _5703_ (.Y(_1928_),
    .A(_1927_),
    .B(net145));
 sg13g2_a21oi_1 _5704_ (.A1(_1925_),
    .A2(net49),
    .Y(_1929_),
    .B1(_1928_));
 sg13g2_nor3_1 _5705_ (.A(_2949_),
    .B(_1923_),
    .C(_1929_),
    .Y(_1930_));
 sg13g2_a21oi_1 _5706_ (.A1(_1917_),
    .A2(net183),
    .Y(_1931_),
    .B1(_1930_));
 sg13g2_nand2_1 _5707_ (.Y(_1932_),
    .A(_1890_),
    .B(_1931_));
 sg13g2_nand2_1 _5708_ (.Y(_1933_),
    .A(_1932_),
    .B(net212));
 sg13g2_nand2_1 _5709_ (.Y(_1934_),
    .A(_0429_),
    .B(net101));
 sg13g2_nand2_1 _5710_ (.Y(_1935_),
    .A(_1934_),
    .B(_2725_));
 sg13g2_nand3_1 _5711_ (.B(_2432_),
    .C(_1244_),
    .A(_1935_),
    .Y(_1936_));
 sg13g2_o21ai_1 _5712_ (.B1(net54),
    .Y(_1938_),
    .A1(_2585_),
    .A2(_2965_));
 sg13g2_a21oi_1 _5713_ (.A1(_2786_),
    .A2(net99),
    .Y(_1939_),
    .B1(net192));
 sg13g2_nand3_1 _5714_ (.B(_1938_),
    .C(_1939_),
    .A(_1936_),
    .Y(_1940_));
 sg13g2_nand3_1 _5715_ (.B(net163),
    .C(net129),
    .A(_1064_),
    .Y(_1941_));
 sg13g2_nand2_1 _5716_ (.Y(_1942_),
    .A(_2560_),
    .B(_2386_));
 sg13g2_nand4_1 _5717_ (.B(net116),
    .C(_1942_),
    .A(_1941_),
    .Y(_1943_),
    .D(_1789_));
 sg13g2_a21oi_1 _5718_ (.A1(_1500_),
    .A2(_2445_),
    .Y(_1944_),
    .B1(_1173_));
 sg13g2_nor2_1 _5719_ (.A(_1944_),
    .B(_1709_),
    .Y(_1945_));
 sg13g2_a21oi_1 _5720_ (.A1(_1943_),
    .A2(_1945_),
    .Y(_1946_),
    .B1(_3041_));
 sg13g2_nand2_1 _5721_ (.Y(_1947_),
    .A(_1940_),
    .B(_1946_));
 sg13g2_nand2_1 _5722_ (.Y(_1949_),
    .A(_1413_),
    .B(_2397_));
 sg13g2_a21oi_1 _5723_ (.A1(_1949_),
    .A2(net85),
    .Y(_1950_),
    .B1(_1368_));
 sg13g2_o21ai_1 _5724_ (.B1(_1950_),
    .Y(_1951_),
    .A1(_2563_),
    .A2(_1375_));
 sg13g2_a21oi_1 _5725_ (.A1(_1951_),
    .A2(net86),
    .Y(_1952_),
    .B1(net218));
 sg13g2_and2_1 _5726_ (.A(_1947_),
    .B(_1952_),
    .X(_1953_));
 sg13g2_a22oi_1 _5727_ (.Y(_1954_),
    .B1(_2490_),
    .B2(_0687_),
    .A2(_1363_),
    .A1(_2488_));
 sg13g2_nand2_1 _5728_ (.Y(_1955_),
    .A(_0635_),
    .B(net104));
 sg13g2_a221oi_1 _5729_ (.B2(_0836_),
    .C1(_2423_),
    .B1(_1955_),
    .A1(net76),
    .Y(_1956_),
    .A2(net117));
 sg13g2_nor2_1 _5730_ (.A(_2469_),
    .B(_1956_),
    .Y(_1957_));
 sg13g2_o21ai_1 _5731_ (.B1(_1957_),
    .Y(_1958_),
    .A1(_0194_),
    .A2(_1954_));
 sg13g2_a21oi_1 _5732_ (.A1(_1953_),
    .A2(_1958_),
    .Y(_1960_),
    .B1(net212));
 sg13g2_nand3_1 _5733_ (.B(net157),
    .C(_2885_),
    .A(_2807_),
    .Y(_1961_));
 sg13g2_nand3_1 _5734_ (.B(net119),
    .C(_2762_),
    .A(_1741_),
    .Y(_1962_));
 sg13g2_nand3_1 _5735_ (.B(_0260_),
    .C(_1962_),
    .A(_1961_),
    .Y(_1963_));
 sg13g2_a21oi_1 _5736_ (.A1(_1347_),
    .A2(_1741_),
    .Y(_1964_),
    .B1(_0140_));
 sg13g2_nand2_1 _5737_ (.Y(_1965_),
    .A(_1157_),
    .B(_0510_));
 sg13g2_nand2_1 _5738_ (.Y(_1966_),
    .A(_1964_),
    .B(_1965_));
 sg13g2_a21oi_1 _5739_ (.A1(_1963_),
    .A2(_1966_),
    .Y(_1967_),
    .B1(_2629_));
 sg13g2_o21ai_1 _5740_ (.B1(_0700_),
    .Y(_1968_),
    .A1(_1308_),
    .A2(_0750_));
 sg13g2_a21oi_1 _5741_ (.A1(_2863_),
    .A2(_2474_),
    .Y(_1969_),
    .B1(_2585_));
 sg13g2_nor3_1 _5742_ (.A(_0149_),
    .B(_3045_),
    .C(_1969_),
    .Y(_1971_));
 sg13g2_a21oi_1 _5743_ (.A1(_1968_),
    .A2(_2406_),
    .Y(_1972_),
    .B1(_1971_));
 sg13g2_nand2b_1 _5744_ (.Y(_1973_),
    .B(_1972_),
    .A_N(_1967_));
 sg13g2_nand2_1 _5745_ (.Y(_1974_),
    .A(_1973_),
    .B(_2414_));
 sg13g2_a21oi_1 _5746_ (.A1(_2434_),
    .A2(net71),
    .Y(_1975_),
    .B1(_1942_));
 sg13g2_a21oi_1 _5747_ (.A1(_0461_),
    .A2(_0662_),
    .Y(_1976_),
    .B1(_2378_));
 sg13g2_nor2_1 _5748_ (.A(_1975_),
    .B(_1976_),
    .Y(_1977_));
 sg13g2_nor2b_1 _5749_ (.A(_1977_),
    .B_N(_0983_),
    .Y(_1978_));
 sg13g2_a22oi_1 _5750_ (.Y(_1979_),
    .B1(_1028_),
    .B2(_1161_),
    .A2(_0177_),
    .A1(_2939_));
 sg13g2_nand2_1 _5751_ (.Y(_1980_),
    .A(_1979_),
    .B(net171));
 sg13g2_nand2_1 _5752_ (.Y(_1982_),
    .A(_1193_),
    .B(_2588_));
 sg13g2_o21ai_1 _5753_ (.B1(_1982_),
    .Y(_1983_),
    .A1(_2628_),
    .A2(_2508_));
 sg13g2_nand2_1 _5754_ (.Y(_1984_),
    .A(_0800_),
    .B(net77));
 sg13g2_nand3_1 _5755_ (.B(_1670_),
    .C(_2727_),
    .A(_1984_),
    .Y(_1985_));
 sg13g2_nand2_1 _5756_ (.Y(_1986_),
    .A(_1983_),
    .B(_1985_));
 sg13g2_a21oi_1 _5757_ (.A1(_1980_),
    .A2(_1986_),
    .Y(_1987_),
    .B1(_2749_));
 sg13g2_nor3_1 _5758_ (.A(net188),
    .B(_1978_),
    .C(_1987_),
    .Y(_1988_));
 sg13g2_nand2_1 _5759_ (.Y(_1989_),
    .A(_1974_),
    .B(_1988_));
 sg13g2_nand2_1 _5760_ (.Y(_1990_),
    .A(_1960_),
    .B(_1989_));
 sg13g2_nand2_1 _5761_ (.Y(_0020_),
    .A(_1933_),
    .B(_1990_));
 sg13g2_buf_2 _5762_ (.A(ui_in[3]),
    .X(_1992_));
 sg13g2_inv_1 _5763_ (.Y(_1993_),
    .A(_1992_));
 sg13g2_buf_2 _5764_ (.A(ui_in[2]),
    .X(_1994_));
 sg13g2_buf_1 _5765_ (.A(_1994_),
    .X(_1995_));
 sg13g2_buf_1 _5766_ (.A(ui_in[1]),
    .X(_1996_));
 sg13g2_nand2_1 _5767_ (.Y(_1997_),
    .A(net20),
    .B(net240));
 sg13g2_inv_1 _5768_ (.Y(_1998_),
    .A(_1997_));
 sg13g2_nor2_1 _5769_ (.A(net237),
    .B(_1998_),
    .Y(_1999_));
 sg13g2_nor2_1 _5770_ (.A(_1993_),
    .B(_1999_),
    .Y(_2000_));
 sg13g2_buf_1 _5771_ (.A(net20),
    .X(_2001_));
 sg13g2_nor2_1 _5772_ (.A(net239),
    .B(_1994_),
    .Y(_2003_));
 sg13g2_inv_2 _5773_ (.Y(_2004_),
    .A(_1994_));
 sg13g2_nor2_1 _5774_ (.A(net240),
    .B(_2004_),
    .Y(_2005_));
 sg13g2_nor2_1 _5775_ (.A(_1992_),
    .B(_2005_),
    .Y(_2006_));
 sg13g2_inv_1 _5776_ (.Y(_2007_),
    .A(_2006_));
 sg13g2_buf_2 _5777_ (.A(ui_in[4]),
    .X(_2008_));
 sg13g2_buf_2 _5778_ (.A(ui_in[5]),
    .X(_2009_));
 sg13g2_inv_2 _5779_ (.Y(_2010_),
    .A(_2009_));
 sg13g2_nor2_1 _5780_ (.A(_2008_),
    .B(_2010_),
    .Y(_2011_));
 sg13g2_buf_2 _5781_ (.A(_2011_),
    .X(_2012_));
 sg13g2_o21ai_1 _5782_ (.B1(_2012_),
    .Y(_2014_),
    .A1(_2003_),
    .A2(_2007_));
 sg13g2_inv_2 _5783_ (.Y(_2015_),
    .A(_2008_));
 sg13g2_nor2_1 _5784_ (.A(net240),
    .B(net237),
    .Y(_2016_));
 sg13g2_nor2_1 _5785_ (.A(_1993_),
    .B(_2016_),
    .Y(_2017_));
 sg13g2_buf_1 _5786_ (.A(_1992_),
    .X(_2018_));
 sg13g2_inv_1 _5787_ (.Y(_2019_),
    .A(_2001_));
 sg13g2_nor2_1 _5788_ (.A(net240),
    .B(_2019_),
    .Y(_2020_));
 sg13g2_nor2_1 _5789_ (.A(_1994_),
    .B(_2020_),
    .Y(_2021_));
 sg13g2_inv_1 _5790_ (.Y(_2022_),
    .A(_2021_));
 sg13g2_nand2_2 _5791_ (.Y(_2023_),
    .A(net239),
    .B(_1994_));
 sg13g2_nand2_1 _5792_ (.Y(_2025_),
    .A(_2022_),
    .B(_2023_));
 sg13g2_nor2_1 _5793_ (.A(net236),
    .B(_2025_),
    .Y(_2026_));
 sg13g2_nor3_1 _5794_ (.A(_2015_),
    .B(_2017_),
    .C(_2026_),
    .Y(_2027_));
 sg13g2_buf_1 _5795_ (.A(_2008_),
    .X(_2028_));
 sg13g2_inv_1 _5796_ (.Y(_2029_),
    .A(_1996_));
 sg13g2_nor2_2 _5797_ (.A(_1994_),
    .B(_2029_),
    .Y(_2030_));
 sg13g2_nor2_1 _5798_ (.A(net236),
    .B(_2030_),
    .Y(_2031_));
 sg13g2_inv_1 _5799_ (.Y(_2032_),
    .A(_2023_));
 sg13g2_nor2_1 _5800_ (.A(_2005_),
    .B(_2032_),
    .Y(_2033_));
 sg13g2_a22oi_1 _5801_ (.Y(_2034_),
    .B1(_2033_),
    .B2(_2000_),
    .A2(_2031_),
    .A1(net239));
 sg13g2_nor2_1 _5802_ (.A(net235),
    .B(_2034_),
    .Y(_2036_));
 sg13g2_o21ai_1 _5803_ (.B1(_2010_),
    .Y(_2037_),
    .A1(_2027_),
    .A2(_2036_));
 sg13g2_o21ai_1 _5804_ (.B1(_2037_),
    .Y(_0000_),
    .A1(_2000_),
    .A2(_2014_));
 sg13g2_nor2_1 _5805_ (.A(net239),
    .B(_2029_),
    .Y(_2038_));
 sg13g2_nor2_1 _5806_ (.A(_2005_),
    .B(_2030_),
    .Y(_2039_));
 sg13g2_nand2_1 _5807_ (.Y(_2040_),
    .A(_1992_),
    .B(net239));
 sg13g2_inv_1 _5808_ (.Y(_2041_),
    .A(_2040_));
 sg13g2_nand2_1 _5809_ (.Y(_2042_),
    .A(_2039_),
    .B(_2041_));
 sg13g2_nand2_1 _5810_ (.Y(_2043_),
    .A(_2042_),
    .B(_2012_));
 sg13g2_nor2_1 _5811_ (.A(net239),
    .B(net240),
    .Y(_2044_));
 sg13g2_nor2_1 _5812_ (.A(_2044_),
    .B(_1998_),
    .Y(_2046_));
 sg13g2_inv_1 _5813_ (.Y(_2047_),
    .A(_2046_));
 sg13g2_nor2_1 _5814_ (.A(_1993_),
    .B(_2047_),
    .Y(_2048_));
 sg13g2_inv_1 _5815_ (.Y(_2049_),
    .A(_2048_));
 sg13g2_nor2_1 _5816_ (.A(_1994_),
    .B(_2019_),
    .Y(_2050_));
 sg13g2_nor3_1 _5817_ (.A(_1992_),
    .B(_2030_),
    .C(_2050_),
    .Y(_2051_));
 sg13g2_nand2_1 _5818_ (.Y(_2052_),
    .A(_2051_),
    .B(_1997_));
 sg13g2_o21ai_1 _5819_ (.B1(_2052_),
    .Y(_2053_),
    .A1(_2003_),
    .A2(_2049_));
 sg13g2_nor2_1 _5820_ (.A(net237),
    .B(_2046_),
    .Y(_2054_));
 sg13g2_buf_1 _5821_ (.A(net236),
    .X(_2055_));
 sg13g2_nand2_1 _5822_ (.Y(_2057_),
    .A(net240),
    .B(net237));
 sg13g2_nand2_1 _5823_ (.Y(_2058_),
    .A(_2023_),
    .B(_2057_));
 sg13g2_a21oi_1 _5824_ (.A1(_2054_),
    .A2(net233),
    .Y(_2059_),
    .B1(_2058_));
 sg13g2_a21oi_1 _5825_ (.A1(_2059_),
    .A2(_2015_),
    .Y(_2060_),
    .B1(_2009_));
 sg13g2_o21ai_1 _5826_ (.B1(_2060_),
    .Y(_2061_),
    .A1(_2015_),
    .A2(_2053_));
 sg13g2_o21ai_1 _5827_ (.B1(_2061_),
    .Y(_0007_),
    .A1(_2038_),
    .A2(_2043_));
 sg13g2_inv_2 _5828_ (.Y(_2062_),
    .A(_2012_));
 sg13g2_nand2_1 _5829_ (.Y(_2063_),
    .A(_2018_),
    .B(_1996_));
 sg13g2_nand2_1 _5830_ (.Y(_2064_),
    .A(_2003_),
    .B(_2063_));
 sg13g2_nand3_1 _5831_ (.B(_2057_),
    .C(_2040_),
    .A(_2064_),
    .Y(_2065_));
 sg13g2_inv_1 _5832_ (.Y(_2067_),
    .A(_2044_));
 sg13g2_nand2_1 _5833_ (.Y(_2068_),
    .A(_2020_),
    .B(_1994_));
 sg13g2_o21ai_1 _5834_ (.B1(_2068_),
    .Y(_2069_),
    .A1(net237),
    .A2(_2067_));
 sg13g2_a21oi_1 _5835_ (.A1(_2069_),
    .A2(_1993_),
    .Y(_2070_),
    .B1(_2008_));
 sg13g2_nor2_1 _5836_ (.A(net237),
    .B(_2038_),
    .Y(_2071_));
 sg13g2_o21ai_1 _5837_ (.B1(net236),
    .Y(_2072_),
    .A1(_2020_),
    .A2(_2071_));
 sg13g2_and2_1 _5838_ (.A(_2070_),
    .B(_2072_),
    .X(_2073_));
 sg13g2_inv_1 _5839_ (.Y(_2074_),
    .A(_2030_));
 sg13g2_nor2_1 _5840_ (.A(net239),
    .B(_2074_),
    .Y(_2075_));
 sg13g2_a21oi_1 _5841_ (.A1(_2047_),
    .A2(net237),
    .Y(_2076_),
    .B1(_2075_));
 sg13g2_buf_1 _5842_ (.A(_1993_),
    .X(_2078_));
 sg13g2_a221oi_1 _5843_ (.B2(net232),
    .C1(_2015_),
    .B1(_2076_),
    .A1(_2019_),
    .Y(_2079_),
    .A2(_2017_));
 sg13g2_o21ai_1 _5844_ (.B1(_2010_),
    .Y(_2080_),
    .A1(_2073_),
    .A2(_2079_));
 sg13g2_o21ai_1 _5845_ (.B1(_2080_),
    .Y(_0008_),
    .A1(_2062_),
    .A2(_2065_));
 sg13g2_nor2_2 _5846_ (.A(_2009_),
    .B(_2015_),
    .Y(_2081_));
 sg13g2_inv_1 _5847_ (.Y(_2082_),
    .A(_2081_));
 sg13g2_inv_1 _5848_ (.Y(_2083_),
    .A(_2054_));
 sg13g2_o21ai_1 _5849_ (.B1(_2083_),
    .Y(_2084_),
    .A1(_2004_),
    .A2(_1998_));
 sg13g2_a22oi_1 _5850_ (.Y(_2085_),
    .B1(_2078_),
    .B2(_2084_),
    .A2(_2048_),
    .A1(_2004_));
 sg13g2_inv_1 _5851_ (.Y(_2086_),
    .A(_2039_));
 sg13g2_nor2_1 _5852_ (.A(_1992_),
    .B(_2003_),
    .Y(_2088_));
 sg13g2_a21o_1 _5853_ (.A2(_2088_),
    .A1(_2086_),
    .B1(_2048_),
    .X(_2089_));
 sg13g2_a21oi_1 _5854_ (.A1(net240),
    .A2(_1995_),
    .Y(_2090_),
    .B1(_1993_));
 sg13g2_inv_1 _5855_ (.Y(_2091_),
    .A(_2050_));
 sg13g2_nor2_1 _5856_ (.A(_2001_),
    .B(_2004_),
    .Y(_2092_));
 sg13g2_nor2_1 _5857_ (.A(_1992_),
    .B(_2092_),
    .Y(_2093_));
 sg13g2_a221oi_1 _5858_ (.B2(_2093_),
    .C1(_2028_),
    .B1(_2039_),
    .A1(_2090_),
    .Y(_2094_),
    .A2(_2091_));
 sg13g2_a22oi_1 _5859_ (.Y(_2095_),
    .B1(_2010_),
    .B2(_2094_),
    .A2(_2012_),
    .A1(_2089_));
 sg13g2_o21ai_1 _5860_ (.B1(_2095_),
    .Y(_0009_),
    .A1(_2082_),
    .A2(_2085_));
 sg13g2_nor2_1 _5861_ (.A(_2029_),
    .B(_2023_),
    .Y(_2096_));
 sg13g2_inv_1 _5862_ (.Y(_2098_),
    .A(_2096_));
 sg13g2_nand2_1 _5863_ (.Y(_2099_),
    .A(_2098_),
    .B(_2018_));
 sg13g2_o21ai_1 _5864_ (.B1(_2099_),
    .Y(_2100_),
    .A1(_2007_),
    .A2(_2075_));
 sg13g2_o21ai_1 _5865_ (.B1(_2093_),
    .Y(_2101_),
    .A1(_1995_),
    .A2(_1998_));
 sg13g2_a21oi_1 _5866_ (.A1(_2049_),
    .A2(_2101_),
    .Y(_2102_),
    .B1(net235));
 sg13g2_a21oi_1 _5867_ (.A1(net235),
    .A2(_2100_),
    .Y(_2103_),
    .B1(_2102_));
 sg13g2_o21ai_1 _5868_ (.B1(_2012_),
    .Y(_2104_),
    .A1(_2020_),
    .A2(_2007_));
 sg13g2_nand3_1 _5869_ (.B(net233),
    .C(_2068_),
    .A(_2083_),
    .Y(_2105_));
 sg13g2_nand2b_1 _5870_ (.Y(_2106_),
    .B(_2105_),
    .A_N(_2104_));
 sg13g2_o21ai_1 _5871_ (.B1(_2106_),
    .Y(_0010_),
    .A1(_2009_),
    .A2(_2103_));
 sg13g2_a21oi_1 _5872_ (.A1(_2017_),
    .A2(_1997_),
    .Y(_2108_),
    .B1(_2008_));
 sg13g2_nor2_1 _5873_ (.A(_2004_),
    .B(_2047_),
    .Y(_2109_));
 sg13g2_nor2_1 _5874_ (.A(net236),
    .B(_2109_),
    .Y(_2110_));
 sg13g2_a21oi_1 _5875_ (.A1(_2110_),
    .A2(_2022_),
    .Y(_2111_),
    .B1(_2041_));
 sg13g2_a22oi_1 _5876_ (.Y(_2112_),
    .B1(net235),
    .B2(_2111_),
    .A2(_2108_),
    .A1(_2007_));
 sg13g2_nand2_1 _5877_ (.Y(_2113_),
    .A(_2091_),
    .B(_2029_));
 sg13g2_a22oi_1 _5878_ (.Y(_2114_),
    .B1(net233),
    .B2(_2113_),
    .A2(_2088_),
    .A1(_2046_));
 sg13g2_nand3_1 _5879_ (.B(_2015_),
    .C(_2009_),
    .A(_2114_),
    .Y(_2115_));
 sg13g2_o21ai_1 _5880_ (.B1(_2115_),
    .Y(_0011_),
    .A1(_2009_),
    .A2(_2112_));
 sg13g2_o21ai_1 _5881_ (.B1(_2055_),
    .Y(_2116_),
    .A1(net239),
    .A2(_2086_));
 sg13g2_nand3_1 _5882_ (.B(_2116_),
    .C(_2009_),
    .A(_2070_),
    .Y(_2118_));
 sg13g2_a21o_1 _5883_ (.A2(_2049_),
    .A1(_2052_),
    .B1(_2082_),
    .X(_2119_));
 sg13g2_nor2_1 _5884_ (.A(_1992_),
    .B(net240),
    .Y(_2120_));
 sg13g2_inv_1 _5885_ (.Y(_2121_),
    .A(_2120_));
 sg13g2_nor2_1 _5886_ (.A(_2008_),
    .B(_2009_),
    .Y(_2122_));
 sg13g2_nand3_1 _5887_ (.B(_2121_),
    .C(_2122_),
    .A(_2074_),
    .Y(_2123_));
 sg13g2_nand3_1 _5888_ (.B(_2119_),
    .C(_2123_),
    .A(_2118_),
    .Y(_0012_));
 sg13g2_a21oi_1 _5889_ (.A1(_2017_),
    .A2(_2010_),
    .Y(_2124_),
    .B1(_2081_));
 sg13g2_o21ai_1 _5890_ (.B1(_1999_),
    .Y(_2125_),
    .A1(net233),
    .A2(_2044_));
 sg13g2_and3_1 _5891_ (.X(_2126_),
    .A(_2125_),
    .B(net235),
    .C(_2098_));
 sg13g2_nand2_1 _5892_ (.Y(_2128_),
    .A(_2004_),
    .B(net236));
 sg13g2_a21oi_1 _5893_ (.A1(_2096_),
    .A2(net236),
    .Y(_2129_),
    .B1(_2062_));
 sg13g2_inv_1 _5894_ (.Y(_2130_),
    .A(_2129_));
 sg13g2_a21oi_1 _5895_ (.A1(net232),
    .A2(_2058_),
    .Y(_2131_),
    .B1(_2130_));
 sg13g2_o21ai_1 _5896_ (.B1(_2131_),
    .Y(_2132_),
    .A1(_2067_),
    .A2(_2128_));
 sg13g2_o21ai_1 _5897_ (.B1(_2132_),
    .Y(_0013_),
    .A1(_2124_),
    .A2(_2126_));
 sg13g2_a21oi_1 _5898_ (.A1(_2058_),
    .A2(_2040_),
    .Y(_2133_),
    .B1(_2090_));
 sg13g2_nor2_1 _5899_ (.A(net237),
    .B(_2067_),
    .Y(_2134_));
 sg13g2_a21oi_1 _5900_ (.A1(_2134_),
    .A2(net232),
    .Y(_2135_),
    .B1(_2082_));
 sg13g2_nand2b_1 _5901_ (.Y(_2136_),
    .B(_2135_),
    .A_N(_2000_));
 sg13g2_o21ai_1 _5902_ (.B1(_2136_),
    .Y(_0014_),
    .A1(_2062_),
    .A2(_2133_));
 sg13g2_a21o_1 _5903_ (.A2(_2081_),
    .A1(_2000_),
    .B1(_2129_),
    .X(_0015_));
 sg13g2_nand2b_1 _5904_ (.Y(_2138_),
    .B(_2091_),
    .A_N(_2063_));
 sg13g2_nor2_1 _5905_ (.A(_2062_),
    .B(_2093_),
    .Y(_2139_));
 sg13g2_nand4_1 _5906_ (.B(_2023_),
    .C(_2057_),
    .A(_2121_),
    .Y(_2140_),
    .D(_2063_));
 sg13g2_o21ai_1 _5907_ (.B1(_2098_),
    .Y(_2141_),
    .A1(_2120_),
    .A2(_2088_));
 sg13g2_nand3_1 _5908_ (.B(net235),
    .C(_2042_),
    .A(_2141_),
    .Y(_2142_));
 sg13g2_o21ai_1 _5909_ (.B1(_2142_),
    .Y(_2143_),
    .A1(_2028_),
    .A2(_2140_));
 sg13g2_a22oi_1 _5910_ (.Y(_0001_),
    .B1(_2010_),
    .B2(_2143_),
    .A2(_2139_),
    .A1(_2138_));
 sg13g2_nor3_1 _5911_ (.A(_2082_),
    .B(_2090_),
    .C(_2110_),
    .Y(_2144_));
 sg13g2_nand2_1 _5912_ (.Y(_2146_),
    .A(_2122_),
    .B(_2040_));
 sg13g2_nor2_1 _5913_ (.A(_2019_),
    .B(_2030_),
    .Y(_2147_));
 sg13g2_nor2_1 _5914_ (.A(_2147_),
    .B(_2007_),
    .Y(_2148_));
 sg13g2_nand3_1 _5915_ (.B(_2044_),
    .C(net233),
    .A(_2081_),
    .Y(_2149_));
 sg13g2_o21ai_1 _5916_ (.B1(_2149_),
    .Y(_2150_),
    .A1(_2146_),
    .A2(_2148_));
 sg13g2_a22oi_1 _5917_ (.Y(_2151_),
    .B1(net233),
    .B2(_2069_),
    .A2(_2031_),
    .A1(_2033_));
 sg13g2_nor2_1 _5918_ (.A(_2062_),
    .B(_2151_),
    .Y(_2152_));
 sg13g2_nor3_1 _5919_ (.A(_2144_),
    .B(_2150_),
    .C(_2152_),
    .Y(_0002_));
 sg13g2_nor2_1 _5920_ (.A(net232),
    .B(_2021_),
    .Y(_2153_));
 sg13g2_inv_1 _5921_ (.Y(_2154_),
    .A(_2109_));
 sg13g2_a22oi_1 _5922_ (.Y(_2156_),
    .B1(_2153_),
    .B2(_2154_),
    .A2(_2032_),
    .A1(net232));
 sg13g2_nand2b_1 _5923_ (.Y(_2157_),
    .B(_2081_),
    .A_N(_2156_));
 sg13g2_nor2_1 _5924_ (.A(net232),
    .B(_2109_),
    .Y(_2158_));
 sg13g2_inv_1 _5925_ (.Y(_2159_),
    .A(_2158_));
 sg13g2_a21oi_1 _5926_ (.A1(_2006_),
    .A2(_1997_),
    .Y(_2160_),
    .B1(_2062_));
 sg13g2_o21ai_1 _5927_ (.B1(_2160_),
    .Y(_2161_),
    .A1(_2134_),
    .A2(_2159_));
 sg13g2_nor2_1 _5928_ (.A(_2153_),
    .B(_2051_),
    .Y(_2162_));
 sg13g2_o21ai_1 _5929_ (.B1(_2122_),
    .Y(_2163_),
    .A1(_2092_),
    .A2(_2162_));
 sg13g2_nand3_1 _5930_ (.B(_2161_),
    .C(_2163_),
    .A(_2157_),
    .Y(_0003_));
 sg13g2_o21ai_1 _5931_ (.B1(_2008_),
    .Y(_2164_),
    .A1(net236),
    .A2(_2004_));
 sg13g2_a21oi_1 _5932_ (.A1(_2025_),
    .A2(net233),
    .Y(_2166_),
    .B1(_2164_));
 sg13g2_nand2b_1 _5933_ (.Y(_2167_),
    .B(_2010_),
    .A_N(_2166_));
 sg13g2_nor3_1 _5934_ (.A(net233),
    .B(_2016_),
    .C(_2109_),
    .Y(_2168_));
 sg13g2_nor3_1 _5935_ (.A(net235),
    .B(_2153_),
    .C(_2168_),
    .Y(_2169_));
 sg13g2_nand3_1 _5936_ (.B(net232),
    .C(_2019_),
    .A(_2039_),
    .Y(_2170_));
 sg13g2_nand3_1 _5937_ (.B(_2170_),
    .C(_2012_),
    .A(_2159_),
    .Y(_2171_));
 sg13g2_o21ai_1 _5938_ (.B1(_2171_),
    .Y(_0004_),
    .A1(_2167_),
    .A2(_2169_));
 sg13g2_nand2_1 _5939_ (.Y(_2172_),
    .A(_2032_),
    .B(_2120_));
 sg13g2_o21ai_1 _5940_ (.B1(_2172_),
    .Y(_2173_),
    .A1(net232),
    .A2(_2067_));
 sg13g2_nand2_1 _5941_ (.Y(_2174_),
    .A(_2173_),
    .B(net235));
 sg13g2_nand3_1 _5942_ (.B(_2015_),
    .C(_2128_),
    .A(_2172_),
    .Y(_2176_));
 sg13g2_nand3_1 _5943_ (.B(_2176_),
    .C(_2010_),
    .A(_2174_),
    .Y(_2177_));
 sg13g2_o21ai_1 _5944_ (.B1(_2055_),
    .Y(_2178_),
    .A1(_2038_),
    .A2(_2147_));
 sg13g2_nand2_1 _5945_ (.Y(_2179_),
    .A(_2113_),
    .B(_2078_));
 sg13g2_nand3_1 _5946_ (.B(_2012_),
    .C(_2179_),
    .A(_2178_),
    .Y(_2180_));
 sg13g2_nand2_1 _5947_ (.Y(_0005_),
    .A(_2177_),
    .B(_2180_));
 sg13g2_o21ai_1 _5948_ (.B1(_2149_),
    .Y(_0006_),
    .A1(_2062_),
    .A2(_2170_));
 sg13g2_inv_1 _5949_ (.Y(_2181_),
    .A(net19));
 sg13g2_buf_1 _5950_ (.A(net238),
    .X(_2182_));
 sg13g2_inv_1 _5951_ (.Y(_2183_),
    .A(\clk_picker.counter[17] ));
 sg13g2_nor3_1 _5952_ (.A(\clk_picker.counter[9] ),
    .B(\clk_picker.counter[10] ),
    .C(\clk_picker.counter[11] ),
    .Y(_2185_));
 sg13g2_inv_1 _5953_ (.Y(_2186_),
    .A(\clk_picker.counter[7] ));
 sg13g2_inv_1 _5954_ (.Y(_2187_),
    .A(\clk_picker.counter[8] ));
 sg13g2_nand3_1 _5955_ (.B(_2186_),
    .C(_2187_),
    .A(_2185_),
    .Y(_2188_));
 sg13g2_inv_1 _5956_ (.Y(_2189_),
    .A(\clk_picker.counter[12] ));
 sg13g2_inv_1 _5957_ (.Y(_2190_),
    .A(\clk_picker.counter[13] ));
 sg13g2_nand2_1 _5958_ (.Y(_2191_),
    .A(\clk_picker.counter[14] ),
    .B(\clk_picker.counter[15] ));
 sg13g2_nor3_1 _5959_ (.A(_2189_),
    .B(_2190_),
    .C(_2191_),
    .Y(_2192_));
 sg13g2_a21oi_1 _5960_ (.A1(_2188_),
    .A2(_2192_),
    .Y(_2193_),
    .B1(\clk_picker.counter[16] ));
 sg13g2_inv_1 _5961_ (.Y(_2194_),
    .A(\clk_picker.counter[18] ));
 sg13g2_o21ai_1 _5962_ (.B1(_2194_),
    .Y(_2196_),
    .A1(_2183_),
    .A2(_2193_));
 sg13g2_nand2_1 _5963_ (.Y(_2197_),
    .A(\clk_picker.counter[20] ),
    .B(\clk_picker.counter[21] ));
 sg13g2_inv_1 _5964_ (.Y(_2198_),
    .A(_2197_));
 sg13g2_and3_1 _5965_ (.X(_2199_),
    .A(_2198_),
    .B(\clk_picker.counter[22] ),
    .C(\clk_picker.counter[23] ));
 sg13g2_nand4_1 _5966_ (.B(\clk_picker.counter[19] ),
    .C(\clk_picker.counter[25] ),
    .A(_2196_),
    .Y(_2200_),
    .D(_2199_));
 sg13g2_inv_1 _5967_ (.Y(_2201_),
    .A(\clk_picker.clk_slow ));
 sg13g2_nand2_1 _5968_ (.Y(_2202_),
    .A(\clk_picker.counter[24] ),
    .B(\clk_picker.counter[25] ));
 sg13g2_and3_1 _5969_ (.X(_2203_),
    .A(_2200_),
    .B(_2201_),
    .C(_2202_));
 sg13g2_and2_1 _5970_ (.A(_2200_),
    .B(_2202_),
    .X(_2204_));
 sg13g2_nor2_1 _5971_ (.A(_0030_),
    .B(_2204_),
    .Y(_2205_));
 sg13g2_nor3_1 _5972_ (.A(_2182_),
    .B(_2203_),
    .C(_2205_),
    .Y(_0040_));
 sg13g2_nand2_1 _5973_ (.Y(_2207_),
    .A(_2204_),
    .B(net19));
 sg13g2_buf_2 _5974_ (.A(_2207_),
    .X(_2208_));
 sg13g2_buf_1 _5975_ (.A(_2208_),
    .X(_2209_));
 sg13g2_nor2b_1 _5976_ (.A(net231),
    .B_N(_0039_),
    .Y(_0041_));
 sg13g2_nand2_1 _5977_ (.Y(_2210_),
    .A(\clk_picker.counter[1] ),
    .B(\clk_picker.counter[0] ));
 sg13g2_nor2b_1 _5978_ (.A(_2210_),
    .B_N(\clk_picker.counter[2] ),
    .Y(_2211_));
 sg13g2_nand2_1 _5979_ (.Y(_2212_),
    .A(_2211_),
    .B(\clk_picker.counter[3] ));
 sg13g2_nor2b_1 _5980_ (.A(_2212_),
    .B_N(\clk_picker.counter[4] ),
    .Y(_2213_));
 sg13g2_nand2_1 _5981_ (.Y(_2214_),
    .A(_2213_),
    .B(\clk_picker.counter[5] ));
 sg13g2_nor2b_1 _5982_ (.A(_2214_),
    .B_N(\clk_picker.counter[6] ),
    .Y(_2216_));
 sg13g2_nand2_1 _5983_ (.Y(_2217_),
    .A(_2216_),
    .B(\clk_picker.counter[7] ));
 sg13g2_nor2_1 _5984_ (.A(_2187_),
    .B(_2217_),
    .Y(_2218_));
 sg13g2_nand2_1 _5985_ (.Y(_2219_),
    .A(_2218_),
    .B(\clk_picker.counter[9] ));
 sg13g2_inv_2 _5986_ (.Y(_2220_),
    .A(_2219_));
 sg13g2_nand2_1 _5987_ (.Y(_2221_),
    .A(_2220_),
    .B(\clk_picker.counter[10] ));
 sg13g2_inv_1 _5988_ (.Y(_2222_),
    .A(_2221_));
 sg13g2_nor2_1 _5989_ (.A(\clk_picker.counter[10] ),
    .B(_2220_),
    .Y(_2223_));
 sg13g2_nor3_1 _5990_ (.A(_2222_),
    .B(_2223_),
    .C(net231),
    .Y(_0042_));
 sg13g2_nor2_1 _5991_ (.A(\clk_picker.counter[11] ),
    .B(_2222_),
    .Y(_2224_));
 sg13g2_nand2_1 _5992_ (.Y(_2226_),
    .A(\clk_picker.counter[10] ),
    .B(\clk_picker.counter[11] ));
 sg13g2_nor2_1 _5993_ (.A(_2226_),
    .B(_2219_),
    .Y(_2227_));
 sg13g2_nor3_1 _5994_ (.A(_2224_),
    .B(_2227_),
    .C(net231),
    .Y(_0043_));
 sg13g2_nor2_1 _5995_ (.A(\clk_picker.counter[12] ),
    .B(_2227_),
    .Y(_2228_));
 sg13g2_nor3_1 _5996_ (.A(_2189_),
    .B(_2226_),
    .C(_2219_),
    .Y(_2229_));
 sg13g2_nor3_1 _5997_ (.A(_2228_),
    .B(_2229_),
    .C(_2209_),
    .Y(_0044_));
 sg13g2_nor2_1 _5998_ (.A(\clk_picker.counter[13] ),
    .B(_2229_),
    .Y(_2230_));
 sg13g2_nand2_1 _5999_ (.Y(_2231_),
    .A(_2229_),
    .B(\clk_picker.counter[13] ));
 sg13g2_inv_1 _6000_ (.Y(_2232_),
    .A(_2231_));
 sg13g2_buf_1 _6001_ (.A(_2208_),
    .X(_2233_));
 sg13g2_nor3_1 _6002_ (.A(_2230_),
    .B(_2232_),
    .C(_2233_),
    .Y(_0045_));
 sg13g2_xor2_1 _6003_ (.B(_2231_),
    .A(\clk_picker.counter[14] ),
    .X(_2235_));
 sg13g2_nor2_1 _6004_ (.A(_2209_),
    .B(_2235_),
    .Y(_0046_));
 sg13g2_and4_1 _6005_ (.A(\clk_picker.counter[11] ),
    .B(\clk_picker.counter[12] ),
    .C(\clk_picker.counter[13] ),
    .D(\clk_picker.counter[14] ),
    .X(_2236_));
 sg13g2_a21oi_1 _6006_ (.A1(_2222_),
    .A2(_2236_),
    .Y(_2237_),
    .B1(\clk_picker.counter[15] ));
 sg13g2_inv_1 _6007_ (.Y(_2238_),
    .A(_2226_));
 sg13g2_nand4_1 _6008_ (.B(\clk_picker.counter[8] ),
    .C(\clk_picker.counter[9] ),
    .A(_2192_),
    .Y(_2239_),
    .D(_2238_));
 sg13g2_nor2_2 _6009_ (.A(_2239_),
    .B(_2217_),
    .Y(_2240_));
 sg13g2_nor3_1 _6010_ (.A(_2237_),
    .B(_2240_),
    .C(net230),
    .Y(_0047_));
 sg13g2_nor2_1 _6011_ (.A(\clk_picker.counter[16] ),
    .B(_2240_),
    .Y(_2241_));
 sg13g2_nand2_1 _6012_ (.Y(_2243_),
    .A(_2240_),
    .B(\clk_picker.counter[16] ));
 sg13g2_inv_1 _6013_ (.Y(_2244_),
    .A(_2243_));
 sg13g2_nor3_1 _6014_ (.A(_2241_),
    .B(_2244_),
    .C(net230),
    .Y(_0048_));
 sg13g2_nor2_1 _6015_ (.A(\clk_picker.counter[17] ),
    .B(_2244_),
    .Y(_2245_));
 sg13g2_nor2_1 _6016_ (.A(_2183_),
    .B(_2243_),
    .Y(_2246_));
 sg13g2_nor3_1 _6017_ (.A(_2245_),
    .B(_2246_),
    .C(_2233_),
    .Y(_0049_));
 sg13g2_nor2_1 _6018_ (.A(\clk_picker.counter[18] ),
    .B(_2246_),
    .Y(_2247_));
 sg13g2_nor3_1 _6019_ (.A(_2183_),
    .B(_2194_),
    .C(_2243_),
    .Y(_2248_));
 sg13g2_nor3_1 _6020_ (.A(_2247_),
    .B(_2248_),
    .C(net230),
    .Y(_0050_));
 sg13g2_xnor2_1 _6021_ (.Y(_2249_),
    .A(\clk_picker.counter[19] ),
    .B(_2248_));
 sg13g2_nor2_1 _6022_ (.A(_2249_),
    .B(net231),
    .Y(_0051_));
 sg13g2_inv_1 _6023_ (.Y(_2251_),
    .A(_2210_));
 sg13g2_nor2_1 _6024_ (.A(\clk_picker.counter[1] ),
    .B(\clk_picker.counter[0] ),
    .Y(_2252_));
 sg13g2_nor3_1 _6025_ (.A(_2251_),
    .B(_2252_),
    .C(net230),
    .Y(_0052_));
 sg13g2_inv_1 _6026_ (.Y(_2253_),
    .A(\clk_picker.counter[16] ));
 sg13g2_nand2_1 _6027_ (.Y(_2254_),
    .A(\clk_picker.counter[18] ),
    .B(\clk_picker.counter[19] ));
 sg13g2_nor3_1 _6028_ (.A(_2253_),
    .B(_2183_),
    .C(_2254_),
    .Y(_2255_));
 sg13g2_a21oi_1 _6029_ (.A1(_2240_),
    .A2(_2255_),
    .Y(_2256_),
    .B1(\clk_picker.counter[20] ));
 sg13g2_nand3_1 _6030_ (.B(\clk_picker.counter[20] ),
    .C(_2255_),
    .A(_2240_),
    .Y(_2257_));
 sg13g2_nand2b_1 _6031_ (.Y(_2258_),
    .B(_2257_),
    .A_N(_2256_));
 sg13g2_nor2_1 _6032_ (.A(_2258_),
    .B(net231),
    .Y(_0053_));
 sg13g2_xor2_1 _6033_ (.B(_2257_),
    .A(\clk_picker.counter[21] ),
    .X(_2260_));
 sg13g2_nor2_1 _6034_ (.A(_2260_),
    .B(net231),
    .Y(_0054_));
 sg13g2_nand3_1 _6035_ (.B(_2198_),
    .C(_2255_),
    .A(_2240_),
    .Y(_2261_));
 sg13g2_nor2b_1 _6036_ (.A(\clk_picker.counter[22] ),
    .B_N(_2261_),
    .Y(_2262_));
 sg13g2_nor2b_1 _6037_ (.A(_2261_),
    .B_N(\clk_picker.counter[22] ),
    .Y(_2263_));
 sg13g2_nor3_1 _6038_ (.A(_2262_),
    .B(_2263_),
    .C(net230),
    .Y(_0055_));
 sg13g2_nand2_1 _6039_ (.Y(_2264_),
    .A(_2263_),
    .B(\clk_picker.counter[23] ));
 sg13g2_inv_2 _6040_ (.Y(_2265_),
    .A(_2264_));
 sg13g2_nor2_1 _6041_ (.A(\clk_picker.counter[23] ),
    .B(_2263_),
    .Y(_2266_));
 sg13g2_nor3_1 _6042_ (.A(_2265_),
    .B(_2266_),
    .C(net230),
    .Y(_0056_));
 sg13g2_xor2_1 _6043_ (.B(_2264_),
    .A(\clk_picker.counter[24] ),
    .X(_2268_));
 sg13g2_nor2_1 _6044_ (.A(net231),
    .B(_2268_),
    .Y(_0057_));
 sg13g2_a21oi_1 _6045_ (.A1(_2265_),
    .A2(\clk_picker.counter[24] ),
    .Y(_2269_),
    .B1(\clk_picker.counter[25] ));
 sg13g2_nor2_1 _6046_ (.A(net231),
    .B(_2269_),
    .Y(_0058_));
 sg13g2_nor2_1 _6047_ (.A(\clk_picker.counter[2] ),
    .B(_2251_),
    .Y(_2270_));
 sg13g2_nor3_1 _6048_ (.A(_2211_),
    .B(_2270_),
    .C(net230),
    .Y(_0059_));
 sg13g2_inv_1 _6049_ (.Y(_2271_),
    .A(_2212_));
 sg13g2_nor2_1 _6050_ (.A(\clk_picker.counter[3] ),
    .B(_2211_),
    .Y(_2272_));
 sg13g2_nor3_1 _6051_ (.A(_2271_),
    .B(_2272_),
    .C(net230),
    .Y(_0060_));
 sg13g2_nor2_1 _6052_ (.A(\clk_picker.counter[4] ),
    .B(_2271_),
    .Y(_2274_));
 sg13g2_nor3_1 _6053_ (.A(_2213_),
    .B(_2274_),
    .C(_2208_),
    .Y(_0061_));
 sg13g2_inv_1 _6054_ (.Y(_2275_),
    .A(_2214_));
 sg13g2_nor2_1 _6055_ (.A(\clk_picker.counter[5] ),
    .B(_2213_),
    .Y(_2276_));
 sg13g2_nor3_1 _6056_ (.A(_2275_),
    .B(_2276_),
    .C(_2208_),
    .Y(_0062_));
 sg13g2_nor2_1 _6057_ (.A(\clk_picker.counter[6] ),
    .B(_2275_),
    .Y(_2277_));
 sg13g2_nor3_1 _6058_ (.A(_2216_),
    .B(_2277_),
    .C(_2208_),
    .Y(_0063_));
 sg13g2_inv_1 _6059_ (.Y(_2278_),
    .A(_2217_));
 sg13g2_nor2_1 _6060_ (.A(\clk_picker.counter[7] ),
    .B(_2216_),
    .Y(_2279_));
 sg13g2_nor3_1 _6061_ (.A(_2278_),
    .B(_2279_),
    .C(_2208_),
    .Y(_0064_));
 sg13g2_nor2_1 _6062_ (.A(\clk_picker.counter[8] ),
    .B(_2278_),
    .Y(_2281_));
 sg13g2_nor3_1 _6063_ (.A(_2218_),
    .B(_2281_),
    .C(_2208_),
    .Y(_0065_));
 sg13g2_nor2_1 _6064_ (.A(\clk_picker.counter[9] ),
    .B(_2218_),
    .Y(_2282_));
 sg13g2_nor3_1 _6065_ (.A(_2220_),
    .B(_2282_),
    .C(_2208_),
    .Y(_0066_));
 sg13g2_nor2_1 _6066_ (.A(net21),
    .B(\transformer_1.started ),
    .Y(_2283_));
 sg13g2_buf_1 _6067_ (.A(_2283_),
    .X(_2284_));
 sg13g2_nor2_1 _6068_ (.A(_0031_),
    .B(_2284_),
    .Y(_2285_));
 sg13g2_inv_1 _6069_ (.Y(_2286_),
    .A(_2284_));
 sg13g2_nor2_1 _6070_ (.A(\line_mapper_1.pointer_addr[10] ),
    .B(_2286_),
    .Y(_2287_));
 sg13g2_or2_1 _6071_ (.X(_2288_),
    .B(\chars_remaining[1] ),
    .A(\chars_remaining[2] ));
 sg13g2_nor2_1 _6072_ (.A(\chars_remaining[0] ),
    .B(_2288_),
    .Y(_2290_));
 sg13g2_inv_2 _6073_ (.Y(_2291_),
    .A(_2290_));
 sg13g2_nor2_1 _6074_ (.A(\chars_remaining[3] ),
    .B(_2291_),
    .Y(_2292_));
 sg13g2_inv_1 _6075_ (.Y(_2293_),
    .A(\chars_remaining[4] ));
 sg13g2_nand2_1 _6076_ (.Y(_2294_),
    .A(_2292_),
    .B(_2293_));
 sg13g2_nor2_1 _6077_ (.A(\chars_remaining[5] ),
    .B(_2294_),
    .Y(_2295_));
 sg13g2_nor4_2 _6078_ (.A(\chars_remaining[9] ),
    .B(\chars_remaining[8] ),
    .C(\chars_remaining[7] ),
    .Y(_2296_),
    .D(\chars_remaining[6] ));
 sg13g2_nand2_1 _6079_ (.Y(_2297_),
    .A(_2295_),
    .B(_2296_));
 sg13g2_nor2_1 _6080_ (.A(net211),
    .B(_2297_),
    .Y(_2298_));
 sg13g2_buf_1 _6081_ (.A(_2298_),
    .X(_2299_));
 sg13g2_nor4_1 _6082_ (.A(net234),
    .B(_2285_),
    .C(_2287_),
    .D(net38),
    .Y(_0067_));
 sg13g2_buf_1 _6083_ (.A(net211),
    .X(_2301_));
 sg13g2_xnor2_1 _6084_ (.Y(_2302_),
    .A(\chars_remaining[0] ),
    .B(\chars_remaining[1] ));
 sg13g2_nand2_2 _6085_ (.Y(_2303_),
    .A(_2297_),
    .B(_2286_));
 sg13g2_inv_1 _6086_ (.Y(_2304_),
    .A(_2303_));
 sg13g2_buf_1 _6087_ (.A(_2304_),
    .X(_2305_));
 sg13g2_a22oi_1 _6088_ (.Y(_2306_),
    .B1(_2302_),
    .B2(net37),
    .A2(_2301_),
    .A1(\line_mapper_1.pointer_addr[11] ));
 sg13g2_nor2_1 _6089_ (.A(net234),
    .B(_2306_),
    .Y(_0068_));
 sg13g2_o21ai_1 _6090_ (.B1(\chars_remaining[2] ),
    .Y(_2307_),
    .A1(\chars_remaining[0] ),
    .A2(\chars_remaining[1] ));
 sg13g2_nand2_1 _6091_ (.Y(_2308_),
    .A(_2291_),
    .B(_2307_));
 sg13g2_a22oi_1 _6092_ (.Y(_2310_),
    .B1(_2308_),
    .B2(net37),
    .A2(_2301_),
    .A1(\line_mapper_1.pointer_addr[12] ));
 sg13g2_nor2_1 _6093_ (.A(net234),
    .B(_2310_),
    .Y(_0069_));
 sg13g2_inv_1 _6094_ (.Y(_2311_),
    .A(\chars_remaining[3] ));
 sg13g2_nor2_1 _6095_ (.A(_2311_),
    .B(_2290_),
    .Y(_2312_));
 sg13g2_o21ai_1 _6096_ (.B1(net37),
    .Y(_2313_),
    .A1(_2292_),
    .A2(_2312_));
 sg13g2_nand2_1 _6097_ (.Y(_2314_),
    .A(net181),
    .B(\line_mapper_1.pointer_addr[13] ));
 sg13g2_a21oi_1 _6098_ (.A1(_2313_),
    .A2(_2314_),
    .Y(_0070_),
    .B1(net234));
 sg13g2_o21ai_1 _6099_ (.B1(\chars_remaining[4] ),
    .Y(_2315_),
    .A1(\chars_remaining[3] ),
    .A2(_2291_));
 sg13g2_a21o_1 _6100_ (.A2(_2315_),
    .A1(_2294_),
    .B1(_2303_),
    .X(_2316_));
 sg13g2_nand2_1 _6101_ (.Y(_2317_),
    .A(net181),
    .B(\line_mapper_1.pointer_addr[14] ));
 sg13g2_a21oi_1 _6102_ (.A1(_2316_),
    .A2(_2317_),
    .Y(_0071_),
    .B1(net234));
 sg13g2_nor3_1 _6103_ (.A(\chars_remaining[4] ),
    .B(\chars_remaining[3] ),
    .C(_2288_),
    .Y(_2319_));
 sg13g2_nand2_1 _6104_ (.Y(_2320_),
    .A(_2319_),
    .B(_0031_));
 sg13g2_xnor2_1 _6105_ (.Y(_2321_),
    .A(\chars_remaining[5] ),
    .B(_2320_));
 sg13g2_a22oi_1 _6106_ (.Y(_2322_),
    .B1(_2321_),
    .B2(net37),
    .A2(net181),
    .A1(\line_mapper_1.pointer_addr[15] ));
 sg13g2_nor2_1 _6107_ (.A(_2182_),
    .B(_2322_),
    .Y(_0072_));
 sg13g2_inv_1 _6108_ (.Y(_2323_),
    .A(_2295_));
 sg13g2_o21ai_1 _6109_ (.B1(\chars_remaining[6] ),
    .Y(_2324_),
    .A1(_2296_),
    .A2(_2323_));
 sg13g2_nor2_1 _6110_ (.A(_2296_),
    .B(_2323_),
    .Y(_2325_));
 sg13g2_nand2b_1 _6111_ (.Y(_2326_),
    .B(_2325_),
    .A_N(\chars_remaining[6] ));
 sg13g2_nor2_1 _6112_ (.A(net238),
    .B(net211),
    .Y(_2328_));
 sg13g2_inv_1 _6113_ (.Y(_2329_),
    .A(_2328_));
 sg13g2_a21oi_1 _6114_ (.A1(_2324_),
    .A2(_2326_),
    .Y(_0073_),
    .B1(_2329_));
 sg13g2_or2_1 _6115_ (.X(_2330_),
    .B(_2326_),
    .A(\chars_remaining[7] ));
 sg13g2_buf_1 _6116_ (.A(_2330_),
    .X(_2331_));
 sg13g2_nand2_1 _6117_ (.Y(_2332_),
    .A(_2326_),
    .B(\chars_remaining[7] ));
 sg13g2_a21oi_1 _6118_ (.A1(_2331_),
    .A2(_2332_),
    .Y(_0074_),
    .B1(_2329_));
 sg13g2_inv_1 _6119_ (.Y(_2333_),
    .A(\chars_remaining[8] ));
 sg13g2_o21ai_1 _6120_ (.B1(_2328_),
    .Y(_2334_),
    .A1(_2333_),
    .A2(_2331_));
 sg13g2_a21oi_1 _6121_ (.A1(_2333_),
    .A2(_2331_),
    .Y(_0075_),
    .B1(_2334_));
 sg13g2_inv_1 _6122_ (.Y(_2336_),
    .A(\chars_remaining[9] ));
 sg13g2_nor4_1 _6123_ (.A(\chars_remaining[8] ),
    .B(\chars_remaining[7] ),
    .C(\chars_remaining[6] ),
    .D(_2323_),
    .Y(_2337_));
 sg13g2_nor3_1 _6124_ (.A(_2336_),
    .B(_2329_),
    .C(_2337_),
    .Y(_0076_));
 sg13g2_nand2_1 _6125_ (.Y(_2338_),
    .A(net37),
    .B(_2300_));
 sg13g2_nand2_1 _6126_ (.Y(_2339_),
    .A(net38),
    .B(net222));
 sg13g2_a21oi_1 _6127_ (.A1(net181),
    .A2(\line_mapper_1.pointer_addr[0] ),
    .Y(_2340_),
    .B1(net238));
 sg13g2_nand3_1 _6128_ (.B(_2339_),
    .C(_2340_),
    .A(_2338_),
    .Y(_0077_));
 sg13g2_a221oi_1 _6129_ (.B2(net200),
    .C1(_2181_),
    .B1(net38),
    .A1(\line_mapper_1.pointer_addr[1] ),
    .Y(_2341_),
    .A2(net211));
 sg13g2_o21ai_1 _6130_ (.B1(_2341_),
    .Y(_0078_),
    .A1(net41),
    .A2(_2303_));
 sg13g2_nand2_1 _6131_ (.Y(_2342_),
    .A(net37),
    .B(_2942_));
 sg13g2_nand2_1 _6132_ (.Y(_2344_),
    .A(net38),
    .B(_2379_));
 sg13g2_a21oi_1 _6133_ (.A1(net181),
    .A2(\line_mapper_1.pointer_addr[2] ),
    .Y(_2345_),
    .B1(net238));
 sg13g2_nand3_1 _6134_ (.B(_2344_),
    .C(_2345_),
    .A(_2342_),
    .Y(_0079_));
 sg13g2_nor2_1 _6135_ (.A(_2300_),
    .B(net175),
    .Y(_2346_));
 sg13g2_xnor2_1 _6136_ (.Y(_2347_),
    .A(net39),
    .B(_2346_));
 sg13g2_a22oi_1 _6137_ (.Y(_2348_),
    .B1(_2347_),
    .B2(_2305_),
    .A2(net71),
    .A1(_2299_));
 sg13g2_a21oi_1 _6138_ (.A1(net181),
    .A2(\line_mapper_1.pointer_addr[3] ),
    .Y(_2349_),
    .B1(net234));
 sg13g2_nand2_1 _6139_ (.Y(_0080_),
    .A(_2348_),
    .B(_2349_));
 sg13g2_xnor2_1 _6140_ (.Y(_2350_),
    .A(net105),
    .B(_1557_));
 sg13g2_nand2_1 _6141_ (.Y(_2351_),
    .A(_2305_),
    .B(_2350_));
 sg13g2_nand2_1 _6142_ (.Y(_2353_),
    .A(_2299_),
    .B(net105));
 sg13g2_a21oi_1 _6143_ (.A1(net211),
    .A2(\line_mapper_1.pointer_addr[4] ),
    .Y(_2354_),
    .B1(net238));
 sg13g2_nand3_1 _6144_ (.B(_2353_),
    .C(_2354_),
    .A(_2351_),
    .Y(_0081_));
 sg13g2_nand2_1 _6145_ (.Y(_2355_),
    .A(_2972_),
    .B(net120));
 sg13g2_nor2_1 _6146_ (.A(net49),
    .B(_2355_),
    .Y(_2356_));
 sg13g2_nand2_1 _6147_ (.Y(_2357_),
    .A(_2355_),
    .B(net49));
 sg13g2_nand3b_1 _6148_ (.B(_2304_),
    .C(_2357_),
    .Y(_2358_),
    .A_N(_2356_));
 sg13g2_nand2_1 _6149_ (.Y(_2359_),
    .A(net38),
    .B(net135));
 sg13g2_a21oi_1 _6150_ (.A1(net211),
    .A2(\line_mapper_1.pointer_addr[5] ),
    .Y(_2360_),
    .B1(net238));
 sg13g2_nand3_1 _6151_ (.B(_2359_),
    .C(_2360_),
    .A(_2358_),
    .Y(_0082_));
 sg13g2_xnor2_1 _6152_ (.Y(_2362_),
    .A(net55),
    .B(_2356_));
 sg13g2_a22oi_1 _6153_ (.Y(_2363_),
    .B1(_2362_),
    .B2(net37),
    .A2(net156),
    .A1(net38));
 sg13g2_a21oi_1 _6154_ (.A1(net181),
    .A2(\line_mapper_1.pointer_addr[6] ),
    .Y(_2364_),
    .B1(net234));
 sg13g2_nand2_1 _6155_ (.Y(_0083_),
    .A(_2363_),
    .B(_2364_));
 sg13g2_nand4_1 _6156_ (.B(_1636_),
    .C(_3014_),
    .A(_2297_),
    .Y(_2365_),
    .D(_2782_));
 sg13g2_nor2b_1 _6157_ (.A(net138),
    .B_N(_2365_),
    .Y(_2366_));
 sg13g2_o21ai_1 _6158_ (.B1(_2286_),
    .Y(_2367_),
    .A1(_2414_),
    .A2(_2365_));
 sg13g2_a21oi_1 _6159_ (.A1(net181),
    .A2(\line_mapper_1.pointer_addr[7] ),
    .Y(_2368_),
    .B1(net238));
 sg13g2_o21ai_1 _6160_ (.B1(_2368_),
    .Y(_0084_),
    .A1(_2366_),
    .A2(_2367_));
 sg13g2_nand2_1 _6161_ (.Y(_2369_),
    .A(_2356_),
    .B(net86));
 sg13g2_xnor2_1 _6162_ (.Y(_2371_),
    .A(net194),
    .B(_2369_));
 sg13g2_a221oi_1 _6163_ (.B2(net190),
    .C1(net238),
    .B1(net38),
    .A1(\line_mapper_1.pointer_addr[8] ),
    .Y(_2372_),
    .A2(net211));
 sg13g2_o21ai_1 _6164_ (.B1(_2372_),
    .Y(_0085_),
    .A1(_2303_),
    .A2(_2371_));
 sg13g2_nand3_1 _6165_ (.B(_2782_),
    .C(_2848_),
    .A(_2972_),
    .Y(_2373_));
 sg13g2_xnor2_1 _6166_ (.Y(_2374_),
    .A(net182),
    .B(_2373_));
 sg13g2_a221oi_1 _6167_ (.B2(net212),
    .C1(_2181_),
    .B1(net38),
    .A1(\line_mapper_1.pointer_addr[9] ),
    .Y(_2375_),
    .A2(net211));
 sg13g2_o21ai_1 _6168_ (.B1(_2375_),
    .Y(_0086_),
    .A1(_2303_),
    .A2(_2374_));
 sg13g2_inv_1 _6169_ (.Y(_2376_),
    .A(\transformer_1.started ));
 sg13g2_a21oi_1 _6170_ (.A1(net37),
    .A2(_2376_),
    .Y(_0087_),
    .B1(net234));
 sg13g2_nand2_1 _6171_ (.Y(_2377_),
    .A(clknet_2_1__leaf_clk),
    .B(net15));
 sg13g2_o21ai_1 _6172_ (.B1(_2377_),
    .Y(clk_buffered),
    .A1(net22),
    .A2(_2201_));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _6175__225 (.L_HI(net243));
 sg13g2_buf_1 _6175_ (.A(net243),
    .X(uio_oe[0]));
 sg13g2_buf_1 _6176_ (.A(net244),
    .X(uio_oe[1]));
 sg13g2_buf_1 _6177_ (.A(net245),
    .X(uio_oe[2]));
 sg13g2_buf_1 _6178_ (.A(net246),
    .X(uio_oe[3]));
 sg13g2_buf_1 _6179_ (.A(net247),
    .X(uio_oe[4]));
 sg13g2_buf_1 _6180_ (.A(net248),
    .X(uio_oe[5]));
 sg13g2_buf_1 _6181_ (.A(net249),
    .X(uio_oe[6]));
 sg13g2_buf_1 _6182_ (.A(net250),
    .X(uio_oe[7]));
 sg13g2_buf_1 _6183_ (.A(net241),
    .X(uio_out[7]));
 sg13g2_buf_1 _6184_ (.A(net242),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \clk_picker.clk_slow$_SDFFE_PN0P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net251),
    .D(_0040_),
    .Q_N(_0030_),
    .Q(\clk_picker.clk_slow ));
 sg13g2_dfrbp_1 \clk_picker.counter[0]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net252),
    .D(_0041_),
    .Q_N(_0039_),
    .Q(\clk_picker.counter[0] ));
 sg13g2_dfrbp_1 \clk_picker.counter[10]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net253),
    .D(_0042_),
    .Q_N(_3093_),
    .Q(\clk_picker.counter[10] ));
 sg13g2_dfrbp_1 \clk_picker.counter[11]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net254),
    .D(_0043_),
    .Q_N(_3092_),
    .Q(\clk_picker.counter[11] ));
 sg13g2_dfrbp_1 \clk_picker.counter[12]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net255),
    .D(_0044_),
    .Q_N(_3091_),
    .Q(\clk_picker.counter[12] ));
 sg13g2_dfrbp_1 \clk_picker.counter[13]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net256),
    .D(_0045_),
    .Q_N(_3090_),
    .Q(\clk_picker.counter[13] ));
 sg13g2_dfrbp_1 \clk_picker.counter[14]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net257),
    .D(_0046_),
    .Q_N(_3089_),
    .Q(\clk_picker.counter[14] ));
 sg13g2_dfrbp_1 \clk_picker.counter[15]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net258),
    .D(_0047_),
    .Q_N(_3088_),
    .Q(\clk_picker.counter[15] ));
 sg13g2_dfrbp_1 \clk_picker.counter[16]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net259),
    .D(_0048_),
    .Q_N(_3087_),
    .Q(\clk_picker.counter[16] ));
 sg13g2_dfrbp_1 \clk_picker.counter[17]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net260),
    .D(_0049_),
    .Q_N(_3086_),
    .Q(\clk_picker.counter[17] ));
 sg13g2_dfrbp_1 \clk_picker.counter[18]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net261),
    .D(_0050_),
    .Q_N(_3085_),
    .Q(\clk_picker.counter[18] ));
 sg13g2_dfrbp_1 \clk_picker.counter[19]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net262),
    .D(_0051_),
    .Q_N(_3084_),
    .Q(\clk_picker.counter[19] ));
 sg13g2_dfrbp_1 \clk_picker.counter[1]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net263),
    .D(_0052_),
    .Q_N(_3083_),
    .Q(\clk_picker.counter[1] ));
 sg13g2_dfrbp_1 \clk_picker.counter[20]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net264),
    .D(_0053_),
    .Q_N(_3082_),
    .Q(\clk_picker.counter[20] ));
 sg13g2_dfrbp_1 \clk_picker.counter[21]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net265),
    .D(_0054_),
    .Q_N(_3081_),
    .Q(\clk_picker.counter[21] ));
 sg13g2_dfrbp_1 \clk_picker.counter[22]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net266),
    .D(_0055_),
    .Q_N(_3080_),
    .Q(\clk_picker.counter[22] ));
 sg13g2_dfrbp_1 \clk_picker.counter[23]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net267),
    .D(_0056_),
    .Q_N(_3079_),
    .Q(\clk_picker.counter[23] ));
 sg13g2_dfrbp_1 \clk_picker.counter[24]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net268),
    .D(_0057_),
    .Q_N(_3078_),
    .Q(\clk_picker.counter[24] ));
 sg13g2_dfrbp_1 \clk_picker.counter[25]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net269),
    .D(_0058_),
    .Q_N(_3077_),
    .Q(\clk_picker.counter[25] ));
 sg13g2_dfrbp_1 \clk_picker.counter[2]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net270),
    .D(_0059_),
    .Q_N(_3076_),
    .Q(\clk_picker.counter[2] ));
 sg13g2_dfrbp_1 \clk_picker.counter[3]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net271),
    .D(_0060_),
    .Q_N(_3075_),
    .Q(\clk_picker.counter[3] ));
 sg13g2_dfrbp_1 \clk_picker.counter[4]$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net272),
    .D(_0061_),
    .Q_N(_3074_),
    .Q(\clk_picker.counter[4] ));
 sg13g2_dfrbp_1 \clk_picker.counter[5]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net273),
    .D(_0062_),
    .Q_N(_3073_),
    .Q(\clk_picker.counter[5] ));
 sg13g2_dfrbp_1 \clk_picker.counter[6]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net274),
    .D(_0063_),
    .Q_N(_3072_),
    .Q(\clk_picker.counter[6] ));
 sg13g2_dfrbp_1 \clk_picker.counter[7]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net275),
    .D(_0064_),
    .Q_N(_3071_),
    .Q(\clk_picker.counter[7] ));
 sg13g2_dfrbp_1 \clk_picker.counter[8]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net276),
    .D(_0065_),
    .Q_N(_3070_),
    .Q(\clk_picker.counter[8] ));
 sg13g2_dfrbp_1 \clk_picker.counter[9]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net277),
    .D(_0066_),
    .Q_N(_3094_),
    .Q(\clk_picker.counter[9] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[0]$_DFF_P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net278),
    .D(_0000_),
    .Q_N(_3095_),
    .Q(\line_mapper_1.pointer_addr[0] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[10]$_DFF_P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net279),
    .D(_0001_),
    .Q_N(_3096_),
    .Q(\line_mapper_1.pointer_addr[10] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[11]$_DFF_P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net280),
    .D(_0002_),
    .Q_N(_3097_),
    .Q(\line_mapper_1.pointer_addr[11] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[12]$_DFF_P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net281),
    .D(_0003_),
    .Q_N(_3098_),
    .Q(\line_mapper_1.pointer_addr[12] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[13]$_DFF_P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net282),
    .D(_0004_),
    .Q_N(_3099_),
    .Q(\line_mapper_1.pointer_addr[13] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[14]$_DFF_P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net283),
    .D(_0005_),
    .Q_N(_3100_),
    .Q(\line_mapper_1.pointer_addr[14] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[15]$_DFF_P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net284),
    .D(_0006_),
    .Q_N(_3101_),
    .Q(\line_mapper_1.pointer_addr[15] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[1]$_DFF_P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net285),
    .D(_0007_),
    .Q_N(_3102_),
    .Q(\line_mapper_1.pointer_addr[1] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[2]$_DFF_P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net286),
    .D(_0008_),
    .Q_N(_3103_),
    .Q(\line_mapper_1.pointer_addr[2] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[3]$_DFF_P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net287),
    .D(_0009_),
    .Q_N(_3104_),
    .Q(\line_mapper_1.pointer_addr[3] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[4]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net288),
    .D(_0010_),
    .Q_N(_3105_),
    .Q(\line_mapper_1.pointer_addr[4] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[5]$_DFF_P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net289),
    .D(_0011_),
    .Q_N(_3106_),
    .Q(\line_mapper_1.pointer_addr[5] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[6]$_DFF_P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net290),
    .D(_0012_),
    .Q_N(_3107_),
    .Q(\line_mapper_1.pointer_addr[6] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[7]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net291),
    .D(_0013_),
    .Q_N(_3108_),
    .Q(\line_mapper_1.pointer_addr[7] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[8]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net292),
    .D(_0014_),
    .Q_N(_3109_),
    .Q(\line_mapper_1.pointer_addr[8] ));
 sg13g2_dfrbp_1 \line_mapper_1.pointer_addr[9]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net293),
    .D(_0015_),
    .Q_N(_3110_),
    .Q(\line_mapper_1.pointer_addr[9] ));
 sg13g2_dfrbp_1 \memory_1.dout[0]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net294),
    .D(_0016_),
    .Q_N(_3111_),
    .Q(net30));
 sg13g2_dfrbp_1 \memory_1.dout[10]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net295),
    .D(_0029_),
    .Q_N(_3112_),
    .Q(net25));
 sg13g2_dfrbp_1 \memory_1.dout[11]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net296),
    .D(_0017_),
    .Q_N(_3113_),
    .Q(net26));
 sg13g2_dfrbp_1 \memory_1.dout[12]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net297),
    .D(_0018_),
    .Q_N(_3114_),
    .Q(net27));
 sg13g2_dfrbp_1 \memory_1.dout[13]$_DFF_P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net298),
    .D(_0019_),
    .Q_N(_3115_),
    .Q(net28));
 sg13g2_dfrbp_1 \memory_1.dout[14]$_DFF_P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net299),
    .D(_0020_),
    .Q_N(_3116_),
    .Q(net29));
 sg13g2_dfrbp_1 \memory_1.dout[1]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net300),
    .D(_0021_),
    .Q_N(_3117_),
    .Q(net31));
 sg13g2_dfrbp_1 \memory_1.dout[2]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net301),
    .D(_0022_),
    .Q_N(_3118_),
    .Q(net32));
 sg13g2_dfrbp_1 \memory_1.dout[3]$_DFF_P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net302),
    .D(_0023_),
    .Q_N(_3119_),
    .Q(net33));
 sg13g2_dfrbp_1 \memory_1.dout[4]$_DFF_P_  (.CLK(clknet_3_2__leaf_clk_buffered),
    .RESET_B(net303),
    .D(_0024_),
    .Q_N(_3120_),
    .Q(net34));
 sg13g2_dfrbp_1 \memory_1.dout[5]$_DFF_P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net304),
    .D(_0025_),
    .Q_N(_3121_),
    .Q(net35));
 sg13g2_dfrbp_1 \memory_1.dout[6]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net305),
    .D(_0026_),
    .Q_N(_3122_),
    .Q(net36));
 sg13g2_dfrbp_1 \memory_1.dout[8]$_DFF_P_  (.CLK(clknet_3_0__leaf_clk_buffered),
    .RESET_B(net306),
    .D(_0027_),
    .Q_N(_3123_),
    .Q(net23));
 sg13g2_dfrbp_1 \memory_1.dout[9]$_DFF_P_  (.CLK(clknet_3_1__leaf_clk_buffered),
    .RESET_B(net307),
    .D(_0028_),
    .Q_N(_3069_),
    .Q(net24));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[0]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net308),
    .D(_0067_),
    .Q_N(_0031_),
    .Q(\chars_remaining[0] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[1]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net309),
    .D(_0068_),
    .Q_N(_3068_),
    .Q(\chars_remaining[1] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[2]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net310),
    .D(_0069_),
    .Q_N(_3067_),
    .Q(\chars_remaining[2] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[3]$_SDFFE_PN0P_  (.CLK(clknet_3_3__leaf_clk_buffered),
    .RESET_B(net311),
    .D(_0070_),
    .Q_N(_3066_),
    .Q(\chars_remaining[3] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[4]$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net312),
    .D(_0071_),
    .Q_N(_3065_),
    .Q(\chars_remaining[4] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[5]$_SDFFE_PN0P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net313),
    .D(_0072_),
    .Q_N(_3064_),
    .Q(\chars_remaining[5] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[6]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net314),
    .D(_0073_),
    .Q_N(_3063_),
    .Q(\chars_remaining[6] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[7]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net315),
    .D(_0074_),
    .Q_N(_3062_),
    .Q(\chars_remaining[7] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[8]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net316),
    .D(_0075_),
    .Q_N(_3061_),
    .Q(\chars_remaining[8] ));
 sg13g2_dfrbp_1 \transformer_1.chars_remaining[9]$_SDFFE_PN0P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net317),
    .D(_0076_),
    .Q_N(_3060_),
    .Q(\chars_remaining[9] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[0]$_SDFFE_PN1P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net318),
    .D(_0077_),
    .Q_N(_0032_),
    .Q(\mem_addr[0] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[1]$_SDFFE_PN1P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net319),
    .D(_0078_),
    .Q_N(_0038_),
    .Q(\mem_addr[1] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[2]$_SDFFE_PN1P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net320),
    .D(_0079_),
    .Q_N(_0037_),
    .Q(\mem_addr[2] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[3]$_SDFFE_PN1P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net321),
    .D(_0080_),
    .Q_N(_0036_),
    .Q(\mem_addr[3] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[4]$_SDFFE_PN1P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net322),
    .D(_0081_),
    .Q_N(_0035_),
    .Q(\mem_addr[4] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[5]$_SDFFE_PN1P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net323),
    .D(_0082_),
    .Q_N(_0034_),
    .Q(\mem_addr[5] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[6]$_SDFFE_PN1P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net324),
    .D(_0083_),
    .Q_N(_0033_),
    .Q(\mem_addr[6] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[7]$_SDFFE_PN1P_  (.CLK(clknet_3_5__leaf_clk_buffered),
    .RESET_B(net325),
    .D(_0084_),
    .Q_N(_3059_),
    .Q(\mem_addr[7] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[8]$_SDFFE_PN1P_  (.CLK(clknet_3_7__leaf_clk_buffered),
    .RESET_B(net326),
    .D(_0085_),
    .Q_N(_3058_),
    .Q(\mem_addr[8] ));
 sg13g2_dfrbp_1 \transformer_1.mem_addr[9]$_SDFFE_PN1P_  (.CLK(clknet_3_4__leaf_clk_buffered),
    .RESET_B(net327),
    .D(_0086_),
    .Q_N(_3057_),
    .Q(\memory_1.mem_addr[9] ));
 sg13g2_dfrbp_1 \transformer_1.started$_SDFFE_PN0P_  (.CLK(clknet_3_6__leaf_clk_buffered),
    .RESET_B(net328),
    .D(_0087_),
    .Q_N(_3056_),
    .Q(\transformer_1.started ));
 sg13g2_dlygate4sd3_1 hold1 (.A(net11),
    .X(net1));
 sg13g2_dlygate4sd3_1 hold2 (.A(net9),
    .X(net2));
 sg13g2_dlygate4sd3_1 hold3 (.A(net13),
    .X(net3));
 sg13g2_dlygate4sd3_1 hold4 (.A(net17),
    .X(net4));
 sg13g2_dlygate4sd3_1 hold5 (.A(net10),
    .X(net5));
 sg13g2_dlygate4sd3_1 hold6 (.A(net12),
    .X(net6));
 sg13g2_dlygate4sd3_1 hold7 (.A(net14),
    .X(net7));
 sg13g2_dlygate4sd3_1 hold8 (.A(net16),
    .X(net8));
 sg13g2_dlygate4sd3_1 hold9 (.A(net18),
    .X(net9));
 sg13g2_dlygate4sd3_1 hold10 (.A(net2),
    .X(net10));
 sg13g2_dlygate4sd3_1 hold11 (.A(net5),
    .X(net11));
 sg13g2_dlygate4sd3_1 hold12 (.A(net1),
    .X(net12));
 sg13g2_dlygate4sd3_1 hold13 (.A(net6),
    .X(net13));
 sg13g2_dlygate4sd3_1 hold14 (.A(net3),
    .X(net14));
 sg13g2_dlygate4sd3_1 hold15 (.A(net7),
    .X(net15));
 sg13g2_dlygate4sd3_1 hold16 (.A(net22),
    .X(net16));
 sg13g2_dlygate4sd3_1 hold17 (.A(net8),
    .X(net17));
 sg13g2_dlygate4sd3_1 hold18 (.A(net4),
    .X(net18));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net19));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net20));
 sg13g2_buf_1 input3 (.A(ui_in[6]),
    .X(net21));
 sg13g2_buf_1 input4 (.A(ui_in[7]),
    .X(net22));
 sg13g2_buf_1 output5 (.A(net23),
    .X(uio_out[0]));
 sg13g2_buf_1 output6 (.A(net24),
    .X(uio_out[1]));
 sg13g2_buf_1 output7 (.A(net25),
    .X(uio_out[2]));
 sg13g2_buf_1 output8 (.A(net26),
    .X(uio_out[3]));
 sg13g2_buf_1 output9 (.A(net27),
    .X(uio_out[4]));
 sg13g2_buf_1 output10 (.A(net28),
    .X(uio_out[5]));
 sg13g2_buf_1 output11 (.A(net29),
    .X(uio_out[6]));
 sg13g2_buf_1 output12 (.A(net30),
    .X(uo_out[0]));
 sg13g2_buf_1 output13 (.A(net31),
    .X(uo_out[1]));
 sg13g2_buf_1 output14 (.A(net32),
    .X(uo_out[2]));
 sg13g2_buf_1 output15 (.A(net33),
    .X(uo_out[3]));
 sg13g2_buf_1 output16 (.A(net34),
    .X(uo_out[4]));
 sg13g2_buf_1 output17 (.A(net35),
    .X(uo_out[5]));
 sg13g2_buf_1 output18 (.A(net36),
    .X(uo_out[6]));
 sg13g2_buf_2 fanout19 (.A(_2305_),
    .X(net37));
 sg13g2_buf_2 fanout20 (.A(_2299_),
    .X(net38));
 sg13g2_buf_2 fanout21 (.A(_0191_),
    .X(net39));
 sg13g2_buf_2 fanout22 (.A(_2845_),
    .X(net40));
 sg13g2_buf_2 fanout23 (.A(_2584_),
    .X(net41));
 sg13g2_buf_2 fanout24 (.A(_2564_),
    .X(net42));
 sg13g2_buf_2 fanout25 (.A(_2527_),
    .X(net43));
 sg13g2_buf_2 fanout26 (.A(_2484_),
    .X(net44));
 sg13g2_buf_2 fanout27 (.A(_2426_),
    .X(net45));
 sg13g2_buf_2 fanout28 (.A(_2424_),
    .X(net46));
 sg13g2_buf_2 fanout29 (.A(_0532_),
    .X(net47));
 sg13g2_buf_2 fanout30 (.A(_0455_),
    .X(net48));
 sg13g2_buf_2 fanout31 (.A(_0297_),
    .X(net49));
 sg13g2_buf_2 fanout32 (.A(_0283_),
    .X(net50));
 sg13g2_buf_2 fanout33 (.A(_0134_),
    .X(net51));
 sg13g2_buf_2 fanout34 (.A(_0114_),
    .X(net52));
 sg13g2_buf_2 fanout35 (.A(_2984_),
    .X(net53));
 sg13g2_buf_2 fanout36 (.A(_2983_),
    .X(net54));
 sg13g2_buf_2 fanout37 (.A(_2947_),
    .X(net55));
 sg13g2_buf_2 fanout38 (.A(_2871_),
    .X(net56));
 sg13g2_buf_2 fanout39 (.A(_2805_),
    .X(net57));
 sg13g2_buf_2 fanout40 (.A(_2771_),
    .X(net58));
 sg13g2_buf_2 fanout41 (.A(_2714_),
    .X(net59));
 sg13g2_buf_2 fanout42 (.A(_2701_),
    .X(net60));
 sg13g2_buf_2 fanout43 (.A(_2700_),
    .X(net61));
 sg13g2_buf_2 fanout44 (.A(_2624_),
    .X(net62));
 sg13g2_buf_2 fanout45 (.A(_2595_),
    .X(net63));
 sg13g2_buf_2 fanout46 (.A(_2555_),
    .X(net64));
 sg13g2_buf_2 fanout47 (.A(_2540_),
    .X(net65));
 sg13g2_buf_2 fanout48 (.A(_2537_),
    .X(net66));
 sg13g2_buf_2 fanout49 (.A(_2529_),
    .X(net67));
 sg13g2_buf_2 fanout50 (.A(_2526_),
    .X(net68));
 sg13g2_buf_2 fanout51 (.A(_2523_),
    .X(net69));
 sg13g2_buf_2 fanout52 (.A(_2521_),
    .X(net70));
 sg13g2_buf_2 fanout53 (.A(_2486_),
    .X(net71));
 sg13g2_buf_2 fanout54 (.A(_2462_),
    .X(net72));
 sg13g2_buf_2 fanout55 (.A(_2441_),
    .X(net73));
 sg13g2_buf_2 fanout56 (.A(_2425_),
    .X(net74));
 sg13g2_buf_2 fanout57 (.A(_2423_),
    .X(net75));
 sg13g2_buf_2 fanout58 (.A(_2378_),
    .X(net76));
 sg13g2_buf_2 fanout59 (.A(_2259_),
    .X(net77));
 sg13g2_buf_2 fanout60 (.A(_1621_),
    .X(net78));
 sg13g2_buf_2 fanout61 (.A(_1523_),
    .X(net79));
 sg13g2_buf_2 fanout62 (.A(_1468_),
    .X(net80));
 sg13g2_buf_2 fanout63 (.A(_1381_),
    .X(net81));
 sg13g2_buf_2 fanout64 (.A(_1064_),
    .X(net82));
 sg13g2_buf_2 fanout65 (.A(_1020_),
    .X(net83));
 sg13g2_buf_2 fanout66 (.A(_0482_),
    .X(net84));
 sg13g2_buf_2 fanout67 (.A(_0381_),
    .X(net85));
 sg13g2_buf_2 fanout68 (.A(_0351_),
    .X(net86));
 sg13g2_buf_2 fanout69 (.A(_0308_),
    .X(net87));
 sg13g2_buf_2 fanout70 (.A(_0304_),
    .X(net88));
 sg13g2_buf_2 fanout71 (.A(_0197_),
    .X(net89));
 sg13g2_buf_2 fanout72 (.A(_0118_),
    .X(net90));
 sg13g2_buf_2 fanout73 (.A(_2971_),
    .X(net91));
 sg13g2_buf_2 fanout74 (.A(_2967_),
    .X(net92));
 sg13g2_buf_2 fanout75 (.A(_2946_),
    .X(net93));
 sg13g2_buf_2 fanout76 (.A(_2904_),
    .X(net94));
 sg13g2_buf_2 fanout77 (.A(_2882_),
    .X(net95));
 sg13g2_buf_2 fanout78 (.A(_2863_),
    .X(net96));
 sg13g2_buf_2 fanout79 (.A(_2860_),
    .X(net97));
 sg13g2_buf_2 fanout80 (.A(_2839_),
    .X(net98));
 sg13g2_buf_2 fanout81 (.A(_2819_),
    .X(net99));
 sg13g2_buf_2 fanout82 (.A(_2808_),
    .X(net100));
 sg13g2_buf_2 fanout83 (.A(_2769_),
    .X(net101));
 sg13g2_buf_2 fanout84 (.A(_2659_),
    .X(net102));
 sg13g2_buf_2 fanout85 (.A(_2648_),
    .X(net103));
 sg13g2_buf_2 fanout86 (.A(_2637_),
    .X(net104));
 sg13g2_buf_2 fanout87 (.A(_2634_),
    .X(net105));
 sg13g2_buf_2 fanout88 (.A(_2606_),
    .X(net106));
 sg13g2_buf_2 fanout89 (.A(_2597_),
    .X(net107));
 sg13g2_buf_2 fanout90 (.A(_2568_),
    .X(net108));
 sg13g2_buf_2 fanout91 (.A(_2566_),
    .X(net109));
 sg13g2_buf_2 fanout92 (.A(_2551_),
    .X(net110));
 sg13g2_buf_2 fanout93 (.A(_2531_),
    .X(net111));
 sg13g2_buf_2 fanout94 (.A(_2479_),
    .X(net112));
 sg13g2_buf_2 fanout95 (.A(_2472_),
    .X(net113));
 sg13g2_buf_2 fanout96 (.A(_2463_),
    .X(net114));
 sg13g2_buf_2 fanout97 (.A(_2459_),
    .X(net115));
 sg13g2_buf_2 fanout98 (.A(_2422_),
    .X(net116));
 sg13g2_buf_2 fanout99 (.A(_2401_),
    .X(net117));
 sg13g2_buf_2 fanout100 (.A(_2391_),
    .X(net118));
 sg13g2_buf_2 fanout101 (.A(_2370_),
    .X(net119));
 sg13g2_buf_2 fanout102 (.A(_2280_),
    .X(net120));
 sg13g2_buf_2 fanout103 (.A(_2225_),
    .X(net121));
 sg13g2_buf_2 fanout104 (.A(_2184_),
    .X(net122));
 sg13g2_buf_4 fanout105 (.X(net123),
    .A(_2066_));
 sg13g2_buf_2 fanout106 (.A(_2056_),
    .X(net124));
 sg13g2_buf_2 fanout107 (.A(_1991_),
    .X(net125));
 sg13g2_buf_2 fanout108 (.A(_1850_),
    .X(net126));
 sg13g2_buf_2 fanout109 (.A(_1796_),
    .X(net127));
 sg13g2_buf_2 fanout110 (.A(_1457_),
    .X(net128));
 sg13g2_buf_2 fanout111 (.A(_1348_),
    .X(net129));
 sg13g2_buf_2 fanout112 (.A(_1304_),
    .X(net130));
 sg13g2_buf_2 fanout113 (.A(_1228_),
    .X(net131));
 sg13g2_buf_2 fanout114 (.A(_1108_),
    .X(net132));
 sg13g2_buf_2 fanout115 (.A(_0896_),
    .X(net133));
 sg13g2_buf_2 fanout116 (.A(_0260_),
    .X(net134));
 sg13g2_buf_2 fanout117 (.A(_0194_),
    .X(net135));
 sg13g2_buf_2 fanout118 (.A(_0141_),
    .X(net136));
 sg13g2_buf_2 fanout119 (.A(_0136_),
    .X(net137));
 sg13g2_buf_2 fanout120 (.A(_3042_),
    .X(net138));
 sg13g2_buf_2 fanout121 (.A(_2999_),
    .X(net139));
 sg13g2_buf_2 fanout122 (.A(_2890_),
    .X(net140));
 sg13g2_buf_2 fanout123 (.A(_2840_),
    .X(net141));
 sg13g2_buf_2 fanout124 (.A(_2793_),
    .X(net142));
 sg13g2_buf_2 fanout125 (.A(_2749_),
    .X(net143));
 sg13g2_buf_2 fanout126 (.A(_2727_),
    .X(net144));
 sg13g2_buf_2 fanout127 (.A(_2711_),
    .X(net145));
 sg13g2_buf_2 fanout128 (.A(_2705_),
    .X(net146));
 sg13g2_buf_2 fanout129 (.A(_2689_),
    .X(net147));
 sg13g2_buf_2 fanout130 (.A(_2665_),
    .X(net148));
 sg13g2_buf_2 fanout131 (.A(_2658_),
    .X(net149));
 sg13g2_buf_2 fanout132 (.A(_2629_),
    .X(net150));
 sg13g2_buf_2 fanout133 (.A(_2594_),
    .X(net151));
 sg13g2_buf_2 fanout134 (.A(_2575_),
    .X(net152));
 sg13g2_buf_2 fanout135 (.A(_2560_),
    .X(net153));
 sg13g2_buf_2 fanout136 (.A(_2553_),
    .X(net154));
 sg13g2_buf_2 fanout137 (.A(_2550_),
    .X(net155));
 sg13g2_buf_2 fanout138 (.A(_2548_),
    .X(net156));
 sg13g2_buf_2 fanout139 (.A(_2501_),
    .X(net157));
 sg13g2_buf_2 fanout140 (.A(_2487_),
    .X(net158));
 sg13g2_buf_2 fanout141 (.A(_2478_),
    .X(net159));
 sg13g2_buf_2 fanout142 (.A(_2474_),
    .X(net160));
 sg13g2_buf_2 fanout143 (.A(_2469_),
    .X(net161));
 sg13g2_buf_2 fanout144 (.A(_2450_),
    .X(net162));
 sg13g2_buf_2 fanout145 (.A(_2431_),
    .X(net163));
 sg13g2_buf_2 fanout146 (.A(_2421_),
    .X(net164));
 sg13g2_buf_2 fanout147 (.A(_2418_),
    .X(net165));
 sg13g2_buf_2 fanout148 (.A(_2414_),
    .X(net166));
 sg13g2_buf_2 fanout149 (.A(_2406_),
    .X(net167));
 sg13g2_buf_2 fanout150 (.A(_2395_),
    .X(net168));
 sg13g2_buf_2 fanout151 (.A(_2390_),
    .X(net169));
 sg13g2_buf_2 fanout152 (.A(_2379_),
    .X(net170));
 sg13g2_buf_2 fanout153 (.A(_2361_),
    .X(net171));
 sg13g2_buf_2 fanout154 (.A(_2175_),
    .X(net172));
 sg13g2_buf_4 fanout155 (.X(net173),
    .A(_2024_));
 sg13g2_buf_2 fanout156 (.A(_1981_),
    .X(net174));
 sg13g2_buf_2 fanout157 (.A(_1719_),
    .X(net175));
 sg13g2_buf_4 fanout158 (.X(net176),
    .A(_1708_));
 sg13g2_buf_2 fanout159 (.A(_1654_),
    .X(net177));
 sg13g2_buf_2 fanout160 (.A(_1599_),
    .X(net178));
 sg13g2_buf_2 fanout161 (.A(_1173_),
    .X(net179));
 sg13g2_buf_4 fanout162 (.X(net180),
    .A(_1097_));
 sg13g2_buf_2 fanout163 (.A(_2301_),
    .X(net181));
 sg13g2_buf_2 fanout164 (.A(_0713_),
    .X(net182));
 sg13g2_buf_2 fanout165 (.A(_0556_),
    .X(net183));
 sg13g2_buf_2 fanout166 (.A(_0272_),
    .X(net184));
 sg13g2_buf_2 fanout167 (.A(_0140_),
    .X(net185));
 sg13g2_buf_2 fanout168 (.A(_3044_),
    .X(net186));
 sg13g2_buf_2 fanout169 (.A(_3041_),
    .X(net187));
 sg13g2_buf_2 fanout170 (.A(_3010_),
    .X(net188));
 sg13g2_buf_2 fanout171 (.A(_2998_),
    .X(net189));
 sg13g2_buf_2 fanout172 (.A(_2751_),
    .X(net190));
 sg13g2_buf_2 fanout173 (.A(_2673_),
    .X(net191));
 sg13g2_buf_2 fanout174 (.A(_2628_),
    .X(net192));
 sg13g2_buf_2 fanout175 (.A(_2547_),
    .X(net193));
 sg13g2_buf_2 fanout176 (.A(_2517_),
    .X(net194));
 sg13g2_buf_2 fanout177 (.A(_2500_),
    .X(net195));
 sg13g2_buf_2 fanout178 (.A(_2492_),
    .X(net196));
 sg13g2_buf_2 fanout179 (.A(_2430_),
    .X(net197));
 sg13g2_buf_2 fanout180 (.A(_2420_),
    .X(net198));
 sg13g2_buf_2 fanout181 (.A(_2413_),
    .X(net199));
 sg13g2_buf_2 fanout182 (.A(_2386_),
    .X(net200));
 sg13g2_buf_2 fanout183 (.A(_2383_),
    .X(net201));
 sg13g2_buf_2 fanout184 (.A(_2165_),
    .X(net202));
 sg13g2_buf_2 fanout185 (.A(_1970_),
    .X(net203));
 sg13g2_buf_2 fanout186 (.A(_1817_),
    .X(net204));
 sg13g2_buf_4 fanout187 (.X(net205),
    .A(_1697_));
 sg13g2_buf_2 fanout188 (.A(_1534_),
    .X(net206));
 sg13g2_buf_4 fanout189 (.X(net207),
    .A(_1086_));
 sg13g2_buf_4 fanout190 (.X(net208),
    .A(_1031_));
 sg13g2_buf_2 fanout191 (.A(_0998_),
    .X(net209));
 sg13g2_buf_2 fanout192 (.A(_0966_),
    .X(net210));
 sg13g2_buf_2 fanout193 (.A(_2284_),
    .X(net211));
 sg13g2_buf_2 fanout194 (.A(_0495_),
    .X(net212));
 sg13g2_buf_2 fanout195 (.A(_2920_),
    .X(net213));
 sg13g2_buf_2 fanout196 (.A(_2779_),
    .X(net214));
 sg13g2_buf_2 fanout197 (.A(_2630_),
    .X(net215));
 sg13g2_buf_2 fanout198 (.A(_2592_),
    .X(net216));
 sg13g2_buf_2 fanout199 (.A(_2546_),
    .X(net217));
 sg13g2_buf_2 fanout200 (.A(_2516_),
    .X(net218));
 sg13g2_buf_2 fanout201 (.A(_2491_),
    .X(net219));
 sg13g2_buf_4 fanout202 (.X(net220),
    .A(_2398_));
 sg13g2_buf_2 fanout203 (.A(_2388_),
    .X(net221));
 sg13g2_buf_4 fanout204 (.X(net222),
    .A(_1239_));
 sg13g2_buf_2 fanout205 (.A(_0987_),
    .X(net223));
 sg13g2_buf_2 fanout206 (.A(_0955_),
    .X(net224));
 sg13g2_buf_4 fanout207 (.X(net225),
    .A(_0878_));
 sg13g2_buf_2 fanout208 (.A(_3002_),
    .X(net226));
 sg13g2_buf_2 fanout209 (.A(_1140_),
    .X(net227));
 sg13g2_buf_2 fanout210 (.A(_0736_),
    .X(net228));
 sg13g2_buf_2 fanout211 (.A(_0725_),
    .X(net229));
 sg13g2_buf_2 fanout212 (.A(_2233_),
    .X(net230));
 sg13g2_buf_2 fanout213 (.A(_2209_),
    .X(net231));
 sg13g2_buf_2 fanout214 (.A(_2078_),
    .X(net232));
 sg13g2_buf_2 fanout215 (.A(_2055_),
    .X(net233));
 sg13g2_buf_2 fanout216 (.A(_2182_),
    .X(net234));
 sg13g2_buf_2 fanout217 (.A(_2028_),
    .X(net235));
 sg13g2_buf_2 fanout218 (.A(_2018_),
    .X(net236));
 sg13g2_buf_2 fanout219 (.A(_1995_),
    .X(net237));
 sg13g2_buf_2 fanout220 (.A(_2181_),
    .X(net238));
 sg13g2_buf_2 fanout221 (.A(_2001_),
    .X(net239));
 sg13g2_buf_2 fanout222 (.A(_1996_),
    .X(net240));
 sg13g2_tielo _6183__223 (.L_LO(net241));
 sg13g2_tielo _6184__224 (.L_LO(net242));
 sg13g2_tiehi _6176__226 (.L_HI(net244));
 sg13g2_tiehi _6177__227 (.L_HI(net245));
 sg13g2_tiehi _6178__228 (.L_HI(net246));
 sg13g2_tiehi _6179__229 (.L_HI(net247));
 sg13g2_tiehi _6180__230 (.L_HI(net248));
 sg13g2_tiehi _6181__231 (.L_HI(net249));
 sg13g2_tiehi _6182__232 (.L_HI(net250));
 sg13g2_tiehi \clk_picker.clk_slow$_SDFFE_PN0P__233  (.L_HI(net251));
 sg13g2_tiehi \clk_picker.counter[0]$_SDFF_PN0__234  (.L_HI(net252));
 sg13g2_tiehi \clk_picker.counter[10]$_SDFF_PN0__235  (.L_HI(net253));
 sg13g2_tiehi \clk_picker.counter[11]$_SDFF_PN0__236  (.L_HI(net254));
 sg13g2_tiehi \clk_picker.counter[12]$_SDFF_PN0__237  (.L_HI(net255));
 sg13g2_tiehi \clk_picker.counter[13]$_SDFF_PN0__238  (.L_HI(net256));
 sg13g2_tiehi \clk_picker.counter[14]$_SDFF_PN0__239  (.L_HI(net257));
 sg13g2_tiehi \clk_picker.counter[15]$_SDFF_PN0__240  (.L_HI(net258));
 sg13g2_tiehi \clk_picker.counter[16]$_SDFF_PN0__241  (.L_HI(net259));
 sg13g2_tiehi \clk_picker.counter[17]$_SDFF_PN0__242  (.L_HI(net260));
 sg13g2_tiehi \clk_picker.counter[18]$_SDFF_PN0__243  (.L_HI(net261));
 sg13g2_tiehi \clk_picker.counter[19]$_SDFF_PN0__244  (.L_HI(net262));
 sg13g2_tiehi \clk_picker.counter[1]$_SDFF_PN0__245  (.L_HI(net263));
 sg13g2_tiehi \clk_picker.counter[20]$_SDFF_PN0__246  (.L_HI(net264));
 sg13g2_tiehi \clk_picker.counter[21]$_SDFF_PN0__247  (.L_HI(net265));
 sg13g2_tiehi \clk_picker.counter[22]$_SDFF_PN0__248  (.L_HI(net266));
 sg13g2_tiehi \clk_picker.counter[23]$_SDFF_PN0__249  (.L_HI(net267));
 sg13g2_tiehi \clk_picker.counter[24]$_SDFF_PN0__250  (.L_HI(net268));
 sg13g2_tiehi \clk_picker.counter[25]$_SDFF_PN0__251  (.L_HI(net269));
 sg13g2_tiehi \clk_picker.counter[2]$_SDFF_PN0__252  (.L_HI(net270));
 sg13g2_tiehi \clk_picker.counter[3]$_SDFF_PN0__253  (.L_HI(net271));
 sg13g2_tiehi \clk_picker.counter[4]$_SDFF_PN0__254  (.L_HI(net272));
 sg13g2_tiehi \clk_picker.counter[5]$_SDFF_PN0__255  (.L_HI(net273));
 sg13g2_tiehi \clk_picker.counter[6]$_SDFF_PN0__256  (.L_HI(net274));
 sg13g2_tiehi \clk_picker.counter[7]$_SDFF_PN0__257  (.L_HI(net275));
 sg13g2_tiehi \clk_picker.counter[8]$_SDFF_PN0__258  (.L_HI(net276));
 sg13g2_tiehi \clk_picker.counter[9]$_SDFF_PN0__259  (.L_HI(net277));
 sg13g2_tiehi \line_mapper_1.pointer_addr[0]$_DFF_P__260  (.L_HI(net278));
 sg13g2_tiehi \line_mapper_1.pointer_addr[10]$_DFF_P__261  (.L_HI(net279));
 sg13g2_tiehi \line_mapper_1.pointer_addr[11]$_DFF_P__262  (.L_HI(net280));
 sg13g2_tiehi \line_mapper_1.pointer_addr[12]$_DFF_P__263  (.L_HI(net281));
 sg13g2_tiehi \line_mapper_1.pointer_addr[13]$_DFF_P__264  (.L_HI(net282));
 sg13g2_tiehi \line_mapper_1.pointer_addr[14]$_DFF_P__265  (.L_HI(net283));
 sg13g2_tiehi \line_mapper_1.pointer_addr[15]$_DFF_P__266  (.L_HI(net284));
 sg13g2_tiehi \line_mapper_1.pointer_addr[1]$_DFF_P__267  (.L_HI(net285));
 sg13g2_tiehi \line_mapper_1.pointer_addr[2]$_DFF_P__268  (.L_HI(net286));
 sg13g2_tiehi \line_mapper_1.pointer_addr[3]$_DFF_P__269  (.L_HI(net287));
 sg13g2_tiehi \line_mapper_1.pointer_addr[4]$_DFF_P__270  (.L_HI(net288));
 sg13g2_tiehi \line_mapper_1.pointer_addr[5]$_DFF_P__271  (.L_HI(net289));
 sg13g2_tiehi \line_mapper_1.pointer_addr[6]$_DFF_P__272  (.L_HI(net290));
 sg13g2_tiehi \line_mapper_1.pointer_addr[7]$_DFF_P__273  (.L_HI(net291));
 sg13g2_tiehi \line_mapper_1.pointer_addr[8]$_DFF_P__274  (.L_HI(net292));
 sg13g2_tiehi \line_mapper_1.pointer_addr[9]$_DFF_P__275  (.L_HI(net293));
 sg13g2_tiehi \memory_1.dout[0]$_DFF_P__276  (.L_HI(net294));
 sg13g2_tiehi \memory_1.dout[10]$_DFF_P__277  (.L_HI(net295));
 sg13g2_tiehi \memory_1.dout[11]$_DFF_P__278  (.L_HI(net296));
 sg13g2_tiehi \memory_1.dout[12]$_DFF_P__279  (.L_HI(net297));
 sg13g2_tiehi \memory_1.dout[13]$_DFF_P__280  (.L_HI(net298));
 sg13g2_tiehi \memory_1.dout[14]$_DFF_P__281  (.L_HI(net299));
 sg13g2_tiehi \memory_1.dout[1]$_DFF_P__282  (.L_HI(net300));
 sg13g2_tiehi \memory_1.dout[2]$_DFF_P__283  (.L_HI(net301));
 sg13g2_tiehi \memory_1.dout[3]$_DFF_P__284  (.L_HI(net302));
 sg13g2_tiehi \memory_1.dout[4]$_DFF_P__285  (.L_HI(net303));
 sg13g2_tiehi \memory_1.dout[5]$_DFF_P__286  (.L_HI(net304));
 sg13g2_tiehi \memory_1.dout[6]$_DFF_P__287  (.L_HI(net305));
 sg13g2_tiehi \memory_1.dout[8]$_DFF_P__288  (.L_HI(net306));
 sg13g2_tiehi \memory_1.dout[9]$_DFF_P__289  (.L_HI(net307));
 sg13g2_tiehi \transformer_1.chars_remaining[0]$_SDFFE_PN0P__290  (.L_HI(net308));
 sg13g2_tiehi \transformer_1.chars_remaining[1]$_SDFFE_PN0P__291  (.L_HI(net309));
 sg13g2_tiehi \transformer_1.chars_remaining[2]$_SDFFE_PN0P__292  (.L_HI(net310));
 sg13g2_tiehi \transformer_1.chars_remaining[3]$_SDFFE_PN0P__293  (.L_HI(net311));
 sg13g2_tiehi \transformer_1.chars_remaining[4]$_SDFFE_PN0P__294  (.L_HI(net312));
 sg13g2_tiehi \transformer_1.chars_remaining[5]$_SDFFE_PN0P__295  (.L_HI(net313));
 sg13g2_tiehi \transformer_1.chars_remaining[6]$_SDFFE_PN0P__296  (.L_HI(net314));
 sg13g2_tiehi \transformer_1.chars_remaining[7]$_SDFFE_PN0P__297  (.L_HI(net315));
 sg13g2_tiehi \transformer_1.chars_remaining[8]$_SDFFE_PN0P__298  (.L_HI(net316));
 sg13g2_tiehi \transformer_1.chars_remaining[9]$_SDFFE_PN0P__299  (.L_HI(net317));
 sg13g2_tiehi \transformer_1.mem_addr[0]$_SDFFE_PN1P__300  (.L_HI(net318));
 sg13g2_tiehi \transformer_1.mem_addr[1]$_SDFFE_PN1P__301  (.L_HI(net319));
 sg13g2_tiehi \transformer_1.mem_addr[2]$_SDFFE_PN1P__302  (.L_HI(net320));
 sg13g2_tiehi \transformer_1.mem_addr[3]$_SDFFE_PN1P__303  (.L_HI(net321));
 sg13g2_tiehi \transformer_1.mem_addr[4]$_SDFFE_PN1P__304  (.L_HI(net322));
 sg13g2_tiehi \transformer_1.mem_addr[5]$_SDFFE_PN1P__305  (.L_HI(net323));
 sg13g2_tiehi \transformer_1.mem_addr[6]$_SDFFE_PN1P__306  (.L_HI(net324));
 sg13g2_tiehi \transformer_1.mem_addr[7]$_SDFFE_PN1P__307  (.L_HI(net325));
 sg13g2_tiehi \transformer_1.mem_addr[8]$_SDFFE_PN1P__308  (.L_HI(net326));
 sg13g2_tiehi \transformer_1.mem_addr[9]$_SDFFE_PN1P__309  (.L_HI(net327));
 sg13g2_tiehi \transformer_1.started$_SDFFE_PN0P__310  (.L_HI(net328));
 sg13g2_buf_2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_2 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_2 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_2 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_2_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_2_2__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_2_3__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk_buffered (.A(clk_buffered),
    .X(clknet_0_clk_buffered));
 sg13g2_buf_2 clkbuf_3_0__f_clk_buffered (.A(clknet_0_clk_buffered),
    .X(clknet_3_0__leaf_clk_buffered));
 sg13g2_buf_2 clkbuf_3_1__f_clk_buffered (.A(clknet_0_clk_buffered),
    .X(clknet_3_1__leaf_clk_buffered));
 sg13g2_buf_2 clkbuf_3_2__f_clk_buffered (.A(clknet_0_clk_buffered),
    .X(clknet_3_2__leaf_clk_buffered));
 sg13g2_buf_2 clkbuf_3_3__f_clk_buffered (.A(clknet_0_clk_buffered),
    .X(clknet_3_3__leaf_clk_buffered));
 sg13g2_buf_2 clkbuf_3_4__f_clk_buffered (.A(clknet_0_clk_buffered),
    .X(clknet_3_4__leaf_clk_buffered));
 sg13g2_buf_2 clkbuf_3_5__f_clk_buffered (.A(clknet_0_clk_buffered),
    .X(clknet_3_5__leaf_clk_buffered));
 sg13g2_buf_2 clkbuf_3_6__f_clk_buffered (.A(clknet_0_clk_buffered),
    .X(clknet_3_6__leaf_clk_buffered));
 sg13g2_buf_2 clkbuf_3_7__f_clk_buffered (.A(clknet_0_clk_buffered),
    .X(clknet_3_7__leaf_clk_buffered));
 sg13g2_inv_1 clkload3 (.A(clknet_3_1__leaf_clk_buffered));
 sg13g2_inv_1 clkload4 (.A(clknet_3_3__leaf_clk_buffered));
 sg13g2_inv_1 clkload5 (.A(clknet_3_5__leaf_clk_buffered));
 sg13g2_inv_1 clkload6 (.A(clknet_3_6__leaf_clk_buffered));
 sg13g2_inv_1 clkload7 (.A(clknet_3_7__leaf_clk_buffered));
 sg13g2_antennanp ANTENNA_1 (.A(_0023_));
 sg13g2_antennanp ANTENNA_2 (.A(_0077_));
 sg13g2_antennanp ANTENNA_3 (.A(_0077_));
 sg13g2_antennanp ANTENNA_4 (.A(_0079_));
 sg13g2_antennanp ANTENNA_5 (.A(_0079_));
 sg13g2_antennanp ANTENNA_6 (.A(_0080_));
 sg13g2_antennanp ANTENNA_7 (.A(_0080_));
 sg13g2_antennanp ANTENNA_8 (.A(_0081_));
 sg13g2_antennanp ANTENNA_9 (.A(_0081_));
 sg13g2_antennanp ANTENNA_10 (.A(_0083_));
 sg13g2_antennanp ANTENNA_11 (.A(_0083_));
 sg13g2_antennanp ANTENNA_12 (.A(_0084_));
 sg13g2_antennanp ANTENNA_13 (.A(_0084_));
 sg13g2_antennanp ANTENNA_14 (.A(_0283_));
 sg13g2_antennanp ANTENNA_15 (.A(_0283_));
 sg13g2_antennanp ANTENNA_16 (.A(_0283_));
 sg13g2_antennanp ANTENNA_17 (.A(_2409_));
 sg13g2_antennanp ANTENNA_18 (.A(_2798_));
 sg13g2_antennanp ANTENNA_19 (.A(\mem_addr[1] ));
 sg13g2_antennanp ANTENNA_20 (.A(_0023_));
 sg13g2_antennanp ANTENNA_21 (.A(_0079_));
 sg13g2_antennanp ANTENNA_22 (.A(_0079_));
 sg13g2_antennanp ANTENNA_23 (.A(_0080_));
 sg13g2_antennanp ANTENNA_24 (.A(_0080_));
 sg13g2_antennanp ANTENNA_25 (.A(_0084_));
 sg13g2_antennanp ANTENNA_26 (.A(_0084_));
 sg13g2_antennanp ANTENNA_27 (.A(_0283_));
 sg13g2_antennanp ANTENNA_28 (.A(_0283_));
 sg13g2_antennanp ANTENNA_29 (.A(_0283_));
 sg13g2_antennanp ANTENNA_30 (.A(_2409_));
 sg13g2_antennanp ANTENNA_31 (.A(_2798_));
 sg13g2_antennanp ANTENNA_32 (.A(\mem_addr[1] ));
 sg13g2_antennanp ANTENNA_33 (.A(_0023_));
 sg13g2_antennanp ANTENNA_34 (.A(_0080_));
 sg13g2_antennanp ANTENNA_35 (.A(_0080_));
 sg13g2_antennanp ANTENNA_36 (.A(_0084_));
 sg13g2_antennanp ANTENNA_37 (.A(_0084_));
 sg13g2_antennanp ANTENNA_38 (.A(_0283_));
 sg13g2_antennanp ANTENNA_39 (.A(_0283_));
 sg13g2_antennanp ANTENNA_40 (.A(_0283_));
 sg13g2_antennanp ANTENNA_41 (.A(_2409_));
 sg13g2_antennanp ANTENNA_42 (.A(_2798_));
 sg13g2_antennanp ANTENNA_43 (.A(\mem_addr[1] ));
 sg13g2_antennanp ANTENNA_44 (.A(_0023_));
 sg13g2_antennanp ANTENNA_45 (.A(_0084_));
 sg13g2_antennanp ANTENNA_46 (.A(_0084_));
 sg13g2_antennanp ANTENNA_47 (.A(_0283_));
 sg13g2_antennanp ANTENNA_48 (.A(_0283_));
 sg13g2_antennanp ANTENNA_49 (.A(_0283_));
 sg13g2_antennanp ANTENNA_50 (.A(_2409_));
 sg13g2_antennanp ANTENNA_51 (.A(_2798_));
 sg13g2_antennanp ANTENNA_52 (.A(\mem_addr[1] ));
 sg13g2_antennanp ANTENNA_53 (.A(_0023_));
 sg13g2_antennanp ANTENNA_54 (.A(_0084_));
 sg13g2_antennanp ANTENNA_55 (.A(_0084_));
 sg13g2_antennanp ANTENNA_56 (.A(_0283_));
 sg13g2_antennanp ANTENNA_57 (.A(_0283_));
 sg13g2_antennanp ANTENNA_58 (.A(_0283_));
 sg13g2_antennanp ANTENNA_59 (.A(_2409_));
 sg13g2_antennanp ANTENNA_60 (.A(_2798_));
 sg13g2_antennanp ANTENNA_61 (.A(\mem_addr[1] ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_fill_2 FILLER_0_875 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_fill_2 FILLER_1_875 ();
 sg13g2_fill_1 FILLER_1_877 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_decap_8 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_2_868 ();
 sg13g2_fill_2 FILLER_2_875 ();
 sg13g2_fill_1 FILLER_2_877 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_fill_2 FILLER_3_875 ();
 sg13g2_fill_1 FILLER_3_877 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_fill_2 FILLER_4_875 ();
 sg13g2_fill_1 FILLER_4_877 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_decap_8 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_5_868 ();
 sg13g2_fill_2 FILLER_5_875 ();
 sg13g2_fill_1 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_decap_8 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_6_868 ();
 sg13g2_fill_2 FILLER_6_875 ();
 sg13g2_fill_1 FILLER_6_877 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_fill_2 FILLER_7_875 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_fill_2 FILLER_8_875 ();
 sg13g2_fill_1 FILLER_8_877 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_fill_2 FILLER_9_875 ();
 sg13g2_fill_1 FILLER_9_877 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_fill_2 FILLER_10_392 ();
 sg13g2_fill_1 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_decap_8 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_10_436 ();
 sg13g2_decap_8 FILLER_10_443 ();
 sg13g2_decap_8 FILLER_10_450 ();
 sg13g2_decap_8 FILLER_10_457 ();
 sg13g2_decap_8 FILLER_10_464 ();
 sg13g2_decap_8 FILLER_10_471 ();
 sg13g2_decap_8 FILLER_10_478 ();
 sg13g2_decap_8 FILLER_10_485 ();
 sg13g2_decap_8 FILLER_10_492 ();
 sg13g2_decap_8 FILLER_10_499 ();
 sg13g2_decap_8 FILLER_10_506 ();
 sg13g2_decap_8 FILLER_10_513 ();
 sg13g2_decap_8 FILLER_10_520 ();
 sg13g2_decap_8 FILLER_10_527 ();
 sg13g2_decap_8 FILLER_10_534 ();
 sg13g2_decap_8 FILLER_10_541 ();
 sg13g2_decap_8 FILLER_10_548 ();
 sg13g2_decap_8 FILLER_10_555 ();
 sg13g2_decap_8 FILLER_10_562 ();
 sg13g2_decap_8 FILLER_10_569 ();
 sg13g2_decap_8 FILLER_10_576 ();
 sg13g2_decap_8 FILLER_10_583 ();
 sg13g2_decap_8 FILLER_10_590 ();
 sg13g2_decap_8 FILLER_10_597 ();
 sg13g2_decap_8 FILLER_10_604 ();
 sg13g2_decap_8 FILLER_10_611 ();
 sg13g2_decap_8 FILLER_10_618 ();
 sg13g2_decap_8 FILLER_10_625 ();
 sg13g2_decap_8 FILLER_10_632 ();
 sg13g2_decap_8 FILLER_10_639 ();
 sg13g2_decap_8 FILLER_10_646 ();
 sg13g2_decap_8 FILLER_10_653 ();
 sg13g2_decap_8 FILLER_10_660 ();
 sg13g2_decap_8 FILLER_10_667 ();
 sg13g2_decap_8 FILLER_10_674 ();
 sg13g2_decap_8 FILLER_10_681 ();
 sg13g2_decap_8 FILLER_10_688 ();
 sg13g2_decap_8 FILLER_10_695 ();
 sg13g2_decap_8 FILLER_10_702 ();
 sg13g2_decap_8 FILLER_10_709 ();
 sg13g2_decap_8 FILLER_10_716 ();
 sg13g2_decap_8 FILLER_10_723 ();
 sg13g2_decap_8 FILLER_10_730 ();
 sg13g2_decap_8 FILLER_10_737 ();
 sg13g2_decap_8 FILLER_10_744 ();
 sg13g2_decap_8 FILLER_10_751 ();
 sg13g2_decap_8 FILLER_10_758 ();
 sg13g2_decap_8 FILLER_10_765 ();
 sg13g2_decap_8 FILLER_10_772 ();
 sg13g2_decap_8 FILLER_10_779 ();
 sg13g2_decap_8 FILLER_10_786 ();
 sg13g2_decap_8 FILLER_10_793 ();
 sg13g2_decap_8 FILLER_10_800 ();
 sg13g2_decap_8 FILLER_10_807 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_8 FILLER_10_828 ();
 sg13g2_decap_8 FILLER_10_835 ();
 sg13g2_decap_8 FILLER_10_842 ();
 sg13g2_decap_8 FILLER_10_849 ();
 sg13g2_decap_8 FILLER_10_856 ();
 sg13g2_decap_8 FILLER_10_863 ();
 sg13g2_decap_8 FILLER_10_870 ();
 sg13g2_fill_1 FILLER_10_877 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_4 FILLER_11_371 ();
 sg13g2_fill_2 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_390 ();
 sg13g2_decap_4 FILLER_11_397 ();
 sg13g2_fill_2 FILLER_11_401 ();
 sg13g2_decap_4 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_419 ();
 sg13g2_decap_4 FILLER_11_431 ();
 sg13g2_decap_8 FILLER_11_457 ();
 sg13g2_decap_8 FILLER_11_464 ();
 sg13g2_decap_8 FILLER_11_471 ();
 sg13g2_fill_2 FILLER_11_478 ();
 sg13g2_fill_1 FILLER_11_480 ();
 sg13g2_decap_8 FILLER_11_486 ();
 sg13g2_decap_8 FILLER_11_493 ();
 sg13g2_decap_4 FILLER_11_500 ();
 sg13g2_fill_1 FILLER_11_504 ();
 sg13g2_fill_1 FILLER_11_523 ();
 sg13g2_decap_8 FILLER_11_528 ();
 sg13g2_decap_8 FILLER_11_535 ();
 sg13g2_fill_2 FILLER_11_542 ();
 sg13g2_decap_4 FILLER_11_557 ();
 sg13g2_fill_2 FILLER_11_561 ();
 sg13g2_decap_8 FILLER_11_576 ();
 sg13g2_decap_8 FILLER_11_583 ();
 sg13g2_decap_8 FILLER_11_590 ();
 sg13g2_decap_8 FILLER_11_597 ();
 sg13g2_decap_8 FILLER_11_604 ();
 sg13g2_decap_8 FILLER_11_611 ();
 sg13g2_fill_2 FILLER_11_618 ();
 sg13g2_fill_1 FILLER_11_620 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_662 ();
 sg13g2_decap_8 FILLER_11_669 ();
 sg13g2_decap_4 FILLER_11_676 ();
 sg13g2_fill_1 FILLER_11_680 ();
 sg13g2_decap_8 FILLER_11_694 ();
 sg13g2_decap_8 FILLER_11_701 ();
 sg13g2_decap_8 FILLER_11_708 ();
 sg13g2_decap_8 FILLER_11_715 ();
 sg13g2_decap_8 FILLER_11_722 ();
 sg13g2_decap_8 FILLER_11_729 ();
 sg13g2_decap_4 FILLER_11_741 ();
 sg13g2_fill_1 FILLER_11_745 ();
 sg13g2_decap_8 FILLER_11_752 ();
 sg13g2_decap_8 FILLER_11_759 ();
 sg13g2_decap_8 FILLER_11_766 ();
 sg13g2_decap_8 FILLER_11_773 ();
 sg13g2_decap_8 FILLER_11_780 ();
 sg13g2_decap_8 FILLER_11_787 ();
 sg13g2_decap_8 FILLER_11_794 ();
 sg13g2_decap_8 FILLER_11_801 ();
 sg13g2_decap_8 FILLER_11_808 ();
 sg13g2_decap_8 FILLER_11_815 ();
 sg13g2_decap_8 FILLER_11_822 ();
 sg13g2_decap_8 FILLER_11_829 ();
 sg13g2_decap_8 FILLER_11_836 ();
 sg13g2_decap_8 FILLER_11_843 ();
 sg13g2_decap_8 FILLER_11_850 ();
 sg13g2_decap_8 FILLER_11_857 ();
 sg13g2_decap_8 FILLER_11_864 ();
 sg13g2_decap_8 FILLER_11_871 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_fill_2 FILLER_12_273 ();
 sg13g2_fill_1 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_285 ();
 sg13g2_decap_4 FILLER_12_292 ();
 sg13g2_decap_8 FILLER_12_304 ();
 sg13g2_decap_8 FILLER_12_311 ();
 sg13g2_decap_8 FILLER_12_318 ();
 sg13g2_decap_8 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_332 ();
 sg13g2_decap_8 FILLER_12_339 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_fill_1 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_379 ();
 sg13g2_decap_4 FILLER_12_386 ();
 sg13g2_fill_2 FILLER_12_394 ();
 sg13g2_fill_1 FILLER_12_396 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_decap_4 FILLER_12_408 ();
 sg13g2_fill_1 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_433 ();
 sg13g2_decap_8 FILLER_12_440 ();
 sg13g2_decap_8 FILLER_12_447 ();
 sg13g2_decap_8 FILLER_12_454 ();
 sg13g2_decap_8 FILLER_12_461 ();
 sg13g2_decap_8 FILLER_12_468 ();
 sg13g2_decap_8 FILLER_12_480 ();
 sg13g2_decap_8 FILLER_12_491 ();
 sg13g2_decap_8 FILLER_12_498 ();
 sg13g2_decap_8 FILLER_12_505 ();
 sg13g2_decap_8 FILLER_12_512 ();
 sg13g2_fill_1 FILLER_12_519 ();
 sg13g2_decap_8 FILLER_12_529 ();
 sg13g2_decap_4 FILLER_12_536 ();
 sg13g2_fill_1 FILLER_12_540 ();
 sg13g2_decap_8 FILLER_12_549 ();
 sg13g2_decap_8 FILLER_12_556 ();
 sg13g2_decap_8 FILLER_12_563 ();
 sg13g2_decap_8 FILLER_12_570 ();
 sg13g2_decap_8 FILLER_12_577 ();
 sg13g2_decap_4 FILLER_12_584 ();
 sg13g2_decap_8 FILLER_12_593 ();
 sg13g2_decap_8 FILLER_12_608 ();
 sg13g2_decap_8 FILLER_12_615 ();
 sg13g2_decap_8 FILLER_12_622 ();
 sg13g2_decap_8 FILLER_12_629 ();
 sg13g2_decap_8 FILLER_12_636 ();
 sg13g2_decap_4 FILLER_12_643 ();
 sg13g2_fill_2 FILLER_12_647 ();
 sg13g2_decap_8 FILLER_12_654 ();
 sg13g2_decap_8 FILLER_12_661 ();
 sg13g2_decap_4 FILLER_12_668 ();
 sg13g2_decap_4 FILLER_12_676 ();
 sg13g2_decap_8 FILLER_12_684 ();
 sg13g2_fill_1 FILLER_12_691 ();
 sg13g2_decap_8 FILLER_12_705 ();
 sg13g2_decap_8 FILLER_12_712 ();
 sg13g2_fill_2 FILLER_12_719 ();
 sg13g2_fill_1 FILLER_12_721 ();
 sg13g2_fill_1 FILLER_12_754 ();
 sg13g2_decap_8 FILLER_12_765 ();
 sg13g2_decap_8 FILLER_12_776 ();
 sg13g2_decap_8 FILLER_12_783 ();
 sg13g2_decap_8 FILLER_12_790 ();
 sg13g2_decap_8 FILLER_12_797 ();
 sg13g2_decap_8 FILLER_12_804 ();
 sg13g2_decap_8 FILLER_12_811 ();
 sg13g2_decap_8 FILLER_12_818 ();
 sg13g2_decap_8 FILLER_12_825 ();
 sg13g2_decap_8 FILLER_12_832 ();
 sg13g2_decap_8 FILLER_12_839 ();
 sg13g2_decap_8 FILLER_12_846 ();
 sg13g2_decap_8 FILLER_12_853 ();
 sg13g2_decap_8 FILLER_12_860 ();
 sg13g2_decap_8 FILLER_12_867 ();
 sg13g2_decap_4 FILLER_12_874 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_4 FILLER_13_238 ();
 sg13g2_fill_2 FILLER_13_242 ();
 sg13g2_decap_4 FILLER_13_251 ();
 sg13g2_fill_1 FILLER_13_255 ();
 sg13g2_decap_8 FILLER_13_260 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_decap_8 FILLER_13_271 ();
 sg13g2_decap_8 FILLER_13_278 ();
 sg13g2_fill_2 FILLER_13_293 ();
 sg13g2_fill_1 FILLER_13_299 ();
 sg13g2_decap_4 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_317 ();
 sg13g2_decap_8 FILLER_13_324 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_fill_2 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_351 ();
 sg13g2_decap_8 FILLER_13_358 ();
 sg13g2_fill_2 FILLER_13_365 ();
 sg13g2_fill_2 FILLER_13_371 ();
 sg13g2_fill_1 FILLER_13_373 ();
 sg13g2_fill_2 FILLER_13_377 ();
 sg13g2_fill_1 FILLER_13_379 ();
 sg13g2_decap_4 FILLER_13_386 ();
 sg13g2_fill_1 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_decap_8 FILLER_13_407 ();
 sg13g2_fill_2 FILLER_13_439 ();
 sg13g2_decap_8 FILLER_13_445 ();
 sg13g2_decap_8 FILLER_13_452 ();
 sg13g2_decap_8 FILLER_13_459 ();
 sg13g2_decap_8 FILLER_13_466 ();
 sg13g2_decap_8 FILLER_13_473 ();
 sg13g2_fill_2 FILLER_13_480 ();
 sg13g2_decap_8 FILLER_13_486 ();
 sg13g2_decap_8 FILLER_13_493 ();
 sg13g2_decap_8 FILLER_13_500 ();
 sg13g2_decap_8 FILLER_13_507 ();
 sg13g2_decap_8 FILLER_13_514 ();
 sg13g2_decap_4 FILLER_13_521 ();
 sg13g2_decap_8 FILLER_13_533 ();
 sg13g2_decap_4 FILLER_13_545 ();
 sg13g2_fill_2 FILLER_13_549 ();
 sg13g2_fill_1 FILLER_13_560 ();
 sg13g2_decap_4 FILLER_13_565 ();
 sg13g2_fill_2 FILLER_13_569 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_fill_1 FILLER_13_581 ();
 sg13g2_fill_2 FILLER_13_599 ();
 sg13g2_fill_1 FILLER_13_605 ();
 sg13g2_decap_4 FILLER_13_610 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_fill_1 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_648 ();
 sg13g2_decap_8 FILLER_13_655 ();
 sg13g2_decap_8 FILLER_13_662 ();
 sg13g2_decap_4 FILLER_13_669 ();
 sg13g2_fill_2 FILLER_13_673 ();
 sg13g2_decap_4 FILLER_13_680 ();
 sg13g2_fill_1 FILLER_13_684 ();
 sg13g2_fill_1 FILLER_13_690 ();
 sg13g2_decap_8 FILLER_13_704 ();
 sg13g2_decap_8 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_718 ();
 sg13g2_decap_8 FILLER_13_730 ();
 sg13g2_fill_1 FILLER_13_737 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_4 FILLER_13_763 ();
 sg13g2_fill_2 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_774 ();
 sg13g2_decap_8 FILLER_13_781 ();
 sg13g2_decap_8 FILLER_13_788 ();
 sg13g2_decap_8 FILLER_13_795 ();
 sg13g2_decap_8 FILLER_13_802 ();
 sg13g2_decap_8 FILLER_13_809 ();
 sg13g2_decap_8 FILLER_13_816 ();
 sg13g2_decap_8 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_8 FILLER_13_844 ();
 sg13g2_decap_8 FILLER_13_851 ();
 sg13g2_decap_8 FILLER_13_858 ();
 sg13g2_decap_8 FILLER_13_865 ();
 sg13g2_decap_4 FILLER_13_872 ();
 sg13g2_fill_2 FILLER_13_876 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_fill_2 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_241 ();
 sg13g2_decap_8 FILLER_14_248 ();
 sg13g2_fill_2 FILLER_14_255 ();
 sg13g2_fill_1 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_4 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_4 FILLER_14_292 ();
 sg13g2_fill_2 FILLER_14_296 ();
 sg13g2_fill_2 FILLER_14_303 ();
 sg13g2_decap_4 FILLER_14_310 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_fill_2 FILLER_14_320 ();
 sg13g2_fill_1 FILLER_14_322 ();
 sg13g2_fill_2 FILLER_14_331 ();
 sg13g2_fill_1 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_decap_4 FILLER_14_349 ();
 sg13g2_decap_4 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_4 FILLER_14_406 ();
 sg13g2_fill_2 FILLER_14_410 ();
 sg13g2_decap_8 FILLER_14_416 ();
 sg13g2_fill_2 FILLER_14_423 ();
 sg13g2_fill_1 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_435 ();
 sg13g2_decap_8 FILLER_14_440 ();
 sg13g2_decap_8 FILLER_14_447 ();
 sg13g2_decap_8 FILLER_14_454 ();
 sg13g2_decap_8 FILLER_14_461 ();
 sg13g2_decap_8 FILLER_14_468 ();
 sg13g2_decap_8 FILLER_14_475 ();
 sg13g2_decap_8 FILLER_14_486 ();
 sg13g2_decap_8 FILLER_14_493 ();
 sg13g2_fill_2 FILLER_14_500 ();
 sg13g2_fill_2 FILLER_14_506 ();
 sg13g2_fill_2 FILLER_14_514 ();
 sg13g2_fill_1 FILLER_14_516 ();
 sg13g2_decap_8 FILLER_14_523 ();
 sg13g2_decap_8 FILLER_14_530 ();
 sg13g2_decap_8 FILLER_14_537 ();
 sg13g2_decap_8 FILLER_14_544 ();
 sg13g2_fill_2 FILLER_14_551 ();
 sg13g2_fill_1 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_562 ();
 sg13g2_fill_2 FILLER_14_569 ();
 sg13g2_decap_8 FILLER_14_575 ();
 sg13g2_decap_8 FILLER_14_582 ();
 sg13g2_decap_4 FILLER_14_589 ();
 sg13g2_fill_2 FILLER_14_593 ();
 sg13g2_decap_4 FILLER_14_599 ();
 sg13g2_fill_2 FILLER_14_603 ();
 sg13g2_decap_8 FILLER_14_613 ();
 sg13g2_decap_8 FILLER_14_620 ();
 sg13g2_decap_8 FILLER_14_627 ();
 sg13g2_decap_4 FILLER_14_634 ();
 sg13g2_fill_1 FILLER_14_638 ();
 sg13g2_decap_4 FILLER_14_644 ();
 sg13g2_fill_2 FILLER_14_648 ();
 sg13g2_decap_4 FILLER_14_663 ();
 sg13g2_fill_2 FILLER_14_667 ();
 sg13g2_decap_8 FILLER_14_678 ();
 sg13g2_decap_8 FILLER_14_685 ();
 sg13g2_decap_8 FILLER_14_692 ();
 sg13g2_decap_4 FILLER_14_699 ();
 sg13g2_fill_2 FILLER_14_703 ();
 sg13g2_decap_8 FILLER_14_709 ();
 sg13g2_decap_4 FILLER_14_716 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_fill_1 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_783 ();
 sg13g2_decap_8 FILLER_14_790 ();
 sg13g2_decap_8 FILLER_14_797 ();
 sg13g2_decap_8 FILLER_14_804 ();
 sg13g2_decap_8 FILLER_14_811 ();
 sg13g2_decap_8 FILLER_14_818 ();
 sg13g2_decap_8 FILLER_14_825 ();
 sg13g2_decap_8 FILLER_14_832 ();
 sg13g2_decap_8 FILLER_14_839 ();
 sg13g2_decap_8 FILLER_14_846 ();
 sg13g2_decap_8 FILLER_14_853 ();
 sg13g2_decap_8 FILLER_14_860 ();
 sg13g2_decap_8 FILLER_14_867 ();
 sg13g2_decap_4 FILLER_14_874 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_4 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_155 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_decap_4 FILLER_15_166 ();
 sg13g2_fill_1 FILLER_15_170 ();
 sg13g2_decap_8 FILLER_15_187 ();
 sg13g2_fill_2 FILLER_15_194 ();
 sg13g2_fill_1 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_202 ();
 sg13g2_fill_2 FILLER_15_209 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_decap_4 FILLER_15_217 ();
 sg13g2_fill_1 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_234 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_4 FILLER_15_255 ();
 sg13g2_fill_1 FILLER_15_259 ();
 sg13g2_decap_4 FILLER_15_271 ();
 sg13g2_fill_2 FILLER_15_275 ();
 sg13g2_decap_8 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_289 ();
 sg13g2_fill_1 FILLER_15_296 ();
 sg13g2_decap_8 FILLER_15_310 ();
 sg13g2_decap_8 FILLER_15_317 ();
 sg13g2_decap_8 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_331 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_decap_8 FILLER_15_342 ();
 sg13g2_fill_2 FILLER_15_349 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_4 FILLER_15_363 ();
 sg13g2_fill_2 FILLER_15_367 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_fill_2 FILLER_15_396 ();
 sg13g2_fill_1 FILLER_15_398 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_fill_1 FILLER_15_409 ();
 sg13g2_decap_8 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_decap_8 FILLER_15_429 ();
 sg13g2_fill_2 FILLER_15_436 ();
 sg13g2_fill_2 FILLER_15_441 ();
 sg13g2_fill_1 FILLER_15_443 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_fill_2 FILLER_15_473 ();
 sg13g2_fill_1 FILLER_15_475 ();
 sg13g2_decap_4 FILLER_15_481 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_509 ();
 sg13g2_decap_8 FILLER_15_516 ();
 sg13g2_decap_8 FILLER_15_523 ();
 sg13g2_decap_8 FILLER_15_530 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_fill_1 FILLER_15_564 ();
 sg13g2_decap_4 FILLER_15_575 ();
 sg13g2_decap_8 FILLER_15_585 ();
 sg13g2_decap_8 FILLER_15_592 ();
 sg13g2_decap_8 FILLER_15_599 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_decap_8 FILLER_15_613 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_8 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_decap_4 FILLER_15_648 ();
 sg13g2_decap_4 FILLER_15_656 ();
 sg13g2_decap_8 FILLER_15_682 ();
 sg13g2_fill_2 FILLER_15_689 ();
 sg13g2_decap_4 FILLER_15_709 ();
 sg13g2_decap_4 FILLER_15_719 ();
 sg13g2_decap_8 FILLER_15_727 ();
 sg13g2_decap_4 FILLER_15_739 ();
 sg13g2_decap_8 FILLER_15_747 ();
 sg13g2_decap_8 FILLER_15_754 ();
 sg13g2_decap_8 FILLER_15_761 ();
 sg13g2_decap_8 FILLER_15_768 ();
 sg13g2_decap_8 FILLER_15_775 ();
 sg13g2_decap_8 FILLER_15_782 ();
 sg13g2_decap_8 FILLER_15_789 ();
 sg13g2_decap_8 FILLER_15_796 ();
 sg13g2_decap_8 FILLER_15_803 ();
 sg13g2_decap_8 FILLER_15_810 ();
 sg13g2_decap_8 FILLER_15_817 ();
 sg13g2_decap_8 FILLER_15_824 ();
 sg13g2_decap_8 FILLER_15_831 ();
 sg13g2_decap_8 FILLER_15_838 ();
 sg13g2_decap_8 FILLER_15_845 ();
 sg13g2_decap_8 FILLER_15_852 ();
 sg13g2_decap_8 FILLER_15_859 ();
 sg13g2_decap_8 FILLER_15_866 ();
 sg13g2_decap_4 FILLER_15_873 ();
 sg13g2_fill_1 FILLER_15_877 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_decap_4 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_decap_4 FILLER_16_194 ();
 sg13g2_fill_2 FILLER_16_202 ();
 sg13g2_fill_1 FILLER_16_204 ();
 sg13g2_fill_1 FILLER_16_209 ();
 sg13g2_decap_4 FILLER_16_214 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_233 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_fill_1 FILLER_16_252 ();
 sg13g2_decap_4 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_decap_8 FILLER_16_281 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_fill_1 FILLER_16_295 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_fill_1 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_4 FILLER_16_387 ();
 sg13g2_fill_1 FILLER_16_391 ();
 sg13g2_fill_2 FILLER_16_409 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_16_424 ();
 sg13g2_fill_2 FILLER_16_431 ();
 sg13g2_fill_1 FILLER_16_433 ();
 sg13g2_fill_2 FILLER_16_459 ();
 sg13g2_fill_2 FILLER_16_469 ();
 sg13g2_fill_1 FILLER_16_471 ();
 sg13g2_fill_2 FILLER_16_483 ();
 sg13g2_fill_2 FILLER_16_491 ();
 sg13g2_decap_4 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_507 ();
 sg13g2_decap_8 FILLER_16_514 ();
 sg13g2_decap_4 FILLER_16_521 ();
 sg13g2_decap_8 FILLER_16_529 ();
 sg13g2_decap_8 FILLER_16_536 ();
 sg13g2_decap_8 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_550 ();
 sg13g2_decap_8 FILLER_16_557 ();
 sg13g2_decap_4 FILLER_16_564 ();
 sg13g2_decap_8 FILLER_16_589 ();
 sg13g2_decap_8 FILLER_16_596 ();
 sg13g2_decap_4 FILLER_16_603 ();
 sg13g2_decap_8 FILLER_16_619 ();
 sg13g2_decap_8 FILLER_16_626 ();
 sg13g2_decap_8 FILLER_16_633 ();
 sg13g2_fill_2 FILLER_16_640 ();
 sg13g2_fill_2 FILLER_16_646 ();
 sg13g2_fill_1 FILLER_16_648 ();
 sg13g2_fill_1 FILLER_16_654 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_4 FILLER_16_672 ();
 sg13g2_fill_1 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_681 ();
 sg13g2_decap_4 FILLER_16_688 ();
 sg13g2_fill_1 FILLER_16_692 ();
 sg13g2_decap_4 FILLER_16_698 ();
 sg13g2_fill_1 FILLER_16_702 ();
 sg13g2_decap_4 FILLER_16_708 ();
 sg13g2_fill_1 FILLER_16_712 ();
 sg13g2_decap_4 FILLER_16_722 ();
 sg13g2_fill_2 FILLER_16_726 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_fill_1 FILLER_16_753 ();
 sg13g2_decap_4 FILLER_16_762 ();
 sg13g2_fill_2 FILLER_16_766 ();
 sg13g2_decap_8 FILLER_16_780 ();
 sg13g2_decap_8 FILLER_16_787 ();
 sg13g2_decap_8 FILLER_16_794 ();
 sg13g2_decap_8 FILLER_16_801 ();
 sg13g2_decap_8 FILLER_16_808 ();
 sg13g2_decap_8 FILLER_16_815 ();
 sg13g2_decap_8 FILLER_16_822 ();
 sg13g2_decap_8 FILLER_16_829 ();
 sg13g2_decap_8 FILLER_16_836 ();
 sg13g2_decap_8 FILLER_16_843 ();
 sg13g2_decap_8 FILLER_16_850 ();
 sg13g2_decap_8 FILLER_16_857 ();
 sg13g2_decap_8 FILLER_16_864 ();
 sg13g2_decap_8 FILLER_16_871 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_132 ();
 sg13g2_decap_4 FILLER_17_139 ();
 sg13g2_fill_1 FILLER_17_143 ();
 sg13g2_decap_4 FILLER_17_149 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_decap_4 FILLER_17_182 ();
 sg13g2_fill_1 FILLER_17_186 ();
 sg13g2_decap_8 FILLER_17_200 ();
 sg13g2_decap_4 FILLER_17_212 ();
 sg13g2_fill_2 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_fill_2 FILLER_17_242 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_fill_2 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_255 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_4 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_fill_2 FILLER_17_331 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_338 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_decap_8 FILLER_17_352 ();
 sg13g2_decap_8 FILLER_17_359 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_17_387 ();
 sg13g2_decap_8 FILLER_17_394 ();
 sg13g2_fill_1 FILLER_17_401 ();
 sg13g2_decap_8 FILLER_17_411 ();
 sg13g2_decap_4 FILLER_17_418 ();
 sg13g2_fill_1 FILLER_17_422 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_fill_2 FILLER_17_436 ();
 sg13g2_fill_1 FILLER_17_438 ();
 sg13g2_fill_2 FILLER_17_442 ();
 sg13g2_fill_1 FILLER_17_449 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_500 ();
 sg13g2_decap_8 FILLER_17_507 ();
 sg13g2_decap_8 FILLER_17_514 ();
 sg13g2_decap_8 FILLER_17_521 ();
 sg13g2_decap_8 FILLER_17_528 ();
 sg13g2_decap_8 FILLER_17_535 ();
 sg13g2_decap_8 FILLER_17_542 ();
 sg13g2_fill_2 FILLER_17_549 ();
 sg13g2_fill_1 FILLER_17_551 ();
 sg13g2_decap_8 FILLER_17_556 ();
 sg13g2_decap_4 FILLER_17_563 ();
 sg13g2_fill_1 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_573 ();
 sg13g2_decap_4 FILLER_17_580 ();
 sg13g2_fill_1 FILLER_17_584 ();
 sg13g2_decap_8 FILLER_17_589 ();
 sg13g2_fill_1 FILLER_17_596 ();
 sg13g2_decap_8 FILLER_17_607 ();
 sg13g2_decap_8 FILLER_17_614 ();
 sg13g2_decap_8 FILLER_17_621 ();
 sg13g2_fill_1 FILLER_17_628 ();
 sg13g2_decap_8 FILLER_17_634 ();
 sg13g2_decap_8 FILLER_17_641 ();
 sg13g2_fill_1 FILLER_17_648 ();
 sg13g2_decap_8 FILLER_17_662 ();
 sg13g2_decap_8 FILLER_17_669 ();
 sg13g2_decap_8 FILLER_17_676 ();
 sg13g2_decap_8 FILLER_17_683 ();
 sg13g2_decap_8 FILLER_17_690 ();
 sg13g2_decap_8 FILLER_17_697 ();
 sg13g2_decap_4 FILLER_17_704 ();
 sg13g2_decap_8 FILLER_17_712 ();
 sg13g2_decap_8 FILLER_17_719 ();
 sg13g2_decap_8 FILLER_17_726 ();
 sg13g2_decap_8 FILLER_17_733 ();
 sg13g2_fill_1 FILLER_17_740 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_fill_1 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_772 ();
 sg13g2_decap_8 FILLER_17_779 ();
 sg13g2_decap_8 FILLER_17_786 ();
 sg13g2_decap_8 FILLER_17_793 ();
 sg13g2_decap_8 FILLER_17_800 ();
 sg13g2_decap_8 FILLER_17_807 ();
 sg13g2_decap_8 FILLER_17_814 ();
 sg13g2_decap_8 FILLER_17_821 ();
 sg13g2_decap_8 FILLER_17_828 ();
 sg13g2_decap_8 FILLER_17_835 ();
 sg13g2_decap_8 FILLER_17_842 ();
 sg13g2_decap_8 FILLER_17_849 ();
 sg13g2_decap_8 FILLER_17_856 ();
 sg13g2_decap_8 FILLER_17_863 ();
 sg13g2_decap_8 FILLER_17_870 ();
 sg13g2_fill_1 FILLER_17_877 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_117 ();
 sg13g2_decap_8 FILLER_18_124 ();
 sg13g2_decap_4 FILLER_18_131 ();
 sg13g2_fill_1 FILLER_18_135 ();
 sg13g2_decap_4 FILLER_18_141 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_decap_8 FILLER_18_173 ();
 sg13g2_decap_4 FILLER_18_180 ();
 sg13g2_decap_4 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_4 FILLER_18_207 ();
 sg13g2_fill_2 FILLER_18_211 ();
 sg13g2_decap_8 FILLER_18_218 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_234 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_decap_4 FILLER_18_263 ();
 sg13g2_fill_2 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_272 ();
 sg13g2_decap_4 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_297 ();
 sg13g2_decap_4 FILLER_18_304 ();
 sg13g2_fill_2 FILLER_18_308 ();
 sg13g2_fill_2 FILLER_18_314 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_4 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_fill_1 FILLER_18_366 ();
 sg13g2_fill_1 FILLER_18_372 ();
 sg13g2_fill_2 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_8 FILLER_18_403 ();
 sg13g2_decap_4 FILLER_18_410 ();
 sg13g2_decap_8 FILLER_18_422 ();
 sg13g2_decap_4 FILLER_18_429 ();
 sg13g2_fill_1 FILLER_18_433 ();
 sg13g2_fill_2 FILLER_18_439 ();
 sg13g2_decap_8 FILLER_18_446 ();
 sg13g2_decap_8 FILLER_18_453 ();
 sg13g2_decap_8 FILLER_18_460 ();
 sg13g2_decap_8 FILLER_18_467 ();
 sg13g2_fill_2 FILLER_18_474 ();
 sg13g2_fill_1 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_481 ();
 sg13g2_decap_8 FILLER_18_488 ();
 sg13g2_decap_4 FILLER_18_495 ();
 sg13g2_fill_2 FILLER_18_499 ();
 sg13g2_decap_4 FILLER_18_510 ();
 sg13g2_decap_4 FILLER_18_518 ();
 sg13g2_fill_2 FILLER_18_522 ();
 sg13g2_decap_4 FILLER_18_528 ();
 sg13g2_fill_1 FILLER_18_537 ();
 sg13g2_decap_8 FILLER_18_542 ();
 sg13g2_fill_1 FILLER_18_549 ();
 sg13g2_decap_4 FILLER_18_562 ();
 sg13g2_decap_4 FILLER_18_576 ();
 sg13g2_decap_4 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_597 ();
 sg13g2_decap_8 FILLER_18_604 ();
 sg13g2_decap_8 FILLER_18_611 ();
 sg13g2_decap_8 FILLER_18_618 ();
 sg13g2_decap_8 FILLER_18_625 ();
 sg13g2_decap_8 FILLER_18_632 ();
 sg13g2_decap_4 FILLER_18_639 ();
 sg13g2_decap_8 FILLER_18_653 ();
 sg13g2_decap_8 FILLER_18_660 ();
 sg13g2_decap_4 FILLER_18_667 ();
 sg13g2_fill_1 FILLER_18_671 ();
 sg13g2_decap_8 FILLER_18_677 ();
 sg13g2_decap_8 FILLER_18_684 ();
 sg13g2_decap_8 FILLER_18_691 ();
 sg13g2_fill_2 FILLER_18_698 ();
 sg13g2_decap_8 FILLER_18_717 ();
 sg13g2_decap_4 FILLER_18_724 ();
 sg13g2_fill_2 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_785 ();
 sg13g2_decap_8 FILLER_18_792 ();
 sg13g2_decap_8 FILLER_18_799 ();
 sg13g2_decap_8 FILLER_18_806 ();
 sg13g2_decap_8 FILLER_18_813 ();
 sg13g2_decap_8 FILLER_18_820 ();
 sg13g2_decap_8 FILLER_18_827 ();
 sg13g2_decap_8 FILLER_18_834 ();
 sg13g2_decap_8 FILLER_18_841 ();
 sg13g2_decap_8 FILLER_18_848 ();
 sg13g2_decap_8 FILLER_18_855 ();
 sg13g2_decap_8 FILLER_18_862 ();
 sg13g2_decap_8 FILLER_18_869 ();
 sg13g2_fill_2 FILLER_18_876 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_117 ();
 sg13g2_decap_8 FILLER_19_124 ();
 sg13g2_fill_1 FILLER_19_131 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_decap_4 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_159 ();
 sg13g2_decap_4 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_decap_4 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_decap_8 FILLER_19_229 ();
 sg13g2_decap_8 FILLER_19_240 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_fill_1 FILLER_19_269 ();
 sg13g2_decap_4 FILLER_19_275 ();
 sg13g2_decap_8 FILLER_19_283 ();
 sg13g2_decap_4 FILLER_19_294 ();
 sg13g2_fill_2 FILLER_19_307 ();
 sg13g2_fill_1 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_fill_2 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_363 ();
 sg13g2_decap_4 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_8 FILLER_19_405 ();
 sg13g2_decap_4 FILLER_19_412 ();
 sg13g2_fill_2 FILLER_19_416 ();
 sg13g2_decap_8 FILLER_19_422 ();
 sg13g2_fill_2 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_19_436 ();
 sg13g2_decap_8 FILLER_19_443 ();
 sg13g2_fill_1 FILLER_19_450 ();
 sg13g2_fill_1 FILLER_19_460 ();
 sg13g2_decap_8 FILLER_19_466 ();
 sg13g2_fill_2 FILLER_19_473 ();
 sg13g2_fill_1 FILLER_19_475 ();
 sg13g2_decap_8 FILLER_19_480 ();
 sg13g2_fill_2 FILLER_19_487 ();
 sg13g2_decap_4 FILLER_19_493 ();
 sg13g2_fill_2 FILLER_19_500 ();
 sg13g2_fill_2 FILLER_19_511 ();
 sg13g2_fill_1 FILLER_19_513 ();
 sg13g2_decap_8 FILLER_19_522 ();
 sg13g2_fill_2 FILLER_19_529 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_4 FILLER_19_546 ();
 sg13g2_fill_2 FILLER_19_550 ();
 sg13g2_fill_1 FILLER_19_556 ();
 sg13g2_decap_8 FILLER_19_561 ();
 sg13g2_fill_2 FILLER_19_568 ();
 sg13g2_fill_2 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_586 ();
 sg13g2_fill_2 FILLER_19_593 ();
 sg13g2_decap_8 FILLER_19_599 ();
 sg13g2_decap_8 FILLER_19_606 ();
 sg13g2_decap_8 FILLER_19_613 ();
 sg13g2_decap_8 FILLER_19_629 ();
 sg13g2_fill_1 FILLER_19_636 ();
 sg13g2_decap_8 FILLER_19_641 ();
 sg13g2_decap_8 FILLER_19_648 ();
 sg13g2_decap_8 FILLER_19_655 ();
 sg13g2_fill_2 FILLER_19_662 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_decap_8 FILLER_19_676 ();
 sg13g2_decap_8 FILLER_19_683 ();
 sg13g2_decap_8 FILLER_19_690 ();
 sg13g2_decap_4 FILLER_19_697 ();
 sg13g2_fill_2 FILLER_19_701 ();
 sg13g2_decap_4 FILLER_19_707 ();
 sg13g2_fill_2 FILLER_19_711 ();
 sg13g2_decap_8 FILLER_19_722 ();
 sg13g2_decap_8 FILLER_19_729 ();
 sg13g2_decap_8 FILLER_19_736 ();
 sg13g2_decap_8 FILLER_19_743 ();
 sg13g2_decap_8 FILLER_19_750 ();
 sg13g2_decap_4 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_778 ();
 sg13g2_decap_8 FILLER_19_785 ();
 sg13g2_decap_8 FILLER_19_792 ();
 sg13g2_decap_8 FILLER_19_799 ();
 sg13g2_decap_8 FILLER_19_806 ();
 sg13g2_decap_8 FILLER_19_813 ();
 sg13g2_decap_8 FILLER_19_820 ();
 sg13g2_decap_8 FILLER_19_827 ();
 sg13g2_decap_8 FILLER_19_834 ();
 sg13g2_decap_8 FILLER_19_841 ();
 sg13g2_decap_8 FILLER_19_848 ();
 sg13g2_decap_8 FILLER_19_855 ();
 sg13g2_decap_8 FILLER_19_862 ();
 sg13g2_decap_8 FILLER_19_869 ();
 sg13g2_fill_2 FILLER_19_876 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_4 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_114 ();
 sg13g2_decap_8 FILLER_20_121 ();
 sg13g2_decap_8 FILLER_20_128 ();
 sg13g2_decap_8 FILLER_20_135 ();
 sg13g2_decap_8 FILLER_20_142 ();
 sg13g2_decap_8 FILLER_20_149 ();
 sg13g2_decap_8 FILLER_20_156 ();
 sg13g2_fill_1 FILLER_20_163 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_177 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_196 ();
 sg13g2_fill_1 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_211 ();
 sg13g2_fill_2 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_220 ();
 sg13g2_fill_2 FILLER_20_225 ();
 sg13g2_decap_8 FILLER_20_232 ();
 sg13g2_decap_4 FILLER_20_244 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_decap_8 FILLER_20_262 ();
 sg13g2_decap_8 FILLER_20_269 ();
 sg13g2_decap_4 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_decap_4 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_decap_8 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_314 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_decap_8 FILLER_20_328 ();
 sg13g2_decap_8 FILLER_20_335 ();
 sg13g2_decap_8 FILLER_20_342 ();
 sg13g2_decap_8 FILLER_20_349 ();
 sg13g2_decap_8 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_363 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_4 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_404 ();
 sg13g2_decap_8 FILLER_20_411 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_fill_2 FILLER_20_425 ();
 sg13g2_decap_8 FILLER_20_436 ();
 sg13g2_fill_1 FILLER_20_443 ();
 sg13g2_fill_2 FILLER_20_449 ();
 sg13g2_fill_1 FILLER_20_456 ();
 sg13g2_decap_8 FILLER_20_481 ();
 sg13g2_fill_1 FILLER_20_488 ();
 sg13g2_decap_8 FILLER_20_506 ();
 sg13g2_decap_8 FILLER_20_513 ();
 sg13g2_decap_8 FILLER_20_520 ();
 sg13g2_fill_1 FILLER_20_527 ();
 sg13g2_decap_4 FILLER_20_533 ();
 sg13g2_fill_1 FILLER_20_541 ();
 sg13g2_decap_4 FILLER_20_549 ();
 sg13g2_decap_8 FILLER_20_557 ();
 sg13g2_decap_8 FILLER_20_564 ();
 sg13g2_fill_2 FILLER_20_571 ();
 sg13g2_decap_8 FILLER_20_593 ();
 sg13g2_decap_8 FILLER_20_600 ();
 sg13g2_fill_2 FILLER_20_607 ();
 sg13g2_fill_1 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_619 ();
 sg13g2_decap_8 FILLER_20_626 ();
 sg13g2_decap_4 FILLER_20_638 ();
 sg13g2_fill_2 FILLER_20_642 ();
 sg13g2_decap_8 FILLER_20_652 ();
 sg13g2_fill_1 FILLER_20_659 ();
 sg13g2_decap_4 FILLER_20_666 ();
 sg13g2_fill_2 FILLER_20_670 ();
 sg13g2_decap_8 FILLER_20_676 ();
 sg13g2_decap_4 FILLER_20_683 ();
 sg13g2_fill_1 FILLER_20_687 ();
 sg13g2_decap_4 FILLER_20_692 ();
 sg13g2_decap_8 FILLER_20_701 ();
 sg13g2_decap_4 FILLER_20_708 ();
 sg13g2_fill_2 FILLER_20_712 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_fill_1 FILLER_20_726 ();
 sg13g2_decap_8 FILLER_20_733 ();
 sg13g2_decap_8 FILLER_20_740 ();
 sg13g2_fill_2 FILLER_20_747 ();
 sg13g2_decap_8 FILLER_20_757 ();
 sg13g2_decap_4 FILLER_20_764 ();
 sg13g2_fill_1 FILLER_20_772 ();
 sg13g2_decap_8 FILLER_20_778 ();
 sg13g2_decap_8 FILLER_20_785 ();
 sg13g2_decap_8 FILLER_20_792 ();
 sg13g2_decap_8 FILLER_20_799 ();
 sg13g2_decap_8 FILLER_20_806 ();
 sg13g2_decap_8 FILLER_20_813 ();
 sg13g2_decap_8 FILLER_20_820 ();
 sg13g2_decap_8 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_decap_8 FILLER_20_841 ();
 sg13g2_decap_8 FILLER_20_848 ();
 sg13g2_decap_8 FILLER_20_855 ();
 sg13g2_decap_8 FILLER_20_862 ();
 sg13g2_decap_8 FILLER_20_869 ();
 sg13g2_fill_2 FILLER_20_876 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_decap_8 FILLER_21_136 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_fill_1 FILLER_21_157 ();
 sg13g2_decap_4 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_decap_8 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_194 ();
 sg13g2_decap_8 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_211 ();
 sg13g2_decap_4 FILLER_21_218 ();
 sg13g2_fill_1 FILLER_21_222 ();
 sg13g2_decap_8 FILLER_21_233 ();
 sg13g2_decap_4 FILLER_21_240 ();
 sg13g2_fill_1 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_254 ();
 sg13g2_decap_8 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_decap_8 FILLER_21_275 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_4 FILLER_21_294 ();
 sg13g2_fill_2 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_4 FILLER_21_319 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_fill_2 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_4 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_366 ();
 sg13g2_decap_4 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_2 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_21_415 ();
 sg13g2_decap_4 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_21_438 ();
 sg13g2_fill_1 FILLER_21_445 ();
 sg13g2_decap_8 FILLER_21_451 ();
 sg13g2_decap_8 FILLER_21_458 ();
 sg13g2_decap_8 FILLER_21_465 ();
 sg13g2_decap_8 FILLER_21_472 ();
 sg13g2_decap_4 FILLER_21_489 ();
 sg13g2_fill_2 FILLER_21_493 ();
 sg13g2_decap_8 FILLER_21_499 ();
 sg13g2_decap_8 FILLER_21_506 ();
 sg13g2_decap_8 FILLER_21_513 ();
 sg13g2_fill_2 FILLER_21_520 ();
 sg13g2_fill_1 FILLER_21_522 ();
 sg13g2_decap_8 FILLER_21_526 ();
 sg13g2_decap_8 FILLER_21_533 ();
 sg13g2_decap_8 FILLER_21_540 ();
 sg13g2_decap_8 FILLER_21_547 ();
 sg13g2_decap_8 FILLER_21_554 ();
 sg13g2_decap_4 FILLER_21_561 ();
 sg13g2_fill_1 FILLER_21_565 ();
 sg13g2_decap_8 FILLER_21_570 ();
 sg13g2_decap_4 FILLER_21_577 ();
 sg13g2_decap_8 FILLER_21_585 ();
 sg13g2_fill_2 FILLER_21_592 ();
 sg13g2_fill_1 FILLER_21_594 ();
 sg13g2_decap_8 FILLER_21_599 ();
 sg13g2_decap_4 FILLER_21_606 ();
 sg13g2_decap_4 FILLER_21_618 ();
 sg13g2_decap_8 FILLER_21_627 ();
 sg13g2_fill_2 FILLER_21_634 ();
 sg13g2_fill_1 FILLER_21_636 ();
 sg13g2_decap_8 FILLER_21_647 ();
 sg13g2_decap_8 FILLER_21_654 ();
 sg13g2_decap_4 FILLER_21_661 ();
 sg13g2_decap_4 FILLER_21_671 ();
 sg13g2_fill_2 FILLER_21_675 ();
 sg13g2_decap_4 FILLER_21_682 ();
 sg13g2_fill_2 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_696 ();
 sg13g2_decap_4 FILLER_21_703 ();
 sg13g2_fill_1 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_718 ();
 sg13g2_decap_8 FILLER_21_725 ();
 sg13g2_decap_8 FILLER_21_732 ();
 sg13g2_decap_8 FILLER_21_739 ();
 sg13g2_fill_2 FILLER_21_746 ();
 sg13g2_fill_1 FILLER_21_748 ();
 sg13g2_decap_8 FILLER_21_773 ();
 sg13g2_decap_8 FILLER_21_793 ();
 sg13g2_decap_8 FILLER_21_800 ();
 sg13g2_decap_8 FILLER_21_807 ();
 sg13g2_decap_8 FILLER_21_814 ();
 sg13g2_decap_8 FILLER_21_821 ();
 sg13g2_decap_8 FILLER_21_828 ();
 sg13g2_decap_8 FILLER_21_835 ();
 sg13g2_decap_8 FILLER_21_842 ();
 sg13g2_decap_8 FILLER_21_849 ();
 sg13g2_decap_8 FILLER_21_856 ();
 sg13g2_decap_8 FILLER_21_863 ();
 sg13g2_decap_8 FILLER_21_870 ();
 sg13g2_fill_1 FILLER_21_877 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_decap_8 FILLER_22_92 ();
 sg13g2_decap_4 FILLER_22_104 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_fill_2 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_decap_8 FILLER_22_132 ();
 sg13g2_decap_4 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_decap_4 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_174 ();
 sg13g2_decap_8 FILLER_22_181 ();
 sg13g2_decap_4 FILLER_22_188 ();
 sg13g2_fill_1 FILLER_22_192 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_decap_4 FILLER_22_205 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_fill_1 FILLER_22_222 ();
 sg13g2_fill_2 FILLER_22_226 ();
 sg13g2_decap_8 FILLER_22_232 ();
 sg13g2_decap_8 FILLER_22_239 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_fill_2 FILLER_22_253 ();
 sg13g2_decap_8 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_271 ();
 sg13g2_fill_2 FILLER_22_278 ();
 sg13g2_decap_8 FILLER_22_285 ();
 sg13g2_decap_8 FILLER_22_292 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_310 ();
 sg13g2_decap_4 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_4 FILLER_22_333 ();
 sg13g2_fill_2 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_4 FILLER_22_361 ();
 sg13g2_decap_4 FILLER_22_370 ();
 sg13g2_fill_1 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_4 FILLER_22_386 ();
 sg13g2_fill_1 FILLER_22_390 ();
 sg13g2_fill_1 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_fill_2 FILLER_22_413 ();
 sg13g2_decap_4 FILLER_22_419 ();
 sg13g2_decap_4 FILLER_22_431 ();
 sg13g2_fill_1 FILLER_22_435 ();
 sg13g2_decap_4 FILLER_22_445 ();
 sg13g2_decap_4 FILLER_22_453 ();
 sg13g2_decap_4 FILLER_22_461 ();
 sg13g2_fill_1 FILLER_22_465 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_4 FILLER_22_490 ();
 sg13g2_fill_2 FILLER_22_494 ();
 sg13g2_decap_8 FILLER_22_501 ();
 sg13g2_fill_2 FILLER_22_508 ();
 sg13g2_fill_1 FILLER_22_510 ();
 sg13g2_decap_8 FILLER_22_516 ();
 sg13g2_fill_2 FILLER_22_523 ();
 sg13g2_decap_4 FILLER_22_531 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_580 ();
 sg13g2_decap_8 FILLER_22_607 ();
 sg13g2_fill_1 FILLER_22_614 ();
 sg13g2_decap_8 FILLER_22_620 ();
 sg13g2_fill_1 FILLER_22_627 ();
 sg13g2_fill_2 FILLER_22_632 ();
 sg13g2_fill_1 FILLER_22_643 ();
 sg13g2_decap_8 FILLER_22_649 ();
 sg13g2_decap_8 FILLER_22_660 ();
 sg13g2_decap_4 FILLER_22_667 ();
 sg13g2_decap_8 FILLER_22_680 ();
 sg13g2_fill_2 FILLER_22_687 ();
 sg13g2_fill_1 FILLER_22_689 ();
 sg13g2_decap_8 FILLER_22_694 ();
 sg13g2_decap_8 FILLER_22_701 ();
 sg13g2_decap_8 FILLER_22_708 ();
 sg13g2_decap_4 FILLER_22_715 ();
 sg13g2_decap_8 FILLER_22_723 ();
 sg13g2_decap_8 FILLER_22_730 ();
 sg13g2_decap_8 FILLER_22_737 ();
 sg13g2_decap_8 FILLER_22_744 ();
 sg13g2_decap_8 FILLER_22_751 ();
 sg13g2_decap_8 FILLER_22_758 ();
 sg13g2_fill_1 FILLER_22_765 ();
 sg13g2_fill_1 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_776 ();
 sg13g2_decap_8 FILLER_22_783 ();
 sg13g2_decap_8 FILLER_22_790 ();
 sg13g2_decap_8 FILLER_22_797 ();
 sg13g2_decap_8 FILLER_22_804 ();
 sg13g2_decap_8 FILLER_22_811 ();
 sg13g2_decap_8 FILLER_22_818 ();
 sg13g2_decap_8 FILLER_22_825 ();
 sg13g2_decap_8 FILLER_22_832 ();
 sg13g2_decap_8 FILLER_22_839 ();
 sg13g2_decap_8 FILLER_22_846 ();
 sg13g2_decap_8 FILLER_22_853 ();
 sg13g2_decap_8 FILLER_22_860 ();
 sg13g2_decap_8 FILLER_22_867 ();
 sg13g2_decap_4 FILLER_22_874 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_72 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_fill_1 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_108 ();
 sg13g2_decap_4 FILLER_23_115 ();
 sg13g2_decap_4 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_131 ();
 sg13g2_fill_1 FILLER_23_133 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_fill_2 FILLER_23_154 ();
 sg13g2_fill_2 FILLER_23_165 ();
 sg13g2_fill_1 FILLER_23_167 ();
 sg13g2_decap_4 FILLER_23_173 ();
 sg13g2_fill_2 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_185 ();
 sg13g2_fill_2 FILLER_23_190 ();
 sg13g2_fill_1 FILLER_23_192 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_decap_4 FILLER_23_205 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_4 FILLER_23_228 ();
 sg13g2_fill_1 FILLER_23_232 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_4 FILLER_23_252 ();
 sg13g2_fill_1 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_262 ();
 sg13g2_decap_8 FILLER_23_269 ();
 sg13g2_decap_4 FILLER_23_276 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_fill_2 FILLER_23_287 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_fill_1 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_8 FILLER_23_356 ();
 sg13g2_decap_4 FILLER_23_363 ();
 sg13g2_fill_1 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_fill_2 FILLER_23_395 ();
 sg13g2_fill_1 FILLER_23_397 ();
 sg13g2_decap_8 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_23_412 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_fill_2 FILLER_23_426 ();
 sg13g2_decap_4 FILLER_23_458 ();
 sg13g2_fill_2 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_467 ();
 sg13g2_decap_8 FILLER_23_474 ();
 sg13g2_decap_8 FILLER_23_481 ();
 sg13g2_decap_4 FILLER_23_488 ();
 sg13g2_fill_2 FILLER_23_492 ();
 sg13g2_decap_8 FILLER_23_499 ();
 sg13g2_decap_8 FILLER_23_506 ();
 sg13g2_decap_8 FILLER_23_513 ();
 sg13g2_fill_2 FILLER_23_529 ();
 sg13g2_fill_2 FILLER_23_545 ();
 sg13g2_fill_1 FILLER_23_547 ();
 sg13g2_decap_8 FILLER_23_552 ();
 sg13g2_decap_8 FILLER_23_559 ();
 sg13g2_decap_4 FILLER_23_566 ();
 sg13g2_decap_4 FILLER_23_574 ();
 sg13g2_fill_2 FILLER_23_586 ();
 sg13g2_fill_1 FILLER_23_608 ();
 sg13g2_decap_8 FILLER_23_619 ();
 sg13g2_decap_8 FILLER_23_626 ();
 sg13g2_decap_8 FILLER_23_633 ();
 sg13g2_fill_1 FILLER_23_640 ();
 sg13g2_decap_4 FILLER_23_645 ();
 sg13g2_fill_1 FILLER_23_649 ();
 sg13g2_decap_4 FILLER_23_654 ();
 sg13g2_fill_1 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_664 ();
 sg13g2_decap_8 FILLER_23_671 ();
 sg13g2_fill_2 FILLER_23_678 ();
 sg13g2_fill_1 FILLER_23_680 ();
 sg13g2_decap_8 FILLER_23_689 ();
 sg13g2_decap_8 FILLER_23_696 ();
 sg13g2_decap_8 FILLER_23_703 ();
 sg13g2_decap_8 FILLER_23_710 ();
 sg13g2_decap_8 FILLER_23_717 ();
 sg13g2_decap_4 FILLER_23_724 ();
 sg13g2_decap_8 FILLER_23_732 ();
 sg13g2_decap_8 FILLER_23_739 ();
 sg13g2_decap_8 FILLER_23_746 ();
 sg13g2_decap_4 FILLER_23_753 ();
 sg13g2_fill_1 FILLER_23_757 ();
 sg13g2_fill_2 FILLER_23_770 ();
 sg13g2_fill_1 FILLER_23_772 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_decap_8 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_fill_2 FILLER_23_875 ();
 sg13g2_fill_1 FILLER_23_877 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_fill_2 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_65 ();
 sg13g2_fill_1 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_75 ();
 sg13g2_decap_8 FILLER_24_82 ();
 sg13g2_decap_8 FILLER_24_89 ();
 sg13g2_decap_4 FILLER_24_96 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_decap_8 FILLER_24_106 ();
 sg13g2_decap_8 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_120 ();
 sg13g2_decap_8 FILLER_24_127 ();
 sg13g2_decap_8 FILLER_24_134 ();
 sg13g2_fill_2 FILLER_24_141 ();
 sg13g2_fill_1 FILLER_24_143 ();
 sg13g2_decap_4 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_153 ();
 sg13g2_decap_4 FILLER_24_160 ();
 sg13g2_fill_1 FILLER_24_164 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_fill_2 FILLER_24_185 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_229 ();
 sg13g2_decap_4 FILLER_24_247 ();
 sg13g2_fill_2 FILLER_24_251 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_4 FILLER_24_273 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_283 ();
 sg13g2_fill_2 FILLER_24_290 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_decap_4 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_358 ();
 sg13g2_decap_4 FILLER_24_363 ();
 sg13g2_fill_2 FILLER_24_367 ();
 sg13g2_fill_1 FILLER_24_381 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_fill_2 FILLER_24_393 ();
 sg13g2_fill_1 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_decap_8 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_24_415 ();
 sg13g2_fill_1 FILLER_24_422 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_4 FILLER_24_469 ();
 sg13g2_fill_1 FILLER_24_473 ();
 sg13g2_fill_1 FILLER_24_483 ();
 sg13g2_decap_4 FILLER_24_493 ();
 sg13g2_fill_2 FILLER_24_501 ();
 sg13g2_fill_1 FILLER_24_503 ();
 sg13g2_decap_8 FILLER_24_509 ();
 sg13g2_decap_4 FILLER_24_516 ();
 sg13g2_fill_2 FILLER_24_520 ();
 sg13g2_fill_1 FILLER_24_526 ();
 sg13g2_decap_8 FILLER_24_533 ();
 sg13g2_decap_8 FILLER_24_540 ();
 sg13g2_fill_2 FILLER_24_547 ();
 sg13g2_fill_1 FILLER_24_549 ();
 sg13g2_decap_4 FILLER_24_556 ();
 sg13g2_fill_2 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_568 ();
 sg13g2_fill_2 FILLER_24_575 ();
 sg13g2_decap_8 FILLER_24_582 ();
 sg13g2_decap_4 FILLER_24_589 ();
 sg13g2_fill_2 FILLER_24_593 ();
 sg13g2_fill_1 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_615 ();
 sg13g2_decap_8 FILLER_24_622 ();
 sg13g2_decap_8 FILLER_24_629 ();
 sg13g2_decap_4 FILLER_24_636 ();
 sg13g2_fill_2 FILLER_24_640 ();
 sg13g2_fill_1 FILLER_24_653 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_fill_1 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_671 ();
 sg13g2_fill_2 FILLER_24_678 ();
 sg13g2_fill_1 FILLER_24_680 ();
 sg13g2_decap_4 FILLER_24_690 ();
 sg13g2_fill_1 FILLER_24_694 ();
 sg13g2_fill_1 FILLER_24_704 ();
 sg13g2_fill_1 FILLER_24_710 ();
 sg13g2_fill_2 FILLER_24_716 ();
 sg13g2_fill_2 FILLER_24_722 ();
 sg13g2_fill_1 FILLER_24_724 ();
 sg13g2_decap_4 FILLER_24_729 ();
 sg13g2_fill_2 FILLER_24_733 ();
 sg13g2_decap_8 FILLER_24_739 ();
 sg13g2_decap_4 FILLER_24_746 ();
 sg13g2_fill_1 FILLER_24_750 ();
 sg13g2_decap_8 FILLER_24_760 ();
 sg13g2_decap_8 FILLER_24_767 ();
 sg13g2_fill_1 FILLER_24_774 ();
 sg13g2_decap_8 FILLER_24_783 ();
 sg13g2_decap_8 FILLER_24_790 ();
 sg13g2_decap_8 FILLER_24_797 ();
 sg13g2_decap_8 FILLER_24_804 ();
 sg13g2_decap_8 FILLER_24_811 ();
 sg13g2_decap_8 FILLER_24_818 ();
 sg13g2_decap_8 FILLER_24_825 ();
 sg13g2_decap_8 FILLER_24_832 ();
 sg13g2_decap_8 FILLER_24_839 ();
 sg13g2_decap_8 FILLER_24_846 ();
 sg13g2_decap_8 FILLER_24_853 ();
 sg13g2_decap_8 FILLER_24_860 ();
 sg13g2_decap_8 FILLER_24_867 ();
 sg13g2_decap_4 FILLER_24_874 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_4 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_75 ();
 sg13g2_fill_2 FILLER_25_85 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_decap_4 FILLER_25_101 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_154 ();
 sg13g2_fill_2 FILLER_25_159 ();
 sg13g2_decap_8 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_173 ();
 sg13g2_decap_8 FILLER_25_179 ();
 sg13g2_decap_4 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_decap_8 FILLER_25_218 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_decap_8 FILLER_25_239 ();
 sg13g2_decap_4 FILLER_25_246 ();
 sg13g2_fill_1 FILLER_25_250 ();
 sg13g2_decap_4 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_265 ();
 sg13g2_fill_1 FILLER_25_267 ();
 sg13g2_decap_4 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_289 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_4 FILLER_25_329 ();
 sg13g2_fill_2 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_fill_2 FILLER_25_387 ();
 sg13g2_fill_1 FILLER_25_389 ();
 sg13g2_fill_2 FILLER_25_395 ();
 sg13g2_fill_1 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_411 ();
 sg13g2_decap_4 FILLER_25_418 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_fill_1 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_460 ();
 sg13g2_decap_8 FILLER_25_467 ();
 sg13g2_decap_8 FILLER_25_474 ();
 sg13g2_fill_2 FILLER_25_481 ();
 sg13g2_decap_8 FILLER_25_492 ();
 sg13g2_decap_4 FILLER_25_508 ();
 sg13g2_fill_2 FILLER_25_512 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_4 FILLER_25_557 ();
 sg13g2_fill_1 FILLER_25_561 ();
 sg13g2_fill_2 FILLER_25_567 ();
 sg13g2_fill_1 FILLER_25_569 ();
 sg13g2_fill_1 FILLER_25_583 ();
 sg13g2_decap_4 FILLER_25_595 ();
 sg13g2_fill_2 FILLER_25_599 ();
 sg13g2_fill_1 FILLER_25_605 ();
 sg13g2_decap_8 FILLER_25_610 ();
 sg13g2_decap_8 FILLER_25_617 ();
 sg13g2_fill_2 FILLER_25_624 ();
 sg13g2_fill_2 FILLER_25_639 ();
 sg13g2_fill_1 FILLER_25_641 ();
 sg13g2_decap_8 FILLER_25_667 ();
 sg13g2_fill_2 FILLER_25_674 ();
 sg13g2_fill_1 FILLER_25_676 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_decap_4 FILLER_25_690 ();
 sg13g2_fill_1 FILLER_25_694 ();
 sg13g2_decap_8 FILLER_25_711 ();
 sg13g2_decap_4 FILLER_25_718 ();
 sg13g2_fill_1 FILLER_25_732 ();
 sg13g2_decap_8 FILLER_25_739 ();
 sg13g2_decap_8 FILLER_25_746 ();
 sg13g2_decap_4 FILLER_25_753 ();
 sg13g2_decap_4 FILLER_25_762 ();
 sg13g2_decap_4 FILLER_25_771 ();
 sg13g2_fill_1 FILLER_25_775 ();
 sg13g2_decap_8 FILLER_25_781 ();
 sg13g2_decap_8 FILLER_25_788 ();
 sg13g2_decap_8 FILLER_25_795 ();
 sg13g2_decap_8 FILLER_25_802 ();
 sg13g2_decap_8 FILLER_25_809 ();
 sg13g2_decap_8 FILLER_25_816 ();
 sg13g2_decap_8 FILLER_25_823 ();
 sg13g2_decap_8 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_8 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_25_865 ();
 sg13g2_decap_4 FILLER_25_872 ();
 sg13g2_fill_2 FILLER_25_876 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_4 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_80 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_119 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_4 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_164 ();
 sg13g2_decap_8 FILLER_26_171 ();
 sg13g2_decap_8 FILLER_26_178 ();
 sg13g2_decap_8 FILLER_26_185 ();
 sg13g2_decap_4 FILLER_26_192 ();
 sg13g2_fill_2 FILLER_26_200 ();
 sg13g2_decap_4 FILLER_26_206 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_227 ();
 sg13g2_decap_4 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_decap_8 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_decap_4 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_271 ();
 sg13g2_decap_4 FILLER_26_276 ();
 sg13g2_decap_4 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_decap_8 FILLER_26_295 ();
 sg13g2_decap_8 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_321 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_fill_2 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_fill_1 FILLER_26_349 ();
 sg13g2_decap_4 FILLER_26_360 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_1 FILLER_26_369 ();
 sg13g2_fill_2 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_fill_2 FILLER_26_403 ();
 sg13g2_decap_4 FILLER_26_412 ();
 sg13g2_fill_1 FILLER_26_416 ();
 sg13g2_fill_1 FILLER_26_421 ();
 sg13g2_decap_8 FILLER_26_426 ();
 sg13g2_decap_4 FILLER_26_433 ();
 sg13g2_fill_1 FILLER_26_437 ();
 sg13g2_decap_4 FILLER_26_442 ();
 sg13g2_fill_2 FILLER_26_446 ();
 sg13g2_decap_8 FILLER_26_472 ();
 sg13g2_decap_8 FILLER_26_479 ();
 sg13g2_decap_8 FILLER_26_486 ();
 sg13g2_decap_4 FILLER_26_493 ();
 sg13g2_fill_2 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_fill_1 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_520 ();
 sg13g2_decap_4 FILLER_26_527 ();
 sg13g2_decap_8 FILLER_26_536 ();
 sg13g2_decap_8 FILLER_26_547 ();
 sg13g2_fill_1 FILLER_26_554 ();
 sg13g2_fill_1 FILLER_26_559 ();
 sg13g2_decap_8 FILLER_26_566 ();
 sg13g2_decap_4 FILLER_26_573 ();
 sg13g2_fill_1 FILLER_26_577 ();
 sg13g2_fill_2 FILLER_26_582 ();
 sg13g2_fill_1 FILLER_26_584 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_4 FILLER_26_602 ();
 sg13g2_fill_2 FILLER_26_606 ();
 sg13g2_decap_8 FILLER_26_612 ();
 sg13g2_decap_8 FILLER_26_619 ();
 sg13g2_decap_8 FILLER_26_626 ();
 sg13g2_fill_1 FILLER_26_633 ();
 sg13g2_decap_4 FILLER_26_638 ();
 sg13g2_fill_2 FILLER_26_642 ();
 sg13g2_decap_4 FILLER_26_648 ();
 sg13g2_fill_1 FILLER_26_652 ();
 sg13g2_decap_4 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_667 ();
 sg13g2_decap_8 FILLER_26_674 ();
 sg13g2_decap_4 FILLER_26_681 ();
 sg13g2_fill_1 FILLER_26_685 ();
 sg13g2_decap_8 FILLER_26_690 ();
 sg13g2_decap_8 FILLER_26_697 ();
 sg13g2_decap_8 FILLER_26_704 ();
 sg13g2_decap_4 FILLER_26_711 ();
 sg13g2_fill_1 FILLER_26_715 ();
 sg13g2_decap_8 FILLER_26_727 ();
 sg13g2_decap_8 FILLER_26_734 ();
 sg13g2_fill_1 FILLER_26_741 ();
 sg13g2_decap_8 FILLER_26_746 ();
 sg13g2_fill_1 FILLER_26_753 ();
 sg13g2_decap_8 FILLER_26_758 ();
 sg13g2_fill_2 FILLER_26_765 ();
 sg13g2_decap_8 FILLER_26_771 ();
 sg13g2_decap_8 FILLER_26_778 ();
 sg13g2_decap_8 FILLER_26_785 ();
 sg13g2_decap_8 FILLER_26_792 ();
 sg13g2_decap_8 FILLER_26_799 ();
 sg13g2_decap_8 FILLER_26_806 ();
 sg13g2_decap_8 FILLER_26_813 ();
 sg13g2_decap_8 FILLER_26_820 ();
 sg13g2_decap_8 FILLER_26_827 ();
 sg13g2_decap_8 FILLER_26_834 ();
 sg13g2_decap_8 FILLER_26_841 ();
 sg13g2_decap_8 FILLER_26_848 ();
 sg13g2_decap_8 FILLER_26_855 ();
 sg13g2_decap_8 FILLER_26_862 ();
 sg13g2_decap_8 FILLER_26_869 ();
 sg13g2_fill_2 FILLER_26_876 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_64 ();
 sg13g2_decap_8 FILLER_27_71 ();
 sg13g2_fill_1 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_97 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_fill_2 FILLER_27_110 ();
 sg13g2_fill_2 FILLER_27_121 ();
 sg13g2_decap_4 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_decap_4 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_150 ();
 sg13g2_decap_4 FILLER_27_155 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_fill_1 FILLER_27_170 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_191 ();
 sg13g2_fill_2 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_206 ();
 sg13g2_decap_8 FILLER_27_213 ();
 sg13g2_decap_8 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_decap_8 FILLER_27_232 ();
 sg13g2_fill_2 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_241 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_4 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_decap_8 FILLER_27_296 ();
 sg13g2_decap_4 FILLER_27_307 ();
 sg13g2_fill_2 FILLER_27_311 ();
 sg13g2_decap_8 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_323 ();
 sg13g2_decap_4 FILLER_27_330 ();
 sg13g2_fill_2 FILLER_27_334 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_fill_2 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_407 ();
 sg13g2_fill_2 FILLER_27_414 ();
 sg13g2_fill_1 FILLER_27_421 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_decap_8 FILLER_27_436 ();
 sg13g2_decap_4 FILLER_27_443 ();
 sg13g2_fill_1 FILLER_27_447 ();
 sg13g2_decap_8 FILLER_27_458 ();
 sg13g2_decap_8 FILLER_27_465 ();
 sg13g2_fill_2 FILLER_27_472 ();
 sg13g2_decap_8 FILLER_27_478 ();
 sg13g2_decap_8 FILLER_27_485 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_fill_1 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_516 ();
 sg13g2_fill_2 FILLER_27_523 ();
 sg13g2_decap_8 FILLER_27_529 ();
 sg13g2_decap_8 FILLER_27_536 ();
 sg13g2_decap_8 FILLER_27_543 ();
 sg13g2_fill_1 FILLER_27_550 ();
 sg13g2_fill_1 FILLER_27_560 ();
 sg13g2_decap_4 FILLER_27_565 ();
 sg13g2_fill_2 FILLER_27_581 ();
 sg13g2_fill_2 FILLER_27_592 ();
 sg13g2_fill_1 FILLER_27_594 ();
 sg13g2_fill_2 FILLER_27_600 ();
 sg13g2_fill_1 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_613 ();
 sg13g2_decap_8 FILLER_27_620 ();
 sg13g2_decap_8 FILLER_27_627 ();
 sg13g2_decap_8 FILLER_27_634 ();
 sg13g2_decap_8 FILLER_27_641 ();
 sg13g2_decap_8 FILLER_27_648 ();
 sg13g2_decap_4 FILLER_27_655 ();
 sg13g2_fill_2 FILLER_27_659 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_fill_2 FILLER_27_672 ();
 sg13g2_fill_1 FILLER_27_674 ();
 sg13g2_decap_8 FILLER_27_683 ();
 sg13g2_fill_2 FILLER_27_690 ();
 sg13g2_decap_8 FILLER_27_697 ();
 sg13g2_decap_4 FILLER_27_713 ();
 sg13g2_fill_1 FILLER_27_717 ();
 sg13g2_decap_8 FILLER_27_722 ();
 sg13g2_decap_8 FILLER_27_729 ();
 sg13g2_decap_4 FILLER_27_736 ();
 sg13g2_fill_1 FILLER_27_740 ();
 sg13g2_decap_8 FILLER_27_754 ();
 sg13g2_decap_8 FILLER_27_761 ();
 sg13g2_decap_4 FILLER_27_768 ();
 sg13g2_fill_1 FILLER_27_772 ();
 sg13g2_fill_1 FILLER_27_781 ();
 sg13g2_decap_8 FILLER_27_786 ();
 sg13g2_decap_8 FILLER_27_793 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_8 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_fill_1 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_4 FILLER_28_63 ();
 sg13g2_decap_4 FILLER_28_75 ();
 sg13g2_fill_2 FILLER_28_79 ();
 sg13g2_decap_8 FILLER_28_86 ();
 sg13g2_decap_8 FILLER_28_93 ();
 sg13g2_decap_8 FILLER_28_100 ();
 sg13g2_decap_8 FILLER_28_107 ();
 sg13g2_decap_8 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_121 ();
 sg13g2_decap_8 FILLER_28_128 ();
 sg13g2_decap_8 FILLER_28_135 ();
 sg13g2_fill_1 FILLER_28_142 ();
 sg13g2_decap_8 FILLER_28_151 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_decap_8 FILLER_28_169 ();
 sg13g2_decap_4 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_decap_8 FILLER_28_204 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_fill_2 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_decap_8 FILLER_28_226 ();
 sg13g2_fill_1 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_245 ();
 sg13g2_fill_1 FILLER_28_254 ();
 sg13g2_decap_8 FILLER_28_260 ();
 sg13g2_decap_8 FILLER_28_267 ();
 sg13g2_decap_8 FILLER_28_274 ();
 sg13g2_fill_2 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_298 ();
 sg13g2_decap_4 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_fill_2 FILLER_28_392 ();
 sg13g2_fill_1 FILLER_28_394 ();
 sg13g2_decap_4 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_414 ();
 sg13g2_decap_8 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_445 ();
 sg13g2_decap_4 FILLER_28_451 ();
 sg13g2_fill_2 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_468 ();
 sg13g2_fill_1 FILLER_28_475 ();
 sg13g2_decap_8 FILLER_28_482 ();
 sg13g2_decap_4 FILLER_28_489 ();
 sg13g2_decap_4 FILLER_28_497 ();
 sg13g2_fill_2 FILLER_28_501 ();
 sg13g2_decap_8 FILLER_28_507 ();
 sg13g2_decap_8 FILLER_28_531 ();
 sg13g2_decap_8 FILLER_28_538 ();
 sg13g2_decap_8 FILLER_28_545 ();
 sg13g2_fill_2 FILLER_28_552 ();
 sg13g2_fill_1 FILLER_28_558 ();
 sg13g2_fill_1 FILLER_28_568 ();
 sg13g2_fill_1 FILLER_28_573 ();
 sg13g2_fill_1 FILLER_28_580 ();
 sg13g2_fill_1 FILLER_28_592 ();
 sg13g2_decap_8 FILLER_28_606 ();
 sg13g2_decap_8 FILLER_28_613 ();
 sg13g2_decap_8 FILLER_28_620 ();
 sg13g2_decap_8 FILLER_28_627 ();
 sg13g2_decap_8 FILLER_28_634 ();
 sg13g2_decap_8 FILLER_28_641 ();
 sg13g2_decap_8 FILLER_28_648 ();
 sg13g2_decap_8 FILLER_28_669 ();
 sg13g2_fill_1 FILLER_28_676 ();
 sg13g2_fill_1 FILLER_28_682 ();
 sg13g2_fill_1 FILLER_28_688 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_4 FILLER_28_714 ();
 sg13g2_fill_1 FILLER_28_718 ();
 sg13g2_decap_8 FILLER_28_723 ();
 sg13g2_decap_8 FILLER_28_730 ();
 sg13g2_decap_8 FILLER_28_741 ();
 sg13g2_decap_4 FILLER_28_748 ();
 sg13g2_decap_4 FILLER_28_764 ();
 sg13g2_fill_2 FILLER_28_768 ();
 sg13g2_decap_8 FILLER_28_782 ();
 sg13g2_decap_8 FILLER_28_789 ();
 sg13g2_decap_8 FILLER_28_796 ();
 sg13g2_decap_8 FILLER_28_803 ();
 sg13g2_decap_8 FILLER_28_810 ();
 sg13g2_decap_8 FILLER_28_817 ();
 sg13g2_decap_8 FILLER_28_824 ();
 sg13g2_decap_8 FILLER_28_831 ();
 sg13g2_decap_8 FILLER_28_838 ();
 sg13g2_decap_8 FILLER_28_845 ();
 sg13g2_decap_8 FILLER_28_852 ();
 sg13g2_decap_8 FILLER_28_859 ();
 sg13g2_decap_8 FILLER_28_866 ();
 sg13g2_decap_4 FILLER_28_873 ();
 sg13g2_fill_1 FILLER_28_877 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_75 ();
 sg13g2_fill_1 FILLER_29_77 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_decap_8 FILLER_29_89 ();
 sg13g2_decap_8 FILLER_29_96 ();
 sg13g2_fill_2 FILLER_29_103 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_125 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_decap_4 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_153 ();
 sg13g2_fill_1 FILLER_29_155 ();
 sg13g2_decap_8 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_184 ();
 sg13g2_decap_4 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_212 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_fill_2 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_decap_8 FILLER_29_246 ();
 sg13g2_decap_8 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_260 ();
 sg13g2_fill_1 FILLER_29_262 ();
 sg13g2_fill_2 FILLER_29_274 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_4 FILLER_29_287 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_decap_4 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_4 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_decap_4 FILLER_29_332 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_4 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_4 FILLER_29_371 ();
 sg13g2_fill_1 FILLER_29_375 ();
 sg13g2_fill_2 FILLER_29_381 ();
 sg13g2_fill_2 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_390 ();
 sg13g2_decap_4 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_411 ();
 sg13g2_decap_8 FILLER_29_418 ();
 sg13g2_decap_8 FILLER_29_425 ();
 sg13g2_decap_8 FILLER_29_432 ();
 sg13g2_decap_8 FILLER_29_439 ();
 sg13g2_fill_2 FILLER_29_446 ();
 sg13g2_decap_4 FILLER_29_453 ();
 sg13g2_fill_1 FILLER_29_457 ();
 sg13g2_decap_8 FILLER_29_473 ();
 sg13g2_fill_1 FILLER_29_480 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_fill_1 FILLER_29_518 ();
 sg13g2_fill_1 FILLER_29_524 ();
 sg13g2_decap_8 FILLER_29_535 ();
 sg13g2_fill_2 FILLER_29_542 ();
 sg13g2_fill_1 FILLER_29_544 ();
 sg13g2_fill_1 FILLER_29_550 ();
 sg13g2_fill_2 FILLER_29_557 ();
 sg13g2_decap_4 FILLER_29_563 ();
 sg13g2_fill_2 FILLER_29_567 ();
 sg13g2_fill_2 FILLER_29_573 ();
 sg13g2_fill_1 FILLER_29_575 ();
 sg13g2_decap_8 FILLER_29_585 ();
 sg13g2_decap_8 FILLER_29_592 ();
 sg13g2_decap_8 FILLER_29_599 ();
 sg13g2_fill_1 FILLER_29_606 ();
 sg13g2_fill_2 FILLER_29_632 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_4 FILLER_29_655 ();
 sg13g2_decap_8 FILLER_29_671 ();
 sg13g2_decap_8 FILLER_29_678 ();
 sg13g2_decap_4 FILLER_29_685 ();
 sg13g2_fill_2 FILLER_29_689 ();
 sg13g2_fill_1 FILLER_29_696 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_fill_1 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_712 ();
 sg13g2_fill_1 FILLER_29_719 ();
 sg13g2_decap_8 FILLER_29_726 ();
 sg13g2_fill_1 FILLER_29_733 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_fill_2 FILLER_29_763 ();
 sg13g2_decap_4 FILLER_29_769 ();
 sg13g2_fill_2 FILLER_29_773 ();
 sg13g2_decap_8 FILLER_29_780 ();
 sg13g2_decap_8 FILLER_29_787 ();
 sg13g2_decap_8 FILLER_29_794 ();
 sg13g2_decap_8 FILLER_29_801 ();
 sg13g2_decap_8 FILLER_29_808 ();
 sg13g2_decap_8 FILLER_29_815 ();
 sg13g2_decap_8 FILLER_29_822 ();
 sg13g2_decap_8 FILLER_29_829 ();
 sg13g2_decap_8 FILLER_29_836 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_decap_8 FILLER_29_850 ();
 sg13g2_decap_8 FILLER_29_857 ();
 sg13g2_decap_8 FILLER_29_864 ();
 sg13g2_decap_8 FILLER_29_871 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_58 ();
 sg13g2_fill_2 FILLER_30_64 ();
 sg13g2_fill_1 FILLER_30_66 ();
 sg13g2_decap_8 FILLER_30_72 ();
 sg13g2_decap_8 FILLER_30_79 ();
 sg13g2_decap_4 FILLER_30_86 ();
 sg13g2_fill_2 FILLER_30_90 ();
 sg13g2_decap_4 FILLER_30_96 ();
 sg13g2_fill_1 FILLER_30_100 ();
 sg13g2_fill_2 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_115 ();
 sg13g2_decap_4 FILLER_30_127 ();
 sg13g2_decap_8 FILLER_30_136 ();
 sg13g2_decap_4 FILLER_30_143 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_decap_8 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_212 ();
 sg13g2_fill_1 FILLER_30_214 ();
 sg13g2_fill_1 FILLER_30_224 ();
 sg13g2_fill_2 FILLER_30_229 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_251 ();
 sg13g2_decap_8 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_fill_1 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_317 ();
 sg13g2_decap_4 FILLER_30_324 ();
 sg13g2_decap_8 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_345 ();
 sg13g2_decap_8 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_fill_1 FILLER_30_373 ();
 sg13g2_decap_4 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_30_409 ();
 sg13g2_decap_4 FILLER_30_416 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_30_433 ();
 sg13g2_decap_4 FILLER_30_440 ();
 sg13g2_fill_1 FILLER_30_444 ();
 sg13g2_decap_4 FILLER_30_449 ();
 sg13g2_decap_8 FILLER_30_457 ();
 sg13g2_decap_4 FILLER_30_464 ();
 sg13g2_fill_1 FILLER_30_468 ();
 sg13g2_decap_8 FILLER_30_474 ();
 sg13g2_decap_8 FILLER_30_481 ();
 sg13g2_decap_8 FILLER_30_488 ();
 sg13g2_decap_8 FILLER_30_500 ();
 sg13g2_decap_8 FILLER_30_507 ();
 sg13g2_fill_2 FILLER_30_514 ();
 sg13g2_decap_8 FILLER_30_529 ();
 sg13g2_decap_8 FILLER_30_536 ();
 sg13g2_decap_8 FILLER_30_543 ();
 sg13g2_decap_4 FILLER_30_554 ();
 sg13g2_fill_2 FILLER_30_558 ();
 sg13g2_decap_8 FILLER_30_565 ();
 sg13g2_decap_8 FILLER_30_572 ();
 sg13g2_decap_4 FILLER_30_579 ();
 sg13g2_fill_1 FILLER_30_583 ();
 sg13g2_fill_2 FILLER_30_588 ();
 sg13g2_fill_1 FILLER_30_590 ();
 sg13g2_decap_8 FILLER_30_606 ();
 sg13g2_fill_1 FILLER_30_613 ();
 sg13g2_decap_8 FILLER_30_627 ();
 sg13g2_decap_8 FILLER_30_634 ();
 sg13g2_decap_4 FILLER_30_641 ();
 sg13g2_fill_1 FILLER_30_645 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_4 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_666 ();
 sg13g2_decap_8 FILLER_30_673 ();
 sg13g2_decap_8 FILLER_30_680 ();
 sg13g2_decap_4 FILLER_30_687 ();
 sg13g2_decap_8 FILLER_30_695 ();
 sg13g2_decap_8 FILLER_30_706 ();
 sg13g2_fill_2 FILLER_30_713 ();
 sg13g2_fill_1 FILLER_30_715 ();
 sg13g2_fill_1 FILLER_30_720 ();
 sg13g2_decap_8 FILLER_30_725 ();
 sg13g2_decap_4 FILLER_30_732 ();
 sg13g2_decap_8 FILLER_30_740 ();
 sg13g2_fill_2 FILLER_30_747 ();
 sg13g2_fill_1 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_decap_8 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_30_868 ();
 sg13g2_fill_2 FILLER_30_875 ();
 sg13g2_fill_1 FILLER_30_877 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_4 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_75 ();
 sg13g2_decap_4 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_86 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_111 ();
 sg13g2_decap_8 FILLER_31_138 ();
 sg13g2_decap_8 FILLER_31_145 ();
 sg13g2_decap_8 FILLER_31_152 ();
 sg13g2_fill_1 FILLER_31_159 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_194 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_decap_8 FILLER_31_214 ();
 sg13g2_fill_2 FILLER_31_221 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_decap_4 FILLER_31_249 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_decap_4 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_decap_8 FILLER_31_267 ();
 sg13g2_decap_8 FILLER_31_274 ();
 sg13g2_decap_8 FILLER_31_281 ();
 sg13g2_decap_8 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_318 ();
 sg13g2_decap_8 FILLER_31_325 ();
 sg13g2_fill_2 FILLER_31_332 ();
 sg13g2_decap_4 FILLER_31_341 ();
 sg13g2_fill_2 FILLER_31_345 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_384 ();
 sg13g2_fill_2 FILLER_31_391 ();
 sg13g2_fill_1 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_fill_2 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_426 ();
 sg13g2_decap_4 FILLER_31_433 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_fill_1 FILLER_31_469 ();
 sg13g2_fill_2 FILLER_31_474 ();
 sg13g2_fill_2 FILLER_31_497 ();
 sg13g2_fill_1 FILLER_31_508 ();
 sg13g2_fill_2 FILLER_31_514 ();
 sg13g2_fill_1 FILLER_31_516 ();
 sg13g2_fill_2 FILLER_31_521 ();
 sg13g2_fill_1 FILLER_31_523 ();
 sg13g2_decap_4 FILLER_31_536 ();
 sg13g2_fill_1 FILLER_31_545 ();
 sg13g2_decap_8 FILLER_31_556 ();
 sg13g2_decap_4 FILLER_31_563 ();
 sg13g2_fill_2 FILLER_31_567 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_decap_4 FILLER_31_586 ();
 sg13g2_fill_1 FILLER_31_590 ();
 sg13g2_fill_1 FILLER_31_596 ();
 sg13g2_fill_2 FILLER_31_601 ();
 sg13g2_decap_8 FILLER_31_608 ();
 sg13g2_decap_8 FILLER_31_615 ();
 sg13g2_decap_4 FILLER_31_622 ();
 sg13g2_fill_2 FILLER_31_626 ();
 sg13g2_decap_4 FILLER_31_632 ();
 sg13g2_fill_2 FILLER_31_636 ();
 sg13g2_fill_2 FILLER_31_647 ();
 sg13g2_decap_8 FILLER_31_653 ();
 sg13g2_decap_8 FILLER_31_660 ();
 sg13g2_decap_8 FILLER_31_667 ();
 sg13g2_decap_4 FILLER_31_674 ();
 sg13g2_decap_8 FILLER_31_684 ();
 sg13g2_decap_8 FILLER_31_691 ();
 sg13g2_decap_4 FILLER_31_698 ();
 sg13g2_decap_8 FILLER_31_706 ();
 sg13g2_decap_8 FILLER_31_713 ();
 sg13g2_fill_1 FILLER_31_720 ();
 sg13g2_decap_8 FILLER_31_725 ();
 sg13g2_decap_8 FILLER_31_732 ();
 sg13g2_decap_8 FILLER_31_739 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_decap_8 FILLER_31_757 ();
 sg13g2_decap_8 FILLER_31_764 ();
 sg13g2_decap_4 FILLER_31_771 ();
 sg13g2_fill_1 FILLER_31_775 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_decap_8 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_31_868 ();
 sg13g2_fill_2 FILLER_31_875 ();
 sg13g2_fill_1 FILLER_31_877 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_58 ();
 sg13g2_fill_2 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_93 ();
 sg13g2_decap_8 FILLER_32_100 ();
 sg13g2_decap_8 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_114 ();
 sg13g2_decap_8 FILLER_32_120 ();
 sg13g2_decap_8 FILLER_32_127 ();
 sg13g2_decap_4 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_fill_2 FILLER_32_159 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_2 FILLER_32_190 ();
 sg13g2_decap_4 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_decap_4 FILLER_32_216 ();
 sg13g2_fill_1 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_decap_8 FILLER_32_246 ();
 sg13g2_decap_8 FILLER_32_253 ();
 sg13g2_fill_1 FILLER_32_260 ();
 sg13g2_fill_2 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_fill_2 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_4 FILLER_32_301 ();
 sg13g2_decap_4 FILLER_32_309 ();
 sg13g2_decap_8 FILLER_32_317 ();
 sg13g2_decap_8 FILLER_32_324 ();
 sg13g2_decap_4 FILLER_32_331 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_fill_2 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_4 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_373 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_decap_8 FILLER_32_393 ();
 sg13g2_decap_8 FILLER_32_400 ();
 sg13g2_decap_8 FILLER_32_407 ();
 sg13g2_decap_8 FILLER_32_414 ();
 sg13g2_decap_8 FILLER_32_421 ();
 sg13g2_decap_4 FILLER_32_428 ();
 sg13g2_fill_2 FILLER_32_432 ();
 sg13g2_fill_1 FILLER_32_447 ();
 sg13g2_decap_8 FILLER_32_452 ();
 sg13g2_decap_8 FILLER_32_459 ();
 sg13g2_decap_4 FILLER_32_466 ();
 sg13g2_fill_2 FILLER_32_475 ();
 sg13g2_fill_1 FILLER_32_477 ();
 sg13g2_decap_8 FILLER_32_486 ();
 sg13g2_decap_4 FILLER_32_493 ();
 sg13g2_fill_2 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_503 ();
 sg13g2_decap_8 FILLER_32_510 ();
 sg13g2_decap_8 FILLER_32_517 ();
 sg13g2_decap_8 FILLER_32_524 ();
 sg13g2_decap_8 FILLER_32_531 ();
 sg13g2_decap_8 FILLER_32_538 ();
 sg13g2_decap_8 FILLER_32_545 ();
 sg13g2_fill_2 FILLER_32_552 ();
 sg13g2_decap_8 FILLER_32_566 ();
 sg13g2_decap_8 FILLER_32_573 ();
 sg13g2_decap_8 FILLER_32_580 ();
 sg13g2_decap_8 FILLER_32_587 ();
 sg13g2_decap_4 FILLER_32_594 ();
 sg13g2_fill_1 FILLER_32_598 ();
 sg13g2_decap_8 FILLER_32_609 ();
 sg13g2_fill_2 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_622 ();
 sg13g2_decap_8 FILLER_32_629 ();
 sg13g2_fill_2 FILLER_32_636 ();
 sg13g2_fill_2 FILLER_32_646 ();
 sg13g2_decap_8 FILLER_32_652 ();
 sg13g2_fill_1 FILLER_32_659 ();
 sg13g2_decap_8 FILLER_32_663 ();
 sg13g2_decap_8 FILLER_32_670 ();
 sg13g2_decap_8 FILLER_32_677 ();
 sg13g2_decap_8 FILLER_32_688 ();
 sg13g2_decap_8 FILLER_32_695 ();
 sg13g2_decap_4 FILLER_32_702 ();
 sg13g2_fill_1 FILLER_32_711 ();
 sg13g2_decap_8 FILLER_32_719 ();
 sg13g2_decap_8 FILLER_32_726 ();
 sg13g2_decap_4 FILLER_32_733 ();
 sg13g2_fill_1 FILLER_32_741 ();
 sg13g2_decap_8 FILLER_32_751 ();
 sg13g2_fill_2 FILLER_32_764 ();
 sg13g2_fill_1 FILLER_32_766 ();
 sg13g2_decap_8 FILLER_32_780 ();
 sg13g2_decap_8 FILLER_32_787 ();
 sg13g2_decap_8 FILLER_32_794 ();
 sg13g2_decap_8 FILLER_32_801 ();
 sg13g2_decap_8 FILLER_32_808 ();
 sg13g2_decap_8 FILLER_32_815 ();
 sg13g2_decap_8 FILLER_32_822 ();
 sg13g2_decap_8 FILLER_32_829 ();
 sg13g2_decap_8 FILLER_32_836 ();
 sg13g2_decap_8 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_850 ();
 sg13g2_decap_8 FILLER_32_857 ();
 sg13g2_decap_8 FILLER_32_864 ();
 sg13g2_decap_8 FILLER_32_871 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_68 ();
 sg13g2_fill_1 FILLER_33_78 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_4 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_116 ();
 sg13g2_decap_8 FILLER_33_127 ();
 sg13g2_decap_8 FILLER_33_134 ();
 sg13g2_decap_8 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_148 ();
 sg13g2_fill_2 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_decap_8 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_187 ();
 sg13g2_decap_8 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_4 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_224 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_decap_8 FILLER_33_267 ();
 sg13g2_decap_8 FILLER_33_274 ();
 sg13g2_decap_8 FILLER_33_281 ();
 sg13g2_decap_8 FILLER_33_288 ();
 sg13g2_decap_8 FILLER_33_295 ();
 sg13g2_decap_4 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_311 ();
 sg13g2_decap_8 FILLER_33_318 ();
 sg13g2_decap_8 FILLER_33_325 ();
 sg13g2_decap_4 FILLER_33_348 ();
 sg13g2_fill_1 FILLER_33_381 ();
 sg13g2_decap_4 FILLER_33_392 ();
 sg13g2_fill_2 FILLER_33_396 ();
 sg13g2_decap_8 FILLER_33_404 ();
 sg13g2_fill_2 FILLER_33_418 ();
 sg13g2_decap_8 FILLER_33_424 ();
 sg13g2_fill_2 FILLER_33_431 ();
 sg13g2_fill_2 FILLER_33_450 ();
 sg13g2_fill_1 FILLER_33_452 ();
 sg13g2_decap_8 FILLER_33_457 ();
 sg13g2_decap_8 FILLER_33_464 ();
 sg13g2_decap_8 FILLER_33_471 ();
 sg13g2_decap_8 FILLER_33_478 ();
 sg13g2_decap_8 FILLER_33_485 ();
 sg13g2_decap_8 FILLER_33_492 ();
 sg13g2_decap_8 FILLER_33_499 ();
 sg13g2_fill_1 FILLER_33_506 ();
 sg13g2_decap_8 FILLER_33_512 ();
 sg13g2_fill_2 FILLER_33_519 ();
 sg13g2_fill_1 FILLER_33_521 ();
 sg13g2_decap_8 FILLER_33_528 ();
 sg13g2_decap_8 FILLER_33_535 ();
 sg13g2_decap_8 FILLER_33_542 ();
 sg13g2_fill_2 FILLER_33_549 ();
 sg13g2_fill_1 FILLER_33_551 ();
 sg13g2_fill_1 FILLER_33_565 ();
 sg13g2_decap_8 FILLER_33_570 ();
 sg13g2_decap_8 FILLER_33_577 ();
 sg13g2_decap_8 FILLER_33_584 ();
 sg13g2_decap_8 FILLER_33_591 ();
 sg13g2_decap_4 FILLER_33_598 ();
 sg13g2_fill_1 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_613 ();
 sg13g2_fill_1 FILLER_33_624 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_fill_1 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_4 FILLER_33_700 ();
 sg13g2_fill_2 FILLER_33_704 ();
 sg13g2_decap_8 FILLER_33_710 ();
 sg13g2_fill_2 FILLER_33_722 ();
 sg13g2_fill_2 FILLER_33_729 ();
 sg13g2_fill_2 FILLER_33_746 ();
 sg13g2_fill_1 FILLER_33_748 ();
 sg13g2_decap_8 FILLER_33_753 ();
 sg13g2_decap_8 FILLER_33_760 ();
 sg13g2_decap_8 FILLER_33_767 ();
 sg13g2_decap_8 FILLER_33_774 ();
 sg13g2_decap_8 FILLER_33_781 ();
 sg13g2_decap_8 FILLER_33_788 ();
 sg13g2_decap_8 FILLER_33_795 ();
 sg13g2_decap_8 FILLER_33_802 ();
 sg13g2_decap_8 FILLER_33_809 ();
 sg13g2_decap_8 FILLER_33_816 ();
 sg13g2_decap_8 FILLER_33_823 ();
 sg13g2_decap_8 FILLER_33_830 ();
 sg13g2_decap_8 FILLER_33_837 ();
 sg13g2_decap_8 FILLER_33_844 ();
 sg13g2_decap_8 FILLER_33_851 ();
 sg13g2_decap_8 FILLER_33_858 ();
 sg13g2_decap_8 FILLER_33_865 ();
 sg13g2_decap_4 FILLER_33_872 ();
 sg13g2_fill_2 FILLER_33_876 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_72 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_fill_2 FILLER_34_154 ();
 sg13g2_decap_4 FILLER_34_161 ();
 sg13g2_fill_2 FILLER_34_169 ();
 sg13g2_fill_1 FILLER_34_171 ();
 sg13g2_decap_8 FILLER_34_177 ();
 sg13g2_fill_1 FILLER_34_184 ();
 sg13g2_decap_8 FILLER_34_190 ();
 sg13g2_fill_2 FILLER_34_197 ();
 sg13g2_fill_1 FILLER_34_199 ();
 sg13g2_decap_8 FILLER_34_204 ();
 sg13g2_decap_8 FILLER_34_211 ();
 sg13g2_decap_8 FILLER_34_218 ();
 sg13g2_decap_8 FILLER_34_225 ();
 sg13g2_fill_2 FILLER_34_232 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_fill_2 FILLER_34_265 ();
 sg13g2_fill_1 FILLER_34_267 ();
 sg13g2_decap_8 FILLER_34_271 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_decap_8 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_307 ();
 sg13g2_decap_4 FILLER_34_314 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_decap_8 FILLER_34_323 ();
 sg13g2_decap_4 FILLER_34_330 ();
 sg13g2_fill_2 FILLER_34_334 ();
 sg13g2_decap_4 FILLER_34_340 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_decap_4 FILLER_34_386 ();
 sg13g2_fill_1 FILLER_34_390 ();
 sg13g2_decap_4 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_417 ();
 sg13g2_decap_8 FILLER_34_424 ();
 sg13g2_decap_8 FILLER_34_431 ();
 sg13g2_fill_2 FILLER_34_438 ();
 sg13g2_decap_8 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_455 ();
 sg13g2_decap_8 FILLER_34_462 ();
 sg13g2_fill_2 FILLER_34_469 ();
 sg13g2_fill_1 FILLER_34_471 ();
 sg13g2_decap_8 FILLER_34_487 ();
 sg13g2_decap_8 FILLER_34_494 ();
 sg13g2_decap_4 FILLER_34_510 ();
 sg13g2_fill_1 FILLER_34_514 ();
 sg13g2_decap_8 FILLER_34_520 ();
 sg13g2_decap_8 FILLER_34_527 ();
 sg13g2_decap_4 FILLER_34_534 ();
 sg13g2_fill_1 FILLER_34_538 ();
 sg13g2_decap_8 FILLER_34_543 ();
 sg13g2_decap_8 FILLER_34_550 ();
 sg13g2_fill_1 FILLER_34_557 ();
 sg13g2_fill_2 FILLER_34_563 ();
 sg13g2_fill_2 FILLER_34_568 ();
 sg13g2_fill_1 FILLER_34_570 ();
 sg13g2_fill_1 FILLER_34_587 ();
 sg13g2_decap_4 FILLER_34_592 ();
 sg13g2_fill_1 FILLER_34_600 ();
 sg13g2_fill_1 FILLER_34_606 ();
 sg13g2_fill_1 FILLER_34_611 ();
 sg13g2_fill_2 FILLER_34_617 ();
 sg13g2_decap_8 FILLER_34_638 ();
 sg13g2_decap_8 FILLER_34_645 ();
 sg13g2_fill_2 FILLER_34_652 ();
 sg13g2_decap_8 FILLER_34_659 ();
 sg13g2_decap_4 FILLER_34_670 ();
 sg13g2_fill_1 FILLER_34_674 ();
 sg13g2_fill_1 FILLER_34_684 ();
 sg13g2_decap_4 FILLER_34_690 ();
 sg13g2_fill_1 FILLER_34_694 ();
 sg13g2_decap_4 FILLER_34_702 ();
 sg13g2_decap_4 FILLER_34_711 ();
 sg13g2_fill_2 FILLER_34_715 ();
 sg13g2_decap_8 FILLER_34_722 ();
 sg13g2_fill_2 FILLER_34_729 ();
 sg13g2_fill_1 FILLER_34_731 ();
 sg13g2_decap_8 FILLER_34_741 ();
 sg13g2_decap_8 FILLER_34_748 ();
 sg13g2_decap_8 FILLER_34_755 ();
 sg13g2_decap_8 FILLER_34_762 ();
 sg13g2_decap_4 FILLER_34_769 ();
 sg13g2_fill_1 FILLER_34_773 ();
 sg13g2_decap_8 FILLER_34_779 ();
 sg13g2_decap_8 FILLER_34_786 ();
 sg13g2_decap_8 FILLER_34_793 ();
 sg13g2_decap_8 FILLER_34_800 ();
 sg13g2_decap_8 FILLER_34_807 ();
 sg13g2_decap_8 FILLER_34_814 ();
 sg13g2_decap_8 FILLER_34_821 ();
 sg13g2_decap_8 FILLER_34_828 ();
 sg13g2_decap_8 FILLER_34_835 ();
 sg13g2_decap_8 FILLER_34_842 ();
 sg13g2_decap_8 FILLER_34_849 ();
 sg13g2_decap_8 FILLER_34_856 ();
 sg13g2_decap_8 FILLER_34_863 ();
 sg13g2_decap_8 FILLER_34_870 ();
 sg13g2_fill_1 FILLER_34_877 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_63 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_fill_1 FILLER_35_71 ();
 sg13g2_fill_1 FILLER_35_83 ();
 sg13g2_fill_2 FILLER_35_104 ();
 sg13g2_fill_2 FILLER_35_111 ();
 sg13g2_decap_8 FILLER_35_118 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_decap_8 FILLER_35_137 ();
 sg13g2_decap_8 FILLER_35_144 ();
 sg13g2_decap_4 FILLER_35_151 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_decap_8 FILLER_35_162 ();
 sg13g2_decap_4 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_179 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_211 ();
 sg13g2_decap_8 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_247 ();
 sg13g2_decap_8 FILLER_35_254 ();
 sg13g2_decap_8 FILLER_35_261 ();
 sg13g2_decap_8 FILLER_35_268 ();
 sg13g2_decap_8 FILLER_35_275 ();
 sg13g2_decap_8 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_fill_2 FILLER_35_296 ();
 sg13g2_decap_4 FILLER_35_304 ();
 sg13g2_fill_1 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_313 ();
 sg13g2_decap_8 FILLER_35_320 ();
 sg13g2_decap_8 FILLER_35_327 ();
 sg13g2_decap_4 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_349 ();
 sg13g2_decap_8 FILLER_35_356 ();
 sg13g2_decap_8 FILLER_35_363 ();
 sg13g2_fill_2 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_372 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_4 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_404 ();
 sg13g2_decap_8 FILLER_35_411 ();
 sg13g2_decap_4 FILLER_35_418 ();
 sg13g2_fill_2 FILLER_35_422 ();
 sg13g2_decap_8 FILLER_35_428 ();
 sg13g2_decap_4 FILLER_35_435 ();
 sg13g2_fill_2 FILLER_35_439 ();
 sg13g2_decap_8 FILLER_35_446 ();
 sg13g2_decap_4 FILLER_35_453 ();
 sg13g2_fill_2 FILLER_35_457 ();
 sg13g2_decap_8 FILLER_35_464 ();
 sg13g2_decap_8 FILLER_35_471 ();
 sg13g2_fill_2 FILLER_35_478 ();
 sg13g2_decap_8 FILLER_35_485 ();
 sg13g2_fill_2 FILLER_35_492 ();
 sg13g2_fill_1 FILLER_35_494 ();
 sg13g2_fill_1 FILLER_35_509 ();
 sg13g2_fill_2 FILLER_35_514 ();
 sg13g2_decap_8 FILLER_35_519 ();
 sg13g2_decap_8 FILLER_35_526 ();
 sg13g2_decap_8 FILLER_35_533 ();
 sg13g2_decap_8 FILLER_35_540 ();
 sg13g2_decap_4 FILLER_35_547 ();
 sg13g2_fill_1 FILLER_35_551 ();
 sg13g2_decap_4 FILLER_35_560 ();
 sg13g2_fill_1 FILLER_35_564 ();
 sg13g2_fill_1 FILLER_35_577 ();
 sg13g2_fill_2 FILLER_35_584 ();
 sg13g2_fill_1 FILLER_35_586 ();
 sg13g2_decap_8 FILLER_35_591 ();
 sg13g2_fill_2 FILLER_35_598 ();
 sg13g2_fill_1 FILLER_35_600 ();
 sg13g2_fill_1 FILLER_35_611 ();
 sg13g2_decap_8 FILLER_35_617 ();
 sg13g2_decap_4 FILLER_35_624 ();
 sg13g2_fill_1 FILLER_35_628 ();
 sg13g2_decap_8 FILLER_35_634 ();
 sg13g2_decap_8 FILLER_35_641 ();
 sg13g2_decap_8 FILLER_35_648 ();
 sg13g2_fill_2 FILLER_35_655 ();
 sg13g2_fill_2 FILLER_35_661 ();
 sg13g2_decap_8 FILLER_35_666 ();
 sg13g2_decap_8 FILLER_35_673 ();
 sg13g2_decap_4 FILLER_35_680 ();
 sg13g2_decap_8 FILLER_35_688 ();
 sg13g2_decap_8 FILLER_35_695 ();
 sg13g2_decap_8 FILLER_35_702 ();
 sg13g2_decap_8 FILLER_35_709 ();
 sg13g2_decap_4 FILLER_35_716 ();
 sg13g2_fill_1 FILLER_35_724 ();
 sg13g2_fill_2 FILLER_35_741 ();
 sg13g2_fill_2 FILLER_35_759 ();
 sg13g2_fill_1 FILLER_35_761 ();
 sg13g2_decap_8 FILLER_35_766 ();
 sg13g2_fill_2 FILLER_35_773 ();
 sg13g2_fill_1 FILLER_35_775 ();
 sg13g2_decap_8 FILLER_35_780 ();
 sg13g2_decap_8 FILLER_35_787 ();
 sg13g2_decap_8 FILLER_35_794 ();
 sg13g2_decap_8 FILLER_35_801 ();
 sg13g2_decap_8 FILLER_35_808 ();
 sg13g2_decap_8 FILLER_35_815 ();
 sg13g2_decap_8 FILLER_35_822 ();
 sg13g2_decap_8 FILLER_35_829 ();
 sg13g2_decap_8 FILLER_35_836 ();
 sg13g2_decap_8 FILLER_35_843 ();
 sg13g2_decap_8 FILLER_35_850 ();
 sg13g2_decap_8 FILLER_35_857 ();
 sg13g2_decap_8 FILLER_35_864 ();
 sg13g2_decap_8 FILLER_35_871 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_65 ();
 sg13g2_decap_8 FILLER_36_79 ();
 sg13g2_decap_8 FILLER_36_86 ();
 sg13g2_decap_8 FILLER_36_93 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_decap_4 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_111 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_fill_2 FILLER_36_147 ();
 sg13g2_fill_1 FILLER_36_149 ();
 sg13g2_decap_4 FILLER_36_159 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_decap_8 FILLER_36_186 ();
 sg13g2_decap_4 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_213 ();
 sg13g2_fill_2 FILLER_36_218 ();
 sg13g2_fill_2 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_decap_8 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_250 ();
 sg13g2_decap_8 FILLER_36_257 ();
 sg13g2_decap_8 FILLER_36_264 ();
 sg13g2_fill_2 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_278 ();
 sg13g2_fill_1 FILLER_36_294 ();
 sg13g2_fill_2 FILLER_36_300 ();
 sg13g2_decap_8 FILLER_36_314 ();
 sg13g2_decap_4 FILLER_36_321 ();
 sg13g2_decap_4 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_decap_8 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_fill_2 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_fill_2 FILLER_36_403 ();
 sg13g2_decap_4 FILLER_36_409 ();
 sg13g2_decap_8 FILLER_36_419 ();
 sg13g2_decap_8 FILLER_36_426 ();
 sg13g2_fill_1 FILLER_36_433 ();
 sg13g2_decap_4 FILLER_36_438 ();
 sg13g2_fill_2 FILLER_36_442 ();
 sg13g2_fill_2 FILLER_36_459 ();
 sg13g2_fill_2 FILLER_36_465 ();
 sg13g2_fill_2 FILLER_36_478 ();
 sg13g2_decap_8 FILLER_36_484 ();
 sg13g2_decap_8 FILLER_36_491 ();
 sg13g2_fill_2 FILLER_36_498 ();
 sg13g2_fill_1 FILLER_36_500 ();
 sg13g2_fill_2 FILLER_36_505 ();
 sg13g2_decap_8 FILLER_36_512 ();
 sg13g2_decap_8 FILLER_36_519 ();
 sg13g2_fill_1 FILLER_36_526 ();
 sg13g2_decap_8 FILLER_36_532 ();
 sg13g2_decap_8 FILLER_36_539 ();
 sg13g2_decap_8 FILLER_36_546 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_fill_2 FILLER_36_560 ();
 sg13g2_fill_1 FILLER_36_562 ();
 sg13g2_fill_2 FILLER_36_572 ();
 sg13g2_decap_4 FILLER_36_579 ();
 sg13g2_fill_1 FILLER_36_583 ();
 sg13g2_decap_8 FILLER_36_593 ();
 sg13g2_fill_2 FILLER_36_604 ();
 sg13g2_decap_8 FILLER_36_610 ();
 sg13g2_decap_8 FILLER_36_617 ();
 sg13g2_fill_2 FILLER_36_628 ();
 sg13g2_decap_4 FILLER_36_636 ();
 sg13g2_fill_2 FILLER_36_640 ();
 sg13g2_decap_8 FILLER_36_646 ();
 sg13g2_decap_8 FILLER_36_653 ();
 sg13g2_decap_4 FILLER_36_660 ();
 sg13g2_fill_1 FILLER_36_664 ();
 sg13g2_decap_4 FILLER_36_678 ();
 sg13g2_decap_8 FILLER_36_687 ();
 sg13g2_decap_8 FILLER_36_694 ();
 sg13g2_decap_8 FILLER_36_701 ();
 sg13g2_fill_2 FILLER_36_708 ();
 sg13g2_fill_2 FILLER_36_719 ();
 sg13g2_decap_4 FILLER_36_727 ();
 sg13g2_decap_4 FILLER_36_740 ();
 sg13g2_fill_1 FILLER_36_744 ();
 sg13g2_decap_8 FILLER_36_750 ();
 sg13g2_fill_2 FILLER_36_757 ();
 sg13g2_decap_4 FILLER_36_763 ();
 sg13g2_fill_1 FILLER_36_767 ();
 sg13g2_decap_8 FILLER_36_773 ();
 sg13g2_decap_8 FILLER_36_780 ();
 sg13g2_decap_8 FILLER_36_787 ();
 sg13g2_decap_8 FILLER_36_794 ();
 sg13g2_decap_8 FILLER_36_801 ();
 sg13g2_decap_8 FILLER_36_808 ();
 sg13g2_decap_8 FILLER_36_815 ();
 sg13g2_decap_8 FILLER_36_822 ();
 sg13g2_decap_8 FILLER_36_829 ();
 sg13g2_decap_8 FILLER_36_836 ();
 sg13g2_decap_8 FILLER_36_843 ();
 sg13g2_decap_8 FILLER_36_850 ();
 sg13g2_decap_8 FILLER_36_857 ();
 sg13g2_decap_8 FILLER_36_864 ();
 sg13g2_decap_8 FILLER_36_871 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_79 ();
 sg13g2_decap_8 FILLER_37_99 ();
 sg13g2_decap_8 FILLER_37_106 ();
 sg13g2_decap_4 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_117 ();
 sg13g2_fill_2 FILLER_37_123 ();
 sg13g2_fill_1 FILLER_37_125 ();
 sg13g2_decap_4 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_139 ();
 sg13g2_decap_8 FILLER_37_145 ();
 sg13g2_decap_4 FILLER_37_152 ();
 sg13g2_fill_1 FILLER_37_156 ();
 sg13g2_fill_1 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_183 ();
 sg13g2_decap_8 FILLER_37_194 ();
 sg13g2_decap_4 FILLER_37_211 ();
 sg13g2_decap_4 FILLER_37_219 ();
 sg13g2_decap_8 FILLER_37_227 ();
 sg13g2_decap_8 FILLER_37_234 ();
 sg13g2_decap_8 FILLER_37_241 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_fill_2 FILLER_37_254 ();
 sg13g2_fill_2 FILLER_37_261 ();
 sg13g2_decap_8 FILLER_37_267 ();
 sg13g2_fill_2 FILLER_37_274 ();
 sg13g2_fill_2 FILLER_37_282 ();
 sg13g2_fill_1 FILLER_37_284 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_310 ();
 sg13g2_fill_1 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_4 FILLER_37_323 ();
 sg13g2_fill_1 FILLER_37_327 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_decap_4 FILLER_37_340 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_decap_4 FILLER_37_351 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_decap_8 FILLER_37_362 ();
 sg13g2_decap_8 FILLER_37_369 ();
 sg13g2_decap_8 FILLER_37_376 ();
 sg13g2_decap_4 FILLER_37_383 ();
 sg13g2_fill_2 FILLER_37_387 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_417 ();
 sg13g2_decap_8 FILLER_37_424 ();
 sg13g2_decap_8 FILLER_37_431 ();
 sg13g2_decap_4 FILLER_37_453 ();
 sg13g2_decap_8 FILLER_37_461 ();
 sg13g2_decap_4 FILLER_37_468 ();
 sg13g2_fill_1 FILLER_37_472 ();
 sg13g2_fill_2 FILLER_37_477 ();
 sg13g2_fill_1 FILLER_37_479 ();
 sg13g2_decap_8 FILLER_37_506 ();
 sg13g2_decap_8 FILLER_37_513 ();
 sg13g2_fill_1 FILLER_37_520 ();
 sg13g2_fill_1 FILLER_37_529 ();
 sg13g2_fill_1 FILLER_37_533 ();
 sg13g2_fill_2 FILLER_37_540 ();
 sg13g2_fill_1 FILLER_37_542 ();
 sg13g2_decap_8 FILLER_37_549 ();
 sg13g2_decap_8 FILLER_37_556 ();
 sg13g2_fill_2 FILLER_37_563 ();
 sg13g2_fill_2 FILLER_37_576 ();
 sg13g2_decap_4 FILLER_37_583 ();
 sg13g2_decap_8 FILLER_37_596 ();
 sg13g2_fill_1 FILLER_37_603 ();
 sg13g2_decap_8 FILLER_37_609 ();
 sg13g2_decap_4 FILLER_37_622 ();
 sg13g2_decap_8 FILLER_37_632 ();
 sg13g2_decap_8 FILLER_37_639 ();
 sg13g2_decap_8 FILLER_37_646 ();
 sg13g2_fill_2 FILLER_37_653 ();
 sg13g2_fill_1 FILLER_37_655 ();
 sg13g2_decap_8 FILLER_37_666 ();
 sg13g2_decap_4 FILLER_37_673 ();
 sg13g2_fill_1 FILLER_37_677 ();
 sg13g2_fill_1 FILLER_37_701 ();
 sg13g2_decap_4 FILLER_37_712 ();
 sg13g2_decap_4 FILLER_37_739 ();
 sg13g2_decap_4 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_759 ();
 sg13g2_decap_8 FILLER_37_766 ();
 sg13g2_decap_8 FILLER_37_773 ();
 sg13g2_decap_8 FILLER_37_780 ();
 sg13g2_decap_8 FILLER_37_787 ();
 sg13g2_decap_8 FILLER_37_794 ();
 sg13g2_decap_8 FILLER_37_801 ();
 sg13g2_decap_8 FILLER_37_808 ();
 sg13g2_decap_8 FILLER_37_815 ();
 sg13g2_decap_8 FILLER_37_822 ();
 sg13g2_decap_8 FILLER_37_829 ();
 sg13g2_decap_8 FILLER_37_836 ();
 sg13g2_decap_8 FILLER_37_843 ();
 sg13g2_decap_8 FILLER_37_850 ();
 sg13g2_decap_8 FILLER_37_857 ();
 sg13g2_decap_8 FILLER_37_864 ();
 sg13g2_decap_8 FILLER_37_871 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_fill_2 FILLER_38_63 ();
 sg13g2_fill_1 FILLER_38_65 ();
 sg13g2_fill_1 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_78 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_98 ();
 sg13g2_decap_4 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_109 ();
 sg13g2_fill_1 FILLER_38_115 ();
 sg13g2_decap_4 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_138 ();
 sg13g2_decap_8 FILLER_38_145 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_160 ();
 sg13g2_decap_8 FILLER_38_167 ();
 sg13g2_decap_8 FILLER_38_174 ();
 sg13g2_decap_8 FILLER_38_181 ();
 sg13g2_decap_8 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_decap_4 FILLER_38_200 ();
 sg13g2_fill_1 FILLER_38_204 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_decap_8 FILLER_38_270 ();
 sg13g2_decap_8 FILLER_38_277 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_decap_8 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_298 ();
 sg13g2_decap_4 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_decap_8 FILLER_38_331 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_fill_1 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_fill_2 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_fill_1 FILLER_38_409 ();
 sg13g2_decap_8 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_425 ();
 sg13g2_decap_8 FILLER_38_432 ();
 sg13g2_decap_8 FILLER_38_439 ();
 sg13g2_decap_8 FILLER_38_446 ();
 sg13g2_decap_8 FILLER_38_453 ();
 sg13g2_decap_8 FILLER_38_460 ();
 sg13g2_decap_4 FILLER_38_467 ();
 sg13g2_fill_2 FILLER_38_471 ();
 sg13g2_decap_4 FILLER_38_477 ();
 sg13g2_fill_2 FILLER_38_489 ();
 sg13g2_fill_1 FILLER_38_491 ();
 sg13g2_fill_2 FILLER_38_496 ();
 sg13g2_decap_8 FILLER_38_505 ();
 sg13g2_decap_8 FILLER_38_512 ();
 sg13g2_decap_8 FILLER_38_519 ();
 sg13g2_decap_8 FILLER_38_526 ();
 sg13g2_decap_8 FILLER_38_533 ();
 sg13g2_decap_8 FILLER_38_540 ();
 sg13g2_decap_8 FILLER_38_553 ();
 sg13g2_decap_4 FILLER_38_560 ();
 sg13g2_fill_1 FILLER_38_564 ();
 sg13g2_decap_8 FILLER_38_574 ();
 sg13g2_decap_8 FILLER_38_581 ();
 sg13g2_decap_8 FILLER_38_588 ();
 sg13g2_decap_4 FILLER_38_595 ();
 sg13g2_fill_2 FILLER_38_599 ();
 sg13g2_decap_8 FILLER_38_610 ();
 sg13g2_decap_4 FILLER_38_626 ();
 sg13g2_fill_2 FILLER_38_630 ();
 sg13g2_decap_8 FILLER_38_670 ();
 sg13g2_decap_8 FILLER_38_677 ();
 sg13g2_fill_2 FILLER_38_684 ();
 sg13g2_decap_8 FILLER_38_695 ();
 sg13g2_decap_8 FILLER_38_702 ();
 sg13g2_decap_8 FILLER_38_709 ();
 sg13g2_decap_8 FILLER_38_716 ();
 sg13g2_decap_8 FILLER_38_723 ();
 sg13g2_decap_4 FILLER_38_730 ();
 sg13g2_fill_1 FILLER_38_734 ();
 sg13g2_decap_8 FILLER_38_744 ();
 sg13g2_decap_8 FILLER_38_751 ();
 sg13g2_decap_8 FILLER_38_758 ();
 sg13g2_fill_2 FILLER_38_765 ();
 sg13g2_decap_8 FILLER_38_776 ();
 sg13g2_decap_8 FILLER_38_783 ();
 sg13g2_decap_8 FILLER_38_790 ();
 sg13g2_decap_8 FILLER_38_797 ();
 sg13g2_decap_8 FILLER_38_804 ();
 sg13g2_decap_8 FILLER_38_811 ();
 sg13g2_decap_8 FILLER_38_818 ();
 sg13g2_decap_8 FILLER_38_825 ();
 sg13g2_decap_8 FILLER_38_832 ();
 sg13g2_decap_8 FILLER_38_839 ();
 sg13g2_decap_8 FILLER_38_846 ();
 sg13g2_decap_8 FILLER_38_853 ();
 sg13g2_decap_8 FILLER_38_860 ();
 sg13g2_decap_8 FILLER_38_867 ();
 sg13g2_decap_4 FILLER_38_874 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_fill_2 FILLER_39_53 ();
 sg13g2_fill_1 FILLER_39_55 ();
 sg13g2_decap_8 FILLER_39_64 ();
 sg13g2_fill_1 FILLER_39_71 ();
 sg13g2_fill_1 FILLER_39_76 ();
 sg13g2_decap_8 FILLER_39_82 ();
 sg13g2_decap_8 FILLER_39_92 ();
 sg13g2_decap_8 FILLER_39_99 ();
 sg13g2_decap_4 FILLER_39_106 ();
 sg13g2_fill_1 FILLER_39_113 ();
 sg13g2_fill_2 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_4 FILLER_39_133 ();
 sg13g2_fill_2 FILLER_39_140 ();
 sg13g2_decap_4 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_163 ();
 sg13g2_decap_4 FILLER_39_170 ();
 sg13g2_decap_4 FILLER_39_178 ();
 sg13g2_fill_1 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_192 ();
 sg13g2_decap_8 FILLER_39_199 ();
 sg13g2_decap_4 FILLER_39_206 ();
 sg13g2_decap_8 FILLER_39_214 ();
 sg13g2_decap_8 FILLER_39_221 ();
 sg13g2_fill_2 FILLER_39_228 ();
 sg13g2_decap_8 FILLER_39_234 ();
 sg13g2_decap_4 FILLER_39_241 ();
 sg13g2_fill_2 FILLER_39_245 ();
 sg13g2_decap_4 FILLER_39_251 ();
 sg13g2_fill_2 FILLER_39_255 ();
 sg13g2_fill_1 FILLER_39_261 ();
 sg13g2_decap_8 FILLER_39_267 ();
 sg13g2_decap_8 FILLER_39_279 ();
 sg13g2_fill_1 FILLER_39_286 ();
 sg13g2_decap_4 FILLER_39_291 ();
 sg13g2_decap_4 FILLER_39_299 ();
 sg13g2_decap_8 FILLER_39_312 ();
 sg13g2_fill_2 FILLER_39_319 ();
 sg13g2_fill_1 FILLER_39_321 ();
 sg13g2_decap_4 FILLER_39_330 ();
 sg13g2_fill_2 FILLER_39_334 ();
 sg13g2_fill_2 FILLER_39_342 ();
 sg13g2_fill_1 FILLER_39_344 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_fill_1 FILLER_39_371 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_decap_4 FILLER_39_383 ();
 sg13g2_fill_2 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_39_414 ();
 sg13g2_decap_8 FILLER_39_421 ();
 sg13g2_fill_2 FILLER_39_428 ();
 sg13g2_fill_1 FILLER_39_430 ();
 sg13g2_decap_4 FILLER_39_436 ();
 sg13g2_fill_1 FILLER_39_440 ();
 sg13g2_decap_8 FILLER_39_449 ();
 sg13g2_decap_8 FILLER_39_456 ();
 sg13g2_decap_8 FILLER_39_463 ();
 sg13g2_decap_8 FILLER_39_470 ();
 sg13g2_decap_8 FILLER_39_477 ();
 sg13g2_decap_8 FILLER_39_484 ();
 sg13g2_decap_4 FILLER_39_491 ();
 sg13g2_fill_2 FILLER_39_500 ();
 sg13g2_fill_1 FILLER_39_502 ();
 sg13g2_decap_8 FILLER_39_507 ();
 sg13g2_decap_4 FILLER_39_514 ();
 sg13g2_fill_2 FILLER_39_518 ();
 sg13g2_fill_2 FILLER_39_523 ();
 sg13g2_decap_8 FILLER_39_531 ();
 sg13g2_fill_1 FILLER_39_538 ();
 sg13g2_decap_4 FILLER_39_547 ();
 sg13g2_fill_2 FILLER_39_551 ();
 sg13g2_fill_1 FILLER_39_557 ();
 sg13g2_decap_8 FILLER_39_584 ();
 sg13g2_decap_8 FILLER_39_591 ();
 sg13g2_decap_8 FILLER_39_615 ();
 sg13g2_decap_8 FILLER_39_622 ();
 sg13g2_decap_8 FILLER_39_629 ();
 sg13g2_decap_8 FILLER_39_636 ();
 sg13g2_fill_1 FILLER_39_647 ();
 sg13g2_fill_2 FILLER_39_653 ();
 sg13g2_fill_1 FILLER_39_655 ();
 sg13g2_decap_8 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_672 ();
 sg13g2_decap_8 FILLER_39_688 ();
 sg13g2_decap_8 FILLER_39_695 ();
 sg13g2_decap_8 FILLER_39_702 ();
 sg13g2_fill_2 FILLER_39_709 ();
 sg13g2_fill_1 FILLER_39_711 ();
 sg13g2_decap_8 FILLER_39_723 ();
 sg13g2_decap_8 FILLER_39_730 ();
 sg13g2_decap_8 FILLER_39_737 ();
 sg13g2_decap_8 FILLER_39_744 ();
 sg13g2_decap_8 FILLER_39_751 ();
 sg13g2_decap_8 FILLER_39_758 ();
 sg13g2_decap_8 FILLER_39_765 ();
 sg13g2_decap_8 FILLER_39_772 ();
 sg13g2_decap_8 FILLER_39_779 ();
 sg13g2_decap_8 FILLER_39_786 ();
 sg13g2_decap_8 FILLER_39_793 ();
 sg13g2_decap_8 FILLER_39_800 ();
 sg13g2_decap_8 FILLER_39_807 ();
 sg13g2_decap_8 FILLER_39_814 ();
 sg13g2_decap_8 FILLER_39_821 ();
 sg13g2_decap_8 FILLER_39_828 ();
 sg13g2_decap_8 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_842 ();
 sg13g2_decap_8 FILLER_39_849 ();
 sg13g2_decap_8 FILLER_39_856 ();
 sg13g2_decap_8 FILLER_39_863 ();
 sg13g2_decap_8 FILLER_39_870 ();
 sg13g2_fill_1 FILLER_39_877 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_fill_2 FILLER_40_63 ();
 sg13g2_decap_4 FILLER_40_69 ();
 sg13g2_decap_8 FILLER_40_78 ();
 sg13g2_decap_8 FILLER_40_85 ();
 sg13g2_decap_8 FILLER_40_92 ();
 sg13g2_decap_8 FILLER_40_99 ();
 sg13g2_decap_8 FILLER_40_106 ();
 sg13g2_decap_8 FILLER_40_113 ();
 sg13g2_decap_8 FILLER_40_120 ();
 sg13g2_decap_8 FILLER_40_127 ();
 sg13g2_decap_8 FILLER_40_134 ();
 sg13g2_decap_8 FILLER_40_141 ();
 sg13g2_decap_8 FILLER_40_148 ();
 sg13g2_decap_8 FILLER_40_155 ();
 sg13g2_fill_2 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_164 ();
 sg13g2_decap_8 FILLER_40_170 ();
 sg13g2_fill_1 FILLER_40_177 ();
 sg13g2_decap_4 FILLER_40_187 ();
 sg13g2_decap_8 FILLER_40_205 ();
 sg13g2_decap_8 FILLER_40_212 ();
 sg13g2_fill_2 FILLER_40_219 ();
 sg13g2_fill_1 FILLER_40_221 ();
 sg13g2_decap_8 FILLER_40_226 ();
 sg13g2_fill_1 FILLER_40_233 ();
 sg13g2_decap_8 FILLER_40_237 ();
 sg13g2_decap_4 FILLER_40_244 ();
 sg13g2_fill_2 FILLER_40_248 ();
 sg13g2_decap_8 FILLER_40_260 ();
 sg13g2_decap_8 FILLER_40_267 ();
 sg13g2_decap_8 FILLER_40_274 ();
 sg13g2_decap_8 FILLER_40_281 ();
 sg13g2_decap_4 FILLER_40_288 ();
 sg13g2_fill_1 FILLER_40_292 ();
 sg13g2_fill_2 FILLER_40_298 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_fill_2 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_4 FILLER_40_364 ();
 sg13g2_fill_2 FILLER_40_368 ();
 sg13g2_fill_1 FILLER_40_379 ();
 sg13g2_decap_8 FILLER_40_386 ();
 sg13g2_fill_1 FILLER_40_393 ();
 sg13g2_decap_8 FILLER_40_398 ();
 sg13g2_decap_8 FILLER_40_405 ();
 sg13g2_decap_8 FILLER_40_412 ();
 sg13g2_decap_8 FILLER_40_419 ();
 sg13g2_decap_8 FILLER_40_442 ();
 sg13g2_decap_8 FILLER_40_449 ();
 sg13g2_decap_8 FILLER_40_456 ();
 sg13g2_decap_8 FILLER_40_463 ();
 sg13g2_fill_2 FILLER_40_470 ();
 sg13g2_fill_1 FILLER_40_472 ();
 sg13g2_decap_8 FILLER_40_477 ();
 sg13g2_decap_8 FILLER_40_484 ();
 sg13g2_decap_4 FILLER_40_491 ();
 sg13g2_fill_1 FILLER_40_495 ();
 sg13g2_decap_4 FILLER_40_500 ();
 sg13g2_decap_4 FILLER_40_514 ();
 sg13g2_fill_1 FILLER_40_518 ();
 sg13g2_fill_2 FILLER_40_524 ();
 sg13g2_fill_2 FILLER_40_529 ();
 sg13g2_decap_4 FILLER_40_535 ();
 sg13g2_decap_4 FILLER_40_543 ();
 sg13g2_fill_1 FILLER_40_547 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_fill_2 FILLER_40_575 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_decap_4 FILLER_40_588 ();
 sg13g2_fill_1 FILLER_40_592 ();
 sg13g2_decap_4 FILLER_40_598 ();
 sg13g2_fill_1 FILLER_40_602 ();
 sg13g2_fill_2 FILLER_40_608 ();
 sg13g2_decap_8 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_4 FILLER_40_644 ();
 sg13g2_fill_1 FILLER_40_648 ();
 sg13g2_decap_8 FILLER_40_653 ();
 sg13g2_fill_2 FILLER_40_660 ();
 sg13g2_fill_1 FILLER_40_662 ();
 sg13g2_decap_8 FILLER_40_668 ();
 sg13g2_fill_2 FILLER_40_675 ();
 sg13g2_fill_1 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_689 ();
 sg13g2_decap_4 FILLER_40_696 ();
 sg13g2_fill_1 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_705 ();
 sg13g2_decap_4 FILLER_40_712 ();
 sg13g2_fill_2 FILLER_40_716 ();
 sg13g2_decap_8 FILLER_40_724 ();
 sg13g2_fill_2 FILLER_40_731 ();
 sg13g2_decap_8 FILLER_40_737 ();
 sg13g2_decap_8 FILLER_40_744 ();
 sg13g2_fill_2 FILLER_40_751 ();
 sg13g2_fill_2 FILLER_40_768 ();
 sg13g2_fill_1 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_775 ();
 sg13g2_decap_8 FILLER_40_782 ();
 sg13g2_decap_8 FILLER_40_789 ();
 sg13g2_decap_8 FILLER_40_796 ();
 sg13g2_decap_8 FILLER_40_803 ();
 sg13g2_decap_8 FILLER_40_810 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_decap_8 FILLER_40_824 ();
 sg13g2_decap_8 FILLER_40_831 ();
 sg13g2_decap_8 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_845 ();
 sg13g2_decap_8 FILLER_40_852 ();
 sg13g2_decap_8 FILLER_40_859 ();
 sg13g2_decap_8 FILLER_40_866 ();
 sg13g2_decap_4 FILLER_40_873 ();
 sg13g2_fill_1 FILLER_40_877 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_fill_1 FILLER_41_70 ();
 sg13g2_decap_4 FILLER_41_76 ();
 sg13g2_decap_8 FILLER_41_85 ();
 sg13g2_decap_8 FILLER_41_92 ();
 sg13g2_decap_4 FILLER_41_99 ();
 sg13g2_fill_2 FILLER_41_103 ();
 sg13g2_decap_8 FILLER_41_111 ();
 sg13g2_decap_8 FILLER_41_118 ();
 sg13g2_decap_8 FILLER_41_125 ();
 sg13g2_decap_4 FILLER_41_132 ();
 sg13g2_fill_1 FILLER_41_136 ();
 sg13g2_decap_8 FILLER_41_141 ();
 sg13g2_decap_8 FILLER_41_148 ();
 sg13g2_decap_8 FILLER_41_155 ();
 sg13g2_decap_4 FILLER_41_162 ();
 sg13g2_decap_8 FILLER_41_170 ();
 sg13g2_decap_4 FILLER_41_181 ();
 sg13g2_decap_8 FILLER_41_197 ();
 sg13g2_decap_8 FILLER_41_204 ();
 sg13g2_decap_8 FILLER_41_211 ();
 sg13g2_decap_8 FILLER_41_218 ();
 sg13g2_decap_8 FILLER_41_225 ();
 sg13g2_decap_8 FILLER_41_232 ();
 sg13g2_decap_8 FILLER_41_239 ();
 sg13g2_decap_8 FILLER_41_255 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_278 ();
 sg13g2_decap_8 FILLER_41_285 ();
 sg13g2_fill_1 FILLER_41_292 ();
 sg13g2_decap_4 FILLER_41_298 ();
 sg13g2_fill_2 FILLER_41_302 ();
 sg13g2_decap_8 FILLER_41_314 ();
 sg13g2_decap_8 FILLER_41_321 ();
 sg13g2_fill_2 FILLER_41_328 ();
 sg13g2_decap_8 FILLER_41_349 ();
 sg13g2_decap_4 FILLER_41_361 ();
 sg13g2_fill_2 FILLER_41_365 ();
 sg13g2_fill_2 FILLER_41_376 ();
 sg13g2_fill_2 FILLER_41_383 ();
 sg13g2_fill_1 FILLER_41_385 ();
 sg13g2_decap_4 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_398 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_fill_1 FILLER_41_427 ();
 sg13g2_decap_4 FILLER_41_437 ();
 sg13g2_decap_8 FILLER_41_446 ();
 sg13g2_decap_4 FILLER_41_462 ();
 sg13g2_fill_1 FILLER_41_466 ();
 sg13g2_decap_8 FILLER_41_472 ();
 sg13g2_fill_2 FILLER_41_479 ();
 sg13g2_decap_8 FILLER_41_485 ();
 sg13g2_decap_8 FILLER_41_492 ();
 sg13g2_fill_1 FILLER_41_499 ();
 sg13g2_fill_2 FILLER_41_507 ();
 sg13g2_decap_4 FILLER_41_519 ();
 sg13g2_decap_4 FILLER_41_529 ();
 sg13g2_fill_2 FILLER_41_533 ();
 sg13g2_decap_8 FILLER_41_542 ();
 sg13g2_decap_4 FILLER_41_549 ();
 sg13g2_fill_1 FILLER_41_553 ();
 sg13g2_decap_8 FILLER_41_562 ();
 sg13g2_decap_4 FILLER_41_569 ();
 sg13g2_fill_2 FILLER_41_578 ();
 sg13g2_fill_1 FILLER_41_580 ();
 sg13g2_decap_4 FILLER_41_591 ();
 sg13g2_fill_2 FILLER_41_600 ();
 sg13g2_decap_8 FILLER_41_610 ();
 sg13g2_decap_8 FILLER_41_617 ();
 sg13g2_decap_8 FILLER_41_624 ();
 sg13g2_decap_8 FILLER_41_631 ();
 sg13g2_fill_2 FILLER_41_638 ();
 sg13g2_fill_1 FILLER_41_640 ();
 sg13g2_fill_2 FILLER_41_646 ();
 sg13g2_fill_1 FILLER_41_667 ();
 sg13g2_decap_8 FILLER_41_674 ();
 sg13g2_decap_8 FILLER_41_681 ();
 sg13g2_decap_4 FILLER_41_688 ();
 sg13g2_fill_2 FILLER_41_692 ();
 sg13g2_fill_2 FILLER_41_698 ();
 sg13g2_fill_1 FILLER_41_700 ();
 sg13g2_fill_1 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_713 ();
 sg13g2_decap_4 FILLER_41_720 ();
 sg13g2_fill_1 FILLER_41_724 ();
 sg13g2_fill_2 FILLER_41_737 ();
 sg13g2_fill_1 FILLER_41_739 ();
 sg13g2_fill_2 FILLER_41_747 ();
 sg13g2_fill_1 FILLER_41_749 ();
 sg13g2_fill_2 FILLER_41_754 ();
 sg13g2_fill_1 FILLER_41_756 ();
 sg13g2_fill_2 FILLER_41_765 ();
 sg13g2_fill_1 FILLER_41_767 ();
 sg13g2_fill_1 FILLER_41_772 ();
 sg13g2_decap_8 FILLER_41_785 ();
 sg13g2_decap_8 FILLER_41_792 ();
 sg13g2_decap_8 FILLER_41_799 ();
 sg13g2_decap_8 FILLER_41_806 ();
 sg13g2_decap_8 FILLER_41_813 ();
 sg13g2_decap_8 FILLER_41_820 ();
 sg13g2_decap_8 FILLER_41_827 ();
 sg13g2_decap_8 FILLER_41_834 ();
 sg13g2_decap_8 FILLER_41_841 ();
 sg13g2_decap_8 FILLER_41_848 ();
 sg13g2_decap_8 FILLER_41_855 ();
 sg13g2_decap_8 FILLER_41_862 ();
 sg13g2_decap_8 FILLER_41_869 ();
 sg13g2_fill_2 FILLER_41_876 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_4 FILLER_42_56 ();
 sg13g2_fill_2 FILLER_42_73 ();
 sg13g2_fill_1 FILLER_42_80 ();
 sg13g2_decap_8 FILLER_42_86 ();
 sg13g2_decap_8 FILLER_42_93 ();
 sg13g2_decap_8 FILLER_42_100 ();
 sg13g2_decap_8 FILLER_42_107 ();
 sg13g2_decap_8 FILLER_42_114 ();
 sg13g2_decap_8 FILLER_42_121 ();
 sg13g2_decap_8 FILLER_42_128 ();
 sg13g2_fill_1 FILLER_42_135 ();
 sg13g2_decap_4 FILLER_42_141 ();
 sg13g2_fill_1 FILLER_42_145 ();
 sg13g2_decap_8 FILLER_42_162 ();
 sg13g2_decap_4 FILLER_42_169 ();
 sg13g2_fill_1 FILLER_42_173 ();
 sg13g2_decap_4 FILLER_42_179 ();
 sg13g2_fill_1 FILLER_42_183 ();
 sg13g2_decap_8 FILLER_42_201 ();
 sg13g2_fill_2 FILLER_42_208 ();
 sg13g2_decap_8 FILLER_42_214 ();
 sg13g2_fill_2 FILLER_42_221 ();
 sg13g2_fill_1 FILLER_42_223 ();
 sg13g2_decap_8 FILLER_42_229 ();
 sg13g2_fill_1 FILLER_42_236 ();
 sg13g2_fill_2 FILLER_42_242 ();
 sg13g2_fill_1 FILLER_42_244 ();
 sg13g2_decap_8 FILLER_42_254 ();
 sg13g2_decap_8 FILLER_42_261 ();
 sg13g2_decap_8 FILLER_42_268 ();
 sg13g2_decap_8 FILLER_42_275 ();
 sg13g2_decap_8 FILLER_42_282 ();
 sg13g2_fill_2 FILLER_42_289 ();
 sg13g2_fill_1 FILLER_42_302 ();
 sg13g2_decap_4 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_316 ();
 sg13g2_decap_8 FILLER_42_323 ();
 sg13g2_decap_4 FILLER_42_335 ();
 sg13g2_fill_2 FILLER_42_339 ();
 sg13g2_fill_2 FILLER_42_346 ();
 sg13g2_decap_8 FILLER_42_352 ();
 sg13g2_fill_2 FILLER_42_359 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_decap_4 FILLER_42_368 ();
 sg13g2_fill_1 FILLER_42_372 ();
 sg13g2_decap_4 FILLER_42_377 ();
 sg13g2_fill_1 FILLER_42_381 ();
 sg13g2_decap_8 FILLER_42_386 ();
 sg13g2_decap_8 FILLER_42_393 ();
 sg13g2_decap_4 FILLER_42_405 ();
 sg13g2_fill_1 FILLER_42_414 ();
 sg13g2_decap_4 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_428 ();
 sg13g2_decap_8 FILLER_42_435 ();
 sg13g2_decap_4 FILLER_42_442 ();
 sg13g2_fill_2 FILLER_42_446 ();
 sg13g2_decap_4 FILLER_42_452 ();
 sg13g2_decap_8 FILLER_42_471 ();
 sg13g2_decap_8 FILLER_42_478 ();
 sg13g2_decap_4 FILLER_42_499 ();
 sg13g2_fill_1 FILLER_42_503 ();
 sg13g2_decap_4 FILLER_42_508 ();
 sg13g2_decap_8 FILLER_42_519 ();
 sg13g2_decap_8 FILLER_42_526 ();
 sg13g2_decap_8 FILLER_42_533 ();
 sg13g2_decap_8 FILLER_42_545 ();
 sg13g2_decap_8 FILLER_42_552 ();
 sg13g2_fill_1 FILLER_42_559 ();
 sg13g2_fill_2 FILLER_42_566 ();
 sg13g2_fill_2 FILLER_42_573 ();
 sg13g2_fill_1 FILLER_42_582 ();
 sg13g2_fill_1 FILLER_42_592 ();
 sg13g2_fill_1 FILLER_42_597 ();
 sg13g2_decap_4 FILLER_42_602 ();
 sg13g2_fill_2 FILLER_42_611 ();
 sg13g2_fill_1 FILLER_42_613 ();
 sg13g2_decap_8 FILLER_42_619 ();
 sg13g2_decap_8 FILLER_42_626 ();
 sg13g2_decap_8 FILLER_42_633 ();
 sg13g2_decap_4 FILLER_42_640 ();
 sg13g2_fill_1 FILLER_42_644 ();
 sg13g2_decap_8 FILLER_42_650 ();
 sg13g2_fill_1 FILLER_42_657 ();
 sg13g2_fill_2 FILLER_42_662 ();
 sg13g2_fill_1 FILLER_42_664 ();
 sg13g2_fill_1 FILLER_42_678 ();
 sg13g2_decap_8 FILLER_42_689 ();
 sg13g2_decap_8 FILLER_42_696 ();
 sg13g2_fill_2 FILLER_42_703 ();
 sg13g2_decap_8 FILLER_42_708 ();
 sg13g2_decap_8 FILLER_42_715 ();
 sg13g2_decap_8 FILLER_42_722 ();
 sg13g2_decap_8 FILLER_42_729 ();
 sg13g2_fill_2 FILLER_42_736 ();
 sg13g2_decap_8 FILLER_42_750 ();
 sg13g2_decap_8 FILLER_42_757 ();
 sg13g2_fill_1 FILLER_42_764 ();
 sg13g2_decap_8 FILLER_42_774 ();
 sg13g2_decap_8 FILLER_42_781 ();
 sg13g2_decap_8 FILLER_42_788 ();
 sg13g2_decap_8 FILLER_42_795 ();
 sg13g2_decap_8 FILLER_42_802 ();
 sg13g2_decap_8 FILLER_42_809 ();
 sg13g2_decap_8 FILLER_42_816 ();
 sg13g2_decap_8 FILLER_42_823 ();
 sg13g2_decap_8 FILLER_42_830 ();
 sg13g2_decap_8 FILLER_42_837 ();
 sg13g2_decap_8 FILLER_42_844 ();
 sg13g2_decap_8 FILLER_42_851 ();
 sg13g2_decap_8 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_42_865 ();
 sg13g2_decap_4 FILLER_42_872 ();
 sg13g2_fill_2 FILLER_42_876 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_fill_1 FILLER_43_56 ();
 sg13g2_decap_4 FILLER_43_70 ();
 sg13g2_fill_1 FILLER_43_78 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_4 FILLER_43_105 ();
 sg13g2_fill_2 FILLER_43_123 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_fill_1 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_146 ();
 sg13g2_fill_1 FILLER_43_153 ();
 sg13g2_decap_8 FILLER_43_158 ();
 sg13g2_fill_1 FILLER_43_165 ();
 sg13g2_decap_4 FILLER_43_171 ();
 sg13g2_fill_1 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_181 ();
 sg13g2_fill_1 FILLER_43_188 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_4 FILLER_43_203 ();
 sg13g2_fill_2 FILLER_43_207 ();
 sg13g2_decap_4 FILLER_43_212 ();
 sg13g2_fill_2 FILLER_43_216 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_decap_4 FILLER_43_228 ();
 sg13g2_fill_1 FILLER_43_236 ();
 sg13g2_decap_4 FILLER_43_242 ();
 sg13g2_decap_8 FILLER_43_250 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_311 ();
 sg13g2_decap_4 FILLER_43_318 ();
 sg13g2_fill_2 FILLER_43_322 ();
 sg13g2_decap_4 FILLER_43_328 ();
 sg13g2_decap_4 FILLER_43_335 ();
 sg13g2_fill_1 FILLER_43_339 ();
 sg13g2_decap_8 FILLER_43_344 ();
 sg13g2_decap_8 FILLER_43_351 ();
 sg13g2_decap_8 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_365 ();
 sg13g2_decap_4 FILLER_43_372 ();
 sg13g2_fill_2 FILLER_43_376 ();
 sg13g2_fill_2 FILLER_43_386 ();
 sg13g2_fill_1 FILLER_43_388 ();
 sg13g2_fill_1 FILLER_43_401 ();
 sg13g2_fill_1 FILLER_43_411 ();
 sg13g2_decap_8 FILLER_43_430 ();
 sg13g2_decap_8 FILLER_43_437 ();
 sg13g2_fill_2 FILLER_43_444 ();
 sg13g2_fill_1 FILLER_43_446 ();
 sg13g2_decap_8 FILLER_43_451 ();
 sg13g2_fill_1 FILLER_43_458 ();
 sg13g2_fill_2 FILLER_43_465 ();
 sg13g2_fill_1 FILLER_43_467 ();
 sg13g2_decap_8 FILLER_43_481 ();
 sg13g2_decap_8 FILLER_43_488 ();
 sg13g2_decap_4 FILLER_43_495 ();
 sg13g2_decap_8 FILLER_43_503 ();
 sg13g2_decap_8 FILLER_43_510 ();
 sg13g2_decap_4 FILLER_43_517 ();
 sg13g2_fill_2 FILLER_43_521 ();
 sg13g2_decap_8 FILLER_43_528 ();
 sg13g2_decap_8 FILLER_43_535 ();
 sg13g2_decap_8 FILLER_43_542 ();
 sg13g2_decap_8 FILLER_43_549 ();
 sg13g2_decap_8 FILLER_43_556 ();
 sg13g2_decap_8 FILLER_43_563 ();
 sg13g2_decap_8 FILLER_43_570 ();
 sg13g2_decap_8 FILLER_43_577 ();
 sg13g2_decap_8 FILLER_43_584 ();
 sg13g2_decap_8 FILLER_43_591 ();
 sg13g2_decap_8 FILLER_43_598 ();
 sg13g2_fill_2 FILLER_43_618 ();
 sg13g2_decap_8 FILLER_43_625 ();
 sg13g2_decap_8 FILLER_43_632 ();
 sg13g2_decap_8 FILLER_43_639 ();
 sg13g2_decap_4 FILLER_43_646 ();
 sg13g2_fill_2 FILLER_43_650 ();
 sg13g2_decap_8 FILLER_43_656 ();
 sg13g2_decap_8 FILLER_43_663 ();
 sg13g2_fill_2 FILLER_43_674 ();
 sg13g2_fill_1 FILLER_43_676 ();
 sg13g2_fill_1 FILLER_43_686 ();
 sg13g2_decap_8 FILLER_43_692 ();
 sg13g2_decap_4 FILLER_43_699 ();
 sg13g2_fill_2 FILLER_43_703 ();
 sg13g2_decap_8 FILLER_43_709 ();
 sg13g2_decap_8 FILLER_43_716 ();
 sg13g2_decap_8 FILLER_43_723 ();
 sg13g2_decap_4 FILLER_43_734 ();
 sg13g2_decap_8 FILLER_43_746 ();
 sg13g2_decap_8 FILLER_43_753 ();
 sg13g2_decap_8 FILLER_43_760 ();
 sg13g2_decap_8 FILLER_43_767 ();
 sg13g2_decap_8 FILLER_43_774 ();
 sg13g2_decap_8 FILLER_43_781 ();
 sg13g2_decap_8 FILLER_43_788 ();
 sg13g2_decap_8 FILLER_43_795 ();
 sg13g2_decap_8 FILLER_43_802 ();
 sg13g2_decap_8 FILLER_43_809 ();
 sg13g2_decap_8 FILLER_43_816 ();
 sg13g2_decap_8 FILLER_43_823 ();
 sg13g2_decap_8 FILLER_43_830 ();
 sg13g2_decap_8 FILLER_43_837 ();
 sg13g2_decap_8 FILLER_43_844 ();
 sg13g2_decap_8 FILLER_43_851 ();
 sg13g2_decap_8 FILLER_43_858 ();
 sg13g2_decap_8 FILLER_43_865 ();
 sg13g2_decap_4 FILLER_43_872 ();
 sg13g2_fill_2 FILLER_43_876 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_4 FILLER_44_49 ();
 sg13g2_fill_1 FILLER_44_53 ();
 sg13g2_decap_8 FILLER_44_62 ();
 sg13g2_decap_4 FILLER_44_69 ();
 sg13g2_fill_2 FILLER_44_73 ();
 sg13g2_decap_8 FILLER_44_79 ();
 sg13g2_decap_4 FILLER_44_86 ();
 sg13g2_fill_1 FILLER_44_90 ();
 sg13g2_fill_2 FILLER_44_105 ();
 sg13g2_fill_1 FILLER_44_107 ();
 sg13g2_decap_4 FILLER_44_116 ();
 sg13g2_fill_1 FILLER_44_120 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_fill_2 FILLER_44_133 ();
 sg13g2_fill_1 FILLER_44_135 ();
 sg13g2_decap_8 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_fill_1 FILLER_44_165 ();
 sg13g2_fill_1 FILLER_44_173 ();
 sg13g2_fill_2 FILLER_44_178 ();
 sg13g2_fill_2 FILLER_44_189 ();
 sg13g2_decap_4 FILLER_44_215 ();
 sg13g2_fill_1 FILLER_44_219 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_4 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_4 FILLER_44_277 ();
 sg13g2_fill_2 FILLER_44_281 ();
 sg13g2_decap_8 FILLER_44_288 ();
 sg13g2_decap_8 FILLER_44_305 ();
 sg13g2_decap_8 FILLER_44_312 ();
 sg13g2_fill_1 FILLER_44_319 ();
 sg13g2_decap_4 FILLER_44_335 ();
 sg13g2_fill_2 FILLER_44_339 ();
 sg13g2_decap_4 FILLER_44_345 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_decap_8 FILLER_44_358 ();
 sg13g2_decap_8 FILLER_44_365 ();
 sg13g2_fill_1 FILLER_44_372 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_4 FILLER_44_411 ();
 sg13g2_fill_2 FILLER_44_415 ();
 sg13g2_fill_2 FILLER_44_420 ();
 sg13g2_fill_1 FILLER_44_422 ();
 sg13g2_decap_8 FILLER_44_428 ();
 sg13g2_decap_4 FILLER_44_435 ();
 sg13g2_fill_1 FILLER_44_439 ();
 sg13g2_decap_8 FILLER_44_450 ();
 sg13g2_decap_8 FILLER_44_457 ();
 sg13g2_decap_8 FILLER_44_464 ();
 sg13g2_decap_8 FILLER_44_475 ();
 sg13g2_decap_8 FILLER_44_482 ();
 sg13g2_decap_8 FILLER_44_489 ();
 sg13g2_decap_8 FILLER_44_496 ();
 sg13g2_decap_8 FILLER_44_503 ();
 sg13g2_decap_8 FILLER_44_510 ();
 sg13g2_fill_2 FILLER_44_517 ();
 sg13g2_decap_4 FILLER_44_524 ();
 sg13g2_decap_4 FILLER_44_537 ();
 sg13g2_fill_1 FILLER_44_541 ();
 sg13g2_decap_4 FILLER_44_546 ();
 sg13g2_fill_1 FILLER_44_550 ();
 sg13g2_decap_8 FILLER_44_560 ();
 sg13g2_decap_8 FILLER_44_567 ();
 sg13g2_decap_8 FILLER_44_574 ();
 sg13g2_decap_8 FILLER_44_581 ();
 sg13g2_decap_4 FILLER_44_594 ();
 sg13g2_fill_2 FILLER_44_598 ();
 sg13g2_decap_8 FILLER_44_606 ();
 sg13g2_decap_8 FILLER_44_613 ();
 sg13g2_decap_8 FILLER_44_620 ();
 sg13g2_fill_2 FILLER_44_627 ();
 sg13g2_fill_2 FILLER_44_633 ();
 sg13g2_fill_1 FILLER_44_635 ();
 sg13g2_decap_4 FILLER_44_641 ();
 sg13g2_decap_8 FILLER_44_649 ();
 sg13g2_decap_4 FILLER_44_660 ();
 sg13g2_fill_1 FILLER_44_669 ();
 sg13g2_fill_2 FILLER_44_675 ();
 sg13g2_fill_1 FILLER_44_684 ();
 sg13g2_decap_8 FILLER_44_689 ();
 sg13g2_fill_2 FILLER_44_700 ();
 sg13g2_fill_1 FILLER_44_702 ();
 sg13g2_decap_4 FILLER_44_707 ();
 sg13g2_decap_4 FILLER_44_721 ();
 sg13g2_fill_2 FILLER_44_725 ();
 sg13g2_fill_2 FILLER_44_731 ();
 sg13g2_fill_1 FILLER_44_733 ();
 sg13g2_decap_4 FILLER_44_738 ();
 sg13g2_decap_8 FILLER_44_751 ();
 sg13g2_decap_8 FILLER_44_758 ();
 sg13g2_decap_8 FILLER_44_765 ();
 sg13g2_decap_8 FILLER_44_772 ();
 sg13g2_decap_8 FILLER_44_779 ();
 sg13g2_decap_8 FILLER_44_786 ();
 sg13g2_decap_8 FILLER_44_793 ();
 sg13g2_decap_8 FILLER_44_800 ();
 sg13g2_decap_8 FILLER_44_807 ();
 sg13g2_decap_8 FILLER_44_814 ();
 sg13g2_decap_8 FILLER_44_821 ();
 sg13g2_decap_8 FILLER_44_828 ();
 sg13g2_decap_8 FILLER_44_835 ();
 sg13g2_decap_8 FILLER_44_842 ();
 sg13g2_decap_8 FILLER_44_849 ();
 sg13g2_decap_8 FILLER_44_856 ();
 sg13g2_decap_8 FILLER_44_863 ();
 sg13g2_decap_8 FILLER_44_870 ();
 sg13g2_fill_1 FILLER_44_877 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_4 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_67 ();
 sg13g2_decap_4 FILLER_45_74 ();
 sg13g2_fill_1 FILLER_45_78 ();
 sg13g2_decap_8 FILLER_45_88 ();
 sg13g2_fill_2 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_104 ();
 sg13g2_fill_1 FILLER_45_106 ();
 sg13g2_decap_8 FILLER_45_113 ();
 sg13g2_fill_2 FILLER_45_120 ();
 sg13g2_fill_1 FILLER_45_122 ();
 sg13g2_decap_4 FILLER_45_127 ();
 sg13g2_fill_2 FILLER_45_131 ();
 sg13g2_decap_4 FILLER_45_137 ();
 sg13g2_fill_2 FILLER_45_141 ();
 sg13g2_fill_1 FILLER_45_147 ();
 sg13g2_fill_1 FILLER_45_153 ();
 sg13g2_fill_1 FILLER_45_166 ();
 sg13g2_fill_1 FILLER_45_171 ();
 sg13g2_fill_1 FILLER_45_177 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_4 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_197 ();
 sg13g2_fill_2 FILLER_45_204 ();
 sg13g2_fill_1 FILLER_45_206 ();
 sg13g2_decap_4 FILLER_45_218 ();
 sg13g2_fill_2 FILLER_45_222 ();
 sg13g2_decap_8 FILLER_45_229 ();
 sg13g2_decap_8 FILLER_45_236 ();
 sg13g2_decap_8 FILLER_45_243 ();
 sg13g2_decap_4 FILLER_45_250 ();
 sg13g2_decap_4 FILLER_45_259 ();
 sg13g2_decap_4 FILLER_45_267 ();
 sg13g2_fill_2 FILLER_45_276 ();
 sg13g2_fill_1 FILLER_45_298 ();
 sg13g2_fill_1 FILLER_45_303 ();
 sg13g2_decap_8 FILLER_45_310 ();
 sg13g2_decap_4 FILLER_45_317 ();
 sg13g2_fill_2 FILLER_45_324 ();
 sg13g2_fill_1 FILLER_45_326 ();
 sg13g2_decap_8 FILLER_45_331 ();
 sg13g2_decap_8 FILLER_45_338 ();
 sg13g2_decap_8 FILLER_45_345 ();
 sg13g2_fill_2 FILLER_45_352 ();
 sg13g2_decap_8 FILLER_45_359 ();
 sg13g2_decap_8 FILLER_45_366 ();
 sg13g2_decap_8 FILLER_45_373 ();
 sg13g2_decap_4 FILLER_45_380 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_422 ();
 sg13g2_fill_2 FILLER_45_429 ();
 sg13g2_fill_1 FILLER_45_431 ();
 sg13g2_decap_8 FILLER_45_442 ();
 sg13g2_decap_8 FILLER_45_449 ();
 sg13g2_decap_8 FILLER_45_456 ();
 sg13g2_decap_8 FILLER_45_463 ();
 sg13g2_decap_8 FILLER_45_470 ();
 sg13g2_decap_8 FILLER_45_477 ();
 sg13g2_decap_8 FILLER_45_484 ();
 sg13g2_decap_4 FILLER_45_491 ();
 sg13g2_fill_2 FILLER_45_505 ();
 sg13g2_fill_1 FILLER_45_507 ();
 sg13g2_fill_1 FILLER_45_516 ();
 sg13g2_decap_8 FILLER_45_521 ();
 sg13g2_decap_8 FILLER_45_533 ();
 sg13g2_decap_4 FILLER_45_540 ();
 sg13g2_fill_1 FILLER_45_557 ();
 sg13g2_decap_8 FILLER_45_562 ();
 sg13g2_decap_8 FILLER_45_569 ();
 sg13g2_fill_1 FILLER_45_576 ();
 sg13g2_decap_8 FILLER_45_582 ();
 sg13g2_decap_8 FILLER_45_589 ();
 sg13g2_decap_4 FILLER_45_596 ();
 sg13g2_fill_1 FILLER_45_600 ();
 sg13g2_decap_4 FILLER_45_605 ();
 sg13g2_decap_8 FILLER_45_619 ();
 sg13g2_decap_4 FILLER_45_626 ();
 sg13g2_fill_1 FILLER_45_630 ();
 sg13g2_decap_8 FILLER_45_637 ();
 sg13g2_decap_8 FILLER_45_644 ();
 sg13g2_decap_4 FILLER_45_651 ();
 sg13g2_fill_2 FILLER_45_660 ();
 sg13g2_fill_1 FILLER_45_662 ();
 sg13g2_fill_2 FILLER_45_668 ();
 sg13g2_decap_8 FILLER_45_676 ();
 sg13g2_fill_1 FILLER_45_683 ();
 sg13g2_fill_2 FILLER_45_696 ();
 sg13g2_decap_8 FILLER_45_704 ();
 sg13g2_decap_4 FILLER_45_714 ();
 sg13g2_decap_4 FILLER_45_721 ();
 sg13g2_decap_4 FILLER_45_729 ();
 sg13g2_fill_1 FILLER_45_733 ();
 sg13g2_fill_1 FILLER_45_738 ();
 sg13g2_decap_8 FILLER_45_744 ();
 sg13g2_decap_8 FILLER_45_751 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_774 ();
 sg13g2_decap_8 FILLER_45_781 ();
 sg13g2_decap_8 FILLER_45_788 ();
 sg13g2_decap_8 FILLER_45_795 ();
 sg13g2_decap_8 FILLER_45_802 ();
 sg13g2_decap_8 FILLER_45_809 ();
 sg13g2_decap_8 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_823 ();
 sg13g2_decap_8 FILLER_45_830 ();
 sg13g2_decap_8 FILLER_45_837 ();
 sg13g2_decap_8 FILLER_45_844 ();
 sg13g2_decap_8 FILLER_45_851 ();
 sg13g2_decap_8 FILLER_45_858 ();
 sg13g2_decap_8 FILLER_45_865 ();
 sg13g2_decap_4 FILLER_45_872 ();
 sg13g2_fill_2 FILLER_45_876 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_fill_1 FILLER_46_81 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_4 FILLER_46_119 ();
 sg13g2_decap_4 FILLER_46_128 ();
 sg13g2_decap_8 FILLER_46_146 ();
 sg13g2_decap_8 FILLER_46_171 ();
 sg13g2_decap_8 FILLER_46_178 ();
 sg13g2_decap_8 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_192 ();
 sg13g2_decap_4 FILLER_46_199 ();
 sg13g2_fill_2 FILLER_46_203 ();
 sg13g2_fill_2 FILLER_46_210 ();
 sg13g2_decap_4 FILLER_46_217 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_decap_8 FILLER_46_227 ();
 sg13g2_decap_8 FILLER_46_234 ();
 sg13g2_decap_8 FILLER_46_241 ();
 sg13g2_decap_8 FILLER_46_248 ();
 sg13g2_decap_8 FILLER_46_255 ();
 sg13g2_fill_1 FILLER_46_262 ();
 sg13g2_decap_8 FILLER_46_267 ();
 sg13g2_decap_4 FILLER_46_274 ();
 sg13g2_fill_2 FILLER_46_278 ();
 sg13g2_decap_4 FILLER_46_284 ();
 sg13g2_fill_1 FILLER_46_288 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_fill_1 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_331 ();
 sg13g2_fill_2 FILLER_46_338 ();
 sg13g2_decap_8 FILLER_46_345 ();
 sg13g2_decap_8 FILLER_46_352 ();
 sg13g2_decap_8 FILLER_46_359 ();
 sg13g2_decap_8 FILLER_46_366 ();
 sg13g2_decap_4 FILLER_46_378 ();
 sg13g2_fill_1 FILLER_46_382 ();
 sg13g2_fill_1 FILLER_46_391 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_decap_8 FILLER_46_403 ();
 sg13g2_decap_8 FILLER_46_410 ();
 sg13g2_decap_8 FILLER_46_417 ();
 sg13g2_decap_8 FILLER_46_424 ();
 sg13g2_fill_2 FILLER_46_431 ();
 sg13g2_fill_1 FILLER_46_433 ();
 sg13g2_decap_4 FILLER_46_439 ();
 sg13g2_fill_1 FILLER_46_443 ();
 sg13g2_decap_8 FILLER_46_463 ();
 sg13g2_decap_8 FILLER_46_470 ();
 sg13g2_decap_8 FILLER_46_477 ();
 sg13g2_decap_4 FILLER_46_484 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_fill_2 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_fill_2 FILLER_46_546 ();
 sg13g2_fill_1 FILLER_46_548 ();
 sg13g2_decap_4 FILLER_46_555 ();
 sg13g2_fill_1 FILLER_46_559 ();
 sg13g2_fill_1 FILLER_46_565 ();
 sg13g2_fill_2 FILLER_46_571 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_fill_1 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_605 ();
 sg13g2_fill_1 FILLER_46_612 ();
 sg13g2_decap_4 FILLER_46_623 ();
 sg13g2_decap_4 FILLER_46_632 ();
 sg13g2_fill_2 FILLER_46_641 ();
 sg13g2_fill_1 FILLER_46_643 ();
 sg13g2_fill_1 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_664 ();
 sg13g2_decap_8 FILLER_46_671 ();
 sg13g2_decap_8 FILLER_46_678 ();
 sg13g2_decap_8 FILLER_46_685 ();
 sg13g2_decap_8 FILLER_46_692 ();
 sg13g2_decap_8 FILLER_46_699 ();
 sg13g2_decap_8 FILLER_46_710 ();
 sg13g2_decap_8 FILLER_46_717 ();
 sg13g2_decap_8 FILLER_46_724 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_738 ();
 sg13g2_decap_4 FILLER_46_745 ();
 sg13g2_fill_2 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_755 ();
 sg13g2_decap_8 FILLER_46_762 ();
 sg13g2_decap_8 FILLER_46_769 ();
 sg13g2_decap_8 FILLER_46_776 ();
 sg13g2_decap_8 FILLER_46_783 ();
 sg13g2_decap_8 FILLER_46_790 ();
 sg13g2_decap_8 FILLER_46_797 ();
 sg13g2_decap_8 FILLER_46_804 ();
 sg13g2_decap_8 FILLER_46_811 ();
 sg13g2_decap_8 FILLER_46_818 ();
 sg13g2_decap_8 FILLER_46_825 ();
 sg13g2_decap_8 FILLER_46_832 ();
 sg13g2_decap_8 FILLER_46_839 ();
 sg13g2_decap_8 FILLER_46_846 ();
 sg13g2_decap_8 FILLER_46_853 ();
 sg13g2_decap_8 FILLER_46_860 ();
 sg13g2_decap_8 FILLER_46_867 ();
 sg13g2_decap_4 FILLER_46_874 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_fill_2 FILLER_47_56 ();
 sg13g2_fill_1 FILLER_47_58 ();
 sg13g2_decap_4 FILLER_47_63 ();
 sg13g2_fill_1 FILLER_47_67 ();
 sg13g2_fill_2 FILLER_47_82 ();
 sg13g2_decap_8 FILLER_47_89 ();
 sg13g2_fill_2 FILLER_47_96 ();
 sg13g2_decap_4 FILLER_47_103 ();
 sg13g2_decap_4 FILLER_47_111 ();
 sg13g2_fill_1 FILLER_47_115 ();
 sg13g2_decap_8 FILLER_47_124 ();
 sg13g2_decap_8 FILLER_47_131 ();
 sg13g2_decap_4 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_142 ();
 sg13g2_fill_1 FILLER_47_148 ();
 sg13g2_decap_8 FILLER_47_157 ();
 sg13g2_decap_4 FILLER_47_164 ();
 sg13g2_fill_2 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_179 ();
 sg13g2_decap_8 FILLER_47_186 ();
 sg13g2_decap_8 FILLER_47_200 ();
 sg13g2_decap_8 FILLER_47_207 ();
 sg13g2_decap_8 FILLER_47_214 ();
 sg13g2_fill_1 FILLER_47_221 ();
 sg13g2_decap_8 FILLER_47_230 ();
 sg13g2_decap_8 FILLER_47_237 ();
 sg13g2_decap_8 FILLER_47_244 ();
 sg13g2_decap_8 FILLER_47_251 ();
 sg13g2_decap_4 FILLER_47_258 ();
 sg13g2_decap_8 FILLER_47_278 ();
 sg13g2_decap_8 FILLER_47_285 ();
 sg13g2_decap_8 FILLER_47_292 ();
 sg13g2_decap_4 FILLER_47_315 ();
 sg13g2_fill_1 FILLER_47_319 ();
 sg13g2_decap_8 FILLER_47_327 ();
 sg13g2_decap_4 FILLER_47_334 ();
 sg13g2_fill_2 FILLER_47_338 ();
 sg13g2_decap_8 FILLER_47_349 ();
 sg13g2_decap_8 FILLER_47_356 ();
 sg13g2_decap_8 FILLER_47_363 ();
 sg13g2_decap_8 FILLER_47_370 ();
 sg13g2_decap_8 FILLER_47_377 ();
 sg13g2_decap_8 FILLER_47_384 ();
 sg13g2_decap_8 FILLER_47_396 ();
 sg13g2_decap_8 FILLER_47_403 ();
 sg13g2_decap_4 FILLER_47_410 ();
 sg13g2_fill_2 FILLER_47_414 ();
 sg13g2_decap_8 FILLER_47_421 ();
 sg13g2_decap_8 FILLER_47_433 ();
 sg13g2_decap_8 FILLER_47_440 ();
 sg13g2_decap_8 FILLER_47_447 ();
 sg13g2_decap_8 FILLER_47_454 ();
 sg13g2_decap_4 FILLER_47_461 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_4 FILLER_47_483 ();
 sg13g2_fill_2 FILLER_47_487 ();
 sg13g2_decap_8 FILLER_47_498 ();
 sg13g2_fill_1 FILLER_47_505 ();
 sg13g2_decap_8 FILLER_47_512 ();
 sg13g2_fill_2 FILLER_47_519 ();
 sg13g2_fill_1 FILLER_47_521 ();
 sg13g2_decap_4 FILLER_47_536 ();
 sg13g2_decap_4 FILLER_47_548 ();
 sg13g2_fill_2 FILLER_47_552 ();
 sg13g2_decap_4 FILLER_47_566 ();
 sg13g2_fill_1 FILLER_47_570 ();
 sg13g2_decap_8 FILLER_47_576 ();
 sg13g2_decap_8 FILLER_47_583 ();
 sg13g2_decap_8 FILLER_47_590 ();
 sg13g2_fill_1 FILLER_47_597 ();
 sg13g2_fill_2 FILLER_47_604 ();
 sg13g2_fill_1 FILLER_47_606 ();
 sg13g2_decap_4 FILLER_47_612 ();
 sg13g2_decap_8 FILLER_47_621 ();
 sg13g2_decap_8 FILLER_47_628 ();
 sg13g2_decap_8 FILLER_47_635 ();
 sg13g2_decap_4 FILLER_47_654 ();
 sg13g2_decap_8 FILLER_47_662 ();
 sg13g2_decap_8 FILLER_47_669 ();
 sg13g2_decap_4 FILLER_47_685 ();
 sg13g2_decap_8 FILLER_47_694 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_4 FILLER_47_718 ();
 sg13g2_fill_2 FILLER_47_722 ();
 sg13g2_fill_1 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_734 ();
 sg13g2_decap_8 FILLER_47_741 ();
 sg13g2_decap_4 FILLER_47_748 ();
 sg13g2_fill_2 FILLER_47_761 ();
 sg13g2_fill_1 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_768 ();
 sg13g2_decap_8 FILLER_47_775 ();
 sg13g2_decap_8 FILLER_47_782 ();
 sg13g2_decap_8 FILLER_47_789 ();
 sg13g2_decap_8 FILLER_47_796 ();
 sg13g2_decap_8 FILLER_47_803 ();
 sg13g2_decap_8 FILLER_47_810 ();
 sg13g2_decap_8 FILLER_47_817 ();
 sg13g2_decap_8 FILLER_47_824 ();
 sg13g2_decap_8 FILLER_47_831 ();
 sg13g2_decap_8 FILLER_47_838 ();
 sg13g2_decap_8 FILLER_47_845 ();
 sg13g2_decap_8 FILLER_47_852 ();
 sg13g2_decap_8 FILLER_47_859 ();
 sg13g2_decap_8 FILLER_47_866 ();
 sg13g2_decap_4 FILLER_47_873 ();
 sg13g2_fill_1 FILLER_47_877 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_4 FILLER_48_56 ();
 sg13g2_decap_4 FILLER_48_64 ();
 sg13g2_fill_2 FILLER_48_68 ();
 sg13g2_decap_8 FILLER_48_86 ();
 sg13g2_decap_8 FILLER_48_93 ();
 sg13g2_fill_2 FILLER_48_100 ();
 sg13g2_fill_1 FILLER_48_102 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_129 ();
 sg13g2_fill_2 FILLER_48_136 ();
 sg13g2_fill_1 FILLER_48_138 ();
 sg13g2_decap_4 FILLER_48_144 ();
 sg13g2_fill_1 FILLER_48_148 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_fill_1 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_172 ();
 sg13g2_decap_8 FILLER_48_179 ();
 sg13g2_decap_8 FILLER_48_186 ();
 sg13g2_decap_8 FILLER_48_193 ();
 sg13g2_fill_2 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_202 ();
 sg13g2_decap_8 FILLER_48_212 ();
 sg13g2_decap_8 FILLER_48_219 ();
 sg13g2_decap_8 FILLER_48_226 ();
 sg13g2_decap_8 FILLER_48_233 ();
 sg13g2_fill_2 FILLER_48_245 ();
 sg13g2_decap_4 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_260 ();
 sg13g2_decap_4 FILLER_48_265 ();
 sg13g2_fill_1 FILLER_48_269 ();
 sg13g2_decap_8 FILLER_48_278 ();
 sg13g2_decap_4 FILLER_48_285 ();
 sg13g2_fill_2 FILLER_48_289 ();
 sg13g2_decap_4 FILLER_48_297 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_decap_4 FILLER_48_317 ();
 sg13g2_fill_2 FILLER_48_321 ();
 sg13g2_decap_4 FILLER_48_333 ();
 sg13g2_decap_8 FILLER_48_342 ();
 sg13g2_decap_8 FILLER_48_349 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_4 FILLER_48_363 ();
 sg13g2_decap_4 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_379 ();
 sg13g2_fill_2 FILLER_48_386 ();
 sg13g2_decap_4 FILLER_48_394 ();
 sg13g2_decap_4 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_48_415 ();
 sg13g2_decap_4 FILLER_48_422 ();
 sg13g2_fill_1 FILLER_48_426 ();
 sg13g2_decap_4 FILLER_48_433 ();
 sg13g2_fill_2 FILLER_48_437 ();
 sg13g2_decap_8 FILLER_48_449 ();
 sg13g2_decap_8 FILLER_48_456 ();
 sg13g2_fill_1 FILLER_48_463 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_fill_1 FILLER_48_476 ();
 sg13g2_decap_4 FILLER_48_481 ();
 sg13g2_decap_8 FILLER_48_492 ();
 sg13g2_fill_2 FILLER_48_499 ();
 sg13g2_decap_8 FILLER_48_510 ();
 sg13g2_decap_4 FILLER_48_517 ();
 sg13g2_decap_4 FILLER_48_524 ();
 sg13g2_fill_1 FILLER_48_528 ();
 sg13g2_decap_4 FILLER_48_538 ();
 sg13g2_decap_8 FILLER_48_547 ();
 sg13g2_decap_4 FILLER_48_554 ();
 sg13g2_decap_4 FILLER_48_562 ();
 sg13g2_fill_1 FILLER_48_566 ();
 sg13g2_decap_8 FILLER_48_575 ();
 sg13g2_decap_4 FILLER_48_582 ();
 sg13g2_fill_2 FILLER_48_586 ();
 sg13g2_decap_8 FILLER_48_593 ();
 sg13g2_fill_2 FILLER_48_600 ();
 sg13g2_decap_8 FILLER_48_617 ();
 sg13g2_decap_8 FILLER_48_624 ();
 sg13g2_decap_8 FILLER_48_631 ();
 sg13g2_fill_1 FILLER_48_642 ();
 sg13g2_decap_8 FILLER_48_648 ();
 sg13g2_fill_2 FILLER_48_655 ();
 sg13g2_fill_1 FILLER_48_657 ();
 sg13g2_decap_4 FILLER_48_666 ();
 sg13g2_fill_2 FILLER_48_670 ();
 sg13g2_fill_2 FILLER_48_677 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_4 FILLER_48_700 ();
 sg13g2_fill_2 FILLER_48_704 ();
 sg13g2_decap_8 FILLER_48_724 ();
 sg13g2_decap_8 FILLER_48_731 ();
 sg13g2_fill_2 FILLER_48_738 ();
 sg13g2_fill_1 FILLER_48_740 ();
 sg13g2_fill_2 FILLER_48_751 ();
 sg13g2_fill_1 FILLER_48_753 ();
 sg13g2_decap_4 FILLER_48_758 ();
 sg13g2_fill_1 FILLER_48_762 ();
 sg13g2_decap_8 FILLER_48_769 ();
 sg13g2_decap_8 FILLER_48_776 ();
 sg13g2_decap_8 FILLER_48_783 ();
 sg13g2_decap_8 FILLER_48_790 ();
 sg13g2_decap_8 FILLER_48_797 ();
 sg13g2_decap_8 FILLER_48_804 ();
 sg13g2_decap_8 FILLER_48_811 ();
 sg13g2_decap_8 FILLER_48_818 ();
 sg13g2_decap_8 FILLER_48_825 ();
 sg13g2_decap_8 FILLER_48_832 ();
 sg13g2_decap_8 FILLER_48_839 ();
 sg13g2_decap_8 FILLER_48_846 ();
 sg13g2_decap_8 FILLER_48_853 ();
 sg13g2_decap_8 FILLER_48_860 ();
 sg13g2_decap_8 FILLER_48_867 ();
 sg13g2_decap_4 FILLER_48_874 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_4 FILLER_49_56 ();
 sg13g2_fill_1 FILLER_49_60 ();
 sg13g2_decap_4 FILLER_49_65 ();
 sg13g2_fill_1 FILLER_49_69 ();
 sg13g2_decap_4 FILLER_49_79 ();
 sg13g2_fill_1 FILLER_49_83 ();
 sg13g2_decap_8 FILLER_49_89 ();
 sg13g2_decap_4 FILLER_49_96 ();
 sg13g2_fill_2 FILLER_49_100 ();
 sg13g2_decap_8 FILLER_49_106 ();
 sg13g2_fill_1 FILLER_49_113 ();
 sg13g2_fill_1 FILLER_49_123 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_fill_2 FILLER_49_140 ();
 sg13g2_fill_1 FILLER_49_142 ();
 sg13g2_decap_8 FILLER_49_152 ();
 sg13g2_decap_8 FILLER_49_159 ();
 sg13g2_fill_1 FILLER_49_166 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_4 FILLER_49_179 ();
 sg13g2_decap_8 FILLER_49_192 ();
 sg13g2_fill_2 FILLER_49_218 ();
 sg13g2_decap_8 FILLER_49_225 ();
 sg13g2_decap_4 FILLER_49_232 ();
 sg13g2_fill_1 FILLER_49_236 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_256 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_fill_2 FILLER_49_277 ();
 sg13g2_decap_8 FILLER_49_284 ();
 sg13g2_decap_4 FILLER_49_291 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_decap_4 FILLER_49_305 ();
 sg13g2_fill_1 FILLER_49_309 ();
 sg13g2_decap_8 FILLER_49_320 ();
 sg13g2_decap_4 FILLER_49_327 ();
 sg13g2_fill_2 FILLER_49_331 ();
 sg13g2_decap_4 FILLER_49_337 ();
 sg13g2_fill_2 FILLER_49_341 ();
 sg13g2_decap_4 FILLER_49_348 ();
 sg13g2_fill_1 FILLER_49_352 ();
 sg13g2_decap_8 FILLER_49_359 ();
 sg13g2_decap_4 FILLER_49_366 ();
 sg13g2_decap_8 FILLER_49_376 ();
 sg13g2_decap_4 FILLER_49_383 ();
 sg13g2_fill_1 FILLER_49_387 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_411 ();
 sg13g2_decap_4 FILLER_49_418 ();
 sg13g2_fill_2 FILLER_49_426 ();
 sg13g2_fill_1 FILLER_49_428 ();
 sg13g2_decap_4 FILLER_49_434 ();
 sg13g2_fill_2 FILLER_49_438 ();
 sg13g2_decap_8 FILLER_49_450 ();
 sg13g2_fill_2 FILLER_49_457 ();
 sg13g2_decap_8 FILLER_49_464 ();
 sg13g2_decap_4 FILLER_49_471 ();
 sg13g2_fill_2 FILLER_49_475 ();
 sg13g2_decap_8 FILLER_49_482 ();
 sg13g2_decap_8 FILLER_49_489 ();
 sg13g2_decap_8 FILLER_49_496 ();
 sg13g2_decap_8 FILLER_49_503 ();
 sg13g2_decap_4 FILLER_49_510 ();
 sg13g2_fill_1 FILLER_49_514 ();
 sg13g2_decap_8 FILLER_49_520 ();
 sg13g2_decap_4 FILLER_49_527 ();
 sg13g2_fill_2 FILLER_49_531 ();
 sg13g2_decap_8 FILLER_49_542 ();
 sg13g2_fill_2 FILLER_49_549 ();
 sg13g2_fill_1 FILLER_49_551 ();
 sg13g2_decap_4 FILLER_49_555 ();
 sg13g2_fill_2 FILLER_49_559 ();
 sg13g2_decap_8 FILLER_49_580 ();
 sg13g2_decap_8 FILLER_49_587 ();
 sg13g2_decap_4 FILLER_49_594 ();
 sg13g2_fill_1 FILLER_49_598 ();
 sg13g2_decap_8 FILLER_49_614 ();
 sg13g2_decap_8 FILLER_49_621 ();
 sg13g2_decap_8 FILLER_49_628 ();
 sg13g2_decap_4 FILLER_49_635 ();
 sg13g2_decap_8 FILLER_49_642 ();
 sg13g2_fill_2 FILLER_49_649 ();
 sg13g2_fill_1 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_fill_1 FILLER_49_672 ();
 sg13g2_fill_2 FILLER_49_678 ();
 sg13g2_fill_1 FILLER_49_680 ();
 sg13g2_fill_2 FILLER_49_684 ();
 sg13g2_decap_8 FILLER_49_691 ();
 sg13g2_decap_4 FILLER_49_698 ();
 sg13g2_fill_2 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_fill_1 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_738 ();
 sg13g2_decap_8 FILLER_49_745 ();
 sg13g2_fill_2 FILLER_49_752 ();
 sg13g2_decap_8 FILLER_49_760 ();
 sg13g2_decap_8 FILLER_49_767 ();
 sg13g2_decap_8 FILLER_49_774 ();
 sg13g2_decap_8 FILLER_49_781 ();
 sg13g2_decap_8 FILLER_49_788 ();
 sg13g2_decap_8 FILLER_49_795 ();
 sg13g2_decap_8 FILLER_49_802 ();
 sg13g2_decap_8 FILLER_49_809 ();
 sg13g2_decap_8 FILLER_49_816 ();
 sg13g2_decap_8 FILLER_49_823 ();
 sg13g2_decap_8 FILLER_49_830 ();
 sg13g2_decap_8 FILLER_49_837 ();
 sg13g2_decap_8 FILLER_49_844 ();
 sg13g2_decap_8 FILLER_49_851 ();
 sg13g2_decap_8 FILLER_49_858 ();
 sg13g2_decap_8 FILLER_49_865 ();
 sg13g2_decap_4 FILLER_49_872 ();
 sg13g2_fill_2 FILLER_49_876 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_68 ();
 sg13g2_decap_4 FILLER_50_75 ();
 sg13g2_fill_1 FILLER_50_79 ();
 sg13g2_decap_8 FILLER_50_90 ();
 sg13g2_decap_8 FILLER_50_97 ();
 sg13g2_decap_4 FILLER_50_104 ();
 sg13g2_fill_1 FILLER_50_108 ();
 sg13g2_decap_4 FILLER_50_113 ();
 sg13g2_fill_1 FILLER_50_117 ();
 sg13g2_decap_8 FILLER_50_131 ();
 sg13g2_decap_4 FILLER_50_138 ();
 sg13g2_fill_2 FILLER_50_147 ();
 sg13g2_fill_1 FILLER_50_149 ();
 sg13g2_decap_4 FILLER_50_167 ();
 sg13g2_fill_2 FILLER_50_171 ();
 sg13g2_decap_4 FILLER_50_184 ();
 sg13g2_decap_8 FILLER_50_193 ();
 sg13g2_decap_8 FILLER_50_200 ();
 sg13g2_decap_8 FILLER_50_207 ();
 sg13g2_decap_4 FILLER_50_214 ();
 sg13g2_fill_2 FILLER_50_218 ();
 sg13g2_fill_2 FILLER_50_224 ();
 sg13g2_fill_1 FILLER_50_226 ();
 sg13g2_decap_8 FILLER_50_236 ();
 sg13g2_decap_4 FILLER_50_243 ();
 sg13g2_decap_8 FILLER_50_252 ();
 sg13g2_decap_8 FILLER_50_259 ();
 sg13g2_decap_4 FILLER_50_266 ();
 sg13g2_fill_2 FILLER_50_270 ();
 sg13g2_decap_8 FILLER_50_276 ();
 sg13g2_decap_8 FILLER_50_283 ();
 sg13g2_decap_4 FILLER_50_290 ();
 sg13g2_fill_2 FILLER_50_294 ();
 sg13g2_decap_8 FILLER_50_301 ();
 sg13g2_decap_4 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_322 ();
 sg13g2_decap_8 FILLER_50_329 ();
 sg13g2_decap_8 FILLER_50_336 ();
 sg13g2_decap_8 FILLER_50_343 ();
 sg13g2_decap_8 FILLER_50_350 ();
 sg13g2_decap_8 FILLER_50_357 ();
 sg13g2_decap_4 FILLER_50_364 ();
 sg13g2_fill_1 FILLER_50_368 ();
 sg13g2_decap_4 FILLER_50_374 ();
 sg13g2_fill_2 FILLER_50_378 ();
 sg13g2_decap_8 FILLER_50_388 ();
 sg13g2_decap_8 FILLER_50_395 ();
 sg13g2_fill_2 FILLER_50_402 ();
 sg13g2_decap_4 FILLER_50_413 ();
 sg13g2_fill_1 FILLER_50_417 ();
 sg13g2_fill_2 FILLER_50_423 ();
 sg13g2_fill_1 FILLER_50_425 ();
 sg13g2_decap_4 FILLER_50_431 ();
 sg13g2_decap_8 FILLER_50_439 ();
 sg13g2_decap_8 FILLER_50_446 ();
 sg13g2_decap_8 FILLER_50_453 ();
 sg13g2_decap_8 FILLER_50_460 ();
 sg13g2_decap_4 FILLER_50_467 ();
 sg13g2_fill_2 FILLER_50_471 ();
 sg13g2_fill_2 FILLER_50_480 ();
 sg13g2_fill_1 FILLER_50_486 ();
 sg13g2_decap_4 FILLER_50_492 ();
 sg13g2_fill_2 FILLER_50_496 ();
 sg13g2_decap_8 FILLER_50_503 ();
 sg13g2_decap_8 FILLER_50_510 ();
 sg13g2_decap_8 FILLER_50_517 ();
 sg13g2_fill_2 FILLER_50_524 ();
 sg13g2_decap_4 FILLER_50_531 ();
 sg13g2_decap_8 FILLER_50_540 ();
 sg13g2_decap_8 FILLER_50_547 ();
 sg13g2_decap_8 FILLER_50_554 ();
 sg13g2_decap_8 FILLER_50_561 ();
 sg13g2_decap_4 FILLER_50_578 ();
 sg13g2_decap_8 FILLER_50_587 ();
 sg13g2_decap_8 FILLER_50_594 ();
 sg13g2_fill_2 FILLER_50_601 ();
 sg13g2_fill_1 FILLER_50_603 ();
 sg13g2_decap_4 FILLER_50_608 ();
 sg13g2_fill_2 FILLER_50_612 ();
 sg13g2_decap_8 FILLER_50_624 ();
 sg13g2_fill_2 FILLER_50_631 ();
 sg13g2_decap_4 FILLER_50_637 ();
 sg13g2_fill_2 FILLER_50_641 ();
 sg13g2_fill_1 FILLER_50_649 ();
 sg13g2_decap_4 FILLER_50_655 ();
 sg13g2_decap_8 FILLER_50_667 ();
 sg13g2_decap_8 FILLER_50_674 ();
 sg13g2_decap_8 FILLER_50_681 ();
 sg13g2_decap_8 FILLER_50_688 ();
 sg13g2_decap_8 FILLER_50_695 ();
 sg13g2_decap_4 FILLER_50_702 ();
 sg13g2_fill_2 FILLER_50_706 ();
 sg13g2_fill_2 FILLER_50_712 ();
 sg13g2_decap_4 FILLER_50_740 ();
 sg13g2_fill_1 FILLER_50_748 ();
 sg13g2_decap_8 FILLER_50_753 ();
 sg13g2_decap_8 FILLER_50_760 ();
 sg13g2_decap_8 FILLER_50_767 ();
 sg13g2_decap_8 FILLER_50_774 ();
 sg13g2_decap_8 FILLER_50_781 ();
 sg13g2_decap_8 FILLER_50_788 ();
 sg13g2_decap_8 FILLER_50_795 ();
 sg13g2_decap_8 FILLER_50_802 ();
 sg13g2_decap_8 FILLER_50_809 ();
 sg13g2_decap_8 FILLER_50_816 ();
 sg13g2_decap_8 FILLER_50_823 ();
 sg13g2_decap_8 FILLER_50_830 ();
 sg13g2_decap_8 FILLER_50_837 ();
 sg13g2_decap_8 FILLER_50_844 ();
 sg13g2_decap_8 FILLER_50_851 ();
 sg13g2_decap_8 FILLER_50_858 ();
 sg13g2_decap_8 FILLER_50_865 ();
 sg13g2_decap_4 FILLER_50_872 ();
 sg13g2_fill_2 FILLER_50_876 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_55 ();
 sg13g2_decap_8 FILLER_51_62 ();
 sg13g2_decap_8 FILLER_51_69 ();
 sg13g2_decap_4 FILLER_51_76 ();
 sg13g2_fill_2 FILLER_51_80 ();
 sg13g2_decap_4 FILLER_51_86 ();
 sg13g2_fill_1 FILLER_51_90 ();
 sg13g2_decap_8 FILLER_51_95 ();
 sg13g2_fill_1 FILLER_51_102 ();
 sg13g2_fill_2 FILLER_51_108 ();
 sg13g2_decap_4 FILLER_51_124 ();
 sg13g2_fill_1 FILLER_51_128 ();
 sg13g2_fill_2 FILLER_51_134 ();
 sg13g2_decap_4 FILLER_51_140 ();
 sg13g2_fill_1 FILLER_51_144 ();
 sg13g2_fill_2 FILLER_51_150 ();
 sg13g2_decap_8 FILLER_51_157 ();
 sg13g2_decap_4 FILLER_51_164 ();
 sg13g2_fill_1 FILLER_51_168 ();
 sg13g2_fill_2 FILLER_51_179 ();
 sg13g2_decap_8 FILLER_51_190 ();
 sg13g2_decap_4 FILLER_51_197 ();
 sg13g2_decap_4 FILLER_51_208 ();
 sg13g2_fill_1 FILLER_51_212 ();
 sg13g2_decap_8 FILLER_51_222 ();
 sg13g2_decap_8 FILLER_51_229 ();
 sg13g2_decap_8 FILLER_51_236 ();
 sg13g2_decap_8 FILLER_51_247 ();
 sg13g2_decap_4 FILLER_51_254 ();
 sg13g2_decap_4 FILLER_51_263 ();
 sg13g2_fill_1 FILLER_51_267 ();
 sg13g2_decap_8 FILLER_51_277 ();
 sg13g2_decap_8 FILLER_51_284 ();
 sg13g2_decap_4 FILLER_51_291 ();
 sg13g2_decap_8 FILLER_51_304 ();
 sg13g2_decap_8 FILLER_51_311 ();
 sg13g2_decap_8 FILLER_51_318 ();
 sg13g2_decap_8 FILLER_51_325 ();
 sg13g2_decap_4 FILLER_51_332 ();
 sg13g2_fill_2 FILLER_51_340 ();
 sg13g2_fill_1 FILLER_51_342 ();
 sg13g2_decap_8 FILLER_51_354 ();
 sg13g2_decap_8 FILLER_51_361 ();
 sg13g2_decap_8 FILLER_51_368 ();
 sg13g2_decap_8 FILLER_51_375 ();
 sg13g2_decap_8 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_4 FILLER_51_403 ();
 sg13g2_fill_1 FILLER_51_407 ();
 sg13g2_decap_4 FILLER_51_413 ();
 sg13g2_decap_4 FILLER_51_422 ();
 sg13g2_fill_1 FILLER_51_426 ();
 sg13g2_fill_2 FILLER_51_431 ();
 sg13g2_decap_4 FILLER_51_444 ();
 sg13g2_fill_2 FILLER_51_455 ();
 sg13g2_decap_8 FILLER_51_467 ();
 sg13g2_decap_8 FILLER_51_474 ();
 sg13g2_fill_1 FILLER_51_481 ();
 sg13g2_decap_4 FILLER_51_488 ();
 sg13g2_fill_2 FILLER_51_492 ();
 sg13g2_decap_8 FILLER_51_498 ();
 sg13g2_fill_2 FILLER_51_505 ();
 sg13g2_fill_1 FILLER_51_507 ();
 sg13g2_decap_8 FILLER_51_513 ();
 sg13g2_decap_8 FILLER_51_520 ();
 sg13g2_decap_4 FILLER_51_527 ();
 sg13g2_fill_1 FILLER_51_531 ();
 sg13g2_decap_8 FILLER_51_542 ();
 sg13g2_decap_8 FILLER_51_549 ();
 sg13g2_decap_4 FILLER_51_556 ();
 sg13g2_fill_2 FILLER_51_584 ();
 sg13g2_decap_4 FILLER_51_591 ();
 sg13g2_decap_8 FILLER_51_605 ();
 sg13g2_decap_4 FILLER_51_616 ();
 sg13g2_fill_1 FILLER_51_620 ();
 sg13g2_fill_1 FILLER_51_630 ();
 sg13g2_decap_4 FILLER_51_639 ();
 sg13g2_decap_8 FILLER_51_653 ();
 sg13g2_decap_8 FILLER_51_660 ();
 sg13g2_decap_8 FILLER_51_667 ();
 sg13g2_fill_2 FILLER_51_681 ();
 sg13g2_decap_8 FILLER_51_688 ();
 sg13g2_decap_8 FILLER_51_695 ();
 sg13g2_decap_8 FILLER_51_716 ();
 sg13g2_decap_4 FILLER_51_723 ();
 sg13g2_fill_2 FILLER_51_727 ();
 sg13g2_decap_8 FILLER_51_738 ();
 sg13g2_decap_8 FILLER_51_745 ();
 sg13g2_decap_8 FILLER_51_752 ();
 sg13g2_decap_8 FILLER_51_759 ();
 sg13g2_decap_8 FILLER_51_766 ();
 sg13g2_decap_8 FILLER_51_773 ();
 sg13g2_decap_8 FILLER_51_780 ();
 sg13g2_decap_8 FILLER_51_787 ();
 sg13g2_decap_8 FILLER_51_794 ();
 sg13g2_decap_8 FILLER_51_801 ();
 sg13g2_decap_8 FILLER_51_808 ();
 sg13g2_decap_8 FILLER_51_815 ();
 sg13g2_decap_8 FILLER_51_822 ();
 sg13g2_decap_8 FILLER_51_829 ();
 sg13g2_decap_8 FILLER_51_836 ();
 sg13g2_decap_8 FILLER_51_843 ();
 sg13g2_decap_8 FILLER_51_850 ();
 sg13g2_decap_8 FILLER_51_857 ();
 sg13g2_decap_8 FILLER_51_864 ();
 sg13g2_decap_8 FILLER_51_871 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_4 FILLER_52_42 ();
 sg13g2_decap_4 FILLER_52_55 ();
 sg13g2_fill_1 FILLER_52_59 ();
 sg13g2_decap_8 FILLER_52_65 ();
 sg13g2_decap_8 FILLER_52_72 ();
 sg13g2_fill_1 FILLER_52_79 ();
 sg13g2_decap_8 FILLER_52_85 ();
 sg13g2_fill_2 FILLER_52_92 ();
 sg13g2_decap_4 FILLER_52_98 ();
 sg13g2_fill_1 FILLER_52_102 ();
 sg13g2_fill_2 FILLER_52_108 ();
 sg13g2_fill_1 FILLER_52_110 ();
 sg13g2_decap_8 FILLER_52_115 ();
 sg13g2_decap_8 FILLER_52_122 ();
 sg13g2_decap_8 FILLER_52_129 ();
 sg13g2_decap_8 FILLER_52_136 ();
 sg13g2_decap_8 FILLER_52_143 ();
 sg13g2_decap_8 FILLER_52_150 ();
 sg13g2_decap_8 FILLER_52_157 ();
 sg13g2_decap_8 FILLER_52_164 ();
 sg13g2_decap_4 FILLER_52_171 ();
 sg13g2_fill_1 FILLER_52_175 ();
 sg13g2_decap_8 FILLER_52_184 ();
 sg13g2_decap_8 FILLER_52_191 ();
 sg13g2_decap_8 FILLER_52_198 ();
 sg13g2_decap_8 FILLER_52_205 ();
 sg13g2_fill_1 FILLER_52_212 ();
 sg13g2_decap_8 FILLER_52_228 ();
 sg13g2_decap_4 FILLER_52_235 ();
 sg13g2_decap_4 FILLER_52_244 ();
 sg13g2_fill_1 FILLER_52_248 ();
 sg13g2_decap_8 FILLER_52_269 ();
 sg13g2_decap_8 FILLER_52_276 ();
 sg13g2_decap_8 FILLER_52_283 ();
 sg13g2_decap_8 FILLER_52_290 ();
 sg13g2_fill_2 FILLER_52_297 ();
 sg13g2_fill_2 FILLER_52_313 ();
 sg13g2_decap_4 FILLER_52_318 ();
 sg13g2_fill_1 FILLER_52_322 ();
 sg13g2_fill_2 FILLER_52_331 ();
 sg13g2_fill_1 FILLER_52_333 ();
 sg13g2_decap_8 FILLER_52_340 ();
 sg13g2_decap_4 FILLER_52_347 ();
 sg13g2_fill_1 FILLER_52_351 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_4 FILLER_52_371 ();
 sg13g2_fill_1 FILLER_52_375 ();
 sg13g2_fill_2 FILLER_52_380 ();
 sg13g2_fill_1 FILLER_52_382 ();
 sg13g2_decap_8 FILLER_52_386 ();
 sg13g2_decap_8 FILLER_52_393 ();
 sg13g2_decap_4 FILLER_52_400 ();
 sg13g2_fill_2 FILLER_52_415 ();
 sg13g2_fill_2 FILLER_52_422 ();
 sg13g2_decap_8 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_52_436 ();
 sg13g2_decap_8 FILLER_52_443 ();
 sg13g2_decap_8 FILLER_52_450 ();
 sg13g2_decap_8 FILLER_52_457 ();
 sg13g2_decap_4 FILLER_52_464 ();
 sg13g2_fill_1 FILLER_52_468 ();
 sg13g2_decap_8 FILLER_52_478 ();
 sg13g2_decap_8 FILLER_52_485 ();
 sg13g2_fill_2 FILLER_52_492 ();
 sg13g2_fill_1 FILLER_52_494 ();
 sg13g2_fill_1 FILLER_52_510 ();
 sg13g2_decap_8 FILLER_52_516 ();
 sg13g2_decap_4 FILLER_52_523 ();
 sg13g2_decap_8 FILLER_52_537 ();
 sg13g2_decap_8 FILLER_52_544 ();
 sg13g2_decap_4 FILLER_52_554 ();
 sg13g2_fill_1 FILLER_52_558 ();
 sg13g2_decap_8 FILLER_52_569 ();
 sg13g2_decap_8 FILLER_52_576 ();
 sg13g2_decap_4 FILLER_52_583 ();
 sg13g2_decap_8 FILLER_52_591 ();
 sg13g2_decap_8 FILLER_52_598 ();
 sg13g2_decap_4 FILLER_52_614 ();
 sg13g2_fill_2 FILLER_52_618 ();
 sg13g2_decap_8 FILLER_52_626 ();
 sg13g2_decap_8 FILLER_52_633 ();
 sg13g2_decap_8 FILLER_52_644 ();
 sg13g2_decap_8 FILLER_52_651 ();
 sg13g2_decap_4 FILLER_52_658 ();
 sg13g2_fill_1 FILLER_52_662 ();
 sg13g2_fill_2 FILLER_52_667 ();
 sg13g2_fill_2 FILLER_52_680 ();
 sg13g2_fill_1 FILLER_52_682 ();
 sg13g2_decap_8 FILLER_52_697 ();
 sg13g2_fill_2 FILLER_52_704 ();
 sg13g2_fill_1 FILLER_52_706 ();
 sg13g2_decap_4 FILLER_52_711 ();
 sg13g2_decap_8 FILLER_52_724 ();
 sg13g2_decap_8 FILLER_52_731 ();
 sg13g2_decap_8 FILLER_52_738 ();
 sg13g2_decap_8 FILLER_52_754 ();
 sg13g2_fill_2 FILLER_52_765 ();
 sg13g2_decap_8 FILLER_52_770 ();
 sg13g2_decap_8 FILLER_52_777 ();
 sg13g2_decap_8 FILLER_52_784 ();
 sg13g2_decap_8 FILLER_52_791 ();
 sg13g2_decap_8 FILLER_52_798 ();
 sg13g2_decap_8 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_decap_8 FILLER_52_840 ();
 sg13g2_decap_8 FILLER_52_847 ();
 sg13g2_decap_8 FILLER_52_854 ();
 sg13g2_decap_8 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_52_868 ();
 sg13g2_fill_2 FILLER_52_875 ();
 sg13g2_fill_1 FILLER_52_877 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_fill_2 FILLER_53_56 ();
 sg13g2_fill_1 FILLER_53_58 ();
 sg13g2_fill_2 FILLER_53_63 ();
 sg13g2_fill_1 FILLER_53_65 ();
 sg13g2_decap_4 FILLER_53_71 ();
 sg13g2_decap_8 FILLER_53_80 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_decap_8 FILLER_53_100 ();
 sg13g2_fill_1 FILLER_53_107 ();
 sg13g2_decap_8 FILLER_53_117 ();
 sg13g2_decap_8 FILLER_53_124 ();
 sg13g2_decap_8 FILLER_53_131 ();
 sg13g2_decap_8 FILLER_53_138 ();
 sg13g2_decap_8 FILLER_53_145 ();
 sg13g2_fill_2 FILLER_53_162 ();
 sg13g2_decap_8 FILLER_53_174 ();
 sg13g2_decap_8 FILLER_53_181 ();
 sg13g2_decap_8 FILLER_53_188 ();
 sg13g2_decap_4 FILLER_53_195 ();
 sg13g2_decap_8 FILLER_53_204 ();
 sg13g2_decap_8 FILLER_53_211 ();
 sg13g2_decap_4 FILLER_53_218 ();
 sg13g2_fill_2 FILLER_53_222 ();
 sg13g2_fill_2 FILLER_53_229 ();
 sg13g2_fill_2 FILLER_53_236 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_decap_4 FILLER_53_255 ();
 sg13g2_decap_8 FILLER_53_264 ();
 sg13g2_decap_8 FILLER_53_271 ();
 sg13g2_decap_8 FILLER_53_281 ();
 sg13g2_fill_1 FILLER_53_288 ();
 sg13g2_decap_4 FILLER_53_297 ();
 sg13g2_decap_8 FILLER_53_306 ();
 sg13g2_decap_8 FILLER_53_313 ();
 sg13g2_fill_2 FILLER_53_320 ();
 sg13g2_fill_1 FILLER_53_322 ();
 sg13g2_decap_8 FILLER_53_337 ();
 sg13g2_decap_8 FILLER_53_344 ();
 sg13g2_decap_8 FILLER_53_351 ();
 sg13g2_decap_8 FILLER_53_358 ();
 sg13g2_decap_4 FILLER_53_365 ();
 sg13g2_fill_1 FILLER_53_369 ();
 sg13g2_fill_1 FILLER_53_375 ();
 sg13g2_decap_4 FILLER_53_381 ();
 sg13g2_decap_8 FILLER_53_389 ();
 sg13g2_decap_8 FILLER_53_396 ();
 sg13g2_decap_8 FILLER_53_403 ();
 sg13g2_fill_2 FILLER_53_410 ();
 sg13g2_fill_1 FILLER_53_412 ();
 sg13g2_decap_8 FILLER_53_418 ();
 sg13g2_decap_8 FILLER_53_425 ();
 sg13g2_decap_8 FILLER_53_432 ();
 sg13g2_fill_2 FILLER_53_439 ();
 sg13g2_decap_8 FILLER_53_446 ();
 sg13g2_decap_8 FILLER_53_453 ();
 sg13g2_decap_4 FILLER_53_460 ();
 sg13g2_fill_2 FILLER_53_469 ();
 sg13g2_fill_1 FILLER_53_471 ();
 sg13g2_decap_8 FILLER_53_481 ();
 sg13g2_decap_8 FILLER_53_488 ();
 sg13g2_decap_8 FILLER_53_495 ();
 sg13g2_fill_2 FILLER_53_502 ();
 sg13g2_decap_8 FILLER_53_513 ();
 sg13g2_decap_8 FILLER_53_520 ();
 sg13g2_decap_8 FILLER_53_527 ();
 sg13g2_decap_8 FILLER_53_542 ();
 sg13g2_decap_8 FILLER_53_549 ();
 sg13g2_decap_8 FILLER_53_556 ();
 sg13g2_fill_2 FILLER_53_563 ();
 sg13g2_fill_2 FILLER_53_570 ();
 sg13g2_decap_8 FILLER_53_577 ();
 sg13g2_decap_8 FILLER_53_584 ();
 sg13g2_decap_8 FILLER_53_591 ();
 sg13g2_decap_4 FILLER_53_603 ();
 sg13g2_fill_1 FILLER_53_607 ();
 sg13g2_decap_8 FILLER_53_612 ();
 sg13g2_decap_8 FILLER_53_619 ();
 sg13g2_decap_8 FILLER_53_626 ();
 sg13g2_fill_2 FILLER_53_633 ();
 sg13g2_decap_8 FILLER_53_639 ();
 sg13g2_decap_4 FILLER_53_646 ();
 sg13g2_fill_1 FILLER_53_655 ();
 sg13g2_decap_4 FILLER_53_660 ();
 sg13g2_fill_2 FILLER_53_669 ();
 sg13g2_decap_4 FILLER_53_681 ();
 sg13g2_fill_1 FILLER_53_685 ();
 sg13g2_decap_8 FILLER_53_696 ();
 sg13g2_decap_4 FILLER_53_703 ();
 sg13g2_fill_1 FILLER_53_707 ();
 sg13g2_fill_2 FILLER_53_718 ();
 sg13g2_fill_1 FILLER_53_720 ();
 sg13g2_decap_8 FILLER_53_726 ();
 sg13g2_decap_8 FILLER_53_733 ();
 sg13g2_decap_8 FILLER_53_740 ();
 sg13g2_decap_8 FILLER_53_747 ();
 sg13g2_decap_8 FILLER_53_754 ();
 sg13g2_decap_8 FILLER_53_761 ();
 sg13g2_decap_8 FILLER_53_768 ();
 sg13g2_decap_8 FILLER_53_775 ();
 sg13g2_decap_8 FILLER_53_782 ();
 sg13g2_decap_8 FILLER_53_789 ();
 sg13g2_decap_8 FILLER_53_796 ();
 sg13g2_decap_8 FILLER_53_803 ();
 sg13g2_decap_8 FILLER_53_810 ();
 sg13g2_decap_8 FILLER_53_817 ();
 sg13g2_decap_8 FILLER_53_824 ();
 sg13g2_decap_8 FILLER_53_831 ();
 sg13g2_decap_8 FILLER_53_838 ();
 sg13g2_decap_8 FILLER_53_845 ();
 sg13g2_decap_8 FILLER_53_852 ();
 sg13g2_decap_8 FILLER_53_859 ();
 sg13g2_decap_8 FILLER_53_866 ();
 sg13g2_decap_4 FILLER_53_873 ();
 sg13g2_fill_1 FILLER_53_877 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_4 FILLER_54_70 ();
 sg13g2_fill_1 FILLER_54_74 ();
 sg13g2_decap_4 FILLER_54_88 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_fill_2 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_118 ();
 sg13g2_decap_4 FILLER_54_129 ();
 sg13g2_decap_4 FILLER_54_137 ();
 sg13g2_decap_4 FILLER_54_145 ();
 sg13g2_fill_2 FILLER_54_149 ();
 sg13g2_decap_4 FILLER_54_161 ();
 sg13g2_decap_4 FILLER_54_170 ();
 sg13g2_decap_8 FILLER_54_178 ();
 sg13g2_decap_8 FILLER_54_185 ();
 sg13g2_decap_4 FILLER_54_192 ();
 sg13g2_fill_1 FILLER_54_196 ();
 sg13g2_decap_8 FILLER_54_201 ();
 sg13g2_decap_8 FILLER_54_208 ();
 sg13g2_decap_4 FILLER_54_215 ();
 sg13g2_fill_1 FILLER_54_219 ();
 sg13g2_decap_8 FILLER_54_228 ();
 sg13g2_decap_4 FILLER_54_235 ();
 sg13g2_fill_1 FILLER_54_239 ();
 sg13g2_fill_2 FILLER_54_245 ();
 sg13g2_fill_1 FILLER_54_247 ();
 sg13g2_fill_2 FILLER_54_253 ();
 sg13g2_fill_1 FILLER_54_255 ();
 sg13g2_decap_8 FILLER_54_261 ();
 sg13g2_decap_8 FILLER_54_268 ();
 sg13g2_decap_8 FILLER_54_275 ();
 sg13g2_decap_8 FILLER_54_282 ();
 sg13g2_fill_1 FILLER_54_289 ();
 sg13g2_decap_8 FILLER_54_295 ();
 sg13g2_fill_1 FILLER_54_302 ();
 sg13g2_decap_4 FILLER_54_313 ();
 sg13g2_fill_2 FILLER_54_317 ();
 sg13g2_fill_2 FILLER_54_324 ();
 sg13g2_fill_1 FILLER_54_326 ();
 sg13g2_decap_8 FILLER_54_339 ();
 sg13g2_decap_8 FILLER_54_346 ();
 sg13g2_fill_1 FILLER_54_353 ();
 sg13g2_fill_2 FILLER_54_362 ();
 sg13g2_decap_8 FILLER_54_369 ();
 sg13g2_decap_8 FILLER_54_376 ();
 sg13g2_fill_1 FILLER_54_383 ();
 sg13g2_fill_1 FILLER_54_389 ();
 sg13g2_decap_8 FILLER_54_394 ();
 sg13g2_decap_8 FILLER_54_401 ();
 sg13g2_decap_4 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_54_417 ();
 sg13g2_decap_8 FILLER_54_424 ();
 sg13g2_fill_2 FILLER_54_431 ();
 sg13g2_fill_1 FILLER_54_433 ();
 sg13g2_fill_1 FILLER_54_449 ();
 sg13g2_decap_8 FILLER_54_453 ();
 sg13g2_decap_8 FILLER_54_460 ();
 sg13g2_fill_1 FILLER_54_467 ();
 sg13g2_decap_8 FILLER_54_473 ();
 sg13g2_fill_2 FILLER_54_480 ();
 sg13g2_decap_8 FILLER_54_487 ();
 sg13g2_decap_8 FILLER_54_494 ();
 sg13g2_decap_8 FILLER_54_501 ();
 sg13g2_decap_8 FILLER_54_513 ();
 sg13g2_decap_8 FILLER_54_520 ();
 sg13g2_fill_2 FILLER_54_527 ();
 sg13g2_decap_8 FILLER_54_534 ();
 sg13g2_decap_8 FILLER_54_541 ();
 sg13g2_decap_8 FILLER_54_548 ();
 sg13g2_decap_8 FILLER_54_555 ();
 sg13g2_fill_2 FILLER_54_562 ();
 sg13g2_fill_1 FILLER_54_564 ();
 sg13g2_fill_2 FILLER_54_570 ();
 sg13g2_fill_1 FILLER_54_572 ();
 sg13g2_decap_4 FILLER_54_577 ();
 sg13g2_fill_2 FILLER_54_593 ();
 sg13g2_decap_8 FILLER_54_600 ();
 sg13g2_fill_2 FILLER_54_607 ();
 sg13g2_fill_1 FILLER_54_609 ();
 sg13g2_decap_8 FILLER_54_613 ();
 sg13g2_decap_8 FILLER_54_620 ();
 sg13g2_decap_4 FILLER_54_627 ();
 sg13g2_decap_8 FILLER_54_640 ();
 sg13g2_decap_4 FILLER_54_647 ();
 sg13g2_fill_1 FILLER_54_651 ();
 sg13g2_decap_8 FILLER_54_666 ();
 sg13g2_decap_4 FILLER_54_673 ();
 sg13g2_fill_2 FILLER_54_677 ();
 sg13g2_decap_8 FILLER_54_684 ();
 sg13g2_fill_2 FILLER_54_691 ();
 sg13g2_decap_8 FILLER_54_697 ();
 sg13g2_decap_8 FILLER_54_704 ();
 sg13g2_decap_8 FILLER_54_711 ();
 sg13g2_decap_8 FILLER_54_718 ();
 sg13g2_decap_4 FILLER_54_729 ();
 sg13g2_decap_8 FILLER_54_737 ();
 sg13g2_decap_8 FILLER_54_744 ();
 sg13g2_decap_8 FILLER_54_751 ();
 sg13g2_decap_8 FILLER_54_758 ();
 sg13g2_decap_8 FILLER_54_765 ();
 sg13g2_decap_8 FILLER_54_772 ();
 sg13g2_decap_8 FILLER_54_779 ();
 sg13g2_decap_8 FILLER_54_786 ();
 sg13g2_decap_8 FILLER_54_793 ();
 sg13g2_decap_8 FILLER_54_800 ();
 sg13g2_decap_8 FILLER_54_807 ();
 sg13g2_decap_8 FILLER_54_814 ();
 sg13g2_decap_8 FILLER_54_821 ();
 sg13g2_decap_8 FILLER_54_828 ();
 sg13g2_decap_8 FILLER_54_835 ();
 sg13g2_decap_8 FILLER_54_842 ();
 sg13g2_decap_8 FILLER_54_849 ();
 sg13g2_decap_8 FILLER_54_856 ();
 sg13g2_decap_8 FILLER_54_863 ();
 sg13g2_decap_8 FILLER_54_870 ();
 sg13g2_fill_1 FILLER_54_877 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_4 FILLER_55_42 ();
 sg13g2_fill_1 FILLER_55_46 ();
 sg13g2_decap_8 FILLER_55_51 ();
 sg13g2_decap_8 FILLER_55_58 ();
 sg13g2_decap_4 FILLER_55_65 ();
 sg13g2_fill_1 FILLER_55_69 ();
 sg13g2_decap_8 FILLER_55_79 ();
 sg13g2_decap_8 FILLER_55_86 ();
 sg13g2_decap_8 FILLER_55_93 ();
 sg13g2_decap_8 FILLER_55_100 ();
 sg13g2_decap_8 FILLER_55_107 ();
 sg13g2_fill_2 FILLER_55_114 ();
 sg13g2_fill_1 FILLER_55_116 ();
 sg13g2_decap_8 FILLER_55_122 ();
 sg13g2_decap_4 FILLER_55_129 ();
 sg13g2_fill_1 FILLER_55_133 ();
 sg13g2_fill_2 FILLER_55_138 ();
 sg13g2_fill_1 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_146 ();
 sg13g2_decap_8 FILLER_55_153 ();
 sg13g2_fill_2 FILLER_55_165 ();
 sg13g2_decap_8 FILLER_55_172 ();
 sg13g2_decap_8 FILLER_55_179 ();
 sg13g2_fill_2 FILLER_55_186 ();
 sg13g2_fill_1 FILLER_55_188 ();
 sg13g2_decap_8 FILLER_55_198 ();
 sg13g2_decap_8 FILLER_55_209 ();
 sg13g2_decap_8 FILLER_55_216 ();
 sg13g2_decap_8 FILLER_55_223 ();
 sg13g2_decap_8 FILLER_55_235 ();
 sg13g2_fill_2 FILLER_55_242 ();
 sg13g2_decap_4 FILLER_55_254 ();
 sg13g2_decap_8 FILLER_55_262 ();
 sg13g2_decap_4 FILLER_55_269 ();
 sg13g2_fill_1 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_279 ();
 sg13g2_decap_8 FILLER_55_286 ();
 sg13g2_decap_4 FILLER_55_293 ();
 sg13g2_fill_1 FILLER_55_297 ();
 sg13g2_decap_8 FILLER_55_302 ();
 sg13g2_decap_8 FILLER_55_309 ();
 sg13g2_fill_2 FILLER_55_316 ();
 sg13g2_fill_1 FILLER_55_318 ();
 sg13g2_fill_2 FILLER_55_324 ();
 sg13g2_decap_8 FILLER_55_329 ();
 sg13g2_decap_8 FILLER_55_336 ();
 sg13g2_fill_2 FILLER_55_343 ();
 sg13g2_decap_8 FILLER_55_354 ();
 sg13g2_decap_8 FILLER_55_361 ();
 sg13g2_decap_4 FILLER_55_368 ();
 sg13g2_fill_2 FILLER_55_372 ();
 sg13g2_decap_4 FILLER_55_379 ();
 sg13g2_fill_1 FILLER_55_383 ();
 sg13g2_decap_8 FILLER_55_390 ();
 sg13g2_decap_8 FILLER_55_397 ();
 sg13g2_decap_4 FILLER_55_404 ();
 sg13g2_fill_2 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_55_419 ();
 sg13g2_decap_8 FILLER_55_426 ();
 sg13g2_decap_8 FILLER_55_433 ();
 sg13g2_decap_4 FILLER_55_440 ();
 sg13g2_fill_2 FILLER_55_444 ();
 sg13g2_decap_8 FILLER_55_462 ();
 sg13g2_decap_4 FILLER_55_469 ();
 sg13g2_fill_1 FILLER_55_473 ();
 sg13g2_fill_1 FILLER_55_479 ();
 sg13g2_decap_8 FILLER_55_489 ();
 sg13g2_decap_8 FILLER_55_496 ();
 sg13g2_fill_1 FILLER_55_503 ();
 sg13g2_decap_8 FILLER_55_518 ();
 sg13g2_decap_8 FILLER_55_525 ();
 sg13g2_fill_1 FILLER_55_532 ();
 sg13g2_fill_1 FILLER_55_537 ();
 sg13g2_decap_8 FILLER_55_543 ();
 sg13g2_decap_8 FILLER_55_550 ();
 sg13g2_decap_4 FILLER_55_557 ();
 sg13g2_fill_1 FILLER_55_561 ();
 sg13g2_fill_2 FILLER_55_567 ();
 sg13g2_fill_2 FILLER_55_574 ();
 sg13g2_decap_8 FILLER_55_585 ();
 sg13g2_decap_8 FILLER_55_592 ();
 sg13g2_decap_4 FILLER_55_604 ();
 sg13g2_fill_1 FILLER_55_608 ();
 sg13g2_decap_8 FILLER_55_613 ();
 sg13g2_decap_4 FILLER_55_647 ();
 sg13g2_fill_1 FILLER_55_651 ();
 sg13g2_decap_8 FILLER_55_655 ();
 sg13g2_decap_8 FILLER_55_662 ();
 sg13g2_decap_8 FILLER_55_669 ();
 sg13g2_fill_2 FILLER_55_676 ();
 sg13g2_fill_2 FILLER_55_682 ();
 sg13g2_fill_1 FILLER_55_684 ();
 sg13g2_fill_2 FILLER_55_689 ();
 sg13g2_fill_1 FILLER_55_699 ();
 sg13g2_fill_2 FILLER_55_705 ();
 sg13g2_fill_1 FILLER_55_707 ();
 sg13g2_fill_2 FILLER_55_713 ();
 sg13g2_fill_2 FILLER_55_729 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_decap_8 FILLER_55_744 ();
 sg13g2_decap_8 FILLER_55_751 ();
 sg13g2_decap_8 FILLER_55_758 ();
 sg13g2_decap_8 FILLER_55_765 ();
 sg13g2_decap_8 FILLER_55_772 ();
 sg13g2_decap_8 FILLER_55_779 ();
 sg13g2_decap_8 FILLER_55_786 ();
 sg13g2_decap_8 FILLER_55_793 ();
 sg13g2_decap_8 FILLER_55_800 ();
 sg13g2_decap_8 FILLER_55_807 ();
 sg13g2_decap_8 FILLER_55_814 ();
 sg13g2_decap_8 FILLER_55_821 ();
 sg13g2_decap_8 FILLER_55_828 ();
 sg13g2_decap_8 FILLER_55_835 ();
 sg13g2_decap_8 FILLER_55_842 ();
 sg13g2_decap_8 FILLER_55_849 ();
 sg13g2_decap_8 FILLER_55_856 ();
 sg13g2_decap_8 FILLER_55_863 ();
 sg13g2_decap_8 FILLER_55_870 ();
 sg13g2_fill_1 FILLER_55_877 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_63 ();
 sg13g2_fill_2 FILLER_56_76 ();
 sg13g2_fill_1 FILLER_56_78 ();
 sg13g2_decap_4 FILLER_56_83 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_4 FILLER_56_105 ();
 sg13g2_fill_2 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_128 ();
 sg13g2_decap_8 FILLER_56_134 ();
 sg13g2_decap_4 FILLER_56_141 ();
 sg13g2_fill_2 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_155 ();
 sg13g2_decap_8 FILLER_56_169 ();
 sg13g2_decap_4 FILLER_56_176 ();
 sg13g2_fill_1 FILLER_56_180 ();
 sg13g2_fill_2 FILLER_56_196 ();
 sg13g2_fill_1 FILLER_56_198 ();
 sg13g2_decap_8 FILLER_56_209 ();
 sg13g2_decap_8 FILLER_56_216 ();
 sg13g2_decap_8 FILLER_56_223 ();
 sg13g2_fill_1 FILLER_56_230 ();
 sg13g2_decap_4 FILLER_56_235 ();
 sg13g2_decap_4 FILLER_56_243 ();
 sg13g2_fill_1 FILLER_56_247 ();
 sg13g2_decap_8 FILLER_56_253 ();
 sg13g2_fill_2 FILLER_56_271 ();
 sg13g2_decap_8 FILLER_56_278 ();
 sg13g2_decap_8 FILLER_56_285 ();
 sg13g2_decap_8 FILLER_56_292 ();
 sg13g2_decap_8 FILLER_56_299 ();
 sg13g2_decap_8 FILLER_56_306 ();
 sg13g2_fill_2 FILLER_56_313 ();
 sg13g2_fill_1 FILLER_56_315 ();
 sg13g2_fill_2 FILLER_56_320 ();
 sg13g2_decap_8 FILLER_56_326 ();
 sg13g2_decap_8 FILLER_56_333 ();
 sg13g2_decap_8 FILLER_56_340 ();
 sg13g2_fill_2 FILLER_56_347 ();
 sg13g2_decap_8 FILLER_56_353 ();
 sg13g2_decap_4 FILLER_56_365 ();
 sg13g2_decap_8 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_385 ();
 sg13g2_decap_8 FILLER_56_392 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_decap_8 FILLER_56_416 ();
 sg13g2_decap_8 FILLER_56_423 ();
 sg13g2_decap_4 FILLER_56_430 ();
 sg13g2_fill_1 FILLER_56_434 ();
 sg13g2_decap_8 FILLER_56_439 ();
 sg13g2_decap_8 FILLER_56_446 ();
 sg13g2_fill_2 FILLER_56_453 ();
 sg13g2_fill_1 FILLER_56_455 ();
 sg13g2_decap_8 FILLER_56_461 ();
 sg13g2_decap_4 FILLER_56_468 ();
 sg13g2_fill_1 FILLER_56_472 ();
 sg13g2_fill_2 FILLER_56_477 ();
 sg13g2_fill_1 FILLER_56_479 ();
 sg13g2_decap_4 FILLER_56_485 ();
 sg13g2_decap_8 FILLER_56_493 ();
 sg13g2_fill_1 FILLER_56_500 ();
 sg13g2_fill_1 FILLER_56_506 ();
 sg13g2_fill_1 FILLER_56_511 ();
 sg13g2_fill_2 FILLER_56_529 ();
 sg13g2_fill_1 FILLER_56_531 ();
 sg13g2_decap_8 FILLER_56_542 ();
 sg13g2_decap_8 FILLER_56_549 ();
 sg13g2_decap_8 FILLER_56_556 ();
 sg13g2_fill_2 FILLER_56_563 ();
 sg13g2_decap_8 FILLER_56_574 ();
 sg13g2_decap_4 FILLER_56_581 ();
 sg13g2_decap_8 FILLER_56_592 ();
 sg13g2_decap_8 FILLER_56_599 ();
 sg13g2_fill_2 FILLER_56_606 ();
 sg13g2_decap_4 FILLER_56_614 ();
 sg13g2_fill_1 FILLER_56_618 ();
 sg13g2_decap_8 FILLER_56_624 ();
 sg13g2_decap_8 FILLER_56_631 ();
 sg13g2_fill_2 FILLER_56_638 ();
 sg13g2_decap_8 FILLER_56_645 ();
 sg13g2_fill_1 FILLER_56_652 ();
 sg13g2_fill_2 FILLER_56_664 ();
 sg13g2_fill_2 FILLER_56_670 ();
 sg13g2_fill_1 FILLER_56_672 ();
 sg13g2_fill_1 FILLER_56_677 ();
 sg13g2_decap_4 FILLER_56_682 ();
 sg13g2_fill_1 FILLER_56_695 ();
 sg13g2_decap_4 FILLER_56_700 ();
 sg13g2_fill_1 FILLER_56_707 ();
 sg13g2_decap_8 FILLER_56_712 ();
 sg13g2_decap_8 FILLER_56_719 ();
 sg13g2_decap_8 FILLER_56_726 ();
 sg13g2_decap_8 FILLER_56_733 ();
 sg13g2_decap_8 FILLER_56_740 ();
 sg13g2_decap_8 FILLER_56_747 ();
 sg13g2_decap_8 FILLER_56_754 ();
 sg13g2_decap_8 FILLER_56_761 ();
 sg13g2_decap_8 FILLER_56_768 ();
 sg13g2_decap_8 FILLER_56_775 ();
 sg13g2_decap_8 FILLER_56_782 ();
 sg13g2_decap_8 FILLER_56_789 ();
 sg13g2_decap_8 FILLER_56_796 ();
 sg13g2_decap_8 FILLER_56_803 ();
 sg13g2_decap_8 FILLER_56_810 ();
 sg13g2_decap_8 FILLER_56_817 ();
 sg13g2_decap_8 FILLER_56_824 ();
 sg13g2_decap_8 FILLER_56_831 ();
 sg13g2_decap_8 FILLER_56_838 ();
 sg13g2_decap_8 FILLER_56_845 ();
 sg13g2_decap_8 FILLER_56_852 ();
 sg13g2_decap_8 FILLER_56_859 ();
 sg13g2_decap_8 FILLER_56_866 ();
 sg13g2_decap_4 FILLER_56_873 ();
 sg13g2_fill_1 FILLER_56_877 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_4 FILLER_57_63 ();
 sg13g2_fill_2 FILLER_57_67 ();
 sg13g2_decap_8 FILLER_57_73 ();
 sg13g2_decap_4 FILLER_57_80 ();
 sg13g2_fill_1 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_93 ();
 sg13g2_decap_8 FILLER_57_100 ();
 sg13g2_decap_8 FILLER_57_107 ();
 sg13g2_fill_2 FILLER_57_114 ();
 sg13g2_decap_8 FILLER_57_124 ();
 sg13g2_decap_8 FILLER_57_131 ();
 sg13g2_decap_4 FILLER_57_138 ();
 sg13g2_fill_2 FILLER_57_142 ();
 sg13g2_decap_4 FILLER_57_150 ();
 sg13g2_decap_4 FILLER_57_162 ();
 sg13g2_fill_1 FILLER_57_166 ();
 sg13g2_fill_1 FILLER_57_170 ();
 sg13g2_decap_4 FILLER_57_185 ();
 sg13g2_decap_8 FILLER_57_198 ();
 sg13g2_fill_2 FILLER_57_205 ();
 sg13g2_fill_1 FILLER_57_207 ();
 sg13g2_decap_8 FILLER_57_213 ();
 sg13g2_decap_8 FILLER_57_220 ();
 sg13g2_decap_4 FILLER_57_227 ();
 sg13g2_fill_1 FILLER_57_231 ();
 sg13g2_decap_8 FILLER_57_241 ();
 sg13g2_decap_8 FILLER_57_248 ();
 sg13g2_decap_4 FILLER_57_255 ();
 sg13g2_fill_2 FILLER_57_259 ();
 sg13g2_decap_8 FILLER_57_266 ();
 sg13g2_decap_8 FILLER_57_273 ();
 sg13g2_decap_8 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_287 ();
 sg13g2_decap_4 FILLER_57_298 ();
 sg13g2_decap_4 FILLER_57_315 ();
 sg13g2_fill_2 FILLER_57_319 ();
 sg13g2_fill_2 FILLER_57_326 ();
 sg13g2_fill_1 FILLER_57_328 ();
 sg13g2_fill_1 FILLER_57_348 ();
 sg13g2_decap_8 FILLER_57_353 ();
 sg13g2_decap_8 FILLER_57_360 ();
 sg13g2_decap_8 FILLER_57_367 ();
 sg13g2_decap_8 FILLER_57_374 ();
 sg13g2_fill_1 FILLER_57_381 ();
 sg13g2_decap_8 FILLER_57_390 ();
 sg13g2_decap_4 FILLER_57_397 ();
 sg13g2_fill_1 FILLER_57_401 ();
 sg13g2_decap_4 FILLER_57_406 ();
 sg13g2_fill_2 FILLER_57_414 ();
 sg13g2_decap_4 FILLER_57_424 ();
 sg13g2_decap_8 FILLER_57_433 ();
 sg13g2_decap_8 FILLER_57_440 ();
 sg13g2_fill_2 FILLER_57_447 ();
 sg13g2_decap_8 FILLER_57_453 ();
 sg13g2_decap_8 FILLER_57_460 ();
 sg13g2_decap_8 FILLER_57_467 ();
 sg13g2_fill_2 FILLER_57_474 ();
 sg13g2_fill_1 FILLER_57_476 ();
 sg13g2_decap_8 FILLER_57_482 ();
 sg13g2_fill_2 FILLER_57_489 ();
 sg13g2_decap_8 FILLER_57_495 ();
 sg13g2_decap_8 FILLER_57_502 ();
 sg13g2_fill_1 FILLER_57_509 ();
 sg13g2_fill_2 FILLER_57_515 ();
 sg13g2_decap_4 FILLER_57_521 ();
 sg13g2_fill_2 FILLER_57_530 ();
 sg13g2_fill_1 FILLER_57_532 ();
 sg13g2_decap_4 FILLER_57_537 ();
 sg13g2_fill_1 FILLER_57_541 ();
 sg13g2_decap_8 FILLER_57_547 ();
 sg13g2_decap_4 FILLER_57_554 ();
 sg13g2_fill_1 FILLER_57_558 ();
 sg13g2_decap_8 FILLER_57_569 ();
 sg13g2_decap_8 FILLER_57_585 ();
 sg13g2_decap_8 FILLER_57_592 ();
 sg13g2_decap_8 FILLER_57_599 ();
 sg13g2_decap_8 FILLER_57_606 ();
 sg13g2_decap_8 FILLER_57_613 ();
 sg13g2_fill_1 FILLER_57_620 ();
 sg13g2_decap_8 FILLER_57_649 ();
 sg13g2_decap_8 FILLER_57_656 ();
 sg13g2_decap_8 FILLER_57_663 ();
 sg13g2_decap_8 FILLER_57_674 ();
 sg13g2_decap_8 FILLER_57_681 ();
 sg13g2_decap_8 FILLER_57_692 ();
 sg13g2_decap_8 FILLER_57_699 ();
 sg13g2_decap_8 FILLER_57_706 ();
 sg13g2_decap_8 FILLER_57_713 ();
 sg13g2_decap_8 FILLER_57_720 ();
 sg13g2_decap_8 FILLER_57_727 ();
 sg13g2_decap_8 FILLER_57_734 ();
 sg13g2_decap_8 FILLER_57_741 ();
 sg13g2_decap_8 FILLER_57_748 ();
 sg13g2_decap_8 FILLER_57_755 ();
 sg13g2_decap_8 FILLER_57_762 ();
 sg13g2_decap_8 FILLER_57_769 ();
 sg13g2_decap_8 FILLER_57_776 ();
 sg13g2_decap_8 FILLER_57_783 ();
 sg13g2_decap_8 FILLER_57_790 ();
 sg13g2_decap_8 FILLER_57_797 ();
 sg13g2_decap_8 FILLER_57_804 ();
 sg13g2_decap_8 FILLER_57_811 ();
 sg13g2_decap_8 FILLER_57_818 ();
 sg13g2_decap_8 FILLER_57_825 ();
 sg13g2_decap_8 FILLER_57_832 ();
 sg13g2_decap_8 FILLER_57_839 ();
 sg13g2_decap_8 FILLER_57_846 ();
 sg13g2_decap_8 FILLER_57_853 ();
 sg13g2_decap_8 FILLER_57_860 ();
 sg13g2_decap_8 FILLER_57_867 ();
 sg13g2_decap_4 FILLER_57_874 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_4 FILLER_58_49 ();
 sg13g2_fill_2 FILLER_58_53 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_4 FILLER_58_105 ();
 sg13g2_fill_2 FILLER_58_109 ();
 sg13g2_decap_8 FILLER_58_116 ();
 sg13g2_decap_8 FILLER_58_123 ();
 sg13g2_decap_8 FILLER_58_130 ();
 sg13g2_decap_8 FILLER_58_137 ();
 sg13g2_decap_8 FILLER_58_144 ();
 sg13g2_decap_8 FILLER_58_151 ();
 sg13g2_decap_8 FILLER_58_158 ();
 sg13g2_fill_1 FILLER_58_165 ();
 sg13g2_decap_8 FILLER_58_170 ();
 sg13g2_decap_8 FILLER_58_177 ();
 sg13g2_decap_8 FILLER_58_184 ();
 sg13g2_decap_8 FILLER_58_191 ();
 sg13g2_decap_4 FILLER_58_198 ();
 sg13g2_fill_2 FILLER_58_206 ();
 sg13g2_decap_8 FILLER_58_220 ();
 sg13g2_fill_1 FILLER_58_227 ();
 sg13g2_decap_8 FILLER_58_232 ();
 sg13g2_decap_8 FILLER_58_239 ();
 sg13g2_decap_8 FILLER_58_246 ();
 sg13g2_decap_8 FILLER_58_253 ();
 sg13g2_decap_8 FILLER_58_260 ();
 sg13g2_decap_8 FILLER_58_267 ();
 sg13g2_decap_8 FILLER_58_274 ();
 sg13g2_decap_8 FILLER_58_281 ();
 sg13g2_fill_2 FILLER_58_288 ();
 sg13g2_fill_1 FILLER_58_290 ();
 sg13g2_decap_4 FILLER_58_299 ();
 sg13g2_decap_8 FILLER_58_311 ();
 sg13g2_decap_8 FILLER_58_318 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_fill_2 FILLER_58_336 ();
 sg13g2_fill_1 FILLER_58_338 ();
 sg13g2_fill_1 FILLER_58_342 ();
 sg13g2_fill_1 FILLER_58_347 ();
 sg13g2_decap_8 FILLER_58_353 ();
 sg13g2_decap_8 FILLER_58_360 ();
 sg13g2_decap_8 FILLER_58_367 ();
 sg13g2_fill_2 FILLER_58_374 ();
 sg13g2_fill_1 FILLER_58_376 ();
 sg13g2_fill_2 FILLER_58_382 ();
 sg13g2_fill_1 FILLER_58_384 ();
 sg13g2_decap_8 FILLER_58_390 ();
 sg13g2_fill_2 FILLER_58_397 ();
 sg13g2_decap_8 FILLER_58_408 ();
 sg13g2_decap_4 FILLER_58_415 ();
 sg13g2_fill_1 FILLER_58_419 ();
 sg13g2_fill_1 FILLER_58_433 ();
 sg13g2_decap_4 FILLER_58_439 ();
 sg13g2_fill_1 FILLER_58_443 ();
 sg13g2_fill_1 FILLER_58_448 ();
 sg13g2_decap_8 FILLER_58_457 ();
 sg13g2_decap_8 FILLER_58_464 ();
 sg13g2_decap_8 FILLER_58_471 ();
 sg13g2_decap_8 FILLER_58_478 ();
 sg13g2_decap_8 FILLER_58_485 ();
 sg13g2_decap_8 FILLER_58_492 ();
 sg13g2_fill_2 FILLER_58_499 ();
 sg13g2_fill_1 FILLER_58_501 ();
 sg13g2_fill_2 FILLER_58_506 ();
 sg13g2_fill_2 FILLER_58_512 ();
 sg13g2_fill_2 FILLER_58_520 ();
 sg13g2_decap_8 FILLER_58_526 ();
 sg13g2_fill_2 FILLER_58_533 ();
 sg13g2_decap_8 FILLER_58_538 ();
 sg13g2_decap_8 FILLER_58_545 ();
 sg13g2_decap_8 FILLER_58_552 ();
 sg13g2_decap_8 FILLER_58_570 ();
 sg13g2_decap_8 FILLER_58_577 ();
 sg13g2_decap_8 FILLER_58_584 ();
 sg13g2_decap_4 FILLER_58_591 ();
 sg13g2_fill_1 FILLER_58_595 ();
 sg13g2_fill_1 FILLER_58_600 ();
 sg13g2_decap_8 FILLER_58_606 ();
 sg13g2_decap_4 FILLER_58_613 ();
 sg13g2_fill_1 FILLER_58_617 ();
 sg13g2_decap_4 FILLER_58_630 ();
 sg13g2_decap_8 FILLER_58_639 ();
 sg13g2_decap_8 FILLER_58_646 ();
 sg13g2_decap_8 FILLER_58_653 ();
 sg13g2_decap_8 FILLER_58_660 ();
 sg13g2_decap_4 FILLER_58_667 ();
 sg13g2_fill_1 FILLER_58_671 ();
 sg13g2_fill_1 FILLER_58_682 ();
 sg13g2_decap_8 FILLER_58_695 ();
 sg13g2_decap_8 FILLER_58_702 ();
 sg13g2_fill_2 FILLER_58_709 ();
 sg13g2_fill_1 FILLER_58_711 ();
 sg13g2_decap_8 FILLER_58_730 ();
 sg13g2_decap_8 FILLER_58_737 ();
 sg13g2_decap_8 FILLER_58_757 ();
 sg13g2_decap_8 FILLER_58_764 ();
 sg13g2_decap_8 FILLER_58_771 ();
 sg13g2_decap_8 FILLER_58_778 ();
 sg13g2_decap_8 FILLER_58_785 ();
 sg13g2_decap_8 FILLER_58_792 ();
 sg13g2_decap_8 FILLER_58_799 ();
 sg13g2_decap_8 FILLER_58_806 ();
 sg13g2_decap_8 FILLER_58_813 ();
 sg13g2_decap_8 FILLER_58_820 ();
 sg13g2_decap_8 FILLER_58_827 ();
 sg13g2_decap_8 FILLER_58_834 ();
 sg13g2_decap_8 FILLER_58_841 ();
 sg13g2_decap_8 FILLER_58_848 ();
 sg13g2_decap_8 FILLER_58_855 ();
 sg13g2_decap_8 FILLER_58_862 ();
 sg13g2_decap_8 FILLER_58_869 ();
 sg13g2_fill_2 FILLER_58_876 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_4 FILLER_59_42 ();
 sg13g2_fill_1 FILLER_59_46 ();
 sg13g2_decap_8 FILLER_59_73 ();
 sg13g2_decap_8 FILLER_59_80 ();
 sg13g2_decap_8 FILLER_59_87 ();
 sg13g2_decap_8 FILLER_59_94 ();
 sg13g2_decap_8 FILLER_59_101 ();
 sg13g2_decap_4 FILLER_59_108 ();
 sg13g2_decap_8 FILLER_59_116 ();
 sg13g2_fill_1 FILLER_59_123 ();
 sg13g2_decap_8 FILLER_59_129 ();
 sg13g2_fill_2 FILLER_59_136 ();
 sg13g2_fill_1 FILLER_59_138 ();
 sg13g2_decap_8 FILLER_59_143 ();
 sg13g2_decap_8 FILLER_59_150 ();
 sg13g2_decap_4 FILLER_59_157 ();
 sg13g2_decap_8 FILLER_59_165 ();
 sg13g2_fill_2 FILLER_59_172 ();
 sg13g2_fill_1 FILLER_59_174 ();
 sg13g2_decap_8 FILLER_59_180 ();
 sg13g2_fill_2 FILLER_59_187 ();
 sg13g2_fill_1 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_194 ();
 sg13g2_decap_8 FILLER_59_201 ();
 sg13g2_fill_1 FILLER_59_208 ();
 sg13g2_decap_8 FILLER_59_213 ();
 sg13g2_decap_8 FILLER_59_220 ();
 sg13g2_decap_8 FILLER_59_227 ();
 sg13g2_decap_8 FILLER_59_234 ();
 sg13g2_decap_8 FILLER_59_241 ();
 sg13g2_decap_8 FILLER_59_248 ();
 sg13g2_decap_8 FILLER_59_255 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_decap_8 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_decap_8 FILLER_59_287 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_4 FILLER_59_301 ();
 sg13g2_fill_1 FILLER_59_309 ();
 sg13g2_decap_8 FILLER_59_314 ();
 sg13g2_decap_8 FILLER_59_321 ();
 sg13g2_decap_8 FILLER_59_328 ();
 sg13g2_decap_8 FILLER_59_335 ();
 sg13g2_decap_4 FILLER_59_342 ();
 sg13g2_fill_2 FILLER_59_346 ();
 sg13g2_decap_8 FILLER_59_353 ();
 sg13g2_decap_8 FILLER_59_360 ();
 sg13g2_decap_8 FILLER_59_367 ();
 sg13g2_fill_2 FILLER_59_374 ();
 sg13g2_decap_8 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_decap_4 FILLER_59_420 ();
 sg13g2_fill_1 FILLER_59_424 ();
 sg13g2_decap_8 FILLER_59_429 ();
 sg13g2_decap_8 FILLER_59_436 ();
 sg13g2_fill_2 FILLER_59_448 ();
 sg13g2_decap_8 FILLER_59_455 ();
 sg13g2_decap_8 FILLER_59_462 ();
 sg13g2_decap_4 FILLER_59_469 ();
 sg13g2_fill_2 FILLER_59_473 ();
 sg13g2_decap_8 FILLER_59_479 ();
 sg13g2_decap_8 FILLER_59_486 ();
 sg13g2_decap_8 FILLER_59_497 ();
 sg13g2_fill_1 FILLER_59_504 ();
 sg13g2_decap_8 FILLER_59_514 ();
 sg13g2_decap_8 FILLER_59_521 ();
 sg13g2_decap_8 FILLER_59_528 ();
 sg13g2_fill_2 FILLER_59_535 ();
 sg13g2_decap_8 FILLER_59_541 ();
 sg13g2_fill_2 FILLER_59_548 ();
 sg13g2_decap_8 FILLER_59_561 ();
 sg13g2_decap_8 FILLER_59_568 ();
 sg13g2_decap_4 FILLER_59_575 ();
 sg13g2_fill_2 FILLER_59_579 ();
 sg13g2_fill_2 FILLER_59_586 ();
 sg13g2_decap_8 FILLER_59_593 ();
 sg13g2_decap_8 FILLER_59_600 ();
 sg13g2_decap_8 FILLER_59_607 ();
 sg13g2_decap_8 FILLER_59_614 ();
 sg13g2_decap_8 FILLER_59_621 ();
 sg13g2_decap_8 FILLER_59_628 ();
 sg13g2_decap_8 FILLER_59_635 ();
 sg13g2_decap_8 FILLER_59_642 ();
 sg13g2_decap_8 FILLER_59_649 ();
 sg13g2_decap_8 FILLER_59_656 ();
 sg13g2_decap_8 FILLER_59_663 ();
 sg13g2_decap_8 FILLER_59_670 ();
 sg13g2_decap_8 FILLER_59_677 ();
 sg13g2_fill_2 FILLER_59_684 ();
 sg13g2_fill_1 FILLER_59_686 ();
 sg13g2_decap_8 FILLER_59_692 ();
 sg13g2_decap_4 FILLER_59_699 ();
 sg13g2_fill_2 FILLER_59_703 ();
 sg13g2_fill_2 FILLER_59_710 ();
 sg13g2_decap_8 FILLER_59_747 ();
 sg13g2_decap_8 FILLER_59_754 ();
 sg13g2_decap_8 FILLER_59_761 ();
 sg13g2_decap_8 FILLER_59_768 ();
 sg13g2_decap_8 FILLER_59_775 ();
 sg13g2_decap_8 FILLER_59_782 ();
 sg13g2_decap_8 FILLER_59_789 ();
 sg13g2_decap_8 FILLER_59_796 ();
 sg13g2_decap_8 FILLER_59_803 ();
 sg13g2_decap_8 FILLER_59_810 ();
 sg13g2_decap_8 FILLER_59_817 ();
 sg13g2_decap_8 FILLER_59_824 ();
 sg13g2_decap_8 FILLER_59_831 ();
 sg13g2_decap_8 FILLER_59_838 ();
 sg13g2_decap_8 FILLER_59_845 ();
 sg13g2_decap_8 FILLER_59_852 ();
 sg13g2_decap_8 FILLER_59_859 ();
 sg13g2_decap_8 FILLER_59_866 ();
 sg13g2_decap_4 FILLER_59_873 ();
 sg13g2_fill_1 FILLER_59_877 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_fill_2 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_fill_2 FILLER_60_98 ();
 sg13g2_fill_1 FILLER_60_100 ();
 sg13g2_fill_1 FILLER_60_131 ();
 sg13g2_decap_8 FILLER_60_158 ();
 sg13g2_decap_8 FILLER_60_165 ();
 sg13g2_decap_8 FILLER_60_172 ();
 sg13g2_decap_8 FILLER_60_179 ();
 sg13g2_decap_8 FILLER_60_186 ();
 sg13g2_decap_8 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_200 ();
 sg13g2_fill_2 FILLER_60_207 ();
 sg13g2_fill_1 FILLER_60_209 ();
 sg13g2_decap_8 FILLER_60_214 ();
 sg13g2_decap_8 FILLER_60_221 ();
 sg13g2_decap_8 FILLER_60_228 ();
 sg13g2_decap_8 FILLER_60_235 ();
 sg13g2_decap_4 FILLER_60_242 ();
 sg13g2_decap_4 FILLER_60_250 ();
 sg13g2_fill_1 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_275 ();
 sg13g2_decap_8 FILLER_60_282 ();
 sg13g2_decap_8 FILLER_60_289 ();
 sg13g2_decap_8 FILLER_60_296 ();
 sg13g2_decap_8 FILLER_60_303 ();
 sg13g2_decap_8 FILLER_60_314 ();
 sg13g2_decap_8 FILLER_60_321 ();
 sg13g2_decap_8 FILLER_60_328 ();
 sg13g2_decap_8 FILLER_60_335 ();
 sg13g2_decap_4 FILLER_60_342 ();
 sg13g2_fill_2 FILLER_60_346 ();
 sg13g2_decap_8 FILLER_60_354 ();
 sg13g2_decap_8 FILLER_60_361 ();
 sg13g2_decap_8 FILLER_60_368 ();
 sg13g2_decap_8 FILLER_60_375 ();
 sg13g2_decap_4 FILLER_60_382 ();
 sg13g2_fill_2 FILLER_60_386 ();
 sg13g2_decap_8 FILLER_60_391 ();
 sg13g2_decap_8 FILLER_60_398 ();
 sg13g2_decap_8 FILLER_60_405 ();
 sg13g2_decap_8 FILLER_60_412 ();
 sg13g2_decap_8 FILLER_60_419 ();
 sg13g2_decap_8 FILLER_60_426 ();
 sg13g2_decap_8 FILLER_60_433 ();
 sg13g2_decap_8 FILLER_60_440 ();
 sg13g2_decap_8 FILLER_60_447 ();
 sg13g2_decap_8 FILLER_60_454 ();
 sg13g2_decap_8 FILLER_60_461 ();
 sg13g2_decap_8 FILLER_60_468 ();
 sg13g2_decap_8 FILLER_60_475 ();
 sg13g2_fill_2 FILLER_60_482 ();
 sg13g2_fill_1 FILLER_60_484 ();
 sg13g2_fill_1 FILLER_60_489 ();
 sg13g2_fill_1 FILLER_60_494 ();
 sg13g2_fill_1 FILLER_60_499 ();
 sg13g2_decap_8 FILLER_60_513 ();
 sg13g2_decap_8 FILLER_60_520 ();
 sg13g2_decap_8 FILLER_60_527 ();
 sg13g2_decap_4 FILLER_60_534 ();
 sg13g2_decap_8 FILLER_60_546 ();
 sg13g2_decap_8 FILLER_60_553 ();
 sg13g2_decap_8 FILLER_60_560 ();
 sg13g2_decap_8 FILLER_60_567 ();
 sg13g2_decap_8 FILLER_60_574 ();
 sg13g2_decap_8 FILLER_60_581 ();
 sg13g2_decap_8 FILLER_60_588 ();
 sg13g2_decap_4 FILLER_60_595 ();
 sg13g2_decap_8 FILLER_60_603 ();
 sg13g2_decap_8 FILLER_60_610 ();
 sg13g2_decap_8 FILLER_60_617 ();
 sg13g2_fill_1 FILLER_60_624 ();
 sg13g2_decap_8 FILLER_60_628 ();
 sg13g2_decap_8 FILLER_60_635 ();
 sg13g2_decap_8 FILLER_60_642 ();
 sg13g2_decap_8 FILLER_60_649 ();
 sg13g2_decap_8 FILLER_60_656 ();
 sg13g2_decap_8 FILLER_60_663 ();
 sg13g2_decap_8 FILLER_60_670 ();
 sg13g2_decap_8 FILLER_60_677 ();
 sg13g2_fill_1 FILLER_60_684 ();
 sg13g2_fill_2 FILLER_60_689 ();
 sg13g2_decap_8 FILLER_60_694 ();
 sg13g2_decap_8 FILLER_60_701 ();
 sg13g2_decap_8 FILLER_60_708 ();
 sg13g2_decap_8 FILLER_60_715 ();
 sg13g2_decap_8 FILLER_60_722 ();
 sg13g2_decap_4 FILLER_60_729 ();
 sg13g2_decap_8 FILLER_60_739 ();
 sg13g2_fill_2 FILLER_60_746 ();
 sg13g2_fill_1 FILLER_60_748 ();
 sg13g2_decap_8 FILLER_60_754 ();
 sg13g2_decap_8 FILLER_60_761 ();
 sg13g2_decap_8 FILLER_60_768 ();
 sg13g2_decap_8 FILLER_60_775 ();
 sg13g2_decap_8 FILLER_60_782 ();
 sg13g2_decap_8 FILLER_60_789 ();
 sg13g2_decap_8 FILLER_60_796 ();
 sg13g2_decap_8 FILLER_60_803 ();
 sg13g2_decap_8 FILLER_60_810 ();
 sg13g2_decap_8 FILLER_60_817 ();
 sg13g2_decap_8 FILLER_60_824 ();
 sg13g2_decap_8 FILLER_60_831 ();
 sg13g2_decap_8 FILLER_60_838 ();
 sg13g2_decap_8 FILLER_60_845 ();
 sg13g2_decap_8 FILLER_60_852 ();
 sg13g2_decap_8 FILLER_60_859 ();
 sg13g2_decap_8 FILLER_60_866 ();
 sg13g2_decap_4 FILLER_60_873 ();
 sg13g2_fill_1 FILLER_60_877 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_fill_1 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_54 ();
 sg13g2_decap_8 FILLER_61_61 ();
 sg13g2_decap_8 FILLER_61_68 ();
 sg13g2_decap_8 FILLER_61_75 ();
 sg13g2_decap_4 FILLER_61_82 ();
 sg13g2_decap_8 FILLER_61_90 ();
 sg13g2_decap_8 FILLER_61_97 ();
 sg13g2_decap_8 FILLER_61_104 ();
 sg13g2_decap_8 FILLER_61_111 ();
 sg13g2_fill_2 FILLER_61_118 ();
 sg13g2_fill_1 FILLER_61_146 ();
 sg13g2_decap_8 FILLER_61_151 ();
 sg13g2_decap_8 FILLER_61_158 ();
 sg13g2_decap_8 FILLER_61_165 ();
 sg13g2_decap_8 FILLER_61_172 ();
 sg13g2_decap_8 FILLER_61_179 ();
 sg13g2_fill_2 FILLER_61_186 ();
 sg13g2_decap_8 FILLER_61_192 ();
 sg13g2_decap_8 FILLER_61_199 ();
 sg13g2_decap_8 FILLER_61_206 ();
 sg13g2_decap_8 FILLER_61_213 ();
 sg13g2_decap_4 FILLER_61_220 ();
 sg13g2_decap_8 FILLER_61_228 ();
 sg13g2_decap_8 FILLER_61_235 ();
 sg13g2_decap_8 FILLER_61_242 ();
 sg13g2_decap_8 FILLER_61_249 ();
 sg13g2_decap_4 FILLER_61_256 ();
 sg13g2_fill_1 FILLER_61_260 ();
 sg13g2_decap_4 FILLER_61_269 ();
 sg13g2_fill_2 FILLER_61_273 ();
 sg13g2_decap_8 FILLER_61_285 ();
 sg13g2_decap_8 FILLER_61_292 ();
 sg13g2_decap_8 FILLER_61_299 ();
 sg13g2_decap_8 FILLER_61_314 ();
 sg13g2_decap_8 FILLER_61_321 ();
 sg13g2_decap_8 FILLER_61_328 ();
 sg13g2_fill_2 FILLER_61_335 ();
 sg13g2_decap_8 FILLER_61_355 ();
 sg13g2_decap_8 FILLER_61_362 ();
 sg13g2_decap_8 FILLER_61_369 ();
 sg13g2_decap_8 FILLER_61_376 ();
 sg13g2_decap_8 FILLER_61_383 ();
 sg13g2_decap_8 FILLER_61_390 ();
 sg13g2_decap_8 FILLER_61_397 ();
 sg13g2_decap_4 FILLER_61_404 ();
 sg13g2_decap_4 FILLER_61_416 ();
 sg13g2_decap_8 FILLER_61_432 ();
 sg13g2_fill_1 FILLER_61_439 ();
 sg13g2_decap_8 FILLER_61_448 ();
 sg13g2_decap_8 FILLER_61_455 ();
 sg13g2_decap_8 FILLER_61_462 ();
 sg13g2_decap_8 FILLER_61_469 ();
 sg13g2_decap_8 FILLER_61_476 ();
 sg13g2_decap_8 FILLER_61_483 ();
 sg13g2_decap_8 FILLER_61_490 ();
 sg13g2_fill_2 FILLER_61_501 ();
 sg13g2_fill_1 FILLER_61_503 ();
 sg13g2_decap_8 FILLER_61_508 ();
 sg13g2_decap_8 FILLER_61_515 ();
 sg13g2_decap_8 FILLER_61_522 ();
 sg13g2_decap_4 FILLER_61_529 ();
 sg13g2_fill_2 FILLER_61_533 ();
 sg13g2_decap_8 FILLER_61_569 ();
 sg13g2_decap_8 FILLER_61_576 ();
 sg13g2_decap_8 FILLER_61_583 ();
 sg13g2_decap_4 FILLER_61_616 ();
 sg13g2_fill_2 FILLER_61_620 ();
 sg13g2_decap_8 FILLER_61_651 ();
 sg13g2_fill_1 FILLER_61_658 ();
 sg13g2_decap_8 FILLER_61_677 ();
 sg13g2_decap_4 FILLER_61_684 ();
 sg13g2_decap_4 FILLER_61_717 ();
 sg13g2_fill_2 FILLER_61_721 ();
 sg13g2_decap_8 FILLER_61_759 ();
 sg13g2_decap_8 FILLER_61_766 ();
 sg13g2_decap_8 FILLER_61_773 ();
 sg13g2_decap_8 FILLER_61_780 ();
 sg13g2_decap_8 FILLER_61_787 ();
 sg13g2_decap_8 FILLER_61_794 ();
 sg13g2_decap_8 FILLER_61_801 ();
 sg13g2_decap_8 FILLER_61_808 ();
 sg13g2_decap_8 FILLER_61_815 ();
 sg13g2_decap_8 FILLER_61_822 ();
 sg13g2_decap_8 FILLER_61_829 ();
 sg13g2_decap_8 FILLER_61_836 ();
 sg13g2_decap_8 FILLER_61_843 ();
 sg13g2_decap_8 FILLER_61_850 ();
 sg13g2_decap_8 FILLER_61_857 ();
 sg13g2_decap_8 FILLER_61_864 ();
 sg13g2_decap_8 FILLER_61_871 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_fill_2 FILLER_62_42 ();
 sg13g2_fill_1 FILLER_62_44 ();
 sg13g2_decap_8 FILLER_62_71 ();
 sg13g2_decap_8 FILLER_62_78 ();
 sg13g2_decap_8 FILLER_62_85 ();
 sg13g2_decap_8 FILLER_62_92 ();
 sg13g2_decap_8 FILLER_62_99 ();
 sg13g2_decap_8 FILLER_62_106 ();
 sg13g2_decap_8 FILLER_62_113 ();
 sg13g2_decap_8 FILLER_62_120 ();
 sg13g2_decap_8 FILLER_62_127 ();
 sg13g2_decap_8 FILLER_62_134 ();
 sg13g2_decap_8 FILLER_62_171 ();
 sg13g2_decap_8 FILLER_62_178 ();
 sg13g2_decap_8 FILLER_62_185 ();
 sg13g2_decap_8 FILLER_62_192 ();
 sg13g2_decap_4 FILLER_62_199 ();
 sg13g2_fill_1 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_230 ();
 sg13g2_decap_8 FILLER_62_237 ();
 sg13g2_decap_8 FILLER_62_244 ();
 sg13g2_decap_8 FILLER_62_251 ();
 sg13g2_decap_4 FILLER_62_258 ();
 sg13g2_fill_2 FILLER_62_278 ();
 sg13g2_decap_8 FILLER_62_285 ();
 sg13g2_decap_8 FILLER_62_292 ();
 sg13g2_fill_2 FILLER_62_299 ();
 sg13g2_decap_8 FILLER_62_332 ();
 sg13g2_decap_4 FILLER_62_339 ();
 sg13g2_fill_1 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_349 ();
 sg13g2_decap_4 FILLER_62_356 ();
 sg13g2_fill_2 FILLER_62_360 ();
 sg13g2_fill_1 FILLER_62_366 ();
 sg13g2_decap_8 FILLER_62_372 ();
 sg13g2_decap_8 FILLER_62_379 ();
 sg13g2_decap_8 FILLER_62_386 ();
 sg13g2_decap_8 FILLER_62_393 ();
 sg13g2_decap_4 FILLER_62_400 ();
 sg13g2_fill_2 FILLER_62_408 ();
 sg13g2_fill_2 FILLER_62_426 ();
 sg13g2_fill_1 FILLER_62_428 ();
 sg13g2_decap_8 FILLER_62_434 ();
 sg13g2_decap_8 FILLER_62_441 ();
 sg13g2_decap_8 FILLER_62_448 ();
 sg13g2_decap_8 FILLER_62_455 ();
 sg13g2_decap_8 FILLER_62_462 ();
 sg13g2_decap_8 FILLER_62_469 ();
 sg13g2_decap_8 FILLER_62_476 ();
 sg13g2_decap_8 FILLER_62_483 ();
 sg13g2_decap_8 FILLER_62_490 ();
 sg13g2_fill_2 FILLER_62_497 ();
 sg13g2_decap_8 FILLER_62_503 ();
 sg13g2_decap_8 FILLER_62_510 ();
 sg13g2_decap_8 FILLER_62_517 ();
 sg13g2_decap_8 FILLER_62_524 ();
 sg13g2_decap_8 FILLER_62_531 ();
 sg13g2_decap_8 FILLER_62_538 ();
 sg13g2_fill_1 FILLER_62_545 ();
 sg13g2_decap_8 FILLER_62_550 ();
 sg13g2_decap_8 FILLER_62_557 ();
 sg13g2_decap_8 FILLER_62_564 ();
 sg13g2_decap_8 FILLER_62_571 ();
 sg13g2_decap_8 FILLER_62_578 ();
 sg13g2_decap_8 FILLER_62_585 ();
 sg13g2_decap_8 FILLER_62_592 ();
 sg13g2_decap_8 FILLER_62_599 ();
 sg13g2_decap_8 FILLER_62_606 ();
 sg13g2_decap_8 FILLER_62_613 ();
 sg13g2_decap_8 FILLER_62_620 ();
 sg13g2_decap_4 FILLER_62_627 ();
 sg13g2_fill_1 FILLER_62_631 ();
 sg13g2_decap_4 FILLER_62_636 ();
 sg13g2_fill_1 FILLER_62_640 ();
 sg13g2_decap_8 FILLER_62_646 ();
 sg13g2_decap_8 FILLER_62_688 ();
 sg13g2_fill_1 FILLER_62_695 ();
 sg13g2_decap_8 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_707 ();
 sg13g2_decap_8 FILLER_62_714 ();
 sg13g2_decap_8 FILLER_62_721 ();
 sg13g2_decap_8 FILLER_62_728 ();
 sg13g2_decap_8 FILLER_62_735 ();
 sg13g2_decap_8 FILLER_62_746 ();
 sg13g2_decap_8 FILLER_62_753 ();
 sg13g2_decap_8 FILLER_62_760 ();
 sg13g2_decap_8 FILLER_62_767 ();
 sg13g2_decap_8 FILLER_62_774 ();
 sg13g2_decap_8 FILLER_62_781 ();
 sg13g2_decap_8 FILLER_62_788 ();
 sg13g2_decap_8 FILLER_62_795 ();
 sg13g2_decap_8 FILLER_62_802 ();
 sg13g2_decap_8 FILLER_62_809 ();
 sg13g2_decap_8 FILLER_62_816 ();
 sg13g2_decap_8 FILLER_62_823 ();
 sg13g2_decap_8 FILLER_62_830 ();
 sg13g2_decap_8 FILLER_62_837 ();
 sg13g2_decap_8 FILLER_62_844 ();
 sg13g2_decap_8 FILLER_62_851 ();
 sg13g2_decap_8 FILLER_62_858 ();
 sg13g2_decap_8 FILLER_62_865 ();
 sg13g2_decap_4 FILLER_62_872 ();
 sg13g2_fill_2 FILLER_62_876 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_fill_2 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_55 ();
 sg13g2_decap_8 FILLER_63_66 ();
 sg13g2_decap_8 FILLER_63_73 ();
 sg13g2_decap_8 FILLER_63_80 ();
 sg13g2_decap_8 FILLER_63_87 ();
 sg13g2_decap_8 FILLER_63_94 ();
 sg13g2_decap_8 FILLER_63_101 ();
 sg13g2_decap_8 FILLER_63_108 ();
 sg13g2_decap_8 FILLER_63_115 ();
 sg13g2_decap_8 FILLER_63_122 ();
 sg13g2_decap_8 FILLER_63_129 ();
 sg13g2_decap_8 FILLER_63_136 ();
 sg13g2_decap_8 FILLER_63_143 ();
 sg13g2_decap_8 FILLER_63_150 ();
 sg13g2_fill_2 FILLER_63_157 ();
 sg13g2_decap_8 FILLER_63_185 ();
 sg13g2_fill_2 FILLER_63_192 ();
 sg13g2_fill_1 FILLER_63_194 ();
 sg13g2_decap_8 FILLER_63_199 ();
 sg13g2_decap_4 FILLER_63_206 ();
 sg13g2_fill_2 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_216 ();
 sg13g2_decap_8 FILLER_63_223 ();
 sg13g2_decap_8 FILLER_63_230 ();
 sg13g2_decap_8 FILLER_63_237 ();
 sg13g2_decap_8 FILLER_63_244 ();
 sg13g2_decap_8 FILLER_63_251 ();
 sg13g2_decap_8 FILLER_63_258 ();
 sg13g2_decap_4 FILLER_63_265 ();
 sg13g2_fill_1 FILLER_63_269 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_decap_4 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_288 ();
 sg13g2_decap_8 FILLER_63_295 ();
 sg13g2_decap_8 FILLER_63_302 ();
 sg13g2_decap_4 FILLER_63_309 ();
 sg13g2_decap_8 FILLER_63_317 ();
 sg13g2_decap_8 FILLER_63_324 ();
 sg13g2_decap_8 FILLER_63_331 ();
 sg13g2_decap_8 FILLER_63_338 ();
 sg13g2_fill_2 FILLER_63_345 ();
 sg13g2_decap_4 FILLER_63_360 ();
 sg13g2_fill_1 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_4 FILLER_63_399 ();
 sg13g2_fill_2 FILLER_63_403 ();
 sg13g2_fill_1 FILLER_63_414 ();
 sg13g2_fill_2 FILLER_63_420 ();
 sg13g2_fill_1 FILLER_63_428 ();
 sg13g2_decap_8 FILLER_63_433 ();
 sg13g2_decap_8 FILLER_63_440 ();
 sg13g2_decap_8 FILLER_63_447 ();
 sg13g2_decap_8 FILLER_63_454 ();
 sg13g2_decap_8 FILLER_63_461 ();
 sg13g2_decap_8 FILLER_63_468 ();
 sg13g2_decap_8 FILLER_63_475 ();
 sg13g2_decap_8 FILLER_63_482 ();
 sg13g2_decap_8 FILLER_63_489 ();
 sg13g2_decap_8 FILLER_63_496 ();
 sg13g2_decap_8 FILLER_63_503 ();
 sg13g2_decap_8 FILLER_63_510 ();
 sg13g2_decap_8 FILLER_63_517 ();
 sg13g2_decap_8 FILLER_63_524 ();
 sg13g2_decap_8 FILLER_63_531 ();
 sg13g2_decap_8 FILLER_63_538 ();
 sg13g2_decap_8 FILLER_63_545 ();
 sg13g2_decap_8 FILLER_63_552 ();
 sg13g2_decap_8 FILLER_63_559 ();
 sg13g2_decap_8 FILLER_63_566 ();
 sg13g2_decap_8 FILLER_63_573 ();
 sg13g2_decap_8 FILLER_63_580 ();
 sg13g2_decap_4 FILLER_63_587 ();
 sg13g2_fill_1 FILLER_63_591 ();
 sg13g2_decap_8 FILLER_63_600 ();
 sg13g2_decap_8 FILLER_63_607 ();
 sg13g2_decap_8 FILLER_63_614 ();
 sg13g2_decap_8 FILLER_63_621 ();
 sg13g2_decap_8 FILLER_63_628 ();
 sg13g2_decap_8 FILLER_63_635 ();
 sg13g2_decap_8 FILLER_63_642 ();
 sg13g2_decap_8 FILLER_63_649 ();
 sg13g2_fill_2 FILLER_63_656 ();
 sg13g2_fill_1 FILLER_63_658 ();
 sg13g2_decap_4 FILLER_63_662 ();
 sg13g2_fill_2 FILLER_63_666 ();
 sg13g2_decap_8 FILLER_63_672 ();
 sg13g2_decap_8 FILLER_63_679 ();
 sg13g2_decap_8 FILLER_63_686 ();
 sg13g2_decap_8 FILLER_63_693 ();
 sg13g2_decap_8 FILLER_63_700 ();
 sg13g2_decap_8 FILLER_63_707 ();
 sg13g2_decap_8 FILLER_63_714 ();
 sg13g2_decap_8 FILLER_63_721 ();
 sg13g2_decap_8 FILLER_63_728 ();
 sg13g2_decap_8 FILLER_63_735 ();
 sg13g2_decap_8 FILLER_63_742 ();
 sg13g2_decap_8 FILLER_63_749 ();
 sg13g2_decap_8 FILLER_63_756 ();
 sg13g2_decap_8 FILLER_63_763 ();
 sg13g2_decap_8 FILLER_63_770 ();
 sg13g2_decap_8 FILLER_63_777 ();
 sg13g2_decap_8 FILLER_63_784 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_decap_8 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_decap_8 FILLER_63_812 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_decap_8 FILLER_63_840 ();
 sg13g2_decap_8 FILLER_63_847 ();
 sg13g2_decap_8 FILLER_63_854 ();
 sg13g2_decap_8 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_63_868 ();
 sg13g2_fill_2 FILLER_63_875 ();
 sg13g2_fill_1 FILLER_63_877 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_4 FILLER_64_49 ();
 sg13g2_fill_2 FILLER_64_53 ();
 sg13g2_decap_8 FILLER_64_81 ();
 sg13g2_decap_4 FILLER_64_88 ();
 sg13g2_fill_1 FILLER_64_92 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_fill_1 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_163 ();
 sg13g2_decap_8 FILLER_64_170 ();
 sg13g2_decap_8 FILLER_64_177 ();
 sg13g2_decap_4 FILLER_64_184 ();
 sg13g2_fill_1 FILLER_64_188 ();
 sg13g2_decap_8 FILLER_64_215 ();
 sg13g2_decap_8 FILLER_64_222 ();
 sg13g2_decap_8 FILLER_64_229 ();
 sg13g2_decap_8 FILLER_64_236 ();
 sg13g2_decap_8 FILLER_64_243 ();
 sg13g2_decap_8 FILLER_64_250 ();
 sg13g2_decap_8 FILLER_64_257 ();
 sg13g2_decap_8 FILLER_64_264 ();
 sg13g2_fill_1 FILLER_64_271 ();
 sg13g2_decap_8 FILLER_64_285 ();
 sg13g2_decap_8 FILLER_64_292 ();
 sg13g2_decap_8 FILLER_64_299 ();
 sg13g2_decap_8 FILLER_64_306 ();
 sg13g2_decap_4 FILLER_64_313 ();
 sg13g2_fill_1 FILLER_64_317 ();
 sg13g2_decap_8 FILLER_64_323 ();
 sg13g2_decap_8 FILLER_64_330 ();
 sg13g2_decap_8 FILLER_64_337 ();
 sg13g2_decap_4 FILLER_64_344 ();
 sg13g2_decap_8 FILLER_64_374 ();
 sg13g2_decap_8 FILLER_64_381 ();
 sg13g2_decap_8 FILLER_64_388 ();
 sg13g2_decap_8 FILLER_64_395 ();
 sg13g2_decap_8 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_64_414 ();
 sg13g2_decap_8 FILLER_64_421 ();
 sg13g2_decap_8 FILLER_64_428 ();
 sg13g2_decap_8 FILLER_64_435 ();
 sg13g2_decap_8 FILLER_64_442 ();
 sg13g2_decap_8 FILLER_64_449 ();
 sg13g2_decap_8 FILLER_64_456 ();
 sg13g2_decap_8 FILLER_64_463 ();
 sg13g2_decap_8 FILLER_64_470 ();
 sg13g2_decap_8 FILLER_64_477 ();
 sg13g2_decap_8 FILLER_64_484 ();
 sg13g2_decap_8 FILLER_64_491 ();
 sg13g2_decap_8 FILLER_64_498 ();
 sg13g2_decap_8 FILLER_64_505 ();
 sg13g2_decap_8 FILLER_64_512 ();
 sg13g2_fill_1 FILLER_64_519 ();
 sg13g2_decap_8 FILLER_64_537 ();
 sg13g2_decap_8 FILLER_64_544 ();
 sg13g2_decap_8 FILLER_64_551 ();
 sg13g2_decap_8 FILLER_64_558 ();
 sg13g2_decap_8 FILLER_64_565 ();
 sg13g2_decap_8 FILLER_64_572 ();
 sg13g2_decap_4 FILLER_64_579 ();
 sg13g2_decap_8 FILLER_64_591 ();
 sg13g2_decap_8 FILLER_64_598 ();
 sg13g2_decap_8 FILLER_64_605 ();
 sg13g2_decap_8 FILLER_64_612 ();
 sg13g2_decap_8 FILLER_64_619 ();
 sg13g2_decap_8 FILLER_64_626 ();
 sg13g2_decap_8 FILLER_64_633 ();
 sg13g2_decap_8 FILLER_64_640 ();
 sg13g2_decap_8 FILLER_64_647 ();
 sg13g2_decap_8 FILLER_64_654 ();
 sg13g2_decap_8 FILLER_64_661 ();
 sg13g2_decap_8 FILLER_64_668 ();
 sg13g2_decap_8 FILLER_64_675 ();
 sg13g2_decap_8 FILLER_64_682 ();
 sg13g2_decap_8 FILLER_64_689 ();
 sg13g2_decap_8 FILLER_64_696 ();
 sg13g2_decap_8 FILLER_64_703 ();
 sg13g2_decap_8 FILLER_64_710 ();
 sg13g2_decap_8 FILLER_64_717 ();
 sg13g2_decap_8 FILLER_64_724 ();
 sg13g2_decap_8 FILLER_64_731 ();
 sg13g2_decap_8 FILLER_64_738 ();
 sg13g2_decap_8 FILLER_64_745 ();
 sg13g2_decap_8 FILLER_64_752 ();
 sg13g2_decap_8 FILLER_64_759 ();
 sg13g2_decap_8 FILLER_64_766 ();
 sg13g2_decap_8 FILLER_64_773 ();
 sg13g2_decap_8 FILLER_64_780 ();
 sg13g2_decap_8 FILLER_64_787 ();
 sg13g2_decap_8 FILLER_64_794 ();
 sg13g2_decap_8 FILLER_64_801 ();
 sg13g2_decap_8 FILLER_64_808 ();
 sg13g2_decap_8 FILLER_64_815 ();
 sg13g2_decap_8 FILLER_64_822 ();
 sg13g2_decap_8 FILLER_64_829 ();
 sg13g2_decap_8 FILLER_64_836 ();
 sg13g2_decap_8 FILLER_64_843 ();
 sg13g2_decap_8 FILLER_64_850 ();
 sg13g2_decap_8 FILLER_64_857 ();
 sg13g2_decap_8 FILLER_64_864 ();
 sg13g2_decap_8 FILLER_64_871 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_fill_1 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_103 ();
 sg13g2_decap_8 FILLER_65_110 ();
 sg13g2_decap_8 FILLER_65_117 ();
 sg13g2_decap_8 FILLER_65_124 ();
 sg13g2_decap_8 FILLER_65_131 ();
 sg13g2_decap_8 FILLER_65_138 ();
 sg13g2_decap_8 FILLER_65_145 ();
 sg13g2_decap_4 FILLER_65_157 ();
 sg13g2_fill_1 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_188 ();
 sg13g2_decap_4 FILLER_65_195 ();
 sg13g2_fill_1 FILLER_65_199 ();
 sg13g2_decap_8 FILLER_65_226 ();
 sg13g2_decap_8 FILLER_65_233 ();
 sg13g2_decap_8 FILLER_65_240 ();
 sg13g2_decap_8 FILLER_65_247 ();
 sg13g2_decap_8 FILLER_65_254 ();
 sg13g2_decap_8 FILLER_65_261 ();
 sg13g2_decap_8 FILLER_65_268 ();
 sg13g2_decap_8 FILLER_65_275 ();
 sg13g2_decap_8 FILLER_65_282 ();
 sg13g2_decap_8 FILLER_65_289 ();
 sg13g2_decap_4 FILLER_65_296 ();
 sg13g2_fill_1 FILLER_65_300 ();
 sg13g2_decap_8 FILLER_65_306 ();
 sg13g2_decap_8 FILLER_65_313 ();
 sg13g2_decap_8 FILLER_65_320 ();
 sg13g2_decap_8 FILLER_65_327 ();
 sg13g2_decap_8 FILLER_65_334 ();
 sg13g2_decap_8 FILLER_65_341 ();
 sg13g2_decap_8 FILLER_65_348 ();
 sg13g2_fill_2 FILLER_65_355 ();
 sg13g2_decap_8 FILLER_65_361 ();
 sg13g2_decap_8 FILLER_65_368 ();
 sg13g2_decap_8 FILLER_65_375 ();
 sg13g2_decap_8 FILLER_65_382 ();
 sg13g2_decap_8 FILLER_65_389 ();
 sg13g2_decap_8 FILLER_65_404 ();
 sg13g2_decap_8 FILLER_65_411 ();
 sg13g2_decap_8 FILLER_65_418 ();
 sg13g2_decap_8 FILLER_65_425 ();
 sg13g2_decap_8 FILLER_65_432 ();
 sg13g2_decap_8 FILLER_65_439 ();
 sg13g2_decap_8 FILLER_65_446 ();
 sg13g2_fill_2 FILLER_65_453 ();
 sg13g2_fill_1 FILLER_65_455 ();
 sg13g2_decap_4 FILLER_65_482 ();
 sg13g2_decap_8 FILLER_65_490 ();
 sg13g2_decap_4 FILLER_65_497 ();
 sg13g2_fill_1 FILLER_65_501 ();
 sg13g2_decap_8 FILLER_65_558 ();
 sg13g2_fill_2 FILLER_65_565 ();
 sg13g2_fill_1 FILLER_65_567 ();
 sg13g2_fill_2 FILLER_65_594 ();
 sg13g2_fill_1 FILLER_65_596 ();
 sg13g2_decap_8 FILLER_65_623 ();
 sg13g2_decap_8 FILLER_65_630 ();
 sg13g2_decap_8 FILLER_65_637 ();
 sg13g2_decap_8 FILLER_65_644 ();
 sg13g2_decap_8 FILLER_65_651 ();
 sg13g2_decap_8 FILLER_65_658 ();
 sg13g2_decap_8 FILLER_65_665 ();
 sg13g2_decap_8 FILLER_65_672 ();
 sg13g2_decap_8 FILLER_65_679 ();
 sg13g2_decap_8 FILLER_65_686 ();
 sg13g2_decap_8 FILLER_65_693 ();
 sg13g2_decap_8 FILLER_65_700 ();
 sg13g2_decap_8 FILLER_65_707 ();
 sg13g2_decap_8 FILLER_65_714 ();
 sg13g2_decap_8 FILLER_65_721 ();
 sg13g2_decap_8 FILLER_65_728 ();
 sg13g2_decap_8 FILLER_65_735 ();
 sg13g2_decap_8 FILLER_65_742 ();
 sg13g2_decap_8 FILLER_65_749 ();
 sg13g2_decap_8 FILLER_65_756 ();
 sg13g2_decap_8 FILLER_65_763 ();
 sg13g2_decap_8 FILLER_65_770 ();
 sg13g2_decap_8 FILLER_65_777 ();
 sg13g2_decap_8 FILLER_65_784 ();
 sg13g2_decap_8 FILLER_65_791 ();
 sg13g2_decap_8 FILLER_65_798 ();
 sg13g2_decap_8 FILLER_65_805 ();
 sg13g2_decap_8 FILLER_65_812 ();
 sg13g2_decap_8 FILLER_65_819 ();
 sg13g2_decap_8 FILLER_65_826 ();
 sg13g2_decap_8 FILLER_65_833 ();
 sg13g2_decap_8 FILLER_65_840 ();
 sg13g2_decap_8 FILLER_65_847 ();
 sg13g2_decap_8 FILLER_65_854 ();
 sg13g2_decap_8 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_65_868 ();
 sg13g2_fill_2 FILLER_65_875 ();
 sg13g2_fill_1 FILLER_65_877 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_4 FILLER_66_35 ();
 sg13g2_fill_1 FILLER_66_43 ();
 sg13g2_decap_8 FILLER_66_61 ();
 sg13g2_decap_8 FILLER_66_68 ();
 sg13g2_fill_1 FILLER_66_75 ();
 sg13g2_decap_4 FILLER_66_81 ();
 sg13g2_fill_1 FILLER_66_85 ();
 sg13g2_decap_8 FILLER_66_96 ();
 sg13g2_decap_8 FILLER_66_103 ();
 sg13g2_decap_4 FILLER_66_110 ();
 sg13g2_decap_8 FILLER_66_117 ();
 sg13g2_decap_8 FILLER_66_124 ();
 sg13g2_decap_8 FILLER_66_131 ();
 sg13g2_decap_8 FILLER_66_138 ();
 sg13g2_decap_8 FILLER_66_145 ();
 sg13g2_decap_8 FILLER_66_152 ();
 sg13g2_decap_8 FILLER_66_159 ();
 sg13g2_fill_2 FILLER_66_166 ();
 sg13g2_fill_1 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_173 ();
 sg13g2_decap_8 FILLER_66_180 ();
 sg13g2_decap_8 FILLER_66_187 ();
 sg13g2_decap_8 FILLER_66_194 ();
 sg13g2_decap_8 FILLER_66_201 ();
 sg13g2_decap_8 FILLER_66_212 ();
 sg13g2_decap_8 FILLER_66_219 ();
 sg13g2_fill_2 FILLER_66_226 ();
 sg13g2_decap_8 FILLER_66_254 ();
 sg13g2_decap_8 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_4 FILLER_66_280 ();
 sg13g2_fill_2 FILLER_66_284 ();
 sg13g2_decap_8 FILLER_66_291 ();
 sg13g2_decap_8 FILLER_66_298 ();
 sg13g2_fill_1 FILLER_66_305 ();
 sg13g2_decap_8 FILLER_66_311 ();
 sg13g2_decap_8 FILLER_66_318 ();
 sg13g2_decap_8 FILLER_66_325 ();
 sg13g2_decap_8 FILLER_66_332 ();
 sg13g2_decap_8 FILLER_66_339 ();
 sg13g2_decap_8 FILLER_66_346 ();
 sg13g2_decap_8 FILLER_66_353 ();
 sg13g2_decap_8 FILLER_66_360 ();
 sg13g2_decap_8 FILLER_66_367 ();
 sg13g2_decap_8 FILLER_66_374 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_4 FILLER_66_392 ();
 sg13g2_fill_2 FILLER_66_396 ();
 sg13g2_decap_8 FILLER_66_424 ();
 sg13g2_decap_8 FILLER_66_431 ();
 sg13g2_decap_8 FILLER_66_438 ();
 sg13g2_decap_8 FILLER_66_445 ();
 sg13g2_decap_4 FILLER_66_452 ();
 sg13g2_fill_2 FILLER_66_456 ();
 sg13g2_decap_8 FILLER_66_498 ();
 sg13g2_decap_8 FILLER_66_505 ();
 sg13g2_decap_4 FILLER_66_512 ();
 sg13g2_fill_2 FILLER_66_516 ();
 sg13g2_decap_4 FILLER_66_523 ();
 sg13g2_fill_2 FILLER_66_530 ();
 sg13g2_fill_1 FILLER_66_532 ();
 sg13g2_fill_1 FILLER_66_538 ();
 sg13g2_decap_8 FILLER_66_543 ();
 sg13g2_decap_8 FILLER_66_550 ();
 sg13g2_decap_8 FILLER_66_557 ();
 sg13g2_decap_8 FILLER_66_564 ();
 sg13g2_decap_4 FILLER_66_571 ();
 sg13g2_fill_1 FILLER_66_575 ();
 sg13g2_fill_1 FILLER_66_580 ();
 sg13g2_decap_4 FILLER_66_586 ();
 sg13g2_fill_1 FILLER_66_593 ();
 sg13g2_fill_1 FILLER_66_603 ();
 sg13g2_fill_1 FILLER_66_609 ();
 sg13g2_decap_8 FILLER_66_614 ();
 sg13g2_decap_8 FILLER_66_621 ();
 sg13g2_fill_2 FILLER_66_628 ();
 sg13g2_decap_8 FILLER_66_660 ();
 sg13g2_decap_8 FILLER_66_667 ();
 sg13g2_decap_8 FILLER_66_674 ();
 sg13g2_decap_8 FILLER_66_681 ();
 sg13g2_decap_8 FILLER_66_688 ();
 sg13g2_decap_8 FILLER_66_695 ();
 sg13g2_decap_8 FILLER_66_702 ();
 sg13g2_decap_8 FILLER_66_709 ();
 sg13g2_decap_8 FILLER_66_716 ();
 sg13g2_decap_8 FILLER_66_723 ();
 sg13g2_decap_8 FILLER_66_730 ();
 sg13g2_decap_8 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_744 ();
 sg13g2_decap_8 FILLER_66_751 ();
 sg13g2_decap_8 FILLER_66_758 ();
 sg13g2_decap_8 FILLER_66_765 ();
 sg13g2_decap_8 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_decap_8 FILLER_66_786 ();
 sg13g2_decap_8 FILLER_66_793 ();
 sg13g2_decap_8 FILLER_66_800 ();
 sg13g2_decap_8 FILLER_66_807 ();
 sg13g2_decap_8 FILLER_66_814 ();
 sg13g2_decap_8 FILLER_66_821 ();
 sg13g2_decap_8 FILLER_66_828 ();
 sg13g2_decap_8 FILLER_66_835 ();
 sg13g2_decap_8 FILLER_66_842 ();
 sg13g2_decap_8 FILLER_66_849 ();
 sg13g2_decap_8 FILLER_66_856 ();
 sg13g2_decap_8 FILLER_66_863 ();
 sg13g2_decap_8 FILLER_66_870 ();
 sg13g2_fill_1 FILLER_66_877 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_fill_2 FILLER_67_42 ();
 sg13g2_fill_2 FILLER_67_60 ();
 sg13g2_fill_1 FILLER_67_70 ();
 sg13g2_fill_1 FILLER_67_88 ();
 sg13g2_fill_2 FILLER_67_123 ();
 sg13g2_fill_1 FILLER_67_125 ();
 sg13g2_decap_8 FILLER_67_129 ();
 sg13g2_fill_2 FILLER_67_136 ();
 sg13g2_decap_8 FILLER_67_150 ();
 sg13g2_decap_8 FILLER_67_157 ();
 sg13g2_decap_8 FILLER_67_164 ();
 sg13g2_decap_8 FILLER_67_171 ();
 sg13g2_decap_8 FILLER_67_178 ();
 sg13g2_decap_8 FILLER_67_185 ();
 sg13g2_decap_8 FILLER_67_192 ();
 sg13g2_decap_8 FILLER_67_199 ();
 sg13g2_decap_8 FILLER_67_206 ();
 sg13g2_decap_8 FILLER_67_213 ();
 sg13g2_decap_8 FILLER_67_220 ();
 sg13g2_decap_8 FILLER_67_227 ();
 sg13g2_fill_2 FILLER_67_234 ();
 sg13g2_fill_1 FILLER_67_236 ();
 sg13g2_decap_8 FILLER_67_241 ();
 sg13g2_decap_4 FILLER_67_248 ();
 sg13g2_fill_1 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_257 ();
 sg13g2_decap_8 FILLER_67_264 ();
 sg13g2_decap_8 FILLER_67_271 ();
 sg13g2_decap_8 FILLER_67_278 ();
 sg13g2_decap_4 FILLER_67_285 ();
 sg13g2_decap_4 FILLER_67_323 ();
 sg13g2_fill_1 FILLER_67_327 ();
 sg13g2_decap_4 FILLER_67_333 ();
 sg13g2_fill_2 FILLER_67_337 ();
 sg13g2_decap_4 FILLER_67_343 ();
 sg13g2_fill_1 FILLER_67_347 ();
 sg13g2_decap_8 FILLER_67_354 ();
 sg13g2_decap_8 FILLER_67_361 ();
 sg13g2_decap_8 FILLER_67_368 ();
 sg13g2_fill_2 FILLER_67_375 ();
 sg13g2_decap_8 FILLER_67_381 ();
 sg13g2_decap_8 FILLER_67_388 ();
 sg13g2_fill_2 FILLER_67_395 ();
 sg13g2_fill_1 FILLER_67_397 ();
 sg13g2_fill_2 FILLER_67_401 ();
 sg13g2_decap_8 FILLER_67_433 ();
 sg13g2_decap_8 FILLER_67_440 ();
 sg13g2_decap_8 FILLER_67_447 ();
 sg13g2_decap_8 FILLER_67_454 ();
 sg13g2_decap_4 FILLER_67_461 ();
 sg13g2_fill_1 FILLER_67_465 ();
 sg13g2_fill_1 FILLER_67_483 ();
 sg13g2_decap_8 FILLER_67_492 ();
 sg13g2_decap_8 FILLER_67_499 ();
 sg13g2_decap_8 FILLER_67_506 ();
 sg13g2_decap_8 FILLER_67_513 ();
 sg13g2_decap_8 FILLER_67_520 ();
 sg13g2_decap_8 FILLER_67_527 ();
 sg13g2_decap_8 FILLER_67_534 ();
 sg13g2_decap_8 FILLER_67_541 ();
 sg13g2_decap_8 FILLER_67_548 ();
 sg13g2_decap_8 FILLER_67_555 ();
 sg13g2_decap_8 FILLER_67_562 ();
 sg13g2_decap_8 FILLER_67_569 ();
 sg13g2_decap_8 FILLER_67_576 ();
 sg13g2_decap_8 FILLER_67_583 ();
 sg13g2_decap_8 FILLER_67_590 ();
 sg13g2_decap_8 FILLER_67_597 ();
 sg13g2_decap_8 FILLER_67_604 ();
 sg13g2_decap_8 FILLER_67_611 ();
 sg13g2_decap_8 FILLER_67_618 ();
 sg13g2_fill_2 FILLER_67_625 ();
 sg13g2_fill_2 FILLER_67_631 ();
 sg13g2_decap_8 FILLER_67_668 ();
 sg13g2_decap_8 FILLER_67_675 ();
 sg13g2_decap_8 FILLER_67_682 ();
 sg13g2_decap_8 FILLER_67_689 ();
 sg13g2_decap_8 FILLER_67_696 ();
 sg13g2_decap_8 FILLER_67_703 ();
 sg13g2_decap_8 FILLER_67_710 ();
 sg13g2_decap_8 FILLER_67_717 ();
 sg13g2_decap_8 FILLER_67_724 ();
 sg13g2_decap_8 FILLER_67_731 ();
 sg13g2_decap_8 FILLER_67_738 ();
 sg13g2_decap_8 FILLER_67_745 ();
 sg13g2_decap_8 FILLER_67_752 ();
 sg13g2_decap_8 FILLER_67_759 ();
 sg13g2_decap_8 FILLER_67_766 ();
 sg13g2_decap_8 FILLER_67_773 ();
 sg13g2_decap_8 FILLER_67_780 ();
 sg13g2_decap_8 FILLER_67_787 ();
 sg13g2_decap_8 FILLER_67_794 ();
 sg13g2_decap_8 FILLER_67_801 ();
 sg13g2_decap_8 FILLER_67_808 ();
 sg13g2_decap_8 FILLER_67_815 ();
 sg13g2_decap_8 FILLER_67_822 ();
 sg13g2_decap_8 FILLER_67_829 ();
 sg13g2_decap_8 FILLER_67_836 ();
 sg13g2_decap_8 FILLER_67_843 ();
 sg13g2_decap_8 FILLER_67_850 ();
 sg13g2_decap_8 FILLER_67_857 ();
 sg13g2_decap_8 FILLER_67_864 ();
 sg13g2_decap_8 FILLER_67_871 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_fill_2 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_37 ();
 sg13g2_fill_2 FILLER_68_59 ();
 sg13g2_decap_4 FILLER_68_79 ();
 sg13g2_fill_1 FILLER_68_88 ();
 sg13g2_decap_8 FILLER_68_106 ();
 sg13g2_decap_4 FILLER_68_113 ();
 sg13g2_decap_4 FILLER_68_122 ();
 sg13g2_decap_8 FILLER_68_162 ();
 sg13g2_decap_8 FILLER_68_169 ();
 sg13g2_decap_8 FILLER_68_176 ();
 sg13g2_decap_8 FILLER_68_183 ();
 sg13g2_decap_8 FILLER_68_190 ();
 sg13g2_fill_1 FILLER_68_197 ();
 sg13g2_decap_8 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_231 ();
 sg13g2_decap_8 FILLER_68_238 ();
 sg13g2_fill_2 FILLER_68_245 ();
 sg13g2_fill_1 FILLER_68_247 ();
 sg13g2_decap_8 FILLER_68_274 ();
 sg13g2_fill_1 FILLER_68_281 ();
 sg13g2_decap_8 FILLER_68_308 ();
 sg13g2_decap_8 FILLER_68_315 ();
 sg13g2_decap_8 FILLER_68_322 ();
 sg13g2_fill_2 FILLER_68_329 ();
 sg13g2_fill_1 FILLER_68_331 ();
 sg13g2_decap_8 FILLER_68_358 ();
 sg13g2_decap_8 FILLER_68_365 ();
 sg13g2_decap_8 FILLER_68_372 ();
 sg13g2_decap_8 FILLER_68_379 ();
 sg13g2_decap_8 FILLER_68_386 ();
 sg13g2_decap_4 FILLER_68_393 ();
 sg13g2_fill_1 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_68_425 ();
 sg13g2_decap_8 FILLER_68_432 ();
 sg13g2_decap_8 FILLER_68_439 ();
 sg13g2_decap_8 FILLER_68_446 ();
 sg13g2_decap_8 FILLER_68_453 ();
 sg13g2_decap_8 FILLER_68_460 ();
 sg13g2_decap_8 FILLER_68_467 ();
 sg13g2_decap_8 FILLER_68_474 ();
 sg13g2_decap_8 FILLER_68_481 ();
 sg13g2_decap_8 FILLER_68_488 ();
 sg13g2_decap_8 FILLER_68_495 ();
 sg13g2_decap_8 FILLER_68_502 ();
 sg13g2_decap_8 FILLER_68_509 ();
 sg13g2_decap_8 FILLER_68_516 ();
 sg13g2_decap_8 FILLER_68_523 ();
 sg13g2_decap_8 FILLER_68_530 ();
 sg13g2_decap_8 FILLER_68_537 ();
 sg13g2_decap_8 FILLER_68_544 ();
 sg13g2_decap_8 FILLER_68_551 ();
 sg13g2_decap_8 FILLER_68_558 ();
 sg13g2_decap_8 FILLER_68_565 ();
 sg13g2_decap_8 FILLER_68_572 ();
 sg13g2_decap_8 FILLER_68_579 ();
 sg13g2_decap_8 FILLER_68_586 ();
 sg13g2_decap_8 FILLER_68_593 ();
 sg13g2_decap_8 FILLER_68_600 ();
 sg13g2_decap_8 FILLER_68_607 ();
 sg13g2_decap_8 FILLER_68_614 ();
 sg13g2_decap_8 FILLER_68_621 ();
 sg13g2_fill_2 FILLER_68_628 ();
 sg13g2_fill_1 FILLER_68_630 ();
 sg13g2_decap_4 FILLER_68_646 ();
 sg13g2_decap_8 FILLER_68_654 ();
 sg13g2_decap_8 FILLER_68_661 ();
 sg13g2_decap_8 FILLER_68_668 ();
 sg13g2_decap_8 FILLER_68_675 ();
 sg13g2_decap_8 FILLER_68_682 ();
 sg13g2_decap_8 FILLER_68_689 ();
 sg13g2_decap_8 FILLER_68_696 ();
 sg13g2_decap_8 FILLER_68_703 ();
 sg13g2_decap_8 FILLER_68_710 ();
 sg13g2_decap_8 FILLER_68_717 ();
 sg13g2_decap_8 FILLER_68_724 ();
 sg13g2_decap_8 FILLER_68_731 ();
 sg13g2_decap_8 FILLER_68_738 ();
 sg13g2_decap_8 FILLER_68_745 ();
 sg13g2_decap_8 FILLER_68_752 ();
 sg13g2_decap_8 FILLER_68_759 ();
 sg13g2_decap_8 FILLER_68_766 ();
 sg13g2_decap_8 FILLER_68_773 ();
 sg13g2_decap_8 FILLER_68_780 ();
 sg13g2_decap_8 FILLER_68_787 ();
 sg13g2_decap_8 FILLER_68_794 ();
 sg13g2_decap_8 FILLER_68_801 ();
 sg13g2_decap_8 FILLER_68_808 ();
 sg13g2_decap_8 FILLER_68_815 ();
 sg13g2_decap_8 FILLER_68_822 ();
 sg13g2_decap_8 FILLER_68_829 ();
 sg13g2_decap_8 FILLER_68_836 ();
 sg13g2_decap_8 FILLER_68_843 ();
 sg13g2_decap_8 FILLER_68_850 ();
 sg13g2_decap_8 FILLER_68_857 ();
 sg13g2_decap_8 FILLER_68_864 ();
 sg13g2_decap_8 FILLER_68_871 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_fill_2 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_58 ();
 sg13g2_fill_1 FILLER_69_65 ();
 sg13g2_fill_1 FILLER_69_69 ();
 sg13g2_fill_2 FILLER_69_74 ();
 sg13g2_fill_2 FILLER_69_81 ();
 sg13g2_decap_8 FILLER_69_102 ();
 sg13g2_decap_8 FILLER_69_109 ();
 sg13g2_decap_8 FILLER_69_116 ();
 sg13g2_fill_2 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_125 ();
 sg13g2_fill_2 FILLER_69_153 ();
 sg13g2_decap_8 FILLER_69_160 ();
 sg13g2_decap_8 FILLER_69_167 ();
 sg13g2_decap_8 FILLER_69_174 ();
 sg13g2_decap_8 FILLER_69_181 ();
 sg13g2_decap_8 FILLER_69_188 ();
 sg13g2_decap_8 FILLER_69_195 ();
 sg13g2_fill_1 FILLER_69_202 ();
 sg13g2_decap_8 FILLER_69_207 ();
 sg13g2_decap_8 FILLER_69_214 ();
 sg13g2_decap_8 FILLER_69_221 ();
 sg13g2_decap_8 FILLER_69_228 ();
 sg13g2_decap_8 FILLER_69_235 ();
 sg13g2_decap_8 FILLER_69_242 ();
 sg13g2_decap_8 FILLER_69_249 ();
 sg13g2_decap_8 FILLER_69_256 ();
 sg13g2_decap_8 FILLER_69_263 ();
 sg13g2_decap_8 FILLER_69_270 ();
 sg13g2_decap_8 FILLER_69_277 ();
 sg13g2_decap_8 FILLER_69_284 ();
 sg13g2_decap_8 FILLER_69_291 ();
 sg13g2_decap_8 FILLER_69_298 ();
 sg13g2_decap_8 FILLER_69_305 ();
 sg13g2_decap_8 FILLER_69_312 ();
 sg13g2_decap_8 FILLER_69_319 ();
 sg13g2_decap_8 FILLER_69_326 ();
 sg13g2_decap_8 FILLER_69_333 ();
 sg13g2_decap_8 FILLER_69_340 ();
 sg13g2_decap_8 FILLER_69_347 ();
 sg13g2_decap_8 FILLER_69_354 ();
 sg13g2_decap_8 FILLER_69_361 ();
 sg13g2_decap_8 FILLER_69_368 ();
 sg13g2_fill_2 FILLER_69_375 ();
 sg13g2_fill_1 FILLER_69_377 ();
 sg13g2_fill_2 FILLER_69_382 ();
 sg13g2_decap_4 FILLER_69_387 ();
 sg13g2_decap_8 FILLER_69_417 ();
 sg13g2_decap_8 FILLER_69_424 ();
 sg13g2_decap_8 FILLER_69_431 ();
 sg13g2_decap_8 FILLER_69_438 ();
 sg13g2_decap_8 FILLER_69_445 ();
 sg13g2_decap_8 FILLER_69_452 ();
 sg13g2_decap_8 FILLER_69_459 ();
 sg13g2_decap_8 FILLER_69_466 ();
 sg13g2_decap_8 FILLER_69_473 ();
 sg13g2_decap_8 FILLER_69_480 ();
 sg13g2_decap_8 FILLER_69_487 ();
 sg13g2_decap_8 FILLER_69_494 ();
 sg13g2_decap_8 FILLER_69_501 ();
 sg13g2_fill_1 FILLER_69_508 ();
 sg13g2_decap_8 FILLER_69_518 ();
 sg13g2_decap_8 FILLER_69_525 ();
 sg13g2_decap_4 FILLER_69_532 ();
 sg13g2_decap_8 FILLER_69_540 ();
 sg13g2_decap_8 FILLER_69_547 ();
 sg13g2_decap_8 FILLER_69_554 ();
 sg13g2_decap_8 FILLER_69_561 ();
 sg13g2_decap_8 FILLER_69_568 ();
 sg13g2_decap_8 FILLER_69_575 ();
 sg13g2_decap_8 FILLER_69_582 ();
 sg13g2_decap_8 FILLER_69_589 ();
 sg13g2_decap_8 FILLER_69_596 ();
 sg13g2_decap_8 FILLER_69_603 ();
 sg13g2_decap_8 FILLER_69_610 ();
 sg13g2_decap_8 FILLER_69_617 ();
 sg13g2_decap_4 FILLER_69_624 ();
 sg13g2_fill_2 FILLER_69_628 ();
 sg13g2_decap_8 FILLER_69_633 ();
 sg13g2_decap_8 FILLER_69_640 ();
 sg13g2_decap_8 FILLER_69_647 ();
 sg13g2_decap_8 FILLER_69_654 ();
 sg13g2_decap_8 FILLER_69_661 ();
 sg13g2_decap_8 FILLER_69_668 ();
 sg13g2_decap_8 FILLER_69_675 ();
 sg13g2_decap_8 FILLER_69_682 ();
 sg13g2_decap_8 FILLER_69_689 ();
 sg13g2_decap_8 FILLER_69_696 ();
 sg13g2_decap_8 FILLER_69_703 ();
 sg13g2_decap_8 FILLER_69_710 ();
 sg13g2_decap_8 FILLER_69_717 ();
 sg13g2_decap_8 FILLER_69_724 ();
 sg13g2_decap_8 FILLER_69_731 ();
 sg13g2_decap_8 FILLER_69_738 ();
 sg13g2_decap_8 FILLER_69_745 ();
 sg13g2_decap_8 FILLER_69_752 ();
 sg13g2_decap_8 FILLER_69_759 ();
 sg13g2_decap_8 FILLER_69_766 ();
 sg13g2_decap_8 FILLER_69_773 ();
 sg13g2_decap_8 FILLER_69_780 ();
 sg13g2_decap_8 FILLER_69_787 ();
 sg13g2_decap_8 FILLER_69_794 ();
 sg13g2_decap_8 FILLER_69_801 ();
 sg13g2_decap_8 FILLER_69_808 ();
 sg13g2_decap_8 FILLER_69_815 ();
 sg13g2_decap_8 FILLER_69_822 ();
 sg13g2_decap_8 FILLER_69_829 ();
 sg13g2_decap_8 FILLER_69_836 ();
 sg13g2_decap_8 FILLER_69_843 ();
 sg13g2_decap_8 FILLER_69_850 ();
 sg13g2_decap_8 FILLER_69_857 ();
 sg13g2_decap_8 FILLER_69_864 ();
 sg13g2_decap_8 FILLER_69_871 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_fill_1 FILLER_70_42 ();
 sg13g2_decap_4 FILLER_70_46 ();
 sg13g2_decap_8 FILLER_70_55 ();
 sg13g2_fill_1 FILLER_70_67 ();
 sg13g2_fill_1 FILLER_70_72 ();
 sg13g2_fill_1 FILLER_70_79 ();
 sg13g2_fill_1 FILLER_70_85 ();
 sg13g2_fill_1 FILLER_70_101 ();
 sg13g2_decap_8 FILLER_70_106 ();
 sg13g2_decap_4 FILLER_70_113 ();
 sg13g2_fill_1 FILLER_70_117 ();
 sg13g2_fill_1 FILLER_70_122 ();
 sg13g2_fill_1 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_145 ();
 sg13g2_fill_2 FILLER_70_156 ();
 sg13g2_decap_8 FILLER_70_162 ();
 sg13g2_decap_8 FILLER_70_169 ();
 sg13g2_decap_8 FILLER_70_176 ();
 sg13g2_decap_8 FILLER_70_183 ();
 sg13g2_decap_8 FILLER_70_190 ();
 sg13g2_decap_8 FILLER_70_197 ();
 sg13g2_decap_8 FILLER_70_204 ();
 sg13g2_decap_4 FILLER_70_211 ();
 sg13g2_fill_2 FILLER_70_215 ();
 sg13g2_decap_8 FILLER_70_243 ();
 sg13g2_decap_4 FILLER_70_250 ();
 sg13g2_fill_1 FILLER_70_254 ();
 sg13g2_fill_2 FILLER_70_259 ();
 sg13g2_fill_1 FILLER_70_261 ();
 sg13g2_decap_8 FILLER_70_267 ();
 sg13g2_decap_8 FILLER_70_281 ();
 sg13g2_decap_8 FILLER_70_288 ();
 sg13g2_decap_8 FILLER_70_295 ();
 sg13g2_decap_8 FILLER_70_302 ();
 sg13g2_decap_8 FILLER_70_309 ();
 sg13g2_decap_8 FILLER_70_316 ();
 sg13g2_decap_8 FILLER_70_323 ();
 sg13g2_fill_1 FILLER_70_330 ();
 sg13g2_decap_8 FILLER_70_334 ();
 sg13g2_decap_8 FILLER_70_341 ();
 sg13g2_decap_4 FILLER_70_352 ();
 sg13g2_fill_1 FILLER_70_356 ();
 sg13g2_fill_2 FILLER_70_361 ();
 sg13g2_fill_1 FILLER_70_363 ();
 sg13g2_decap_4 FILLER_70_369 ();
 sg13g2_decap_4 FILLER_70_377 ();
 sg13g2_fill_1 FILLER_70_381 ();
 sg13g2_fill_2 FILLER_70_395 ();
 sg13g2_decap_8 FILLER_70_416 ();
 sg13g2_decap_4 FILLER_70_423 ();
 sg13g2_fill_2 FILLER_70_427 ();
 sg13g2_decap_8 FILLER_70_433 ();
 sg13g2_decap_8 FILLER_70_440 ();
 sg13g2_decap_8 FILLER_70_447 ();
 sg13g2_decap_8 FILLER_70_480 ();
 sg13g2_decap_8 FILLER_70_487 ();
 sg13g2_decap_8 FILLER_70_494 ();
 sg13g2_decap_8 FILLER_70_501 ();
 sg13g2_decap_4 FILLER_70_508 ();
 sg13g2_fill_2 FILLER_70_543 ();
 sg13g2_fill_1 FILLER_70_545 ();
 sg13g2_decap_8 FILLER_70_588 ();
 sg13g2_fill_2 FILLER_70_595 ();
 sg13g2_decap_4 FILLER_70_601 ();
 sg13g2_fill_1 FILLER_70_605 ();
 sg13g2_decap_8 FILLER_70_610 ();
 sg13g2_decap_8 FILLER_70_617 ();
 sg13g2_decap_4 FILLER_70_624 ();
 sg13g2_fill_2 FILLER_70_628 ();
 sg13g2_fill_1 FILLER_70_639 ();
 sg13g2_fill_1 FILLER_70_644 ();
 sg13g2_decap_8 FILLER_70_650 ();
 sg13g2_decap_8 FILLER_70_657 ();
 sg13g2_fill_1 FILLER_70_664 ();
 sg13g2_decap_8 FILLER_70_691 ();
 sg13g2_decap_8 FILLER_70_698 ();
 sg13g2_decap_8 FILLER_70_705 ();
 sg13g2_decap_8 FILLER_70_712 ();
 sg13g2_decap_8 FILLER_70_719 ();
 sg13g2_decap_8 FILLER_70_726 ();
 sg13g2_decap_8 FILLER_70_733 ();
 sg13g2_decap_8 FILLER_70_740 ();
 sg13g2_decap_8 FILLER_70_747 ();
 sg13g2_decap_8 FILLER_70_754 ();
 sg13g2_decap_8 FILLER_70_761 ();
 sg13g2_decap_8 FILLER_70_768 ();
 sg13g2_decap_8 FILLER_70_775 ();
 sg13g2_decap_8 FILLER_70_782 ();
 sg13g2_decap_8 FILLER_70_789 ();
 sg13g2_decap_8 FILLER_70_796 ();
 sg13g2_decap_8 FILLER_70_803 ();
 sg13g2_decap_8 FILLER_70_810 ();
 sg13g2_decap_8 FILLER_70_817 ();
 sg13g2_decap_8 FILLER_70_824 ();
 sg13g2_decap_8 FILLER_70_831 ();
 sg13g2_decap_8 FILLER_70_838 ();
 sg13g2_decap_8 FILLER_70_845 ();
 sg13g2_decap_8 FILLER_70_852 ();
 sg13g2_decap_8 FILLER_70_859 ();
 sg13g2_decap_8 FILLER_70_866 ();
 sg13g2_decap_4 FILLER_70_873 ();
 sg13g2_fill_1 FILLER_70_877 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_4 FILLER_71_35 ();
 sg13g2_fill_2 FILLER_71_39 ();
 sg13g2_fill_2 FILLER_71_61 ();
 sg13g2_fill_1 FILLER_71_63 ();
 sg13g2_fill_2 FILLER_71_68 ();
 sg13g2_fill_2 FILLER_71_74 ();
 sg13g2_fill_1 FILLER_71_76 ();
 sg13g2_fill_2 FILLER_71_82 ();
 sg13g2_fill_1 FILLER_71_84 ();
 sg13g2_fill_2 FILLER_71_93 ();
 sg13g2_fill_2 FILLER_71_100 ();
 sg13g2_fill_1 FILLER_71_102 ();
 sg13g2_fill_1 FILLER_71_116 ();
 sg13g2_fill_1 FILLER_71_121 ();
 sg13g2_fill_1 FILLER_71_144 ();
 sg13g2_decap_8 FILLER_71_149 ();
 sg13g2_decap_8 FILLER_71_156 ();
 sg13g2_decap_8 FILLER_71_163 ();
 sg13g2_decap_8 FILLER_71_170 ();
 sg13g2_decap_8 FILLER_71_177 ();
 sg13g2_decap_8 FILLER_71_184 ();
 sg13g2_decap_8 FILLER_71_191 ();
 sg13g2_decap_8 FILLER_71_198 ();
 sg13g2_decap_4 FILLER_71_205 ();
 sg13g2_fill_2 FILLER_71_209 ();
 sg13g2_decap_8 FILLER_71_215 ();
 sg13g2_fill_2 FILLER_71_222 ();
 sg13g2_decap_8 FILLER_71_228 ();
 sg13g2_decap_8 FILLER_71_235 ();
 sg13g2_decap_8 FILLER_71_242 ();
 sg13g2_decap_8 FILLER_71_249 ();
 sg13g2_decap_4 FILLER_71_256 ();
 sg13g2_decap_8 FILLER_71_286 ();
 sg13g2_decap_8 FILLER_71_293 ();
 sg13g2_decap_8 FILLER_71_300 ();
 sg13g2_decap_8 FILLER_71_307 ();
 sg13g2_decap_8 FILLER_71_314 ();
 sg13g2_decap_8 FILLER_71_321 ();
 sg13g2_decap_8 FILLER_71_333 ();
 sg13g2_decap_8 FILLER_71_340 ();
 sg13g2_decap_8 FILLER_71_347 ();
 sg13g2_decap_8 FILLER_71_354 ();
 sg13g2_decap_8 FILLER_71_361 ();
 sg13g2_decap_8 FILLER_71_368 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_decap_4 FILLER_71_382 ();
 sg13g2_fill_2 FILLER_71_391 ();
 sg13g2_fill_1 FILLER_71_393 ();
 sg13g2_decap_8 FILLER_71_397 ();
 sg13g2_decap_8 FILLER_71_404 ();
 sg13g2_decap_8 FILLER_71_411 ();
 sg13g2_decap_4 FILLER_71_418 ();
 sg13g2_decap_8 FILLER_71_448 ();
 sg13g2_decap_8 FILLER_71_455 ();
 sg13g2_fill_1 FILLER_71_462 ();
 sg13g2_decap_4 FILLER_71_467 ();
 sg13g2_fill_2 FILLER_71_471 ();
 sg13g2_decap_8 FILLER_71_483 ();
 sg13g2_decap_8 FILLER_71_490 ();
 sg13g2_fill_2 FILLER_71_497 ();
 sg13g2_fill_1 FILLER_71_499 ();
 sg13g2_fill_2 FILLER_71_513 ();
 sg13g2_fill_1 FILLER_71_547 ();
 sg13g2_fill_1 FILLER_71_554 ();
 sg13g2_fill_2 FILLER_71_559 ();
 sg13g2_fill_1 FILLER_71_565 ();
 sg13g2_fill_2 FILLER_71_575 ();
 sg13g2_decap_8 FILLER_71_613 ();
 sg13g2_fill_1 FILLER_71_626 ();
 sg13g2_fill_2 FILLER_71_633 ();
 sg13g2_decap_8 FILLER_71_652 ();
 sg13g2_decap_4 FILLER_71_659 ();
 sg13g2_fill_1 FILLER_71_663 ();
 sg13g2_decap_4 FILLER_71_668 ();
 sg13g2_fill_2 FILLER_71_672 ();
 sg13g2_decap_8 FILLER_71_678 ();
 sg13g2_decap_8 FILLER_71_685 ();
 sg13g2_decap_8 FILLER_71_692 ();
 sg13g2_decap_8 FILLER_71_699 ();
 sg13g2_decap_8 FILLER_71_706 ();
 sg13g2_decap_8 FILLER_71_713 ();
 sg13g2_decap_8 FILLER_71_720 ();
 sg13g2_decap_8 FILLER_71_727 ();
 sg13g2_decap_8 FILLER_71_734 ();
 sg13g2_decap_8 FILLER_71_741 ();
 sg13g2_decap_8 FILLER_71_748 ();
 sg13g2_decap_8 FILLER_71_755 ();
 sg13g2_decap_8 FILLER_71_762 ();
 sg13g2_decap_8 FILLER_71_769 ();
 sg13g2_decap_8 FILLER_71_776 ();
 sg13g2_decap_8 FILLER_71_783 ();
 sg13g2_decap_8 FILLER_71_790 ();
 sg13g2_decap_8 FILLER_71_797 ();
 sg13g2_decap_8 FILLER_71_804 ();
 sg13g2_decap_8 FILLER_71_811 ();
 sg13g2_decap_8 FILLER_71_818 ();
 sg13g2_decap_8 FILLER_71_825 ();
 sg13g2_decap_8 FILLER_71_832 ();
 sg13g2_decap_8 FILLER_71_839 ();
 sg13g2_decap_8 FILLER_71_846 ();
 sg13g2_decap_8 FILLER_71_853 ();
 sg13g2_decap_8 FILLER_71_860 ();
 sg13g2_decap_8 FILLER_71_867 ();
 sg13g2_decap_4 FILLER_71_874 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_4 FILLER_72_35 ();
 sg13g2_fill_2 FILLER_72_39 ();
 sg13g2_fill_1 FILLER_72_52 ();
 sg13g2_fill_2 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_90 ();
 sg13g2_decap_8 FILLER_72_97 ();
 sg13g2_decap_8 FILLER_72_104 ();
 sg13g2_fill_2 FILLER_72_111 ();
 sg13g2_fill_1 FILLER_72_113 ();
 sg13g2_fill_2 FILLER_72_118 ();
 sg13g2_fill_2 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_144 ();
 sg13g2_decap_8 FILLER_72_151 ();
 sg13g2_decap_8 FILLER_72_158 ();
 sg13g2_decap_8 FILLER_72_165 ();
 sg13g2_decap_8 FILLER_72_172 ();
 sg13g2_decap_8 FILLER_72_179 ();
 sg13g2_decap_8 FILLER_72_186 ();
 sg13g2_decap_8 FILLER_72_193 ();
 sg13g2_decap_4 FILLER_72_200 ();
 sg13g2_decap_8 FILLER_72_230 ();
 sg13g2_decap_8 FILLER_72_237 ();
 sg13g2_decap_8 FILLER_72_244 ();
 sg13g2_decap_8 FILLER_72_251 ();
 sg13g2_decap_8 FILLER_72_258 ();
 sg13g2_fill_2 FILLER_72_265 ();
 sg13g2_fill_1 FILLER_72_267 ();
 sg13g2_decap_8 FILLER_72_272 ();
 sg13g2_fill_1 FILLER_72_279 ();
 sg13g2_fill_1 FILLER_72_288 ();
 sg13g2_decap_8 FILLER_72_293 ();
 sg13g2_decap_8 FILLER_72_300 ();
 sg13g2_decap_4 FILLER_72_307 ();
 sg13g2_fill_1 FILLER_72_321 ();
 sg13g2_decap_8 FILLER_72_334 ();
 sg13g2_fill_1 FILLER_72_341 ();
 sg13g2_decap_8 FILLER_72_346 ();
 sg13g2_decap_8 FILLER_72_353 ();
 sg13g2_decap_8 FILLER_72_360 ();
 sg13g2_decap_4 FILLER_72_367 ();
 sg13g2_fill_1 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_72_409 ();
 sg13g2_decap_8 FILLER_72_416 ();
 sg13g2_decap_8 FILLER_72_423 ();
 sg13g2_decap_8 FILLER_72_430 ();
 sg13g2_decap_8 FILLER_72_437 ();
 sg13g2_decap_8 FILLER_72_444 ();
 sg13g2_decap_8 FILLER_72_451 ();
 sg13g2_decap_8 FILLER_72_458 ();
 sg13g2_decap_8 FILLER_72_465 ();
 sg13g2_decap_8 FILLER_72_472 ();
 sg13g2_decap_8 FILLER_72_479 ();
 sg13g2_decap_8 FILLER_72_486 ();
 sg13g2_decap_4 FILLER_72_493 ();
 sg13g2_decap_8 FILLER_72_523 ();
 sg13g2_decap_8 FILLER_72_530 ();
 sg13g2_fill_1 FILLER_72_537 ();
 sg13g2_decap_4 FILLER_72_543 ();
 sg13g2_decap_8 FILLER_72_552 ();
 sg13g2_decap_8 FILLER_72_559 ();
 sg13g2_decap_8 FILLER_72_566 ();
 sg13g2_decap_8 FILLER_72_573 ();
 sg13g2_decap_8 FILLER_72_580 ();
 sg13g2_decap_8 FILLER_72_587 ();
 sg13g2_decap_8 FILLER_72_594 ();
 sg13g2_decap_8 FILLER_72_601 ();
 sg13g2_decap_8 FILLER_72_608 ();
 sg13g2_decap_8 FILLER_72_615 ();
 sg13g2_decap_4 FILLER_72_622 ();
 sg13g2_decap_8 FILLER_72_629 ();
 sg13g2_fill_2 FILLER_72_636 ();
 sg13g2_fill_2 FILLER_72_654 ();
 sg13g2_decap_8 FILLER_72_682 ();
 sg13g2_decap_8 FILLER_72_689 ();
 sg13g2_decap_8 FILLER_72_696 ();
 sg13g2_decap_8 FILLER_72_703 ();
 sg13g2_decap_8 FILLER_72_710 ();
 sg13g2_decap_8 FILLER_72_717 ();
 sg13g2_decap_8 FILLER_72_724 ();
 sg13g2_decap_8 FILLER_72_731 ();
 sg13g2_decap_8 FILLER_72_738 ();
 sg13g2_decap_8 FILLER_72_745 ();
 sg13g2_decap_8 FILLER_72_752 ();
 sg13g2_decap_8 FILLER_72_759 ();
 sg13g2_decap_8 FILLER_72_766 ();
 sg13g2_decap_8 FILLER_72_773 ();
 sg13g2_decap_8 FILLER_72_780 ();
 sg13g2_decap_8 FILLER_72_787 ();
 sg13g2_decap_8 FILLER_72_794 ();
 sg13g2_decap_8 FILLER_72_801 ();
 sg13g2_decap_8 FILLER_72_808 ();
 sg13g2_decap_8 FILLER_72_815 ();
 sg13g2_decap_8 FILLER_72_822 ();
 sg13g2_decap_8 FILLER_72_829 ();
 sg13g2_decap_8 FILLER_72_836 ();
 sg13g2_decap_8 FILLER_72_843 ();
 sg13g2_decap_8 FILLER_72_850 ();
 sg13g2_decap_8 FILLER_72_857 ();
 sg13g2_decap_8 FILLER_72_864 ();
 sg13g2_decap_8 FILLER_72_871 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_fill_2 FILLER_73_42 ();
 sg13g2_fill_1 FILLER_73_44 ();
 sg13g2_fill_2 FILLER_73_49 ();
 sg13g2_fill_2 FILLER_73_54 ();
 sg13g2_decap_4 FILLER_73_62 ();
 sg13g2_fill_1 FILLER_73_66 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_108 ();
 sg13g2_decap_4 FILLER_73_115 ();
 sg13g2_fill_2 FILLER_73_119 ();
 sg13g2_fill_2 FILLER_73_146 ();
 sg13g2_fill_2 FILLER_73_153 ();
 sg13g2_fill_1 FILLER_73_155 ();
 sg13g2_decap_8 FILLER_73_162 ();
 sg13g2_decap_8 FILLER_73_169 ();
 sg13g2_decap_8 FILLER_73_176 ();
 sg13g2_decap_8 FILLER_73_183 ();
 sg13g2_decap_8 FILLER_73_190 ();
 sg13g2_decap_8 FILLER_73_197 ();
 sg13g2_decap_8 FILLER_73_204 ();
 sg13g2_decap_8 FILLER_73_211 ();
 sg13g2_decap_8 FILLER_73_218 ();
 sg13g2_decap_8 FILLER_73_225 ();
 sg13g2_decap_8 FILLER_73_232 ();
 sg13g2_decap_8 FILLER_73_239 ();
 sg13g2_decap_8 FILLER_73_246 ();
 sg13g2_decap_4 FILLER_73_253 ();
 sg13g2_fill_1 FILLER_73_257 ();
 sg13g2_decap_8 FILLER_73_263 ();
 sg13g2_fill_2 FILLER_73_270 ();
 sg13g2_fill_1 FILLER_73_272 ();
 sg13g2_fill_2 FILLER_73_285 ();
 sg13g2_decap_8 FILLER_73_296 ();
 sg13g2_fill_2 FILLER_73_303 ();
 sg13g2_decap_8 FILLER_73_361 ();
 sg13g2_decap_8 FILLER_73_368 ();
 sg13g2_decap_8 FILLER_73_375 ();
 sg13g2_decap_8 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_73_389 ();
 sg13g2_fill_1 FILLER_73_396 ();
 sg13g2_decap_8 FILLER_73_400 ();
 sg13g2_decap_8 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_73_414 ();
 sg13g2_decap_8 FILLER_73_421 ();
 sg13g2_decap_8 FILLER_73_428 ();
 sg13g2_decap_8 FILLER_73_435 ();
 sg13g2_decap_8 FILLER_73_442 ();
 sg13g2_decap_8 FILLER_73_449 ();
 sg13g2_decap_8 FILLER_73_456 ();
 sg13g2_decap_8 FILLER_73_463 ();
 sg13g2_decap_8 FILLER_73_470 ();
 sg13g2_decap_8 FILLER_73_477 ();
 sg13g2_decap_8 FILLER_73_484 ();
 sg13g2_decap_8 FILLER_73_491 ();
 sg13g2_decap_8 FILLER_73_498 ();
 sg13g2_decap_8 FILLER_73_505 ();
 sg13g2_decap_8 FILLER_73_512 ();
 sg13g2_decap_8 FILLER_73_519 ();
 sg13g2_decap_8 FILLER_73_526 ();
 sg13g2_fill_1 FILLER_73_533 ();
 sg13g2_decap_8 FILLER_73_539 ();
 sg13g2_decap_8 FILLER_73_546 ();
 sg13g2_decap_8 FILLER_73_553 ();
 sg13g2_decap_8 FILLER_73_560 ();
 sg13g2_decap_8 FILLER_73_567 ();
 sg13g2_decap_4 FILLER_73_574 ();
 sg13g2_fill_1 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_584 ();
 sg13g2_decap_8 FILLER_73_591 ();
 sg13g2_decap_8 FILLER_73_598 ();
 sg13g2_decap_8 FILLER_73_605 ();
 sg13g2_decap_8 FILLER_73_612 ();
 sg13g2_decap_8 FILLER_73_619 ();
 sg13g2_decap_8 FILLER_73_626 ();
 sg13g2_decap_8 FILLER_73_633 ();
 sg13g2_decap_8 FILLER_73_640 ();
 sg13g2_decap_8 FILLER_73_647 ();
 sg13g2_decap_8 FILLER_73_654 ();
 sg13g2_decap_8 FILLER_73_661 ();
 sg13g2_decap_8 FILLER_73_668 ();
 sg13g2_decap_8 FILLER_73_675 ();
 sg13g2_decap_8 FILLER_73_682 ();
 sg13g2_decap_8 FILLER_73_689 ();
 sg13g2_decap_8 FILLER_73_696 ();
 sg13g2_decap_8 FILLER_73_703 ();
 sg13g2_decap_8 FILLER_73_710 ();
 sg13g2_decap_8 FILLER_73_717 ();
 sg13g2_decap_8 FILLER_73_724 ();
 sg13g2_decap_8 FILLER_73_731 ();
 sg13g2_decap_8 FILLER_73_738 ();
 sg13g2_decap_8 FILLER_73_745 ();
 sg13g2_decap_8 FILLER_73_752 ();
 sg13g2_decap_8 FILLER_73_759 ();
 sg13g2_decap_8 FILLER_73_766 ();
 sg13g2_decap_8 FILLER_73_773 ();
 sg13g2_decap_8 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_787 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_8 FILLER_73_857 ();
 sg13g2_decap_8 FILLER_73_864 ();
 sg13g2_decap_8 FILLER_73_871 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_4 FILLER_74_42 ();
 sg13g2_decap_4 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_78 ();
 sg13g2_fill_2 FILLER_74_85 ();
 sg13g2_fill_1 FILLER_74_87 ();
 sg13g2_decap_4 FILLER_74_93 ();
 sg13g2_fill_1 FILLER_74_97 ();
 sg13g2_decap_8 FILLER_74_102 ();
 sg13g2_decap_8 FILLER_74_109 ();
 sg13g2_decap_8 FILLER_74_124 ();
 sg13g2_decap_4 FILLER_74_131 ();
 sg13g2_decap_8 FILLER_74_138 ();
 sg13g2_decap_8 FILLER_74_145 ();
 sg13g2_decap_8 FILLER_74_152 ();
 sg13g2_decap_8 FILLER_74_159 ();
 sg13g2_decap_8 FILLER_74_166 ();
 sg13g2_decap_8 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_180 ();
 sg13g2_decap_8 FILLER_74_207 ();
 sg13g2_fill_2 FILLER_74_214 ();
 sg13g2_decap_8 FILLER_74_220 ();
 sg13g2_decap_8 FILLER_74_227 ();
 sg13g2_decap_8 FILLER_74_234 ();
 sg13g2_decap_8 FILLER_74_241 ();
 sg13g2_fill_2 FILLER_74_248 ();
 sg13g2_fill_1 FILLER_74_250 ();
 sg13g2_fill_1 FILLER_74_277 ();
 sg13g2_fill_2 FILLER_74_286 ();
 sg13g2_fill_1 FILLER_74_288 ();
 sg13g2_fill_2 FILLER_74_293 ();
 sg13g2_fill_1 FILLER_74_295 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_fill_2 FILLER_74_308 ();
 sg13g2_decap_4 FILLER_74_314 ();
 sg13g2_fill_1 FILLER_74_318 ();
 sg13g2_fill_1 FILLER_74_324 ();
 sg13g2_decap_8 FILLER_74_335 ();
 sg13g2_decap_8 FILLER_74_342 ();
 sg13g2_decap_8 FILLER_74_349 ();
 sg13g2_decap_8 FILLER_74_356 ();
 sg13g2_decap_8 FILLER_74_363 ();
 sg13g2_decap_8 FILLER_74_370 ();
 sg13g2_decap_8 FILLER_74_377 ();
 sg13g2_decap_8 FILLER_74_384 ();
 sg13g2_decap_8 FILLER_74_391 ();
 sg13g2_fill_2 FILLER_74_398 ();
 sg13g2_fill_1 FILLER_74_400 ();
 sg13g2_fill_1 FILLER_74_405 ();
 sg13g2_fill_1 FILLER_74_411 ();
 sg13g2_fill_1 FILLER_74_416 ();
 sg13g2_decap_8 FILLER_74_426 ();
 sg13g2_decap_8 FILLER_74_433 ();
 sg13g2_decap_8 FILLER_74_440 ();
 sg13g2_decap_8 FILLER_74_447 ();
 sg13g2_decap_8 FILLER_74_454 ();
 sg13g2_decap_4 FILLER_74_461 ();
 sg13g2_decap_8 FILLER_74_495 ();
 sg13g2_decap_8 FILLER_74_502 ();
 sg13g2_decap_8 FILLER_74_509 ();
 sg13g2_fill_2 FILLER_74_516 ();
 sg13g2_fill_1 FILLER_74_518 ();
 sg13g2_decap_8 FILLER_74_525 ();
 sg13g2_decap_8 FILLER_74_532 ();
 sg13g2_decap_8 FILLER_74_539 ();
 sg13g2_decap_8 FILLER_74_546 ();
 sg13g2_decap_8 FILLER_74_553 ();
 sg13g2_fill_1 FILLER_74_560 ();
 sg13g2_decap_8 FILLER_74_571 ();
 sg13g2_decap_8 FILLER_74_578 ();
 sg13g2_decap_8 FILLER_74_585 ();
 sg13g2_fill_2 FILLER_74_592 ();
 sg13g2_decap_8 FILLER_74_598 ();
 sg13g2_decap_8 FILLER_74_605 ();
 sg13g2_decap_8 FILLER_74_612 ();
 sg13g2_decap_8 FILLER_74_619 ();
 sg13g2_fill_2 FILLER_74_626 ();
 sg13g2_fill_1 FILLER_74_633 ();
 sg13g2_decap_8 FILLER_74_650 ();
 sg13g2_decap_8 FILLER_74_657 ();
 sg13g2_decap_8 FILLER_74_664 ();
 sg13g2_fill_1 FILLER_74_671 ();
 sg13g2_decap_8 FILLER_74_676 ();
 sg13g2_decap_8 FILLER_74_683 ();
 sg13g2_decap_8 FILLER_74_690 ();
 sg13g2_decap_8 FILLER_74_697 ();
 sg13g2_decap_8 FILLER_74_704 ();
 sg13g2_decap_8 FILLER_74_711 ();
 sg13g2_decap_8 FILLER_74_718 ();
 sg13g2_decap_8 FILLER_74_725 ();
 sg13g2_decap_8 FILLER_74_732 ();
 sg13g2_decap_8 FILLER_74_739 ();
 sg13g2_decap_8 FILLER_74_746 ();
 sg13g2_decap_8 FILLER_74_753 ();
 sg13g2_decap_8 FILLER_74_760 ();
 sg13g2_decap_8 FILLER_74_767 ();
 sg13g2_decap_8 FILLER_74_774 ();
 sg13g2_decap_8 FILLER_74_781 ();
 sg13g2_decap_8 FILLER_74_788 ();
 sg13g2_decap_8 FILLER_74_795 ();
 sg13g2_decap_8 FILLER_74_802 ();
 sg13g2_decap_8 FILLER_74_809 ();
 sg13g2_decap_8 FILLER_74_816 ();
 sg13g2_decap_8 FILLER_74_823 ();
 sg13g2_decap_8 FILLER_74_830 ();
 sg13g2_decap_8 FILLER_74_837 ();
 sg13g2_decap_8 FILLER_74_844 ();
 sg13g2_decap_8 FILLER_74_851 ();
 sg13g2_decap_8 FILLER_74_858 ();
 sg13g2_decap_8 FILLER_74_865 ();
 sg13g2_decap_4 FILLER_74_872 ();
 sg13g2_fill_2 FILLER_74_876 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_4 FILLER_75_40 ();
 sg13g2_fill_1 FILLER_75_44 ();
 sg13g2_fill_2 FILLER_75_50 ();
 sg13g2_fill_1 FILLER_75_52 ();
 sg13g2_fill_1 FILLER_75_59 ();
 sg13g2_decap_8 FILLER_75_64 ();
 sg13g2_fill_2 FILLER_75_71 ();
 sg13g2_decap_4 FILLER_75_77 ();
 sg13g2_fill_1 FILLER_75_85 ();
 sg13g2_decap_8 FILLER_75_100 ();
 sg13g2_fill_1 FILLER_75_116 ();
 sg13g2_fill_2 FILLER_75_120 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_137 ();
 sg13g2_decap_8 FILLER_75_148 ();
 sg13g2_decap_8 FILLER_75_155 ();
 sg13g2_fill_2 FILLER_75_162 ();
 sg13g2_fill_1 FILLER_75_164 ();
 sg13g2_decap_8 FILLER_75_170 ();
 sg13g2_decap_8 FILLER_75_177 ();
 sg13g2_fill_2 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_186 ();
 sg13g2_decap_8 FILLER_75_191 ();
 sg13g2_decap_8 FILLER_75_198 ();
 sg13g2_decap_4 FILLER_75_205 ();
 sg13g2_fill_2 FILLER_75_209 ();
 sg13g2_decap_8 FILLER_75_237 ();
 sg13g2_decap_8 FILLER_75_244 ();
 sg13g2_fill_2 FILLER_75_251 ();
 sg13g2_decap_8 FILLER_75_261 ();
 sg13g2_decap_8 FILLER_75_268 ();
 sg13g2_decap_4 FILLER_75_275 ();
 sg13g2_fill_1 FILLER_75_279 ();
 sg13g2_decap_8 FILLER_75_284 ();
 sg13g2_decap_8 FILLER_75_291 ();
 sg13g2_decap_8 FILLER_75_298 ();
 sg13g2_decap_8 FILLER_75_305 ();
 sg13g2_decap_8 FILLER_75_312 ();
 sg13g2_decap_8 FILLER_75_319 ();
 sg13g2_decap_8 FILLER_75_326 ();
 sg13g2_decap_8 FILLER_75_333 ();
 sg13g2_decap_8 FILLER_75_340 ();
 sg13g2_decap_8 FILLER_75_347 ();
 sg13g2_decap_8 FILLER_75_354 ();
 sg13g2_decap_8 FILLER_75_361 ();
 sg13g2_decap_8 FILLER_75_368 ();
 sg13g2_decap_8 FILLER_75_375 ();
 sg13g2_decap_8 FILLER_75_382 ();
 sg13g2_decap_4 FILLER_75_389 ();
 sg13g2_fill_1 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_427 ();
 sg13g2_decap_8 FILLER_75_434 ();
 sg13g2_decap_8 FILLER_75_441 ();
 sg13g2_decap_8 FILLER_75_448 ();
 sg13g2_decap_8 FILLER_75_455 ();
 sg13g2_decap_8 FILLER_75_462 ();
 sg13g2_fill_2 FILLER_75_469 ();
 sg13g2_fill_1 FILLER_75_471 ();
 sg13g2_fill_2 FILLER_75_476 ();
 sg13g2_fill_1 FILLER_75_478 ();
 sg13g2_decap_4 FILLER_75_484 ();
 sg13g2_fill_1 FILLER_75_488 ();
 sg13g2_fill_1 FILLER_75_493 ();
 sg13g2_decap_8 FILLER_75_499 ();
 sg13g2_decap_8 FILLER_75_506 ();
 sg13g2_decap_8 FILLER_75_513 ();
 sg13g2_decap_8 FILLER_75_520 ();
 sg13g2_decap_8 FILLER_75_527 ();
 sg13g2_decap_8 FILLER_75_534 ();
 sg13g2_decap_8 FILLER_75_541 ();
 sg13g2_decap_4 FILLER_75_548 ();
 sg13g2_fill_1 FILLER_75_552 ();
 sg13g2_decap_4 FILLER_75_583 ();
 sg13g2_fill_2 FILLER_75_587 ();
 sg13g2_fill_2 FILLER_75_625 ();
 sg13g2_fill_2 FILLER_75_639 ();
 sg13g2_fill_1 FILLER_75_641 ();
 sg13g2_fill_1 FILLER_75_646 ();
 sg13g2_decap_8 FILLER_75_652 ();
 sg13g2_decap_4 FILLER_75_659 ();
 sg13g2_fill_2 FILLER_75_663 ();
 sg13g2_decap_8 FILLER_75_691 ();
 sg13g2_decap_8 FILLER_75_698 ();
 sg13g2_decap_8 FILLER_75_705 ();
 sg13g2_decap_8 FILLER_75_712 ();
 sg13g2_decap_8 FILLER_75_719 ();
 sg13g2_decap_8 FILLER_75_726 ();
 sg13g2_decap_8 FILLER_75_733 ();
 sg13g2_decap_8 FILLER_75_740 ();
 sg13g2_decap_8 FILLER_75_747 ();
 sg13g2_decap_8 FILLER_75_754 ();
 sg13g2_decap_8 FILLER_75_761 ();
 sg13g2_decap_8 FILLER_75_768 ();
 sg13g2_decap_8 FILLER_75_775 ();
 sg13g2_decap_8 FILLER_75_782 ();
 sg13g2_decap_8 FILLER_75_789 ();
 sg13g2_decap_8 FILLER_75_796 ();
 sg13g2_decap_8 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_810 ();
 sg13g2_decap_8 FILLER_75_817 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_decap_8 FILLER_75_859 ();
 sg13g2_decap_8 FILLER_75_866 ();
 sg13g2_decap_4 FILLER_75_873 ();
 sg13g2_fill_1 FILLER_75_877 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_fill_2 FILLER_76_35 ();
 sg13g2_fill_1 FILLER_76_37 ();
 sg13g2_fill_2 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_69 ();
 sg13g2_decap_8 FILLER_76_96 ();
 sg13g2_decap_4 FILLER_76_103 ();
 sg13g2_fill_1 FILLER_76_107 ();
 sg13g2_fill_1 FILLER_76_112 ();
 sg13g2_fill_2 FILLER_76_117 ();
 sg13g2_fill_2 FILLER_76_123 ();
 sg13g2_fill_1 FILLER_76_125 ();
 sg13g2_decap_8 FILLER_76_135 ();
 sg13g2_decap_8 FILLER_76_142 ();
 sg13g2_fill_1 FILLER_76_149 ();
 sg13g2_decap_8 FILLER_76_159 ();
 sg13g2_decap_4 FILLER_76_166 ();
 sg13g2_fill_1 FILLER_76_170 ();
 sg13g2_decap_8 FILLER_76_197 ();
 sg13g2_decap_8 FILLER_76_204 ();
 sg13g2_decap_4 FILLER_76_211 ();
 sg13g2_fill_1 FILLER_76_215 ();
 sg13g2_decap_8 FILLER_76_220 ();
 sg13g2_decap_8 FILLER_76_227 ();
 sg13g2_decap_8 FILLER_76_234 ();
 sg13g2_decap_8 FILLER_76_241 ();
 sg13g2_decap_8 FILLER_76_248 ();
 sg13g2_decap_4 FILLER_76_255 ();
 sg13g2_fill_1 FILLER_76_259 ();
 sg13g2_fill_1 FILLER_76_276 ();
 sg13g2_decap_8 FILLER_76_295 ();
 sg13g2_decap_8 FILLER_76_302 ();
 sg13g2_decap_8 FILLER_76_309 ();
 sg13g2_decap_8 FILLER_76_316 ();
 sg13g2_fill_1 FILLER_76_323 ();
 sg13g2_fill_1 FILLER_76_329 ();
 sg13g2_decap_4 FILLER_76_334 ();
 sg13g2_fill_1 FILLER_76_338 ();
 sg13g2_decap_8 FILLER_76_346 ();
 sg13g2_decap_8 FILLER_76_353 ();
 sg13g2_decap_8 FILLER_76_360 ();
 sg13g2_decap_8 FILLER_76_367 ();
 sg13g2_decap_8 FILLER_76_374 ();
 sg13g2_decap_8 FILLER_76_381 ();
 sg13g2_decap_8 FILLER_76_388 ();
 sg13g2_decap_8 FILLER_76_395 ();
 sg13g2_decap_8 FILLER_76_402 ();
 sg13g2_decap_8 FILLER_76_409 ();
 sg13g2_decap_4 FILLER_76_416 ();
 sg13g2_decap_8 FILLER_76_423 ();
 sg13g2_decap_8 FILLER_76_430 ();
 sg13g2_decap_8 FILLER_76_437 ();
 sg13g2_decap_8 FILLER_76_444 ();
 sg13g2_decap_8 FILLER_76_451 ();
 sg13g2_decap_8 FILLER_76_458 ();
 sg13g2_decap_8 FILLER_76_465 ();
 sg13g2_decap_8 FILLER_76_472 ();
 sg13g2_decap_8 FILLER_76_483 ();
 sg13g2_fill_1 FILLER_76_490 ();
 sg13g2_fill_2 FILLER_76_499 ();
 sg13g2_fill_1 FILLER_76_501 ();
 sg13g2_decap_8 FILLER_76_506 ();
 sg13g2_decap_8 FILLER_76_513 ();
 sg13g2_decap_4 FILLER_76_520 ();
 sg13g2_fill_1 FILLER_76_524 ();
 sg13g2_fill_2 FILLER_76_546 ();
 sg13g2_fill_2 FILLER_76_553 ();
 sg13g2_fill_1 FILLER_76_555 ();
 sg13g2_decap_8 FILLER_76_572 ();
 sg13g2_decap_8 FILLER_76_579 ();
 sg13g2_decap_8 FILLER_76_586 ();
 sg13g2_decap_8 FILLER_76_593 ();
 sg13g2_decap_8 FILLER_76_600 ();
 sg13g2_decap_8 FILLER_76_611 ();
 sg13g2_decap_8 FILLER_76_618 ();
 sg13g2_decap_4 FILLER_76_625 ();
 sg13g2_fill_1 FILLER_76_629 ();
 sg13g2_decap_4 FILLER_76_643 ();
 sg13g2_fill_2 FILLER_76_647 ();
 sg13g2_decap_8 FILLER_76_653 ();
 sg13g2_decap_8 FILLER_76_660 ();
 sg13g2_decap_8 FILLER_76_667 ();
 sg13g2_decap_8 FILLER_76_674 ();
 sg13g2_decap_8 FILLER_76_681 ();
 sg13g2_decap_8 FILLER_76_688 ();
 sg13g2_decap_8 FILLER_76_695 ();
 sg13g2_decap_8 FILLER_76_702 ();
 sg13g2_decap_8 FILLER_76_709 ();
 sg13g2_decap_8 FILLER_76_716 ();
 sg13g2_decap_8 FILLER_76_723 ();
 sg13g2_decap_8 FILLER_76_730 ();
 sg13g2_decap_8 FILLER_76_737 ();
 sg13g2_decap_8 FILLER_76_744 ();
 sg13g2_decap_8 FILLER_76_751 ();
 sg13g2_decap_8 FILLER_76_758 ();
 sg13g2_decap_8 FILLER_76_765 ();
 sg13g2_decap_8 FILLER_76_772 ();
 sg13g2_decap_8 FILLER_76_779 ();
 sg13g2_decap_8 FILLER_76_786 ();
 sg13g2_decap_8 FILLER_76_793 ();
 sg13g2_decap_8 FILLER_76_800 ();
 sg13g2_decap_8 FILLER_76_807 ();
 sg13g2_decap_8 FILLER_76_814 ();
 sg13g2_decap_8 FILLER_76_821 ();
 sg13g2_decap_8 FILLER_76_828 ();
 sg13g2_decap_8 FILLER_76_835 ();
 sg13g2_decap_8 FILLER_76_842 ();
 sg13g2_decap_8 FILLER_76_849 ();
 sg13g2_decap_8 FILLER_76_856 ();
 sg13g2_decap_8 FILLER_76_863 ();
 sg13g2_decap_8 FILLER_76_870 ();
 sg13g2_fill_1 FILLER_76_877 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_fill_1 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_61 ();
 sg13g2_fill_1 FILLER_77_68 ();
 sg13g2_decap_8 FILLER_77_86 ();
 sg13g2_decap_8 FILLER_77_93 ();
 sg13g2_decap_8 FILLER_77_100 ();
 sg13g2_fill_2 FILLER_77_125 ();
 sg13g2_fill_1 FILLER_77_127 ();
 sg13g2_decap_8 FILLER_77_132 ();
 sg13g2_decap_8 FILLER_77_139 ();
 sg13g2_decap_8 FILLER_77_146 ();
 sg13g2_decap_8 FILLER_77_153 ();
 sg13g2_decap_8 FILLER_77_160 ();
 sg13g2_decap_8 FILLER_77_167 ();
 sg13g2_decap_4 FILLER_77_174 ();
 sg13g2_fill_1 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_235 ();
 sg13g2_decap_8 FILLER_77_242 ();
 sg13g2_decap_8 FILLER_77_249 ();
 sg13g2_fill_2 FILLER_77_256 ();
 sg13g2_fill_1 FILLER_77_262 ();
 sg13g2_decap_8 FILLER_77_289 ();
 sg13g2_decap_8 FILLER_77_296 ();
 sg13g2_decap_8 FILLER_77_303 ();
 sg13g2_decap_8 FILLER_77_310 ();
 sg13g2_decap_4 FILLER_77_317 ();
 sg13g2_decap_8 FILLER_77_347 ();
 sg13g2_decap_4 FILLER_77_354 ();
 sg13g2_fill_2 FILLER_77_358 ();
 sg13g2_fill_2 FILLER_77_369 ();
 sg13g2_decap_8 FILLER_77_389 ();
 sg13g2_decap_8 FILLER_77_396 ();
 sg13g2_decap_8 FILLER_77_403 ();
 sg13g2_decap_8 FILLER_77_410 ();
 sg13g2_decap_4 FILLER_77_417 ();
 sg13g2_fill_1 FILLER_77_421 ();
 sg13g2_decap_4 FILLER_77_449 ();
 sg13g2_fill_2 FILLER_77_462 ();
 sg13g2_fill_1 FILLER_77_464 ();
 sg13g2_fill_1 FILLER_77_535 ();
 sg13g2_decap_8 FILLER_77_541 ();
 sg13g2_decap_8 FILLER_77_548 ();
 sg13g2_decap_4 FILLER_77_555 ();
 sg13g2_fill_2 FILLER_77_559 ();
 sg13g2_decap_8 FILLER_77_573 ();
 sg13g2_decap_8 FILLER_77_580 ();
 sg13g2_decap_8 FILLER_77_587 ();
 sg13g2_decap_8 FILLER_77_594 ();
 sg13g2_decap_8 FILLER_77_601 ();
 sg13g2_decap_4 FILLER_77_608 ();
 sg13g2_fill_1 FILLER_77_612 ();
 sg13g2_fill_1 FILLER_77_618 ();
 sg13g2_fill_2 FILLER_77_622 ();
 sg13g2_fill_1 FILLER_77_624 ();
 sg13g2_fill_2 FILLER_77_633 ();
 sg13g2_decap_8 FILLER_77_669 ();
 sg13g2_decap_8 FILLER_77_676 ();
 sg13g2_decap_8 FILLER_77_683 ();
 sg13g2_decap_8 FILLER_77_690 ();
 sg13g2_decap_8 FILLER_77_697 ();
 sg13g2_decap_8 FILLER_77_704 ();
 sg13g2_decap_8 FILLER_77_711 ();
 sg13g2_decap_8 FILLER_77_718 ();
 sg13g2_decap_8 FILLER_77_725 ();
 sg13g2_decap_8 FILLER_77_732 ();
 sg13g2_decap_8 FILLER_77_739 ();
 sg13g2_decap_8 FILLER_77_746 ();
 sg13g2_decap_8 FILLER_77_753 ();
 sg13g2_decap_8 FILLER_77_760 ();
 sg13g2_decap_8 FILLER_77_767 ();
 sg13g2_decap_8 FILLER_77_774 ();
 sg13g2_decap_8 FILLER_77_781 ();
 sg13g2_decap_8 FILLER_77_788 ();
 sg13g2_decap_8 FILLER_77_795 ();
 sg13g2_decap_8 FILLER_77_802 ();
 sg13g2_decap_8 FILLER_77_809 ();
 sg13g2_decap_8 FILLER_77_816 ();
 sg13g2_decap_8 FILLER_77_823 ();
 sg13g2_decap_8 FILLER_77_830 ();
 sg13g2_decap_8 FILLER_77_837 ();
 sg13g2_decap_8 FILLER_77_844 ();
 sg13g2_decap_8 FILLER_77_851 ();
 sg13g2_decap_8 FILLER_77_858 ();
 sg13g2_decap_8 FILLER_77_865 ();
 sg13g2_decap_4 FILLER_77_872 ();
 sg13g2_fill_2 FILLER_77_876 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_fill_1 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_41 ();
 sg13g2_decap_8 FILLER_78_50 ();
 sg13g2_decap_8 FILLER_78_57 ();
 sg13g2_fill_2 FILLER_78_64 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_4 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_128 ();
 sg13g2_decap_8 FILLER_78_135 ();
 sg13g2_decap_8 FILLER_78_142 ();
 sg13g2_decap_8 FILLER_78_149 ();
 sg13g2_decap_8 FILLER_78_156 ();
 sg13g2_decap_8 FILLER_78_163 ();
 sg13g2_decap_8 FILLER_78_170 ();
 sg13g2_decap_8 FILLER_78_177 ();
 sg13g2_decap_8 FILLER_78_184 ();
 sg13g2_decap_8 FILLER_78_195 ();
 sg13g2_decap_8 FILLER_78_202 ();
 sg13g2_fill_2 FILLER_78_209 ();
 sg13g2_fill_1 FILLER_78_211 ();
 sg13g2_decap_8 FILLER_78_216 ();
 sg13g2_decap_8 FILLER_78_223 ();
 sg13g2_decap_8 FILLER_78_230 ();
 sg13g2_decap_8 FILLER_78_237 ();
 sg13g2_decap_4 FILLER_78_244 ();
 sg13g2_fill_2 FILLER_78_248 ();
 sg13g2_fill_1 FILLER_78_258 ();
 sg13g2_decap_8 FILLER_78_289 ();
 sg13g2_decap_8 FILLER_78_296 ();
 sg13g2_decap_4 FILLER_78_303 ();
 sg13g2_fill_1 FILLER_78_307 ();
 sg13g2_decap_8 FILLER_78_312 ();
 sg13g2_decap_8 FILLER_78_319 ();
 sg13g2_fill_1 FILLER_78_326 ();
 sg13g2_decap_4 FILLER_78_331 ();
 sg13g2_fill_2 FILLER_78_335 ();
 sg13g2_fill_1 FILLER_78_364 ();
 sg13g2_fill_1 FILLER_78_374 ();
 sg13g2_fill_2 FILLER_78_384 ();
 sg13g2_decap_4 FILLER_78_395 ();
 sg13g2_fill_2 FILLER_78_399 ();
 sg13g2_fill_2 FILLER_78_419 ();
 sg13g2_fill_1 FILLER_78_421 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_4 FILLER_78_434 ();
 sg13g2_fill_2 FILLER_78_438 ();
 sg13g2_decap_8 FILLER_78_448 ();
 sg13g2_decap_4 FILLER_78_455 ();
 sg13g2_fill_2 FILLER_78_459 ();
 sg13g2_fill_2 FILLER_78_470 ();
 sg13g2_fill_1 FILLER_78_472 ();
 sg13g2_decap_8 FILLER_78_486 ();
 sg13g2_decap_8 FILLER_78_493 ();
 sg13g2_decap_8 FILLER_78_500 ();
 sg13g2_decap_4 FILLER_78_507 ();
 sg13g2_fill_1 FILLER_78_511 ();
 sg13g2_decap_8 FILLER_78_516 ();
 sg13g2_decap_8 FILLER_78_553 ();
 sg13g2_fill_2 FILLER_78_560 ();
 sg13g2_decap_8 FILLER_78_588 ();
 sg13g2_decap_8 FILLER_78_595 ();
 sg13g2_fill_2 FILLER_78_602 ();
 sg13g2_fill_1 FILLER_78_604 ();
 sg13g2_decap_4 FILLER_78_631 ();
 sg13g2_fill_2 FILLER_78_639 ();
 sg13g2_fill_1 FILLER_78_641 ();
 sg13g2_decap_8 FILLER_78_646 ();
 sg13g2_decap_8 FILLER_78_653 ();
 sg13g2_decap_8 FILLER_78_660 ();
 sg13g2_decap_8 FILLER_78_667 ();
 sg13g2_decap_8 FILLER_78_674 ();
 sg13g2_decap_8 FILLER_78_681 ();
 sg13g2_decap_8 FILLER_78_688 ();
 sg13g2_decap_8 FILLER_78_695 ();
 sg13g2_decap_8 FILLER_78_702 ();
 sg13g2_decap_8 FILLER_78_709 ();
 sg13g2_decap_8 FILLER_78_716 ();
 sg13g2_decap_8 FILLER_78_723 ();
 sg13g2_decap_8 FILLER_78_730 ();
 sg13g2_decap_8 FILLER_78_737 ();
 sg13g2_decap_8 FILLER_78_744 ();
 sg13g2_decap_8 FILLER_78_751 ();
 sg13g2_decap_8 FILLER_78_758 ();
 sg13g2_decap_8 FILLER_78_765 ();
 sg13g2_decap_8 FILLER_78_772 ();
 sg13g2_decap_8 FILLER_78_779 ();
 sg13g2_decap_8 FILLER_78_786 ();
 sg13g2_decap_8 FILLER_78_793 ();
 sg13g2_decap_8 FILLER_78_800 ();
 sg13g2_decap_8 FILLER_78_807 ();
 sg13g2_decap_8 FILLER_78_814 ();
 sg13g2_decap_8 FILLER_78_821 ();
 sg13g2_decap_8 FILLER_78_828 ();
 sg13g2_decap_8 FILLER_78_835 ();
 sg13g2_decap_8 FILLER_78_842 ();
 sg13g2_decap_8 FILLER_78_849 ();
 sg13g2_decap_8 FILLER_78_856 ();
 sg13g2_decap_8 FILLER_78_863 ();
 sg13g2_decap_8 FILLER_78_870 ();
 sg13g2_fill_1 FILLER_78_877 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_fill_2 FILLER_79_35 ();
 sg13g2_fill_1 FILLER_79_37 ();
 sg13g2_decap_8 FILLER_79_64 ();
 sg13g2_decap_8 FILLER_79_71 ();
 sg13g2_decap_8 FILLER_79_78 ();
 sg13g2_fill_2 FILLER_79_85 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_4 FILLER_79_98 ();
 sg13g2_fill_1 FILLER_79_102 ();
 sg13g2_decap_8 FILLER_79_107 ();
 sg13g2_decap_8 FILLER_79_114 ();
 sg13g2_decap_8 FILLER_79_121 ();
 sg13g2_decap_8 FILLER_79_128 ();
 sg13g2_decap_8 FILLER_79_135 ();
 sg13g2_decap_8 FILLER_79_142 ();
 sg13g2_decap_8 FILLER_79_149 ();
 sg13g2_fill_1 FILLER_79_156 ();
 sg13g2_decap_4 FILLER_79_161 ();
 sg13g2_fill_1 FILLER_79_165 ();
 sg13g2_fill_1 FILLER_79_171 ();
 sg13g2_decap_8 FILLER_79_176 ();
 sg13g2_decap_8 FILLER_79_183 ();
 sg13g2_decap_8 FILLER_79_190 ();
 sg13g2_decap_8 FILLER_79_197 ();
 sg13g2_fill_2 FILLER_79_204 ();
 sg13g2_decap_8 FILLER_79_232 ();
 sg13g2_decap_8 FILLER_79_239 ();
 sg13g2_decap_8 FILLER_79_246 ();
 sg13g2_decap_8 FILLER_79_253 ();
 sg13g2_decap_8 FILLER_79_260 ();
 sg13g2_fill_2 FILLER_79_267 ();
 sg13g2_fill_1 FILLER_79_269 ();
 sg13g2_decap_8 FILLER_79_274 ();
 sg13g2_decap_8 FILLER_79_281 ();
 sg13g2_decap_8 FILLER_79_288 ();
 sg13g2_decap_8 FILLER_79_295 ();
 sg13g2_decap_8 FILLER_79_328 ();
 sg13g2_decap_8 FILLER_79_335 ();
 sg13g2_decap_8 FILLER_79_342 ();
 sg13g2_decap_8 FILLER_79_349 ();
 sg13g2_decap_8 FILLER_79_356 ();
 sg13g2_decap_8 FILLER_79_363 ();
 sg13g2_decap_8 FILLER_79_370 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_decap_8 FILLER_79_384 ();
 sg13g2_decap_8 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_decap_8 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_79_412 ();
 sg13g2_decap_8 FILLER_79_419 ();
 sg13g2_decap_8 FILLER_79_426 ();
 sg13g2_decap_8 FILLER_79_459 ();
 sg13g2_decap_8 FILLER_79_466 ();
 sg13g2_decap_8 FILLER_79_473 ();
 sg13g2_decap_8 FILLER_79_480 ();
 sg13g2_decap_8 FILLER_79_487 ();
 sg13g2_decap_8 FILLER_79_494 ();
 sg13g2_decap_8 FILLER_79_501 ();
 sg13g2_decap_8 FILLER_79_508 ();
 sg13g2_decap_8 FILLER_79_515 ();
 sg13g2_decap_8 FILLER_79_522 ();
 sg13g2_decap_8 FILLER_79_529 ();
 sg13g2_decap_8 FILLER_79_536 ();
 sg13g2_decap_8 FILLER_79_543 ();
 sg13g2_decap_8 FILLER_79_550 ();
 sg13g2_decap_8 FILLER_79_557 ();
 sg13g2_decap_4 FILLER_79_564 ();
 sg13g2_decap_8 FILLER_79_572 ();
 sg13g2_decap_8 FILLER_79_579 ();
 sg13g2_decap_8 FILLER_79_586 ();
 sg13g2_decap_8 FILLER_79_593 ();
 sg13g2_decap_8 FILLER_79_600 ();
 sg13g2_decap_4 FILLER_79_607 ();
 sg13g2_fill_1 FILLER_79_611 ();
 sg13g2_decap_8 FILLER_79_616 ();
 sg13g2_decap_8 FILLER_79_623 ();
 sg13g2_decap_4 FILLER_79_630 ();
 sg13g2_fill_2 FILLER_79_634 ();
 sg13g2_decap_8 FILLER_79_662 ();
 sg13g2_decap_8 FILLER_79_669 ();
 sg13g2_decap_8 FILLER_79_676 ();
 sg13g2_decap_8 FILLER_79_683 ();
 sg13g2_decap_8 FILLER_79_690 ();
 sg13g2_decap_8 FILLER_79_697 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_8 FILLER_79_711 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_decap_8 FILLER_79_725 ();
 sg13g2_decap_8 FILLER_79_732 ();
 sg13g2_decap_8 FILLER_79_739 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_decap_8 FILLER_79_753 ();
 sg13g2_decap_8 FILLER_79_760 ();
 sg13g2_decap_8 FILLER_79_767 ();
 sg13g2_decap_8 FILLER_79_774 ();
 sg13g2_decap_8 FILLER_79_781 ();
 sg13g2_decap_8 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_8 FILLER_79_858 ();
 sg13g2_decap_8 FILLER_79_865 ();
 sg13g2_decap_4 FILLER_79_872 ();
 sg13g2_fill_2 FILLER_79_876 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_4 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_67 ();
 sg13g2_fill_1 FILLER_80_73 ();
 sg13g2_fill_1 FILLER_80_78 ();
 sg13g2_fill_1 FILLER_80_83 ();
 sg13g2_fill_1 FILLER_80_88 ();
 sg13g2_fill_2 FILLER_80_93 ();
 sg13g2_fill_1 FILLER_80_99 ();
 sg13g2_fill_2 FILLER_80_104 ();
 sg13g2_decap_4 FILLER_80_126 ();
 sg13g2_fill_2 FILLER_80_130 ();
 sg13g2_fill_2 FILLER_80_140 ();
 sg13g2_fill_1 FILLER_80_142 ();
 sg13g2_fill_1 FILLER_80_156 ();
 sg13g2_fill_2 FILLER_80_170 ();
 sg13g2_fill_1 FILLER_80_189 ();
 sg13g2_decap_4 FILLER_80_194 ();
 sg13g2_fill_2 FILLER_80_202 ();
 sg13g2_fill_2 FILLER_80_208 ();
 sg13g2_fill_1 FILLER_80_210 ();
 sg13g2_decap_4 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_227 ();
 sg13g2_fill_1 FILLER_80_237 ();
 sg13g2_decap_4 FILLER_80_242 ();
 sg13g2_fill_1 FILLER_80_246 ();
 sg13g2_decap_8 FILLER_80_251 ();
 sg13g2_decap_8 FILLER_80_258 ();
 sg13g2_decap_8 FILLER_80_265 ();
 sg13g2_decap_8 FILLER_80_272 ();
 sg13g2_decap_8 FILLER_80_279 ();
 sg13g2_decap_8 FILLER_80_286 ();
 sg13g2_decap_8 FILLER_80_293 ();
 sg13g2_decap_8 FILLER_80_300 ();
 sg13g2_decap_8 FILLER_80_307 ();
 sg13g2_decap_8 FILLER_80_314 ();
 sg13g2_decap_8 FILLER_80_321 ();
 sg13g2_decap_8 FILLER_80_328 ();
 sg13g2_fill_1 FILLER_80_335 ();
 sg13g2_fill_2 FILLER_80_340 ();
 sg13g2_fill_1 FILLER_80_342 ();
 sg13g2_decap_8 FILLER_80_347 ();
 sg13g2_decap_8 FILLER_80_354 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_4 FILLER_80_368 ();
 sg13g2_fill_2 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_378 ();
 sg13g2_decap_8 FILLER_80_385 ();
 sg13g2_decap_4 FILLER_80_392 ();
 sg13g2_fill_2 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_402 ();
 sg13g2_decap_8 FILLER_80_409 ();
 sg13g2_decap_8 FILLER_80_416 ();
 sg13g2_decap_8 FILLER_80_423 ();
 sg13g2_decap_8 FILLER_80_430 ();
 sg13g2_decap_8 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_444 ();
 sg13g2_decap_8 FILLER_80_451 ();
 sg13g2_decap_8 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_decap_8 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_479 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_decap_8 FILLER_80_493 ();
 sg13g2_decap_8 FILLER_80_500 ();
 sg13g2_decap_8 FILLER_80_507 ();
 sg13g2_decap_8 FILLER_80_514 ();
 sg13g2_decap_8 FILLER_80_521 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_decap_8 FILLER_80_535 ();
 sg13g2_decap_8 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_549 ();
 sg13g2_decap_8 FILLER_80_556 ();
 sg13g2_decap_8 FILLER_80_563 ();
 sg13g2_decap_8 FILLER_80_570 ();
 sg13g2_decap_8 FILLER_80_577 ();
 sg13g2_decap_8 FILLER_80_584 ();
 sg13g2_decap_8 FILLER_80_591 ();
 sg13g2_decap_8 FILLER_80_598 ();
 sg13g2_decap_8 FILLER_80_605 ();
 sg13g2_decap_8 FILLER_80_612 ();
 sg13g2_decap_8 FILLER_80_619 ();
 sg13g2_decap_8 FILLER_80_626 ();
 sg13g2_decap_8 FILLER_80_633 ();
 sg13g2_decap_8 FILLER_80_640 ();
 sg13g2_decap_8 FILLER_80_647 ();
 sg13g2_decap_8 FILLER_80_654 ();
 sg13g2_decap_8 FILLER_80_661 ();
 sg13g2_decap_8 FILLER_80_668 ();
 sg13g2_decap_8 FILLER_80_675 ();
 sg13g2_decap_8 FILLER_80_682 ();
 sg13g2_decap_8 FILLER_80_689 ();
 sg13g2_decap_8 FILLER_80_696 ();
 sg13g2_decap_8 FILLER_80_703 ();
 sg13g2_decap_8 FILLER_80_710 ();
 sg13g2_decap_8 FILLER_80_717 ();
 sg13g2_decap_8 FILLER_80_724 ();
 sg13g2_decap_8 FILLER_80_731 ();
 sg13g2_decap_8 FILLER_80_738 ();
 sg13g2_decap_8 FILLER_80_745 ();
 sg13g2_decap_8 FILLER_80_752 ();
 sg13g2_decap_8 FILLER_80_759 ();
 sg13g2_decap_8 FILLER_80_766 ();
 sg13g2_decap_8 FILLER_80_773 ();
 sg13g2_decap_8 FILLER_80_780 ();
 sg13g2_decap_8 FILLER_80_787 ();
 sg13g2_decap_8 FILLER_80_794 ();
 sg13g2_decap_8 FILLER_80_801 ();
 sg13g2_decap_8 FILLER_80_808 ();
 sg13g2_decap_8 FILLER_80_815 ();
 sg13g2_decap_8 FILLER_80_822 ();
 sg13g2_decap_8 FILLER_80_829 ();
 sg13g2_decap_8 FILLER_80_836 ();
 sg13g2_decap_8 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_850 ();
 sg13g2_decap_8 FILLER_80_857 ();
 sg13g2_decap_8 FILLER_80_864 ();
 sg13g2_decap_8 FILLER_80_871 ();
endmodule
