module tt_um_pulse_generator (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire clknet_0_clk;
 wire \pulse_gen_inst.count_counter[0] ;
 wire \pulse_gen_inst.count_counter[10] ;
 wire \pulse_gen_inst.count_counter[11] ;
 wire \pulse_gen_inst.count_counter[12] ;
 wire \pulse_gen_inst.count_counter[13] ;
 wire \pulse_gen_inst.count_counter[14] ;
 wire \pulse_gen_inst.count_counter[15] ;
 wire \pulse_gen_inst.count_counter[1] ;
 wire \pulse_gen_inst.count_counter[2] ;
 wire \pulse_gen_inst.count_counter[3] ;
 wire \pulse_gen_inst.count_counter[4] ;
 wire \pulse_gen_inst.count_counter[5] ;
 wire \pulse_gen_inst.count_counter[6] ;
 wire \pulse_gen_inst.count_counter[7] ;
 wire \pulse_gen_inst.count_counter[8] ;
 wire \pulse_gen_inst.count_counter[9] ;
 wire \pulse_gen_inst.period_counter[0] ;
 wire \pulse_gen_inst.period_counter[10] ;
 wire \pulse_gen_inst.period_counter[11] ;
 wire \pulse_gen_inst.period_counter[12] ;
 wire \pulse_gen_inst.period_counter[13] ;
 wire \pulse_gen_inst.period_counter[14] ;
 wire \pulse_gen_inst.period_counter[15] ;
 wire \pulse_gen_inst.period_counter[16] ;
 wire \pulse_gen_inst.period_counter[17] ;
 wire \pulse_gen_inst.period_counter[18] ;
 wire \pulse_gen_inst.period_counter[19] ;
 wire \pulse_gen_inst.period_counter[1] ;
 wire \pulse_gen_inst.period_counter[20] ;
 wire \pulse_gen_inst.period_counter[21] ;
 wire \pulse_gen_inst.period_counter[22] ;
 wire \pulse_gen_inst.period_counter[23] ;
 wire \pulse_gen_inst.period_counter[24] ;
 wire \pulse_gen_inst.period_counter[25] ;
 wire \pulse_gen_inst.period_counter[26] ;
 wire \pulse_gen_inst.period_counter[27] ;
 wire \pulse_gen_inst.period_counter[28] ;
 wire \pulse_gen_inst.period_counter[29] ;
 wire \pulse_gen_inst.period_counter[2] ;
 wire \pulse_gen_inst.period_counter[30] ;
 wire \pulse_gen_inst.period_counter[31] ;
 wire \pulse_gen_inst.period_counter[3] ;
 wire \pulse_gen_inst.period_counter[4] ;
 wire \pulse_gen_inst.period_counter[5] ;
 wire \pulse_gen_inst.period_counter[6] ;
 wire \pulse_gen_inst.period_counter[7] ;
 wire \pulse_gen_inst.period_counter[8] ;
 wire \pulse_gen_inst.period_counter[9] ;
 wire \pulse_gen_inst.pulse_active ;
 wire \pulse_gen_inst.pulse_counter[0] ;
 wire \pulse_gen_inst.pulse_counter[10] ;
 wire \pulse_gen_inst.pulse_counter[11] ;
 wire \pulse_gen_inst.pulse_counter[12] ;
 wire \pulse_gen_inst.pulse_counter[13] ;
 wire \pulse_gen_inst.pulse_counter[14] ;
 wire \pulse_gen_inst.pulse_counter[15] ;
 wire \pulse_gen_inst.pulse_counter[16] ;
 wire \pulse_gen_inst.pulse_counter[17] ;
 wire \pulse_gen_inst.pulse_counter[18] ;
 wire \pulse_gen_inst.pulse_counter[19] ;
 wire \pulse_gen_inst.pulse_counter[1] ;
 wire \pulse_gen_inst.pulse_counter[20] ;
 wire \pulse_gen_inst.pulse_counter[21] ;
 wire \pulse_gen_inst.pulse_counter[22] ;
 wire \pulse_gen_inst.pulse_counter[23] ;
 wire \pulse_gen_inst.pulse_counter[24] ;
 wire \pulse_gen_inst.pulse_counter[25] ;
 wire \pulse_gen_inst.pulse_counter[26] ;
 wire \pulse_gen_inst.pulse_counter[27] ;
 wire \pulse_gen_inst.pulse_counter[28] ;
 wire \pulse_gen_inst.pulse_counter[29] ;
 wire \pulse_gen_inst.pulse_counter[2] ;
 wire \pulse_gen_inst.pulse_counter[30] ;
 wire \pulse_gen_inst.pulse_counter[31] ;
 wire \pulse_gen_inst.pulse_counter[3] ;
 wire \pulse_gen_inst.pulse_counter[4] ;
 wire \pulse_gen_inst.pulse_counter[5] ;
 wire \pulse_gen_inst.pulse_counter[6] ;
 wire \pulse_gen_inst.pulse_counter[7] ;
 wire \pulse_gen_inst.pulse_counter[8] ;
 wire \pulse_gen_inst.pulse_counter[9] ;
 wire \pulse_gen_inst.ttl_out ;
 wire \reg_sequence_select[0] ;
 wire \reg_sequence_select[1] ;
 wire \reg_sequence_select[2] ;
 wire \reg_sequence_select[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _0647_ (.A(\pulse_gen_inst.pulse_active ),
    .X(_0100_));
 sg13g2_buf_1 _0648_ (.A(net36),
    .X(_0101_));
 sg13g2_buf_2 _0649_ (.A(\pulse_gen_inst.period_counter[11] ),
    .X(_0102_));
 sg13g2_inv_1 _0650_ (.Y(_0103_),
    .A(_0102_));
 sg13g2_buf_1 _0651_ (.A(\reg_sequence_select[1] ),
    .X(_0104_));
 sg13g2_nor2b_1 _0652_ (.A(_0002_),
    .B_N(net35),
    .Y(_0105_));
 sg13g2_buf_2 _0653_ (.A(\reg_sequence_select[0] ),
    .X(_0106_));
 sg13g2_buf_8 _0654_ (.A(\reg_sequence_select[3] ),
    .X(_0107_));
 sg13g2_buf_8 _0655_ (.A(_0107_),
    .X(_0108_));
 sg13g2_nor2_1 _0656_ (.A(_0106_),
    .B(_0108_),
    .Y(_0109_));
 sg13g2_nor2b_1 _0657_ (.A(_0106_),
    .B_N(_0107_),
    .Y(_0110_));
 sg13g2_buf_8 _0658_ (.A(\reg_sequence_select[2] ),
    .X(_0111_));
 sg13g2_nand2_1 _0659_ (.Y(_0112_),
    .A(net35),
    .B(net34));
 sg13g2_a22oi_1 _0660_ (.Y(_0113_),
    .B1(_0110_),
    .B2(_0112_),
    .A2(_0109_),
    .A1(_0105_));
 sg13g2_inv_1 _0661_ (.Y(_0114_),
    .A(_0113_));
 sg13g2_buf_8 _0662_ (.A(_0106_),
    .X(_0115_));
 sg13g2_inv_1 _0663_ (.Y(_0116_),
    .A(net35));
 sg13g2_and2_1 _0664_ (.A(net34),
    .B(_0107_),
    .X(_0117_));
 sg13g2_nor3_1 _0665_ (.A(net29),
    .B(_0116_),
    .C(_0117_),
    .Y(_0118_));
 sg13g2_nand3b_1 _0666_ (.B(net34),
    .C(net30),
    .Y(_0119_),
    .A_N(net35));
 sg13g2_nand2b_1 _0667_ (.Y(_0120_),
    .B(_0002_),
    .A_N(net30));
 sg13g2_inv_2 _0668_ (.Y(_0121_),
    .A(_0106_));
 sg13g2_a21oi_1 _0669_ (.A1(_0119_),
    .A2(_0120_),
    .Y(_0122_),
    .B1(_0121_));
 sg13g2_o21ai_1 _0670_ (.B1(\pulse_gen_inst.period_counter[9] ),
    .Y(_0123_),
    .A1(_0118_),
    .A2(_0122_));
 sg13g2_inv_1 _0671_ (.Y(_0124_),
    .A(_0005_));
 sg13g2_nor3_1 _0672_ (.A(_0124_),
    .B(_0118_),
    .C(_0122_),
    .Y(_0125_));
 sg13g2_o21ai_1 _0673_ (.B1(_0124_),
    .Y(_0126_),
    .A1(_0118_),
    .A2(_0122_));
 sg13g2_buf_1 _0674_ (.A(_0107_),
    .X(_0127_));
 sg13g2_nor2b_1 _0675_ (.A(net28),
    .B_N(_0002_),
    .Y(_0128_));
 sg13g2_buf_8 _0676_ (.A(net35),
    .X(_0129_));
 sg13g2_nor2b_1 _0677_ (.A(net27),
    .B_N(net29),
    .Y(_0130_));
 sg13g2_a22oi_1 _0678_ (.Y(_0131_),
    .B1(_0128_),
    .B2(_0130_),
    .A2(_0117_),
    .A1(_0004_));
 sg13g2_nor2b_1 _0679_ (.A(net34),
    .B_N(net30),
    .Y(_0132_));
 sg13g2_nor2b_1 _0680_ (.A(net29),
    .B_N(net27),
    .Y(_0133_));
 sg13g2_o21ai_1 _0681_ (.B1(_0133_),
    .Y(_0134_),
    .A1(_0132_),
    .A2(_0128_));
 sg13g2_a21oi_1 _0682_ (.A1(_0131_),
    .A2(_0134_),
    .Y(_0135_),
    .B1(_0006_));
 sg13g2_nand3b_1 _0683_ (.B(_0126_),
    .C(_0135_),
    .Y(_0136_),
    .A_N(_0125_));
 sg13g2_nand2b_1 _0684_ (.Y(_0137_),
    .B(_0127_),
    .A_N(net34));
 sg13g2_a21oi_1 _0685_ (.A1(_0115_),
    .A2(_0129_),
    .Y(_0138_),
    .B1(_0137_));
 sg13g2_nor2b_2 _0686_ (.A(_0107_),
    .B_N(_0111_),
    .Y(_0139_));
 sg13g2_or2_1 _0687_ (.X(_0140_),
    .B(_0104_),
    .A(_0106_));
 sg13g2_xnor2_1 _0688_ (.Y(_0141_),
    .A(_0139_),
    .B(_0140_));
 sg13g2_nor2_2 _0689_ (.A(_0138_),
    .B(_0141_),
    .Y(_0142_));
 sg13g2_xnor2_1 _0690_ (.Y(_0143_),
    .A(_0003_),
    .B(_0142_));
 sg13g2_a221oi_1 _0691_ (.B2(_0136_),
    .C1(_0143_),
    .B1(_0123_),
    .A1(_0103_),
    .Y(_0144_),
    .A2(_0114_));
 sg13g2_nand2_1 _0692_ (.Y(_0145_),
    .A(_0102_),
    .B(_0113_));
 sg13g2_nor2b_1 _0693_ (.A(_0142_),
    .B_N(\pulse_gen_inst.period_counter[10] ),
    .Y(_0146_));
 sg13g2_o21ai_1 _0694_ (.B1(_0146_),
    .Y(_0147_),
    .A1(_0102_),
    .A2(_0113_));
 sg13g2_nand3b_1 _0695_ (.B(_0145_),
    .C(_0147_),
    .Y(_0148_),
    .A_N(_0144_));
 sg13g2_buf_2 _0696_ (.A(_0148_),
    .X(_0149_));
 sg13g2_nor4_1 _0697_ (.A(\pulse_gen_inst.period_counter[31] ),
    .B(\pulse_gen_inst.period_counter[18] ),
    .C(\pulse_gen_inst.period_counter[17] ),
    .D(\pulse_gen_inst.period_counter[16] ),
    .Y(_0150_));
 sg13g2_nor4_1 _0698_ (.A(\pulse_gen_inst.period_counter[15] ),
    .B(\pulse_gen_inst.period_counter[14] ),
    .C(\pulse_gen_inst.period_counter[13] ),
    .D(\pulse_gen_inst.period_counter[12] ),
    .Y(_0151_));
 sg13g2_nor4_1 _0699_ (.A(\pulse_gen_inst.period_counter[30] ),
    .B(\pulse_gen_inst.period_counter[21] ),
    .C(\pulse_gen_inst.period_counter[20] ),
    .D(\pulse_gen_inst.period_counter[19] ),
    .Y(_0152_));
 sg13g2_nand3_1 _0700_ (.B(_0151_),
    .C(_0152_),
    .A(_0150_),
    .Y(_0153_));
 sg13g2_nor4_1 _0701_ (.A(\pulse_gen_inst.period_counter[29] ),
    .B(\pulse_gen_inst.period_counter[28] ),
    .C(\pulse_gen_inst.period_counter[27] ),
    .D(\pulse_gen_inst.period_counter[22] ),
    .Y(_0154_));
 sg13g2_nor4_1 _0702_ (.A(\pulse_gen_inst.period_counter[26] ),
    .B(\pulse_gen_inst.period_counter[25] ),
    .C(\pulse_gen_inst.period_counter[24] ),
    .D(\pulse_gen_inst.period_counter[23] ),
    .Y(_0155_));
 sg13g2_nand2_1 _0703_ (.Y(_0156_),
    .A(_0154_),
    .B(_0155_));
 sg13g2_nor2_1 _0704_ (.A(_0153_),
    .B(_0156_),
    .Y(_0157_));
 sg13g2_nor2b_1 _0705_ (.A(_0125_),
    .B_N(_0126_),
    .Y(_0158_));
 sg13g2_xor2_1 _0706_ (.B(_0142_),
    .A(_0003_),
    .X(_0159_));
 sg13g2_nand2_1 _0707_ (.Y(_0160_),
    .A(_0131_),
    .B(_0134_));
 sg13g2_xnor2_1 _0708_ (.Y(_0161_),
    .A(_0006_),
    .B(_0160_));
 sg13g2_nand2b_1 _0709_ (.Y(_0162_),
    .B(_0103_),
    .A_N(_0113_));
 sg13g2_and3_1 _0710_ (.X(_0163_),
    .A(_0145_),
    .B(_0151_),
    .C(_0162_));
 sg13g2_nand4_1 _0711_ (.B(_0159_),
    .C(_0161_),
    .A(_0158_),
    .Y(_0164_),
    .D(_0163_));
 sg13g2_nor2_2 _0712_ (.A(\reg_sequence_select[2] ),
    .B(_0107_),
    .Y(_0165_));
 sg13g2_xor2_1 _0713_ (.B(_0107_),
    .A(net34),
    .X(_0166_));
 sg13g2_and2_1 _0714_ (.A(net35),
    .B(_0111_),
    .X(_0167_));
 sg13g2_a221oi_1 _0715_ (.B2(_0115_),
    .C1(_0167_),
    .B1(_0166_),
    .A1(_0004_),
    .Y(_0168_),
    .A2(_0165_));
 sg13g2_and2_1 _0716_ (.A(_0009_),
    .B(_0168_),
    .X(_0169_));
 sg13g2_inv_1 _0717_ (.Y(_0170_),
    .A(_0010_));
 sg13g2_inv_2 _0718_ (.Y(_0171_),
    .A(_0107_));
 sg13g2_inv_1 _0719_ (.Y(_0172_),
    .A(_0011_));
 sg13g2_nor2b_1 _0720_ (.A(_0002_),
    .B_N(net30),
    .Y(_0173_));
 sg13g2_a22oi_1 _0721_ (.Y(_0174_),
    .B1(_0140_),
    .B2(_0173_),
    .A2(_0172_),
    .A1(_0171_));
 sg13g2_buf_1 _0722_ (.A(net29),
    .X(_0175_));
 sg13g2_inv_2 _0723_ (.Y(_0176_),
    .A(net34));
 sg13g2_a21oi_1 _0724_ (.A1(_0175_),
    .A2(net28),
    .Y(_0177_),
    .B1(_0176_));
 sg13g2_nand2b_1 _0725_ (.Y(_0178_),
    .B(net29),
    .A_N(net28));
 sg13g2_a21oi_1 _0726_ (.A1(_0176_),
    .A2(_0178_),
    .Y(_0179_),
    .B1(net27));
 sg13g2_nor4_1 _0727_ (.A(_0170_),
    .B(_0174_),
    .C(_0177_),
    .D(_0179_),
    .Y(_0180_));
 sg13g2_buf_2 _0728_ (.A(\pulse_gen_inst.period_counter[3] ),
    .X(_0181_));
 sg13g2_nor3_1 _0729_ (.A(_0181_),
    .B(_0177_),
    .C(_0179_),
    .Y(_0182_));
 sg13g2_nor3_1 _0730_ (.A(_0181_),
    .B(_0170_),
    .C(_0174_),
    .Y(_0183_));
 sg13g2_nor4_1 _0731_ (.A(_0169_),
    .B(_0180_),
    .C(_0182_),
    .D(_0183_),
    .Y(_0184_));
 sg13g2_nor2_1 _0732_ (.A(_0009_),
    .B(_0168_),
    .Y(_0185_));
 sg13g2_buf_1 _0733_ (.A(net27),
    .X(_0186_));
 sg13g2_buf_1 _0734_ (.A(net34),
    .X(_0187_));
 sg13g2_nand2_1 _0735_ (.Y(_0188_),
    .A(_0187_),
    .B(net28));
 sg13g2_nand3b_1 _0736_ (.B(net30),
    .C(net29),
    .Y(_0189_),
    .A_N(net35));
 sg13g2_nand2b_1 _0737_ (.Y(_0190_),
    .B(_0189_),
    .A_N(_0109_));
 sg13g2_buf_1 _0738_ (.A(net26),
    .X(_0191_));
 sg13g2_a22oi_1 _0739_ (.Y(_0192_),
    .B1(_0190_),
    .B2(net23),
    .A2(_0188_),
    .A1(net24));
 sg13g2_xor2_1 _0740_ (.B(_0192_),
    .A(_0008_),
    .X(_0193_));
 sg13g2_o21ai_1 _0741_ (.B1(_0193_),
    .Y(_0194_),
    .A1(_0184_),
    .A2(_0185_));
 sg13g2_buf_1 _0742_ (.A(\pulse_gen_inst.period_counter[7] ),
    .X(_0195_));
 sg13g2_nand2_1 _0743_ (.Y(_0196_),
    .A(net27),
    .B(net28));
 sg13g2_buf_1 _0744_ (.A(\pulse_gen_inst.period_counter[6] ),
    .X(_0197_));
 sg13g2_nor2_1 _0745_ (.A(net29),
    .B(_0197_),
    .Y(_0198_));
 sg13g2_nor2b_1 _0746_ (.A(net30),
    .B_N(net35),
    .Y(_0199_));
 sg13g2_and2_1 _0747_ (.A(net30),
    .B(_0197_),
    .X(_0200_));
 sg13g2_nor2_1 _0748_ (.A(net29),
    .B(_0187_),
    .Y(_0201_));
 sg13g2_o21ai_1 _0749_ (.B1(_0201_),
    .Y(_0202_),
    .A1(_0199_),
    .A2(_0200_));
 sg13g2_o21ai_1 _0750_ (.B1(_0202_),
    .Y(_0203_),
    .A1(_0196_),
    .A2(_0198_));
 sg13g2_a21oi_1 _0751_ (.A1(_0171_),
    .A2(_0197_),
    .Y(_0204_),
    .B1(net26));
 sg13g2_nand2_1 _0752_ (.Y(_0205_),
    .A(net26),
    .B(_0197_));
 sg13g2_o21ai_1 _0753_ (.B1(_0205_),
    .Y(_0206_),
    .A1(net24),
    .A2(_0204_));
 sg13g2_and2_1 _0754_ (.A(net25),
    .B(net33),
    .X(_0207_));
 sg13g2_nand3b_1 _0755_ (.B(net28),
    .C(net27),
    .Y(_0208_),
    .A_N(net26));
 sg13g2_nand2b_1 _0756_ (.Y(_0209_),
    .B(net26),
    .A_N(net27));
 sg13g2_nand2_1 _0757_ (.Y(_0210_),
    .A(net25),
    .B(_0197_));
 sg13g2_a21oi_1 _0758_ (.A1(_0208_),
    .A2(_0209_),
    .Y(_0211_),
    .B1(_0210_));
 sg13g2_a221oi_1 _0759_ (.B2(_0207_),
    .C1(_0211_),
    .B1(_0206_),
    .A1(net33),
    .Y(_0212_),
    .A2(_0203_));
 sg13g2_inv_1 _0760_ (.Y(_0213_),
    .A(\pulse_gen_inst.period_counter[5] ));
 sg13g2_or2_1 _0761_ (.X(_0214_),
    .B(_0192_),
    .A(_0213_));
 sg13g2_and3_1 _0762_ (.X(_0215_),
    .A(_0157_),
    .B(_0212_),
    .C(_0214_));
 sg13g2_buf_1 _0763_ (.A(_0175_),
    .X(_0216_));
 sg13g2_buf_2 _0764_ (.A(_0007_),
    .X(_0217_));
 sg13g2_nor2b_1 _0765_ (.A(net33),
    .B_N(_0217_),
    .Y(_0218_));
 sg13g2_xor2_1 _0766_ (.B(_0217_),
    .A(_0108_),
    .X(_0219_));
 sg13g2_and2_1 _0767_ (.A(net33),
    .B(_0219_),
    .X(_0220_));
 sg13g2_nor2_1 _0768_ (.A(\pulse_gen_inst.period_counter[7] ),
    .B(_0217_),
    .Y(_0221_));
 sg13g2_and2_1 _0769_ (.A(\pulse_gen_inst.period_counter[7] ),
    .B(_0217_),
    .X(_0222_));
 sg13g2_mux2_1 _0770_ (.A0(_0221_),
    .A1(_0222_),
    .S(_0171_),
    .X(_0223_));
 sg13g2_nor2b_1 _0771_ (.A(_0217_),
    .B_N(\pulse_gen_inst.period_counter[7] ),
    .Y(_0224_));
 sg13g2_mux2_1 _0772_ (.A0(_0218_),
    .A1(_0224_),
    .S(_0171_),
    .X(_0225_));
 sg13g2_mux4_1 _0773_ (.S0(_0176_),
    .A0(_0218_),
    .A1(_0220_),
    .A2(_0223_),
    .A3(_0225_),
    .S1(_0186_),
    .X(_0226_));
 sg13g2_nand2_1 _0774_ (.Y(_0227_),
    .A(net19),
    .B(_0226_));
 sg13g2_buf_1 _0775_ (.A(_0127_),
    .X(_0228_));
 sg13g2_nand4_1 _0776_ (.B(_0228_),
    .C(net33),
    .A(_0176_),
    .Y(_0229_),
    .D(_0217_));
 sg13g2_and3_1 _0777_ (.X(_0230_),
    .A(net30),
    .B(_0195_),
    .C(_0217_));
 sg13g2_a21o_1 _0778_ (.A2(_0165_),
    .A1(_0221_),
    .B1(_0230_),
    .X(_0231_));
 sg13g2_nand2b_1 _0779_ (.Y(_0232_),
    .B(net26),
    .A_N(net28));
 sg13g2_o21ai_1 _0780_ (.B1(_0232_),
    .Y(_0233_),
    .A1(net27),
    .A2(_0132_));
 sg13g2_a22oi_1 _0781_ (.Y(_0234_),
    .B1(_0233_),
    .B2(_0224_),
    .A2(_0231_),
    .A1(_0186_));
 sg13g2_a21o_1 _0782_ (.A2(_0234_),
    .A1(_0229_),
    .B1(net19),
    .X(_0235_));
 sg13g2_and4_1 _0783_ (.A(_0157_),
    .B(_0212_),
    .C(_0227_),
    .D(_0235_),
    .X(_0236_));
 sg13g2_a221oi_1 _0784_ (.B2(_0215_),
    .C1(_0236_),
    .B1(_0194_),
    .A1(_0157_),
    .Y(_0237_),
    .A2(_0164_));
 sg13g2_buf_2 _0785_ (.A(_0237_),
    .X(_0238_));
 sg13g2_or2_1 _0786_ (.X(_0239_),
    .B(_0238_),
    .A(_0149_));
 sg13g2_buf_1 _0787_ (.A(_0239_),
    .X(_0240_));
 sg13g2_buf_1 _0788_ (.A(_0240_),
    .X(_0241_));
 sg13g2_buf_1 _0789_ (.A(\pulse_gen_inst.count_counter[2] ),
    .X(_0242_));
 sg13g2_nor2_1 _0790_ (.A(\pulse_gen_inst.count_counter[6] ),
    .B(\pulse_gen_inst.count_counter[5] ),
    .Y(_0243_));
 sg13g2_nor4_1 _0791_ (.A(\pulse_gen_inst.count_counter[9] ),
    .B(\pulse_gen_inst.count_counter[8] ),
    .C(\pulse_gen_inst.count_counter[7] ),
    .D(\pulse_gen_inst.count_counter[4] ),
    .Y(_0244_));
 sg13g2_nor4_1 _0792_ (.A(\pulse_gen_inst.count_counter[14] ),
    .B(\pulse_gen_inst.count_counter[13] ),
    .C(\pulse_gen_inst.count_counter[12] ),
    .D(\pulse_gen_inst.count_counter[11] ),
    .Y(_0245_));
 sg13g2_nor2_1 _0793_ (.A(\pulse_gen_inst.count_counter[15] ),
    .B(\pulse_gen_inst.count_counter[10] ),
    .Y(_0246_));
 sg13g2_nand4_1 _0794_ (.B(_0244_),
    .C(_0245_),
    .A(_0243_),
    .Y(_0247_),
    .D(_0246_));
 sg13g2_nor3_1 _0795_ (.A(\pulse_gen_inst.count_counter[3] ),
    .B(_0242_),
    .C(_0247_),
    .Y(_0248_));
 sg13g2_nand3b_1 _0796_ (.B(net12),
    .C(_0248_),
    .Y(_0249_),
    .A_N(\pulse_gen_inst.count_counter[1] ));
 sg13g2_or4_1 _0797_ (.A(\pulse_gen_inst.count_counter[3] ),
    .B(_0242_),
    .C(\pulse_gen_inst.count_counter[0] ),
    .D(\pulse_gen_inst.count_counter[1] ),
    .X(_0250_));
 sg13g2_nor2_1 _0798_ (.A(_0250_),
    .B(_0247_),
    .Y(_0251_));
 sg13g2_a21o_1 _0799_ (.A2(_0249_),
    .A1(net31),
    .B1(_0251_),
    .X(_0000_));
 sg13g2_inv_1 _0800_ (.Y(_0252_),
    .A(net36));
 sg13g2_buf_1 _0801_ (.A(_0252_),
    .X(_0253_));
 sg13g2_buf_1 _0802_ (.A(net21),
    .X(_0254_));
 sg13g2_buf_1 _0803_ (.A(_0017_),
    .X(_0255_));
 sg13g2_inv_1 _0804_ (.Y(_0256_),
    .A(net32));
 sg13g2_nand2_1 _0805_ (.Y(_0257_),
    .A(_0256_),
    .B(_0018_));
 sg13g2_inv_1 _0806_ (.Y(_0258_),
    .A(\pulse_gen_inst.count_counter[0] ));
 sg13g2_or2_1 _0807_ (.X(_0259_),
    .B(_0247_),
    .A(_0250_));
 sg13g2_buf_2 _0808_ (.A(_0259_),
    .X(_0260_));
 sg13g2_o21ai_1 _0809_ (.B1(_0260_),
    .Y(_0261_),
    .A1(_0149_),
    .A2(_0238_));
 sg13g2_mux2_1 _0810_ (.A0(_0257_),
    .A1(_0258_),
    .S(_0261_),
    .X(_0262_));
 sg13g2_a21oi_2 _0811_ (.B1(net36),
    .Y(_0263_),
    .A2(_0260_),
    .A1(net32));
 sg13g2_buf_1 _0812_ (.A(_0263_),
    .X(_0264_));
 sg13g2_buf_1 _0813_ (.A(_0129_),
    .X(_0265_));
 sg13g2_nand2_1 _0814_ (.Y(_0266_),
    .A(net19),
    .B(net20));
 sg13g2_or2_1 _0815_ (.X(_0267_),
    .B(_0004_),
    .A(net22));
 sg13g2_nand2_1 _0816_ (.Y(_0268_),
    .A(net23),
    .B(_0267_));
 sg13g2_a21oi_1 _0817_ (.A1(_0171_),
    .A2(_0004_),
    .Y(_0269_),
    .B1(_0266_));
 sg13g2_a22oi_1 _0818_ (.Y(_0270_),
    .B1(_0269_),
    .B2(net23),
    .A2(_0268_),
    .A1(_0266_));
 sg13g2_a22oi_1 _0819_ (.Y(_0271_),
    .B1(net16),
    .B2(_0270_),
    .A2(net32),
    .A1(\pulse_gen_inst.count_counter[0] ));
 sg13g2_o21ai_1 _0820_ (.B1(_0271_),
    .Y(_0019_),
    .A1(net18),
    .A2(_0262_));
 sg13g2_buf_1 _0821_ (.A(net21),
    .X(_0272_));
 sg13g2_nand2_2 _0822_ (.Y(_0273_),
    .A(net32),
    .B(_0260_));
 sg13g2_buf_1 _0823_ (.A(_0261_),
    .X(_0274_));
 sg13g2_inv_1 _0824_ (.Y(_0275_),
    .A(_0250_));
 sg13g2_nand4_1 _0825_ (.B(_0243_),
    .C(_0244_),
    .A(_0275_),
    .Y(_0276_),
    .D(_0273_));
 sg13g2_buf_1 _0826_ (.A(_0276_),
    .X(_0277_));
 sg13g2_a21o_1 _0827_ (.A2(net15),
    .A1(net31),
    .B1(_0277_),
    .X(_0278_));
 sg13g2_inv_1 _0828_ (.Y(_0279_),
    .A(\pulse_gen_inst.count_counter[10] ));
 sg13g2_nor3_1 _0829_ (.A(_0279_),
    .B(net15),
    .C(_0277_),
    .Y(_0280_));
 sg13g2_a221oi_1 _0830_ (.B2(_0279_),
    .C1(_0280_),
    .B1(_0278_),
    .A1(_0272_),
    .Y(_0020_),
    .A2(_0273_));
 sg13g2_nor2b_1 _0831_ (.A(net16),
    .B_N(\pulse_gen_inst.count_counter[11] ),
    .Y(_0281_));
 sg13g2_nor2_1 _0832_ (.A(\pulse_gen_inst.count_counter[11] ),
    .B(_0263_),
    .Y(_0282_));
 sg13g2_nor2_1 _0833_ (.A(\pulse_gen_inst.count_counter[10] ),
    .B(_0277_),
    .Y(_0283_));
 sg13g2_inv_1 _0834_ (.Y(_0284_),
    .A(_0283_));
 sg13g2_a21oi_1 _0835_ (.A1(net36),
    .A2(_0261_),
    .Y(_0285_),
    .B1(_0284_));
 sg13g2_mux2_1 _0836_ (.A0(_0281_),
    .A1(_0282_),
    .S(_0285_),
    .X(_0021_));
 sg13g2_nor4_1 _0837_ (.A(\pulse_gen_inst.count_counter[11] ),
    .B(\pulse_gen_inst.count_counter[10] ),
    .C(_0251_),
    .D(_0277_),
    .Y(_0286_));
 sg13g2_o21ai_1 _0838_ (.B1(_0286_),
    .Y(_0287_),
    .A1(_0149_),
    .A2(_0238_));
 sg13g2_or4_1 _0839_ (.A(net36),
    .B(\pulse_gen_inst.count_counter[11] ),
    .C(\pulse_gen_inst.count_counter[10] ),
    .D(_0277_),
    .X(_0288_));
 sg13g2_nand3_1 _0840_ (.B(_0287_),
    .C(_0288_),
    .A(\pulse_gen_inst.count_counter[12] ),
    .Y(_0289_));
 sg13g2_a21o_1 _0841_ (.A2(_0288_),
    .A1(_0287_),
    .B1(\pulse_gen_inst.count_counter[12] ),
    .X(_0290_));
 sg13g2_a21oi_1 _0842_ (.A1(_0289_),
    .A2(_0290_),
    .Y(_0022_),
    .B1(net16));
 sg13g2_nor2_1 _0843_ (.A(\pulse_gen_inst.count_counter[13] ),
    .B(_0263_),
    .Y(_0291_));
 sg13g2_nor2b_1 _0844_ (.A(_0263_),
    .B_N(\pulse_gen_inst.count_counter[13] ),
    .Y(_0292_));
 sg13g2_mux2_1 _0845_ (.A0(_0291_),
    .A1(_0292_),
    .S(_0290_),
    .X(_0023_));
 sg13g2_nor2b_1 _0846_ (.A(_0263_),
    .B_N(\pulse_gen_inst.count_counter[14] ),
    .Y(_0293_));
 sg13g2_nor2_1 _0847_ (.A(\pulse_gen_inst.count_counter[14] ),
    .B(_0263_),
    .Y(_0294_));
 sg13g2_nor3_1 _0848_ (.A(\pulse_gen_inst.count_counter[13] ),
    .B(\pulse_gen_inst.count_counter[12] ),
    .C(\pulse_gen_inst.count_counter[11] ),
    .Y(_0295_));
 sg13g2_nand2_1 _0849_ (.Y(_0296_),
    .A(_0295_),
    .B(_0283_));
 sg13g2_a21oi_1 _0850_ (.A1(net36),
    .A2(_0261_),
    .Y(_0297_),
    .B1(_0296_));
 sg13g2_mux2_1 _0851_ (.A0(_0293_),
    .A1(_0294_),
    .S(_0297_),
    .X(_0024_));
 sg13g2_o21ai_1 _0852_ (.B1(\pulse_gen_inst.count_counter[15] ),
    .Y(_0298_),
    .A1(net31),
    .A2(net32));
 sg13g2_a21oi_1 _0853_ (.A1(_0245_),
    .A2(_0285_),
    .Y(_0025_),
    .B1(_0298_));
 sg13g2_buf_1 _0854_ (.A(_0240_),
    .X(_0299_));
 sg13g2_nor3_1 _0855_ (.A(\pulse_gen_inst.count_counter[0] ),
    .B(\pulse_gen_inst.count_counter[1] ),
    .C(_0248_),
    .Y(_0300_));
 sg13g2_and2_1 _0856_ (.A(_0256_),
    .B(_0300_),
    .X(_0301_));
 sg13g2_o21ai_1 _0857_ (.B1(_0258_),
    .Y(_0302_),
    .A1(_0149_),
    .A2(_0238_));
 sg13g2_a22oi_1 _0858_ (.Y(_0303_),
    .B1(_0302_),
    .B2(\pulse_gen_inst.count_counter[1] ),
    .A2(_0301_),
    .A1(net11));
 sg13g2_nor2_1 _0859_ (.A(net28),
    .B(_0004_),
    .Y(_0304_));
 sg13g2_xnor2_1 _0860_ (.Y(_0305_),
    .A(_0116_),
    .B(_0110_));
 sg13g2_nor2_1 _0861_ (.A(_0011_),
    .B(_0188_),
    .Y(_0306_));
 sg13g2_a221oi_1 _0862_ (.B2(_0176_),
    .C1(_0306_),
    .B1(_0305_),
    .A1(_0116_),
    .Y(_0307_),
    .A2(_0304_));
 sg13g2_a22oi_1 _0863_ (.Y(_0308_),
    .B1(net16),
    .B2(_0307_),
    .A2(net32),
    .A1(\pulse_gen_inst.count_counter[1] ));
 sg13g2_o21ai_1 _0864_ (.B1(_0308_),
    .Y(_0026_),
    .A1(_0254_),
    .A2(_0303_));
 sg13g2_and4_1 _0865_ (.A(net36),
    .B(_0242_),
    .C(_0240_),
    .D(_0301_),
    .X(_0309_));
 sg13g2_nand2b_1 _0866_ (.Y(_0310_),
    .B(_0100_),
    .A_N(_0242_));
 sg13g2_a21oi_1 _0867_ (.A1(net11),
    .A2(_0300_),
    .Y(_0311_),
    .B1(_0310_));
 sg13g2_inv_1 _0868_ (.Y(_0312_),
    .A(_0004_));
 sg13g2_a22oi_1 _0869_ (.Y(_0313_),
    .B1(_0139_),
    .B2(_0216_),
    .A2(_0312_),
    .A1(net22));
 sg13g2_nor3_1 _0870_ (.A(net20),
    .B(_0165_),
    .C(_0173_),
    .Y(_0314_));
 sg13g2_a21oi_1 _0871_ (.A1(net20),
    .A2(_0313_),
    .Y(_0315_),
    .B1(_0314_));
 sg13g2_nand2_1 _0872_ (.Y(_0316_),
    .A(_0263_),
    .B(_0315_));
 sg13g2_o21ai_1 _0873_ (.B1(_0316_),
    .Y(_0317_),
    .A1(_0242_),
    .A2(_0273_));
 sg13g2_nor3_1 _0874_ (.A(_0309_),
    .B(_0311_),
    .C(_0317_),
    .Y(_0027_));
 sg13g2_a21oi_1 _0875_ (.A1(_0299_),
    .A2(_0301_),
    .Y(_0318_),
    .B1(\pulse_gen_inst.count_counter[3] ));
 sg13g2_inv_1 _0876_ (.Y(_0319_),
    .A(\pulse_gen_inst.count_counter[3] ));
 sg13g2_nor4_1 _0877_ (.A(_0319_),
    .B(_0242_),
    .C(\pulse_gen_inst.count_counter[0] ),
    .D(\pulse_gen_inst.count_counter[1] ),
    .Y(_0320_));
 sg13g2_o21ai_1 _0878_ (.B1(_0320_),
    .Y(_0321_),
    .A1(_0149_),
    .A2(_0238_));
 sg13g2_a21oi_1 _0879_ (.A1(_0319_),
    .A2(_0242_),
    .Y(_0322_),
    .B1(net21));
 sg13g2_nand2_1 _0880_ (.Y(_0323_),
    .A(_0321_),
    .B(_0322_));
 sg13g2_nand2_1 _0881_ (.Y(_0324_),
    .A(_0121_),
    .B(_0139_));
 sg13g2_o21ai_1 _0882_ (.B1(_0324_),
    .Y(_0325_),
    .A1(_0121_),
    .A2(_0166_));
 sg13g2_a21oi_1 _0883_ (.A1(_0216_),
    .A2(_0139_),
    .Y(_0326_),
    .B1(_0110_));
 sg13g2_nor2_1 _0884_ (.A(_0265_),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_a221oi_1 _0885_ (.B2(_0265_),
    .C1(_0327_),
    .B1(_0325_),
    .A1(_0121_),
    .Y(_0328_),
    .A2(_0132_));
 sg13g2_a22oi_1 _0886_ (.Y(_0329_),
    .B1(_0264_),
    .B2(_0328_),
    .A2(_0255_),
    .A1(\pulse_gen_inst.count_counter[3] ));
 sg13g2_o21ai_1 _0887_ (.B1(_0329_),
    .Y(_0028_),
    .A1(_0318_),
    .A2(_0323_));
 sg13g2_inv_1 _0888_ (.Y(_0330_),
    .A(\pulse_gen_inst.count_counter[4] ));
 sg13g2_nor2_1 _0889_ (.A(_0330_),
    .B(net32),
    .Y(_0331_));
 sg13g2_and2_1 _0890_ (.A(_0275_),
    .B(_0247_),
    .X(_0332_));
 sg13g2_o21ai_1 _0891_ (.B1(_0332_),
    .Y(_0333_),
    .A1(_0149_),
    .A2(_0238_));
 sg13g2_mux2_1 _0892_ (.A0(_0331_),
    .A1(_0330_),
    .S(_0333_),
    .X(_0334_));
 sg13g2_a22oi_1 _0893_ (.Y(_0335_),
    .B1(_0139_),
    .B2(_0116_),
    .A2(_0105_),
    .A1(_0228_));
 sg13g2_nand2b_1 _0894_ (.Y(_0336_),
    .B(net19),
    .A_N(_0335_));
 sg13g2_nor2_1 _0895_ (.A(\pulse_gen_inst.count_counter[4] ),
    .B(_0273_),
    .Y(_0337_));
 sg13g2_a221oi_1 _0896_ (.B2(_0264_),
    .C1(_0337_),
    .B1(_0336_),
    .A1(net31),
    .Y(_0029_),
    .A2(_0334_));
 sg13g2_nor2_1 _0897_ (.A(\pulse_gen_inst.count_counter[4] ),
    .B(_0250_),
    .Y(_0338_));
 sg13g2_nand2_1 _0898_ (.Y(_0339_),
    .A(_0273_),
    .B(_0338_));
 sg13g2_o21ai_1 _0899_ (.B1(\pulse_gen_inst.count_counter[5] ),
    .Y(_0340_),
    .A1(_0274_),
    .A2(_0339_));
 sg13g2_or3_1 _0900_ (.A(\pulse_gen_inst.count_counter[5] ),
    .B(net15),
    .C(_0339_),
    .X(_0341_));
 sg13g2_a21oi_1 _0901_ (.A1(_0340_),
    .A2(_0341_),
    .Y(_0030_),
    .B1(net16));
 sg13g2_inv_1 _0902_ (.Y(_0342_),
    .A(\pulse_gen_inst.count_counter[6] ));
 sg13g2_nor4_1 _0903_ (.A(_0342_),
    .B(\pulse_gen_inst.count_counter[5] ),
    .C(net15),
    .D(_0339_),
    .Y(_0343_));
 sg13g2_and2_1 _0904_ (.A(_0342_),
    .B(net15),
    .X(_0344_));
 sg13g2_a21oi_1 _0905_ (.A1(_0273_),
    .A2(_0338_),
    .Y(_0345_),
    .B1(\pulse_gen_inst.count_counter[6] ));
 sg13g2_a22oi_1 _0906_ (.Y(_0346_),
    .B1(_0256_),
    .B2(net21),
    .A2(\pulse_gen_inst.count_counter[5] ),
    .A1(_0342_));
 sg13g2_o21ai_1 _0907_ (.B1(_0346_),
    .Y(_0347_),
    .A1(_0101_),
    .A2(\pulse_gen_inst.count_counter[6] ));
 sg13g2_nor4_1 _0908_ (.A(_0343_),
    .B(_0344_),
    .C(_0345_),
    .D(_0347_),
    .Y(_0031_));
 sg13g2_nand2_1 _0909_ (.Y(_0348_),
    .A(_0243_),
    .B(_0338_));
 sg13g2_a21oi_1 _0910_ (.A1(net32),
    .A2(_0247_),
    .Y(_0349_),
    .B1(_0348_));
 sg13g2_nand2_1 _0911_ (.Y(_0350_),
    .A(\pulse_gen_inst.count_counter[7] ),
    .B(_0349_));
 sg13g2_nor2_1 _0912_ (.A(_0274_),
    .B(_0350_),
    .Y(_0351_));
 sg13g2_nor2_1 _0913_ (.A(net21),
    .B(\pulse_gen_inst.count_counter[7] ),
    .Y(_0352_));
 sg13g2_and2_1 _0914_ (.A(net15),
    .B(_0352_),
    .X(_0353_));
 sg13g2_nor2_1 _0915_ (.A(\pulse_gen_inst.count_counter[7] ),
    .B(_0349_),
    .Y(_0354_));
 sg13g2_nor4_1 _0916_ (.A(net16),
    .B(_0351_),
    .C(_0353_),
    .D(_0354_),
    .Y(_0032_));
 sg13g2_inv_1 _0917_ (.Y(_0355_),
    .A(\pulse_gen_inst.count_counter[8] ));
 sg13g2_nor2b_1 _0918_ (.A(\pulse_gen_inst.count_counter[7] ),
    .B_N(_0349_),
    .Y(_0356_));
 sg13g2_and2_1 _0919_ (.A(_0260_),
    .B(_0356_),
    .X(_0357_));
 sg13g2_o21ai_1 _0920_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_0253_),
    .A2(net12));
 sg13g2_and2_1 _0921_ (.A(\pulse_gen_inst.count_counter[8] ),
    .B(_0356_),
    .X(_0359_));
 sg13g2_a221oi_1 _0922_ (.B2(_0299_),
    .C1(net16),
    .B1(_0359_),
    .A1(_0355_),
    .Y(_0033_),
    .A2(_0358_));
 sg13g2_or2_1 _0923_ (.X(_0360_),
    .B(_0277_),
    .A(net15));
 sg13g2_nand2_1 _0924_ (.Y(_0361_),
    .A(_0355_),
    .B(_0356_));
 sg13g2_o21ai_1 _0925_ (.B1(\pulse_gen_inst.count_counter[9] ),
    .Y(_0362_),
    .A1(net15),
    .A2(_0361_));
 sg13g2_a21oi_1 _0926_ (.A1(_0360_),
    .A2(_0362_),
    .Y(_0034_),
    .B1(net16));
 sg13g2_inv_1 _0927_ (.Y(_0363_),
    .A(\pulse_gen_inst.period_counter[0] ));
 sg13g2_nor2_2 _0928_ (.A(_0149_),
    .B(_0238_),
    .Y(_0364_));
 sg13g2_nand3_1 _0929_ (.B(_0363_),
    .C(_0364_),
    .A(net31),
    .Y(_0365_));
 sg13g2_o21ai_1 _0930_ (.B1(_0365_),
    .Y(_0035_),
    .A1(net31),
    .A2(_0363_));
 sg13g2_and3_1 _0931_ (.X(_0366_),
    .A(\pulse_gen_inst.period_counter[0] ),
    .B(\pulse_gen_inst.period_counter[1] ),
    .C(\pulse_gen_inst.period_counter[2] ));
 sg13g2_buf_8 _0932_ (.A(_0366_),
    .X(_0367_));
 sg13g2_and2_1 _0933_ (.A(_0181_),
    .B(\pulse_gen_inst.period_counter[4] ),
    .X(_0368_));
 sg13g2_and4_1 _0934_ (.A(_0197_),
    .B(\pulse_gen_inst.period_counter[5] ),
    .C(_0367_),
    .D(_0368_),
    .X(_0369_));
 sg13g2_buf_2 _0935_ (.A(_0369_),
    .X(_0370_));
 sg13g2_and2_1 _0936_ (.A(net33),
    .B(_0370_),
    .X(_0371_));
 sg13g2_buf_1 _0937_ (.A(_0371_),
    .X(_0372_));
 sg13g2_nand3_1 _0938_ (.B(\pulse_gen_inst.period_counter[8] ),
    .C(_0372_),
    .A(\pulse_gen_inst.period_counter[9] ),
    .Y(_0373_));
 sg13g2_xnor2_1 _0939_ (.Y(_0374_),
    .A(_0003_),
    .B(_0373_));
 sg13g2_nor3_1 _0940_ (.A(net17),
    .B(net11),
    .C(_0374_),
    .Y(_0375_));
 sg13g2_a21o_1 _0941_ (.A2(net18),
    .A1(\pulse_gen_inst.period_counter[10] ),
    .B1(_0375_),
    .X(_0036_));
 sg13g2_nor2_2 _0942_ (.A(net21),
    .B(_0364_),
    .Y(_0376_));
 sg13g2_buf_1 _0943_ (.A(_0376_),
    .X(_0377_));
 sg13g2_nand2_1 _0944_ (.Y(_0378_),
    .A(\pulse_gen_inst.period_counter[8] ),
    .B(_0372_));
 sg13g2_nand3_1 _0945_ (.B(\pulse_gen_inst.period_counter[9] ),
    .C(net36),
    .A(\pulse_gen_inst.period_counter[10] ),
    .Y(_0379_));
 sg13g2_nor2_1 _0946_ (.A(_0378_),
    .B(_0379_),
    .Y(_0380_));
 sg13g2_xnor2_1 _0947_ (.Y(_0381_),
    .A(_0102_),
    .B(_0380_));
 sg13g2_nor2_1 _0948_ (.A(net10),
    .B(_0381_),
    .Y(_0037_));
 sg13g2_nand2_1 _0949_ (.Y(_0382_),
    .A(_0102_),
    .B(_0380_));
 sg13g2_xor2_1 _0950_ (.B(_0382_),
    .A(\pulse_gen_inst.period_counter[12] ),
    .X(_0383_));
 sg13g2_nor2_1 _0951_ (.A(net10),
    .B(_0383_),
    .Y(_0038_));
 sg13g2_nand3_1 _0952_ (.B(_0102_),
    .C(_0380_),
    .A(\pulse_gen_inst.period_counter[12] ),
    .Y(_0384_));
 sg13g2_xor2_1 _0953_ (.B(_0384_),
    .A(\pulse_gen_inst.period_counter[13] ),
    .X(_0385_));
 sg13g2_nor2_1 _0954_ (.A(net10),
    .B(_0385_),
    .Y(_0039_));
 sg13g2_nand4_1 _0955_ (.B(\pulse_gen_inst.period_counter[12] ),
    .C(_0102_),
    .A(\pulse_gen_inst.period_counter[13] ),
    .Y(_0386_),
    .D(\pulse_gen_inst.period_counter[8] ));
 sg13g2_nor2_1 _0956_ (.A(_0379_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_nand2_1 _0957_ (.Y(_0388_),
    .A(_0372_),
    .B(_0387_));
 sg13g2_xor2_1 _0958_ (.B(_0388_),
    .A(\pulse_gen_inst.period_counter[14] ),
    .X(_0389_));
 sg13g2_nor2_1 _0959_ (.A(_0377_),
    .B(_0389_),
    .Y(_0040_));
 sg13g2_and2_1 _0960_ (.A(\pulse_gen_inst.period_counter[14] ),
    .B(net33),
    .X(_0390_));
 sg13g2_nand3_1 _0961_ (.B(_0387_),
    .C(_0390_),
    .A(_0370_),
    .Y(_0391_));
 sg13g2_xor2_1 _0962_ (.B(_0391_),
    .A(\pulse_gen_inst.period_counter[15] ),
    .X(_0392_));
 sg13g2_nor2_1 _0963_ (.A(_0377_),
    .B(_0392_),
    .Y(_0041_));
 sg13g2_inv_1 _0964_ (.Y(_0393_),
    .A(\pulse_gen_inst.period_counter[16] ));
 sg13g2_nand4_1 _0965_ (.B(_0370_),
    .C(_0387_),
    .A(\pulse_gen_inst.period_counter[15] ),
    .Y(_0394_),
    .D(_0390_));
 sg13g2_xnor2_1 _0966_ (.Y(_0395_),
    .A(_0393_),
    .B(_0394_));
 sg13g2_nor2_1 _0967_ (.A(net10),
    .B(_0395_),
    .Y(_0042_));
 sg13g2_inv_1 _0968_ (.Y(_0396_),
    .A(\pulse_gen_inst.period_counter[17] ));
 sg13g2_or2_1 _0969_ (.X(_0397_),
    .B(_0394_),
    .A(_0393_));
 sg13g2_buf_1 _0970_ (.A(_0397_),
    .X(_0398_));
 sg13g2_xnor2_1 _0971_ (.Y(_0399_),
    .A(_0396_),
    .B(_0398_));
 sg13g2_nor2_1 _0972_ (.A(net10),
    .B(_0399_),
    .Y(_0043_));
 sg13g2_nor2_1 _0973_ (.A(_0396_),
    .B(_0398_),
    .Y(_0400_));
 sg13g2_xnor2_1 _0974_ (.Y(_0401_),
    .A(\pulse_gen_inst.period_counter[18] ),
    .B(_0400_));
 sg13g2_nor2_1 _0975_ (.A(net10),
    .B(_0401_),
    .Y(_0044_));
 sg13g2_nand2_1 _0976_ (.Y(_0402_),
    .A(\pulse_gen_inst.period_counter[18] ),
    .B(\pulse_gen_inst.period_counter[17] ));
 sg13g2_nor2_1 _0977_ (.A(_0398_),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_xnor2_1 _0978_ (.Y(_0404_),
    .A(\pulse_gen_inst.period_counter[19] ),
    .B(_0403_));
 sg13g2_nor2_1 _0979_ (.A(net10),
    .B(_0404_),
    .Y(_0045_));
 sg13g2_o21ai_1 _0980_ (.B1(net31),
    .Y(_0405_),
    .A1(\pulse_gen_inst.period_counter[0] ),
    .A2(net12));
 sg13g2_nor4_1 _0981_ (.A(net21),
    .B(_0363_),
    .C(\pulse_gen_inst.period_counter[1] ),
    .D(net12),
    .Y(_0406_));
 sg13g2_a21o_1 _0982_ (.A2(_0405_),
    .A1(\pulse_gen_inst.period_counter[1] ),
    .B1(_0406_),
    .X(_0046_));
 sg13g2_a21oi_1 _0983_ (.A1(\pulse_gen_inst.period_counter[19] ),
    .A2(_0403_),
    .Y(_0407_),
    .B1(\pulse_gen_inst.period_counter[20] ));
 sg13g2_nor2_1 _0984_ (.A(net10),
    .B(_0407_),
    .Y(_0047_));
 sg13g2_buf_1 _0985_ (.A(_0376_),
    .X(_0408_));
 sg13g2_and3_1 _0986_ (.X(_0409_),
    .A(\pulse_gen_inst.period_counter[20] ),
    .B(\pulse_gen_inst.period_counter[19] ),
    .C(_0403_));
 sg13g2_xnor2_1 _0987_ (.Y(_0410_),
    .A(\pulse_gen_inst.period_counter[21] ),
    .B(_0409_));
 sg13g2_nor2_1 _0988_ (.A(net9),
    .B(_0410_),
    .Y(_0048_));
 sg13g2_nand2_1 _0989_ (.Y(_0411_),
    .A(\pulse_gen_inst.period_counter[21] ),
    .B(_0409_));
 sg13g2_xor2_1 _0990_ (.B(_0411_),
    .A(\pulse_gen_inst.period_counter[22] ),
    .X(_0412_));
 sg13g2_nor2_1 _0991_ (.A(net9),
    .B(_0412_),
    .Y(_0049_));
 sg13g2_nand3_1 _0992_ (.B(\pulse_gen_inst.period_counter[21] ),
    .C(_0409_),
    .A(\pulse_gen_inst.period_counter[22] ),
    .Y(_0413_));
 sg13g2_xor2_1 _0993_ (.B(_0413_),
    .A(\pulse_gen_inst.period_counter[23] ),
    .X(_0414_));
 sg13g2_nor2_1 _0994_ (.A(net9),
    .B(_0414_),
    .Y(_0050_));
 sg13g2_inv_1 _0995_ (.Y(_0415_),
    .A(\pulse_gen_inst.period_counter[24] ));
 sg13g2_nand2_1 _0996_ (.Y(_0416_),
    .A(\pulse_gen_inst.period_counter[23] ),
    .B(\pulse_gen_inst.period_counter[22] ));
 sg13g2_or2_1 _0997_ (.X(_0417_),
    .B(_0416_),
    .A(_0411_));
 sg13g2_a21oi_1 _0998_ (.A1(_0415_),
    .A2(_0417_),
    .Y(_0051_),
    .B1(net9));
 sg13g2_nand4_1 _0999_ (.B(\pulse_gen_inst.period_counter[21] ),
    .C(\pulse_gen_inst.period_counter[20] ),
    .A(\pulse_gen_inst.period_counter[24] ),
    .Y(_0418_),
    .D(\pulse_gen_inst.period_counter[19] ));
 sg13g2_nor4_2 _1000_ (.A(_0398_),
    .B(_0402_),
    .C(_0416_),
    .Y(_0419_),
    .D(_0418_));
 sg13g2_xnor2_1 _1001_ (.Y(_0420_),
    .A(\pulse_gen_inst.period_counter[25] ),
    .B(_0419_));
 sg13g2_nor2_1 _1002_ (.A(net9),
    .B(_0420_),
    .Y(_0052_));
 sg13g2_a21oi_1 _1003_ (.A1(\pulse_gen_inst.period_counter[25] ),
    .A2(_0419_),
    .Y(_0421_),
    .B1(\pulse_gen_inst.period_counter[26] ));
 sg13g2_nor2_1 _1004_ (.A(net9),
    .B(_0421_),
    .Y(_0053_));
 sg13g2_and3_1 _1005_ (.X(_0422_),
    .A(\pulse_gen_inst.period_counter[26] ),
    .B(\pulse_gen_inst.period_counter[25] ),
    .C(_0419_));
 sg13g2_xnor2_1 _1006_ (.Y(_0423_),
    .A(\pulse_gen_inst.period_counter[27] ),
    .B(_0422_));
 sg13g2_nor2_1 _1007_ (.A(net9),
    .B(_0423_),
    .Y(_0054_));
 sg13g2_a21oi_1 _1008_ (.A1(\pulse_gen_inst.period_counter[27] ),
    .A2(_0422_),
    .Y(_0424_),
    .B1(\pulse_gen_inst.period_counter[28] ));
 sg13g2_nor2_1 _1009_ (.A(net9),
    .B(_0424_),
    .Y(_0055_));
 sg13g2_and3_1 _1010_ (.X(_0425_),
    .A(\pulse_gen_inst.period_counter[28] ),
    .B(\pulse_gen_inst.period_counter[27] ),
    .C(_0422_));
 sg13g2_xnor2_1 _1011_ (.Y(_0426_),
    .A(\pulse_gen_inst.period_counter[29] ),
    .B(_0425_));
 sg13g2_nor2_1 _1012_ (.A(_0408_),
    .B(_0426_),
    .Y(_0056_));
 sg13g2_nand2_1 _1013_ (.Y(_0427_),
    .A(\pulse_gen_inst.period_counter[0] ),
    .B(\pulse_gen_inst.period_counter[1] ));
 sg13g2_xnor2_1 _1014_ (.Y(_0428_),
    .A(_0010_),
    .B(_0427_));
 sg13g2_nor3_1 _1015_ (.A(net17),
    .B(net11),
    .C(_0428_),
    .Y(_0429_));
 sg13g2_a21o_1 _1016_ (.A2(\pulse_gen_inst.period_counter[2] ),
    .A1(net18),
    .B1(_0429_),
    .X(_0057_));
 sg13g2_a21oi_1 _1017_ (.A1(\pulse_gen_inst.period_counter[29] ),
    .A2(_0425_),
    .Y(_0430_),
    .B1(\pulse_gen_inst.period_counter[30] ));
 sg13g2_nor2_1 _1018_ (.A(_0408_),
    .B(_0430_),
    .Y(_0058_));
 sg13g2_inv_1 _1019_ (.Y(_0431_),
    .A(\pulse_gen_inst.period_counter[31] ));
 sg13g2_nand3_1 _1020_ (.B(\pulse_gen_inst.period_counter[29] ),
    .C(_0425_),
    .A(\pulse_gen_inst.period_counter[30] ),
    .Y(_0432_));
 sg13g2_a21oi_1 _1021_ (.A1(_0431_),
    .A2(_0432_),
    .Y(_0059_),
    .B1(_0376_));
 sg13g2_o21ai_1 _1022_ (.B1(_0101_),
    .Y(_0433_),
    .A1(_0241_),
    .A2(_0367_));
 sg13g2_inv_1 _1023_ (.Y(_0434_),
    .A(_0367_));
 sg13g2_nor4_1 _1024_ (.A(_0181_),
    .B(net17),
    .C(_0241_),
    .D(_0434_),
    .Y(_0435_));
 sg13g2_a21o_1 _1025_ (.A2(_0433_),
    .A1(_0181_),
    .B1(_0435_),
    .X(_0060_));
 sg13g2_nand2_1 _1026_ (.Y(_0436_),
    .A(_0181_),
    .B(_0367_));
 sg13g2_xnor2_1 _1027_ (.Y(_0437_),
    .A(_0009_),
    .B(_0436_));
 sg13g2_nor3_1 _1028_ (.A(net17),
    .B(net11),
    .C(_0437_),
    .Y(_0438_));
 sg13g2_a21o_1 _1029_ (.A2(\pulse_gen_inst.period_counter[4] ),
    .A1(_0254_),
    .B1(_0438_),
    .X(_0061_));
 sg13g2_nand3_1 _1030_ (.B(\pulse_gen_inst.period_counter[4] ),
    .C(_0367_),
    .A(_0181_),
    .Y(_0439_));
 sg13g2_xnor2_1 _1031_ (.Y(_0440_),
    .A(_0008_),
    .B(_0439_));
 sg13g2_nor3_1 _1032_ (.A(net17),
    .B(net11),
    .C(_0440_),
    .Y(_0441_));
 sg13g2_a21o_1 _1033_ (.A2(net18),
    .A1(\pulse_gen_inst.period_counter[5] ),
    .B1(_0441_),
    .X(_0062_));
 sg13g2_nand3_1 _1034_ (.B(_0367_),
    .C(_0368_),
    .A(\pulse_gen_inst.period_counter[5] ),
    .Y(_0442_));
 sg13g2_xnor2_1 _1035_ (.Y(_0443_),
    .A(_0217_),
    .B(_0442_));
 sg13g2_nor3_1 _1036_ (.A(_0272_),
    .B(net11),
    .C(_0443_),
    .Y(_0444_));
 sg13g2_a21o_1 _1037_ (.A2(net18),
    .A1(_0197_),
    .B1(_0444_),
    .X(_0063_));
 sg13g2_o21ai_1 _1038_ (.B1(net31),
    .Y(_0445_),
    .A1(net12),
    .A2(_0370_));
 sg13g2_inv_1 _1039_ (.Y(_0446_),
    .A(_0370_));
 sg13g2_nor4_1 _1040_ (.A(net33),
    .B(_0253_),
    .C(net12),
    .D(_0446_),
    .Y(_0447_));
 sg13g2_a21o_1 _1041_ (.A2(_0445_),
    .A1(_0195_),
    .B1(_0447_),
    .X(_0064_));
 sg13g2_xor2_1 _1042_ (.B(_0372_),
    .A(_0006_),
    .X(_0448_));
 sg13g2_nor3_1 _1043_ (.A(net17),
    .B(net12),
    .C(_0448_),
    .Y(_0449_));
 sg13g2_a21o_1 _1044_ (.A2(\pulse_gen_inst.period_counter[8] ),
    .A1(net18),
    .B1(_0449_),
    .X(_0065_));
 sg13g2_xnor2_1 _1045_ (.Y(_0450_),
    .A(_0005_),
    .B(_0378_));
 sg13g2_nor3_1 _1046_ (.A(net17),
    .B(net12),
    .C(_0450_),
    .Y(_0451_));
 sg13g2_a21o_1 _1047_ (.A2(net18),
    .A1(\pulse_gen_inst.period_counter[9] ),
    .B1(_0451_),
    .X(_0066_));
 sg13g2_nand2b_1 _1048_ (.Y(_0452_),
    .B(net20),
    .A_N(net22));
 sg13g2_nor2b_1 _1049_ (.A(net24),
    .B_N(net22),
    .Y(_0453_));
 sg13g2_a21oi_1 _1050_ (.A1(net19),
    .A2(_0452_),
    .Y(_0454_),
    .B1(_0453_));
 sg13g2_mux2_1 _1051_ (.A0(_0011_),
    .A1(_0454_),
    .S(net23),
    .X(_0455_));
 sg13g2_inv_1 _1052_ (.Y(_0456_),
    .A(_0001_));
 sg13g2_mux2_1 _1053_ (.A0(net25),
    .A1(net24),
    .S(net23),
    .X(_0457_));
 sg13g2_inv_1 _1054_ (.Y(_0458_),
    .A(\pulse_gen_inst.pulse_counter[0] ));
 sg13g2_a21oi_1 _1055_ (.A1(_0456_),
    .A2(_0457_),
    .Y(_0459_),
    .B1(_0458_));
 sg13g2_buf_1 _1056_ (.A(\pulse_gen_inst.pulse_counter[1] ),
    .X(_0460_));
 sg13g2_a21oi_1 _1057_ (.A1(_0455_),
    .A2(_0459_),
    .Y(_0461_),
    .B1(_0460_));
 sg13g2_nor2_1 _1058_ (.A(_0455_),
    .B(_0459_),
    .Y(_0462_));
 sg13g2_a21oi_1 _1059_ (.A1(net20),
    .A2(_0139_),
    .Y(_0463_),
    .B1(_0453_));
 sg13g2_o21ai_1 _1060_ (.B1(net23),
    .Y(_0464_),
    .A1(net24),
    .A2(net22));
 sg13g2_nor2_1 _1061_ (.A(net19),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_a21oi_1 _1062_ (.A1(net19),
    .A2(_0463_),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_xor2_1 _1063_ (.B(_0466_),
    .A(_0016_),
    .X(_0467_));
 sg13g2_o21ai_1 _1064_ (.B1(_0467_),
    .Y(_0468_),
    .A1(_0461_),
    .A2(_0462_));
 sg13g2_inv_1 _1065_ (.Y(_0469_),
    .A(\pulse_gen_inst.pulse_counter[3] ));
 sg13g2_o21ai_1 _1066_ (.B1(_0208_),
    .Y(_0470_),
    .A1(net20),
    .A2(_0232_));
 sg13g2_a21oi_1 _1067_ (.A1(_0189_),
    .A2(_0267_),
    .Y(_0471_),
    .B1(_0191_));
 sg13g2_a21o_1 _1068_ (.A2(_0470_),
    .A1(_0121_),
    .B1(_0471_),
    .X(_0472_));
 sg13g2_inv_1 _1069_ (.Y(_0473_),
    .A(\pulse_gen_inst.pulse_counter[2] ));
 sg13g2_a22oi_1 _1070_ (.Y(_0474_),
    .B1(_0466_),
    .B2(_0473_),
    .A2(_0472_),
    .A1(_0469_));
 sg13g2_xnor2_1 _1071_ (.Y(_0475_),
    .A(net19),
    .B(_0199_));
 sg13g2_a22oi_1 _1072_ (.Y(_0476_),
    .B1(_0475_),
    .B2(_0191_),
    .A2(_0165_),
    .A1(_0011_));
 sg13g2_xor2_1 _1073_ (.B(_0476_),
    .A(_0015_),
    .X(_0477_));
 sg13g2_nor2_1 _1074_ (.A(net24),
    .B(net26),
    .Y(_0478_));
 sg13g2_a221oi_1 _1075_ (.B2(net20),
    .C1(_0478_),
    .B1(_0304_),
    .A1(_0121_),
    .Y(_0479_),
    .A2(net22));
 sg13g2_xnor2_1 _1076_ (.Y(_0480_),
    .A(_0013_),
    .B(_0479_));
 sg13g2_inv_1 _1077_ (.Y(_0481_),
    .A(\pulse_gen_inst.pulse_counter[7] ));
 sg13g2_a21oi_1 _1078_ (.A1(net20),
    .A2(_0176_),
    .Y(_0482_),
    .B1(net25));
 sg13g2_nand2_1 _1079_ (.Y(_0483_),
    .A(net22),
    .B(_0209_));
 sg13g2_mux2_1 _1080_ (.A0(_0011_),
    .A1(net23),
    .S(net25),
    .X(_0484_));
 sg13g2_nand2_1 _1081_ (.Y(_0485_),
    .A(_0171_),
    .B(_0484_));
 sg13g2_o21ai_1 _1082_ (.B1(_0485_),
    .Y(_0486_),
    .A1(_0482_),
    .A2(_0483_));
 sg13g2_xnor2_1 _1083_ (.Y(_0487_),
    .A(_0481_),
    .B(_0486_));
 sg13g2_a21oi_1 _1084_ (.A1(_0121_),
    .A2(_0470_),
    .Y(_0488_),
    .B1(_0471_));
 sg13g2_o21ai_1 _1085_ (.B1(net25),
    .Y(_0489_),
    .A1(net24),
    .A2(net23));
 sg13g2_nand3_1 _1086_ (.B(_0140_),
    .C(_0489_),
    .A(_0171_),
    .Y(_0490_));
 sg13g2_nand3b_1 _1087_ (.B(net24),
    .C(net26),
    .Y(_0491_),
    .A_N(net25));
 sg13g2_nand3b_1 _1088_ (.B(_0491_),
    .C(net22),
    .Y(_0492_),
    .A_N(_0478_));
 sg13g2_inv_1 _1089_ (.Y(_0493_),
    .A(_0014_));
 sg13g2_a21o_1 _1090_ (.A2(_0492_),
    .A1(_0490_),
    .B1(_0493_),
    .X(_0494_));
 sg13g2_nand3_1 _1091_ (.B(_0490_),
    .C(_0492_),
    .A(_0493_),
    .Y(_0495_));
 sg13g2_a22oi_1 _1092_ (.Y(_0496_),
    .B1(_0494_),
    .B2(_0495_),
    .A2(_0488_),
    .A1(\pulse_gen_inst.pulse_counter[3] ));
 sg13g2_nand4_1 _1093_ (.B(_0480_),
    .C(_0487_),
    .A(_0477_),
    .Y(_0497_),
    .D(_0496_));
 sg13g2_a21o_1 _1094_ (.A2(_0474_),
    .A1(_0468_),
    .B1(_0497_),
    .X(_0498_));
 sg13g2_a221oi_1 _1095_ (.B2(net25),
    .C1(_0165_),
    .B1(_0196_),
    .A1(_0117_),
    .Y(_0499_),
    .A2(_0133_));
 sg13g2_buf_1 _1096_ (.A(_0499_),
    .X(_0500_));
 sg13g2_or4_1 _1097_ (.A(\pulse_gen_inst.pulse_counter[12] ),
    .B(\pulse_gen_inst.pulse_counter[11] ),
    .C(\pulse_gen_inst.pulse_counter[10] ),
    .D(\pulse_gen_inst.pulse_counter[9] ),
    .X(_0501_));
 sg13g2_nor4_2 _1098_ (.A(\pulse_gen_inst.pulse_counter[14] ),
    .B(\pulse_gen_inst.pulse_counter[15] ),
    .C(\pulse_gen_inst.pulse_counter[13] ),
    .Y(_0502_),
    .D(_0501_));
 sg13g2_nor2b_1 _1099_ (.A(\pulse_gen_inst.pulse_counter[8] ),
    .B_N(_0502_),
    .Y(_0503_));
 sg13g2_nand2_1 _1100_ (.Y(_0504_),
    .A(_0015_),
    .B(_0476_));
 sg13g2_and2_1 _1101_ (.A(_0494_),
    .B(_0495_),
    .X(_0505_));
 sg13g2_nand3b_1 _1102_ (.B(_0490_),
    .C(_0492_),
    .Y(_0506_),
    .A_N(\pulse_gen_inst.pulse_counter[5] ));
 sg13g2_o21ai_1 _1103_ (.B1(_0506_),
    .Y(_0507_),
    .A1(_0504_),
    .A2(_0505_));
 sg13g2_and2_1 _1104_ (.A(_0480_),
    .B(_0487_),
    .X(_0508_));
 sg13g2_or2_1 _1105_ (.X(_0509_),
    .B(_0479_),
    .A(\pulse_gen_inst.pulse_counter[6] ));
 sg13g2_o21ai_1 _1106_ (.B1(_0486_),
    .Y(_0510_),
    .A1(\pulse_gen_inst.pulse_counter[7] ),
    .A2(_0509_));
 sg13g2_nand2_1 _1107_ (.Y(_0511_),
    .A(\pulse_gen_inst.pulse_counter[7] ),
    .B(_0509_));
 sg13g2_and2_1 _1108_ (.A(_0510_),
    .B(_0511_),
    .X(_0512_));
 sg13g2_a221oi_1 _1109_ (.B2(_0508_),
    .C1(_0512_),
    .B1(_0507_),
    .A1(_0500_),
    .Y(_0513_),
    .A2(_0503_));
 sg13g2_xor2_1 _1110_ (.B(_0455_),
    .A(_0460_),
    .X(_0514_));
 sg13g2_nand2b_1 _1111_ (.Y(_0515_),
    .B(_0012_),
    .A_N(_0500_));
 sg13g2_nand2b_1 _1112_ (.Y(_0516_),
    .B(_0500_),
    .A_N(_0012_));
 sg13g2_nand3_1 _1113_ (.B(_0458_),
    .C(_0457_),
    .A(_0456_),
    .Y(_0517_));
 sg13g2_nand3b_1 _1114_ (.B(_0502_),
    .C(_0517_),
    .Y(_0518_),
    .A_N(_0459_));
 sg13g2_a221oi_1 _1115_ (.B2(_0516_),
    .C1(_0518_),
    .B1(_0515_),
    .A1(_0469_),
    .Y(_0519_),
    .A2(_0472_));
 sg13g2_nand3_1 _1116_ (.B(_0514_),
    .C(_0519_),
    .A(_0467_),
    .Y(_0520_));
 sg13g2_and3_1 _1117_ (.X(_0521_),
    .A(\pulse_gen_inst.pulse_counter[8] ),
    .B(_0012_),
    .C(_0500_));
 sg13g2_nor2_1 _1118_ (.A(_0012_),
    .B(_0500_),
    .Y(_0522_));
 sg13g2_nor4_1 _1119_ (.A(\pulse_gen_inst.pulse_counter[31] ),
    .B(\pulse_gen_inst.pulse_counter[29] ),
    .C(\pulse_gen_inst.pulse_counter[28] ),
    .D(\pulse_gen_inst.pulse_counter[27] ),
    .Y(_0523_));
 sg13g2_nor2_1 _1120_ (.A(\pulse_gen_inst.pulse_counter[26] ),
    .B(\pulse_gen_inst.pulse_counter[21] ),
    .Y(_0524_));
 sg13g2_nand3_1 _1121_ (.B(_0523_),
    .C(_0524_),
    .A(_0502_),
    .Y(_0525_));
 sg13g2_nor4_1 _1122_ (.A(\pulse_gen_inst.pulse_counter[25] ),
    .B(\pulse_gen_inst.pulse_counter[24] ),
    .C(\pulse_gen_inst.pulse_counter[23] ),
    .D(\pulse_gen_inst.pulse_counter[22] ),
    .Y(_0526_));
 sg13g2_nor4_1 _1123_ (.A(\pulse_gen_inst.pulse_counter[30] ),
    .B(\pulse_gen_inst.pulse_counter[20] ),
    .C(\pulse_gen_inst.pulse_counter[19] ),
    .D(\pulse_gen_inst.pulse_counter[18] ),
    .Y(_0527_));
 sg13g2_nor3_1 _1124_ (.A(\pulse_gen_inst.pulse_counter[17] ),
    .B(\pulse_gen_inst.pulse_counter[16] ),
    .C(net21),
    .Y(_0528_));
 sg13g2_nand3_1 _1125_ (.B(_0527_),
    .C(_0528_),
    .A(_0526_),
    .Y(_0529_));
 sg13g2_nor4_1 _1126_ (.A(_0521_),
    .B(_0522_),
    .C(_0525_),
    .D(_0529_),
    .Y(_0530_));
 sg13g2_o21ai_1 _1127_ (.B1(_0530_),
    .Y(_0531_),
    .A1(_0497_),
    .A2(_0520_));
 sg13g2_a21oi_2 _1128_ (.B1(_0531_),
    .Y(_0532_),
    .A2(_0513_),
    .A1(_0498_));
 sg13g2_nand2_2 _1129_ (.Y(_0533_),
    .A(_0364_),
    .B(_0532_));
 sg13g2_o21ai_1 _1130_ (.B1(_0100_),
    .Y(_0534_),
    .A1(_0149_),
    .A2(_0238_));
 sg13g2_buf_1 _1131_ (.A(_0534_),
    .X(_0535_));
 sg13g2_a221oi_1 _1132_ (.B2(_0516_),
    .C1(_0518_),
    .B1(_0515_),
    .A1(_0469_),
    .Y(_0536_),
    .A2(_0472_));
 sg13g2_nand3_1 _1133_ (.B(_0514_),
    .C(_0536_),
    .A(_0467_),
    .Y(_0537_));
 sg13g2_nor4_1 _1134_ (.A(\pulse_gen_inst.pulse_counter[24] ),
    .B(\pulse_gen_inst.pulse_counter[23] ),
    .C(\pulse_gen_inst.pulse_counter[22] ),
    .D(\pulse_gen_inst.pulse_counter[21] ),
    .Y(_0538_));
 sg13g2_nor4_1 _1135_ (.A(\pulse_gen_inst.pulse_counter[31] ),
    .B(\pulse_gen_inst.pulse_counter[19] ),
    .C(\pulse_gen_inst.pulse_counter[18] ),
    .D(\pulse_gen_inst.pulse_counter[17] ),
    .Y(_0539_));
 sg13g2_nor3_1 _1136_ (.A(\pulse_gen_inst.pulse_counter[30] ),
    .B(\pulse_gen_inst.pulse_counter[16] ),
    .C(_0252_),
    .Y(_0540_));
 sg13g2_nand3_1 _1137_ (.B(_0539_),
    .C(_0540_),
    .A(_0538_),
    .Y(_0541_));
 sg13g2_nor2_1 _1138_ (.A(\pulse_gen_inst.pulse_counter[29] ),
    .B(\pulse_gen_inst.pulse_counter[20] ),
    .Y(_0542_));
 sg13g2_nor4_1 _1139_ (.A(\pulse_gen_inst.pulse_counter[28] ),
    .B(\pulse_gen_inst.pulse_counter[27] ),
    .C(\pulse_gen_inst.pulse_counter[26] ),
    .D(\pulse_gen_inst.pulse_counter[25] ),
    .Y(_0543_));
 sg13g2_nand3_1 _1140_ (.B(_0542_),
    .C(_0543_),
    .A(_0502_),
    .Y(_0544_));
 sg13g2_nor4_1 _1141_ (.A(_0521_),
    .B(_0522_),
    .C(_0541_),
    .D(_0544_),
    .Y(_0545_));
 sg13g2_o21ai_1 _1142_ (.B1(_0545_),
    .Y(_0546_),
    .A1(_0497_),
    .A2(_0537_));
 sg13g2_a21o_1 _1143_ (.A2(_0513_),
    .A1(_0498_),
    .B1(_0546_),
    .X(_0547_));
 sg13g2_buf_1 _1144_ (.A(_0547_),
    .X(_0548_));
 sg13g2_nand3_1 _1145_ (.B(net14),
    .C(net13),
    .A(\pulse_gen_inst.pulse_counter[0] ),
    .Y(_0549_));
 sg13g2_o21ai_1 _1146_ (.B1(_0549_),
    .Y(_0067_),
    .A1(\pulse_gen_inst.pulse_counter[0] ),
    .A2(_0533_));
 sg13g2_buf_1 _1147_ (.A(net14),
    .X(_0550_));
 sg13g2_and2_1 _1148_ (.A(\pulse_gen_inst.pulse_counter[10] ),
    .B(net8),
    .X(_0068_));
 sg13g2_and2_1 _1149_ (.A(\pulse_gen_inst.pulse_counter[11] ),
    .B(_0550_),
    .X(_0069_));
 sg13g2_and2_1 _1150_ (.A(\pulse_gen_inst.pulse_counter[12] ),
    .B(net8),
    .X(_0070_));
 sg13g2_and2_1 _1151_ (.A(\pulse_gen_inst.pulse_counter[13] ),
    .B(net8),
    .X(_0071_));
 sg13g2_and2_1 _1152_ (.A(\pulse_gen_inst.pulse_counter[14] ),
    .B(net8),
    .X(_0072_));
 sg13g2_and2_1 _1153_ (.A(\pulse_gen_inst.pulse_counter[15] ),
    .B(net8),
    .X(_0073_));
 sg13g2_and2_1 _1154_ (.A(\pulse_gen_inst.pulse_counter[16] ),
    .B(_0550_),
    .X(_0074_));
 sg13g2_and2_1 _1155_ (.A(\pulse_gen_inst.pulse_counter[17] ),
    .B(net8),
    .X(_0075_));
 sg13g2_and2_1 _1156_ (.A(\pulse_gen_inst.pulse_counter[18] ),
    .B(net8),
    .X(_0076_));
 sg13g2_and2_1 _1157_ (.A(\pulse_gen_inst.pulse_counter[19] ),
    .B(net8),
    .X(_0077_));
 sg13g2_o21ai_1 _1158_ (.B1(_0460_),
    .Y(_0551_),
    .A1(_0458_),
    .A2(net13));
 sg13g2_nand3b_1 _1159_ (.B(\pulse_gen_inst.pulse_counter[0] ),
    .C(_0532_),
    .Y(_0552_),
    .A_N(_0460_));
 sg13g2_a21oi_1 _1160_ (.A1(_0551_),
    .A2(_0552_),
    .Y(_0078_),
    .B1(_0376_));
 sg13g2_buf_1 _1161_ (.A(net14),
    .X(_0553_));
 sg13g2_and2_1 _1162_ (.A(\pulse_gen_inst.pulse_counter[20] ),
    .B(net7),
    .X(_0079_));
 sg13g2_and2_1 _1163_ (.A(\pulse_gen_inst.pulse_counter[21] ),
    .B(net7),
    .X(_0080_));
 sg13g2_and2_1 _1164_ (.A(\pulse_gen_inst.pulse_counter[22] ),
    .B(_0553_),
    .X(_0081_));
 sg13g2_and2_1 _1165_ (.A(\pulse_gen_inst.pulse_counter[23] ),
    .B(net7),
    .X(_0082_));
 sg13g2_and2_1 _1166_ (.A(\pulse_gen_inst.pulse_counter[24] ),
    .B(net7),
    .X(_0083_));
 sg13g2_and2_1 _1167_ (.A(\pulse_gen_inst.pulse_counter[25] ),
    .B(net7),
    .X(_0084_));
 sg13g2_and2_1 _1168_ (.A(\pulse_gen_inst.pulse_counter[26] ),
    .B(net7),
    .X(_0085_));
 sg13g2_and2_1 _1169_ (.A(\pulse_gen_inst.pulse_counter[27] ),
    .B(_0553_),
    .X(_0086_));
 sg13g2_and2_1 _1170_ (.A(\pulse_gen_inst.pulse_counter[28] ),
    .B(net7),
    .X(_0087_));
 sg13g2_and2_1 _1171_ (.A(\pulse_gen_inst.pulse_counter[29] ),
    .B(net7),
    .X(_0088_));
 sg13g2_nand2_1 _1172_ (.Y(_0554_),
    .A(_0460_),
    .B(\pulse_gen_inst.pulse_counter[0] ));
 sg13g2_xnor2_1 _1173_ (.Y(_0555_),
    .A(_0016_),
    .B(_0554_));
 sg13g2_nand3_1 _1174_ (.B(net14),
    .C(net13),
    .A(\pulse_gen_inst.pulse_counter[2] ),
    .Y(_0556_));
 sg13g2_o21ai_1 _1175_ (.B1(_0556_),
    .Y(_0089_),
    .A1(_0533_),
    .A2(_0555_));
 sg13g2_and2_1 _1176_ (.A(\pulse_gen_inst.pulse_counter[30] ),
    .B(net14),
    .X(_0090_));
 sg13g2_and2_1 _1177_ (.A(\pulse_gen_inst.pulse_counter[31] ),
    .B(net14),
    .X(_0091_));
 sg13g2_nand3_1 _1178_ (.B(_0460_),
    .C(\pulse_gen_inst.pulse_counter[0] ),
    .A(\pulse_gen_inst.pulse_counter[2] ),
    .Y(_0557_));
 sg13g2_o21ai_1 _1179_ (.B1(\pulse_gen_inst.pulse_counter[3] ),
    .Y(_0558_),
    .A1(net13),
    .A2(_0557_));
 sg13g2_or3_1 _1180_ (.A(\pulse_gen_inst.pulse_counter[3] ),
    .B(net13),
    .C(_0557_),
    .X(_0559_));
 sg13g2_a21oi_1 _1181_ (.A1(_0558_),
    .A2(_0559_),
    .Y(_0092_),
    .B1(_0376_));
 sg13g2_nor2_1 _1182_ (.A(_0469_),
    .B(_0557_),
    .Y(_0560_));
 sg13g2_xor2_1 _1183_ (.B(_0560_),
    .A(_0015_),
    .X(_0561_));
 sg13g2_nand3_1 _1184_ (.B(net14),
    .C(net13),
    .A(\pulse_gen_inst.pulse_counter[4] ),
    .Y(_0562_));
 sg13g2_o21ai_1 _1185_ (.B1(_0562_),
    .Y(_0093_),
    .A1(_0533_),
    .A2(_0561_));
 sg13g2_and2_1 _1186_ (.A(\pulse_gen_inst.pulse_counter[4] ),
    .B(_0560_),
    .X(_0563_));
 sg13g2_xnor2_1 _1187_ (.Y(_0564_),
    .A(_0493_),
    .B(_0563_));
 sg13g2_nand3_1 _1188_ (.B(_0535_),
    .C(net13),
    .A(\pulse_gen_inst.pulse_counter[5] ),
    .Y(_0565_));
 sg13g2_o21ai_1 _1189_ (.B1(_0565_),
    .Y(_0094_),
    .A1(_0533_),
    .A2(_0564_));
 sg13g2_nand2_1 _1190_ (.Y(_0566_),
    .A(\pulse_gen_inst.pulse_counter[5] ),
    .B(_0563_));
 sg13g2_xnor2_1 _1191_ (.Y(_0567_),
    .A(_0013_),
    .B(_0566_));
 sg13g2_nand3_1 _1192_ (.B(_0535_),
    .C(_0548_),
    .A(\pulse_gen_inst.pulse_counter[6] ),
    .Y(_0568_));
 sg13g2_o21ai_1 _1193_ (.B1(_0568_),
    .Y(_0095_),
    .A1(_0533_),
    .A2(_0567_));
 sg13g2_and3_1 _1194_ (.X(_0569_),
    .A(\pulse_gen_inst.pulse_counter[6] ),
    .B(\pulse_gen_inst.pulse_counter[5] ),
    .C(_0563_));
 sg13g2_nand3_1 _1195_ (.B(_0532_),
    .C(_0569_),
    .A(_0364_),
    .Y(_0570_));
 sg13g2_nor2_1 _1196_ (.A(_0481_),
    .B(net17),
    .Y(_0571_));
 sg13g2_a21o_1 _1197_ (.A2(_0569_),
    .A1(_0532_),
    .B1(net11),
    .X(_0572_));
 sg13g2_a22oi_1 _1198_ (.Y(_0096_),
    .B1(_0571_),
    .B2(_0572_),
    .A2(_0570_),
    .A1(_0481_));
 sg13g2_nand2_1 _1199_ (.Y(_0573_),
    .A(\pulse_gen_inst.pulse_counter[7] ),
    .B(_0569_));
 sg13g2_xnor2_1 _1200_ (.Y(_0574_),
    .A(_0012_),
    .B(_0573_));
 sg13g2_nand3_1 _1201_ (.B(net14),
    .C(net13),
    .A(\pulse_gen_inst.pulse_counter[8] ),
    .Y(_0575_));
 sg13g2_o21ai_1 _1202_ (.B1(_0575_),
    .Y(_0097_),
    .A1(_0533_),
    .A2(_0574_));
 sg13g2_inv_1 _1203_ (.Y(_0576_),
    .A(\pulse_gen_inst.pulse_counter[9] ));
 sg13g2_nand4_1 _1204_ (.B(\pulse_gen_inst.pulse_counter[7] ),
    .C(_0532_),
    .A(\pulse_gen_inst.pulse_counter[8] ),
    .Y(_0577_),
    .D(_0569_));
 sg13g2_a21oi_1 _1205_ (.A1(_0576_),
    .A2(_0577_),
    .Y(_0098_),
    .B1(_0376_));
 sg13g2_a21o_1 _1206_ (.A2(\pulse_gen_inst.ttl_out ),
    .A1(net18),
    .B1(_0532_),
    .X(_0099_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _1208_ (.A(net53),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1209_ (.A(net54),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1210_ (.A(net55),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1211_ (.A(net56),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1212_ (.A(net57),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1213_ (.A(net58),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1214_ (.A(net59),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1215_ (.A(net60),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1216_ (.A(net61),
    .X(uio_out[0]));
 sg13g2_buf_1 _1217_ (.A(net62),
    .X(uio_out[1]));
 sg13g2_buf_1 _1218_ (.A(net63),
    .X(uio_out[2]));
 sg13g2_buf_1 _1219_ (.A(net64),
    .X(uio_out[3]));
 sg13g2_buf_1 _1220_ (.A(net65),
    .X(uio_out[4]));
 sg13g2_buf_1 _1221_ (.A(net66),
    .X(uio_out[5]));
 sg13g2_buf_1 _1222_ (.A(net67),
    .X(uio_out[6]));
 sg13g2_buf_1 _1223_ (.A(net68),
    .X(uio_out[7]));
 sg13g2_buf_1 _1224_ (.A(\pulse_gen_inst.ttl_out ),
    .X(net6));
 sg13g2_buf_1 _1225_ (.A(net69),
    .X(uo_out[1]));
 sg13g2_buf_1 _1226_ (.A(net70),
    .X(uo_out[2]));
 sg13g2_buf_1 _1227_ (.A(net71),
    .X(uo_out[3]));
 sg13g2_buf_1 _1228_ (.A(net72),
    .X(uo_out[4]));
 sg13g2_buf_1 _1229_ (.A(net73),
    .X(uo_out[5]));
 sg13g2_buf_1 _1230_ (.A(net74),
    .X(uo_out[6]));
 sg13g2_buf_1 _1231_ (.A(net75),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[0]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net46),
    .D(_0019_),
    .Q_N(_0018_),
    .Q(\pulse_gen_inst.count_counter[0] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[10]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net46),
    .D(_0020_),
    .Q_N(_0644_),
    .Q(\pulse_gen_inst.count_counter[10] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[11]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net46),
    .D(_0021_),
    .Q_N(_0643_),
    .Q(\pulse_gen_inst.count_counter[11] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[12]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net46),
    .D(_0022_),
    .Q_N(_0642_),
    .Q(\pulse_gen_inst.count_counter[12] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[13]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net39),
    .D(_0023_),
    .Q_N(_0641_),
    .Q(\pulse_gen_inst.count_counter[13] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[14]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net39),
    .D(_0024_),
    .Q_N(_0640_),
    .Q(\pulse_gen_inst.count_counter[14] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[15]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net46),
    .D(_0025_),
    .Q_N(_0639_),
    .Q(\pulse_gen_inst.count_counter[15] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[1]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net48),
    .D(_0026_),
    .Q_N(_0638_),
    .Q(\pulse_gen_inst.count_counter[1] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[2]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(_0027_),
    .Q_N(_0637_),
    .Q(\pulse_gen_inst.count_counter[2] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[3]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(_0028_),
    .Q_N(_0636_),
    .Q(\pulse_gen_inst.count_counter[3] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[4]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(_0029_),
    .Q_N(_0635_),
    .Q(\pulse_gen_inst.count_counter[4] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[5]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net48),
    .D(_0030_),
    .Q_N(_0634_),
    .Q(\pulse_gen_inst.count_counter[5] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[6]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net46),
    .D(_0031_),
    .Q_N(_0633_),
    .Q(\pulse_gen_inst.count_counter[6] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[7]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net48),
    .D(_0032_),
    .Q_N(_0632_),
    .Q(\pulse_gen_inst.count_counter[7] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[8]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net48),
    .D(_0033_),
    .Q_N(_0631_),
    .Q(\pulse_gen_inst.count_counter[8] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.count_counter[9]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net48),
    .D(_0034_),
    .Q_N(_0630_),
    .Q(\pulse_gen_inst.count_counter[9] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[0]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net47),
    .D(_0035_),
    .Q_N(_0629_),
    .Q(\pulse_gen_inst.period_counter[0] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[10]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net51),
    .D(_0036_),
    .Q_N(_0003_),
    .Q(\pulse_gen_inst.period_counter[10] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[11]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net45),
    .D(_0037_),
    .Q_N(_0628_),
    .Q(\pulse_gen_inst.period_counter[11] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[12]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net39),
    .D(_0038_),
    .Q_N(_0627_),
    .Q(\pulse_gen_inst.period_counter[12] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[13]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net39),
    .D(_0039_),
    .Q_N(_0626_),
    .Q(\pulse_gen_inst.period_counter[13] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[14]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net40),
    .D(_0040_),
    .Q_N(_0625_),
    .Q(\pulse_gen_inst.period_counter[14] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[15]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net40),
    .D(_0041_),
    .Q_N(_0624_),
    .Q(\pulse_gen_inst.period_counter[15] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[16]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net46),
    .D(_0042_),
    .Q_N(_0623_),
    .Q(\pulse_gen_inst.period_counter[16] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[17]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net39),
    .D(_0043_),
    .Q_N(_0622_),
    .Q(\pulse_gen_inst.period_counter[17] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[18]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net39),
    .D(_0044_),
    .Q_N(_0621_),
    .Q(\pulse_gen_inst.period_counter[18] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[19]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net39),
    .D(_0045_),
    .Q_N(_0620_),
    .Q(\pulse_gen_inst.period_counter[19] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[1]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net40),
    .D(_0046_),
    .Q_N(_0619_),
    .Q(\pulse_gen_inst.period_counter[1] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[20]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net39),
    .D(_0047_),
    .Q_N(_0618_),
    .Q(\pulse_gen_inst.period_counter[20] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[21]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net37),
    .D(_0048_),
    .Q_N(_0617_),
    .Q(\pulse_gen_inst.period_counter[21] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[22]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net37),
    .D(_0049_),
    .Q_N(_0616_),
    .Q(\pulse_gen_inst.period_counter[22] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[23]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net37),
    .D(_0050_),
    .Q_N(_0615_),
    .Q(\pulse_gen_inst.period_counter[23] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[24]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net37),
    .D(_0051_),
    .Q_N(_0614_),
    .Q(\pulse_gen_inst.period_counter[24] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[25]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net37),
    .D(_0052_),
    .Q_N(_0613_),
    .Q(\pulse_gen_inst.period_counter[25] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[26]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net37),
    .D(_0053_),
    .Q_N(_0612_),
    .Q(\pulse_gen_inst.period_counter[26] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[27]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net37),
    .D(_0054_),
    .Q_N(_0611_),
    .Q(\pulse_gen_inst.period_counter[27] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[28]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net37),
    .D(_0055_),
    .Q_N(_0610_),
    .Q(\pulse_gen_inst.period_counter[28] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[29]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net38),
    .D(_0056_),
    .Q_N(_0609_),
    .Q(\pulse_gen_inst.period_counter[29] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[2]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net47),
    .D(_0057_),
    .Q_N(_0010_),
    .Q(\pulse_gen_inst.period_counter[2] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[30]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net40),
    .D(_0058_),
    .Q_N(_0608_),
    .Q(\pulse_gen_inst.period_counter[30] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[31]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net40),
    .D(_0059_),
    .Q_N(_0607_),
    .Q(\pulse_gen_inst.period_counter[31] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[3]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net49),
    .D(_0060_),
    .Q_N(_0606_),
    .Q(\pulse_gen_inst.period_counter[3] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[4]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net49),
    .D(_0061_),
    .Q_N(_0009_),
    .Q(\pulse_gen_inst.period_counter[4] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[5]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net49),
    .D(_0062_),
    .Q_N(_0008_),
    .Q(\pulse_gen_inst.period_counter[5] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[6]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net51),
    .D(_0063_),
    .Q_N(_0007_),
    .Q(\pulse_gen_inst.period_counter[6] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[7]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net49),
    .D(_0064_),
    .Q_N(_0605_),
    .Q(\pulse_gen_inst.period_counter[7] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[8]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net47),
    .D(_0065_),
    .Q_N(_0006_),
    .Q(\pulse_gen_inst.period_counter[8] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.period_counter[9]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net47),
    .D(_0066_),
    .Q_N(_0005_),
    .Q(\pulse_gen_inst.period_counter[9] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_active$_DFF_PN0_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net46),
    .D(_0000_),
    .Q_N(_0017_),
    .Q(\pulse_gen_inst.pulse_active ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[0]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net43),
    .D(_0067_),
    .Q_N(_0604_),
    .Q(\pulse_gen_inst.pulse_counter[0] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[10]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net38),
    .D(_0068_),
    .Q_N(_0603_),
    .Q(\pulse_gen_inst.pulse_counter[10] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[11]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net38),
    .D(_0069_),
    .Q_N(_0602_),
    .Q(\pulse_gen_inst.pulse_counter[11] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[12]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net38),
    .D(_0070_),
    .Q_N(_0601_),
    .Q(\pulse_gen_inst.pulse_counter[12] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[13]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net38),
    .D(_0071_),
    .Q_N(_0600_),
    .Q(\pulse_gen_inst.pulse_counter[13] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[14]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net38),
    .D(_0072_),
    .Q_N(_0599_),
    .Q(\pulse_gen_inst.pulse_counter[14] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[15]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net42),
    .D(_0073_),
    .Q_N(_0598_),
    .Q(\pulse_gen_inst.pulse_counter[15] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[16]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net42),
    .D(_0074_),
    .Q_N(_0597_),
    .Q(\pulse_gen_inst.pulse_counter[16] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[17]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net42),
    .D(_0075_),
    .Q_N(_0596_),
    .Q(\pulse_gen_inst.pulse_counter[17] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[18]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net42),
    .D(_0076_),
    .Q_N(_0595_),
    .Q(\pulse_gen_inst.pulse_counter[18] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[19]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net42),
    .D(_0077_),
    .Q_N(_0594_),
    .Q(\pulse_gen_inst.pulse_counter[19] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[1]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net43),
    .D(_0078_),
    .Q_N(_0593_),
    .Q(\pulse_gen_inst.pulse_counter[1] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[20]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net43),
    .D(_0079_),
    .Q_N(_0592_),
    .Q(\pulse_gen_inst.pulse_counter[20] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[21]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net43),
    .D(_0080_),
    .Q_N(_0591_),
    .Q(\pulse_gen_inst.pulse_counter[21] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[22]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net42),
    .D(_0081_),
    .Q_N(_0590_),
    .Q(\pulse_gen_inst.pulse_counter[22] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[23]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net42),
    .D(_0082_),
    .Q_N(_0589_),
    .Q(\pulse_gen_inst.pulse_counter[23] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[24]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net42),
    .D(_0083_),
    .Q_N(_0588_),
    .Q(\pulse_gen_inst.pulse_counter[24] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[25]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net43),
    .D(_0084_),
    .Q_N(_0587_),
    .Q(\pulse_gen_inst.pulse_counter[25] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[26]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net44),
    .D(_0085_),
    .Q_N(_0586_),
    .Q(\pulse_gen_inst.pulse_counter[26] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[27]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net44),
    .D(_0086_),
    .Q_N(_0585_),
    .Q(\pulse_gen_inst.pulse_counter[27] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[28]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net44),
    .D(_0087_),
    .Q_N(_0584_),
    .Q(\pulse_gen_inst.pulse_counter[28] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[29]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net44),
    .D(_0088_),
    .Q_N(_0583_),
    .Q(\pulse_gen_inst.pulse_counter[29] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[2]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net45),
    .D(_0089_),
    .Q_N(_0016_),
    .Q(\pulse_gen_inst.pulse_counter[2] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[30]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net43),
    .D(_0090_),
    .Q_N(_0582_),
    .Q(\pulse_gen_inst.pulse_counter[30] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[31]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net43),
    .D(_0091_),
    .Q_N(_0581_),
    .Q(\pulse_gen_inst.pulse_counter[31] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[3]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net45),
    .D(_0092_),
    .Q_N(_0580_),
    .Q(\pulse_gen_inst.pulse_counter[3] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[4]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net51),
    .D(_0093_),
    .Q_N(_0015_),
    .Q(\pulse_gen_inst.pulse_counter[4] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[5]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net51),
    .D(_0094_),
    .Q_N(_0014_),
    .Q(\pulse_gen_inst.pulse_counter[5] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[6]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net51),
    .D(_0095_),
    .Q_N(_0013_),
    .Q(\pulse_gen_inst.pulse_counter[6] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[7]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net45),
    .D(_0096_),
    .Q_N(_0579_),
    .Q(\pulse_gen_inst.pulse_counter[7] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[8]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net45),
    .D(_0097_),
    .Q_N(_0012_),
    .Q(\pulse_gen_inst.pulse_counter[8] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.pulse_counter[9]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net45),
    .D(_0098_),
    .Q_N(_0578_),
    .Q(\pulse_gen_inst.pulse_counter[9] ));
 sg13g2_dfrbp_1 \pulse_gen_inst.ttl_out$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net51),
    .D(_0099_),
    .Q_N(_0645_),
    .Q(\pulse_gen_inst.ttl_out ));
 sg13g2_dfrbp_1 \reg_sequence_select[0]$_DFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net51),
    .D(net2),
    .Q_N(_0004_),
    .Q(\reg_sequence_select[0] ));
 sg13g2_dfrbp_1 \reg_sequence_select[1]$_DFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net52),
    .D(net3),
    .Q_N(_0011_),
    .Q(\reg_sequence_select[1] ));
 sg13g2_dfrbp_1 \reg_sequence_select[2]$_DFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net52),
    .D(net4),
    .Q_N(_0002_),
    .Q(\reg_sequence_select[2] ));
 sg13g2_dfrbp_1 \reg_sequence_select[3]$_DFF_PN0_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net51),
    .D(net5),
    .Q_N(_0001_),
    .Q(\reg_sequence_select[3] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[0]));
 sg13g2_buf_2 fanout7 (.A(_0553_),
    .X(net7));
 sg13g2_buf_2 fanout8 (.A(_0550_),
    .X(net8));
 sg13g2_buf_2 fanout9 (.A(_0408_),
    .X(net9));
 sg13g2_buf_2 fanout10 (.A(_0377_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_0299_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0241_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0548_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0535_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0274_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0264_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0272_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0254_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0216_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0265_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0253_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0228_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0191_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0186_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0175_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0187_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0129_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0127_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0115_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0108_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0101_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0255_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0195_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0111_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0104_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0100_),
    .X(net36));
 sg13g2_buf_4 fanout37 (.X(net37),
    .A(net41));
 sg13g2_buf_2 fanout38 (.A(net41),
    .X(net38));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(net41));
 sg13g2_buf_2 fanout40 (.A(net41),
    .X(net40));
 sg13g2_buf_1 fanout41 (.A(net1),
    .X(net41));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(net43));
 sg13g2_buf_4 fanout43 (.X(net43),
    .A(net45));
 sg13g2_buf_2 fanout44 (.A(net45),
    .X(net44));
 sg13g2_buf_4 fanout45 (.X(net45),
    .A(net1));
 sg13g2_buf_4 fanout46 (.X(net46),
    .A(net50));
 sg13g2_buf_2 fanout47 (.A(net50),
    .X(net47));
 sg13g2_buf_4 fanout48 (.X(net48),
    .A(net50));
 sg13g2_buf_2 fanout49 (.A(net50),
    .X(net49));
 sg13g2_buf_1 fanout50 (.A(net52),
    .X(net50));
 sg13g2_buf_4 fanout51 (.X(net51),
    .A(net52));
 sg13g2_buf_1 fanout52 (.A(net1),
    .X(net52));
 sg13g2_tielo _1208__53 (.L_LO(net53));
 sg13g2_tielo _1209__54 (.L_LO(net54));
 sg13g2_tielo _1210__55 (.L_LO(net55));
 sg13g2_tielo _1211__56 (.L_LO(net56));
 sg13g2_tielo _1212__57 (.L_LO(net57));
 sg13g2_tielo _1213__58 (.L_LO(net58));
 sg13g2_tielo _1214__59 (.L_LO(net59));
 sg13g2_tielo _1215__60 (.L_LO(net60));
 sg13g2_tielo _1216__61 (.L_LO(net61));
 sg13g2_tielo _1217__62 (.L_LO(net62));
 sg13g2_tielo _1218__63 (.L_LO(net63));
 sg13g2_tielo _1219__64 (.L_LO(net64));
 sg13g2_tielo _1220__65 (.L_LO(net65));
 sg13g2_tielo _1221__66 (.L_LO(net66));
 sg13g2_tielo _1222__67 (.L_LO(net67));
 sg13g2_tielo _1223__68 (.L_LO(net68));
 sg13g2_tielo _1225__69 (.L_LO(net69));
 sg13g2_tielo _1226__70 (.L_LO(net70));
 sg13g2_tielo _1227__71 (.L_LO(net71));
 sg13g2_tielo _1228__72 (.L_LO(net72));
 sg13g2_tielo _1229__73 (.L_LO(net73));
 sg13g2_tielo _1230__74 (.L_LO(net74));
 sg13g2_tielo _1231__75 (.L_LO(net75));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_266 ();
 sg13g2_fill_1 FILLER_13_268 ();
 sg13g2_decap_8 FILLER_13_295 ();
 sg13g2_decap_8 FILLER_13_302 ();
 sg13g2_decap_8 FILLER_13_309 ();
 sg13g2_decap_8 FILLER_13_316 ();
 sg13g2_decap_4 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_327 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_fill_1 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_360 ();
 sg13g2_decap_8 FILLER_13_367 ();
 sg13g2_decap_8 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_fill_2 FILLER_13_388 ();
 sg13g2_decap_8 FILLER_13_416 ();
 sg13g2_decap_8 FILLER_13_423 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_152 ();
 sg13g2_decap_8 FILLER_14_159 ();
 sg13g2_decap_8 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_173 ();
 sg13g2_decap_8 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_decap_8 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_fill_2 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_fill_1 FILLER_14_279 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_fill_2 FILLER_14_299 ();
 sg13g2_fill_2 FILLER_14_344 ();
 sg13g2_fill_1 FILLER_14_346 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_4 FILLER_14_378 ();
 sg13g2_fill_1 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_8 FILLER_14_404 ();
 sg13g2_decap_8 FILLER_14_411 ();
 sg13g2_decap_8 FILLER_14_418 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_decap_8 FILLER_15_142 ();
 sg13g2_decap_4 FILLER_15_149 ();
 sg13g2_fill_2 FILLER_15_153 ();
 sg13g2_decap_8 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_188 ();
 sg13g2_decap_8 FILLER_15_195 ();
 sg13g2_decap_8 FILLER_15_202 ();
 sg13g2_decap_8 FILLER_15_209 ();
 sg13g2_decap_4 FILLER_15_251 ();
 sg13g2_decap_4 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_276 ();
 sg13g2_decap_8 FILLER_15_318 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_fill_1 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_4 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_4 FILLER_16_84 ();
 sg13g2_decap_4 FILLER_16_118 ();
 sg13g2_fill_2 FILLER_16_122 ();
 sg13g2_decap_8 FILLER_16_136 ();
 sg13g2_fill_2 FILLER_16_143 ();
 sg13g2_fill_1 FILLER_16_145 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_163 ();
 sg13g2_fill_2 FILLER_16_195 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_230 ();
 sg13g2_fill_2 FILLER_16_237 ();
 sg13g2_fill_1 FILLER_16_254 ();
 sg13g2_fill_2 FILLER_16_261 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_fill_1 FILLER_16_281 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_fill_1 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_fill_2 FILLER_16_314 ();
 sg13g2_fill_1 FILLER_16_320 ();
 sg13g2_fill_1 FILLER_16_342 ();
 sg13g2_fill_2 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_4 FILLER_16_377 ();
 sg13g2_fill_1 FILLER_16_396 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_4 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_88 ();
 sg13g2_decap_4 FILLER_17_115 ();
 sg13g2_fill_2 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_131 ();
 sg13g2_decap_8 FILLER_17_138 ();
 sg13g2_decap_8 FILLER_17_145 ();
 sg13g2_fill_2 FILLER_17_158 ();
 sg13g2_fill_1 FILLER_17_160 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_decap_8 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_190 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_decap_8 FILLER_17_211 ();
 sg13g2_fill_2 FILLER_17_218 ();
 sg13g2_fill_1 FILLER_17_220 ();
 sg13g2_decap_8 FILLER_17_261 ();
 sg13g2_fill_1 FILLER_17_268 ();
 sg13g2_fill_1 FILLER_17_274 ();
 sg13g2_decap_4 FILLER_17_285 ();
 sg13g2_fill_1 FILLER_17_289 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_332 ();
 sg13g2_decap_4 FILLER_17_339 ();
 sg13g2_fill_1 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_fill_2 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_403 ();
 sg13g2_decap_8 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_4 FILLER_17_424 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_4 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_fill_2 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_120 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_decap_8 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_fill_2 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_226 ();
 sg13g2_decap_8 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_4 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_fill_2 FILLER_18_294 ();
 sg13g2_fill_1 FILLER_18_296 ();
 sg13g2_fill_1 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_1 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_366 ();
 sg13g2_fill_1 FILLER_18_368 ();
 sg13g2_decap_4 FILLER_18_379 ();
 sg13g2_fill_2 FILLER_18_383 ();
 sg13g2_decap_4 FILLER_18_398 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_fill_1 FILLER_19_89 ();
 sg13g2_fill_2 FILLER_19_99 ();
 sg13g2_fill_2 FILLER_19_108 ();
 sg13g2_fill_1 FILLER_19_110 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_fill_2 FILLER_19_158 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_decap_4 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_decap_8 FILLER_19_276 ();
 sg13g2_decap_8 FILLER_19_283 ();
 sg13g2_decap_4 FILLER_19_290 ();
 sg13g2_fill_1 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_299 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_fill_2 FILLER_19_327 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_fill_2 FILLER_19_337 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_fill_1 FILLER_19_351 ();
 sg13g2_fill_2 FILLER_19_360 ();
 sg13g2_fill_1 FILLER_19_367 ();
 sg13g2_fill_2 FILLER_19_372 ();
 sg13g2_fill_1 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_fill_2 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_423 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_fill_2 FILLER_20_63 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_decap_8 FILLER_20_117 ();
 sg13g2_decap_8 FILLER_20_124 ();
 sg13g2_fill_2 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_4 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_decap_8 FILLER_20_215 ();
 sg13g2_decap_8 FILLER_20_222 ();
 sg13g2_decap_8 FILLER_20_229 ();
 sg13g2_decap_4 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_240 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_fill_2 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_304 ();
 sg13g2_decap_4 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_337 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_4 FILLER_20_355 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_369 ();
 sg13g2_decap_4 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_411 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_decap_4 FILLER_20_425 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_4 FILLER_21_84 ();
 sg13g2_fill_1 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_106 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_fill_2 FILLER_21_162 ();
 sg13g2_fill_2 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_227 ();
 sg13g2_fill_2 FILLER_21_254 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_4 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_fill_2 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_4 FILLER_21_345 ();
 sg13g2_fill_2 FILLER_21_349 ();
 sg13g2_decap_8 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_416 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_86 ();
 sg13g2_decap_4 FILLER_22_145 ();
 sg13g2_decap_8 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_decap_4 FILLER_22_194 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_decap_4 FILLER_22_216 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_decap_8 FILLER_22_229 ();
 sg13g2_decap_8 FILLER_22_236 ();
 sg13g2_fill_2 FILLER_22_243 ();
 sg13g2_fill_1 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_267 ();
 sg13g2_fill_1 FILLER_22_274 ();
 sg13g2_decap_4 FILLER_22_293 ();
 sg13g2_fill_2 FILLER_22_297 ();
 sg13g2_decap_4 FILLER_22_304 ();
 sg13g2_fill_1 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_fill_1 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_fill_2 FILLER_22_384 ();
 sg13g2_fill_2 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_fill_1 FILLER_23_63 ();
 sg13g2_decap_4 FILLER_23_90 ();
 sg13g2_decap_4 FILLER_23_120 ();
 sg13g2_decap_8 FILLER_23_129 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_decap_8 FILLER_23_142 ();
 sg13g2_decap_4 FILLER_23_149 ();
 sg13g2_fill_1 FILLER_23_153 ();
 sg13g2_decap_4 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_4 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_242 ();
 sg13g2_decap_4 FILLER_23_250 ();
 sg13g2_fill_1 FILLER_23_254 ();
 sg13g2_decap_4 FILLER_23_263 ();
 sg13g2_fill_2 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_355 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_404 ();
 sg13g2_decap_8 FILLER_23_411 ();
 sg13g2_decap_8 FILLER_23_418 ();
 sg13g2_decap_4 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_4 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_101 ();
 sg13g2_decap_8 FILLER_24_108 ();
 sg13g2_decap_4 FILLER_24_115 ();
 sg13g2_decap_8 FILLER_24_127 ();
 sg13g2_decap_8 FILLER_24_134 ();
 sg13g2_decap_8 FILLER_24_141 ();
 sg13g2_decap_8 FILLER_24_148 ();
 sg13g2_decap_8 FILLER_24_155 ();
 sg13g2_decap_8 FILLER_24_162 ();
 sg13g2_decap_8 FILLER_24_169 ();
 sg13g2_decap_4 FILLER_24_176 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_decap_8 FILLER_24_230 ();
 sg13g2_decap_4 FILLER_24_237 ();
 sg13g2_decap_8 FILLER_24_267 ();
 sg13g2_decap_4 FILLER_24_274 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_decap_4 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_302 ();
 sg13g2_fill_2 FILLER_24_309 ();
 sg13g2_fill_1 FILLER_24_311 ();
 sg13g2_fill_1 FILLER_24_321 ();
 sg13g2_decap_4 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_337 ();
 sg13g2_fill_2 FILLER_24_344 ();
 sg13g2_fill_1 FILLER_24_346 ();
 sg13g2_fill_1 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_383 ();
 sg13g2_fill_2 FILLER_24_392 ();
 sg13g2_fill_2 FILLER_24_398 ();
 sg13g2_fill_1 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_65 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_decap_8 FILLER_25_104 ();
 sg13g2_decap_8 FILLER_25_111 ();
 sg13g2_fill_1 FILLER_25_118 ();
 sg13g2_decap_8 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_decap_8 FILLER_25_205 ();
 sg13g2_decap_4 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_222 ();
 sg13g2_decap_4 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_240 ();
 sg13g2_decap_4 FILLER_25_251 ();
 sg13g2_decap_4 FILLER_25_260 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_fill_2 FILLER_25_309 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_1 FILLER_25_383 ();
 sg13g2_fill_1 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_4 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_49 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_83 ();
 sg13g2_fill_2 FILLER_26_96 ();
 sg13g2_fill_1 FILLER_26_98 ();
 sg13g2_fill_2 FILLER_26_125 ();
 sg13g2_fill_1 FILLER_26_127 ();
 sg13g2_fill_1 FILLER_26_158 ();
 sg13g2_fill_2 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_fill_1 FILLER_26_227 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_253 ();
 sg13g2_decap_8 FILLER_26_260 ();
 sg13g2_decap_4 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_271 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_fill_1 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_334 ();
 sg13g2_fill_2 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_347 ();
 sg13g2_decap_4 FILLER_26_354 ();
 sg13g2_fill_2 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_decap_8 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_26_415 ();
 sg13g2_decap_8 FILLER_26_422 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_decap_8 FILLER_27_97 ();
 sg13g2_fill_2 FILLER_27_104 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_121 ();
 sg13g2_fill_1 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_137 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_225 ();
 sg13g2_decap_8 FILLER_27_232 ();
 sg13g2_decap_4 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_283 ();
 sg13g2_fill_2 FILLER_27_307 ();
 sg13g2_decap_8 FILLER_27_314 ();
 sg13g2_decap_4 FILLER_27_321 ();
 sg13g2_fill_2 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_decap_8 FILLER_27_383 ();
 sg13g2_fill_2 FILLER_27_390 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_2 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_27_410 ();
 sg13g2_decap_8 FILLER_27_416 ();
 sg13g2_decap_8 FILLER_27_423 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_fill_2 FILLER_28_78 ();
 sg13g2_fill_1 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_120 ();
 sg13g2_fill_2 FILLER_28_134 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_decap_8 FILLER_28_163 ();
 sg13g2_decap_8 FILLER_28_170 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_decap_4 FILLER_28_183 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_201 ();
 sg13g2_fill_2 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_fill_2 FILLER_28_229 ();
 sg13g2_fill_2 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_286 ();
 sg13g2_decap_4 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_decap_8 FILLER_28_316 ();
 sg13g2_decap_8 FILLER_28_323 ();
 sg13g2_decap_4 FILLER_28_330 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_fill_1 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_361 ();
 sg13g2_fill_2 FILLER_28_368 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_4 FILLER_28_393 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_107 ();
 sg13g2_fill_2 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_116 ();
 sg13g2_decap_8 FILLER_29_122 ();
 sg13g2_decap_8 FILLER_29_139 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_decap_8 FILLER_29_153 ();
 sg13g2_decap_4 FILLER_29_160 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_decap_8 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_fill_2 FILLER_29_225 ();
 sg13g2_fill_1 FILLER_29_227 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_fill_2 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_251 ();
 sg13g2_decap_4 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_277 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_312 ();
 sg13g2_decap_4 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_344 ();
 sg13g2_fill_1 FILLER_29_360 ();
 sg13g2_fill_1 FILLER_29_366 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_412 ();
 sg13g2_decap_8 FILLER_29_422 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_4 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_72 ();
 sg13g2_fill_1 FILLER_30_79 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_decap_8 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_160 ();
 sg13g2_decap_8 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_30_206 ();
 sg13g2_fill_1 FILLER_30_208 ();
 sg13g2_decap_8 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_decap_4 FILLER_30_239 ();
 sg13g2_fill_2 FILLER_30_243 ();
 sg13g2_decap_8 FILLER_30_271 ();
 sg13g2_decap_8 FILLER_30_278 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_decap_8 FILLER_30_292 ();
 sg13g2_decap_4 FILLER_30_299 ();
 sg13g2_fill_2 FILLER_30_303 ();
 sg13g2_decap_8 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_337 ();
 sg13g2_fill_2 FILLER_30_348 ();
 sg13g2_fill_1 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_30_373 ();
 sg13g2_fill_2 FILLER_30_380 ();
 sg13g2_fill_2 FILLER_30_388 ();
 sg13g2_fill_2 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_425 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_4 FILLER_31_63 ();
 sg13g2_fill_1 FILLER_31_67 ();
 sg13g2_decap_4 FILLER_31_73 ();
 sg13g2_decap_8 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_89 ();
 sg13g2_decap_8 FILLER_31_96 ();
 sg13g2_decap_8 FILLER_31_103 ();
 sg13g2_decap_8 FILLER_31_110 ();
 sg13g2_decap_4 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_121 ();
 sg13g2_decap_4 FILLER_31_153 ();
 sg13g2_fill_1 FILLER_31_157 ();
 sg13g2_decap_4 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_172 ();
 sg13g2_decap_8 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_fill_2 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_fill_2 FILLER_31_231 ();
 sg13g2_fill_2 FILLER_31_270 ();
 sg13g2_decap_8 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_decap_4 FILLER_31_293 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_fill_1 FILLER_31_326 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_357 ();
 sg13g2_decap_4 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_fill_1 FILLER_31_380 ();
 sg13g2_decap_4 FILLER_31_386 ();
 sg13g2_fill_1 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_decap_8 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_31_414 ();
 sg13g2_decap_8 FILLER_31_421 ();
 sg13g2_fill_2 FILLER_31_428 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_4 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_46 ();
 sg13g2_fill_1 FILLER_32_74 ();
 sg13g2_fill_2 FILLER_32_107 ();
 sg13g2_fill_1 FILLER_32_124 ();
 sg13g2_decap_8 FILLER_32_134 ();
 sg13g2_decap_8 FILLER_32_141 ();
 sg13g2_fill_2 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_171 ();
 sg13g2_fill_2 FILLER_32_178 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_decap_4 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_212 ();
 sg13g2_fill_1 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_decap_8 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_fill_2 FILLER_32_244 ();
 sg13g2_decap_4 FILLER_32_252 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_269 ();
 sg13g2_decap_4 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_304 ();
 sg13g2_decap_8 FILLER_32_311 ();
 sg13g2_decap_4 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_fill_1 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_fill_1 FILLER_32_355 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_401 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_4 FILLER_33_56 ();
 sg13g2_fill_2 FILLER_33_60 ();
 sg13g2_decap_4 FILLER_33_93 ();
 sg13g2_fill_2 FILLER_33_97 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_fill_1 FILLER_33_106 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_4 FILLER_33_161 ();
 sg13g2_fill_2 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_decap_4 FILLER_33_188 ();
 sg13g2_fill_1 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_215 ();
 sg13g2_decap_4 FILLER_33_222 ();
 sg13g2_fill_1 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_239 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_decap_4 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_275 ();
 sg13g2_fill_1 FILLER_33_287 ();
 sg13g2_fill_1 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_315 ();
 sg13g2_fill_2 FILLER_33_321 ();
 sg13g2_decap_8 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_360 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_decap_4 FILLER_33_426 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_123 ();
 sg13g2_fill_2 FILLER_34_130 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_4 FILLER_34_182 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_decap_8 FILLER_34_215 ();
 sg13g2_decap_8 FILLER_34_222 ();
 sg13g2_decap_4 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_265 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_decap_8 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_decap_4 FILLER_34_299 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_1 FILLER_34_324 ();
 sg13g2_decap_4 FILLER_34_347 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_372 ();
 sg13g2_fill_2 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_416 ();
 sg13g2_decap_8 FILLER_34_423 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_84 ();
 sg13g2_decap_4 FILLER_35_122 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_153 ();
 sg13g2_decap_4 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_1 FILLER_35_211 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_4 FILLER_35_224 ();
 sg13g2_decap_4 FILLER_35_246 ();
 sg13g2_decap_8 FILLER_35_262 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_decap_8 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_decap_4 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_2 FILLER_35_319 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_decap_4 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_fill_2 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_fill_1 FILLER_35_409 ();
 sg13g2_decap_8 FILLER_35_423 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_4 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_185 ();
 sg13g2_decap_8 FILLER_36_192 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_fill_2 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_224 ();
 sg13g2_decap_4 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_234 ();
 sg13g2_decap_8 FILLER_36_240 ();
 sg13g2_decap_4 FILLER_36_247 ();
 sg13g2_fill_1 FILLER_36_251 ();
 sg13g2_decap_4 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_267 ();
 sg13g2_decap_8 FILLER_36_274 ();
 sg13g2_decap_4 FILLER_36_281 ();
 sg13g2_fill_2 FILLER_36_300 ();
 sg13g2_decap_4 FILLER_36_312 ();
 sg13g2_fill_1 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_372 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_decap_4 FILLER_36_386 ();
 sg13g2_fill_2 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_160 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_decap_8 FILLER_37_218 ();
 sg13g2_decap_8 FILLER_37_225 ();
 sg13g2_decap_4 FILLER_37_232 ();
 sg13g2_fill_2 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_decap_8 FILLER_37_309 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_decap_8 FILLER_37_323 ();
 sg13g2_fill_2 FILLER_37_330 ();
 sg13g2_fill_1 FILLER_37_332 ();
 sg13g2_decap_8 FILLER_37_338 ();
 sg13g2_decap_4 FILLER_37_345 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_4 FILLER_37_375 ();
 sg13g2_fill_1 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_410 ();
 sg13g2_fill_1 FILLER_37_417 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_4 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_decap_4 FILLER_38_345 ();
 sg13g2_decap_8 FILLER_38_353 ();
 sg13g2_fill_2 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_362 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_decap_8 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_38_415 ();
 sg13g2_decap_8 FILLER_38_422 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
