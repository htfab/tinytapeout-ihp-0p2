module tt_um_tomkeddie_b (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire clknet_0_clk;
 wire net35;
 wire tx_pin0;
 wire tx_pin1;
 wire tx_pin2;
 wire tx_pin3;
 wire tx_pin4;
 wire \uart_tx.bit_counter[0] ;
 wire \uart_tx.bit_counter[1] ;
 wire \uart_tx.bit_counter[2] ;
 wire \uart_tx.bit_counter[3] ;
 wire \uart_tx.text_index[0] ;
 wire \uart_tx.text_index[1] ;
 wire \uart_tx.text_index[2] ;
 wire \uart_tx.text_index[3] ;
 wire \uart_tx.text_index[4] ;
 wire \uart_tx.text_index[5] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_buf_2 _0567_ (.A(\uart_tx.bit_counter[2] ),
    .X(_0206_));
 sg13g2_inv_1 _0568_ (.Y(_0217_),
    .A(_0206_));
 sg13g2_nand2_1 _0569_ (.Y(_0228_),
    .A(_0217_),
    .B(\uart_tx.bit_counter[3] ));
 sg13g2_buf_2 _0570_ (.A(\uart_tx.bit_counter[0] ),
    .X(_0239_));
 sg13g2_buf_2 _0571_ (.A(\uart_tx.bit_counter[1] ),
    .X(_0250_));
 sg13g2_inv_2 _0572_ (.Y(_0261_),
    .A(_0250_));
 sg13g2_nor2_1 _0573_ (.A(_0239_),
    .B(_0261_),
    .Y(_0272_));
 sg13g2_nor2b_1 _0574_ (.A(_0228_),
    .B_N(_0272_),
    .Y(_0283_));
 sg13g2_inv_1 _0575_ (.Y(_0294_),
    .A(_0283_));
 sg13g2_nand2_2 _0576_ (.Y(_0305_),
    .A(_0294_),
    .B(net1));
 sg13g2_nor2b_1 _0577_ (.A(_0305_),
    .B_N(_0001_),
    .Y(_0002_));
 sg13g2_buf_1 _0578_ (.A(_0239_),
    .X(_0325_));
 sg13g2_nand2_1 _0579_ (.Y(_0336_),
    .A(_0250_),
    .B(net14));
 sg13g2_inv_1 _0580_ (.Y(_0347_),
    .A(_0336_));
 sg13g2_nor2_2 _0581_ (.A(_0250_),
    .B(_0239_),
    .Y(_0358_));
 sg13g2_nor3_1 _0582_ (.A(_0347_),
    .B(_0358_),
    .C(_0305_),
    .Y(_0003_));
 sg13g2_inv_1 _0583_ (.Y(_0379_),
    .A(_0239_));
 sg13g2_buf_1 _0584_ (.A(_0379_),
    .X(_0390_));
 sg13g2_nand2_1 _0585_ (.Y(_0401_),
    .A(_0250_),
    .B(_0206_));
 sg13g2_nor2_1 _0586_ (.A(net13),
    .B(_0401_),
    .Y(_0411_));
 sg13g2_nor2_1 _0587_ (.A(_0206_),
    .B(_0347_),
    .Y(_0422_));
 sg13g2_nor3_1 _0588_ (.A(_0411_),
    .B(_0422_),
    .C(_0305_),
    .Y(_0004_));
 sg13g2_inv_1 _0589_ (.Y(_0443_),
    .A(\uart_tx.bit_counter[3] ));
 sg13g2_nand2_1 _0590_ (.Y(_0454_),
    .A(_0411_),
    .B(_0443_));
 sg13g2_o21ai_1 _0591_ (.B1(\uart_tx.bit_counter[3] ),
    .Y(_0465_),
    .A1(net13),
    .A2(_0401_));
 sg13g2_a21oi_1 _0592_ (.A1(_0454_),
    .A2(_0465_),
    .Y(_0005_),
    .B1(_0305_));
 sg13g2_buf_8 _0593_ (.A(\uart_tx.text_index[0] ),
    .X(_0485_));
 sg13g2_inv_4 _0594_ (.A(_0485_),
    .Y(_0496_));
 sg13g2_nand2_1 _0595_ (.Y(_0507_),
    .A(_0283_),
    .B(_0485_));
 sg13g2_nand2_1 _0596_ (.Y(_0516_),
    .A(_0507_),
    .B(net1));
 sg13g2_a21oi_1 _0597_ (.A1(_0496_),
    .A2(_0294_),
    .Y(_0006_),
    .B1(_0516_));
 sg13g2_buf_8 _0598_ (.A(\uart_tx.text_index[1] ),
    .X(_0517_));
 sg13g2_inv_4 _0599_ (.A(_0517_),
    .Y(_0518_));
 sg13g2_nor2_1 _0600_ (.A(_0518_),
    .B(_0507_),
    .Y(_0519_));
 sg13g2_a21oi_1 _0601_ (.A1(_0283_),
    .A2(_0485_),
    .Y(_0520_),
    .B1(_0517_));
 sg13g2_buf_8 _0602_ (.A(\uart_tx.text_index[4] ),
    .X(_0521_));
 sg13g2_buf_8 _0603_ (.A(\uart_tx.text_index[5] ),
    .X(_0522_));
 sg13g2_nand2_1 _0604_ (.Y(_0523_),
    .A(_0521_),
    .B(net15));
 sg13g2_nor2_2 _0605_ (.A(_0517_),
    .B(_0496_),
    .Y(_0524_));
 sg13g2_buf_8 _0606_ (.A(\uart_tx.text_index[2] ),
    .X(_0525_));
 sg13g2_buf_8 _0607_ (.A(\uart_tx.text_index[3] ),
    .X(_0526_));
 sg13g2_nor2_1 _0608_ (.A(_0525_),
    .B(_0526_),
    .Y(_0527_));
 sg13g2_buf_8 _0609_ (.A(_0527_),
    .X(_0528_));
 sg13g2_nand2_1 _0610_ (.Y(_0529_),
    .A(_0524_),
    .B(net12));
 sg13g2_nor2_1 _0611_ (.A(_0523_),
    .B(_0529_),
    .Y(_0530_));
 sg13g2_inv_1 _0612_ (.Y(_0531_),
    .A(_0530_));
 sg13g2_o21ai_1 _0613_ (.B1(net1),
    .Y(_0532_),
    .A1(_0294_),
    .A2(_0531_));
 sg13g2_nor3_1 _0614_ (.A(_0519_),
    .B(_0520_),
    .C(_0532_),
    .Y(_0007_));
 sg13g2_inv_4 _0615_ (.A(_0525_),
    .Y(_0533_));
 sg13g2_nand2_2 _0616_ (.Y(_0534_),
    .A(_0485_),
    .B(_0517_));
 sg13g2_nor2_1 _0617_ (.A(_0533_),
    .B(_0534_),
    .Y(_0535_));
 sg13g2_nand2_1 _0618_ (.Y(_0536_),
    .A(_0283_),
    .B(_0535_));
 sg13g2_inv_1 _0619_ (.Y(_0537_),
    .A(_0536_));
 sg13g2_nor2_1 _0620_ (.A(_0525_),
    .B(_0519_),
    .Y(_0538_));
 sg13g2_nor3_1 _0621_ (.A(_0537_),
    .B(_0532_),
    .C(_0538_),
    .Y(_0008_));
 sg13g2_nor2_1 _0622_ (.A(_0526_),
    .B(_0537_),
    .Y(_0539_));
 sg13g2_inv_4 _0623_ (.A(_0526_),
    .Y(_0540_));
 sg13g2_nor2_1 _0624_ (.A(_0540_),
    .B(_0536_),
    .Y(_0541_));
 sg13g2_nor3_1 _0625_ (.A(_0539_),
    .B(_0541_),
    .C(_0532_),
    .Y(_0009_));
 sg13g2_nor2_1 _0626_ (.A(_0521_),
    .B(_0541_),
    .Y(_0542_));
 sg13g2_nand2_1 _0627_ (.Y(_0543_),
    .A(_0541_),
    .B(_0521_));
 sg13g2_inv_1 _0628_ (.Y(_0544_),
    .A(_0543_));
 sg13g2_nor3_1 _0629_ (.A(_0532_),
    .B(_0542_),
    .C(_0544_),
    .Y(_0010_));
 sg13g2_inv_2 _0630_ (.Y(_0545_),
    .A(net15));
 sg13g2_nor2_1 _0631_ (.A(_0545_),
    .B(_0543_),
    .Y(_0546_));
 sg13g2_nor2_1 _0632_ (.A(net15),
    .B(_0544_),
    .Y(_0547_));
 sg13g2_nor3_1 _0633_ (.A(_0532_),
    .B(_0546_),
    .C(_0547_),
    .Y(_0011_));
 sg13g2_nor2_2 _0634_ (.A(_0521_),
    .B(net15),
    .Y(_0548_));
 sg13g2_inv_2 _0635_ (.Y(_0549_),
    .A(_0548_));
 sg13g2_nor2_2 _0636_ (.A(_0525_),
    .B(_0540_),
    .Y(_0550_));
 sg13g2_nand2_1 _0637_ (.Y(_0551_),
    .A(_0524_),
    .B(_0550_));
 sg13g2_nor2_1 _0638_ (.A(_0549_),
    .B(_0551_),
    .Y(_0017_));
 sg13g2_nor2_2 _0639_ (.A(_0526_),
    .B(_0533_),
    .Y(_0018_));
 sg13g2_nand2_1 _0640_ (.Y(_0019_),
    .A(_0524_),
    .B(_0018_));
 sg13g2_nor2_1 _0641_ (.A(_0549_),
    .B(_0019_),
    .Y(_0020_));
 sg13g2_nor2_1 _0642_ (.A(_0017_),
    .B(_0020_),
    .Y(_0021_));
 sg13g2_inv_2 _0643_ (.Y(_0022_),
    .A(_0534_));
 sg13g2_buf_8 _0644_ (.A(_0548_),
    .X(_0023_));
 sg13g2_nand3_1 _0645_ (.B(net12),
    .C(net11),
    .A(_0022_),
    .Y(_0024_));
 sg13g2_buf_2 _0646_ (.A(_0024_),
    .X(_0025_));
 sg13g2_nand2_1 _0647_ (.Y(_0026_),
    .A(_0021_),
    .B(_0025_));
 sg13g2_nand2_2 _0648_ (.Y(_0027_),
    .A(_0525_),
    .B(_0526_));
 sg13g2_nand2_2 _0649_ (.Y(_0028_),
    .A(_0496_),
    .B(_0517_));
 sg13g2_nor2_1 _0650_ (.A(_0027_),
    .B(_0028_),
    .Y(_0029_));
 sg13g2_inv_8 _0651_ (.Y(_0030_),
    .A(_0521_));
 sg13g2_nor2_2 _0652_ (.A(_0522_),
    .B(_0030_),
    .Y(_0031_));
 sg13g2_nand2_1 _0653_ (.Y(_0032_),
    .A(_0029_),
    .B(_0031_));
 sg13g2_nor2_2 _0654_ (.A(_0534_),
    .B(_0027_),
    .Y(_0033_));
 sg13g2_buf_8 _0655_ (.A(_0031_),
    .X(_0034_));
 sg13g2_nand2_1 _0656_ (.Y(_0035_),
    .A(_0033_),
    .B(net9));
 sg13g2_nand2_1 _0657_ (.Y(_0036_),
    .A(_0032_),
    .B(_0035_));
 sg13g2_nor2_2 _0658_ (.A(_0549_),
    .B(_0529_),
    .Y(_0037_));
 sg13g2_nor2_2 _0659_ (.A(_0521_),
    .B(_0545_),
    .Y(_0038_));
 sg13g2_nand2_2 _0660_ (.Y(_0039_),
    .A(_0038_),
    .B(net12));
 sg13g2_nor2_1 _0661_ (.A(_0534_),
    .B(_0039_),
    .Y(_0040_));
 sg13g2_nor2_1 _0662_ (.A(_0037_),
    .B(_0040_),
    .Y(_0041_));
 sg13g2_nand2b_1 _0663_ (.Y(_0042_),
    .B(_0041_),
    .A_N(_0036_));
 sg13g2_nor2_1 _0664_ (.A(_0026_),
    .B(_0042_),
    .Y(_0043_));
 sg13g2_nand2_1 _0665_ (.Y(_0044_),
    .A(_0518_),
    .B(_0485_));
 sg13g2_nand2_1 _0666_ (.Y(_0045_),
    .A(_0540_),
    .B(_0525_));
 sg13g2_nor2_1 _0667_ (.A(_0044_),
    .B(_0045_),
    .Y(_0046_));
 sg13g2_nand2_2 _0668_ (.Y(_0047_),
    .A(_0046_),
    .B(net9));
 sg13g2_nor2_1 _0669_ (.A(_0027_),
    .B(_0044_),
    .Y(_0048_));
 sg13g2_nand2_1 _0670_ (.Y(_0049_),
    .A(_0048_),
    .B(net9));
 sg13g2_nand2_1 _0671_ (.Y(_0050_),
    .A(_0047_),
    .B(_0049_));
 sg13g2_inv_1 _0672_ (.Y(_0051_),
    .A(_0027_));
 sg13g2_nor2_1 _0673_ (.A(_0485_),
    .B(_0517_),
    .Y(_0052_));
 sg13g2_buf_8 _0674_ (.A(_0052_),
    .X(_0053_));
 sg13g2_nand3_1 _0675_ (.B(net11),
    .C(net10),
    .A(_0051_),
    .Y(_0054_));
 sg13g2_nand3_1 _0676_ (.B(_0548_),
    .C(net10),
    .A(_0550_),
    .Y(_0055_));
 sg13g2_buf_2 _0677_ (.A(_0055_),
    .X(_0056_));
 sg13g2_nand2_1 _0678_ (.Y(_0057_),
    .A(_0054_),
    .B(_0056_));
 sg13g2_nand2_1 _0679_ (.Y(_0058_),
    .A(_0030_),
    .B(net15));
 sg13g2_buf_8 _0680_ (.A(_0058_),
    .X(_0059_));
 sg13g2_nand2_2 _0681_ (.Y(_0060_),
    .A(_0528_),
    .B(net10));
 sg13g2_nor2_2 _0682_ (.A(net8),
    .B(_0060_),
    .Y(_0061_));
 sg13g2_nand2_2 _0683_ (.Y(_0062_),
    .A(_0018_),
    .B(net10));
 sg13g2_nor2_1 _0684_ (.A(net8),
    .B(_0062_),
    .Y(_0063_));
 sg13g2_nand2_2 _0685_ (.Y(_0064_),
    .A(_0022_),
    .B(_0018_));
 sg13g2_nor2_1 _0686_ (.A(_0549_),
    .B(_0064_),
    .Y(_0065_));
 sg13g2_nor3_1 _0687_ (.A(_0061_),
    .B(_0063_),
    .C(_0065_),
    .Y(_0066_));
 sg13g2_nand3b_1 _0688_ (.B(_0528_),
    .C(_0053_),
    .Y(_0067_),
    .A_N(_0523_));
 sg13g2_nand2_1 _0689_ (.Y(_0068_),
    .A(_0066_),
    .B(_0067_));
 sg13g2_nor4_1 _0690_ (.A(net14),
    .B(_0050_),
    .C(_0057_),
    .D(_0068_),
    .Y(_0069_));
 sg13g2_inv_1 _0691_ (.Y(_0070_),
    .A(_0031_));
 sg13g2_nor2_1 _0692_ (.A(_0070_),
    .B(_0064_),
    .Y(_0071_));
 sg13g2_nand3_1 _0693_ (.B(_0031_),
    .C(_0550_),
    .A(_0524_),
    .Y(_0072_));
 sg13g2_nor2_2 _0694_ (.A(_0485_),
    .B(_0518_),
    .Y(_0073_));
 sg13g2_nand3_1 _0695_ (.B(_0031_),
    .C(net12),
    .A(_0073_),
    .Y(_0074_));
 sg13g2_nand2_1 _0696_ (.Y(_0075_),
    .A(_0072_),
    .B(_0074_));
 sg13g2_nor2_1 _0697_ (.A(_0070_),
    .B(_0062_),
    .Y(_0076_));
 sg13g2_inv_1 _0698_ (.Y(_0077_),
    .A(_0076_));
 sg13g2_nand3_1 _0699_ (.B(_0018_),
    .C(net9),
    .A(_0073_),
    .Y(_0078_));
 sg13g2_buf_8 _0700_ (.A(_0078_),
    .X(_0079_));
 sg13g2_nand2_1 _0701_ (.Y(_0080_),
    .A(_0077_),
    .B(_0079_));
 sg13g2_nand3_1 _0702_ (.B(_0049_),
    .C(_0056_),
    .A(_0047_),
    .Y(_0081_));
 sg13g2_inv_1 _0703_ (.Y(_0082_),
    .A(_0081_));
 sg13g2_nand4_1 _0704_ (.B(net14),
    .C(_0531_),
    .A(_0082_),
    .Y(_0083_),
    .D(_0035_));
 sg13g2_nor4_1 _0705_ (.A(_0071_),
    .B(_0075_),
    .C(_0080_),
    .D(_0083_),
    .Y(_0084_));
 sg13g2_nor2_1 _0706_ (.A(_0071_),
    .B(_0075_),
    .Y(_0085_));
 sg13g2_nand3_1 _0707_ (.B(net12),
    .C(net10),
    .A(_0031_),
    .Y(_0086_));
 sg13g2_inv_1 _0708_ (.Y(_0087_),
    .A(_0086_));
 sg13g2_nand3_1 _0709_ (.B(_0550_),
    .C(net10),
    .A(net9),
    .Y(_0088_));
 sg13g2_buf_1 _0710_ (.A(_0088_),
    .X(_0089_));
 sg13g2_nand2_1 _0711_ (.Y(_0090_),
    .A(_0079_),
    .B(_0089_));
 sg13g2_nor2_1 _0712_ (.A(_0087_),
    .B(_0090_),
    .Y(_0091_));
 sg13g2_nor2_1 _0713_ (.A(_0070_),
    .B(_0529_),
    .Y(_0092_));
 sg13g2_nand3_1 _0714_ (.B(_0018_),
    .C(net11),
    .A(_0073_),
    .Y(_0093_));
 sg13g2_inv_2 _0715_ (.Y(_0094_),
    .A(_0093_));
 sg13g2_nor2_1 _0716_ (.A(_0092_),
    .B(_0094_),
    .Y(_0095_));
 sg13g2_nand3_1 _0717_ (.B(_0034_),
    .C(_0550_),
    .A(_0073_),
    .Y(_0096_));
 sg13g2_buf_2 _0718_ (.A(_0096_),
    .X(_0097_));
 sg13g2_nand4_1 _0719_ (.B(_0091_),
    .C(_0095_),
    .A(_0085_),
    .Y(_0098_),
    .D(_0097_));
 sg13g2_nor2_1 _0720_ (.A(_0523_),
    .B(_0060_),
    .Y(_0099_));
 sg13g2_nor2_1 _0721_ (.A(_0099_),
    .B(_0530_),
    .Y(_0100_));
 sg13g2_inv_1 _0722_ (.Y(_0101_),
    .A(_0100_));
 sg13g2_nor2_1 _0723_ (.A(_0076_),
    .B(_0101_),
    .Y(_0102_));
 sg13g2_nor2b_1 _0724_ (.A(_0098_),
    .B_N(_0102_),
    .Y(_0103_));
 sg13g2_inv_1 _0725_ (.Y(_0104_),
    .A(_0062_));
 sg13g2_nand2_1 _0726_ (.Y(_0105_),
    .A(_0104_),
    .B(net11));
 sg13g2_inv_1 _0727_ (.Y(_0106_),
    .A(_0105_));
 sg13g2_nand3_1 _0728_ (.B(_0034_),
    .C(net10),
    .A(_0051_),
    .Y(_0107_));
 sg13g2_buf_2 _0729_ (.A(_0107_),
    .X(_0108_));
 sg13g2_o21ai_1 _0730_ (.B1(_0108_),
    .Y(_0109_),
    .A1(_0549_),
    .A2(_0060_));
 sg13g2_nor3_1 _0731_ (.A(_0106_),
    .B(_0109_),
    .C(_0081_),
    .Y(_0110_));
 sg13g2_a21oi_1 _0732_ (.A1(_0044_),
    .A2(_0028_),
    .Y(_0111_),
    .B1(_0039_));
 sg13g2_nand2_2 _0733_ (.Y(_0112_),
    .A(_0048_),
    .B(_0023_));
 sg13g2_nand2_1 _0734_ (.Y(_0113_),
    .A(_0112_),
    .B(_0054_));
 sg13g2_nand3_1 _0735_ (.B(_0550_),
    .C(net11),
    .A(_0073_),
    .Y(_0114_));
 sg13g2_nand2_2 _0736_ (.Y(_0115_),
    .A(_0029_),
    .B(net11));
 sg13g2_nand2_1 _0737_ (.Y(_0116_),
    .A(_0114_),
    .B(_0115_));
 sg13g2_nor3_1 _0738_ (.A(_0111_),
    .B(_0113_),
    .C(_0116_),
    .Y(_0117_));
 sg13g2_nand3_1 _0739_ (.B(_0043_),
    .C(_0117_),
    .A(_0110_),
    .Y(_0118_));
 sg13g2_inv_2 _0740_ (.Y(_0119_),
    .A(_0118_));
 sg13g2_nand3_1 _0741_ (.B(net9),
    .C(net12),
    .A(_0022_),
    .Y(_0120_));
 sg13g2_inv_2 _0742_ (.Y(_0121_),
    .A(_0120_));
 sg13g2_nand2_1 _0743_ (.Y(_0122_),
    .A(_0533_),
    .B(_0526_));
 sg13g2_nor2_1 _0744_ (.A(_0534_),
    .B(_0122_),
    .Y(_0123_));
 sg13g2_nand2_1 _0745_ (.Y(_0124_),
    .A(_0123_),
    .B(net9));
 sg13g2_inv_1 _0746_ (.Y(_0125_),
    .A(_0124_));
 sg13g2_nand2_2 _0747_ (.Y(_0126_),
    .A(_0123_),
    .B(net11));
 sg13g2_nand2_2 _0748_ (.Y(_0127_),
    .A(_0033_),
    .B(_0023_));
 sg13g2_nand2_1 _0749_ (.Y(_0128_),
    .A(_0126_),
    .B(_0127_));
 sg13g2_nor3_1 _0750_ (.A(_0121_),
    .B(_0125_),
    .C(_0128_),
    .Y(_0129_));
 sg13g2_nor2_1 _0751_ (.A(_0534_),
    .B(_0045_),
    .Y(_0130_));
 sg13g2_nand2_1 _0752_ (.Y(_0131_),
    .A(_0130_),
    .B(_0038_));
 sg13g2_nand3_1 _0753_ (.B(_0038_),
    .C(_0053_),
    .A(_0550_),
    .Y(_0132_));
 sg13g2_nand2_1 _0754_ (.Y(_0133_),
    .A(_0123_),
    .B(_0038_));
 sg13g2_nand3_1 _0755_ (.B(_0132_),
    .C(_0133_),
    .A(_0131_),
    .Y(_0134_));
 sg13g2_inv_1 _0756_ (.Y(_0135_),
    .A(_0134_));
 sg13g2_nand3_1 _0757_ (.B(_0135_),
    .C(_0066_),
    .A(_0129_),
    .Y(_0136_));
 sg13g2_nor2_1 _0758_ (.A(net8),
    .B(_0019_),
    .Y(_0137_));
 sg13g2_nor2_1 _0759_ (.A(net8),
    .B(_0551_),
    .Y(_0138_));
 sg13g2_nor3_1 _0760_ (.A(_0028_),
    .B(_0045_),
    .C(net8),
    .Y(_0139_));
 sg13g2_nor2_1 _0761_ (.A(_0138_),
    .B(_0139_),
    .Y(_0140_));
 sg13g2_nor2_1 _0762_ (.A(_0027_),
    .B(_0058_),
    .Y(_0141_));
 sg13g2_inv_1 _0763_ (.Y(_0142_),
    .A(_0141_));
 sg13g2_nand2_1 _0764_ (.Y(_0143_),
    .A(_0073_),
    .B(_0550_));
 sg13g2_nor2_1 _0765_ (.A(net8),
    .B(_0143_),
    .Y(_0144_));
 sg13g2_inv_1 _0766_ (.Y(_0145_),
    .A(_0144_));
 sg13g2_nand3_1 _0767_ (.B(_0142_),
    .C(_0145_),
    .A(_0140_),
    .Y(_0146_));
 sg13g2_nor2_1 _0768_ (.A(_0137_),
    .B(_0146_),
    .Y(_0147_));
 sg13g2_nor2b_1 _0769_ (.A(_0136_),
    .B_N(_0147_),
    .Y(_0148_));
 sg13g2_nand3_1 _0770_ (.B(_0119_),
    .C(_0148_),
    .A(_0103_),
    .Y(_0149_));
 sg13g2_a22oi_1 _0771_ (.Y(_0150_),
    .B1(_0084_),
    .B2(_0149_),
    .A2(_0069_),
    .A1(_0043_));
 sg13g2_nor2_1 _0772_ (.A(_0206_),
    .B(_0261_),
    .Y(_0151_));
 sg13g2_nor2b_1 _0773_ (.A(_0150_),
    .B_N(_0151_),
    .Y(_0152_));
 sg13g2_nand2_2 _0774_ (.Y(_0153_),
    .A(_0261_),
    .B(_0206_));
 sg13g2_inv_1 _0775_ (.Y(_0154_),
    .A(_0025_));
 sg13g2_nor2_1 _0776_ (.A(_0379_),
    .B(_0154_),
    .Y(_0155_));
 sg13g2_inv_1 _0777_ (.Y(_0156_),
    .A(_0155_));
 sg13g2_nor3_1 _0778_ (.A(_0113_),
    .B(_0156_),
    .C(_0042_),
    .Y(_0157_));
 sg13g2_nor3_1 _0779_ (.A(_0101_),
    .B(_0076_),
    .C(_0081_),
    .Y(_0158_));
 sg13g2_inv_2 _0780_ (.Y(_0159_),
    .A(_0032_));
 sg13g2_inv_1 _0781_ (.Y(_0160_),
    .A(_0114_));
 sg13g2_nor2_1 _0782_ (.A(_0159_),
    .B(_0160_),
    .Y(_0161_));
 sg13g2_inv_1 _0783_ (.Y(_0162_),
    .A(_0111_));
 sg13g2_nand3_1 _0784_ (.B(_0162_),
    .C(_0097_),
    .A(_0161_),
    .Y(_0163_));
 sg13g2_nor2_1 _0785_ (.A(_0106_),
    .B(_0109_),
    .Y(_0164_));
 sg13g2_nand2_1 _0786_ (.Y(_0165_),
    .A(_0164_),
    .B(_0082_));
 sg13g2_nor2_1 _0787_ (.A(_0163_),
    .B(_0165_),
    .Y(_0166_));
 sg13g2_inv_1 _0788_ (.Y(_0167_),
    .A(_0017_));
 sg13g2_nand2_1 _0789_ (.Y(_0168_),
    .A(_0167_),
    .B(_0379_));
 sg13g2_nor3_1 _0790_ (.A(_0080_),
    .B(_0168_),
    .C(_0068_),
    .Y(_0169_));
 sg13g2_a22oi_1 _0791_ (.Y(_0170_),
    .B1(_0166_),
    .B2(_0169_),
    .A2(_0158_),
    .A1(_0157_));
 sg13g2_nor2_1 _0792_ (.A(_0153_),
    .B(_0170_),
    .Y(_0171_));
 sg13g2_inv_1 _0793_ (.Y(_0172_),
    .A(_0358_));
 sg13g2_nand2_1 _0794_ (.Y(_0173_),
    .A(_0261_),
    .B(_0217_));
 sg13g2_nand2_1 _0795_ (.Y(_0174_),
    .A(_0173_),
    .B(_0443_));
 sg13g2_o21ai_1 _0796_ (.B1(_0174_),
    .Y(_0175_),
    .A1(_0228_),
    .A2(_0172_));
 sg13g2_nor2_1 _0797_ (.A(\uart_tx.bit_counter[3] ),
    .B(_0206_),
    .Y(_0176_));
 sg13g2_nand2_1 _0798_ (.Y(_0177_),
    .A(_0176_),
    .B(_0000_));
 sg13g2_nand2_1 _0799_ (.Y(_0178_),
    .A(_0175_),
    .B(_0177_));
 sg13g2_a21oi_1 _0800_ (.A1(_0171_),
    .A2(_0149_),
    .Y(_0179_),
    .B1(_0178_));
 sg13g2_inv_1 _0801_ (.Y(_0180_),
    .A(_0151_));
 sg13g2_nand2_2 _0802_ (.Y(_0181_),
    .A(_0180_),
    .B(_0153_));
 sg13g2_nand4_1 _0803_ (.B(_0167_),
    .C(_0114_),
    .A(_0164_),
    .Y(_0182_),
    .D(_0115_));
 sg13g2_nor3_1 _0804_ (.A(_0181_),
    .B(_0098_),
    .C(_0182_),
    .Y(_0183_));
 sg13g2_nand2_1 _0805_ (.Y(_0184_),
    .A(_0183_),
    .B(_0025_));
 sg13g2_nand2_1 _0806_ (.Y(_0185_),
    .A(_0184_),
    .B(_0149_));
 sg13g2_nand2_1 _0807_ (.Y(_0186_),
    .A(_0185_),
    .B(_0272_));
 sg13g2_nand2_1 _0808_ (.Y(_0187_),
    .A(_0179_),
    .B(_0186_));
 sg13g2_nor2_1 _0809_ (.A(_0152_),
    .B(_0187_),
    .Y(_0188_));
 sg13g2_nand3_1 _0810_ (.B(_0095_),
    .C(_0077_),
    .A(_0066_),
    .Y(_0189_));
 sg13g2_nor2_1 _0811_ (.A(_0189_),
    .B(_0118_),
    .Y(_0190_));
 sg13g2_inv_1 _0812_ (.Y(_0191_),
    .A(_0079_));
 sg13g2_nor2_1 _0813_ (.A(_0250_),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_nand3_1 _0814_ (.B(_0190_),
    .C(_0192_),
    .A(_0149_),
    .Y(_0193_));
 sg13g2_nand2_1 _0815_ (.Y(_0194_),
    .A(_0261_),
    .B(net14));
 sg13g2_nand2_1 _0816_ (.Y(_0195_),
    .A(_0103_),
    .B(_0119_));
 sg13g2_nand4_1 _0817_ (.B(_0041_),
    .C(_0239_),
    .A(_0021_),
    .Y(_0196_),
    .D(_0025_));
 sg13g2_nand3_1 _0818_ (.B(_0162_),
    .C(_0161_),
    .A(_0082_),
    .Y(_0197_));
 sg13g2_nor3_1 _0819_ (.A(_0196_),
    .B(_0197_),
    .C(_0098_),
    .Y(_0198_));
 sg13g2_nand3_1 _0820_ (.B(_0198_),
    .C(_0148_),
    .A(_0195_),
    .Y(_0199_));
 sg13g2_nand3_1 _0821_ (.B(_0194_),
    .C(_0199_),
    .A(_0193_),
    .Y(_0200_));
 sg13g2_inv_2 _0822_ (.Y(_0201_),
    .A(_0181_));
 sg13g2_nand2_1 _0823_ (.Y(_0202_),
    .A(_0200_),
    .B(_0201_));
 sg13g2_nand2_1 _0824_ (.Y(_0203_),
    .A(_0188_),
    .B(_0202_));
 sg13g2_a21oi_2 _0825_ (.B1(_0305_),
    .Y(_0204_),
    .A2(_0176_),
    .A1(_0358_));
 sg13g2_nand2_1 _0826_ (.Y(_0012_),
    .A(_0203_),
    .B(_0204_));
 sg13g2_inv_4 _0827_ (.A(_0056_),
    .Y(_0205_));
 sg13g2_nor2_1 _0828_ (.A(_0037_),
    .B(_0205_),
    .Y(_0207_));
 sg13g2_nand2_1 _0829_ (.Y(_0208_),
    .A(_0207_),
    .B(_0054_));
 sg13g2_inv_1 _0830_ (.Y(_0209_),
    .A(_0115_));
 sg13g2_inv_1 _0831_ (.Y(_0210_),
    .A(_0020_));
 sg13g2_nand2_1 _0832_ (.Y(_0211_),
    .A(_0210_),
    .B(_0127_));
 sg13g2_nor2_1 _0833_ (.A(_0209_),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_nand2b_1 _0834_ (.Y(_0213_),
    .B(_0212_),
    .A_N(_0208_));
 sg13g2_nand2_1 _0835_ (.Y(_0214_),
    .A(_0100_),
    .B(_0108_));
 sg13g2_nand2_1 _0836_ (.Y(_0215_),
    .A(_0130_),
    .B(net11));
 sg13g2_nand3_1 _0837_ (.B(net12),
    .C(_0548_),
    .A(_0073_),
    .Y(_0216_));
 sg13g2_nand3_1 _0838_ (.B(_0215_),
    .C(_0216_),
    .A(_0105_),
    .Y(_0218_));
 sg13g2_nor2_1 _0839_ (.A(_0214_),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_a21oi_1 _0840_ (.A1(_0064_),
    .A2(_0062_),
    .Y(_0220_),
    .B1(_0070_));
 sg13g2_nand3_1 _0841_ (.B(_0097_),
    .C(_0126_),
    .A(_0047_),
    .Y(_0221_));
 sg13g2_nor2_1 _0842_ (.A(_0220_),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_nand2_1 _0843_ (.Y(_0223_),
    .A(_0219_),
    .B(_0222_));
 sg13g2_nor2_1 _0844_ (.A(_0213_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_nand3_1 _0845_ (.B(net9),
    .C(net12),
    .A(_0524_),
    .Y(_0225_));
 sg13g2_nand3_1 _0846_ (.B(_0112_),
    .C(_0035_),
    .A(_0225_),
    .Y(_0226_));
 sg13g2_nand3_1 _0847_ (.B(_0089_),
    .C(_0124_),
    .A(_0079_),
    .Y(_0227_));
 sg13g2_nor2_1 _0848_ (.A(_0226_),
    .B(_0227_),
    .Y(_0229_));
 sg13g2_a21oi_1 _0849_ (.A1(_0019_),
    .A2(_0062_),
    .Y(_0230_),
    .B1(net8));
 sg13g2_nand2_1 _0850_ (.Y(_0231_),
    .A(_0141_),
    .B(_0517_));
 sg13g2_nand3_1 _0851_ (.B(_0231_),
    .C(_0025_),
    .A(_0114_),
    .Y(_0232_));
 sg13g2_nor2_1 _0852_ (.A(_0230_),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_nand2_1 _0853_ (.Y(_0234_),
    .A(_0229_),
    .B(_0233_));
 sg13g2_nor3_1 _0854_ (.A(_0517_),
    .B(_0027_),
    .C(_0059_),
    .Y(_0235_));
 sg13g2_nor2_1 _0855_ (.A(_0235_),
    .B(_0144_),
    .Y(_0236_));
 sg13g2_nand2_1 _0856_ (.Y(_0237_),
    .A(_0140_),
    .B(_0236_));
 sg13g2_nor2_1 _0857_ (.A(_0134_),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_nor2b_1 _0858_ (.A(_0234_),
    .B_N(_0238_),
    .Y(_0240_));
 sg13g2_nand2_1 _0859_ (.Y(_0241_),
    .A(_0093_),
    .B(_0086_));
 sg13g2_nor3_1 _0860_ (.A(_0017_),
    .B(_0159_),
    .C(_0241_),
    .Y(_0242_));
 sg13g2_nand2_1 _0861_ (.Y(_0243_),
    .A(_0242_),
    .B(_0049_));
 sg13g2_nor2_1 _0862_ (.A(_0061_),
    .B(_0075_),
    .Y(_0244_));
 sg13g2_inv_1 _0863_ (.Y(_0245_),
    .A(_0040_));
 sg13g2_nor2_1 _0864_ (.A(_0121_),
    .B(_0111_),
    .Y(_0246_));
 sg13g2_nand3_1 _0865_ (.B(_0245_),
    .C(_0246_),
    .A(_0244_),
    .Y(_0247_));
 sg13g2_nor2_1 _0866_ (.A(_0243_),
    .B(_0247_),
    .Y(_0248_));
 sg13g2_nand3_1 _0867_ (.B(_0240_),
    .C(_0248_),
    .A(_0224_),
    .Y(_0249_));
 sg13g2_buf_1 _0868_ (.A(_0249_),
    .X(_0251_));
 sg13g2_nand2_1 _0869_ (.Y(_0252_),
    .A(_0074_),
    .B(_0120_));
 sg13g2_nor2_1 _0870_ (.A(_0160_),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_nand3_1 _0871_ (.B(_0225_),
    .C(_0126_),
    .A(_0253_),
    .Y(_0254_));
 sg13g2_inv_1 _0872_ (.Y(_0255_),
    .A(_0037_));
 sg13g2_nand3_1 _0873_ (.B(_0077_),
    .C(_0127_),
    .A(_0255_),
    .Y(_0256_));
 sg13g2_nand2_1 _0874_ (.Y(_0257_),
    .A(_0215_),
    .B(_0216_));
 sg13g2_nor2_1 _0875_ (.A(_0209_),
    .B(_0257_),
    .Y(_0258_));
 sg13g2_inv_1 _0876_ (.Y(_0259_),
    .A(_0112_));
 sg13g2_nor2_1 _0877_ (.A(_0017_),
    .B(_0259_),
    .Y(_0260_));
 sg13g2_nand3b_1 _0878_ (.B(_0258_),
    .C(_0260_),
    .Y(_0262_),
    .A_N(_0256_));
 sg13g2_nor2_1 _0879_ (.A(_0254_),
    .B(_0262_),
    .Y(_0263_));
 sg13g2_nand2_1 _0880_ (.Y(_0264_),
    .A(_0210_),
    .B(_0025_));
 sg13g2_nand4_1 _0881_ (.B(_0072_),
    .C(_0097_),
    .A(_0047_),
    .Y(_0265_),
    .D(_0089_));
 sg13g2_nor3_1 _0882_ (.A(_0264_),
    .B(_0094_),
    .C(_0265_),
    .Y(_0266_));
 sg13g2_nand3_1 _0883_ (.B(_0263_),
    .C(_0266_),
    .A(net7),
    .Y(_0267_));
 sg13g2_nand2_1 _0884_ (.Y(_0268_),
    .A(_0267_),
    .B(_0358_));
 sg13g2_nor4_1 _0885_ (.A(_0125_),
    .B(_0106_),
    .C(_0050_),
    .D(_0057_),
    .Y(_0269_));
 sg13g2_nand2_1 _0886_ (.Y(_0270_),
    .A(_0269_),
    .B(_0238_));
 sg13g2_nand4_1 _0887_ (.B(_0079_),
    .C(_0231_),
    .A(_0108_),
    .Y(_0271_),
    .D(_0086_));
 sg13g2_nand3_1 _0888_ (.B(_0093_),
    .C(_0025_),
    .A(_0210_),
    .Y(_0273_));
 sg13g2_nor2_1 _0889_ (.A(_0230_),
    .B(_0273_),
    .Y(_0274_));
 sg13g2_inv_1 _0890_ (.Y(_0275_),
    .A(_0039_));
 sg13g2_nor3_1 _0891_ (.A(_0275_),
    .B(_0071_),
    .C(_0036_),
    .Y(_0276_));
 sg13g2_nand3b_1 _0892_ (.B(_0274_),
    .C(_0276_),
    .Y(_0277_),
    .A_N(_0271_));
 sg13g2_nor2_1 _0893_ (.A(_0270_),
    .B(_0277_),
    .Y(_0278_));
 sg13g2_a21oi_1 _0894_ (.A1(_0278_),
    .A2(_0263_),
    .Y(_0279_),
    .B1(_0336_));
 sg13g2_o21ai_1 _0895_ (.B1(_0167_),
    .Y(_0280_),
    .A1(net15),
    .A2(_0019_));
 sg13g2_o21ai_1 _0896_ (.B1(_0272_),
    .Y(_0281_),
    .A1(_0280_),
    .A2(_0256_));
 sg13g2_nor2b_1 _0897_ (.A(_0279_),
    .B_N(_0281_),
    .Y(_0282_));
 sg13g2_nand2_1 _0898_ (.Y(_0284_),
    .A(_0268_),
    .B(_0282_));
 sg13g2_nand2_1 _0899_ (.Y(_0285_),
    .A(_0284_),
    .B(_0177_));
 sg13g2_nand2_1 _0900_ (.Y(_0286_),
    .A(_0285_),
    .B(_0201_));
 sg13g2_inv_1 _0901_ (.Y(_0287_),
    .A(_0127_));
 sg13g2_nor3_1 _0902_ (.A(_0160_),
    .B(_0287_),
    .C(_0252_),
    .Y(_0288_));
 sg13g2_inv_1 _0903_ (.Y(_0289_),
    .A(_0072_));
 sg13g2_inv_1 _0904_ (.Y(_0290_),
    .A(_0047_));
 sg13g2_nor2_1 _0905_ (.A(_0289_),
    .B(_0290_),
    .Y(_0291_));
 sg13g2_nand2_1 _0906_ (.Y(_0292_),
    .A(_0067_),
    .B(_0379_));
 sg13g2_inv_1 _0907_ (.Y(_0293_),
    .A(_0292_));
 sg13g2_nand4_1 _0908_ (.B(_0258_),
    .C(_0291_),
    .A(_0288_),
    .Y(_0295_),
    .D(_0293_));
 sg13g2_nand2_1 _0909_ (.Y(_0296_),
    .A(_0531_),
    .B(_0239_));
 sg13g2_nor2_1 _0910_ (.A(_0259_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_nor3_1 _0911_ (.A(_0076_),
    .B(_0154_),
    .C(_0290_),
    .Y(_0298_));
 sg13g2_nand3_1 _0912_ (.B(_0298_),
    .C(_0253_),
    .A(_0297_),
    .Y(_0299_));
 sg13g2_a21oi_1 _0913_ (.A1(_0295_),
    .A2(_0299_),
    .Y(_0300_),
    .B1(_0261_));
 sg13g2_nand2_1 _0914_ (.Y(_0301_),
    .A(_0100_),
    .B(_0097_));
 sg13g2_nor4_1 _0915_ (.A(_0090_),
    .B(_0094_),
    .C(_0156_),
    .D(_0301_),
    .Y(_0302_));
 sg13g2_nand2_1 _0916_ (.Y(_0303_),
    .A(_0302_),
    .B(_0288_));
 sg13g2_nand2_1 _0917_ (.Y(_0304_),
    .A(_0079_),
    .B(_0097_));
 sg13g2_nor4_1 _0918_ (.A(_0257_),
    .B(_0292_),
    .C(_0304_),
    .D(_0264_),
    .Y(_0306_));
 sg13g2_nand2b_1 _0919_ (.Y(_0307_),
    .B(_0306_),
    .A_N(_0254_));
 sg13g2_a21oi_1 _0920_ (.A1(_0303_),
    .A2(_0307_),
    .Y(_0308_),
    .B1(_0250_));
 sg13g2_o21ai_1 _0921_ (.B1(net7),
    .Y(_0309_),
    .A1(_0300_),
    .A2(_0308_));
 sg13g2_inv_1 _0922_ (.Y(_0310_),
    .A(_0178_));
 sg13g2_nand2_1 _0923_ (.Y(_0311_),
    .A(_0309_),
    .B(_0310_));
 sg13g2_nand2_1 _0924_ (.Y(_0312_),
    .A(_0175_),
    .B(_0201_));
 sg13g2_nand2_1 _0925_ (.Y(_0313_),
    .A(_0311_),
    .B(_0312_));
 sg13g2_nand2_1 _0926_ (.Y(_0314_),
    .A(_0286_),
    .B(_0313_));
 sg13g2_nand2_1 _0927_ (.Y(_0013_),
    .A(_0314_),
    .B(_0204_));
 sg13g2_nand2_1 _0928_ (.Y(_0315_),
    .A(_0077_),
    .B(_0124_));
 sg13g2_nor2_1 _0929_ (.A(_0315_),
    .B(_0232_),
    .Y(_0316_));
 sg13g2_nor3_1 _0930_ (.A(_0235_),
    .B(_0040_),
    .C(_0087_),
    .Y(_0317_));
 sg13g2_nand2_1 _0931_ (.Y(_0318_),
    .A(_0133_),
    .B(_0127_));
 sg13g2_nand3_1 _0932_ (.B(_0018_),
    .C(_0038_),
    .A(_0073_),
    .Y(_0319_));
 sg13g2_nand2_1 _0933_ (.Y(_0320_),
    .A(_0319_),
    .B(_0049_));
 sg13g2_nor2_1 _0934_ (.A(_0318_),
    .B(_0320_),
    .Y(_0321_));
 sg13g2_nand3_1 _0935_ (.B(_0317_),
    .C(_0321_),
    .A(_0316_),
    .Y(_0322_));
 sg13g2_nand3_1 _0936_ (.B(_0089_),
    .C(_0035_),
    .A(_0047_),
    .Y(_0323_));
 sg13g2_nand2_1 _0937_ (.Y(_0324_),
    .A(_0051_),
    .B(net10));
 sg13g2_nor2_1 _0938_ (.A(_0549_),
    .B(_0324_),
    .Y(_0326_));
 sg13g2_nor2_1 _0939_ (.A(_0326_),
    .B(_0138_),
    .Y(_0327_));
 sg13g2_nor2b_1 _0940_ (.A(_0323_),
    .B_N(_0327_),
    .Y(_0328_));
 sg13g2_nor2_1 _0941_ (.A(_0028_),
    .B(_0039_),
    .Y(_0329_));
 sg13g2_nand3b_1 _0942_ (.B(_0145_),
    .C(_0131_),
    .Y(_0330_),
    .A_N(_0329_));
 sg13g2_inv_1 _0943_ (.Y(_0331_),
    .A(_0330_));
 sg13g2_nand2_1 _0944_ (.Y(_0332_),
    .A(_0046_),
    .B(_0030_));
 sg13g2_and2_1 _0945_ (.A(_0332_),
    .B(_0132_),
    .X(_0333_));
 sg13g2_nand3_1 _0946_ (.B(_0331_),
    .C(_0333_),
    .A(_0328_),
    .Y(_0334_));
 sg13g2_nor2_1 _0947_ (.A(_0322_),
    .B(_0334_),
    .Y(_0335_));
 sg13g2_inv_2 _0948_ (.Y(_0337_),
    .A(_0216_));
 sg13g2_nor2_1 _0949_ (.A(_0337_),
    .B(_0121_),
    .Y(_0338_));
 sg13g2_nand2_1 _0950_ (.Y(_0339_),
    .A(_0338_),
    .B(_0115_));
 sg13g2_nor2_1 _0951_ (.A(_0259_),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_nand2_1 _0952_ (.Y(_0341_),
    .A(_0340_),
    .B(_0126_));
 sg13g2_nor2_1 _0953_ (.A(net15),
    .B(_0064_),
    .Y(_0342_));
 sg13g2_nor2_1 _0954_ (.A(_0342_),
    .B(_0094_),
    .Y(_0343_));
 sg13g2_nand2_1 _0955_ (.Y(_0344_),
    .A(_0343_),
    .B(_0079_));
 sg13g2_inv_1 _0956_ (.Y(_0345_),
    .A(_0344_));
 sg13g2_nand2_1 _0957_ (.Y(_0346_),
    .A(_0072_),
    .B(_0225_));
 sg13g2_nor2_1 _0958_ (.A(_0346_),
    .B(_0109_),
    .Y(_0348_));
 sg13g2_nand2_1 _0959_ (.Y(_0349_),
    .A(_0167_),
    .B(_0056_));
 sg13g2_nor2_1 _0960_ (.A(_0101_),
    .B(_0349_),
    .Y(_0350_));
 sg13g2_nand3_1 _0961_ (.B(_0348_),
    .C(_0350_),
    .A(_0345_),
    .Y(_0351_));
 sg13g2_nor2_1 _0962_ (.A(_0341_),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_nor2_1 _0963_ (.A(_0061_),
    .B(_0159_),
    .Y(_0353_));
 sg13g2_inv_1 _0964_ (.Y(_0354_),
    .A(_0353_));
 sg13g2_inv_1 _0965_ (.Y(_0355_),
    .A(_0063_));
 sg13g2_nand2_1 _0966_ (.Y(_0356_),
    .A(_0355_),
    .B(_0097_));
 sg13g2_inv_1 _0967_ (.Y(_0357_),
    .A(_0074_));
 sg13g2_nor2_1 _0968_ (.A(_0037_),
    .B(_0357_),
    .Y(_0359_));
 sg13g2_nor2_1 _0969_ (.A(_0044_),
    .B(_0039_),
    .Y(_0360_));
 sg13g2_inv_1 _0970_ (.Y(_0361_),
    .A(_0360_));
 sg13g2_nand2_1 _0971_ (.Y(_0362_),
    .A(_0359_),
    .B(_0361_));
 sg13g2_nor3_1 _0972_ (.A(_0354_),
    .B(_0356_),
    .C(_0362_),
    .Y(_0363_));
 sg13g2_nand3_1 _0973_ (.B(_0352_),
    .C(_0363_),
    .A(_0335_),
    .Y(_0364_));
 sg13g2_nor2_1 _0974_ (.A(_0545_),
    .B(_0060_),
    .Y(_0365_));
 sg13g2_nand3_1 _0975_ (.B(_0133_),
    .C(_0127_),
    .A(_0332_),
    .Y(_0366_));
 sg13g2_nor4_1 _0976_ (.A(_0191_),
    .B(_0365_),
    .C(_0168_),
    .D(_0366_),
    .Y(_0367_));
 sg13g2_nor3_1 _0977_ (.A(_0356_),
    .B(_0362_),
    .C(_0330_),
    .Y(_0368_));
 sg13g2_nand4_1 _0978_ (.B(_0368_),
    .C(_0126_),
    .A(_0367_),
    .Y(_0369_),
    .D(_0340_));
 sg13g2_nand2_1 _0979_ (.Y(_0370_),
    .A(_0364_),
    .B(_0369_));
 sg13g2_inv_1 _0980_ (.Y(_0371_),
    .A(_0348_));
 sg13g2_nor2_1 _0981_ (.A(_0318_),
    .B(_0349_),
    .Y(_0372_));
 sg13g2_nand3_1 _0982_ (.B(_0333_),
    .C(_0338_),
    .A(_0372_),
    .Y(_0373_));
 sg13g2_nor4_1 _0983_ (.A(_0296_),
    .B(_0365_),
    .C(_0371_),
    .D(_0373_),
    .Y(_0374_));
 sg13g2_a21oi_1 _0984_ (.A1(_0370_),
    .A2(_0206_),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_nor4_1 _0985_ (.A(_0205_),
    .B(_0159_),
    .C(_0061_),
    .D(_0356_),
    .Y(_0376_));
 sg13g2_nor2_1 _0986_ (.A(_0344_),
    .B(_0371_),
    .Y(_0377_));
 sg13g2_nand2_1 _0987_ (.Y(_0378_),
    .A(_0376_),
    .B(_0377_));
 sg13g2_nor3_1 _0988_ (.A(_0341_),
    .B(_0334_),
    .C(_0378_),
    .Y(_0380_));
 sg13g2_nand2_1 _0989_ (.Y(_0381_),
    .A(_0364_),
    .B(_0380_));
 sg13g2_nand2_1 _0990_ (.Y(_0382_),
    .A(_0381_),
    .B(_0390_));
 sg13g2_nand2_1 _0991_ (.Y(_0383_),
    .A(_0382_),
    .B(_0201_));
 sg13g2_nand2_1 _0992_ (.Y(_0384_),
    .A(_0375_),
    .B(_0383_));
 sg13g2_nand2_1 _0993_ (.Y(_0385_),
    .A(_0384_),
    .B(_0261_));
 sg13g2_nor3_1 _0994_ (.A(_0379_),
    .B(_0289_),
    .C(_0349_),
    .Y(_0386_));
 sg13g2_nor2b_1 _0995_ (.A(_0344_),
    .B_N(_0386_),
    .Y(_0387_));
 sg13g2_nand4_1 _0996_ (.B(_0363_),
    .C(_0340_),
    .A(_0335_),
    .Y(_0388_),
    .D(_0387_));
 sg13g2_inv_1 _0997_ (.Y(_0389_),
    .A(_0343_));
 sg13g2_nor4_1 _0998_ (.A(net14),
    .B(_0205_),
    .C(_0259_),
    .D(_0389_),
    .Y(_0391_));
 sg13g2_a21oi_1 _0999_ (.A1(_0391_),
    .A2(_0331_),
    .Y(_0392_),
    .B1(_0181_));
 sg13g2_nand2_1 _1000_ (.Y(_0393_),
    .A(_0364_),
    .B(_0250_));
 sg13g2_a21oi_1 _1001_ (.A1(_0388_),
    .A2(_0392_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_nand4_1 _1002_ (.B(_0056_),
    .C(_0032_),
    .A(_0293_),
    .Y(_0395_),
    .D(_0332_));
 sg13g2_nor3_1 _1003_ (.A(_0339_),
    .B(_0371_),
    .C(_0395_),
    .Y(_0396_));
 sg13g2_nand2_1 _1004_ (.Y(_0397_),
    .A(_0297_),
    .B(_0353_));
 sg13g2_nor3_1 _1005_ (.A(_0344_),
    .B(_0366_),
    .C(_0397_),
    .Y(_0398_));
 sg13g2_a21oi_1 _1006_ (.A1(_0396_),
    .A2(_0328_),
    .Y(_0399_),
    .B1(_0398_));
 sg13g2_o21ai_1 _1007_ (.B1(_0181_),
    .Y(_0400_),
    .A1(_0362_),
    .A2(_0399_));
 sg13g2_a21oi_1 _1008_ (.A1(_0394_),
    .A2(_0400_),
    .Y(_0402_),
    .B1(_0178_));
 sg13g2_nand2_1 _1009_ (.Y(_0403_),
    .A(_0385_),
    .B(_0402_));
 sg13g2_nand2_1 _1010_ (.Y(_0014_),
    .A(_0403_),
    .B(_0204_));
 sg13g2_nor3_1 _1011_ (.A(_0235_),
    .B(_0071_),
    .C(_0205_),
    .Y(_0404_));
 sg13g2_nand2_1 _1012_ (.Y(_0405_),
    .A(_0135_),
    .B(_0404_));
 sg13g2_nand3b_1 _1013_ (.B(_0291_),
    .C(_0108_),
    .Y(_0406_),
    .A_N(_0304_));
 sg13g2_nor2_1 _1014_ (.A(_0405_),
    .B(_0406_),
    .Y(_0407_));
 sg13g2_nand2_1 _1015_ (.Y(_0408_),
    .A(_0245_),
    .B(_0089_));
 sg13g2_nor2_1 _1016_ (.A(_0036_),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_nand2_1 _1017_ (.Y(_0410_),
    .A(_0409_),
    .B(_0361_));
 sg13g2_nand2_1 _1018_ (.Y(_0412_),
    .A(_0105_),
    .B(_0126_));
 sg13g2_nor2_1 _1019_ (.A(_0320_),
    .B(_0412_),
    .Y(_0413_));
 sg13g2_nor3_1 _1020_ (.A(_0061_),
    .B(_0144_),
    .C(_0209_),
    .Y(_0414_));
 sg13g2_nand2_1 _1021_ (.Y(_0415_),
    .A(_0413_),
    .B(_0414_));
 sg13g2_nor2_1 _1022_ (.A(_0410_),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_nand2_1 _1023_ (.Y(_0417_),
    .A(_0407_),
    .B(_0416_));
 sg13g2_nor2_1 _1024_ (.A(_0154_),
    .B(_0160_),
    .Y(_0418_));
 sg13g2_nor2_1 _1025_ (.A(_0092_),
    .B(_0065_),
    .Y(_0419_));
 sg13g2_nand3_1 _1026_ (.B(_0327_),
    .C(_0419_),
    .A(_0418_),
    .Y(_0420_));
 sg13g2_nor2_1 _1027_ (.A(_0230_),
    .B(_0315_),
    .Y(_0421_));
 sg13g2_nor2b_1 _1028_ (.A(_0420_),
    .B_N(_0421_),
    .Y(_0423_));
 sg13g2_nand2_1 _1029_ (.Y(_0424_),
    .A(_0112_),
    .B(_0127_));
 sg13g2_nor2_1 _1030_ (.A(_0337_),
    .B(_0424_),
    .Y(_0425_));
 sg13g2_nand2_1 _1031_ (.Y(_0426_),
    .A(_0425_),
    .B(_0021_));
 sg13g2_nor2_1 _1032_ (.A(_0037_),
    .B(_0252_),
    .Y(_0427_));
 sg13g2_nor2b_1 _1033_ (.A(_0426_),
    .B_N(_0427_),
    .Y(_0428_));
 sg13g2_inv_1 _1034_ (.Y(_0429_),
    .A(_0033_));
 sg13g2_nor2_1 _1035_ (.A(net8),
    .B(_0429_),
    .Y(_0430_));
 sg13g2_nor2_1 _1036_ (.A(_0329_),
    .B(_0241_),
    .Y(_0431_));
 sg13g2_nor3_1 _1037_ (.A(_0027_),
    .B(_0028_),
    .C(_0059_),
    .Y(_0432_));
 sg13g2_inv_1 _1038_ (.Y(_0433_),
    .A(_0432_));
 sg13g2_nand2_1 _1039_ (.Y(_0434_),
    .A(_0431_),
    .B(_0433_));
 sg13g2_nor2_1 _1040_ (.A(_0430_),
    .B(_0434_),
    .Y(_0435_));
 sg13g2_nand3_1 _1041_ (.B(_0428_),
    .C(_0435_),
    .A(_0423_),
    .Y(_0436_));
 sg13g2_nor3_1 _1042_ (.A(net13),
    .B(_0417_),
    .C(_0436_),
    .Y(_0437_));
 sg13g2_nor2_1 _1043_ (.A(_0217_),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_inv_1 _1044_ (.Y(_0439_),
    .A(_0409_));
 sg13g2_nor4_1 _1045_ (.A(_0337_),
    .B(_0439_),
    .C(_0211_),
    .D(_0406_),
    .Y(_0440_));
 sg13g2_nand3_1 _1046_ (.B(net13),
    .C(_0440_),
    .A(_0249_),
    .Y(_0441_));
 sg13g2_nand2_1 _1047_ (.Y(_0442_),
    .A(_0438_),
    .B(_0441_));
 sg13g2_nor3_1 _1048_ (.A(_0329_),
    .B(_0432_),
    .C(_0241_),
    .Y(_0444_));
 sg13g2_nor3_1 _1049_ (.A(_0099_),
    .B(_0337_),
    .C(_0259_),
    .Y(_0445_));
 sg13g2_nand2_1 _1050_ (.Y(_0446_),
    .A(_0255_),
    .B(_0074_));
 sg13g2_nor2_1 _1051_ (.A(_0304_),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_nand4_1 _1052_ (.B(_0445_),
    .C(_0447_),
    .A(_0444_),
    .Y(_0448_),
    .D(_0404_));
 sg13g2_nor2b_1 _1053_ (.A(_0448_),
    .B_N(_0416_),
    .Y(_0449_));
 sg13g2_nand3_1 _1054_ (.B(net13),
    .C(_0449_),
    .A(net7),
    .Y(_0450_));
 sg13g2_nand2_1 _1055_ (.Y(_0451_),
    .A(_0427_),
    .B(_0079_));
 sg13g2_a221oi_1 _1056_ (.B2(_0141_),
    .C1(_0530_),
    .B1(_0524_),
    .A1(_0033_),
    .Y(_0452_),
    .A2(_0030_));
 sg13g2_nand2_1 _1057_ (.Y(_0453_),
    .A(_0452_),
    .B(_0021_));
 sg13g2_nor3_1 _1058_ (.A(_0410_),
    .B(_0451_),
    .C(_0453_),
    .Y(_0455_));
 sg13g2_a21oi_1 _1059_ (.A1(_0455_),
    .A2(net14),
    .Y(_0456_),
    .B1(_0201_));
 sg13g2_nand2_1 _1060_ (.Y(_0457_),
    .A(_0450_),
    .B(_0456_));
 sg13g2_nand2_1 _1061_ (.Y(_0458_),
    .A(_0442_),
    .B(_0457_));
 sg13g2_nand2_1 _1062_ (.Y(_0459_),
    .A(_0458_),
    .B(_0250_));
 sg13g2_nand2b_1 _1063_ (.Y(_0460_),
    .B(_0100_),
    .A_N(_0430_));
 sg13g2_nand4_1 _1064_ (.B(_0167_),
    .C(_0112_),
    .A(_0359_),
    .Y(_0461_),
    .D(_0127_));
 sg13g2_nor4_1 _1065_ (.A(_0356_),
    .B(_0460_),
    .C(_0405_),
    .D(_0461_),
    .Y(_0462_));
 sg13g2_nand2_1 _1066_ (.Y(_0463_),
    .A(net7),
    .B(_0462_));
 sg13g2_nand2_1 _1067_ (.Y(_0464_),
    .A(_0463_),
    .B(net14));
 sg13g2_nand2_1 _1068_ (.Y(_0466_),
    .A(_0291_),
    .B(_0260_));
 sg13g2_nand4_1 _1069_ (.B(_0355_),
    .C(_0067_),
    .A(_0361_),
    .Y(_0467_),
    .D(_0216_));
 sg13g2_nor3_1 _1070_ (.A(_0134_),
    .B(_0466_),
    .C(_0467_),
    .Y(_0468_));
 sg13g2_nor3_1 _1071_ (.A(_0430_),
    .B(_0434_),
    .C(_0451_),
    .Y(_0469_));
 sg13g2_nand2_1 _1072_ (.Y(_0470_),
    .A(_0468_),
    .B(_0469_));
 sg13g2_nand3_1 _1073_ (.B(net13),
    .C(_0470_),
    .A(net7),
    .Y(_0471_));
 sg13g2_nand3_1 _1074_ (.B(_0471_),
    .C(_0181_),
    .A(_0464_),
    .Y(_0472_));
 sg13g2_nand2_1 _1075_ (.Y(_0473_),
    .A(_0428_),
    .B(_0444_));
 sg13g2_nor2_1 _1076_ (.A(_0473_),
    .B(_0417_),
    .Y(_0474_));
 sg13g2_nand2_1 _1077_ (.Y(_0475_),
    .A(net7),
    .B(_0474_));
 sg13g2_nand2_1 _1078_ (.Y(_0476_),
    .A(_0475_),
    .B(_0358_));
 sg13g2_nand2_1 _1079_ (.Y(_0477_),
    .A(_0476_),
    .B(_0153_));
 sg13g2_nand2_1 _1080_ (.Y(_0478_),
    .A(_0472_),
    .B(_0477_));
 sg13g2_nand2_1 _1081_ (.Y(_0479_),
    .A(_0459_),
    .B(_0478_));
 sg13g2_nand2_1 _1082_ (.Y(_0480_),
    .A(_0479_),
    .B(_0310_));
 sg13g2_nand2_1 _1083_ (.Y(_0015_),
    .A(_0480_),
    .B(_0204_));
 sg13g2_nand2_1 _1084_ (.Y(_0481_),
    .A(_0245_),
    .B(_0067_));
 sg13g2_nand3_1 _1085_ (.B(_0115_),
    .C(_0216_),
    .A(_0207_),
    .Y(_0482_));
 sg13g2_nor3_1 _1086_ (.A(_0220_),
    .B(_0481_),
    .C(_0482_),
    .Y(_0483_));
 sg13g2_nand3_1 _1087_ (.B(net13),
    .C(_0483_),
    .A(_0251_),
    .Y(_0484_));
 sg13g2_nor3_1 _1088_ (.A(_0209_),
    .B(_0342_),
    .C(_0101_),
    .Y(_0486_));
 sg13g2_nand3_1 _1089_ (.B(net14),
    .C(_0246_),
    .A(_0486_),
    .Y(_0487_));
 sg13g2_a21oi_1 _1090_ (.A1(_0484_),
    .A2(_0487_),
    .Y(_0488_),
    .B1(_0153_));
 sg13g2_nor2_1 _1091_ (.A(_0522_),
    .B(_0062_),
    .Y(_0489_));
 sg13g2_nor2_1 _1092_ (.A(_0326_),
    .B(_0221_),
    .Y(_0490_));
 sg13g2_inv_1 _1093_ (.Y(_0491_),
    .A(_0490_));
 sg13g2_nor2_1 _1094_ (.A(_0489_),
    .B(_0491_),
    .Y(_0492_));
 sg13g2_nand4_1 _1095_ (.B(net13),
    .C(_0248_),
    .A(_0251_),
    .Y(_0493_),
    .D(_0492_));
 sg13g2_nand3_1 _1096_ (.B(_0248_),
    .C(_0325_),
    .A(_0240_),
    .Y(_0494_));
 sg13g2_nor3_1 _1097_ (.A(_0257_),
    .B(_0211_),
    .C(_0208_),
    .Y(_0495_));
 sg13g2_nand3b_1 _1098_ (.B(_0222_),
    .C(_0495_),
    .Y(_0497_),
    .A_N(_0494_));
 sg13g2_a21oi_1 _1099_ (.A1(_0493_),
    .A2(_0497_),
    .Y(_0498_),
    .B1(_0401_));
 sg13g2_nor2_1 _1100_ (.A(_0488_),
    .B(_0498_),
    .Y(_0499_));
 sg13g2_nand3_1 _1101_ (.B(_0108_),
    .C(_0207_),
    .A(_0212_),
    .Y(_0500_));
 sg13g2_nor3_1 _1102_ (.A(_0218_),
    .B(_0243_),
    .C(_0500_),
    .Y(_0501_));
 sg13g2_nand2_1 _1103_ (.Y(_0502_),
    .A(net7),
    .B(_0501_));
 sg13g2_a21oi_1 _1104_ (.A1(_0502_),
    .A2(_0001_),
    .Y(_0503_),
    .B1(_0173_));
 sg13g2_inv_1 _1105_ (.Y(_0504_),
    .A(_0213_));
 sg13g2_o21ai_1 _1106_ (.B1(_0108_),
    .Y(_0505_),
    .A1(net15),
    .A2(_0064_));
 sg13g2_nor2_1 _1107_ (.A(_0481_),
    .B(_0505_),
    .Y(_0506_));
 sg13g2_nand4_1 _1108_ (.B(_0246_),
    .C(_0244_),
    .A(_0504_),
    .Y(_0508_),
    .D(_0506_));
 sg13g2_nand3_1 _1109_ (.B(_0508_),
    .C(_0390_),
    .A(net7),
    .Y(_0509_));
 sg13g2_nand3_1 _1110_ (.B(_0531_),
    .C(_0215_),
    .A(_0242_),
    .Y(_0510_));
 sg13g2_o21ai_1 _1111_ (.B1(_0325_),
    .Y(_0511_),
    .A1(_0491_),
    .A2(_0510_));
 sg13g2_nand3_1 _1112_ (.B(_0151_),
    .C(_0511_),
    .A(_0509_),
    .Y(_0512_));
 sg13g2_nand2_1 _1113_ (.Y(_0513_),
    .A(_0512_),
    .B(_0310_));
 sg13g2_nor2_1 _1114_ (.A(_0503_),
    .B(_0513_),
    .Y(_0514_));
 sg13g2_nand2_1 _1115_ (.Y(_0515_),
    .A(_0499_),
    .B(_0514_));
 sg13g2_nand2_1 _1116_ (.Y(_0016_),
    .A(_0515_),
    .B(_0204_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \uart_tx.bit_counter[0]$_SDFF_PP0__35  (.L_HI(net35));
 sg13g2_buf_1 _1119_ (.A(net16),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1120_ (.A(net17),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1121_ (.A(net18),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1122_ (.A(net19),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1123_ (.A(net20),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1124_ (.A(net21),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1125_ (.A(net22),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1126_ (.A(net23),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1127_ (.A(net24),
    .X(uio_out[0]));
 sg13g2_buf_1 _1128_ (.A(net25),
    .X(uio_out[1]));
 sg13g2_buf_1 _1129_ (.A(net26),
    .X(uio_out[2]));
 sg13g2_buf_1 _1130_ (.A(net27),
    .X(uio_out[3]));
 sg13g2_buf_1 _1131_ (.A(net28),
    .X(uio_out[4]));
 sg13g2_buf_1 _1132_ (.A(net29),
    .X(uio_out[5]));
 sg13g2_buf_1 _1133_ (.A(net30),
    .X(uio_out[6]));
 sg13g2_buf_1 _1134_ (.A(net31),
    .X(uio_out[7]));
 sg13g2_buf_1 _1135_ (.A(tx_pin0),
    .X(net2));
 sg13g2_buf_1 _1136_ (.A(tx_pin1),
    .X(net3));
 sg13g2_buf_1 _1137_ (.A(tx_pin2),
    .X(net4));
 sg13g2_buf_1 _1138_ (.A(tx_pin3),
    .X(net5));
 sg13g2_buf_1 _1139_ (.A(tx_pin4),
    .X(net6));
 sg13g2_buf_1 _1140_ (.A(net32),
    .X(uo_out[5]));
 sg13g2_buf_1 _1141_ (.A(net33),
    .X(uo_out[6]));
 sg13g2_buf_1 _1142_ (.A(net34),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \uart_tx.bit_counter[0]$_SDFF_PP0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net35),
    .D(_0002_),
    .Q_N(_0001_),
    .Q(\uart_tx.bit_counter[0] ));
 sg13g2_dfrbp_1 \uart_tx.bit_counter[1]$_SDFF_PP0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net36),
    .D(_0003_),
    .Q_N(_0000_),
    .Q(\uart_tx.bit_counter[1] ));
 sg13g2_dfrbp_1 \uart_tx.bit_counter[2]$_SDFF_PP0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net37),
    .D(_0004_),
    .Q_N(_0564_),
    .Q(\uart_tx.bit_counter[2] ));
 sg13g2_dfrbp_1 \uart_tx.bit_counter[3]$_SDFF_PP0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net38),
    .D(_0005_),
    .Q_N(_0563_),
    .Q(\uart_tx.bit_counter[3] ));
 sg13g2_dfrbp_1 \uart_tx.text_index[0]$_SDFFE_PN0P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net39),
    .D(_0006_),
    .Q_N(_0562_),
    .Q(\uart_tx.text_index[0] ));
 sg13g2_dfrbp_1 \uart_tx.text_index[1]$_SDFFE_PN0P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net40),
    .D(_0007_),
    .Q_N(_0561_),
    .Q(\uart_tx.text_index[1] ));
 sg13g2_dfrbp_1 \uart_tx.text_index[2]$_SDFFE_PN0P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net41),
    .D(_0008_),
    .Q_N(_0560_),
    .Q(\uart_tx.text_index[2] ));
 sg13g2_dfrbp_1 \uart_tx.text_index[3]$_SDFFE_PN0P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net42),
    .D(_0009_),
    .Q_N(_0559_),
    .Q(\uart_tx.text_index[3] ));
 sg13g2_dfrbp_1 \uart_tx.text_index[4]$_SDFFE_PN0P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net43),
    .D(_0010_),
    .Q_N(_0558_),
    .Q(\uart_tx.text_index[4] ));
 sg13g2_dfrbp_1 \uart_tx.text_index[5]$_SDFFE_PN0P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net44),
    .D(_0011_),
    .Q_N(_0557_),
    .Q(\uart_tx.text_index[5] ));
 sg13g2_dfrbp_1 \uart_tx.tx_pin0_int$_SDFF_PN1_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net45),
    .D(_0012_),
    .Q_N(_0556_),
    .Q(tx_pin0));
 sg13g2_dfrbp_1 \uart_tx.tx_pin1_int$_SDFF_PN1_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net46),
    .D(_0013_),
    .Q_N(_0555_),
    .Q(tx_pin1));
 sg13g2_dfrbp_1 \uart_tx.tx_pin2_int$_SDFF_PN1_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net47),
    .D(_0014_),
    .Q_N(_0554_),
    .Q(tx_pin2));
 sg13g2_dfrbp_1 \uart_tx.tx_pin3_int$_SDFF_PN1_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net48),
    .D(_0015_),
    .Q_N(_0553_),
    .Q(tx_pin3));
 sg13g2_dfrbp_1 \uart_tx.tx_pin4_int$_SDFF_PN1_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net49),
    .D(_0016_),
    .Q_N(_0552_),
    .Q(tx_pin4));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_2 fanout7 (.A(_0251_),
    .X(net7));
 sg13g2_buf_2 fanout8 (.A(_0059_),
    .X(net8));
 sg13g2_buf_2 fanout9 (.A(_0034_),
    .X(net9));
 sg13g2_buf_2 fanout10 (.A(_0053_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_0023_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0528_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0390_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0325_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0522_),
    .X(net15));
 sg13g2_tielo _1119__16 (.L_LO(net16));
 sg13g2_tielo _1120__17 (.L_LO(net17));
 sg13g2_tielo _1121__18 (.L_LO(net18));
 sg13g2_tielo _1122__19 (.L_LO(net19));
 sg13g2_tielo _1123__20 (.L_LO(net20));
 sg13g2_tielo _1124__21 (.L_LO(net21));
 sg13g2_tielo _1125__22 (.L_LO(net22));
 sg13g2_tielo _1126__23 (.L_LO(net23));
 sg13g2_tielo _1127__24 (.L_LO(net24));
 sg13g2_tielo _1128__25 (.L_LO(net25));
 sg13g2_tielo _1129__26 (.L_LO(net26));
 sg13g2_tielo _1130__27 (.L_LO(net27));
 sg13g2_tielo _1131__28 (.L_LO(net28));
 sg13g2_tielo _1132__29 (.L_LO(net29));
 sg13g2_tielo _1133__30 (.L_LO(net30));
 sg13g2_tielo _1134__31 (.L_LO(net31));
 sg13g2_tielo _1140__32 (.L_LO(net32));
 sg13g2_tielo _1141__33 (.L_LO(net33));
 sg13g2_tielo _1142__34 (.L_LO(net34));
 sg13g2_tiehi \uart_tx.bit_counter[1]$_SDFF_PP0__36  (.L_HI(net36));
 sg13g2_tiehi \uart_tx.bit_counter[2]$_SDFF_PP0__37  (.L_HI(net37));
 sg13g2_tiehi \uart_tx.bit_counter[3]$_SDFF_PP0__38  (.L_HI(net38));
 sg13g2_tiehi \uart_tx.text_index[0]$_SDFFE_PN0P__39  (.L_HI(net39));
 sg13g2_tiehi \uart_tx.text_index[1]$_SDFFE_PN0P__40  (.L_HI(net40));
 sg13g2_tiehi \uart_tx.text_index[2]$_SDFFE_PN0P__41  (.L_HI(net41));
 sg13g2_tiehi \uart_tx.text_index[3]$_SDFFE_PN0P__42  (.L_HI(net42));
 sg13g2_tiehi \uart_tx.text_index[4]$_SDFFE_PN0P__43  (.L_HI(net43));
 sg13g2_tiehi \uart_tx.text_index[5]$_SDFFE_PN0P__44  (.L_HI(net44));
 sg13g2_tiehi \uart_tx.tx_pin0_int$_SDFF_PN1__45  (.L_HI(net45));
 sg13g2_tiehi \uart_tx.tx_pin1_int$_SDFF_PN1__46  (.L_HI(net46));
 sg13g2_tiehi \uart_tx.tx_pin2_int$_SDFF_PN1__47  (.L_HI(net47));
 sg13g2_tiehi \uart_tx.tx_pin3_int$_SDFF_PN1__48  (.L_HI(net48));
 sg13g2_tiehi \uart_tx.tx_pin4_int$_SDFF_PN1__49  (.L_HI(net49));
 sg13g2_buf_1 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_1 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_1 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_1 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_3__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_fill_2 FILLER_20_427 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_4 FILLER_22_301 ();
 sg13g2_fill_2 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_decap_8 FILLER_22_327 ();
 sg13g2_decap_8 FILLER_22_334 ();
 sg13g2_decap_8 FILLER_22_341 ();
 sg13g2_decap_8 FILLER_22_348 ();
 sg13g2_decap_8 FILLER_22_355 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_8 FILLER_22_404 ();
 sg13g2_decap_8 FILLER_22_411 ();
 sg13g2_decap_8 FILLER_22_418 ();
 sg13g2_decap_4 FILLER_22_425 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_4 FILLER_23_287 ();
 sg13g2_fill_1 FILLER_23_291 ();
 sg13g2_fill_2 FILLER_23_301 ();
 sg13g2_decap_4 FILLER_23_307 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_fill_1 FILLER_23_322 ();
 sg13g2_decap_4 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_332 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_23_409 ();
 sg13g2_decap_8 FILLER_23_416 ();
 sg13g2_decap_8 FILLER_23_423 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_decap_4 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_216 ();
 sg13g2_decap_4 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_280 ();
 sg13g2_fill_1 FILLER_24_298 ();
 sg13g2_fill_1 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_335 ();
 sg13g2_fill_2 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_fill_2 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_2 FILLER_25_217 ();
 sg13g2_fill_1 FILLER_25_219 ();
 sg13g2_decap_4 FILLER_25_250 ();
 sg13g2_fill_2 FILLER_25_262 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_311 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_4 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_2 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_fill_1 FILLER_26_240 ();
 sg13g2_fill_2 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_259 ();
 sg13g2_fill_1 FILLER_26_275 ();
 sg13g2_fill_2 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_347 ();
 sg13g2_fill_1 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_368 ();
 sg13g2_fill_2 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_decap_8 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_26_414 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_fill_1 FILLER_27_196 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_219 ();
 sg13g2_fill_1 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_fill_1 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_304 ();
 sg13g2_fill_2 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_fill_2 FILLER_27_353 ();
 sg13g2_fill_1 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_decap_8 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_27_414 ();
 sg13g2_decap_8 FILLER_27_421 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_fill_2 FILLER_28_196 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_fill_1 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_236 ();
 sg13g2_fill_1 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_1 FILLER_28_293 ();
 sg13g2_fill_2 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_340 ();
 sg13g2_fill_2 FILLER_28_392 ();
 sg13g2_fill_2 FILLER_28_400 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_4 FILLER_28_426 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_4 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_245 ();
 sg13g2_fill_2 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_337 ();
 sg13g2_fill_1 FILLER_29_375 ();
 sg13g2_fill_2 FILLER_29_381 ();
 sg13g2_fill_1 FILLER_29_387 ();
 sg13g2_fill_2 FILLER_29_414 ();
 sg13g2_fill_1 FILLER_29_416 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_4 FILLER_30_161 ();
 sg13g2_fill_1 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_245 ();
 sg13g2_fill_1 FILLER_30_250 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_fill_1 FILLER_30_264 ();
 sg13g2_fill_1 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_fill_1 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_401 ();
 sg13g2_fill_2 FILLER_30_408 ();
 sg13g2_fill_1 FILLER_30_410 ();
 sg13g2_fill_2 FILLER_30_415 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_4 FILLER_31_161 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_277 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_fill_2 FILLER_31_355 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_decap_4 FILLER_31_425 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_175 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_decap_4 FILLER_32_229 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_fill_1 FILLER_32_261 ();
 sg13g2_fill_2 FILLER_32_267 ();
 sg13g2_fill_1 FILLER_32_275 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_1 FILLER_32_327 ();
 sg13g2_fill_2 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_375 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_175 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_2 FILLER_33_190 ();
 sg13g2_fill_1 FILLER_33_206 ();
 sg13g2_decap_4 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_fill_1 FILLER_33_246 ();
 sg13g2_fill_1 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_267 ();
 sg13g2_fill_2 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_fill_1 FILLER_33_359 ();
 sg13g2_fill_1 FILLER_33_364 ();
 sg13g2_fill_1 FILLER_33_370 ();
 sg13g2_fill_1 FILLER_33_379 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_4 FILLER_34_189 ();
 sg13g2_fill_2 FILLER_34_193 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_fill_1 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_233 ();
 sg13g2_fill_1 FILLER_34_251 ();
 sg13g2_fill_1 FILLER_34_255 ();
 sg13g2_fill_2 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_300 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_318 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_fill_2 FILLER_34_427 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_215 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_decap_4 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_248 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_fill_2 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_fill_2 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_fill_2 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_331 ();
 sg13g2_fill_1 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_410 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_4 FILLER_36_424 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_decap_4 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_fill_1 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_4 FILLER_37_365 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_decap_4 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_8 FILLER_37_404 ();
 sg13g2_decap_8 FILLER_37_411 ();
 sg13g2_decap_8 FILLER_37_418 ();
 sg13g2_decap_4 FILLER_37_425 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_298 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_decap_4 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_377 ();
 sg13g2_decap_8 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_391 ();
 sg13g2_decap_8 FILLER_38_398 ();
 sg13g2_decap_8 FILLER_38_405 ();
 sg13g2_decap_8 FILLER_38_412 ();
 sg13g2_decap_8 FILLER_38_419 ();
 sg13g2_decap_4 FILLER_38_426 ();
endmodule
