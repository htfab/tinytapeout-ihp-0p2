module tt_um_cejmu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire clknet_0_clk;
 wire net73;
 wire \cla_z[0] ;
 wire \cla_z[10] ;
 wire \cla_z[11] ;
 wire \cla_z[12] ;
 wire \cla_z[13] ;
 wire \cla_z[14] ;
 wire \cla_z[15] ;
 wire \cla_z[16] ;
 wire \cla_z[17] ;
 wire \cla_z[18] ;
 wire \cla_z[19] ;
 wire \cla_z[1] ;
 wire \cla_z[20] ;
 wire \cla_z[21] ;
 wire \cla_z[22] ;
 wire \cla_z[23] ;
 wire \cla_z[2] ;
 wire \cla_z[3] ;
 wire \cla_z[4] ;
 wire \cla_z[5] ;
 wire \cla_z[6] ;
 wire \cla_z[7] ;
 wire \cla_z[8] ;
 wire \cla_z[9] ;
 wire \io_sd._052_[0] ;
 wire \io_sd._052_[10] ;
 wire \io_sd._052_[11] ;
 wire \io_sd._052_[12] ;
 wire \io_sd._052_[13] ;
 wire \io_sd._052_[14] ;
 wire \io_sd._052_[15] ;
 wire \io_sd._052_[16] ;
 wire \io_sd._052_[17] ;
 wire \io_sd._052_[18] ;
 wire \io_sd._052_[19] ;
 wire \io_sd._052_[1] ;
 wire \io_sd._052_[20] ;
 wire \io_sd._052_[21] ;
 wire \io_sd._052_[22] ;
 wire \io_sd._052_[23] ;
 wire \io_sd._052_[2] ;
 wire \io_sd._052_[3] ;
 wire \io_sd._052_[4] ;
 wire \io_sd._052_[5] ;
 wire \io_sd._052_[6] ;
 wire \io_sd._052_[7] ;
 wire \io_sd._052_[8] ;
 wire \io_sd._052_[9] ;
 wire \io_sd._053_[0] ;
 wire \io_sd._053_[10] ;
 wire \io_sd._053_[11] ;
 wire \io_sd._053_[12] ;
 wire \io_sd._053_[13] ;
 wire \io_sd._053_[14] ;
 wire \io_sd._053_[15] ;
 wire \io_sd._053_[16] ;
 wire \io_sd._053_[17] ;
 wire \io_sd._053_[18] ;
 wire \io_sd._053_[19] ;
 wire \io_sd._053_[1] ;
 wire \io_sd._053_[20] ;
 wire \io_sd._053_[21] ;
 wire \io_sd._053_[22] ;
 wire \io_sd._053_[23] ;
 wire \io_sd._053_[2] ;
 wire \io_sd._053_[3] ;
 wire \io_sd._053_[4] ;
 wire \io_sd._053_[5] ;
 wire \io_sd._053_[6] ;
 wire \io_sd._053_[7] ;
 wire \io_sd._053_[8] ;
 wire \io_sd._053_[9] ;
 wire \io_sd._068_ ;
 wire \io_sd._092_ ;
 wire \io_sd._209_[0] ;
 wire \io_sd._210_[0] ;
 wire \io_sd.input_index[3] ;
 wire \io_sd.input_index[4] ;
 wire \io_sd.input_index[5] ;
 wire \io_sd.output_index[3] ;
 wire \io_sd.output_index[4] ;
 wire \io_sd.output_index[5] ;
 wire \rca.generate_adder_modules[0].fa.a ;
 wire \rca.generate_adder_modules[0].fa.b ;
 wire \rca.generate_adder_modules[10].fa.a ;
 wire \rca.generate_adder_modules[10].fa.b ;
 wire \rca.generate_adder_modules[11].fa.a ;
 wire \rca.generate_adder_modules[11].fa.b ;
 wire \rca.generate_adder_modules[12].fa.a ;
 wire \rca.generate_adder_modules[12].fa.b ;
 wire \rca.generate_adder_modules[13].fa.a ;
 wire \rca.generate_adder_modules[13].fa.b ;
 wire \rca.generate_adder_modules[14].fa.a ;
 wire \rca.generate_adder_modules[14].fa.b ;
 wire \rca.generate_adder_modules[15].fa.a ;
 wire \rca.generate_adder_modules[15].fa.b ;
 wire \rca.generate_adder_modules[16].fa.a ;
 wire \rca.generate_adder_modules[16].fa.b ;
 wire \rca.generate_adder_modules[17].fa.a ;
 wire \rca.generate_adder_modules[17].fa.b ;
 wire \rca.generate_adder_modules[18].fa.a ;
 wire \rca.generate_adder_modules[18].fa.b ;
 wire \rca.generate_adder_modules[19].fa.a ;
 wire \rca.generate_adder_modules[19].fa.b ;
 wire \rca.generate_adder_modules[1].fa.a ;
 wire \rca.generate_adder_modules[1].fa.b ;
 wire \rca.generate_adder_modules[20].fa.a ;
 wire \rca.generate_adder_modules[20].fa.b ;
 wire \rca.generate_adder_modules[21].fa.a ;
 wire \rca.generate_adder_modules[21].fa.b ;
 wire \rca.generate_adder_modules[22].fa.a ;
 wire \rca.generate_adder_modules[22].fa.b ;
 wire \rca.generate_adder_modules[23].fa.a ;
 wire \rca.generate_adder_modules[23].fa.b ;
 wire \rca.generate_adder_modules[23].fa.c_out ;
 wire \rca.generate_adder_modules[2].fa.a ;
 wire \rca.generate_adder_modules[2].fa.b ;
 wire \rca.generate_adder_modules[3].fa.a ;
 wire \rca.generate_adder_modules[3].fa.b ;
 wire \rca.generate_adder_modules[4].fa.a ;
 wire \rca.generate_adder_modules[4].fa.b ;
 wire \rca.generate_adder_modules[5].fa.a ;
 wire \rca.generate_adder_modules[5].fa.b ;
 wire \rca.generate_adder_modules[6].fa.a ;
 wire \rca.generate_adder_modules[6].fa.b ;
 wire \rca.generate_adder_modules[7].fa.a ;
 wire \rca.generate_adder_modules[7].fa.b ;
 wire \rca.generate_adder_modules[8].fa.a ;
 wire \rca.generate_adder_modules[8].fa.b ;
 wire \rca.generate_adder_modules[9].fa.a ;
 wire \rca.generate_adder_modules[9].fa.b ;
 wire \cla/_0341_ ;
 wire \cla/_0342_ ;
 wire \cla/_0343_ ;
 wire \cla/_0344_ ;
 wire \cla/_0345_ ;
 wire \cla/_0346_ ;
 wire \cla/_0347_ ;
 wire \cla/_0348_ ;
 wire \cla/_0349_ ;
 wire \cla/_0350_ ;
 wire \cla/_0351_ ;
 wire \cla/_0352_ ;
 wire \cla/_0353_ ;
 wire \cla/_0354_ ;
 wire \cla/_0355_ ;
 wire \cla/_0356_ ;
 wire \cla/_0357_ ;
 wire \cla/_0358_ ;
 wire \cla/_0359_ ;
 wire \cla/_0360_ ;
 wire \cla/_0361_ ;
 wire \cla/_0362_ ;
 wire \cla/_0363_ ;
 wire \cla/_0364_ ;
 wire \cla/_0365_ ;
 wire \cla/_0366_ ;
 wire \cla/_0367_ ;
 wire \cla/_0368_ ;
 wire \cla/_0369_ ;
 wire \cla/_0370_ ;
 wire \cla/_0371_ ;
 wire \cla/_0372_ ;
 wire \cla/_0373_ ;
 wire \cla/_0374_ ;
 wire \cla/_0375_ ;
 wire \cla/_0376_ ;
 wire \cla/_0377_ ;
 wire \cla/_0378_ ;
 wire \cla/_0379_ ;
 wire \cla/_0380_ ;
 wire \cla/_0381_ ;
 wire \cla/_0382_ ;
 wire \cla/_0383_ ;
 wire \cla/_0384_ ;
 wire \cla/_0385_ ;
 wire \cla/_0386_ ;
 wire \cla/_0387_ ;
 wire \cla/_0388_ ;
 wire \cla/_0389_ ;
 wire \cla/_0390_ ;
 wire \cla/_0391_ ;
 wire \cla/_0392_ ;
 wire \cla/_0393_ ;
 wire \cla/_0394_ ;
 wire \cla/_0395_ ;
 wire \cla/_0396_ ;
 wire \cla/_0397_ ;
 wire \cla/_0398_ ;
 wire \cla/_0399_ ;
 wire \cla/_0400_ ;
 wire \cla/_0401_ ;
 wire \cla/_0402_ ;
 wire \cla/_0403_ ;
 wire \cla/_0404_ ;
 wire \cla/_0405_ ;
 wire \cla/_0406_ ;
 wire \cla/_0407_ ;
 wire \cla/_0408_ ;
 wire \cla/_0409_ ;
 wire \cla/_0410_ ;
 wire \cla/_0411_ ;
 wire \cla/_0412_ ;
 wire \cla/_0413_ ;
 wire \cla/_0414_ ;
 wire \cla/_0415_ ;
 wire \cla/_0416_ ;
 wire \cla/_0417_ ;
 wire \cla/_0418_ ;
 wire \cla/_0419_ ;
 wire \cla/_0420_ ;
 wire \cla/_0421_ ;
 wire \cla/_0422_ ;
 wire \cla/_0423_ ;
 wire \cla/_0424_ ;
 wire \cla/_0425_ ;
 wire \cla/_0426_ ;
 wire \cla/_0427_ ;
 wire \cla/_0428_ ;
 wire \cla/_0429_ ;
 wire \cla/_0430_ ;
 wire \cla/_0431_ ;
 wire \cla/_0432_ ;
 wire \cla/_0433_ ;
 wire \cla/_0434_ ;
 wire \cla/_0435_ ;
 wire \cla/_0436_ ;
 wire \cla/_0437_ ;
 wire \cla/_0438_ ;
 wire \cla/_0439_ ;
 wire \cla/_0440_ ;
 wire \cla/_0441_ ;
 wire \cla/_0442_ ;
 wire \cla/_0443_ ;
 wire \cla/_0444_ ;
 wire \cla/_0445_ ;
 wire \cla/_0446_ ;
 wire \cla/_0447_ ;
 wire \cla/_0448_ ;
 wire \cla/_0449_ ;
 wire \cla/_0450_ ;
 wire \cla/_0451_ ;
 wire \cla/_0452_ ;
 wire \cla/_0453_ ;
 wire \cla/_0454_ ;
 wire \cla/_0455_ ;
 wire \cla/_0456_ ;
 wire \cla/_0457_ ;
 wire \cla/_0458_ ;
 wire \cla/_0459_ ;
 wire \cla/_0460_ ;
 wire \cla/_0461_ ;
 wire \cla/_0462_ ;
 wire \cla/_0463_ ;
 wire \cla/_0464_ ;
 wire \cla/_0465_ ;
 wire \cla/_0466_ ;
 wire \cla/_0467_ ;
 wire \cla/_0468_ ;
 wire \cla/_0469_ ;
 wire \cla/_0470_ ;
 wire \cla/_0471_ ;
 wire \cla/_0472_ ;
 wire \cla/_0473_ ;
 wire \cla/_0474_ ;
 wire \cla/_0475_ ;
 wire \cla/_0476_ ;
 wire \cla/_0477_ ;
 wire \cla/_0478_ ;
 wire \cla/_0479_ ;
 wire \cla/_0480_ ;
 wire \cla/_0481_ ;
 wire \cla/_0482_ ;
 wire \cla/_0483_ ;
 wire \cla/_0484_ ;
 wire \cla/_0485_ ;
 wire \cla/_0486_ ;
 wire \cla/_0487_ ;
 wire \cla/_0488_ ;
 wire \cla/_0489_ ;
 wire \cla/_0490_ ;
 wire \cla/_0491_ ;
 wire \cla/_0492_ ;
 wire \cla/_0493_ ;
 wire \cla/_0494_ ;
 wire \cla/_0495_ ;
 wire \cla/_0496_ ;
 wire \cla/_0497_ ;
 wire \cla/_0498_ ;
 wire \cla/_0499_ ;
 wire \cla/_0500_ ;
 wire \cla/_0501_ ;
 wire \cla/_0502_ ;
 wire \cla/_0503_ ;
 wire \cla/_0504_ ;
 wire \cla/_0505_ ;
 wire \cla/_0506_ ;
 wire \cla/_0507_ ;
 wire \cla/_0508_ ;
 wire \cla/_0509_ ;
 wire \cla/_0510_ ;
 wire \cla/_0511_ ;
 wire \cla/_0512_ ;
 wire \cla/_0513_ ;
 wire \cla/_0514_ ;
 wire \cla/_0515_ ;
 wire \cla/_0516_ ;
 wire \cla/_0517_ ;
 wire \cla/_0518_ ;
 wire \cla/_0519_ ;
 wire \cla/_0520_ ;
 wire \cla/_0521_ ;
 wire \cla/_0522_ ;
 wire \cla/_0523_ ;
 wire \cla/_0524_ ;
 wire \cla/_0525_ ;
 wire \cla/_0526_ ;
 wire \cla/_0527_ ;
 wire \cla/_0528_ ;
 wire \cla/_0529_ ;
 wire \cla/_0530_ ;
 wire \cla/_0531_ ;
 wire \cla/_0532_ ;
 wire \cla/_0533_ ;
 wire \cla/_0534_ ;
 wire \cla/_0535_ ;
 wire \cla/_0536_ ;
 wire \cla/_0537_ ;
 wire \cla/_0538_ ;
 wire \cla/_0539_ ;
 wire \cla/_0540_ ;
 wire \cla/_0541_ ;
 wire \cla/_0542_ ;
 wire \cla/_0543_ ;
 wire \cla/_0544_ ;
 wire \cla/_0545_ ;
 wire \cla/_0546_ ;
 wire \cla/_0547_ ;
 wire \cla/_0548_ ;
 wire \cla/_0549_ ;
 wire \cla/_0550_ ;
 wire \cla/_0551_ ;
 wire \cla/_0552_ ;
 wire \cla/_0553_ ;
 wire \cla/_0554_ ;
 wire \cla/_0555_ ;
 wire \cla/_0556_ ;
 wire \cla/_0557_ ;
 wire \cla/_0558_ ;
 wire \cla/_0559_ ;
 wire \cla/_0560_ ;
 wire \cla/_0561_ ;
 wire \cla/_0562_ ;
 wire \cla/_0563_ ;
 wire \cla/_0564_ ;
 wire \cla/_0565_ ;
 wire \cla/_0566_ ;
 wire \cla/_0567_ ;
 wire \cla/_0568_ ;
 wire \cla/_0569_ ;
 wire \cla/_0570_ ;
 wire \cla/_0571_ ;
 wire \cla/_0572_ ;
 wire \cla/_0573_ ;
 wire \cla/_0574_ ;
 wire \cla/_0575_ ;
 wire \cla/_0576_ ;
 wire \cla/_0577_ ;
 wire \cla/_0578_ ;
 wire \cla/_0579_ ;
 wire \cla/_0580_ ;
 wire \cla/_0581_ ;
 wire \cla/_0582_ ;
 wire \cla/_0583_ ;
 wire \cla/_0584_ ;
 wire \cla/_0585_ ;
 wire \cla/_0586_ ;
 wire \cla/_0587_ ;
 wire \cla/_0588_ ;
 wire \cla/_0589_ ;
 wire \cla/_0590_ ;
 wire \cla/_0591_ ;
 wire \cla/_0592_ ;
 wire \cla/_0593_ ;
 wire \cla/_0594_ ;
 wire \cla/_0595_ ;
 wire \cla/_0596_ ;
 wire \cla/_0597_ ;
 wire \cla/_0598_ ;
 wire \cla/_0599_ ;
 wire \cla/_0600_ ;
 wire \cla/_0601_ ;
 wire \cla/_0602_ ;
 wire \cla/_0603_ ;
 wire \cla/_0604_ ;
 wire \cla/_0605_ ;
 wire \cla/_0606_ ;
 wire \cla/_0607_ ;
 wire \cla/_0608_ ;
 wire \cla/_0609_ ;
 wire \cla/_0610_ ;
 wire \cla/_0611_ ;
 wire \cla/_0612_ ;
 wire \cla/_0613_ ;
 wire \cla/_0614_ ;
 wire \cla/_0615_ ;
 wire \cla/_0616_ ;
 wire \cla/_0617_ ;
 wire \cla/_0618_ ;
 wire \cla/_0619_ ;
 wire \cla/_0620_ ;
 wire \cla/_0621_ ;
 wire \cla/_0622_ ;
 wire \cla/_0623_ ;
 wire \cla/_0624_ ;
 wire \cla/_0625_ ;
 wire \cla/_0626_ ;
 wire \cla/_0627_ ;
 wire \cla/_0628_ ;
 wire \cla/_0629_ ;
 wire \cla/_0630_ ;
 wire \cla/_0631_ ;
 wire \cla/_0632_ ;
 wire \cla/_0633_ ;
 wire \cla/_0634_ ;
 wire \cla/_0635_ ;
 wire \cla/_0636_ ;
 wire \cla/_0637_ ;
 wire \cla/_0638_ ;
 wire \cla/_0639_ ;
 wire \cla/_0640_ ;
 wire \cla/_0641_ ;
 wire \cla/_0642_ ;
 wire \cla/_0643_ ;
 wire \cla/_0644_ ;
 wire \cla/_0645_ ;
 wire \cla/_0646_ ;
 wire \cla/_0647_ ;
 wire \cla/_0648_ ;
 wire \cla/_0649_ ;
 wire \cla/_0650_ ;
 wire \cla/_0651_ ;
 wire \cla/_0652_ ;
 wire \cla/_0653_ ;
 wire \cla/_0654_ ;
 wire \cla/_0655_ ;
 wire \cla/_0656_ ;
 wire \cla/_0657_ ;
 wire \cla/_0658_ ;
 wire \cla/_0659_ ;
 wire \cla/_0660_ ;
 wire \cla/_0661_ ;
 wire \cla/_0662_ ;
 wire \cla/_0663_ ;
 wire \cla/_0664_ ;
 wire \cla/_0665_ ;
 wire \cla/_0666_ ;
 wire \cla/_0667_ ;
 wire \cla/_0668_ ;
 wire \cla/_0669_ ;
 wire \cla/_0670_ ;
 wire \cla/_0671_ ;
 wire \cla/_0672_ ;
 wire \cla/_0673_ ;
 wire \cla/_0674_ ;
 wire \cla/_0675_ ;
 wire \cla/_0676_ ;
 wire \cla/_0677_ ;
 wire \cla/_0678_ ;
 wire \cla/_0679_ ;
 wire \cla/_0680_ ;
 wire \cla/_0681_ ;
 wire \cla/_0682_ ;
 wire \cla/_0683_ ;
 wire \cla/generate_adder_modules[0].fa_i._2_ ;
 wire \cla/generate_adder_modules[10].fa_i.s ;
 wire \cla/generate_adder_modules[11].fa_i.s ;
 wire \cla/generate_adder_modules[12].fa_i.s ;
 wire \cla/generate_adder_modules[13].fa_i.s ;
 wire \cla/generate_adder_modules[14].fa_i.s ;
 wire \cla/generate_adder_modules[15].fa_i.s ;
 wire \cla/generate_adder_modules[16].fa_i.s ;
 wire \cla/generate_adder_modules[17].fa_i.s ;
 wire \cla/generate_adder_modules[18].fa_i.s ;
 wire \cla/generate_adder_modules[19].fa_i.s ;
 wire \cla/generate_adder_modules[1].fa_i.s ;
 wire \cla/generate_adder_modules[20].fa_i.s ;
 wire \cla/generate_adder_modules[21].fa_i.s ;
 wire \cla/generate_adder_modules[22].fa_i.s ;
 wire \cla/generate_adder_modules[23].fa_i.s ;
 wire \cla/generate_adder_modules[2].fa_i.s ;
 wire \cla/generate_adder_modules[3].fa_i.s ;
 wire \cla/generate_adder_modules[4].fa_i.s ;
 wire \cla/generate_adder_modules[5].fa_i.s ;
 wire \cla/generate_adder_modules[6].fa_i.s ;
 wire \cla/generate_adder_modules[7].fa_i.s ;
 wire \cla/generate_adder_modules[8].fa_i.s ;
 wire \cla/generate_adder_modules[9].fa_i.s ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_1 _0760_ (.A(rst_n),
    .X(_0070_));
 sg13g2_buf_1 _0761_ (.A(_0070_),
    .X(_0071_));
 sg13g2_buf_1 _0762_ (.A(uio_in[3]),
    .X(_0072_));
 sg13g2_buf_2 _0763_ (.A(\io_sd.input_index[3] ),
    .X(_0073_));
 sg13g2_buf_1 _0764_ (.A(\io_sd.input_index[4] ),
    .X(_0074_));
 sg13g2_nor2_2 _0765_ (.A(_0073_),
    .B(_0074_),
    .Y(_0075_));
 sg13g2_nand2b_1 _0766_ (.Y(_0076_),
    .B(_0075_),
    .A_N(\io_sd.input_index[5] ));
 sg13g2_buf_1 _0767_ (.A(_0073_),
    .X(_0077_));
 sg13g2_nor3_1 _0768_ (.A(net42),
    .B(\io_sd.input_index[5] ),
    .C(net58),
    .Y(_0078_));
 sg13g2_and2_1 _0769_ (.A(\io_sd._068_ ),
    .B(_0078_),
    .X(_0079_));
 sg13g2_a21oi_1 _0770_ (.A1(\io_sd._092_ ),
    .A2(_0076_),
    .Y(_0080_),
    .B1(_0079_));
 sg13g2_buf_1 _0771_ (.A(\io_sd.output_index[4] ),
    .X(_0081_));
 sg13g2_buf_1 _0772_ (.A(_0081_),
    .X(_0082_));
 sg13g2_buf_1 _0773_ (.A(\io_sd.output_index[3] ),
    .X(_0083_));
 sg13g2_buf_1 _0774_ (.A(_0083_),
    .X(_0084_));
 sg13g2_nor3_1 _0775_ (.A(\io_sd.output_index[5] ),
    .B(_0082_),
    .C(net40),
    .Y(_0085_));
 sg13g2_nand3b_1 _0776_ (.B(\io_sd._092_ ),
    .C(net60),
    .Y(_0086_),
    .A_N(_0085_));
 sg13g2_o21ai_1 _0777_ (.B1(_0086_),
    .Y(_0087_),
    .A1(net60),
    .A2(_0080_));
 sg13g2_and2_1 _0778_ (.A(_0071_),
    .B(_0087_),
    .X(_0001_));
 sg13g2_and2_1 _0779_ (.A(net60),
    .B(_0085_),
    .X(_0088_));
 sg13g2_o21ai_1 _0780_ (.B1(\io_sd._068_ ),
    .Y(_0089_),
    .A1(net60),
    .A2(_0076_));
 sg13g2_buf_1 _0781_ (.A(_0070_),
    .X(_0090_));
 sg13g2_o21ai_1 _0782_ (.B1(net57),
    .Y(_0000_),
    .A1(_0088_),
    .A2(_0089_));
 sg13g2_buf_8 _0783_ (.A(uio_in[2]),
    .X(_0091_));
 sg13g2_inv_2 _0784_ (.Y(_0092_),
    .A(_0091_));
 sg13g2_buf_1 _0785_ (.A(_0092_),
    .X(_0093_));
 sg13g2_inv_1 _0786_ (.Y(_0094_),
    .A(\io_sd._052_[9] ));
 sg13g2_nor2_2 _0787_ (.A(net39),
    .B(_0094_),
    .Y(\rca.generate_adder_modules[9].fa.a ));
 sg13g2_inv_1 _0788_ (.Y(_0095_),
    .A(\io_sd._053_[9] ));
 sg13g2_nor2_2 _0789_ (.A(net39),
    .B(_0095_),
    .Y(\rca.generate_adder_modules[9].fa.b ));
 sg13g2_buf_1 _0790_ (.A(_0091_),
    .X(_0096_));
 sg13g2_buf_1 _0791_ (.A(_0096_),
    .X(_0097_));
 sg13g2_buf_1 _0792_ (.A(net38),
    .X(_0098_));
 sg13g2_buf_1 _0793_ (.A(\io_sd._052_[8] ),
    .X(_0099_));
 sg13g2_and2_1 _0794_ (.A(net31),
    .B(net55),
    .X(\rca.generate_adder_modules[8].fa.a ));
 sg13g2_buf_1 _0795_ (.A(\io_sd._053_[8] ),
    .X(_0100_));
 sg13g2_and2_1 _0796_ (.A(net31),
    .B(net54),
    .X(\rca.generate_adder_modules[8].fa.b ));
 sg13g2_and2_1 _0797_ (.A(net56),
    .B(\io_sd._052_[7] ),
    .X(\rca.generate_adder_modules[7].fa.a ));
 sg13g2_buf_8 _0798_ (.A(\io_sd._053_[7] ),
    .X(_0101_));
 sg13g2_and2_1 _0799_ (.A(net31),
    .B(_0101_),
    .X(\rca.generate_adder_modules[7].fa.b ));
 sg13g2_buf_2 _0800_ (.A(\io_sd._052_[6] ),
    .X(_0102_));
 sg13g2_and2_1 _0801_ (.A(net31),
    .B(_0102_),
    .X(\rca.generate_adder_modules[6].fa.a ));
 sg13g2_buf_2 _0802_ (.A(\io_sd._053_[6] ),
    .X(_0103_));
 sg13g2_and2_1 _0803_ (.A(net31),
    .B(_0103_),
    .X(\rca.generate_adder_modules[6].fa.b ));
 sg13g2_buf_2 _0804_ (.A(\io_sd._052_[5] ),
    .X(_0104_));
 sg13g2_and2_1 _0805_ (.A(net31),
    .B(_0104_),
    .X(\rca.generate_adder_modules[5].fa.a ));
 sg13g2_buf_2 _0806_ (.A(\io_sd._053_[5] ),
    .X(_0105_));
 sg13g2_and2_1 _0807_ (.A(net31),
    .B(_0105_),
    .X(\rca.generate_adder_modules[5].fa.b ));
 sg13g2_and2_1 _0808_ (.A(_0098_),
    .B(\io_sd._052_[4] ),
    .X(\rca.generate_adder_modules[4].fa.a ));
 sg13g2_and2_1 _0809_ (.A(_0098_),
    .B(\io_sd._053_[4] ),
    .X(\rca.generate_adder_modules[4].fa.b ));
 sg13g2_and2_1 _0810_ (.A(net31),
    .B(\io_sd._052_[3] ),
    .X(\rca.generate_adder_modules[3].fa.a ));
 sg13g2_buf_2 _0811_ (.A(\io_sd._052_[2] ),
    .X(_0106_));
 sg13g2_inv_1 _0812_ (.Y(_0107_),
    .A(_0106_));
 sg13g2_nor2_1 _0813_ (.A(net39),
    .B(_0107_),
    .Y(\rca.generate_adder_modules[2].fa.a ));
 sg13g2_buf_2 _0814_ (.A(\io_sd._053_[2] ),
    .X(_0108_));
 sg13g2_inv_1 _0815_ (.Y(_0109_),
    .A(_0108_));
 sg13g2_nor2_1 _0816_ (.A(_0093_),
    .B(_0109_),
    .Y(\rca.generate_adder_modules[2].fa.b ));
 sg13g2_buf_1 _0817_ (.A(_0097_),
    .X(_0110_));
 sg13g2_and2_1 _0818_ (.A(_0110_),
    .B(\io_sd._052_[1] ),
    .X(\rca.generate_adder_modules[1].fa.a ));
 sg13g2_buf_2 _0819_ (.A(\io_sd._053_[0] ),
    .X(_0111_));
 sg13g2_and2_1 _0820_ (.A(_0110_),
    .B(_0111_),
    .X(\rca.generate_adder_modules[0].fa.b ));
 sg13g2_and2_1 _0821_ (.A(net30),
    .B(\io_sd._052_[17] ),
    .X(\rca.generate_adder_modules[17].fa.a ));
 sg13g2_and2_1 _0822_ (.A(net30),
    .B(\io_sd._053_[17] ),
    .X(\rca.generate_adder_modules[17].fa.b ));
 sg13g2_buf_1 _0823_ (.A(\io_sd._052_[16] ),
    .X(_0112_));
 sg13g2_and2_1 _0824_ (.A(net30),
    .B(net53),
    .X(\rca.generate_adder_modules[16].fa.a ));
 sg13g2_buf_2 _0825_ (.A(\io_sd._053_[16] ),
    .X(_0113_));
 sg13g2_and2_1 _0826_ (.A(net30),
    .B(_0113_),
    .X(\rca.generate_adder_modules[16].fa.b ));
 sg13g2_buf_2 _0827_ (.A(\io_sd._052_[15] ),
    .X(_0114_));
 sg13g2_and2_2 _0828_ (.A(_0091_),
    .B(_0114_),
    .X(\rca.generate_adder_modules[15].fa.a ));
 sg13g2_buf_2 _0829_ (.A(\io_sd._053_[15] ),
    .X(_0115_));
 sg13g2_and2_1 _0830_ (.A(net30),
    .B(_0115_),
    .X(\rca.generate_adder_modules[15].fa.b ));
 sg13g2_buf_2 _0831_ (.A(\io_sd._052_[14] ),
    .X(_0116_));
 sg13g2_and2_1 _0832_ (.A(net30),
    .B(_0116_),
    .X(\rca.generate_adder_modules[14].fa.a ));
 sg13g2_buf_2 _0833_ (.A(\io_sd._053_[14] ),
    .X(_0117_));
 sg13g2_and2_1 _0834_ (.A(net30),
    .B(_0117_),
    .X(\rca.generate_adder_modules[14].fa.b ));
 sg13g2_buf_2 _0835_ (.A(\io_sd._052_[13] ),
    .X(_0118_));
 sg13g2_inv_1 _0836_ (.Y(_0119_),
    .A(_0118_));
 sg13g2_nor2_1 _0837_ (.A(net39),
    .B(_0119_),
    .Y(\rca.generate_adder_modules[13].fa.a ));
 sg13g2_buf_2 _0838_ (.A(\io_sd._053_[13] ),
    .X(_0120_));
 sg13g2_inv_1 _0839_ (.Y(_0121_),
    .A(_0120_));
 sg13g2_nor2_2 _0840_ (.A(net39),
    .B(_0121_),
    .Y(\rca.generate_adder_modules[13].fa.b ));
 sg13g2_and2_1 _0841_ (.A(net30),
    .B(\io_sd._052_[12] ),
    .X(\rca.generate_adder_modules[12].fa.a ));
 sg13g2_buf_1 _0842_ (.A(net38),
    .X(_0122_));
 sg13g2_and2_2 _0843_ (.A(net29),
    .B(\io_sd._053_[12] ),
    .X(\rca.generate_adder_modules[12].fa.b ));
 sg13g2_buf_2 _0844_ (.A(\io_sd._052_[11] ),
    .X(_0123_));
 sg13g2_and2_1 _0845_ (.A(net29),
    .B(_0123_),
    .X(\rca.generate_adder_modules[11].fa.a ));
 sg13g2_buf_2 _0846_ (.A(\io_sd._053_[11] ),
    .X(_0124_));
 sg13g2_and2_1 _0847_ (.A(net29),
    .B(_0124_),
    .X(\rca.generate_adder_modules[11].fa.b ));
 sg13g2_buf_1 _0848_ (.A(\io_sd._052_[10] ),
    .X(_0125_));
 sg13g2_and2_1 _0849_ (.A(_0122_),
    .B(net52),
    .X(\rca.generate_adder_modules[10].fa.a ));
 sg13g2_buf_1 _0850_ (.A(\io_sd._053_[10] ),
    .X(_0126_));
 sg13g2_and2_1 _0851_ (.A(_0122_),
    .B(_0126_),
    .X(\rca.generate_adder_modules[10].fa.b ));
 sg13g2_inv_1 _0852_ (.Y(_0127_),
    .A(\io_sd._052_[18] ));
 sg13g2_nor2_2 _0853_ (.A(_0092_),
    .B(_0127_),
    .Y(\rca.generate_adder_modules[18].fa.a ));
 sg13g2_buf_1 _0854_ (.A(\io_sd._053_[18] ),
    .X(_0128_));
 sg13g2_inv_1 _0855_ (.Y(_0129_),
    .A(_0128_));
 sg13g2_nor2_1 _0856_ (.A(net39),
    .B(_0129_),
    .Y(\rca.generate_adder_modules[18].fa.b ));
 sg13g2_and2_1 _0857_ (.A(net29),
    .B(\io_sd._052_[19] ),
    .X(\rca.generate_adder_modules[19].fa.a ));
 sg13g2_and2_1 _0858_ (.A(net29),
    .B(\io_sd._053_[19] ),
    .X(\rca.generate_adder_modules[19].fa.b ));
 sg13g2_buf_1 _0859_ (.A(\io_sd._052_[20] ),
    .X(_0130_));
 sg13g2_and2_1 _0860_ (.A(net29),
    .B(_0130_),
    .X(\rca.generate_adder_modules[20].fa.a ));
 sg13g2_buf_1 _0861_ (.A(\io_sd._053_[20] ),
    .X(_0131_));
 sg13g2_and2_1 _0862_ (.A(net29),
    .B(_0131_),
    .X(\rca.generate_adder_modules[20].fa.b ));
 sg13g2_buf_2 _0863_ (.A(\io_sd._052_[21] ),
    .X(_0132_));
 sg13g2_and2_1 _0864_ (.A(net29),
    .B(_0132_),
    .X(\rca.generate_adder_modules[21].fa.a ));
 sg13g2_buf_2 _0865_ (.A(\io_sd._053_[21] ),
    .X(_0133_));
 sg13g2_and2_1 _0866_ (.A(net38),
    .B(_0133_),
    .X(\rca.generate_adder_modules[21].fa.b ));
 sg13g2_buf_2 _0867_ (.A(\io_sd._052_[22] ),
    .X(_0134_));
 sg13g2_and2_1 _0868_ (.A(net38),
    .B(_0134_),
    .X(\rca.generate_adder_modules[22].fa.a ));
 sg13g2_buf_2 _0869_ (.A(\io_sd._053_[22] ),
    .X(_0135_));
 sg13g2_and2_1 _0870_ (.A(net38),
    .B(_0135_),
    .X(\rca.generate_adder_modules[22].fa.b ));
 sg13g2_and2_1 _0871_ (.A(net38),
    .B(\io_sd._052_[23] ),
    .X(\rca.generate_adder_modules[23].fa.a ));
 sg13g2_and2_1 _0872_ (.A(net38),
    .B(\io_sd._053_[23] ),
    .X(\rca.generate_adder_modules[23].fa.b ));
 sg13g2_buf_2 _0873_ (.A(\io_sd._052_[0] ),
    .X(_0136_));
 sg13g2_inv_2 _0874_ (.Y(_0137_),
    .A(net60));
 sg13g2_nand2_2 _0875_ (.Y(_0138_),
    .A(\io_sd._068_ ),
    .B(_0137_));
 sg13g2_buf_1 _0876_ (.A(\io_sd._210_[0] ),
    .X(_0139_));
 sg13g2_buf_1 _0877_ (.A(_0002_),
    .X(_0140_));
 sg13g2_nand3_1 _0878_ (.B(net47),
    .C(_0075_),
    .A(_0139_),
    .Y(_0141_));
 sg13g2_or2_1 _0879_ (.X(_0142_),
    .B(_0141_),
    .A(_0138_));
 sg13g2_buf_1 _0880_ (.A(_0139_),
    .X(_0143_));
 sg13g2_inv_1 _0881_ (.Y(_0144_),
    .A(net42));
 sg13g2_nor3_1 _0882_ (.A(_0143_),
    .B(_0144_),
    .C(_0005_),
    .Y(_0145_));
 sg13g2_a21oi_1 _0883_ (.A1(_0143_),
    .A2(_0144_),
    .Y(_0146_),
    .B1(_0145_));
 sg13g2_nand2_1 _0884_ (.Y(_0147_),
    .A(net47),
    .B(net1));
 sg13g2_nor3_1 _0885_ (.A(net58),
    .B(_0146_),
    .C(_0147_),
    .Y(_0148_));
 sg13g2_nor2b_1 _0886_ (.A(_0072_),
    .B_N(\io_sd._068_ ),
    .Y(_0149_));
 sg13g2_buf_1 _0887_ (.A(_0149_),
    .X(_0150_));
 sg13g2_a22oi_1 _0888_ (.Y(_0151_),
    .B1(_0148_),
    .B2(_0150_),
    .A2(_0142_),
    .A1(_0136_));
 sg13g2_nor2b_1 _0889_ (.A(_0151_),
    .B_N(_0090_),
    .Y(_0006_));
 sg13g2_mux2_1 _0890_ (.A0(net2),
    .A1(net3),
    .S(net37),
    .X(_0152_));
 sg13g2_nor2b_2 _0891_ (.A(net58),
    .B_N(_0073_),
    .Y(_0153_));
 sg13g2_nor2_1 _0892_ (.A(\io_sd._210_[0] ),
    .B(_0073_),
    .Y(_0154_));
 sg13g2_a22oi_1 _0893_ (.Y(_0155_),
    .B1(_0154_),
    .B2(net58),
    .A2(_0153_),
    .A1(\io_sd._210_[0] ));
 sg13g2_nand2b_1 _0894_ (.Y(_0156_),
    .B(net47),
    .A_N(_0155_));
 sg13g2_or2_1 _0895_ (.X(_0157_),
    .B(_0156_),
    .A(_0138_));
 sg13g2_buf_1 _0896_ (.A(_0157_),
    .X(_0158_));
 sg13g2_mux2_1 _0897_ (.A0(_0152_),
    .A1(net52),
    .S(net22),
    .X(_0159_));
 sg13g2_and2_1 _0898_ (.A(net59),
    .B(_0159_),
    .X(_0007_));
 sg13g2_mux2_1 _0899_ (.A0(net3),
    .A1(net4),
    .S(net48),
    .X(_0160_));
 sg13g2_mux2_1 _0900_ (.A0(_0160_),
    .A1(_0123_),
    .S(net22),
    .X(_0161_));
 sg13g2_and2_1 _0901_ (.A(net59),
    .B(_0161_),
    .X(_0008_));
 sg13g2_mux2_1 _0902_ (.A0(net4),
    .A1(net5),
    .S(net37),
    .X(_0162_));
 sg13g2_mux2_1 _0903_ (.A0(_0162_),
    .A1(\io_sd._052_[12] ),
    .S(net22),
    .X(_0163_));
 sg13g2_and2_1 _0904_ (.A(net59),
    .B(_0163_),
    .X(_0009_));
 sg13g2_mux2_2 _0905_ (.A0(net5),
    .A1(net6),
    .S(net48),
    .X(_0164_));
 sg13g2_nor2_1 _0906_ (.A(net22),
    .B(_0164_),
    .Y(_0165_));
 sg13g2_a21oi_1 _0907_ (.A1(_0119_),
    .A2(net22),
    .Y(_0166_),
    .B1(_0165_));
 sg13g2_and2_1 _0908_ (.A(net59),
    .B(_0166_),
    .X(_0010_));
 sg13g2_mux2_1 _0909_ (.A0(net6),
    .A1(net7),
    .S(net48),
    .X(_0167_));
 sg13g2_mux2_1 _0910_ (.A0(_0167_),
    .A1(_0116_),
    .S(net22),
    .X(_0168_));
 sg13g2_and2_1 _0911_ (.A(net59),
    .B(_0168_),
    .X(_0011_));
 sg13g2_mux2_1 _0912_ (.A0(net7),
    .A1(net8),
    .S(net48),
    .X(_0169_));
 sg13g2_mux2_1 _0913_ (.A0(_0169_),
    .A1(_0114_),
    .S(net22),
    .X(_0170_));
 sg13g2_and2_1 _0914_ (.A(net59),
    .B(_0170_),
    .X(_0012_));
 sg13g2_buf_1 _0915_ (.A(_0070_),
    .X(_0171_));
 sg13g2_nand2_1 _0916_ (.Y(_0172_),
    .A(net58),
    .B(net47));
 sg13g2_nor2b_1 _0917_ (.A(_0005_),
    .B_N(net1),
    .Y(_0173_));
 sg13g2_nor2b_1 _0918_ (.A(net42),
    .B_N(net8),
    .Y(_0174_));
 sg13g2_a21oi_1 _0919_ (.A1(net42),
    .A2(_0173_),
    .Y(_0175_),
    .B1(_0174_));
 sg13g2_nand3b_1 _0920_ (.B(_0173_),
    .C(net48),
    .Y(_0176_),
    .A_N(_0077_));
 sg13g2_o21ai_1 _0921_ (.B1(_0176_),
    .Y(_0177_),
    .A1(net37),
    .A2(_0175_));
 sg13g2_nand2b_1 _0922_ (.Y(_0178_),
    .B(_0177_),
    .A_N(_0172_));
 sg13g2_nand3_1 _0923_ (.B(_0140_),
    .C(_0149_),
    .A(net58),
    .Y(_0179_));
 sg13g2_o21ai_1 _0924_ (.B1(_0112_),
    .Y(_0180_),
    .A1(net42),
    .A2(_0179_));
 sg13g2_o21ai_1 _0925_ (.B1(_0180_),
    .Y(_0181_),
    .A1(_0138_),
    .A2(_0178_));
 sg13g2_and2_1 _0926_ (.A(net46),
    .B(_0181_),
    .X(_0013_));
 sg13g2_mux2_2 _0927_ (.A0(net1),
    .A1(net2),
    .S(net48),
    .X(_0182_));
 sg13g2_xnor2_1 _0928_ (.Y(_0183_),
    .A(net48),
    .B(_0073_));
 sg13g2_nor2_1 _0929_ (.A(_0179_),
    .B(_0183_),
    .Y(_0184_));
 sg13g2_buf_2 _0930_ (.A(_0184_),
    .X(_0185_));
 sg13g2_mux2_1 _0931_ (.A0(\io_sd._052_[17] ),
    .A1(_0182_),
    .S(_0185_),
    .X(_0186_));
 sg13g2_and2_1 _0932_ (.A(net46),
    .B(_0186_),
    .X(_0014_));
 sg13g2_nand2_1 _0933_ (.Y(_0187_),
    .A(_0152_),
    .B(_0185_));
 sg13g2_o21ai_1 _0934_ (.B1(_0187_),
    .Y(_0188_),
    .A1(_0127_),
    .A2(_0185_));
 sg13g2_and2_1 _0935_ (.A(net46),
    .B(_0188_),
    .X(_0015_));
 sg13g2_mux2_1 _0936_ (.A0(\io_sd._052_[19] ),
    .A1(_0160_),
    .S(_0185_),
    .X(_0189_));
 sg13g2_and2_1 _0937_ (.A(net46),
    .B(_0189_),
    .X(_0016_));
 sg13g2_nor2_2 _0938_ (.A(_0005_),
    .B(_0141_),
    .Y(_0190_));
 sg13g2_nand2_2 _0939_ (.Y(_0191_),
    .A(net47),
    .B(_0153_));
 sg13g2_nor2_2 _0940_ (.A(net48),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_and2_1 _0941_ (.A(_0182_),
    .B(_0192_),
    .X(_0193_));
 sg13g2_a21o_1 _0942_ (.A2(_0190_),
    .A1(net2),
    .B1(_0193_),
    .X(_0194_));
 sg13g2_o21ai_1 _0943_ (.B1(net36),
    .Y(_0195_),
    .A1(_0190_),
    .A2(_0192_));
 sg13g2_buf_2 _0944_ (.A(_0195_),
    .X(_0196_));
 sg13g2_a22oi_1 _0945_ (.Y(_0197_),
    .B1(_0196_),
    .B2(\io_sd._052_[1] ),
    .A2(_0194_),
    .A1(net36));
 sg13g2_nor2b_1 _0946_ (.A(_0197_),
    .B_N(net57),
    .Y(_0017_));
 sg13g2_mux2_1 _0947_ (.A0(net50),
    .A1(_0162_),
    .S(_0185_),
    .X(_0198_));
 sg13g2_and2_1 _0948_ (.A(net46),
    .B(_0198_),
    .X(_0018_));
 sg13g2_mux2_1 _0949_ (.A0(_0132_),
    .A1(_0164_),
    .S(_0185_),
    .X(_0199_));
 sg13g2_and2_1 _0950_ (.A(net46),
    .B(_0199_),
    .X(_0019_));
 sg13g2_mux2_1 _0951_ (.A0(_0134_),
    .A1(_0167_),
    .S(_0185_),
    .X(_0200_));
 sg13g2_and2_1 _0952_ (.A(net46),
    .B(_0200_),
    .X(_0020_));
 sg13g2_mux2_1 _0953_ (.A0(\io_sd._052_[23] ),
    .A1(_0169_),
    .S(_0185_),
    .X(_0201_));
 sg13g2_and2_1 _0954_ (.A(net46),
    .B(_0201_),
    .X(_0021_));
 sg13g2_and2_1 _0955_ (.A(net3),
    .B(_0190_),
    .X(_0202_));
 sg13g2_a21o_1 _0956_ (.A2(_0192_),
    .A1(net2),
    .B1(_0202_),
    .X(_0203_));
 sg13g2_a22oi_1 _0957_ (.Y(_0204_),
    .B1(_0203_),
    .B2(net36),
    .A2(_0196_),
    .A1(_0106_));
 sg13g2_nor2b_1 _0958_ (.A(_0204_),
    .B_N(net57),
    .Y(_0022_));
 sg13g2_and2_1 _0959_ (.A(_0160_),
    .B(_0192_),
    .X(_0205_));
 sg13g2_a21o_1 _0960_ (.A2(_0190_),
    .A1(net4),
    .B1(_0205_),
    .X(_0206_));
 sg13g2_a22oi_1 _0961_ (.Y(_0207_),
    .B1(_0206_),
    .B2(net36),
    .A2(_0196_),
    .A1(\io_sd._052_[3] ));
 sg13g2_nor2b_1 _0962_ (.A(_0207_),
    .B_N(net57),
    .Y(_0023_));
 sg13g2_and2_1 _0963_ (.A(net5),
    .B(_0190_),
    .X(_0208_));
 sg13g2_a21o_1 _0964_ (.A2(_0192_),
    .A1(net4),
    .B1(_0208_),
    .X(_0209_));
 sg13g2_a22oi_1 _0965_ (.Y(_0210_),
    .B1(_0209_),
    .B2(net36),
    .A2(_0196_),
    .A1(\io_sd._052_[4] ));
 sg13g2_nor2b_1 _0966_ (.A(_0210_),
    .B_N(net57),
    .Y(_0024_));
 sg13g2_and2_1 _0967_ (.A(_0164_),
    .B(_0192_),
    .X(_0211_));
 sg13g2_a21o_1 _0968_ (.A2(_0190_),
    .A1(net6),
    .B1(_0211_),
    .X(_0212_));
 sg13g2_a22oi_1 _0969_ (.Y(_0213_),
    .B1(_0212_),
    .B2(net36),
    .A2(_0196_),
    .A1(_0104_));
 sg13g2_nor2b_1 _0970_ (.A(_0213_),
    .B_N(net57),
    .Y(_0025_));
 sg13g2_and2_1 _0971_ (.A(_0167_),
    .B(_0192_),
    .X(_0214_));
 sg13g2_a21o_1 _0972_ (.A2(_0190_),
    .A1(net7),
    .B1(_0214_),
    .X(_0215_));
 sg13g2_a22oi_1 _0973_ (.Y(_0216_),
    .B1(_0215_),
    .B2(net36),
    .A2(_0196_),
    .A1(_0102_));
 sg13g2_buf_1 _0974_ (.A(_0070_),
    .X(_0217_));
 sg13g2_buf_1 _0975_ (.A(net45),
    .X(_0218_));
 sg13g2_nor2b_1 _0976_ (.A(_0216_),
    .B_N(net35),
    .Y(_0026_));
 sg13g2_nand4_1 _0977_ (.B(net47),
    .C(net8),
    .A(net37),
    .Y(_0219_),
    .D(_0075_));
 sg13g2_o21ai_1 _0978_ (.B1(_0219_),
    .Y(_0220_),
    .A1(net37),
    .A2(_0191_));
 sg13g2_and2_1 _0979_ (.A(_0169_),
    .B(_0220_),
    .X(_0221_));
 sg13g2_a22oi_1 _0980_ (.Y(_0222_),
    .B1(_0221_),
    .B2(net36),
    .A2(_0196_),
    .A1(\io_sd._052_[7] ));
 sg13g2_nor2b_1 _0981_ (.A(_0222_),
    .B_N(net35),
    .Y(_0027_));
 sg13g2_nor2b_1 _0982_ (.A(_0073_),
    .B_N(net58),
    .Y(_0223_));
 sg13g2_a22oi_1 _0983_ (.Y(_0224_),
    .B1(_0223_),
    .B2(_0173_),
    .A2(_0153_),
    .A1(net8));
 sg13g2_nand3_1 _0984_ (.B(_0153_),
    .C(_0173_),
    .A(net37),
    .Y(_0225_));
 sg13g2_o21ai_1 _0985_ (.B1(_0225_),
    .Y(_0226_),
    .A1(net37),
    .A2(_0224_));
 sg13g2_nand2_1 _0986_ (.Y(_0227_),
    .A(net47),
    .B(_0226_));
 sg13g2_o21ai_1 _0987_ (.B1(_0099_),
    .Y(_0228_),
    .A1(_0138_),
    .A2(_0191_));
 sg13g2_o21ai_1 _0988_ (.B1(_0228_),
    .Y(_0229_),
    .A1(_0138_),
    .A2(_0227_));
 sg13g2_and2_1 _0989_ (.A(_0171_),
    .B(_0229_),
    .X(_0028_));
 sg13g2_nor2_1 _0990_ (.A(net22),
    .B(_0182_),
    .Y(_0230_));
 sg13g2_a21oi_1 _0991_ (.A1(_0094_),
    .A2(_0158_),
    .Y(_0231_),
    .B1(_0230_));
 sg13g2_and2_1 _0992_ (.A(_0171_),
    .B(_0231_),
    .X(_0029_));
 sg13g2_nor2b_2 _0993_ (.A(_0072_),
    .B_N(\io_sd._092_ ),
    .Y(_0232_));
 sg13g2_buf_1 _0994_ (.A(_0232_),
    .X(_0233_));
 sg13g2_nand2b_1 _0995_ (.Y(_0234_),
    .B(_0233_),
    .A_N(_0141_));
 sg13g2_a22oi_1 _0996_ (.Y(_0235_),
    .B1(_0234_),
    .B2(_0111_),
    .A2(net34),
    .A1(_0148_));
 sg13g2_nor2b_1 _0997_ (.A(_0235_),
    .B_N(net35),
    .Y(_0030_));
 sg13g2_buf_1 _0998_ (.A(_0070_),
    .X(_0236_));
 sg13g2_nand2b_1 _0999_ (.Y(_0237_),
    .B(_0232_),
    .A_N(_0156_));
 sg13g2_buf_1 _1000_ (.A(_0237_),
    .X(_0238_));
 sg13g2_mux2_1 _1001_ (.A0(_0152_),
    .A1(net51),
    .S(net21),
    .X(_0239_));
 sg13g2_and2_1 _1002_ (.A(net44),
    .B(_0239_),
    .X(_0031_));
 sg13g2_mux2_1 _1003_ (.A0(_0160_),
    .A1(_0124_),
    .S(net21),
    .X(_0240_));
 sg13g2_and2_1 _1004_ (.A(net44),
    .B(_0240_),
    .X(_0032_));
 sg13g2_mux2_1 _1005_ (.A0(_0162_),
    .A1(\io_sd._053_[12] ),
    .S(net21),
    .X(_0241_));
 sg13g2_and2_1 _1006_ (.A(net44),
    .B(_0241_),
    .X(_0033_));
 sg13g2_nor2_1 _1007_ (.A(_0164_),
    .B(net21),
    .Y(_0242_));
 sg13g2_a21oi_1 _1008_ (.A1(_0121_),
    .A2(net21),
    .Y(_0243_),
    .B1(_0242_));
 sg13g2_and2_1 _1009_ (.A(_0236_),
    .B(_0243_),
    .X(_0034_));
 sg13g2_mux2_1 _1010_ (.A0(_0167_),
    .A1(_0117_),
    .S(net21),
    .X(_0244_));
 sg13g2_and2_1 _1011_ (.A(net44),
    .B(_0244_),
    .X(_0035_));
 sg13g2_mux2_1 _1012_ (.A0(_0169_),
    .A1(_0115_),
    .S(net21),
    .X(_0245_));
 sg13g2_and2_1 _1013_ (.A(net44),
    .B(_0245_),
    .X(_0036_));
 sg13g2_nand2_1 _1014_ (.Y(_0246_),
    .A(_0137_),
    .B(\io_sd._092_ ));
 sg13g2_nand2b_1 _1015_ (.Y(_0247_),
    .B(_0232_),
    .A_N(_0172_));
 sg13g2_o21ai_1 _1016_ (.B1(_0113_),
    .Y(_0248_),
    .A1(net42),
    .A2(_0247_));
 sg13g2_o21ai_1 _1017_ (.B1(_0248_),
    .Y(_0249_),
    .A1(_0178_),
    .A2(_0246_));
 sg13g2_and2_1 _1018_ (.A(_0236_),
    .B(_0249_),
    .X(_0037_));
 sg13g2_nor2_1 _1019_ (.A(_0183_),
    .B(_0247_),
    .Y(_0250_));
 sg13g2_buf_2 _1020_ (.A(_0250_),
    .X(_0251_));
 sg13g2_mux2_1 _1021_ (.A0(\io_sd._053_[17] ),
    .A1(_0182_),
    .S(_0251_),
    .X(_0252_));
 sg13g2_and2_1 _1022_ (.A(net44),
    .B(_0252_),
    .X(_0038_));
 sg13g2_nand2_1 _1023_ (.Y(_0253_),
    .A(_0152_),
    .B(_0251_));
 sg13g2_o21ai_1 _1024_ (.B1(_0253_),
    .Y(_0254_),
    .A1(_0129_),
    .A2(_0251_));
 sg13g2_and2_1 _1025_ (.A(net44),
    .B(_0254_),
    .X(_0039_));
 sg13g2_mux2_1 _1026_ (.A0(\io_sd._053_[19] ),
    .A1(_0160_),
    .S(_0251_),
    .X(_0255_));
 sg13g2_and2_1 _1027_ (.A(net44),
    .B(_0255_),
    .X(_0040_));
 sg13g2_o21ai_1 _1028_ (.B1(_0233_),
    .Y(_0256_),
    .A1(_0190_),
    .A2(_0192_));
 sg13g2_buf_2 _1029_ (.A(_0256_),
    .X(_0257_));
 sg13g2_a22oi_1 _1030_ (.Y(_0258_),
    .B1(_0257_),
    .B2(\io_sd._053_[1] ),
    .A2(net34),
    .A1(_0194_));
 sg13g2_nor2b_1 _1031_ (.A(_0258_),
    .B_N(_0218_),
    .Y(_0041_));
 sg13g2_mux2_1 _1032_ (.A0(net49),
    .A1(_0162_),
    .S(_0251_),
    .X(_0259_));
 sg13g2_and2_1 _1033_ (.A(net45),
    .B(_0259_),
    .X(_0042_));
 sg13g2_mux2_1 _1034_ (.A0(_0133_),
    .A1(_0164_),
    .S(_0251_),
    .X(_0260_));
 sg13g2_and2_1 _1035_ (.A(net45),
    .B(_0260_),
    .X(_0043_));
 sg13g2_mux2_1 _1036_ (.A0(_0135_),
    .A1(_0167_),
    .S(_0251_),
    .X(_0261_));
 sg13g2_and2_1 _1037_ (.A(net45),
    .B(_0261_),
    .X(_0044_));
 sg13g2_mux2_1 _1038_ (.A0(\io_sd._053_[23] ),
    .A1(_0169_),
    .S(_0251_),
    .X(_0262_));
 sg13g2_and2_1 _1039_ (.A(net45),
    .B(_0262_),
    .X(_0045_));
 sg13g2_a22oi_1 _1040_ (.Y(_0263_),
    .B1(_0257_),
    .B2(_0108_),
    .A2(net34),
    .A1(_0203_));
 sg13g2_nor2b_1 _1041_ (.A(_0263_),
    .B_N(_0218_),
    .Y(_0046_));
 sg13g2_a22oi_1 _1042_ (.Y(_0264_),
    .B1(_0257_),
    .B2(\io_sd._053_[3] ),
    .A2(net34),
    .A1(_0206_));
 sg13g2_nor2b_1 _1043_ (.A(_0264_),
    .B_N(net35),
    .Y(_0047_));
 sg13g2_a22oi_1 _1044_ (.Y(_0265_),
    .B1(_0257_),
    .B2(\io_sd._053_[4] ),
    .A2(net34),
    .A1(_0209_));
 sg13g2_nor2b_1 _1045_ (.A(_0265_),
    .B_N(net35),
    .Y(_0048_));
 sg13g2_a22oi_1 _1046_ (.Y(_0266_),
    .B1(_0257_),
    .B2(_0105_),
    .A2(net34),
    .A1(_0212_));
 sg13g2_nor2b_1 _1047_ (.A(_0266_),
    .B_N(net35),
    .Y(_0049_));
 sg13g2_a22oi_1 _1048_ (.Y(_0267_),
    .B1(_0257_),
    .B2(_0103_),
    .A2(net34),
    .A1(_0215_));
 sg13g2_nor2b_1 _1049_ (.A(_0267_),
    .B_N(net35),
    .Y(_0050_));
 sg13g2_a22oi_1 _1050_ (.Y(_0268_),
    .B1(_0257_),
    .B2(_0101_),
    .A2(net34),
    .A1(_0221_));
 sg13g2_nor2b_1 _1051_ (.A(_0268_),
    .B_N(net35),
    .Y(_0051_));
 sg13g2_o21ai_1 _1052_ (.B1(_0100_),
    .Y(_0269_),
    .A1(_0191_),
    .A2(_0246_));
 sg13g2_o21ai_1 _1053_ (.B1(_0269_),
    .Y(_0270_),
    .A1(_0227_),
    .A2(_0246_));
 sg13g2_and2_1 _1054_ (.A(net45),
    .B(_0270_),
    .X(_0052_));
 sg13g2_nor2_1 _1055_ (.A(_0182_),
    .B(net21),
    .Y(_0271_));
 sg13g2_a21oi_1 _1056_ (.A1(_0095_),
    .A2(_0238_),
    .Y(_0272_),
    .B1(_0271_));
 sg13g2_and2_1 _1057_ (.A(_0217_),
    .B(_0272_),
    .X(_0053_));
 sg13g2_nor2_2 _1058_ (.A(_0150_),
    .B(_0232_),
    .Y(_0273_));
 sg13g2_nor2b_1 _1059_ (.A(net37),
    .B_N(_0217_),
    .Y(_0274_));
 sg13g2_o21ai_1 _1060_ (.B1(_0274_),
    .Y(_0054_),
    .A1(_0076_),
    .A2(_0273_));
 sg13g2_nor3_1 _1061_ (.A(net42),
    .B(_0078_),
    .C(_0273_),
    .Y(_0275_));
 sg13g2_a21oi_1 _1062_ (.A1(net42),
    .A2(_0273_),
    .Y(_0276_),
    .B1(_0275_));
 sg13g2_nor2b_1 _1063_ (.A(_0276_),
    .B_N(net59),
    .Y(_0055_));
 sg13g2_nor2_1 _1064_ (.A(_0077_),
    .B(_0273_),
    .Y(_0277_));
 sg13g2_xnor2_1 _1065_ (.Y(_0278_),
    .A(net58),
    .B(_0277_));
 sg13g2_nand2_1 _1066_ (.Y(_0056_),
    .A(_0090_),
    .B(_0278_));
 sg13g2_a21o_1 _1067_ (.A2(_0075_),
    .A1(_0140_),
    .B1(_0273_),
    .X(_0279_));
 sg13g2_nor3_1 _1068_ (.A(net47),
    .B(_0075_),
    .C(_0273_),
    .Y(_0280_));
 sg13g2_a21oi_1 _1069_ (.A1(\io_sd.input_index[5] ),
    .A2(_0279_),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_nor2b_1 _1070_ (.A(_0281_),
    .B_N(_0071_),
    .Y(_0057_));
 sg13g2_buf_2 _1071_ (.A(\io_sd._209_[0] ),
    .X(_0282_));
 sg13g2_inv_1 _1072_ (.Y(_0283_),
    .A(_0282_));
 sg13g2_buf_1 _1073_ (.A(_0283_),
    .X(_0284_));
 sg13g2_nand3b_1 _1074_ (.B(net57),
    .C(_0284_),
    .Y(_0058_),
    .A_N(_0088_));
 sg13g2_buf_1 _1075_ (.A(_0084_),
    .X(_0285_));
 sg13g2_nor3_1 _1076_ (.A(_0137_),
    .B(_0285_),
    .C(_0085_),
    .Y(_0286_));
 sg13g2_a21o_1 _1077_ (.A2(_0285_),
    .A1(_0137_),
    .B1(_0286_),
    .X(_0287_));
 sg13g2_and2_1 _1078_ (.A(net45),
    .B(_0287_),
    .X(_0059_));
 sg13g2_nor2_1 _1079_ (.A(_0137_),
    .B(net27),
    .Y(_0288_));
 sg13g2_xnor2_1 _1080_ (.Y(_0289_),
    .A(_0082_),
    .B(_0288_));
 sg13g2_nand2_1 _1081_ (.Y(_0060_),
    .A(net57),
    .B(_0289_));
 sg13g2_nor2_1 _1082_ (.A(_0081_),
    .B(_0083_),
    .Y(_0290_));
 sg13g2_a21o_1 _1083_ (.A2(_0290_),
    .A1(_0003_),
    .B1(_0137_),
    .X(_0291_));
 sg13g2_nor3_1 _1084_ (.A(_0137_),
    .B(_0003_),
    .C(_0290_),
    .Y(_0292_));
 sg13g2_a21oi_1 _1085_ (.A1(\io_sd.output_index[5] ),
    .A2(_0291_),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_nor2b_1 _1086_ (.A(_0293_),
    .B_N(net59),
    .Y(_0061_));
 sg13g2_nand2_1 _1087_ (.Y(_0294_),
    .A(net60),
    .B(_0070_));
 sg13g2_or2_1 _1088_ (.X(_0295_),
    .B(_0282_),
    .A(_0083_));
 sg13g2_buf_1 _1089_ (.A(_0295_),
    .X(_0296_));
 sg13g2_nor2_1 _1090_ (.A(_0081_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_xnor2_1 _1091_ (.Y(_0298_),
    .A(_0003_),
    .B(_0297_));
 sg13g2_nor2_2 _1092_ (.A(_0294_),
    .B(_0298_),
    .Y(_0299_));
 sg13g2_nand3_1 _1093_ (.B(_0003_),
    .C(_0290_),
    .A(_0283_),
    .Y(_0300_));
 sg13g2_xnor2_1 _1094_ (.Y(_0301_),
    .A(\io_sd.output_index[5] ),
    .B(_0003_));
 sg13g2_and2_1 _1095_ (.A(_0083_),
    .B(_0282_),
    .X(_0302_));
 sg13g2_buf_2 _1096_ (.A(_0302_),
    .X(_0303_));
 sg13g2_nand3_1 _1097_ (.B(_0301_),
    .C(_0303_),
    .A(_0081_),
    .Y(_0304_));
 sg13g2_and2_1 _1098_ (.A(_0300_),
    .B(_0304_),
    .X(_0305_));
 sg13g2_buf_2 _1099_ (.A(_0305_),
    .X(_0306_));
 sg13g2_buf_1 _1100_ (.A(uio_in[0]),
    .X(_0307_));
 sg13g2_buf_1 _1101_ (.A(_0307_),
    .X(_0308_));
 sg13g2_nand2_1 _1102_ (.Y(_0309_),
    .A(_0108_),
    .B(_0106_));
 sg13g2_a21oi_1 _1103_ (.A1(_0136_),
    .A2(_0111_),
    .Y(_0310_),
    .B1(\io_sd._052_[1] ));
 sg13g2_nand3_1 _1104_ (.B(_0111_),
    .C(\io_sd._052_[1] ),
    .A(_0136_),
    .Y(_0311_));
 sg13g2_a21oi_1 _1105_ (.A1(_0108_),
    .A2(_0106_),
    .Y(_0312_),
    .B1(\io_sd._053_[1] ));
 sg13g2_a22oi_1 _1106_ (.Y(_0313_),
    .B1(_0311_),
    .B2(_0312_),
    .A2(_0310_),
    .A1(_0309_));
 sg13g2_nand2_1 _1107_ (.Y(_0314_),
    .A(\io_sd._053_[4] ),
    .B(\io_sd._052_[4] ));
 sg13g2_nor2_1 _1108_ (.A(\io_sd._053_[3] ),
    .B(\io_sd._052_[3] ),
    .Y(_0315_));
 sg13g2_nor2_1 _1109_ (.A(\io_sd._053_[4] ),
    .B(\io_sd._052_[4] ),
    .Y(_0316_));
 sg13g2_a221oi_1 _1110_ (.B2(_0315_),
    .C1(_0316_),
    .B1(_0314_),
    .A1(_0109_),
    .Y(_0317_),
    .A2(_0107_));
 sg13g2_nand2_1 _1111_ (.Y(_0318_),
    .A(\io_sd._053_[3] ),
    .B(\io_sd._052_[3] ));
 sg13g2_a21oi_1 _1112_ (.A1(_0314_),
    .A2(_0318_),
    .Y(_0319_),
    .B1(_0316_));
 sg13g2_a21o_1 _1113_ (.A2(_0317_),
    .A1(_0313_),
    .B1(_0319_),
    .X(_0320_));
 sg13g2_buf_2 _1114_ (.A(_0320_),
    .X(_0321_));
 sg13g2_xnor2_1 _1115_ (.Y(_0322_),
    .A(_0101_),
    .B(\io_sd._052_[7] ));
 sg13g2_xnor2_1 _1116_ (.Y(_0323_),
    .A(_0103_),
    .B(_0102_));
 sg13g2_xnor2_1 _1117_ (.Y(_0324_),
    .A(_0105_),
    .B(_0104_));
 sg13g2_nor4_2 _1118_ (.A(_0092_),
    .B(_0322_),
    .C(_0323_),
    .Y(_0325_),
    .D(_0324_));
 sg13g2_nor2_1 _1119_ (.A(_0103_),
    .B(_0102_),
    .Y(_0326_));
 sg13g2_a22oi_1 _1120_ (.Y(_0327_),
    .B1(_0102_),
    .B2(_0103_),
    .A2(_0104_),
    .A1(_0105_));
 sg13g2_nor2_1 _1121_ (.A(_0326_),
    .B(_0327_),
    .Y(_0328_));
 sg13g2_nor2_1 _1122_ (.A(_0092_),
    .B(_0322_),
    .Y(_0329_));
 sg13g2_and2_1 _1123_ (.A(_0328_),
    .B(_0329_),
    .X(_0330_));
 sg13g2_a221oi_1 _1124_ (.B2(_0325_),
    .C1(_0330_),
    .B1(_0321_),
    .A1(_0101_),
    .Y(_0331_),
    .A2(\rca.generate_adder_modules[7].fa.a ));
 sg13g2_xor2_1 _1125_ (.B(net55),
    .A(net54),
    .X(_0332_));
 sg13g2_nand2_1 _1126_ (.Y(_0333_),
    .A(net56),
    .B(_0332_));
 sg13g2_xnor2_1 _1127_ (.Y(_0334_),
    .A(_0331_),
    .B(_0333_));
 sg13g2_nor2_1 _1128_ (.A(net43),
    .B(\cla_z[8] ),
    .Y(_0335_));
 sg13g2_a21oi_1 _1129_ (.A1(net43),
    .A2(_0334_),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_nand2_1 _1130_ (.Y(_0337_),
    .A(_0306_),
    .B(_0336_));
 sg13g2_nor2b_1 _1131_ (.A(_0282_),
    .B_N(net40),
    .Y(_0338_));
 sg13g2_buf_2 _1132_ (.A(_0338_),
    .X(_0339_));
 sg13g2_nand2_1 _1133_ (.Y(_0340_),
    .A(net56),
    .B(_0307_));
 sg13g2_buf_1 _1134_ (.A(_0340_),
    .X(_0341_));
 sg13g2_nand2_1 _1135_ (.Y(_0342_),
    .A(_0136_),
    .B(_0111_));
 sg13g2_xnor2_1 _1136_ (.Y(_0343_),
    .A(\io_sd._053_[1] ),
    .B(\io_sd._052_[1] ));
 sg13g2_xnor2_1 _1137_ (.Y(_0344_),
    .A(_0342_),
    .B(_0343_));
 sg13g2_inv_2 _1138_ (.Y(_0345_),
    .A(_0307_));
 sg13g2_nand2_1 _1139_ (.Y(_0346_),
    .A(_0345_),
    .B(\cla_z[1] ));
 sg13g2_o21ai_1 _1140_ (.B1(_0346_),
    .Y(_0347_),
    .A1(net26),
    .A2(_0344_));
 sg13g2_nand2_1 _1141_ (.Y(_0348_),
    .A(_0339_),
    .B(_0347_));
 sg13g2_nand3_1 _1142_ (.B(_0337_),
    .C(_0348_),
    .A(net27),
    .Y(_0349_));
 sg13g2_nor2_1 _1143_ (.A(_0083_),
    .B(_0282_),
    .Y(_0350_));
 sg13g2_nor2_1 _1144_ (.A(_0092_),
    .B(_0345_),
    .Y(_0351_));
 sg13g2_buf_2 _1145_ (.A(_0351_),
    .X(_0352_));
 sg13g2_nand2_2 _1146_ (.Y(_0353_),
    .A(_0352_),
    .B(_0306_));
 sg13g2_xnor2_1 _1147_ (.Y(_0354_),
    .A(\io_sd._053_[9] ),
    .B(\io_sd._052_[9] ));
 sg13g2_nor3_1 _1148_ (.A(net55),
    .B(_0353_),
    .C(_0354_),
    .Y(_0355_));
 sg13g2_nor3_1 _1149_ (.A(_0100_),
    .B(_0353_),
    .C(_0354_),
    .Y(_0356_));
 sg13g2_o21ai_1 _1150_ (.B1(_0331_),
    .Y(_0357_),
    .A1(_0355_),
    .A2(_0356_));
 sg13g2_nand2_1 _1151_ (.Y(_0358_),
    .A(_0300_),
    .B(_0304_));
 sg13g2_nor2_1 _1152_ (.A(net26),
    .B(_0358_),
    .Y(_0359_));
 sg13g2_nand3_1 _1153_ (.B(_0359_),
    .C(_0354_),
    .A(net55),
    .Y(_0360_));
 sg13g2_nand3_1 _1154_ (.B(_0359_),
    .C(_0354_),
    .A(net54),
    .Y(_0361_));
 sg13g2_a21o_1 _1155_ (.A2(_0361_),
    .A1(_0360_),
    .B1(_0331_),
    .X(_0362_));
 sg13g2_nor2_2 _1156_ (.A(_0307_),
    .B(_0358_),
    .Y(_0363_));
 sg13g2_nor3_1 _1157_ (.A(net54),
    .B(_0099_),
    .C(_0354_),
    .Y(_0364_));
 sg13g2_and4_1 _1158_ (.A(net54),
    .B(net55),
    .C(_0359_),
    .D(_0354_),
    .X(_0365_));
 sg13g2_a221oi_1 _1159_ (.B2(_0359_),
    .C1(_0365_),
    .B1(_0364_),
    .A1(\cla_z[9] ),
    .Y(_0366_),
    .A2(_0363_));
 sg13g2_and3_1 _1160_ (.X(_0367_),
    .A(_0357_),
    .B(_0362_),
    .C(_0366_));
 sg13g2_buf_1 _1161_ (.A(_0345_),
    .X(_0368_));
 sg13g2_buf_1 _1162_ (.A(_0352_),
    .X(_0369_));
 sg13g2_xor2_1 _1163_ (.B(_0111_),
    .A(_0136_),
    .X(_0370_));
 sg13g2_a22oi_1 _1164_ (.Y(_0371_),
    .B1(net25),
    .B2(_0370_),
    .A2(\cla_z[0] ),
    .A1(net33));
 sg13g2_nor2_2 _1165_ (.A(_0084_),
    .B(_0283_),
    .Y(_0372_));
 sg13g2_a22oi_1 _1166_ (.Y(_0373_),
    .B1(_0371_),
    .B2(_0372_),
    .A2(_0367_),
    .A1(_0350_));
 sg13g2_buf_1 _1167_ (.A(_0282_),
    .X(_0374_));
 sg13g2_nor2_1 _1168_ (.A(net41),
    .B(net32),
    .Y(_0375_));
 sg13g2_a22oi_1 _1169_ (.Y(_0376_),
    .B1(_0348_),
    .B2(_0375_),
    .A2(_0296_),
    .A1(net41));
 sg13g2_nand4_1 _1170_ (.B(_0349_),
    .C(_0373_),
    .A(_0299_),
    .Y(_0377_),
    .D(_0376_));
 sg13g2_nor2b_1 _1171_ (.A(net60),
    .B_N(_0070_),
    .Y(_0378_));
 sg13g2_buf_2 _1172_ (.A(_0378_),
    .X(_0379_));
 sg13g2_nand2_1 _1173_ (.Y(_0380_),
    .A(net11),
    .B(_0379_));
 sg13g2_nand2_1 _1174_ (.Y(_0381_),
    .A(_0081_),
    .B(_0299_));
 sg13g2_nand2_1 _1175_ (.Y(_0382_),
    .A(net40),
    .B(net28));
 sg13g2_nor2_1 _1176_ (.A(net20),
    .B(_0382_),
    .Y(_0383_));
 sg13g2_and3_1 _1177_ (.X(_0384_),
    .A(\cla_z[17] ),
    .B(_0363_),
    .C(_0383_));
 sg13g2_xor2_1 _1178_ (.B(\io_sd._052_[17] ),
    .A(\io_sd._053_[17] ),
    .X(_0385_));
 sg13g2_inv_1 _1179_ (.Y(_0386_),
    .A(_0385_));
 sg13g2_nor3_1 _1180_ (.A(net54),
    .B(\io_sd._053_[9] ),
    .C(net55),
    .Y(_0387_));
 sg13g2_o21ai_1 _1181_ (.B1(\io_sd._053_[9] ),
    .Y(_0388_),
    .A1(net54),
    .A2(net55));
 sg13g2_o21ai_1 _1182_ (.B1(_0388_),
    .Y(_0389_),
    .A1(_0094_),
    .A2(_0387_));
 sg13g2_and2_1 _1183_ (.A(net56),
    .B(_0389_),
    .X(_0390_));
 sg13g2_or2_1 _1184_ (.X(_0391_),
    .B(\io_sd._052_[7] ),
    .A(_0101_));
 sg13g2_nand2_1 _1185_ (.Y(_0392_),
    .A(_0101_),
    .B(\io_sd._052_[7] ));
 sg13g2_o21ai_1 _1186_ (.B1(_0392_),
    .Y(_0393_),
    .A1(_0326_),
    .A2(_0327_));
 sg13g2_nand2_1 _1187_ (.Y(_0394_),
    .A(net54),
    .B(net55));
 sg13g2_o21ai_1 _1188_ (.B1(_0394_),
    .Y(_0395_),
    .A1(_0095_),
    .A2(_0094_));
 sg13g2_a21o_1 _1189_ (.A2(_0393_),
    .A1(_0391_),
    .B1(_0395_),
    .X(_0396_));
 sg13g2_and3_1 _1190_ (.X(_0397_),
    .A(net56),
    .B(_0389_),
    .C(_0325_));
 sg13g2_a22oi_1 _1191_ (.Y(_0398_),
    .B1(_0321_),
    .B2(_0397_),
    .A2(_0396_),
    .A1(_0390_));
 sg13g2_buf_2 _1192_ (.A(_0398_),
    .X(_0399_));
 sg13g2_xor2_1 _1193_ (.B(net52),
    .A(net51),
    .X(_0400_));
 sg13g2_nand2_1 _1194_ (.Y(_0401_),
    .A(_0091_),
    .B(_0400_));
 sg13g2_xnor2_1 _1195_ (.Y(_0402_),
    .A(_0124_),
    .B(_0123_));
 sg13g2_xnor2_1 _1196_ (.Y(_0403_),
    .A(\io_sd._053_[12] ),
    .B(\io_sd._052_[12] ));
 sg13g2_nor3_2 _1197_ (.A(_0401_),
    .B(_0402_),
    .C(_0403_),
    .Y(_0404_));
 sg13g2_nand2_1 _1198_ (.Y(_0405_),
    .A(_0117_),
    .B(_0116_));
 sg13g2_nor2_1 _1199_ (.A(_0120_),
    .B(_0118_),
    .Y(_0406_));
 sg13g2_nor2_1 _1200_ (.A(_0117_),
    .B(_0116_),
    .Y(_0407_));
 sg13g2_a21oi_1 _1201_ (.A1(_0405_),
    .A2(_0406_),
    .Y(_0408_),
    .B1(_0407_));
 sg13g2_or2_1 _1202_ (.X(_0409_),
    .B(_0114_),
    .A(_0115_));
 sg13g2_and2_1 _1203_ (.A(_0408_),
    .B(_0409_),
    .X(_0410_));
 sg13g2_nand2_1 _1204_ (.Y(_0411_),
    .A(_0404_),
    .B(_0410_));
 sg13g2_nor2_1 _1205_ (.A(\io_sd._053_[12] ),
    .B(\io_sd._052_[12] ),
    .Y(_0412_));
 sg13g2_and3_1 _1206_ (.X(_0413_),
    .A(_0091_),
    .B(net51),
    .C(net52));
 sg13g2_or2_1 _1207_ (.X(_0414_),
    .B(_0123_),
    .A(_0124_));
 sg13g2_and2_1 _1208_ (.A(_0124_),
    .B(_0123_),
    .X(_0415_));
 sg13g2_a221oi_1 _1209_ (.B2(_0414_),
    .C1(_0415_),
    .B1(_0413_),
    .A1(\io_sd._053_[12] ),
    .Y(_0416_),
    .A2(\io_sd._052_[12] ));
 sg13g2_a22oi_1 _1210_ (.Y(_0417_),
    .B1(_0116_),
    .B2(_0117_),
    .A2(_0118_),
    .A1(_0120_));
 sg13g2_o21ai_1 _1211_ (.B1(_0417_),
    .Y(_0418_),
    .A1(_0412_),
    .A2(_0416_));
 sg13g2_buf_2 _1212_ (.A(_0418_),
    .X(_0419_));
 sg13g2_a22oi_1 _1213_ (.Y(_0420_),
    .B1(_0419_),
    .B2(_0410_),
    .A2(_0114_),
    .A1(_0115_));
 sg13g2_o21ai_1 _1214_ (.B1(_0420_),
    .Y(_0421_),
    .A1(_0399_),
    .A2(_0411_));
 sg13g2_a21oi_1 _1215_ (.A1(net53),
    .A2(_0421_),
    .Y(_0422_),
    .B1(_0113_));
 sg13g2_nor2_1 _1216_ (.A(net53),
    .B(_0421_),
    .Y(_0423_));
 sg13g2_nor3_1 _1217_ (.A(_0386_),
    .B(_0422_),
    .C(_0423_),
    .Y(_0424_));
 sg13g2_nor2_1 _1218_ (.A(_0113_),
    .B(net53),
    .Y(_0425_));
 sg13g2_nor2_1 _1219_ (.A(net39),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_a221oi_1 _1220_ (.B2(_0426_),
    .C1(_0385_),
    .B1(_0421_),
    .A1(_0113_),
    .Y(_0427_),
    .A2(net53));
 sg13g2_inv_1 _1221_ (.Y(_0428_),
    .A(net41));
 sg13g2_nor3_1 _1222_ (.A(_0428_),
    .B(_0294_),
    .C(_0298_),
    .Y(_0429_));
 sg13g2_nand2_1 _1223_ (.Y(_0430_),
    .A(_0429_),
    .B(_0339_));
 sg13g2_nor4_1 _1224_ (.A(_0353_),
    .B(_0424_),
    .C(_0427_),
    .D(_0430_),
    .Y(_0431_));
 sg13g2_nand2b_1 _1225_ (.Y(_0432_),
    .B(_0282_),
    .A_N(net40));
 sg13g2_xnor2_1 _1226_ (.Y(_0433_),
    .A(_0113_),
    .B(net53));
 sg13g2_xnor2_1 _1227_ (.Y(_0434_),
    .A(_0421_),
    .B(_0433_));
 sg13g2_a22oi_1 _1228_ (.Y(_0435_),
    .B1(net25),
    .B2(_0434_),
    .A2(\cla_z[16] ),
    .A1(net33));
 sg13g2_nor3_1 _1229_ (.A(net20),
    .B(_0432_),
    .C(_0435_),
    .Y(_0436_));
 sg13g2_nor3_1 _1230_ (.A(_0384_),
    .B(_0431_),
    .C(_0436_),
    .Y(_0437_));
 sg13g2_nand3_1 _1231_ (.B(_0380_),
    .C(_0437_),
    .A(_0377_),
    .Y(_0062_));
 sg13g2_buf_8 _1232_ (.A(_0399_),
    .X(_0438_));
 sg13g2_xnor2_1 _1233_ (.Y(_0439_),
    .A(net19),
    .B(_0401_));
 sg13g2_o21ai_1 _1234_ (.B1(_0306_),
    .Y(_0440_),
    .A1(net43),
    .A2(\cla_z[10] ));
 sg13g2_a21oi_1 _1235_ (.A1(_0308_),
    .A2(_0439_),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_nor2_1 _1236_ (.A(_0296_),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_a21oi_1 _1237_ (.A1(_0303_),
    .A2(_0367_),
    .Y(_0443_),
    .B1(_0442_));
 sg13g2_or3_1 _1238_ (.A(_0353_),
    .B(_0424_),
    .C(_0427_),
    .X(_0444_));
 sg13g2_nand2_1 _1239_ (.Y(_0445_),
    .A(net41),
    .B(net32));
 sg13g2_a21oi_1 _1240_ (.A1(\cla_z[17] ),
    .A2(_0363_),
    .Y(_0446_),
    .B1(_0445_));
 sg13g2_xor2_1 _1241_ (.B(\io_sd._052_[18] ),
    .A(_0128_),
    .X(_0447_));
 sg13g2_nand2_1 _1242_ (.Y(_0448_),
    .A(net56),
    .B(_0447_));
 sg13g2_nor2_1 _1243_ (.A(\io_sd._053_[17] ),
    .B(\io_sd._052_[17] ),
    .Y(_0449_));
 sg13g2_nor2_1 _1244_ (.A(_0092_),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_xor2_1 _1245_ (.B(_0114_),
    .A(_0115_),
    .X(_0451_));
 sg13g2_nand2_1 _1246_ (.Y(_0452_),
    .A(\io_sd._053_[17] ),
    .B(\io_sd._052_[17] ));
 sg13g2_nand2_1 _1247_ (.Y(_0453_),
    .A(_0425_),
    .B(_0452_));
 sg13g2_and4_1 _1248_ (.A(_0408_),
    .B(_0450_),
    .C(_0451_),
    .D(_0453_),
    .X(_0454_));
 sg13g2_buf_2 _1249_ (.A(_0454_),
    .X(_0455_));
 sg13g2_nand2_1 _1250_ (.Y(_0456_),
    .A(_0404_),
    .B(_0455_));
 sg13g2_nand4_1 _1251_ (.B(_0115_),
    .C(_0114_),
    .A(_0091_),
    .Y(_0457_),
    .D(net53));
 sg13g2_nor2b_1 _1252_ (.A(_0113_),
    .B_N(_0457_),
    .Y(_0458_));
 sg13g2_a21oi_1 _1253_ (.A1(_0115_),
    .A2(\rca.generate_adder_modules[15].fa.a ),
    .Y(_0459_),
    .B1(net53));
 sg13g2_o21ai_1 _1254_ (.B1(_0452_),
    .Y(_0460_),
    .A1(_0458_),
    .A2(_0459_));
 sg13g2_a22oi_1 _1255_ (.Y(_0461_),
    .B1(_0455_),
    .B2(_0419_),
    .A2(_0460_),
    .A1(_0450_));
 sg13g2_o21ai_1 _1256_ (.B1(_0461_),
    .Y(_0462_),
    .A1(net19),
    .A2(_0456_));
 sg13g2_xnor2_1 _1257_ (.Y(_0463_),
    .A(_0448_),
    .B(_0462_));
 sg13g2_nand2_1 _1258_ (.Y(_0464_),
    .A(net43),
    .B(_0463_));
 sg13g2_nand2_1 _1259_ (.Y(_0465_),
    .A(\cla_z[18] ),
    .B(_0363_));
 sg13g2_a21o_1 _1260_ (.A2(_0465_),
    .A1(_0464_),
    .B1(net32),
    .X(_0466_));
 sg13g2_and2_1 _1261_ (.A(net41),
    .B(net27),
    .X(_0467_));
 sg13g2_inv_1 _1262_ (.Y(_0468_),
    .A(\io_sd._053_[1] ));
 sg13g2_a21oi_1 _1263_ (.A1(_0468_),
    .A2(_0311_),
    .Y(_0469_),
    .B1(_0310_));
 sg13g2_xnor2_1 _1264_ (.Y(_0470_),
    .A(_0108_),
    .B(_0106_));
 sg13g2_xnor2_1 _1265_ (.Y(_0471_),
    .A(_0469_),
    .B(_0470_));
 sg13g2_a22oi_1 _1266_ (.Y(_0472_),
    .B1(net25),
    .B2(_0471_),
    .A2(\cla_z[2] ),
    .A1(_0345_));
 sg13g2_a21oi_1 _1267_ (.A1(_0282_),
    .A2(_0347_),
    .Y(_0473_),
    .B1(net40));
 sg13g2_a21oi_1 _1268_ (.A1(net28),
    .A2(_0472_),
    .Y(_0474_),
    .B1(_0473_));
 sg13g2_o21ai_1 _1269_ (.B1(_0299_),
    .Y(_0475_),
    .A1(net41),
    .A2(_0474_));
 sg13g2_a221oi_1 _1270_ (.B2(_0467_),
    .C1(_0475_),
    .B1(_0466_),
    .A1(_0444_),
    .Y(_0476_),
    .A2(_0446_));
 sg13g2_and2_1 _1271_ (.A(net12),
    .B(_0379_),
    .X(_0477_));
 sg13g2_a21o_1 _1272_ (.A2(_0476_),
    .A1(_0443_),
    .B1(_0477_),
    .X(_0063_));
 sg13g2_nand2_1 _1273_ (.Y(_0478_),
    .A(net33),
    .B(\cla_z[18] ));
 sg13g2_a21oi_1 _1274_ (.A1(_0464_),
    .A2(_0478_),
    .Y(_0479_),
    .B1(_0358_));
 sg13g2_o21ai_1 _1275_ (.B1(_0429_),
    .Y(_0480_),
    .A1(net27),
    .A2(_0479_));
 sg13g2_a21oi_1 _1276_ (.A1(_0129_),
    .A2(_0127_),
    .Y(_0481_),
    .B1(_0461_));
 sg13g2_nand3_1 _1277_ (.B(_0404_),
    .C(_0455_),
    .A(\io_sd._052_[18] ),
    .Y(_0482_));
 sg13g2_nor2_1 _1278_ (.A(net19),
    .B(_0482_),
    .Y(_0483_));
 sg13g2_nand3_1 _1279_ (.B(_0404_),
    .C(_0455_),
    .A(_0128_),
    .Y(_0484_));
 sg13g2_nand2_1 _1280_ (.Y(_0485_),
    .A(_0128_),
    .B(\rca.generate_adder_modules[18].fa.a ));
 sg13g2_o21ai_1 _1281_ (.B1(_0485_),
    .Y(_0486_),
    .A1(net19),
    .A2(_0484_));
 sg13g2_nor3_1 _1282_ (.A(_0481_),
    .B(_0483_),
    .C(_0486_),
    .Y(_0487_));
 sg13g2_nand2_1 _1283_ (.Y(_0488_),
    .A(\io_sd._053_[19] ),
    .B(\io_sd._052_[19] ));
 sg13g2_or2_1 _1284_ (.X(_0489_),
    .B(\io_sd._052_[19] ),
    .A(\io_sd._053_[19] ));
 sg13g2_buf_1 _1285_ (.A(_0489_),
    .X(_0490_));
 sg13g2_nand2_1 _1286_ (.Y(_0491_),
    .A(_0488_),
    .B(_0490_));
 sg13g2_xnor2_1 _1287_ (.Y(_0492_),
    .A(_0487_),
    .B(_0491_));
 sg13g2_nand2_1 _1288_ (.Y(_0493_),
    .A(\cla_z[19] ),
    .B(_0363_));
 sg13g2_o21ai_1 _1289_ (.B1(_0493_),
    .Y(_0494_),
    .A1(_0353_),
    .A2(_0492_));
 sg13g2_a21oi_1 _1290_ (.A1(_0339_),
    .A2(_0494_),
    .Y(_0495_),
    .B1(_0372_));
 sg13g2_xnor2_1 _1291_ (.Y(_0496_),
    .A(_0081_),
    .B(_0350_));
 sg13g2_and2_1 _1292_ (.A(_0299_),
    .B(_0496_),
    .X(_0497_));
 sg13g2_and2_1 _1293_ (.A(net40),
    .B(_0497_),
    .X(_0498_));
 sg13g2_buf_1 _1294_ (.A(net26),
    .X(_0499_));
 sg13g2_o21ai_1 _1295_ (.B1(_0313_),
    .Y(_0500_),
    .A1(_0108_),
    .A2(_0106_));
 sg13g2_xnor2_1 _1296_ (.Y(_0501_),
    .A(\io_sd._053_[3] ),
    .B(\io_sd._052_[3] ));
 sg13g2_xnor2_1 _1297_ (.Y(_0502_),
    .A(_0500_),
    .B(_0501_));
 sg13g2_nand2_1 _1298_ (.Y(_0503_),
    .A(net33),
    .B(\cla_z[3] ));
 sg13g2_o21ai_1 _1299_ (.B1(_0503_),
    .Y(_0504_),
    .A1(_0499_),
    .A2(_0502_));
 sg13g2_mux2_1 _1300_ (.A0(_0441_),
    .A1(_0504_),
    .S(net28),
    .X(_0505_));
 sg13g2_nand2_1 _1301_ (.Y(_0506_),
    .A(_0299_),
    .B(_0496_));
 sg13g2_nand2_1 _1302_ (.Y(_0507_),
    .A(_0345_),
    .B(\cla_z[11] ));
 sg13g2_nor3_1 _1303_ (.A(net52),
    .B(net26),
    .C(_0402_),
    .Y(_0508_));
 sg13g2_nor3_1 _1304_ (.A(net51),
    .B(net26),
    .C(_0402_),
    .Y(_0509_));
 sg13g2_o21ai_1 _1305_ (.B1(net19),
    .Y(_0510_),
    .A1(_0508_),
    .A2(_0509_));
 sg13g2_nand3_1 _1306_ (.B(_0352_),
    .C(_0402_),
    .A(net52),
    .Y(_0511_));
 sg13g2_nand3_1 _1307_ (.B(_0352_),
    .C(_0402_),
    .A(net51),
    .Y(_0512_));
 sg13g2_a21o_1 _1308_ (.A2(_0512_),
    .A1(_0511_),
    .B1(net19),
    .X(_0513_));
 sg13g2_or2_1 _1309_ (.X(_0514_),
    .B(net52),
    .A(net51));
 sg13g2_nor3_1 _1310_ (.A(net26),
    .B(_0402_),
    .C(_0514_),
    .Y(_0515_));
 sg13g2_nand4_1 _1311_ (.B(_0125_),
    .C(_0352_),
    .A(net51),
    .Y(_0516_),
    .D(_0402_));
 sg13g2_nor2b_1 _1312_ (.A(_0515_),
    .B_N(_0516_),
    .Y(_0517_));
 sg13g2_nand4_1 _1313_ (.B(_0510_),
    .C(_0513_),
    .A(_0507_),
    .Y(_0518_),
    .D(_0517_));
 sg13g2_nor2_1 _1314_ (.A(net28),
    .B(_0472_),
    .Y(_0519_));
 sg13g2_a21oi_1 _1315_ (.A1(net28),
    .A2(_0518_),
    .Y(_0520_),
    .B1(_0519_));
 sg13g2_nor3_1 _1316_ (.A(net27),
    .B(_0506_),
    .C(_0520_),
    .Y(_0521_));
 sg13g2_a221oi_1 _1317_ (.B2(_0505_),
    .C1(_0521_),
    .B1(_0498_),
    .A1(net13),
    .Y(_0522_),
    .A2(_0379_));
 sg13g2_o21ai_1 _1318_ (.B1(_0522_),
    .Y(_0064_),
    .A1(_0480_),
    .A2(_0495_));
 sg13g2_or2_1 _1319_ (.X(_0523_),
    .B(\io_sd._052_[18] ),
    .A(_0128_));
 sg13g2_and2_1 _1320_ (.A(\io_sd._053_[19] ),
    .B(\io_sd._052_[19] ),
    .X(_0524_));
 sg13g2_a21oi_1 _1321_ (.A1(_0490_),
    .A2(_0523_),
    .Y(_0525_),
    .B1(_0524_));
 sg13g2_nand2_1 _1322_ (.Y(_0526_),
    .A(_0129_),
    .B(_0488_));
 sg13g2_a221oi_1 _1323_ (.B2(_0419_),
    .C1(_0526_),
    .B1(_0455_),
    .A1(_0450_),
    .Y(_0527_),
    .A2(_0460_));
 sg13g2_o21ai_1 _1324_ (.B1(_0527_),
    .Y(_0528_),
    .A1(_0399_),
    .A2(_0456_));
 sg13g2_nand2_1 _1325_ (.Y(_0529_),
    .A(_0127_),
    .B(_0488_));
 sg13g2_a221oi_1 _1326_ (.B2(_0419_),
    .C1(_0529_),
    .B1(_0455_),
    .A1(_0450_),
    .Y(_0530_),
    .A2(_0460_));
 sg13g2_o21ai_1 _1327_ (.B1(_0530_),
    .Y(_0531_),
    .A1(_0399_),
    .A2(_0456_));
 sg13g2_nand3b_1 _1328_ (.B(_0528_),
    .C(_0531_),
    .Y(_0532_),
    .A_N(_0525_));
 sg13g2_buf_2 _1329_ (.A(_0532_),
    .X(_0533_));
 sg13g2_xnor2_1 _1330_ (.Y(_0534_),
    .A(net49),
    .B(net50));
 sg13g2_xnor2_1 _1331_ (.Y(_0535_),
    .A(_0533_),
    .B(_0534_));
 sg13g2_nand2_1 _1332_ (.Y(_0536_),
    .A(\cla_z[20] ),
    .B(_0363_));
 sg13g2_o21ai_1 _1333_ (.B1(_0536_),
    .Y(_0537_),
    .A1(_0353_),
    .A2(_0535_));
 sg13g2_a22oi_1 _1334_ (.Y(_0538_),
    .B1(_0537_),
    .B2(_0339_),
    .A2(_0494_),
    .A1(_0372_));
 sg13g2_nand2_1 _1335_ (.Y(_0539_),
    .A(_0124_),
    .B(_0123_));
 sg13g2_nand2b_1 _1336_ (.Y(_0540_),
    .B(_0539_),
    .A_N(net52));
 sg13g2_a221oi_1 _1337_ (.B2(_0397_),
    .C1(_0540_),
    .B1(_0321_),
    .A1(_0390_),
    .Y(_0541_),
    .A2(_0396_));
 sg13g2_nand2b_1 _1338_ (.Y(_0542_),
    .B(_0539_),
    .A_N(net51));
 sg13g2_a221oi_1 _1339_ (.B2(_0397_),
    .C1(_0542_),
    .B1(_0321_),
    .A1(_0390_),
    .Y(_0543_),
    .A2(_0396_));
 sg13g2_o21ai_1 _1340_ (.B1(_0414_),
    .Y(_0544_),
    .A1(_0415_),
    .A2(_0514_));
 sg13g2_nor3_1 _1341_ (.A(_0541_),
    .B(_0543_),
    .C(_0544_),
    .Y(_0545_));
 sg13g2_xnor2_1 _1342_ (.Y(_0546_),
    .A(_0403_),
    .B(_0545_));
 sg13g2_nor2b_1 _1343_ (.A(_0308_),
    .B_N(\cla_z[12] ),
    .Y(_0547_));
 sg13g2_a21o_1 _1344_ (.A2(_0546_),
    .A1(net25),
    .B1(_0547_),
    .X(_0548_));
 sg13g2_a21oi_1 _1345_ (.A1(_0500_),
    .A2(_0318_),
    .Y(_0549_),
    .B1(_0315_));
 sg13g2_xor2_1 _1346_ (.B(\io_sd._052_[4] ),
    .A(\io_sd._053_[4] ),
    .X(_0550_));
 sg13g2_xnor2_1 _1347_ (.Y(_0551_),
    .A(_0549_),
    .B(_0550_));
 sg13g2_nand2_1 _1348_ (.Y(_0552_),
    .A(net33),
    .B(\cla_z[4] ));
 sg13g2_o21ai_1 _1349_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0499_),
    .A2(_0551_));
 sg13g2_mux4_1 _1350_ (.S0(net28),
    .A0(_0504_),
    .A1(_0548_),
    .A2(_0518_),
    .A3(_0553_),
    .S1(net27),
    .X(_0554_));
 sg13g2_a22oi_1 _1351_ (.Y(_0555_),
    .B1(_0497_),
    .B2(_0554_),
    .A2(_0379_),
    .A1(net14));
 sg13g2_o21ai_1 _1352_ (.B1(_0555_),
    .Y(_0065_),
    .A1(_0381_),
    .A2(_0538_));
 sg13g2_nor2_1 _1353_ (.A(net24),
    .B(_0382_),
    .Y(_0556_));
 sg13g2_nand2_1 _1354_ (.Y(_0557_),
    .A(_0131_),
    .B(net50));
 sg13g2_nor2_1 _1355_ (.A(net49),
    .B(_0130_),
    .Y(_0558_));
 sg13g2_a21oi_1 _1356_ (.A1(_0533_),
    .A2(_0557_),
    .Y(_0559_),
    .B1(_0558_));
 sg13g2_xnor2_1 _1357_ (.Y(_0560_),
    .A(_0133_),
    .B(_0132_));
 sg13g2_xnor2_1 _1358_ (.Y(_0561_),
    .A(_0559_),
    .B(_0560_));
 sg13g2_a22oi_1 _1359_ (.Y(_0562_),
    .B1(_0556_),
    .B2(_0561_),
    .A2(_0537_),
    .A1(_0372_));
 sg13g2_nor2b_1 _1360_ (.A(net43),
    .B_N(\cla_z[13] ),
    .Y(_0563_));
 sg13g2_xor2_1 _1361_ (.B(_0118_),
    .A(_0120_),
    .X(_0564_));
 sg13g2_nand2_1 _1362_ (.Y(_0565_),
    .A(net56),
    .B(_0564_));
 sg13g2_or3_1 _1363_ (.A(_0401_),
    .B(_0402_),
    .C(_0403_),
    .X(_0566_));
 sg13g2_or3_1 _1364_ (.A(_0092_),
    .B(_0412_),
    .C(_0416_),
    .X(_0567_));
 sg13g2_o21ai_1 _1365_ (.B1(_0567_),
    .Y(_0568_),
    .A1(net19),
    .A2(_0566_));
 sg13g2_nand2b_1 _1366_ (.Y(_0569_),
    .B(_0568_),
    .A_N(_0565_));
 sg13g2_and2_1 _1367_ (.A(_0567_),
    .B(_0565_),
    .X(_0570_));
 sg13g2_o21ai_1 _1368_ (.B1(_0570_),
    .Y(_0571_),
    .A1(_0438_),
    .A2(_0566_));
 sg13g2_and3_1 _1369_ (.X(_0572_),
    .A(net43),
    .B(_0306_),
    .C(_0571_));
 sg13g2_a22oi_1 _1370_ (.Y(_0573_),
    .B1(_0569_),
    .B2(_0572_),
    .A2(_0563_),
    .A1(_0306_));
 sg13g2_nor3_1 _1371_ (.A(_0296_),
    .B(net20),
    .C(_0573_),
    .Y(_0574_));
 sg13g2_and4_1 _1372_ (.A(_0374_),
    .B(net25),
    .C(_0498_),
    .D(_0546_),
    .X(_0575_));
 sg13g2_nand2_1 _1373_ (.Y(_0576_),
    .A(_0096_),
    .B(_0321_));
 sg13g2_xor2_1 _1374_ (.B(_0576_),
    .A(_0324_),
    .X(_0577_));
 sg13g2_a22oi_1 _1375_ (.Y(_0578_),
    .B1(net25),
    .B2(_0577_),
    .A2(\cla_z[5] ),
    .A1(net33));
 sg13g2_nand2_1 _1376_ (.Y(_0579_),
    .A(net28),
    .B(_0498_));
 sg13g2_nand3_1 _1377_ (.B(_0498_),
    .C(_0547_),
    .A(net32),
    .Y(_0580_));
 sg13g2_o21ai_1 _1378_ (.B1(_0580_),
    .Y(_0581_),
    .A1(_0578_),
    .A2(_0579_));
 sg13g2_nand4_1 _1379_ (.B(_0290_),
    .C(_0299_),
    .A(_0374_),
    .Y(_0582_),
    .D(_0553_));
 sg13g2_nor2b_1 _1380_ (.A(net43),
    .B_N(\cla_z[21] ),
    .Y(_0583_));
 sg13g2_a22oi_1 _1381_ (.Y(_0584_),
    .B1(_0383_),
    .B2(_0583_),
    .A2(_0379_),
    .A1(net15));
 sg13g2_nand2_1 _1382_ (.Y(_0585_),
    .A(_0582_),
    .B(_0584_));
 sg13g2_nor4_1 _1383_ (.A(_0574_),
    .B(_0575_),
    .C(_0581_),
    .D(_0585_),
    .Y(_0586_));
 sg13g2_o21ai_1 _1384_ (.B1(_0586_),
    .Y(_0066_),
    .A1(net20),
    .A2(_0562_));
 sg13g2_and2_1 _1385_ (.A(net16),
    .B(_0379_),
    .X(_0587_));
 sg13g2_a221oi_1 _1386_ (.B2(_0317_),
    .C1(_0319_),
    .B1(_0313_),
    .A1(_0105_),
    .Y(_0588_),
    .A2(_0104_));
 sg13g2_or2_1 _1387_ (.X(_0589_),
    .B(_0104_),
    .A(_0105_));
 sg13g2_nor2b_1 _1388_ (.A(_0588_),
    .B_N(_0589_),
    .Y(_0590_));
 sg13g2_xnor2_1 _1389_ (.Y(_0591_),
    .A(_0323_),
    .B(_0590_));
 sg13g2_a221oi_1 _1390_ (.B2(_0591_),
    .C1(net32),
    .B1(_0369_),
    .A1(_0368_),
    .Y(_0592_),
    .A2(\cla_z[6] ));
 sg13g2_a21o_1 _1391_ (.A2(_0573_),
    .A1(net32),
    .B1(_0592_),
    .X(_0593_));
 sg13g2_nand2_1 _1392_ (.Y(_0594_),
    .A(_0118_),
    .B(_0404_));
 sg13g2_nand2_1 _1393_ (.Y(_0595_),
    .A(_0120_),
    .B(_0404_));
 sg13g2_a21oi_1 _1394_ (.A1(_0594_),
    .A2(_0595_),
    .Y(_0596_),
    .B1(net19));
 sg13g2_a21oi_1 _1395_ (.A1(_0121_),
    .A2(_0119_),
    .Y(_0597_),
    .B1(_0567_));
 sg13g2_a21o_1 _1396_ (.A2(_0118_),
    .A1(_0120_),
    .B1(_0597_),
    .X(_0598_));
 sg13g2_xor2_1 _1397_ (.B(_0116_),
    .A(_0117_),
    .X(_0599_));
 sg13g2_nand2_1 _1398_ (.Y(_0600_),
    .A(_0352_),
    .B(_0599_));
 sg13g2_nor3_1 _1399_ (.A(_0596_),
    .B(_0598_),
    .C(_0600_),
    .Y(_0601_));
 sg13g2_nor2_1 _1400_ (.A(net26),
    .B(_0599_),
    .Y(_0602_));
 sg13g2_o21ai_1 _1401_ (.B1(_0602_),
    .Y(_0603_),
    .A1(_0596_),
    .A2(_0598_));
 sg13g2_nor2b_1 _1402_ (.A(_0601_),
    .B_N(_0603_),
    .Y(_0604_));
 sg13g2_nand2_1 _1403_ (.Y(_0605_),
    .A(net33),
    .B(\cla_z[14] ));
 sg13g2_nand2_1 _1404_ (.Y(_0606_),
    .A(net28),
    .B(_0300_));
 sg13g2_a21o_1 _1405_ (.A2(_0605_),
    .A1(_0604_),
    .B1(_0606_),
    .X(_0607_));
 sg13g2_nor2_1 _1406_ (.A(_0284_),
    .B(_0578_),
    .Y(_0608_));
 sg13g2_nor2_1 _1407_ (.A(net27),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_a221oi_1 _1408_ (.B2(_0609_),
    .C1(_0506_),
    .B1(_0607_),
    .A1(net27),
    .Y(_0610_),
    .A2(_0593_));
 sg13g2_o21ai_1 _1409_ (.B1(_0488_),
    .Y(_0611_),
    .A1(_0129_),
    .A2(_0127_));
 sg13g2_nand2_1 _1410_ (.Y(_0612_),
    .A(_0133_),
    .B(_0132_));
 sg13g2_nand2_1 _1411_ (.Y(_0613_),
    .A(_0557_),
    .B(_0612_));
 sg13g2_a21oi_1 _1412_ (.A1(_0490_),
    .A2(_0611_),
    .Y(_0614_),
    .B1(_0613_));
 sg13g2_nor2_1 _1413_ (.A(_0133_),
    .B(_0132_),
    .Y(_0615_));
 sg13g2_a221oi_1 _1414_ (.B2(_0523_),
    .C1(_0524_),
    .B1(_0490_),
    .A1(net49),
    .Y(_0616_),
    .A2(net50));
 sg13g2_nor3_1 _1415_ (.A(_0558_),
    .B(_0615_),
    .C(_0616_),
    .Y(_0617_));
 sg13g2_a21oi_1 _1416_ (.A1(_0133_),
    .A2(_0132_),
    .Y(_0618_),
    .B1(_0617_));
 sg13g2_a21o_1 _1417_ (.A2(_0614_),
    .A1(_0461_),
    .B1(_0618_),
    .X(_0619_));
 sg13g2_or3_1 _1418_ (.A(_0399_),
    .B(_0456_),
    .C(_0618_),
    .X(_0620_));
 sg13g2_nand2_2 _1419_ (.Y(_0621_),
    .A(_0619_),
    .B(_0620_));
 sg13g2_xor2_1 _1420_ (.B(_0134_),
    .A(_0135_),
    .X(_0622_));
 sg13g2_xnor2_1 _1421_ (.Y(_0623_),
    .A(_0621_),
    .B(_0622_));
 sg13g2_nand2_1 _1422_ (.Y(_0624_),
    .A(_0345_),
    .B(\cla_z[22] ));
 sg13g2_and2_1 _1423_ (.A(_0432_),
    .B(_0624_),
    .X(_0625_));
 sg13g2_o21ai_1 _1424_ (.B1(_0625_),
    .Y(_0626_),
    .A1(net24),
    .A2(_0623_));
 sg13g2_nor2_1 _1425_ (.A(_0372_),
    .B(_0339_),
    .Y(_0627_));
 sg13g2_nor2_1 _1426_ (.A(net20),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nor3_1 _1427_ (.A(net50),
    .B(net24),
    .C(_0560_),
    .Y(_0629_));
 sg13g2_nor3_1 _1428_ (.A(net49),
    .B(net24),
    .C(_0560_),
    .Y(_0630_));
 sg13g2_o21ai_1 _1429_ (.B1(_0533_),
    .Y(_0631_),
    .A1(_0629_),
    .A2(_0630_));
 sg13g2_nand3_1 _1430_ (.B(net25),
    .C(_0560_),
    .A(net50),
    .Y(_0632_));
 sg13g2_nand3_1 _1431_ (.B(_0352_),
    .C(_0560_),
    .A(net49),
    .Y(_0633_));
 sg13g2_a21o_1 _1432_ (.A2(_0633_),
    .A1(_0632_),
    .B1(_0533_),
    .X(_0634_));
 sg13g2_nor4_1 _1433_ (.A(net49),
    .B(net50),
    .C(net26),
    .D(_0560_),
    .Y(_0635_));
 sg13g2_and4_1 _1434_ (.A(net49),
    .B(net50),
    .C(_0352_),
    .D(_0560_),
    .X(_0636_));
 sg13g2_nor4_1 _1435_ (.A(net40),
    .B(_0583_),
    .C(_0635_),
    .D(_0636_),
    .Y(_0637_));
 sg13g2_nand3_1 _1436_ (.B(_0634_),
    .C(_0637_),
    .A(_0631_),
    .Y(_0638_));
 sg13g2_and3_1 _1437_ (.X(_0639_),
    .A(_0626_),
    .B(_0628_),
    .C(_0638_));
 sg13g2_or3_1 _1438_ (.A(_0587_),
    .B(_0610_),
    .C(_0639_),
    .X(_0067_));
 sg13g2_nor2_1 _1439_ (.A(net24),
    .B(_0623_),
    .Y(_0640_));
 sg13g2_nor2_1 _1440_ (.A(_0135_),
    .B(_0134_),
    .Y(_0641_));
 sg13g2_a21oi_1 _1441_ (.A1(_0619_),
    .A2(_0620_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_a21o_1 _1442_ (.A2(_0134_),
    .A1(_0135_),
    .B1(_0642_),
    .X(_0643_));
 sg13g2_xor2_1 _1443_ (.B(\io_sd._052_[23] ),
    .A(\io_sd._053_[23] ),
    .X(_0644_));
 sg13g2_xor2_1 _1444_ (.B(_0644_),
    .A(_0643_),
    .X(_0645_));
 sg13g2_a21oi_1 _1445_ (.A1(net32),
    .A2(_0624_),
    .Y(_0646_),
    .B1(net40));
 sg13g2_nand2_1 _1446_ (.Y(_0647_),
    .A(net33),
    .B(\cla_z[23] ));
 sg13g2_o21ai_1 _1447_ (.B1(net41),
    .Y(_0648_),
    .A1(net32),
    .A2(_0647_));
 sg13g2_nor2_1 _1448_ (.A(_0646_),
    .B(_0648_),
    .Y(_0649_));
 sg13g2_nor2_1 _1449_ (.A(_0297_),
    .B(_0649_),
    .Y(_0650_));
 sg13g2_a221oi_1 _1450_ (.B2(_0556_),
    .C1(_0650_),
    .B1(_0645_),
    .A1(_0372_),
    .Y(_0651_),
    .A2(_0640_));
 sg13g2_a221oi_1 _1451_ (.B2(_0591_),
    .C1(_0432_),
    .B1(_0369_),
    .A1(_0368_),
    .Y(_0652_),
    .A2(\cla_z[6] ));
 sg13g2_and2_1 _1452_ (.A(_0299_),
    .B(_0304_),
    .X(_0653_));
 sg13g2_a221oi_1 _1453_ (.B2(_0325_),
    .C1(_0341_),
    .B1(_0321_),
    .A1(_0328_),
    .Y(_0654_),
    .A2(_0329_));
 sg13g2_nand3b_1 _1454_ (.B(_0589_),
    .C(net56),
    .Y(_0655_),
    .A_N(_0326_));
 sg13g2_nand2_1 _1455_ (.Y(_0656_),
    .A(_0103_),
    .B(_0102_));
 sg13g2_and2_1 _1456_ (.A(_0656_),
    .B(_0322_),
    .X(_0657_));
 sg13g2_o21ai_1 _1457_ (.B1(_0657_),
    .Y(_0658_),
    .A1(_0588_),
    .A2(_0655_));
 sg13g2_a22oi_1 _1458_ (.Y(_0659_),
    .B1(_0654_),
    .B2(_0658_),
    .A2(\cla_z[7] ),
    .A1(_0345_));
 sg13g2_nand2_1 _1459_ (.Y(_0660_),
    .A(_0339_),
    .B(_0659_));
 sg13g2_nand3b_1 _1460_ (.B(_0653_),
    .C(_0660_),
    .Y(_0661_),
    .A_N(_0652_));
 sg13g2_and3_1 _1461_ (.X(_0662_),
    .A(net20),
    .B(_0303_),
    .C(_0605_));
 sg13g2_a22oi_1 _1462_ (.Y(_0663_),
    .B1(_0662_),
    .B2(_0604_),
    .A2(_0661_),
    .A1(net20));
 sg13g2_inv_1 _1463_ (.Y(_0664_),
    .A(_0419_));
 sg13g2_o21ai_1 _1464_ (.B1(_0664_),
    .Y(_0665_),
    .A1(_0438_),
    .A2(_0566_));
 sg13g2_a21oi_1 _1465_ (.A1(_0408_),
    .A2(_0665_),
    .Y(_0666_),
    .B1(_0451_));
 sg13g2_and3_1 _1466_ (.X(_0667_),
    .A(_0408_),
    .B(_0665_),
    .C(_0451_));
 sg13g2_or2_1 _1467_ (.X(_0668_),
    .B(_0667_),
    .A(_0666_));
 sg13g2_nor2b_1 _1468_ (.A(net43),
    .B_N(\cla_z[15] ),
    .Y(_0669_));
 sg13g2_nor3_1 _1469_ (.A(_0428_),
    .B(_0296_),
    .C(_0669_),
    .Y(_0670_));
 sg13g2_o21ai_1 _1470_ (.B1(_0670_),
    .Y(_0671_),
    .A1(net24),
    .A2(_0668_));
 sg13g2_nand2_1 _1471_ (.Y(_0672_),
    .A(_0663_),
    .B(_0671_));
 sg13g2_nand2_1 _1472_ (.Y(_0673_),
    .A(net17),
    .B(_0379_));
 sg13g2_o21ai_1 _1473_ (.B1(_0673_),
    .Y(_0068_),
    .A1(_0651_),
    .A2(_0672_));
 sg13g2_nand2_1 _1474_ (.Y(_0674_),
    .A(_0303_),
    .B(_0306_));
 sg13g2_nor4_1 _1475_ (.A(net24),
    .B(_0666_),
    .C(_0667_),
    .D(_0674_),
    .Y(_0675_));
 sg13g2_o21ai_1 _1476_ (.B1(_0428_),
    .Y(_0676_),
    .A1(_0432_),
    .A2(_0659_));
 sg13g2_and3_1 _1477_ (.X(_0677_),
    .A(_0303_),
    .B(_0306_),
    .C(_0669_));
 sg13g2_and3_1 _1478_ (.X(_0678_),
    .A(_0339_),
    .B(_0306_),
    .C(_0336_));
 sg13g2_or4_1 _1479_ (.A(_0675_),
    .B(_0676_),
    .C(_0677_),
    .D(_0678_),
    .X(_0679_));
 sg13g2_o21ai_1 _1480_ (.B1(net41),
    .Y(_0680_),
    .A1(_0296_),
    .A2(_0435_));
 sg13g2_nand3_1 _1481_ (.B(_0679_),
    .C(_0680_),
    .A(_0299_),
    .Y(_0681_));
 sg13g2_nor2_1 _1482_ (.A(net24),
    .B(_0644_),
    .Y(_0682_));
 sg13g2_nand2_1 _1483_ (.Y(_0683_),
    .A(net25),
    .B(_0644_));
 sg13g2_a21oi_1 _1484_ (.A1(_0134_),
    .A2(_0621_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_o21ai_1 _1485_ (.B1(_0135_),
    .Y(_0685_),
    .A1(_0134_),
    .A2(_0621_));
 sg13g2_mux2_1 _1486_ (.A0(_0682_),
    .A1(_0684_),
    .S(_0685_),
    .X(_0686_));
 sg13g2_nand3_1 _1487_ (.B(_0621_),
    .C(_0682_),
    .A(_0134_),
    .Y(_0687_));
 sg13g2_nand2_1 _1488_ (.Y(_0688_),
    .A(_0647_),
    .B(_0687_));
 sg13g2_nor3_1 _1489_ (.A(_0004_),
    .B(net20),
    .C(_0627_),
    .Y(_0689_));
 sg13g2_o21ai_1 _1490_ (.B1(_0689_),
    .Y(_0690_),
    .A1(_0686_),
    .A2(_0688_));
 sg13g2_nor2b_1 _1491_ (.A(net60),
    .B_N(net18),
    .Y(_0691_));
 sg13g2_nor3_1 _1492_ (.A(_0137_),
    .B(_0300_),
    .C(_0371_),
    .Y(_0692_));
 sg13g2_o21ai_1 _1493_ (.B1(net45),
    .Y(_0693_),
    .A1(_0691_),
    .A2(_0692_));
 sg13g2_nand3_1 _1494_ (.B(_0690_),
    .C(_0693_),
    .A(_0681_),
    .Y(_0069_));
 sg13g2_and2_1 _1495_ (.A(_0097_),
    .B(_0136_),
    .X(\rca.generate_adder_modules[0].fa.a ));
 sg13g2_nor2_1 _1496_ (.A(_0468_),
    .B(_0093_),
    .Y(\rca.generate_adder_modules[1].fa.b ));
 sg13g2_o21ai_1 _1497_ (.B1(_0643_),
    .Y(_0694_),
    .A1(\io_sd._053_[23] ),
    .A2(\io_sd._052_[23] ));
 sg13g2_nand2_1 _1498_ (.Y(_0695_),
    .A(\io_sd._053_[23] ),
    .B(\io_sd._052_[23] ));
 sg13g2_a21oi_1 _1499_ (.A1(_0694_),
    .A2(_0695_),
    .Y(\rca.generate_adder_modules[23].fa.c_out ),
    .B1(net39));
 sg13g2_and2_1 _1500_ (.A(net38),
    .B(\io_sd._053_[3] ),
    .X(\rca.generate_adder_modules[3].fa.b ));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _1509__73 (.L_HI(net73));
 sg13g2_buf_1 _1503_ (.A(net61),
    .X(uio_oe[0]));
 sg13g2_buf_1 _1504_ (.A(net62),
    .X(uio_oe[1]));
 sg13g2_buf_1 _1505_ (.A(net63),
    .X(uio_oe[2]));
 sg13g2_buf_1 _1506_ (.A(net64),
    .X(uio_oe[3]));
 sg13g2_buf_1 _1507_ (.A(net65),
    .X(uio_oe[4]));
 sg13g2_buf_1 _1508_ (.A(net66),
    .X(uio_oe[5]));
 sg13g2_buf_1 _1509_ (.A(net73),
    .X(uio_oe[6]));
 sg13g2_buf_1 _1510_ (.A(net74),
    .X(uio_oe[7]));
 sg13g2_buf_1 _1511_ (.A(net67),
    .X(uio_out[0]));
 sg13g2_buf_1 _1512_ (.A(net68),
    .X(uio_out[1]));
 sg13g2_buf_1 _1513_ (.A(net69),
    .X(uio_out[2]));
 sg13g2_buf_1 _1514_ (.A(net70),
    .X(uio_out[3]));
 sg13g2_buf_1 _1515_ (.A(net71),
    .X(uio_out[4]));
 sg13g2_buf_1 _1516_ (.A(net72),
    .X(uio_out[5]));
 sg13g2_buf_1 _1517_ (.A(\rca.generate_adder_modules[23].fa.c_out ),
    .X(net9));
 sg13g2_buf_1 \cla/_0684_  (.A(\rca.generate_adder_modules[22].fa.b ),
    .X(\cla/_0658_ ));
 sg13g2_buf_2 \cla/_0685_  (.A(\rca.generate_adder_modules[22].fa.a ),
    .X(\cla/_0659_ ));
 sg13g2_xnor2_1 \cla/_0686_  (.Y(\cla/_0660_ ),
    .A(\rca.generate_adder_modules[19].fa.b ),
    .B(\rca.generate_adder_modules[19].fa.a ));
 sg13g2_xnor2_1 \cla/_0687_  (.Y(\cla/_0661_ ),
    .A(\rca.generate_adder_modules[18].fa.b ),
    .B(\rca.generate_adder_modules[18].fa.a ));
 sg13g2_buf_2 \cla/_0688_  (.A(\rca.generate_adder_modules[17].fa.b ),
    .X(\cla/_0662_ ));
 sg13g2_buf_2 \cla/_0689_  (.A(\rca.generate_adder_modules[17].fa.a ),
    .X(\cla/_0663_ ));
 sg13g2_xnor2_1 \cla/_0690_  (.Y(\cla/_0664_ ),
    .A(\cla/_0662_ ),
    .B(\cla/_0663_ ));
 sg13g2_or3_1 \cla/_0691_  (.A(\cla/_0660_ ),
    .B(\cla/_0661_ ),
    .C(\cla/_0664_ ),
    .X(\cla/_0665_ ));
 sg13g2_buf_2 \cla/_0692_  (.A(\rca.generate_adder_modules[16].fa.b ),
    .X(\cla/_0666_ ));
 sg13g2_buf_2 \cla/_0693_  (.A(\rca.generate_adder_modules[16].fa.a ),
    .X(\cla/_0667_ ));
 sg13g2_xor2_1 \cla/_0694_  (.B(\cla/_0667_ ),
    .A(\cla/_0666_ ),
    .X(\cla/_0668_ ));
 sg13g2_buf_2 \cla/_0695_  (.A(\rca.generate_adder_modules[15].fa.b ),
    .X(\cla/_0669_ ));
 sg13g2_xor2_1 \cla/_0696_  (.B(\rca.generate_adder_modules[15].fa.a ),
    .A(\cla/_0669_ ),
    .X(\cla/_0670_ ));
 sg13g2_and2_1 \cla/_0697_  (.A(\cla/_0668_ ),
    .B(\cla/_0670_ ),
    .X(\cla/_0671_ ));
 sg13g2_buf_8 \cla/_0698_  (.A(\rca.generate_adder_modules[13].fa.a ),
    .X(\cla/_0672_ ));
 sg13g2_xnor2_1 \cla/_0699_  (.Y(\cla/_0673_ ),
    .A(\rca.generate_adder_modules[13].fa.b ),
    .B(\cla/_0672_ ));
 sg13g2_buf_2 \cla/_0700_  (.A(\rca.generate_adder_modules[11].fa.b ),
    .X(\cla/_0674_ ));
 sg13g2_buf_1 \cla/_0701_  (.A(\rca.generate_adder_modules[11].fa.a ),
    .X(\cla/_0675_ ));
 sg13g2_xnor2_1 \cla/_0702_  (.Y(\cla/_0676_ ),
    .A(\cla/_0674_ ),
    .B(\cla/_0675_ ));
 sg13g2_xnor2_1 \cla/_0703_  (.Y(\cla/_0677_ ),
    .A(\rca.generate_adder_modules[12].fa.b ),
    .B(\rca.generate_adder_modules[12].fa.a ));
 sg13g2_buf_2 \cla/_0704_  (.A(\rca.generate_adder_modules[10].fa.a ),
    .X(\cla/_0678_ ));
 sg13g2_nand2_1 \cla/_0705_  (.Y(\cla/_0679_ ),
    .A(\rca.generate_adder_modules[10].fa.b ),
    .B(\cla/_0678_ ));
 sg13g2_or4_1 \cla/_0706_  (.A(\cla/_0673_ ),
    .B(\cla/_0676_ ),
    .C(\cla/_0677_ ),
    .D(\cla/_0679_ ),
    .X(\cla/_0680_ ));
 sg13g2_nor2_1 \cla/_0707_  (.A(\rca.generate_adder_modules[14].fa.b ),
    .B(\rca.generate_adder_modules[14].fa.a ),
    .Y(\cla/_0681_ ));
 sg13g2_nand2_1 \cla/_0708_  (.Y(\cla/_0682_ ),
    .A(\rca.generate_adder_modules[14].fa.b ),
    .B(\rca.generate_adder_modules[14].fa.a ));
 sg13g2_o21ai_1 \cla/_0709_  (.B1(\cla/_0682_ ),
    .Y(\cla/_0683_ ),
    .A1(\cla/_0680_ ),
    .A2(\cla/_0681_ ));
 sg13g2_nand2_1 \cla/_0710_  (.Y(\cla/_0342_ ),
    .A(\cla/_0671_ ),
    .B(\cla/_0683_ ));
 sg13g2_xnor2_1 \cla/_0711_  (.Y(\cla/_0343_ ),
    .A(\cla/_0658_ ),
    .B(\cla/_0659_ ));
 sg13g2_buf_2 \cla/_0712_  (.A(\rca.generate_adder_modules[20].fa.b ),
    .X(\cla/_0344_ ));
 sg13g2_buf_2 \cla/_0713_  (.A(\rca.generate_adder_modules[20].fa.a ),
    .X(\cla/_0345_ ));
 sg13g2_xor2_1 \cla/_0714_  (.B(\cla/_0345_ ),
    .A(\cla/_0344_ ),
    .X(\cla/_0346_ ));
 sg13g2_buf_1 \cla/_0715_  (.A(\rca.generate_adder_modules[21].fa.b ),
    .X(\cla/_0347_ ));
 sg13g2_buf_1 \cla/_0716_  (.A(\rca.generate_adder_modules[21].fa.a ),
    .X(\cla/_0348_ ));
 sg13g2_xor2_1 \cla/_0717_  (.B(\cla/_0348_ ),
    .A(\cla/_0347_ ),
    .X(\cla/_0349_ ));
 sg13g2_and2_1 \cla/_0718_  (.A(\cla/_0346_ ),
    .B(\cla/_0349_ ),
    .X(\cla/_0350_ ));
 sg13g2_nand2b_1 \cla/_0719_  (.Y(\cla/_0351_ ),
    .B(\cla/_0350_ ),
    .A_N(\cla/_0343_ ));
 sg13g2_nor3_1 \cla/_0720_  (.A(\cla/_0665_ ),
    .B(\cla/_0342_ ),
    .C(\cla/_0351_ ),
    .Y(\cla/_0352_ ));
 sg13g2_xnor2_1 \cla/_0721_  (.Y(\cla/_0353_ ),
    .A(\rca.generate_adder_modules[10].fa.b ),
    .B(\cla/_0678_ ));
 sg13g2_xnor2_1 \cla/_0722_  (.Y(\cla/_0354_ ),
    .A(\rca.generate_adder_modules[9].fa.b ),
    .B(\rca.generate_adder_modules[9].fa.a ));
 sg13g2_buf_2 \cla/_0723_  (.A(\rca.generate_adder_modules[8].fa.a ),
    .X(\cla/_0355_ ));
 sg13g2_xnor2_1 \cla/_0724_  (.Y(\cla/_0356_ ),
    .A(\rca.generate_adder_modules[8].fa.b ),
    .B(\cla/_0355_ ));
 sg13g2_nor3_2 \cla/_0725_  (.A(\cla/_0353_ ),
    .B(\cla/_0354_ ),
    .C(\cla/_0356_ ),
    .Y(\cla/_0357_ ));
 sg13g2_nor3_2 \cla/_0726_  (.A(\cla/_0673_ ),
    .B(\cla/_0676_ ),
    .C(\cla/_0677_ ),
    .Y(\cla/_0358_ ));
 sg13g2_nor3_2 \cla/_0727_  (.A(\cla/_0660_ ),
    .B(\cla/_0661_ ),
    .C(\cla/_0664_ ),
    .Y(\cla/_0359_ ));
 sg13g2_xor2_1 \cla/_0728_  (.B(\rca.generate_adder_modules[14].fa.a ),
    .A(\rca.generate_adder_modules[14].fa.b ),
    .X(\cla/_0360_ ));
 sg13g2_and3_1 \cla/_0729_  (.X(\cla/_0361_ ),
    .A(\cla/_0360_ ),
    .B(\cla/_0668_ ),
    .C(\cla/_0670_ ));
 sg13g2_buf_2 \cla/_0730_  (.A(\cla/_0361_ ),
    .X(\cla/_0362_ ));
 sg13g2_nand4_1 \cla/_0731_  (.B(\cla/_0358_ ),
    .C(\cla/_0359_ ),
    .A(\cla/_0357_ ),
    .Y(\cla/_0363_ ),
    .D(\cla/_0362_ ));
 sg13g2_xnor2_1 \cla/_0732_  (.Y(\cla/_0364_ ),
    .A(\rca.generate_adder_modules[7].fa.b ),
    .B(\rca.generate_adder_modules[7].fa.a ));
 sg13g2_xnor2_1 \cla/_0733_  (.Y(\cla/_0365_ ),
    .A(\rca.generate_adder_modules[6].fa.b ),
    .B(\rca.generate_adder_modules[6].fa.a ));
 sg13g2_xnor2_1 \cla/_0734_  (.Y(\cla/_0366_ ),
    .A(\rca.generate_adder_modules[5].fa.b ),
    .B(\rca.generate_adder_modules[5].fa.a ));
 sg13g2_buf_2 \cla/_0735_  (.A(\rca.generate_adder_modules[4].fa.b ),
    .X(\cla/_0367_ ));
 sg13g2_buf_2 \cla/_0736_  (.A(\rca.generate_adder_modules[4].fa.a ),
    .X(\cla/_0368_ ));
 sg13g2_nand2_1 \cla/_0737_  (.Y(\cla/_0369_ ),
    .A(\cla/_0367_ ),
    .B(\cla/_0368_ ));
 sg13g2_nor4_1 \cla/_0738_  (.A(\cla/_0364_ ),
    .B(\cla/_0365_ ),
    .C(\cla/_0366_ ),
    .D(\cla/_0369_ ),
    .Y(\cla/_0370_ ));
 sg13g2_nand2b_1 \cla/_0739_  (.Y(\cla/_0371_ ),
    .B(\cla/_0370_ ),
    .A_N(\cla/_0363_ ));
 sg13g2_xnor2_1 \cla/_0740_  (.Y(\cla/_0372_ ),
    .A(\cla/_0367_ ),
    .B(\cla/_0368_ ));
 sg13g2_nor4_2 \cla/_0741_  (.A(\cla/_0364_ ),
    .B(\cla/_0365_ ),
    .C(\cla/_0366_ ),
    .Y(\cla/_0373_ ),
    .D(\cla/_0372_ ));
 sg13g2_and2_1 \cla/_0742_  (.A(\rca.generate_adder_modules[3].fa.b ),
    .B(\rca.generate_adder_modules[3].fa.a ),
    .X(\cla/_0374_ ));
 sg13g2_buf_1 \cla/_0743_  (.A(\cla/_0374_ ),
    .X(\cla/_0375_ ));
 sg13g2_nand2_1 \cla/_0744_  (.Y(\cla/_0376_ ),
    .A(\cla/_0373_ ),
    .B(\cla/_0375_ ));
 sg13g2_xnor2_1 \cla/_0745_  (.Y(\cla/_0377_ ),
    .A(\rca.generate_adder_modules[3].fa.b ),
    .B(\rca.generate_adder_modules[3].fa.a ));
 sg13g2_nand2_1 \cla/_0746_  (.Y(\cla/_0378_ ),
    .A(\rca.generate_adder_modules[2].fa.b ),
    .B(\rca.generate_adder_modules[2].fa.a ));
 sg13g2_nor2_1 \cla/_0747_  (.A(\cla/_0377_ ),
    .B(\cla/_0378_ ),
    .Y(\cla/_0379_ ));
 sg13g2_xnor2_1 \cla/_0748_  (.Y(\cla/_0380_ ),
    .A(\rca.generate_adder_modules[2].fa.b ),
    .B(\rca.generate_adder_modules[2].fa.a ));
 sg13g2_nor2_1 \cla/_0749_  (.A(\rca.generate_adder_modules[1].fa.b ),
    .B(\rca.generate_adder_modules[1].fa.a ),
    .Y(\cla/_0381_ ));
 sg13g2_a22oi_1 \cla/_0750_  (.Y(\cla/_0382_ ),
    .B1(\rca.generate_adder_modules[1].fa.b ),
    .B2(\rca.generate_adder_modules[1].fa.a ),
    .A2(\rca.generate_adder_modules[0].fa.a ),
    .A1(\rca.generate_adder_modules[0].fa.b ));
 sg13g2_nor4_1 \cla/_0751_  (.A(\cla/_0377_ ),
    .B(\cla/_0380_ ),
    .C(\cla/_0381_ ),
    .D(\cla/_0382_ ),
    .Y(\cla/_0383_ ));
 sg13g2_o21ai_1 \cla/_0752_  (.B1(\cla/_0373_ ),
    .Y(\cla/_0384_ ),
    .A1(\cla/_0379_ ),
    .A2(\cla/_0383_ ));
 sg13g2_a21o_1 \cla/_0753_  (.A2(\cla/_0384_ ),
    .A1(\cla/_0376_ ),
    .B1(\cla/_0363_ ),
    .X(\cla/_0385_ ));
 sg13g2_nand2_1 \cla/_0754_  (.Y(\cla/_0386_ ),
    .A(\cla/_0346_ ),
    .B(\cla/_0349_ ));
 sg13g2_a21oi_1 \cla/_0755_  (.A1(\cla/_0371_ ),
    .A2(\cla/_0385_ ),
    .Y(\cla/_0387_ ),
    .B1(\cla/_0386_ ));
 sg13g2_xnor2_1 \cla/_0756_  (.Y(\cla/_0388_ ),
    .A(\cla/_0666_ ),
    .B(\cla/_0667_ ));
 sg13g2_nor2_1 \cla/_0757_  (.A(\cla/_0665_ ),
    .B(\cla/_0388_ ),
    .Y(\cla/_0389_ ));
 sg13g2_and2_1 \cla/_0758_  (.A(\cla/_0669_ ),
    .B(\rca.generate_adder_modules[15].fa.a ),
    .X(\cla/_0390_ ));
 sg13g2_nor2_1 \cla/_0759_  (.A(\rca.generate_adder_modules[19].fa.b ),
    .B(\rca.generate_adder_modules[19].fa.a ),
    .Y(\cla/_0391_ ));
 sg13g2_nand2_1 \cla/_0760_  (.Y(\cla/_0392_ ),
    .A(\rca.generate_adder_modules[18].fa.b ),
    .B(\rca.generate_adder_modules[18].fa.a ));
 sg13g2_nand2_1 \cla/_0761_  (.Y(\cla/_0393_ ),
    .A(\rca.generate_adder_modules[19].fa.b ),
    .B(\rca.generate_adder_modules[19].fa.a ));
 sg13g2_o21ai_1 \cla/_0762_  (.B1(\cla/_0393_ ),
    .Y(\cla/_0394_ ),
    .A1(\cla/_0391_ ),
    .A2(\cla/_0392_ ));
 sg13g2_a221oi_1 \cla/_0763_  (.B2(\cla/_0390_ ),
    .C1(\cla/_0394_ ),
    .B1(\cla/_0389_ ),
    .A1(\cla/_0347_ ),
    .Y(\cla/_0395_ ),
    .A2(\cla/_0348_ ));
 sg13g2_a21oi_1 \cla/_0764_  (.A1(\cla/_0347_ ),
    .A2(\cla/_0348_ ),
    .Y(\cla/_0396_ ),
    .B1(\cla/_0346_ ));
 sg13g2_nor2_1 \cla/_0765_  (.A(\cla/_0347_ ),
    .B(\cla/_0348_ ),
    .Y(\cla/_0397_ ));
 sg13g2_nor3_1 \cla/_0766_  (.A(\cla/_0395_ ),
    .B(\cla/_0396_ ),
    .C(\cla/_0397_ ),
    .Y(\cla/_0398_ ));
 sg13g2_or3_1 \cla/_0767_  (.A(\cla/_0352_ ),
    .B(\cla/_0387_ ),
    .C(\cla/_0398_ ),
    .X(\cla/_0399_ ));
 sg13g2_a21oi_1 \cla/_0768_  (.A1(\cla/_0658_ ),
    .A2(\cla/_0659_ ),
    .Y(\cla/_0400_ ),
    .B1(\cla/_0399_ ));
 sg13g2_nor2_1 \cla/_0769_  (.A(\rca.generate_adder_modules[23].fa.b ),
    .B(\rca.generate_adder_modules[23].fa.a ),
    .Y(\cla/_0401_ ));
 sg13g2_nor2_1 \cla/_0770_  (.A(\cla/_0658_ ),
    .B(\cla/_0659_ ),
    .Y(\cla/_0402_ ));
 sg13g2_or2_1 \cla/_0771_  (.X(\cla/_0403_ ),
    .B(\cla/_0402_ ),
    .A(\cla/_0401_ ));
 sg13g2_inv_1 \cla/_0772_  (.Y(\cla/_0404_ ),
    .A(\cla/_0349_ ));
 sg13g2_xnor2_1 \cla/_0773_  (.Y(\cla/_0405_ ),
    .A(\rca.generate_adder_modules[23].fa.b ),
    .B(\rca.generate_adder_modules[23].fa.a ));
 sg13g2_nor3_1 \cla/_0774_  (.A(\cla/_0404_ ),
    .B(\cla/_0343_ ),
    .C(\cla/_0405_ ),
    .Y(\cla/_0406_ ));
 sg13g2_inv_1 \cla/_0775_  (.Y(\cla/_0407_ ),
    .A(\cla/_0345_ ));
 sg13g2_and2_1 \cla/_0776_  (.A(\rca.generate_adder_modules[8].fa.b ),
    .B(\cla/_0355_ ),
    .X(\cla/_0408_ ));
 sg13g2_buf_1 \cla/_0777_  (.A(\cla/_0408_ ),
    .X(\cla/_0409_ ));
 sg13g2_nor4_2 \cla/_0778_  (.A(\cla/_0353_ ),
    .B(\cla/_0354_ ),
    .C(\cla/_0676_ ),
    .Y(\cla/_0410_ ),
    .D(\cla/_0677_ ));
 sg13g2_and2_1 \cla/_0779_  (.A(\rca.generate_adder_modules[12].fa.b ),
    .B(\rca.generate_adder_modules[12].fa.a ),
    .X(\cla/_0411_ ));
 sg13g2_buf_1 \cla/_0780_  (.A(\cla/_0411_ ),
    .X(\cla/_0412_ ));
 sg13g2_a21oi_1 \cla/_0781_  (.A1(\cla/_0409_ ),
    .A2(\cla/_0410_ ),
    .Y(\cla/_0413_ ),
    .B1(\cla/_0412_ ));
 sg13g2_xor2_1 \cla/_0782_  (.B(\cla/_0672_ ),
    .A(\rca.generate_adder_modules[13].fa.b ),
    .X(\cla/_0414_ ));
 sg13g2_nand2_1 \cla/_0783_  (.Y(\cla/_0415_ ),
    .A(\cla/_0414_ ),
    .B(\cla/_0362_ ));
 sg13g2_nor3_1 \cla/_0784_  (.A(\cla/_0665_ ),
    .B(\cla/_0413_ ),
    .C(\cla/_0415_ ),
    .Y(\cla/_0416_ ));
 sg13g2_nand2_1 \cla/_0785_  (.Y(\cla/_0417_ ),
    .A(\cla/_0359_ ),
    .B(\cla/_0362_ ));
 sg13g2_nor2_2 \cla/_0786_  (.A(\cla/_0673_ ),
    .B(\cla/_0677_ ),
    .Y(\cla/_0418_ ));
 sg13g2_xor2_1 \cla/_0787_  (.B(\cla/_0678_ ),
    .A(\rca.generate_adder_modules[10].fa.b ),
    .X(\cla/_0419_ ));
 sg13g2_xor2_1 \cla/_0788_  (.B(net23),
    .A(\cla/_0674_ ),
    .X(\cla/_0420_ ));
 sg13g2_and4_1 \cla/_0789_  (.A(\rca.generate_adder_modules[9].fa.b ),
    .B(\rca.generate_adder_modules[9].fa.a ),
    .C(\cla/_0419_ ),
    .D(\cla/_0420_ ),
    .X(\cla/_0421_ ));
 sg13g2_buf_1 \cla/_0790_  (.A(\cla/_0421_ ),
    .X(\cla/_0422_ ));
 sg13g2_and2_1 \cla/_0791_  (.A(\rca.generate_adder_modules[13].fa.b ),
    .B(\cla/_0672_ ),
    .X(\cla/_0423_ ));
 sg13g2_buf_1 \cla/_0792_  (.A(\cla/_0423_ ),
    .X(\cla/_0424_ ));
 sg13g2_a21oi_1 \cla/_0793_  (.A1(\cla/_0418_ ),
    .A2(\cla/_0422_ ),
    .Y(\cla/_0425_ ),
    .B1(\cla/_0424_ ));
 sg13g2_nor2_2 \cla/_0794_  (.A(\cla/_0660_ ),
    .B(\cla/_0661_ ),
    .Y(\cla/_0426_ ));
 sg13g2_nand2_1 \cla/_0795_  (.Y(\cla/_0427_ ),
    .A(\cla/_0666_ ),
    .B(\cla/_0667_ ));
 sg13g2_nor2_1 \cla/_0796_  (.A(\cla/_0662_ ),
    .B(\cla/_0663_ ),
    .Y(\cla/_0428_ ));
 sg13g2_nand2_1 \cla/_0797_  (.Y(\cla/_0429_ ),
    .A(\cla/_0662_ ),
    .B(\cla/_0663_ ));
 sg13g2_o21ai_1 \cla/_0798_  (.B1(\cla/_0429_ ),
    .Y(\cla/_0430_ ),
    .A1(\cla/_0427_ ),
    .A2(\cla/_0428_ ));
 sg13g2_nand2_1 \cla/_0799_  (.Y(\cla/_0431_ ),
    .A(\cla/_0426_ ),
    .B(\cla/_0430_ ));
 sg13g2_o21ai_1 \cla/_0800_  (.B1(\cla/_0431_ ),
    .Y(\cla/_0432_ ),
    .A1(\cla/_0417_ ),
    .A2(\cla/_0425_ ));
 sg13g2_xor2_1 \cla/_0801_  (.B(\rca.generate_adder_modules[12].fa.a ),
    .A(\rca.generate_adder_modules[12].fa.b ),
    .X(\cla/_0433_ ));
 sg13g2_nand4_1 \cla/_0802_  (.B(net23),
    .C(\cla/_0414_ ),
    .A(\cla/_0674_ ),
    .Y(\cla/_0434_ ),
    .D(\cla/_0433_ ));
 sg13g2_nor2_1 \cla/_0803_  (.A(\cla/_0417_ ),
    .B(\cla/_0434_ ),
    .Y(\cla/_0435_ ));
 sg13g2_or2_1 \cla/_0804_  (.X(\cla/_0436_ ),
    .B(\rca.generate_adder_modules[7].fa.a ),
    .A(\rca.generate_adder_modules[7].fa.b ));
 sg13g2_nor2_1 \cla/_0805_  (.A(\rca.generate_adder_modules[6].fa.b ),
    .B(\rca.generate_adder_modules[6].fa.a ),
    .Y(\cla/_0437_ ));
 sg13g2_nand2_1 \cla/_0806_  (.Y(\cla/_0438_ ),
    .A(\rca.generate_adder_modules[5].fa.b ),
    .B(\rca.generate_adder_modules[5].fa.a ));
 sg13g2_a22oi_1 \cla/_0807_  (.Y(\cla/_0439_ ),
    .B1(\rca.generate_adder_modules[7].fa.b ),
    .B2(\rca.generate_adder_modules[7].fa.a ),
    .A2(\rca.generate_adder_modules[6].fa.a ),
    .A1(\rca.generate_adder_modules[6].fa.b ));
 sg13g2_o21ai_1 \cla/_0808_  (.B1(\cla/_0439_ ),
    .Y(\cla/_0440_ ),
    .A1(\cla/_0437_ ),
    .A2(\cla/_0438_ ));
 sg13g2_nand2_1 \cla/_0809_  (.Y(\cla/_0441_ ),
    .A(\cla/_0436_ ),
    .B(\cla/_0440_ ));
 sg13g2_nor2_1 \cla/_0810_  (.A(\cla/_0363_ ),
    .B(\cla/_0441_ ),
    .Y(\cla/_0442_ ));
 sg13g2_nor4_1 \cla/_0811_  (.A(\cla/_0416_ ),
    .B(\cla/_0432_ ),
    .C(\cla/_0435_ ),
    .D(\cla/_0442_ ),
    .Y(\cla/_0443_ ));
 sg13g2_inv_1 \cla/_0812_  (.Y(\cla/_0444_ ),
    .A(\cla/_0344_ ));
 sg13g2_a21oi_1 \cla/_0813_  (.A1(\cla/_0407_ ),
    .A2(\cla/_0443_ ),
    .Y(\cla/_0445_ ),
    .B1(\cla/_0444_ ));
 sg13g2_inv_1 \cla/_0814_  (.Y(\cla/_0446_ ),
    .A(\cla/_0406_ ));
 sg13g2_nor3_1 \cla/_0815_  (.A(\cla/_0407_ ),
    .B(\cla/_0446_ ),
    .C(\cla/_0443_ ),
    .Y(\cla/_0447_ ));
 sg13g2_a221oi_1 \cla/_0816_  (.B2(\cla/_0445_ ),
    .C1(\cla/_0447_ ),
    .B1(\cla/_0406_ ),
    .A1(\rca.generate_adder_modules[23].fa.b ),
    .Y(\cla/_0448_ ),
    .A2(\rca.generate_adder_modules[23].fa.a ));
 sg13g2_o21ai_1 \cla/_0817_  (.B1(\cla/_0448_ ),
    .Y(\cla/_0341_ ),
    .A1(\cla/_0400_ ),
    .A2(\cla/_0403_ ));
 sg13g2_xor2_1 \cla/_0818_  (.B(\rca.generate_adder_modules[0].fa.a ),
    .A(\rca.generate_adder_modules[0].fa.b ),
    .X(\cla/generate_adder_modules[0].fa_i._2_ ));
 sg13g2_inv_1 \cla/_0819_  (.Y(\cla/_0449_ ),
    .A(\rca.generate_adder_modules[9].fa.a ));
 sg13g2_nor2_1 \cla/_0820_  (.A(\cla/_0377_ ),
    .B(\cla/_0380_ ),
    .Y(\cla/_0450_ ));
 sg13g2_nor2_1 \cla/_0821_  (.A(\cla/_0381_ ),
    .B(\cla/_0382_ ),
    .Y(\cla/_0451_ ));
 sg13g2_nand3_1 \cla/_0822_  (.B(\cla/_0450_ ),
    .C(\cla/_0451_ ),
    .A(\cla/_0373_ ),
    .Y(\cla/_0452_ ));
 sg13g2_nor2_1 \cla/_0823_  (.A(\rca.generate_adder_modules[3].fa.b ),
    .B(\rca.generate_adder_modules[3].fa.a ),
    .Y(\cla/_0453_ ));
 sg13g2_a22oi_1 \cla/_0824_  (.Y(\cla/_0454_ ),
    .B1(\cla/_0367_ ),
    .B2(\cla/_0368_ ),
    .A2(\rca.generate_adder_modules[3].fa.a ),
    .A1(\rca.generate_adder_modules[3].fa.b ));
 sg13g2_o21ai_1 \cla/_0825_  (.B1(\cla/_0454_ ),
    .Y(\cla/_0455_ ),
    .A1(\cla/_0378_ ),
    .A2(\cla/_0453_ ));
 sg13g2_nor2_1 \cla/_0826_  (.A(\cla/_0367_ ),
    .B(\cla/_0368_ ),
    .Y(\cla/_0456_ ));
 sg13g2_nor4_1 \cla/_0827_  (.A(\cla/_0364_ ),
    .B(\cla/_0365_ ),
    .C(\cla/_0366_ ),
    .D(\cla/_0456_ ),
    .Y(\cla/_0457_ ));
 sg13g2_a22oi_1 \cla/_0828_  (.Y(\cla/_0458_ ),
    .B1(\cla/_0455_ ),
    .B2(\cla/_0457_ ),
    .A2(\cla/_0440_ ),
    .A1(\cla/_0436_ ));
 sg13g2_nand2_2 \cla/_0829_  (.Y(\cla/_0459_ ),
    .A(\cla/_0452_ ),
    .B(\cla/_0458_ ));
 sg13g2_nand2_1 \cla/_0830_  (.Y(\cla/_0460_ ),
    .A(\cla/_0355_ ),
    .B(\cla/_0459_ ));
 sg13g2_o21ai_1 \cla/_0831_  (.B1(\rca.generate_adder_modules[8].fa.b ),
    .Y(\cla/_0461_ ),
    .A1(\cla/_0355_ ),
    .A2(\cla/_0459_ ));
 sg13g2_nand3_1 \cla/_0832_  (.B(\cla/_0460_ ),
    .C(\cla/_0461_ ),
    .A(\cla/_0449_ ),
    .Y(\cla/_0462_ ));
 sg13g2_a21oi_1 \cla/_0833_  (.A1(\cla/_0460_ ),
    .A2(\cla/_0461_ ),
    .Y(\cla/_0463_ ),
    .B1(\cla/_0449_ ));
 sg13g2_a21oi_1 \cla/_0834_  (.A1(\rca.generate_adder_modules[9].fa.b ),
    .A2(\cla/_0462_ ),
    .Y(\cla/_0464_ ),
    .B1(\cla/_0463_ ));
 sg13g2_xnor2_1 \cla/_0835_  (.Y(\cla/generate_adder_modules[10].fa_i.s ),
    .A(\cla/_0419_ ),
    .B(\cla/_0464_ ));
 sg13g2_or2_1 \cla/_0836_  (.X(\cla/_0465_ ),
    .B(\cla/_0678_ ),
    .A(\rca.generate_adder_modules[10].fa.b ));
 sg13g2_nand2_1 \cla/_0837_  (.Y(\cla/_0466_ ),
    .A(\rca.generate_adder_modules[9].fa.a ),
    .B(\cla/_0409_ ));
 sg13g2_o21ai_1 \cla/_0838_  (.B1(\rca.generate_adder_modules[9].fa.b ),
    .Y(\cla/_0467_ ),
    .A1(\rca.generate_adder_modules[9].fa.a ),
    .A2(\cla/_0409_ ));
 sg13g2_nand3_1 \cla/_0839_  (.B(\cla/_0466_ ),
    .C(\cla/_0467_ ),
    .A(\cla/_0679_ ),
    .Y(\cla/_0468_ ));
 sg13g2_a22oi_1 \cla/_0840_  (.Y(\cla/_0469_ ),
    .B1(\cla/_0465_ ),
    .B2(\cla/_0468_ ),
    .A2(\cla/_0459_ ),
    .A1(\cla/_0357_ ));
 sg13g2_xnor2_1 \cla/_0841_  (.Y(\cla/generate_adder_modules[11].fa_i.s ),
    .A(\cla/_0420_ ),
    .B(\cla/_0469_ ));
 sg13g2_inv_1 \cla/_0842_  (.Y(\cla/_0470_ ),
    .A(\cla/_0674_ ));
 sg13g2_inv_1 \cla/_0843_  (.Y(\cla/_0471_ ),
    .A(net23));
 sg13g2_a21oi_1 \cla/_0844_  (.A1(\cla/_0470_ ),
    .A2(\cla/_0471_ ),
    .Y(\cla/_0472_ ),
    .B1(\cla/_0469_ ));
 sg13g2_a21oi_1 \cla/_0845_  (.A1(\cla/_0674_ ),
    .A2(net23),
    .Y(\cla/_0473_ ),
    .B1(\cla/_0472_ ));
 sg13g2_xnor2_1 \cla/_0846_  (.Y(\cla/generate_adder_modules[12].fa_i.s ),
    .A(\cla/_0433_ ),
    .B(\cla/_0473_ ));
 sg13g2_inv_1 \cla/_0847_  (.Y(\cla/_0474_ ),
    .A(\cla/_0355_ ));
 sg13g2_inv_1 \cla/_0848_  (.Y(\cla/_0475_ ),
    .A(\cla/_0452_ ));
 sg13g2_o21ai_1 \cla/_0849_  (.B1(\rca.generate_adder_modules[8].fa.b ),
    .Y(\cla/_0476_ ),
    .A1(\cla/_0355_ ),
    .A2(\cla/_0475_ ));
 sg13g2_o21ai_1 \cla/_0850_  (.B1(\cla/_0476_ ),
    .Y(\cla/_0477_ ),
    .A1(\cla/_0474_ ),
    .A2(\cla/_0452_ ));
 sg13g2_or3_1 \cla/_0851_  (.A(\cla/_0353_ ),
    .B(\cla/_0354_ ),
    .C(\cla/_0356_ ),
    .X(\cla/_0478_ ));
 sg13g2_buf_1 \cla/_0852_  (.A(\cla/_0478_ ),
    .X(\cla/_0479_ ));
 sg13g2_o21ai_1 \cla/_0853_  (.B1(\cla/_0679_ ),
    .Y(\cla/_0480_ ),
    .A1(\cla/_0479_ ),
    .A2(\cla/_0458_ ));
 sg13g2_nor3_1 \cla/_0854_  (.A(\cla/_0412_ ),
    .B(\cla/_0422_ ),
    .C(\cla/_0480_ ),
    .Y(\cla/_0481_ ));
 sg13g2_nor2_1 \cla/_0855_  (.A(\rca.generate_adder_modules[12].fa.b ),
    .B(\rca.generate_adder_modules[12].fa.a ),
    .Y(\cla/_0482_ ));
 sg13g2_a21oi_1 \cla/_0856_  (.A1(\cla/_0471_ ),
    .A2(\cla/_0481_ ),
    .Y(\cla/_0483_ ),
    .B1(\cla/_0482_ ));
 sg13g2_o21ai_1 \cla/_0857_  (.B1(\rca.generate_adder_modules[12].fa.b ),
    .Y(\cla/_0484_ ),
    .A1(\rca.generate_adder_modules[12].fa.a ),
    .A2(\cla/_0422_ ));
 sg13g2_and2_1 \cla/_0858_  (.A(\cla/_0471_ ),
    .B(\cla/_0484_ ),
    .X(\cla/_0485_ ));
 sg13g2_o21ai_1 \cla/_0859_  (.B1(\cla/_0470_ ),
    .Y(\cla/_0486_ ),
    .A1(\cla/_0481_ ),
    .A2(\cla/_0485_ ));
 sg13g2_a22oi_1 \cla/_0860_  (.Y(\cla/_0487_ ),
    .B1(\cla/_0483_ ),
    .B2(\cla/_0486_ ),
    .A2(\cla/_0477_ ),
    .A1(\cla/_0410_ ));
 sg13g2_xnor2_1 \cla/_0861_  (.Y(\cla/generate_adder_modules[13].fa_i.s ),
    .A(\cla/_0414_ ),
    .B(\cla/_0487_ ));
 sg13g2_xnor2_1 \cla/_0862_  (.Y(\cla/_0488_ ),
    .A(\rca.generate_adder_modules[14].fa.b ),
    .B(\rca.generate_adder_modules[14].fa.a ));
 sg13g2_o21ai_1 \cla/_0863_  (.B1(\cla/_0418_ ),
    .Y(\cla/_0489_ ),
    .A1(net23),
    .A2(\cla/_0480_ ));
 sg13g2_a21oi_1 \cla/_0864_  (.A1(net23),
    .A2(\cla/_0480_ ),
    .Y(\cla/_0490_ ),
    .B1(\cla/_0674_ ));
 sg13g2_a21o_1 \cla/_0865_  (.A2(\cla/_0410_ ),
    .A1(\cla/_0409_ ),
    .B1(\cla/_0412_ ),
    .X(\cla/_0491_ ));
 sg13g2_a21o_1 \cla/_0866_  (.A2(\cla/_0491_ ),
    .A1(\cla/_0672_ ),
    .B1(\rca.generate_adder_modules[13].fa.b ),
    .X(\cla/_0492_ ));
 sg13g2_nand2b_1 \cla/_0867_  (.Y(\cla/_0493_ ),
    .B(\cla/_0413_ ),
    .A_N(\cla/_0672_ ));
 sg13g2_nand2_1 \cla/_0868_  (.Y(\cla/_0494_ ),
    .A(\cla/_0418_ ),
    .B(\cla/_0422_ ));
 sg13g2_nand4_1 \cla/_0869_  (.B(\cla/_0358_ ),
    .C(\cla/_0373_ ),
    .A(\cla/_0357_ ),
    .Y(\cla/_0495_ ),
    .D(\cla/_0383_ ));
 sg13g2_nand2_1 \cla/_0870_  (.Y(\cla/_0496_ ),
    .A(\cla/_0494_ ),
    .B(\cla/_0495_ ));
 sg13g2_a21oi_1 \cla/_0871_  (.A1(\cla/_0492_ ),
    .A2(\cla/_0493_ ),
    .Y(\cla/_0497_ ),
    .B1(\cla/_0496_ ));
 sg13g2_o21ai_1 \cla/_0872_  (.B1(\cla/_0497_ ),
    .Y(\cla/_0498_ ),
    .A1(\cla/_0489_ ),
    .A2(\cla/_0490_ ));
 sg13g2_xnor2_1 \cla/_0873_  (.Y(\cla/generate_adder_modules[14].fa_i.s ),
    .A(\cla/_0488_ ),
    .B(\cla/_0498_ ));
 sg13g2_nand3_1 \cla/_0874_  (.B(\cla/_0420_ ),
    .C(\cla/_0433_ ),
    .A(\cla/_0414_ ),
    .Y(\cla/_0499_ ));
 sg13g2_nor3_1 \cla/_0875_  (.A(\cla/_0479_ ),
    .B(\cla/_0499_ ),
    .C(\cla/_0458_ ),
    .Y(\cla/_0500_ ));
 sg13g2_nand2b_1 \cla/_0876_  (.Y(\cla/_0501_ ),
    .B(\cla/_0497_ ),
    .A_N(\cla/_0500_ ));
 sg13g2_and3_1 \cla/_0877_  (.X(\cla/_0502_ ),
    .A(\cla/_0682_ ),
    .B(\cla/_0680_ ),
    .C(\cla/_0434_ ));
 sg13g2_nor2_1 \cla/_0878_  (.A(\cla/_0681_ ),
    .B(\cla/_0502_ ),
    .Y(\cla/_0503_ ));
 sg13g2_a21oi_1 \cla/_0879_  (.A1(\cla/_0360_ ),
    .A2(\cla/_0501_ ),
    .Y(\cla/_0504_ ),
    .B1(\cla/_0503_ ));
 sg13g2_xnor2_1 \cla/_0880_  (.Y(\cla/generate_adder_modules[15].fa_i.s ),
    .A(\cla/_0670_ ),
    .B(\cla/_0504_ ));
 sg13g2_nand2_2 \cla/_0881_  (.Y(\cla/_0505_ ),
    .A(\cla/_0360_ ),
    .B(\cla/_0670_ ));
 sg13g2_and2_1 \cla/_0882_  (.A(\cla/_0360_ ),
    .B(\cla/_0670_ ),
    .X(\cla/_0506_ ));
 sg13g2_inv_1 \cla/_0883_  (.Y(\cla/_0507_ ),
    .A(\rca.generate_adder_modules[15].fa.a ));
 sg13g2_o21ai_1 \cla/_0884_  (.B1(\cla/_0507_ ),
    .Y(\cla/_0508_ ),
    .A1(\cla/_0681_ ),
    .A2(\cla/_0502_ ));
 sg13g2_nor3_1 \cla/_0885_  (.A(\cla/_0507_ ),
    .B(\cla/_0681_ ),
    .C(\cla/_0502_ ),
    .Y(\cla/_0509_ ));
 sg13g2_a221oi_1 \cla/_0886_  (.B2(\cla/_0669_ ),
    .C1(\cla/_0509_ ),
    .B1(\cla/_0508_ ),
    .A1(\cla/_0506_ ),
    .Y(\cla/_0510_ ),
    .A2(\cla/_0500_ ));
 sg13g2_o21ai_1 \cla/_0887_  (.B1(\cla/_0510_ ),
    .Y(\cla/_0511_ ),
    .A1(\cla/_0505_ ),
    .A2(\cla/_0497_ ));
 sg13g2_xnor2_1 \cla/_0888_  (.Y(\cla/generate_adder_modules[16].fa_i.s ),
    .A(\cla/_0388_ ),
    .B(\cla/_0511_ ));
 sg13g2_inv_1 \cla/_0889_  (.Y(\cla/_0512_ ),
    .A(\cla/_0666_ ));
 sg13g2_inv_1 \cla/_0890_  (.Y(\cla/_0513_ ),
    .A(\cla/_0667_ ));
 sg13g2_o21ai_1 \cla/_0891_  (.B1(\cla/_0506_ ),
    .Y(\cla/_0514_ ),
    .A1(\cla/_0424_ ),
    .A2(\cla/_0496_ ));
 sg13g2_a221oi_1 \cla/_0892_  (.B2(\cla/_0514_ ),
    .C1(\cla/_0664_ ),
    .B1(\cla/_0510_ ),
    .A1(\cla/_0512_ ),
    .Y(\cla/_0515_ ),
    .A2(\cla/_0513_ ));
 sg13g2_and2_1 \cla/_0893_  (.A(\cla/_0414_ ),
    .B(\cla/_0362_ ),
    .X(\cla/_0516_ ));
 sg13g2_nand2_1 \cla/_0894_  (.Y(\cla/_0517_ ),
    .A(\cla/_0513_ ),
    .B(\cla/_0664_ ));
 sg13g2_nand2_1 \cla/_0895_  (.Y(\cla/_0518_ ),
    .A(\cla/_0512_ ),
    .B(\cla/_0664_ ));
 sg13g2_nand2_1 \cla/_0896_  (.Y(\cla/_0519_ ),
    .A(\cla/_0510_ ),
    .B(\cla/_0514_ ));
 sg13g2_a221oi_1 \cla/_0897_  (.B2(\cla/_0518_ ),
    .C1(\cla/_0519_ ),
    .B1(\cla/_0517_ ),
    .A1(\cla/_0491_ ),
    .Y(\cla/_0520_ ),
    .A2(\cla/_0516_ ));
 sg13g2_xor2_1 \cla/_0898_  (.B(\cla/_0663_ ),
    .A(\cla/_0662_ ),
    .X(\cla/_0521_ ));
 sg13g2_nor3_1 \cla/_0899_  (.A(\cla/_0666_ ),
    .B(\cla/_0667_ ),
    .C(\cla/_0521_ ),
    .Y(\cla/_0522_ ));
 sg13g2_nor3_1 \cla/_0900_  (.A(\cla/_0664_ ),
    .B(\cla/_0413_ ),
    .C(\cla/_0415_ ),
    .Y(\cla/_0523_ ));
 sg13g2_nor2_1 \cla/_0901_  (.A(\cla/_0522_ ),
    .B(\cla/_0523_ ),
    .Y(\cla/_0524_ ));
 sg13g2_o21ai_1 \cla/_0902_  (.B1(\cla/_0524_ ),
    .Y(\cla/_0525_ ),
    .A1(\cla/_0664_ ),
    .A2(\cla/_0427_ ));
 sg13g2_nor3_1 \cla/_0903_  (.A(\cla/_0515_ ),
    .B(\cla/_0520_ ),
    .C(\cla/_0525_ ),
    .Y(\cla/generate_adder_modules[17].fa_i.s ));
 sg13g2_inv_1 \cla/_0904_  (.Y(\cla/_0526_ ),
    .A(\cla/_0663_ ));
 sg13g2_a221oi_1 \cla/_0905_  (.B2(\cla/_0457_ ),
    .C1(\cla/_0424_ ),
    .B1(\cla/_0455_ ),
    .A1(\cla/_0436_ ),
    .Y(\cla/_0527_ ),
    .A2(\cla/_0440_ ));
 sg13g2_a21oi_1 \cla/_0906_  (.A1(\cla/_0357_ ),
    .A2(\cla/_0358_ ),
    .Y(\cla/_0528_ ),
    .B1(\cla/_0424_ ));
 sg13g2_or4_1 \cla/_0907_  (.A(\cla/_0513_ ),
    .B(\cla/_0505_ ),
    .C(\cla/_0527_ ),
    .D(\cla/_0528_ ),
    .X(\cla/_0529_ ));
 sg13g2_nand2_1 \cla/_0908_  (.Y(\cla/_0530_ ),
    .A(\cla/_0669_ ),
    .B(\rca.generate_adder_modules[15].fa.a ));
 sg13g2_and3_1 \cla/_0909_  (.X(\cla/_0531_ ),
    .A(\cla/_0674_ ),
    .B(net23),
    .C(\rca.generate_adder_modules[15].fa.a ));
 sg13g2_nand4_1 \cla/_0910_  (.B(\cla/_0433_ ),
    .C(\cla/_0360_ ),
    .A(\cla/_0414_ ),
    .Y(\cla/_0532_ ),
    .D(\cla/_0531_ ));
 sg13g2_and3_1 \cla/_0911_  (.X(\cla/_0533_ ),
    .A(\cla/_0674_ ),
    .B(net23),
    .C(\cla/_0669_ ));
 sg13g2_nand4_1 \cla/_0912_  (.B(\cla/_0433_ ),
    .C(\cla/_0360_ ),
    .A(\cla/_0414_ ),
    .Y(\cla/_0534_ ),
    .D(\cla/_0533_ ));
 sg13g2_nand3_1 \cla/_0913_  (.B(\cla/_0532_ ),
    .C(\cla/_0534_ ),
    .A(\cla/_0530_ ),
    .Y(\cla/_0535_ ));
 sg13g2_a21oi_1 \cla/_0914_  (.A1(\cla/_0667_ ),
    .A2(\cla/_0535_ ),
    .Y(\cla/_0536_ ),
    .B1(\cla/_0666_ ));
 sg13g2_nand2_1 \cla/_0915_  (.Y(\cla/_0537_ ),
    .A(\rca.generate_adder_modules[13].fa.b ),
    .B(\cla/_0672_ ));
 sg13g2_o21ai_1 \cla/_0916_  (.B1(\cla/_0513_ ),
    .Y(\cla/_0538_ ),
    .A1(\cla/_0505_ ),
    .A2(\cla/_0537_ ));
 sg13g2_nor2_1 \cla/_0917_  (.A(\cla/_0535_ ),
    .B(\cla/_0538_ ),
    .Y(\cla/_0539_ ));
 sg13g2_or4_1 \cla/_0918_  (.A(\cla/_0479_ ),
    .B(\cla/_0499_ ),
    .C(\cla/_0505_ ),
    .D(\cla/_0458_ ),
    .X(\cla/_0540_ ));
 sg13g2_a22oi_1 \cla/_0919_  (.Y(\cla/_0541_ ),
    .B1(\cla/_0539_ ),
    .B2(\cla/_0540_ ),
    .A2(\cla/_0536_ ),
    .A1(\cla/_0529_ ));
 sg13g2_nand2_1 \cla/_0920_  (.Y(\cla/_0542_ ),
    .A(\cla/_0521_ ),
    .B(\cla/_0362_ ));
 sg13g2_a21o_1 \cla/_0921_  (.A2(\cla/_0495_ ),
    .A1(\cla/_0494_ ),
    .B1(\cla/_0542_ ),
    .X(\cla/_0543_ ));
 sg13g2_a22oi_1 \cla/_0922_  (.Y(\cla/_0544_ ),
    .B1(\cla/_0491_ ),
    .B2(\cla/_0516_ ),
    .A2(\cla/_0683_ ),
    .A1(\cla/_0671_ ));
 sg13g2_nand2_1 \cla/_0923_  (.Y(\cla/_0545_ ),
    .A(\cla/_0543_ ),
    .B(\cla/_0544_ ));
 sg13g2_nor2_1 \cla/_0924_  (.A(\cla/_0541_ ),
    .B(\cla/_0545_ ),
    .Y(\cla/_0546_ ));
 sg13g2_nand3_1 \cla/_0925_  (.B(\cla/_0543_ ),
    .C(\cla/_0544_ ),
    .A(\cla/_0526_ ),
    .Y(\cla/_0547_ ));
 sg13g2_o21ai_1 \cla/_0926_  (.B1(\cla/_0662_ ),
    .Y(\cla/_0548_ ),
    .A1(\cla/_0541_ ),
    .A2(\cla/_0547_ ));
 sg13g2_o21ai_1 \cla/_0927_  (.B1(\cla/_0548_ ),
    .Y(\cla/_0549_ ),
    .A1(\cla/_0526_ ),
    .A2(\cla/_0546_ ));
 sg13g2_xnor2_1 \cla/_0928_  (.Y(\cla/generate_adder_modules[18].fa_i.s ),
    .A(\cla/_0661_ ),
    .B(\cla/_0549_ ));
 sg13g2_nand3b_1 \cla/_0929_  (.B(\cla/_0543_ ),
    .C(\cla/_0544_ ),
    .Y(\cla/_0550_ ),
    .A_N(\cla/_0662_ ));
 sg13g2_a21oi_1 \cla/_0930_  (.A1(\cla/_0547_ ),
    .A2(\cla/_0550_ ),
    .Y(\cla/_0551_ ),
    .B1(\cla/_0541_ ));
 sg13g2_or2_1 \cla/_0931_  (.X(\cla/_0552_ ),
    .B(\rca.generate_adder_modules[18].fa.a ),
    .A(\rca.generate_adder_modules[18].fa.b ));
 sg13g2_nand2b_1 \cla/_0932_  (.Y(\cla/_0553_ ),
    .B(\cla/_0552_ ),
    .A_N(\cla/_0428_ ));
 sg13g2_o21ai_1 \cla/_0933_  (.B1(\cla/_0392_ ),
    .Y(\cla/_0554_ ),
    .A1(\cla/_0551_ ),
    .A2(\cla/_0553_ ));
 sg13g2_xnor2_1 \cla/_0934_  (.Y(\cla/generate_adder_modules[19].fa_i.s ),
    .A(\cla/_0660_ ),
    .B(\cla/_0554_ ));
 sg13g2_nand2_1 \cla/_0935_  (.Y(\cla/_0555_ ),
    .A(\rca.generate_adder_modules[0].fa.b ),
    .B(\rca.generate_adder_modules[0].fa.a ));
 sg13g2_xor2_1 \cla/_0936_  (.B(\rca.generate_adder_modules[1].fa.a ),
    .A(\rca.generate_adder_modules[1].fa.b ),
    .X(\cla/_0556_ ));
 sg13g2_xnor2_1 \cla/_0937_  (.Y(\cla/generate_adder_modules[1].fa_i.s ),
    .A(\cla/_0555_ ),
    .B(\cla/_0556_ ));
 sg13g2_o21ai_1 \cla/_0938_  (.B1(\cla/_0385_ ),
    .Y(\cla/_0557_ ),
    .A1(\cla/_0665_ ),
    .A2(\cla/_0544_ ));
 sg13g2_nor3_1 \cla/_0939_  (.A(\cla/_0479_ ),
    .B(\cla/_0499_ ),
    .C(\cla/_0488_ ),
    .Y(\cla/_0558_ ));
 sg13g2_a21o_1 \cla/_0940_  (.A2(\cla/_0440_ ),
    .A1(\cla/_0436_ ),
    .B1(\cla/_0370_ ),
    .X(\cla/_0559_ ));
 sg13g2_nor2_1 \cla/_0941_  (.A(\cla/_0505_ ),
    .B(\cla/_0434_ ),
    .Y(\cla/_0560_ ));
 sg13g2_a21oi_1 \cla/_0942_  (.A1(\cla/_0558_ ),
    .A2(\cla/_0559_ ),
    .Y(\cla/_0561_ ),
    .B1(\cla/_0560_ ));
 sg13g2_nand2_1 \cla/_0943_  (.Y(\cla/_0562_ ),
    .A(\rca.generate_adder_modules[15].fa.a ),
    .B(\cla/_0389_ ));
 sg13g2_a21o_1 \cla/_0944_  (.A2(\cla/_0422_ ),
    .A1(\cla/_0418_ ),
    .B1(\cla/_0424_ ),
    .X(\cla/_0563_ ));
 sg13g2_and2_1 \cla/_0945_  (.A(\cla/_0359_ ),
    .B(\cla/_0362_ ),
    .X(\cla/_0564_ ));
 sg13g2_a221oi_1 \cla/_0946_  (.B2(\cla/_0564_ ),
    .C1(\cla/_0394_ ),
    .B1(\cla/_0563_ ),
    .A1(\cla/_0426_ ),
    .Y(\cla/_0565_ ),
    .A2(\cla/_0430_ ));
 sg13g2_o21ai_1 \cla/_0947_  (.B1(\cla/_0565_ ),
    .Y(\cla/_0566_ ),
    .A1(\cla/_0561_ ),
    .A2(\cla/_0562_ ));
 sg13g2_nand2_1 \cla/_0948_  (.Y(\cla/_0567_ ),
    .A(\cla/_0669_ ),
    .B(\cla/_0389_ ));
 sg13g2_nand2_1 \cla/_0949_  (.Y(\cla/_0568_ ),
    .A(\cla/_0389_ ),
    .B(\cla/_0390_ ));
 sg13g2_o21ai_1 \cla/_0950_  (.B1(\cla/_0568_ ),
    .Y(\cla/_0569_ ),
    .A1(\cla/_0561_ ),
    .A2(\cla/_0567_ ));
 sg13g2_nor3_1 \cla/_0951_  (.A(\cla/_0557_ ),
    .B(\cla/_0566_ ),
    .C(\cla/_0569_ ),
    .Y(\cla/_0570_ ));
 sg13g2_xnor2_1 \cla/_0952_  (.Y(\cla/generate_adder_modules[20].fa_i.s ),
    .A(\cla/_0346_ ),
    .B(\cla/_0570_ ));
 sg13g2_nor2_1 \cla/_0953_  (.A(\cla/_0407_ ),
    .B(\cla/_0404_ ),
    .Y(\cla/_0571_ ));
 sg13g2_o21ai_1 \cla/_0954_  (.B1(\cla/_0571_ ),
    .Y(\cla/_0572_ ),
    .A1(\cla/_0566_ ),
    .A2(\cla/_0569_ ));
 sg13g2_nor2_1 \cla/_0955_  (.A(\cla/_0444_ ),
    .B(\cla/_0404_ ),
    .Y(\cla/_0573_ ));
 sg13g2_o21ai_1 \cla/_0956_  (.B1(\cla/_0573_ ),
    .Y(\cla/_0574_ ),
    .A1(\cla/_0566_ ),
    .A2(\cla/_0569_ ));
 sg13g2_nand2_1 \cla/_0957_  (.Y(\cla/_0575_ ),
    .A(\cla/_0407_ ),
    .B(\cla/_0404_ ));
 sg13g2_nor4_1 \cla/_0958_  (.A(\cla/_0557_ ),
    .B(\cla/_0566_ ),
    .C(\cla/_0569_ ),
    .D(\cla/_0575_ ),
    .Y(\cla/_0576_ ));
 sg13g2_nand2_1 \cla/_0959_  (.Y(\cla/_0577_ ),
    .A(\cla/_0444_ ),
    .B(\cla/_0404_ ));
 sg13g2_nor4_1 \cla/_0960_  (.A(\cla/_0557_ ),
    .B(\cla/_0566_ ),
    .C(\cla/_0569_ ),
    .D(\cla/_0577_ ),
    .Y(\cla/_0578_ ));
 sg13g2_nor2_1 \cla/_0961_  (.A(\cla/_0576_ ),
    .B(\cla/_0578_ ),
    .Y(\cla/_0579_ ));
 sg13g2_o21ai_1 \cla/_0962_  (.B1(\cla/_0557_ ),
    .Y(\cla/_0580_ ),
    .A1(\cla/_0571_ ),
    .A2(\cla/_0573_ ));
 sg13g2_nand3_1 \cla/_0963_  (.B(\cla/_0345_ ),
    .C(\cla/_0349_ ),
    .A(\cla/_0344_ ),
    .Y(\cla/_0581_ ));
 sg13g2_nor2_1 \cla/_0964_  (.A(\cla/_0344_ ),
    .B(\cla/_0345_ ),
    .Y(\cla/_0582_ ));
 sg13g2_nand2_1 \cla/_0965_  (.Y(\cla/_0583_ ),
    .A(\cla/_0404_ ),
    .B(\cla/_0582_ ));
 sg13g2_and3_1 \cla/_0966_  (.X(\cla/_0584_ ),
    .A(\cla/_0580_ ),
    .B(\cla/_0581_ ),
    .C(\cla/_0583_ ));
 sg13g2_and4_1 \cla/_0967_  (.A(\cla/_0572_ ),
    .B(\cla/_0574_ ),
    .C(\cla/_0579_ ),
    .D(\cla/_0584_ ),
    .X(\cla/generate_adder_modules[21].fa_i.s ));
 sg13g2_and3_1 \cla/_0968_  (.X(\cla/_0585_ ),
    .A(\cla/_0530_ ),
    .B(\cla/_0532_ ),
    .C(\cla/_0534_ ));
 sg13g2_or4_1 \cla/_0969_  (.A(\cla/_0364_ ),
    .B(\cla/_0365_ ),
    .C(\cla/_0366_ ),
    .D(\cla/_0369_ ),
    .X(\cla/_0586_ ));
 sg13g2_nor3_1 \cla/_0970_  (.A(\cla/_0479_ ),
    .B(\cla/_0499_ ),
    .C(\cla/_0586_ ),
    .Y(\cla/_0587_ ));
 sg13g2_o21ai_1 \cla/_0971_  (.B1(\cla/_0506_ ),
    .Y(\cla/_0588_ ),
    .A1(\cla/_0424_ ),
    .A2(\cla/_0587_ ));
 sg13g2_nand2_1 \cla/_0972_  (.Y(\cla/_0589_ ),
    .A(\cla/_0359_ ),
    .B(\cla/_0668_ ));
 sg13g2_a21oi_1 \cla/_0973_  (.A1(\cla/_0585_ ),
    .A2(\cla/_0588_ ),
    .Y(\cla/_0590_ ),
    .B1(\cla/_0589_ ));
 sg13g2_o21ai_1 \cla/_0974_  (.B1(\cla/_0431_ ),
    .Y(\cla/_0591_ ),
    .A1(\cla/_0417_ ),
    .A2(\cla/_0494_ ));
 sg13g2_nor4_1 \cla/_0975_  (.A(\cla/_0442_ ),
    .B(\cla/_0557_ ),
    .C(\cla/_0590_ ),
    .D(\cla/_0591_ ),
    .Y(\cla/_0592_ ));
 sg13g2_nand2_1 \cla/_0976_  (.Y(\cla/_0593_ ),
    .A(\cla/_0345_ ),
    .B(\cla/_0394_ ));
 sg13g2_o21ai_1 \cla/_0977_  (.B1(\cla/_0344_ ),
    .Y(\cla/_0594_ ),
    .A1(\cla/_0345_ ),
    .A2(\cla/_0394_ ));
 sg13g2_a21oi_1 \cla/_0978_  (.A1(\cla/_0593_ ),
    .A2(\cla/_0594_ ),
    .Y(\cla/_0595_ ),
    .B1(\cla/_0397_ ));
 sg13g2_a21oi_1 \cla/_0979_  (.A1(\cla/_0347_ ),
    .A2(\cla/_0348_ ),
    .Y(\cla/_0596_ ),
    .B1(\cla/_0595_ ));
 sg13g2_o21ai_1 \cla/_0980_  (.B1(\cla/_0596_ ),
    .Y(\cla/_0597_ ),
    .A1(\cla/_0386_ ),
    .A2(\cla/_0592_ ));
 sg13g2_xnor2_1 \cla/_0981_  (.Y(\cla/generate_adder_modules[22].fa_i.s ),
    .A(\cla/_0343_ ),
    .B(\cla/_0597_ ));
 sg13g2_inv_1 \cla/_0982_  (.Y(\cla/_0598_ ),
    .A(\rca.generate_adder_modules[14].fa.b ));
 sg13g2_inv_1 \cla/_0983_  (.Y(\cla/_0599_ ),
    .A(\rca.generate_adder_modules[14].fa.a ));
 sg13g2_nor2_1 \cla/_0984_  (.A(\cla/_0598_ ),
    .B(\cla/_0599_ ),
    .Y(\cla/_0600_ ));
 sg13g2_nor2b_1 \cla/_0985_  (.A(\cla/_0354_ ),
    .B_N(\cla/_0409_ ),
    .Y(\cla/_0601_ ));
 sg13g2_nand2_1 \cla/_0986_  (.Y(\cla/_0602_ ),
    .A(\cla/_0678_ ),
    .B(\cla/_0601_ ));
 sg13g2_o21ai_1 \cla/_0987_  (.B1(\rca.generate_adder_modules[10].fa.b ),
    .Y(\cla/_0603_ ),
    .A1(\cla/_0678_ ),
    .A2(\cla/_0601_ ));
 sg13g2_a221oi_1 \cla/_0988_  (.B2(\cla/_0603_ ),
    .C1(\cla/_0499_ ),
    .B1(\cla/_0602_ ),
    .A1(\cla/_0598_ ),
    .Y(\cla/_0604_ ),
    .A2(\cla/_0599_ ));
 sg13g2_and2_1 \cla/_0989_  (.A(\cla/_0359_ ),
    .B(\cla/_0671_ ),
    .X(\cla/_0605_ ));
 sg13g2_o21ai_1 \cla/_0990_  (.B1(\cla/_0605_ ),
    .Y(\cla/_0606_ ),
    .A1(\cla/_0600_ ),
    .A2(\cla/_0604_ ));
 sg13g2_and4_1 \cla/_0991_  (.A(\cla/_0373_ ),
    .B(\cla/_0375_ ),
    .C(\cla/_0605_ ),
    .D(\cla/_0558_ ),
    .X(\cla/_0607_ ));
 sg13g2_nand4_1 \cla/_0992_  (.B(\cla/_0358_ ),
    .C(\cla/_0373_ ),
    .A(\cla/_0357_ ),
    .Y(\cla/_0608_ ),
    .D(\cla/_0379_ ));
 sg13g2_a21oi_1 \cla/_0993_  (.A1(\cla/_0537_ ),
    .A2(\cla/_0608_ ),
    .Y(\cla/_0609_ ),
    .B1(\cla/_0417_ ));
 sg13g2_a21oi_1 \cla/_0994_  (.A1(\cla/_0452_ ),
    .A2(\cla/_0441_ ),
    .Y(\cla/_0610_ ),
    .B1(\cla/_0363_ ));
 sg13g2_nand3_1 \cla/_0995_  (.B(\cla/_0418_ ),
    .C(\cla/_0422_ ),
    .A(\cla/_0506_ ),
    .Y(\cla/_0611_ ));
 sg13g2_a21oi_1 \cla/_0996_  (.A1(\cla/_0585_ ),
    .A2(\cla/_0611_ ),
    .Y(\cla/_0612_ ),
    .B1(\cla/_0589_ ));
 sg13g2_nor4_1 \cla/_0997_  (.A(\cla/_0607_ ),
    .B(\cla/_0609_ ),
    .C(\cla/_0610_ ),
    .D(\cla/_0612_ ),
    .Y(\cla/_0613_ ));
 sg13g2_a21oi_1 \cla/_0998_  (.A1(\cla/_0606_ ),
    .A2(\cla/_0613_ ),
    .Y(\cla/_0614_ ),
    .B1(\cla/_0351_ ));
 sg13g2_o21ai_1 \cla/_0999_  (.B1(\cla/_0405_ ),
    .Y(\cla/_0615_ ),
    .A1(\cla/_0402_ ),
    .A2(\cla/_0596_ ));
 sg13g2_inv_1 \cla/_1000_  (.Y(\cla/_0616_ ),
    .A(\cla/_0659_ ));
 sg13g2_nand3_1 \cla/_1001_  (.B(\cla/_0426_ ),
    .C(\cla/_0412_ ),
    .A(\cla/_0663_ ),
    .Y(\cla/_0617_ ));
 sg13g2_nand3_1 \cla/_1002_  (.B(\cla/_0426_ ),
    .C(\cla/_0412_ ),
    .A(\cla/_0662_ ),
    .Y(\cla/_0618_ ));
 sg13g2_a21oi_1 \cla/_1003_  (.A1(\cla/_0617_ ),
    .A2(\cla/_0618_ ),
    .Y(\cla/_0619_ ),
    .B1(\cla/_0415_ ));
 sg13g2_a221oi_1 \cla/_1004_  (.B2(\cla/_0564_ ),
    .C1(\cla/_0619_ ),
    .B1(\cla/_0587_ ),
    .A1(\cla/_0426_ ),
    .Y(\cla/_0620_ ),
    .A2(\cla/_0430_ ));
 sg13g2_nor3_1 \cla/_1005_  (.A(\cla/_0616_ ),
    .B(\cla/_0386_ ),
    .C(\cla/_0620_ ),
    .Y(\cla/_0621_ ));
 sg13g2_nand2_1 \cla/_1006_  (.Y(\cla/_0622_ ),
    .A(\cla/_0658_ ),
    .B(\cla/_0350_ ));
 sg13g2_nand2_1 \cla/_1007_  (.Y(\cla/_0623_ ),
    .A(\cla/_0658_ ),
    .B(\cla/_0659_ ));
 sg13g2_o21ai_1 \cla/_1008_  (.B1(\cla/_0623_ ),
    .Y(\cla/_0624_ ),
    .A1(\cla/_0620_ ),
    .A2(\cla/_0622_ ));
 sg13g2_nor4_1 \cla/_1009_  (.A(\cla/_0614_ ),
    .B(\cla/_0615_ ),
    .C(\cla/_0621_ ),
    .D(\cla/_0624_ ),
    .Y(\cla/_0625_ ));
 sg13g2_nor3_1 \cla/_1010_  (.A(\cla/_0660_ ),
    .B(\cla/_0351_ ),
    .C(\cla/_0405_ ),
    .Y(\cla/_0626_ ));
 sg13g2_nand3_1 \cla/_1011_  (.B(\cla/_0552_ ),
    .C(\cla/_0626_ ),
    .A(\cla/_0663_ ),
    .Y(\cla/_0627_ ));
 sg13g2_nand2b_1 \cla/_1012_  (.Y(\cla/_0628_ ),
    .B(\cla/_0626_ ),
    .A_N(\cla/_0392_ ));
 sg13g2_o21ai_1 \cla/_1013_  (.B1(\cla/_0628_ ),
    .Y(\cla/_0629_ ),
    .A1(\cla/_0546_ ),
    .A2(\cla/_0627_ ));
 sg13g2_a22oi_1 \cla/_1014_  (.Y(\cla/_0630_ ),
    .B1(\cla/_0344_ ),
    .B2(\cla/_0345_ ),
    .A2(\rca.generate_adder_modules[19].fa.a ),
    .A1(\rca.generate_adder_modules[19].fa.b ));
 sg13g2_nor3_1 \cla/_1015_  (.A(\cla/_0397_ ),
    .B(\cla/_0582_ ),
    .C(\cla/_0630_ ),
    .Y(\cla/_0631_ ));
 sg13g2_a21o_1 \cla/_1016_  (.A2(\cla/_0348_ ),
    .A1(\cla/_0347_ ),
    .B1(\cla/_0631_ ),
    .X(\cla/_0632_ ));
 sg13g2_o21ai_1 \cla/_1017_  (.B1(\cla/_0658_ ),
    .Y(\cla/_0633_ ),
    .A1(\cla/_0659_ ),
    .A2(\cla/_0632_ ));
 sg13g2_nand2_1 \cla/_1018_  (.Y(\cla/_0634_ ),
    .A(\cla/_0659_ ),
    .B(\cla/_0632_ ));
 sg13g2_a21oi_1 \cla/_1019_  (.A1(\cla/_0633_ ),
    .A2(\cla/_0634_ ),
    .Y(\cla/_0635_ ),
    .B1(\cla/_0405_ ));
 sg13g2_nand2_1 \cla/_1020_  (.Y(\cla/_0636_ ),
    .A(\cla/_0552_ ),
    .B(\cla/_0626_ ));
 sg13g2_nor2_1 \cla/_1021_  (.A(\cla/_0548_ ),
    .B(\cla/_0636_ ),
    .Y(\cla/_0637_ ));
 sg13g2_nor4_1 \cla/_1022_  (.A(\cla/_0625_ ),
    .B(\cla/_0629_ ),
    .C(\cla/_0635_ ),
    .D(\cla/_0637_ ),
    .Y(\cla/generate_adder_modules[23].fa_i.s ));
 sg13g2_xnor2_1 \cla/_1023_  (.Y(\cla/generate_adder_modules[2].fa_i.s ),
    .A(\cla/_0380_ ),
    .B(\cla/_0451_ ));
 sg13g2_inv_1 \cla/_1024_  (.Y(\cla/_0638_ ),
    .A(\rca.generate_adder_modules[2].fa.a ));
 sg13g2_o21ai_1 \cla/_1025_  (.B1(\cla/_0638_ ),
    .Y(\cla/_0639_ ),
    .A1(\cla/_0381_ ),
    .A2(\cla/_0382_ ));
 sg13g2_nor3_1 \cla/_1026_  (.A(\cla/_0638_ ),
    .B(\cla/_0381_ ),
    .C(\cla/_0382_ ),
    .Y(\cla/_0640_ ));
 sg13g2_a21o_1 \cla/_1027_  (.A2(\cla/_0639_ ),
    .A1(\rca.generate_adder_modules[2].fa.b ),
    .B1(\cla/_0640_ ),
    .X(\cla/_0641_ ));
 sg13g2_xnor2_1 \cla/_1028_  (.Y(\cla/generate_adder_modules[3].fa_i.s ),
    .A(\cla/_0377_ ),
    .B(\cla/_0641_ ));
 sg13g2_or2_1 \cla/_1029_  (.X(\cla/_0642_ ),
    .B(\rca.generate_adder_modules[3].fa.a ),
    .A(\rca.generate_adder_modules[3].fa.b ));
 sg13g2_and2_1 \cla/_1030_  (.A(\cla/_0642_ ),
    .B(\cla/_0641_ ),
    .X(\cla/_0643_ ));
 sg13g2_nor2_1 \cla/_1031_  (.A(\cla/_0375_ ),
    .B(\cla/_0643_ ),
    .Y(\cla/_0644_ ));
 sg13g2_xor2_1 \cla/_1032_  (.B(\cla/_0644_ ),
    .A(\cla/_0372_ ),
    .X(\cla/generate_adder_modules[4].fa_i.s ));
 sg13g2_inv_1 \cla/_1033_  (.Y(\cla/_0645_ ),
    .A(\cla/_0367_ ));
 sg13g2_o21ai_1 \cla/_1034_  (.B1(\cla/_0368_ ),
    .Y(\cla/_0646_ ),
    .A1(\cla/_0375_ ),
    .A2(\cla/_0643_ ));
 sg13g2_nor3_1 \cla/_1035_  (.A(\cla/_0368_ ),
    .B(\cla/_0375_ ),
    .C(\cla/_0643_ ),
    .Y(\cla/_0647_ ));
 sg13g2_a21oi_1 \cla/_1036_  (.A1(\cla/_0645_ ),
    .A2(\cla/_0646_ ),
    .Y(\cla/_0648_ ),
    .B1(\cla/_0647_ ));
 sg13g2_xnor2_1 \cla/_1037_  (.Y(\cla/generate_adder_modules[5].fa_i.s ),
    .A(\cla/_0366_ ),
    .B(\cla/_0648_ ));
 sg13g2_nand2b_1 \cla/_1038_  (.Y(\cla/_0649_ ),
    .B(\cla/_0438_ ),
    .A_N(\cla/_0375_ ));
 sg13g2_a221oi_1 \cla/_1039_  (.B2(\cla/_0641_ ),
    .C1(\cla/_0649_ ),
    .B1(\cla/_0642_ ),
    .A1(\cla/_0367_ ),
    .Y(\cla/_0650_ ),
    .A2(\cla/_0368_ ));
 sg13g2_nor2_1 \cla/_1040_  (.A(\rca.generate_adder_modules[5].fa.b ),
    .B(\rca.generate_adder_modules[5].fa.a ),
    .Y(\cla/_0651_ ));
 sg13g2_a21oi_1 \cla/_1041_  (.A1(\cla/_0438_ ),
    .A2(\cla/_0456_ ),
    .Y(\cla/_0652_ ),
    .B1(\cla/_0651_ ));
 sg13g2_nor2b_1 \cla/_1042_  (.A(\cla/_0650_ ),
    .B_N(\cla/_0652_ ),
    .Y(\cla/_0653_ ));
 sg13g2_xnor2_1 \cla/_1043_  (.Y(\cla/generate_adder_modules[6].fa_i.s ),
    .A(\cla/_0365_ ),
    .B(\cla/_0653_ ));
 sg13g2_a21oi_1 \cla/_1044_  (.A1(\rca.generate_adder_modules[6].fa.a ),
    .A2(\cla/_0653_ ),
    .Y(\cla/_0654_ ),
    .B1(\rca.generate_adder_modules[6].fa.b ));
 sg13g2_nor2_1 \cla/_1045_  (.A(\rca.generate_adder_modules[6].fa.a ),
    .B(\cla/_0653_ ),
    .Y(\cla/_0655_ ));
 sg13g2_nor2_1 \cla/_1046_  (.A(\cla/_0654_ ),
    .B(\cla/_0655_ ),
    .Y(\cla/_0656_ ));
 sg13g2_xnor2_1 \cla/_1047_  (.Y(\cla/generate_adder_modules[7].fa_i.s ),
    .A(\cla/_0364_ ),
    .B(\cla/_0656_ ));
 sg13g2_xnor2_1 \cla/_1048_  (.Y(\cla/generate_adder_modules[8].fa_i.s ),
    .A(\cla/_0356_ ),
    .B(\cla/_0459_ ));
 sg13g2_and2_1 \cla/_1049_  (.A(\cla/_0460_ ),
    .B(\cla/_0461_ ),
    .X(\cla/_0657_ ));
 sg13g2_xor2_1 \cla/_1050_  (.B(\cla/_0657_ ),
    .A(\cla/_0354_ ),
    .X(\cla/generate_adder_modules[9].fa_i.s ));
 sg13g2_buf_1 \cla/_1051_  (.A(\cla/generate_adder_modules[0].fa_i._2_ ),
    .X(\cla_z[0] ));
 sg13g2_buf_1 \cla/_1052_  (.A(\cla/generate_adder_modules[1].fa_i.s ),
    .X(\cla_z[1] ));
 sg13g2_buf_1 \cla/_1053_  (.A(\cla/generate_adder_modules[2].fa_i.s ),
    .X(\cla_z[2] ));
 sg13g2_buf_1 \cla/_1054_  (.A(\cla/generate_adder_modules[3].fa_i.s ),
    .X(\cla_z[3] ));
 sg13g2_buf_1 \cla/_1055_  (.A(\cla/generate_adder_modules[4].fa_i.s ),
    .X(\cla_z[4] ));
 sg13g2_buf_1 \cla/_1056_  (.A(\cla/generate_adder_modules[5].fa_i.s ),
    .X(\cla_z[5] ));
 sg13g2_buf_1 \cla/_1057_  (.A(\cla/generate_adder_modules[6].fa_i.s ),
    .X(\cla_z[6] ));
 sg13g2_buf_1 \cla/_1058_  (.A(\cla/generate_adder_modules[7].fa_i.s ),
    .X(\cla_z[7] ));
 sg13g2_buf_1 \cla/_1059_  (.A(\cla/generate_adder_modules[8].fa_i.s ),
    .X(\cla_z[8] ));
 sg13g2_buf_1 \cla/_1060_  (.A(\cla/generate_adder_modules[9].fa_i.s ),
    .X(\cla_z[9] ));
 sg13g2_buf_1 \cla/_1061_  (.A(\cla/generate_adder_modules[10].fa_i.s ),
    .X(\cla_z[10] ));
 sg13g2_buf_1 \cla/_1062_  (.A(\cla/generate_adder_modules[11].fa_i.s ),
    .X(\cla_z[11] ));
 sg13g2_buf_1 \cla/_1063_  (.A(\cla/generate_adder_modules[12].fa_i.s ),
    .X(\cla_z[12] ));
 sg13g2_buf_1 \cla/_1064_  (.A(\cla/generate_adder_modules[13].fa_i.s ),
    .X(\cla_z[13] ));
 sg13g2_buf_1 \cla/_1065_  (.A(\cla/generate_adder_modules[14].fa_i.s ),
    .X(\cla_z[14] ));
 sg13g2_buf_1 \cla/_1066_  (.A(\cla/generate_adder_modules[15].fa_i.s ),
    .X(\cla_z[15] ));
 sg13g2_buf_1 \cla/_1067_  (.A(\cla/generate_adder_modules[16].fa_i.s ),
    .X(\cla_z[16] ));
 sg13g2_buf_1 \cla/_1068_  (.A(\cla/generate_adder_modules[17].fa_i.s ),
    .X(\cla_z[17] ));
 sg13g2_buf_1 \cla/_1069_  (.A(\cla/generate_adder_modules[18].fa_i.s ),
    .X(\cla_z[18] ));
 sg13g2_buf_1 \cla/_1070_  (.A(\cla/generate_adder_modules[19].fa_i.s ),
    .X(\cla_z[19] ));
 sg13g2_buf_1 \cla/_1071_  (.A(\cla/generate_adder_modules[20].fa_i.s ),
    .X(\cla_z[20] ));
 sg13g2_buf_1 \cla/_1072_  (.A(\cla/generate_adder_modules[21].fa_i.s ),
    .X(\cla_z[21] ));
 sg13g2_buf_1 \cla/_1073_  (.A(\cla/generate_adder_modules[22].fa_i.s ),
    .X(\cla_z[22] ));
 sg13g2_buf_1 \cla/_1074_  (.A(\cla/generate_adder_modules[23].fa_i.s ),
    .X(\cla_z[23] ));
 sg13g2_buf_1 \cla/_1075_  (.A(\cla/_0341_ ),
    .X(net10));
 sg13g2_dfrbp_1 \io_sd.a_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net75),
    .D(_0006_),
    .Q_N(_0755_),
    .Q(\io_sd._052_[0] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[10]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net76),
    .D(_0007_),
    .Q_N(_0754_),
    .Q(\io_sd._052_[10] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[11]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net77),
    .D(_0008_),
    .Q_N(_0753_),
    .Q(\io_sd._052_[11] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[12]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net78),
    .D(_0009_),
    .Q_N(_0752_),
    .Q(\io_sd._052_[12] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[13]$_SDFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net79),
    .D(_0010_),
    .Q_N(_0751_),
    .Q(\io_sd._052_[13] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[14]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net80),
    .D(_0011_),
    .Q_N(_0750_),
    .Q(\io_sd._052_[14] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[15]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net81),
    .D(_0012_),
    .Q_N(_0749_),
    .Q(\io_sd._052_[15] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[16]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net82),
    .D(_0013_),
    .Q_N(_0748_),
    .Q(\io_sd._052_[16] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[17]$_SDFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net83),
    .D(_0014_),
    .Q_N(_0747_),
    .Q(\io_sd._052_[17] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[18]$_SDFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net84),
    .D(_0015_),
    .Q_N(_0746_),
    .Q(\io_sd._052_[18] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[19]$_SDFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net85),
    .D(_0016_),
    .Q_N(_0745_),
    .Q(\io_sd._052_[19] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net86),
    .D(_0017_),
    .Q_N(_0744_),
    .Q(\io_sd._052_[1] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[20]$_SDFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net87),
    .D(_0018_),
    .Q_N(_0743_),
    .Q(\io_sd._052_[20] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[21]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net88),
    .D(_0019_),
    .Q_N(_0742_),
    .Q(\io_sd._052_[21] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[22]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net89),
    .D(_0020_),
    .Q_N(_0741_),
    .Q(\io_sd._052_[22] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[23]$_SDFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net90),
    .D(_0021_),
    .Q_N(_0740_),
    .Q(\io_sd._052_[23] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(_0022_),
    .Q_N(_0739_),
    .Q(\io_sd._052_[2] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net92),
    .D(_0023_),
    .Q_N(_0738_),
    .Q(\io_sd._052_[3] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net93),
    .D(_0024_),
    .Q_N(_0737_),
    .Q(\io_sd._052_[4] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net94),
    .D(_0025_),
    .Q_N(_0736_),
    .Q(\io_sd._052_[5] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[6]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net95),
    .D(_0026_),
    .Q_N(_0735_),
    .Q(\io_sd._052_[6] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[7]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net96),
    .D(_0027_),
    .Q_N(_0734_),
    .Q(\io_sd._052_[7] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[8]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net97),
    .D(_0028_),
    .Q_N(_0733_),
    .Q(\io_sd._052_[8] ));
 sg13g2_dfrbp_1 \io_sd.a_reg[9]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net98),
    .D(_0029_),
    .Q_N(_0732_),
    .Q(\io_sd._052_[9] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[0]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net99),
    .D(_0030_),
    .Q_N(_0731_),
    .Q(\io_sd._053_[0] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[10]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net100),
    .D(_0031_),
    .Q_N(_0730_),
    .Q(\io_sd._053_[10] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[11]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net101),
    .D(_0032_),
    .Q_N(_0729_),
    .Q(\io_sd._053_[11] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[12]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net102),
    .D(_0033_),
    .Q_N(_0728_),
    .Q(\io_sd._053_[12] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[13]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(_0034_),
    .Q_N(_0727_),
    .Q(\io_sd._053_[13] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[14]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net104),
    .D(_0035_),
    .Q_N(_0726_),
    .Q(\io_sd._053_[14] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[15]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net105),
    .D(_0036_),
    .Q_N(_0725_),
    .Q(\io_sd._053_[15] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[16]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net106),
    .D(_0037_),
    .Q_N(_0724_),
    .Q(\io_sd._053_[16] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[17]$_SDFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net107),
    .D(_0038_),
    .Q_N(_0723_),
    .Q(\io_sd._053_[17] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[18]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net108),
    .D(_0039_),
    .Q_N(_0722_),
    .Q(\io_sd._053_[18] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[19]$_SDFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net109),
    .D(_0040_),
    .Q_N(_0721_),
    .Q(\io_sd._053_[19] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[1]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net110),
    .D(_0041_),
    .Q_N(_0720_),
    .Q(\io_sd._053_[1] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[20]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net111),
    .D(_0042_),
    .Q_N(_0719_),
    .Q(\io_sd._053_[20] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[21]$_SDFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net112),
    .D(_0043_),
    .Q_N(_0718_),
    .Q(\io_sd._053_[21] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[22]$_SDFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net113),
    .D(_0044_),
    .Q_N(_0717_),
    .Q(\io_sd._053_[22] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[23]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net114),
    .D(_0045_),
    .Q_N(_0716_),
    .Q(\io_sd._053_[23] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[2]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net115),
    .D(_0046_),
    .Q_N(_0715_),
    .Q(\io_sd._053_[2] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[3]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net116),
    .D(_0047_),
    .Q_N(_0714_),
    .Q(\io_sd._053_[3] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[4]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net117),
    .D(_0048_),
    .Q_N(_0713_),
    .Q(\io_sd._053_[4] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[5]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net118),
    .D(_0049_),
    .Q_N(_0712_),
    .Q(\io_sd._053_[5] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[6]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net119),
    .D(_0050_),
    .Q_N(_0711_),
    .Q(\io_sd._053_[6] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[7]$_SDFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net120),
    .D(_0051_),
    .Q_N(_0710_),
    .Q(\io_sd._053_[7] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[8]$_SDFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net121),
    .D(_0052_),
    .Q_N(_0709_),
    .Q(\io_sd._053_[8] ));
 sg13g2_dfrbp_1 \io_sd.b_reg[9]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net122),
    .D(_0053_),
    .Q_N(_0708_),
    .Q(\io_sd._053_[9] ));
 sg13g2_dfrbp_1 \io_sd.input_index[1]$_SDFFE_PN1P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net123),
    .D(_0054_),
    .Q_N(_0005_),
    .Q(\io_sd._210_[0] ));
 sg13g2_dfrbp_1 \io_sd.input_index[3]$_SDFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net124),
    .D(_0055_),
    .Q_N(_0707_),
    .Q(\io_sd.input_index[3] ));
 sg13g2_dfrbp_1 \io_sd.input_index[4]$_SDFFE_PN1P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net125),
    .D(_0056_),
    .Q_N(_0706_),
    .Q(\io_sd.input_index[4] ));
 sg13g2_dfrbp_1 \io_sd.input_index[5]$_SDFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net126),
    .D(_0057_),
    .Q_N(_0002_),
    .Q(\io_sd.input_index[5] ));
 sg13g2_dfrbp_1 \io_sd.output_index[1]$_SDFFE_PN1P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net127),
    .D(_0058_),
    .Q_N(_0004_),
    .Q(\io_sd._209_[0] ));
 sg13g2_dfrbp_1 \io_sd.output_index[3]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net128),
    .D(_0059_),
    .Q_N(_0705_),
    .Q(\io_sd.output_index[3] ));
 sg13g2_dfrbp_1 \io_sd.output_index[4]$_SDFFE_PN1P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net129),
    .D(_0060_),
    .Q_N(_0704_),
    .Q(\io_sd.output_index[4] ));
 sg13g2_dfrbp_1 \io_sd.output_index[5]$_SDFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net130),
    .D(_0061_),
    .Q_N(_0003_),
    .Q(\io_sd.output_index[5] ));
 sg13g2_dfrbp_1 \io_sd.outputs[0]$_SDFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net131),
    .D(_0062_),
    .Q_N(_0703_),
    .Q(net11));
 sg13g2_dfrbp_1 \io_sd.outputs[1]$_SDFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net132),
    .D(_0063_),
    .Q_N(_0702_),
    .Q(net12));
 sg13g2_dfrbp_1 \io_sd.outputs[2]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net133),
    .D(_0064_),
    .Q_N(_0701_),
    .Q(net13));
 sg13g2_dfrbp_1 \io_sd.outputs[3]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net134),
    .D(_0065_),
    .Q_N(_0700_),
    .Q(net14));
 sg13g2_dfrbp_1 \io_sd.outputs[4]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net135),
    .D(_0066_),
    .Q_N(_0699_),
    .Q(net15));
 sg13g2_dfrbp_1 \io_sd.outputs[5]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net136),
    .D(_0067_),
    .Q_N(_0698_),
    .Q(net16));
 sg13g2_dfrbp_1 \io_sd.outputs[6]$_SDFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net137),
    .D(_0068_),
    .Q_N(_0697_),
    .Q(net17));
 sg13g2_dfrbp_1 \io_sd.outputs[7]$_SDFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net138),
    .D(_0069_),
    .Q_N(_0756_),
    .Q(net18));
 sg13g2_dfrbp_1 \io_sd.state[0]$_DFF_P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net139),
    .D(_0000_),
    .Q_N(_0757_),
    .Q(\io_sd._068_ ));
 sg13g2_dfrbp_1 \io_sd.state[2]$_DFF_P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net140),
    .D(_0001_),
    .Q_N(_0696_),
    .Q(\io_sd._092_ ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout19 (.A(_0438_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0381_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0238_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0158_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(\cla/_0675_ ),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0499_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0369_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0341_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0285_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0284_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0122_),
    .X(net29));
 sg13g2_buf_1 fanout30 (.A(_0110_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0098_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0374_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0368_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0233_),
    .X(net34));
 sg13g2_buf_1 fanout35 (.A(_0218_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0150_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0143_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0097_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0093_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0084_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0082_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0077_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0308_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0236_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0217_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0171_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0140_),
    .X(net47));
 sg13g2_buf_4 fanout48 (.X(net48),
    .A(_0139_));
 sg13g2_buf_2 fanout49 (.A(_0131_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0130_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0126_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0125_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0112_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0100_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0099_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0096_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0090_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0074_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0071_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0072_),
    .X(net60));
 sg13g2_tielo _1503__61 (.L_LO(net61));
 sg13g2_tielo _1504__62 (.L_LO(net62));
 sg13g2_tielo _1505__63 (.L_LO(net63));
 sg13g2_tielo _1506__64 (.L_LO(net64));
 sg13g2_tielo _1507__65 (.L_LO(net65));
 sg13g2_tielo _1508__66 (.L_LO(net66));
 sg13g2_tielo _1511__67 (.L_LO(net67));
 sg13g2_tielo _1512__68 (.L_LO(net68));
 sg13g2_tielo _1513__69 (.L_LO(net69));
 sg13g2_tielo _1514__70 (.L_LO(net70));
 sg13g2_tielo _1515__71 (.L_LO(net71));
 sg13g2_tielo _1516__72 (.L_LO(net72));
 sg13g2_tiehi _1510__74 (.L_HI(net74));
 sg13g2_tiehi \io_sd.a_reg[0]$_SDFFE_PN0P__75  (.L_HI(net75));
 sg13g2_tiehi \io_sd.a_reg[10]$_SDFFE_PN0P__76  (.L_HI(net76));
 sg13g2_tiehi \io_sd.a_reg[11]$_SDFFE_PN0P__77  (.L_HI(net77));
 sg13g2_tiehi \io_sd.a_reg[12]$_SDFFE_PN0P__78  (.L_HI(net78));
 sg13g2_tiehi \io_sd.a_reg[13]$_SDFFE_PN0P__79  (.L_HI(net79));
 sg13g2_tiehi \io_sd.a_reg[14]$_SDFFE_PN0P__80  (.L_HI(net80));
 sg13g2_tiehi \io_sd.a_reg[15]$_SDFFE_PN0P__81  (.L_HI(net81));
 sg13g2_tiehi \io_sd.a_reg[16]$_SDFFE_PN0P__82  (.L_HI(net82));
 sg13g2_tiehi \io_sd.a_reg[17]$_SDFFE_PN0P__83  (.L_HI(net83));
 sg13g2_tiehi \io_sd.a_reg[18]$_SDFFE_PN0P__84  (.L_HI(net84));
 sg13g2_tiehi \io_sd.a_reg[19]$_SDFFE_PN0P__85  (.L_HI(net85));
 sg13g2_tiehi \io_sd.a_reg[1]$_SDFFE_PN0P__86  (.L_HI(net86));
 sg13g2_tiehi \io_sd.a_reg[20]$_SDFFE_PN0P__87  (.L_HI(net87));
 sg13g2_tiehi \io_sd.a_reg[21]$_SDFFE_PN0P__88  (.L_HI(net88));
 sg13g2_tiehi \io_sd.a_reg[22]$_SDFFE_PN0P__89  (.L_HI(net89));
 sg13g2_tiehi \io_sd.a_reg[23]$_SDFFE_PN0P__90  (.L_HI(net90));
 sg13g2_tiehi \io_sd.a_reg[2]$_SDFFE_PN0P__91  (.L_HI(net91));
 sg13g2_tiehi \io_sd.a_reg[3]$_SDFFE_PN0P__92  (.L_HI(net92));
 sg13g2_tiehi \io_sd.a_reg[4]$_SDFFE_PN0P__93  (.L_HI(net93));
 sg13g2_tiehi \io_sd.a_reg[5]$_SDFFE_PN0P__94  (.L_HI(net94));
 sg13g2_tiehi \io_sd.a_reg[6]$_SDFFE_PN0P__95  (.L_HI(net95));
 sg13g2_tiehi \io_sd.a_reg[7]$_SDFFE_PN0P__96  (.L_HI(net96));
 sg13g2_tiehi \io_sd.a_reg[8]$_SDFFE_PN0P__97  (.L_HI(net97));
 sg13g2_tiehi \io_sd.a_reg[9]$_SDFFE_PN0P__98  (.L_HI(net98));
 sg13g2_tiehi \io_sd.b_reg[0]$_SDFFE_PN0P__99  (.L_HI(net99));
 sg13g2_tiehi \io_sd.b_reg[10]$_SDFFE_PN0P__100  (.L_HI(net100));
 sg13g2_tiehi \io_sd.b_reg[11]$_SDFFE_PN0P__101  (.L_HI(net101));
 sg13g2_tiehi \io_sd.b_reg[12]$_SDFFE_PN0P__102  (.L_HI(net102));
 sg13g2_tiehi \io_sd.b_reg[13]$_SDFFE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \io_sd.b_reg[14]$_SDFFE_PN0P__104  (.L_HI(net104));
 sg13g2_tiehi \io_sd.b_reg[15]$_SDFFE_PN0P__105  (.L_HI(net105));
 sg13g2_tiehi \io_sd.b_reg[16]$_SDFFE_PN0P__106  (.L_HI(net106));
 sg13g2_tiehi \io_sd.b_reg[17]$_SDFFE_PN0P__107  (.L_HI(net107));
 sg13g2_tiehi \io_sd.b_reg[18]$_SDFFE_PN0P__108  (.L_HI(net108));
 sg13g2_tiehi \io_sd.b_reg[19]$_SDFFE_PN0P__109  (.L_HI(net109));
 sg13g2_tiehi \io_sd.b_reg[1]$_SDFFE_PN0P__110  (.L_HI(net110));
 sg13g2_tiehi \io_sd.b_reg[20]$_SDFFE_PN0P__111  (.L_HI(net111));
 sg13g2_tiehi \io_sd.b_reg[21]$_SDFFE_PN0P__112  (.L_HI(net112));
 sg13g2_tiehi \io_sd.b_reg[22]$_SDFFE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \io_sd.b_reg[23]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \io_sd.b_reg[2]$_SDFFE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \io_sd.b_reg[3]$_SDFFE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \io_sd.b_reg[4]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \io_sd.b_reg[5]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \io_sd.b_reg[6]$_SDFFE_PN0P__119  (.L_HI(net119));
 sg13g2_tiehi \io_sd.b_reg[7]$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi \io_sd.b_reg[8]$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \io_sd.b_reg[9]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \io_sd.input_index[1]$_SDFFE_PN1P__123  (.L_HI(net123));
 sg13g2_tiehi \io_sd.input_index[3]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \io_sd.input_index[4]$_SDFFE_PN1P__125  (.L_HI(net125));
 sg13g2_tiehi \io_sd.input_index[5]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_tiehi \io_sd.output_index[1]$_SDFFE_PN1P__127  (.L_HI(net127));
 sg13g2_tiehi \io_sd.output_index[3]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \io_sd.output_index[4]$_SDFFE_PN1P__129  (.L_HI(net129));
 sg13g2_tiehi \io_sd.output_index[5]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \io_sd.outputs[0]$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_tiehi \io_sd.outputs[1]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_tiehi \io_sd.outputs[2]$_SDFFE_PN0P__133  (.L_HI(net133));
 sg13g2_tiehi \io_sd.outputs[3]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_tiehi \io_sd.outputs[4]$_SDFFE_PN0P__135  (.L_HI(net135));
 sg13g2_tiehi \io_sd.outputs[5]$_SDFFE_PN0P__136  (.L_HI(net136));
 sg13g2_tiehi \io_sd.outputs[6]$_SDFFE_PN0P__137  (.L_HI(net137));
 sg13g2_tiehi \io_sd.outputs[7]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \io_sd.state[0]$_DFF_P__139  (.L_HI(net139));
 sg13g2_tiehi \io_sd.state[2]$_DFF_P__140  (.L_HI(net140));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_155 ();
 sg13g2_decap_8 FILLER_0_162 ();
 sg13g2_decap_8 FILLER_0_169 ();
 sg13g2_decap_8 FILLER_0_176 ();
 sg13g2_decap_8 FILLER_0_183 ();
 sg13g2_decap_8 FILLER_0_190 ();
 sg13g2_decap_8 FILLER_0_197 ();
 sg13g2_decap_8 FILLER_0_204 ();
 sg13g2_decap_8 FILLER_0_211 ();
 sg13g2_decap_8 FILLER_0_218 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_253 ();
 sg13g2_decap_8 FILLER_0_260 ();
 sg13g2_decap_4 FILLER_0_267 ();
 sg13g2_fill_2 FILLER_0_271 ();
 sg13g2_fill_1 FILLER_0_277 ();
 sg13g2_fill_1 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_4 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_4 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_fill_2 FILLER_1_112 ();
 sg13g2_fill_1 FILLER_1_114 ();
 sg13g2_decap_8 FILLER_1_124 ();
 sg13g2_decap_8 FILLER_1_151 ();
 sg13g2_fill_1 FILLER_1_158 ();
 sg13g2_decap_4 FILLER_1_175 ();
 sg13g2_fill_2 FILLER_1_179 ();
 sg13g2_fill_1 FILLER_1_185 ();
 sg13g2_decap_4 FILLER_1_194 ();
 sg13g2_fill_1 FILLER_1_203 ();
 sg13g2_fill_1 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_214 ();
 sg13g2_decap_8 FILLER_1_219 ();
 sg13g2_decap_8 FILLER_1_226 ();
 sg13g2_decap_8 FILLER_1_233 ();
 sg13g2_decap_8 FILLER_1_240 ();
 sg13g2_decap_4 FILLER_1_247 ();
 sg13g2_fill_1 FILLER_1_251 ();
 sg13g2_decap_4 FILLER_1_256 ();
 sg13g2_fill_2 FILLER_1_260 ();
 sg13g2_decap_4 FILLER_1_283 ();
 sg13g2_fill_2 FILLER_1_287 ();
 sg13g2_fill_2 FILLER_1_293 ();
 sg13g2_fill_1 FILLER_1_295 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_4 FILLER_1_315 ();
 sg13g2_fill_2 FILLER_1_335 ();
 sg13g2_fill_1 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_346 ();
 sg13g2_decap_8 FILLER_1_353 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_1_409 ();
 sg13g2_decap_8 FILLER_1_416 ();
 sg13g2_decap_8 FILLER_1_423 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_fill_2 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_128 ();
 sg13g2_decap_4 FILLER_2_135 ();
 sg13g2_decap_4 FILLER_2_143 ();
 sg13g2_decap_4 FILLER_2_151 ();
 sg13g2_fill_1 FILLER_2_155 ();
 sg13g2_decap_4 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_185 ();
 sg13g2_fill_2 FILLER_2_193 ();
 sg13g2_fill_1 FILLER_2_195 ();
 sg13g2_decap_8 FILLER_2_206 ();
 sg13g2_decap_8 FILLER_2_213 ();
 sg13g2_decap_4 FILLER_2_220 ();
 sg13g2_fill_1 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_240 ();
 sg13g2_decap_8 FILLER_2_261 ();
 sg13g2_decap_4 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_276 ();
 sg13g2_fill_1 FILLER_2_283 ();
 sg13g2_decap_8 FILLER_2_304 ();
 sg13g2_decap_4 FILLER_2_311 ();
 sg13g2_fill_2 FILLER_2_320 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_fill_1 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_344 ();
 sg13g2_decap_8 FILLER_2_351 ();
 sg13g2_decap_8 FILLER_2_358 ();
 sg13g2_decap_8 FILLER_2_365 ();
 sg13g2_decap_8 FILLER_2_372 ();
 sg13g2_decap_8 FILLER_2_379 ();
 sg13g2_decap_8 FILLER_2_386 ();
 sg13g2_decap_8 FILLER_2_393 ();
 sg13g2_decap_8 FILLER_2_400 ();
 sg13g2_decap_8 FILLER_2_407 ();
 sg13g2_decap_8 FILLER_2_414 ();
 sg13g2_decap_8 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_428 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_fill_2 FILLER_3_84 ();
 sg13g2_fill_1 FILLER_3_86 ();
 sg13g2_fill_1 FILLER_3_111 ();
 sg13g2_decap_4 FILLER_3_124 ();
 sg13g2_fill_2 FILLER_3_128 ();
 sg13g2_decap_4 FILLER_3_134 ();
 sg13g2_decap_8 FILLER_3_143 ();
 sg13g2_decap_4 FILLER_3_150 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_181 ();
 sg13g2_decap_4 FILLER_3_192 ();
 sg13g2_fill_1 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_202 ();
 sg13g2_fill_2 FILLER_3_209 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_fill_2 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_258 ();
 sg13g2_decap_4 FILLER_3_265 ();
 sg13g2_fill_2 FILLER_3_269 ();
 sg13g2_decap_8 FILLER_3_289 ();
 sg13g2_decap_8 FILLER_3_296 ();
 sg13g2_fill_1 FILLER_3_303 ();
 sg13g2_fill_1 FILLER_3_344 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_4 FILLER_3_361 ();
 sg13g2_fill_2 FILLER_3_365 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_4 FILLER_3_392 ();
 sg13g2_fill_2 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_4 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_94 ();
 sg13g2_fill_2 FILLER_4_101 ();
 sg13g2_fill_1 FILLER_4_103 ();
 sg13g2_fill_1 FILLER_4_108 ();
 sg13g2_decap_4 FILLER_4_113 ();
 sg13g2_fill_1 FILLER_4_122 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_decap_8 FILLER_4_141 ();
 sg13g2_decap_8 FILLER_4_148 ();
 sg13g2_fill_2 FILLER_4_163 ();
 sg13g2_decap_4 FILLER_4_184 ();
 sg13g2_fill_1 FILLER_4_188 ();
 sg13g2_decap_8 FILLER_4_198 ();
 sg13g2_fill_2 FILLER_4_205 ();
 sg13g2_fill_2 FILLER_4_220 ();
 sg13g2_fill_1 FILLER_4_222 ();
 sg13g2_fill_2 FILLER_4_229 ();
 sg13g2_decap_4 FILLER_4_240 ();
 sg13g2_fill_2 FILLER_4_244 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_fill_2 FILLER_4_298 ();
 sg13g2_fill_1 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_313 ();
 sg13g2_decap_8 FILLER_4_320 ();
 sg13g2_decap_4 FILLER_4_327 ();
 sg13g2_fill_1 FILLER_4_342 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_decap_4 FILLER_4_355 ();
 sg13g2_fill_1 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_decap_4 FILLER_5_23 ();
 sg13g2_decap_8 FILLER_5_48 ();
 sg13g2_decap_8 FILLER_5_55 ();
 sg13g2_fill_2 FILLER_5_62 ();
 sg13g2_fill_1 FILLER_5_64 ();
 sg13g2_decap_8 FILLER_5_79 ();
 sg13g2_decap_4 FILLER_5_117 ();
 sg13g2_fill_1 FILLER_5_121 ();
 sg13g2_decap_4 FILLER_5_149 ();
 sg13g2_fill_1 FILLER_5_153 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_4 FILLER_5_168 ();
 sg13g2_fill_1 FILLER_5_172 ();
 sg13g2_decap_4 FILLER_5_188 ();
 sg13g2_fill_2 FILLER_5_192 ();
 sg13g2_decap_8 FILLER_5_205 ();
 sg13g2_decap_8 FILLER_5_212 ();
 sg13g2_decap_4 FILLER_5_219 ();
 sg13g2_fill_1 FILLER_5_232 ();
 sg13g2_fill_1 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_257 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_decap_4 FILLER_5_271 ();
 sg13g2_fill_2 FILLER_5_275 ();
 sg13g2_fill_2 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_4 FILLER_5_299 ();
 sg13g2_fill_1 FILLER_5_303 ();
 sg13g2_decap_8 FILLER_5_313 ();
 sg13g2_fill_1 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_fill_1 FILLER_5_332 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_decap_8 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_fill_2 FILLER_5_367 ();
 sg13g2_fill_1 FILLER_5_369 ();
 sg13g2_fill_2 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_fill_2 FILLER_5_413 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_9 ();
 sg13g2_fill_2 FILLER_6_19 ();
 sg13g2_fill_1 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_38 ();
 sg13g2_decap_8 FILLER_6_45 ();
 sg13g2_decap_4 FILLER_6_52 ();
 sg13g2_fill_2 FILLER_6_68 ();
 sg13g2_decap_8 FILLER_6_79 ();
 sg13g2_decap_8 FILLER_6_86 ();
 sg13g2_decap_8 FILLER_6_93 ();
 sg13g2_fill_2 FILLER_6_100 ();
 sg13g2_fill_1 FILLER_6_102 ();
 sg13g2_fill_2 FILLER_6_112 ();
 sg13g2_fill_2 FILLER_6_119 ();
 sg13g2_fill_1 FILLER_6_121 ();
 sg13g2_decap_8 FILLER_6_127 ();
 sg13g2_decap_4 FILLER_6_134 ();
 sg13g2_fill_2 FILLER_6_138 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_4 FILLER_6_158 ();
 sg13g2_fill_2 FILLER_6_162 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_fill_2 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_fill_1 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_fill_1 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_4 FILLER_6_252 ();
 sg13g2_fill_2 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_264 ();
 sg13g2_fill_1 FILLER_6_271 ();
 sg13g2_fill_1 FILLER_6_289 ();
 sg13g2_decap_4 FILLER_6_295 ();
 sg13g2_fill_1 FILLER_6_299 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_fill_2 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_fill_1 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_11 ();
 sg13g2_decap_8 FILLER_7_23 ();
 sg13g2_decap_4 FILLER_7_30 ();
 sg13g2_fill_1 FILLER_7_50 ();
 sg13g2_fill_2 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_58 ();
 sg13g2_decap_8 FILLER_7_64 ();
 sg13g2_decap_8 FILLER_7_71 ();
 sg13g2_fill_2 FILLER_7_78 ();
 sg13g2_decap_8 FILLER_7_87 ();
 sg13g2_decap_8 FILLER_7_94 ();
 sg13g2_decap_4 FILLER_7_101 ();
 sg13g2_decap_8 FILLER_7_110 ();
 sg13g2_decap_8 FILLER_7_117 ();
 sg13g2_decap_8 FILLER_7_124 ();
 sg13g2_decap_8 FILLER_7_131 ();
 sg13g2_decap_8 FILLER_7_138 ();
 sg13g2_fill_2 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_152 ();
 sg13g2_decap_4 FILLER_7_161 ();
 sg13g2_fill_1 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_184 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_fill_1 FILLER_7_203 ();
 sg13g2_decap_4 FILLER_7_215 ();
 sg13g2_fill_1 FILLER_7_232 ();
 sg13g2_decap_4 FILLER_7_245 ();
 sg13g2_fill_1 FILLER_7_249 ();
 sg13g2_decap_4 FILLER_7_270 ();
 sg13g2_fill_1 FILLER_7_274 ();
 sg13g2_decap_8 FILLER_7_283 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_fill_1 FILLER_7_318 ();
 sg13g2_fill_1 FILLER_7_327 ();
 sg13g2_decap_4 FILLER_7_349 ();
 sg13g2_fill_1 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_1 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_7_417 ();
 sg13g2_decap_4 FILLER_7_424 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_7 ();
 sg13g2_fill_2 FILLER_8_11 ();
 sg13g2_fill_2 FILLER_8_24 ();
 sg13g2_decap_8 FILLER_8_59 ();
 sg13g2_decap_4 FILLER_8_74 ();
 sg13g2_fill_1 FILLER_8_78 ();
 sg13g2_fill_1 FILLER_8_87 ();
 sg13g2_decap_4 FILLER_8_101 ();
 sg13g2_decap_8 FILLER_8_114 ();
 sg13g2_decap_8 FILLER_8_121 ();
 sg13g2_decap_8 FILLER_8_128 ();
 sg13g2_decap_8 FILLER_8_135 ();
 sg13g2_fill_2 FILLER_8_142 ();
 sg13g2_fill_1 FILLER_8_144 ();
 sg13g2_fill_1 FILLER_8_152 ();
 sg13g2_fill_1 FILLER_8_158 ();
 sg13g2_fill_2 FILLER_8_163 ();
 sg13g2_fill_1 FILLER_8_169 ();
 sg13g2_decap_4 FILLER_8_182 ();
 sg13g2_fill_1 FILLER_8_186 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_fill_2 FILLER_8_199 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_decap_4 FILLER_8_214 ();
 sg13g2_fill_1 FILLER_8_223 ();
 sg13g2_fill_2 FILLER_8_236 ();
 sg13g2_fill_1 FILLER_8_238 ();
 sg13g2_decap_4 FILLER_8_252 ();
 sg13g2_fill_1 FILLER_8_256 ();
 sg13g2_fill_2 FILLER_8_263 ();
 sg13g2_fill_1 FILLER_8_265 ();
 sg13g2_decap_4 FILLER_8_274 ();
 sg13g2_fill_2 FILLER_8_278 ();
 sg13g2_fill_1 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_4 FILLER_8_312 ();
 sg13g2_fill_1 FILLER_8_316 ();
 sg13g2_decap_4 FILLER_8_325 ();
 sg13g2_fill_2 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_1 FILLER_8_375 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_18 ();
 sg13g2_fill_2 FILLER_9_24 ();
 sg13g2_fill_1 FILLER_9_30 ();
 sg13g2_fill_2 FILLER_9_40 ();
 sg13g2_fill_1 FILLER_9_42 ();
 sg13g2_fill_2 FILLER_9_48 ();
 sg13g2_decap_8 FILLER_9_58 ();
 sg13g2_decap_8 FILLER_9_65 ();
 sg13g2_decap_8 FILLER_9_72 ();
 sg13g2_fill_1 FILLER_9_79 ();
 sg13g2_fill_1 FILLER_9_85 ();
 sg13g2_fill_2 FILLER_9_91 ();
 sg13g2_fill_2 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_decap_4 FILLER_9_126 ();
 sg13g2_decap_4 FILLER_9_135 ();
 sg13g2_decap_4 FILLER_9_144 ();
 sg13g2_fill_2 FILLER_9_148 ();
 sg13g2_decap_4 FILLER_9_158 ();
 sg13g2_fill_1 FILLER_9_162 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_fill_1 FILLER_9_203 ();
 sg13g2_fill_2 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_215 ();
 sg13g2_decap_8 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_decap_4 FILLER_9_253 ();
 sg13g2_fill_2 FILLER_9_257 ();
 sg13g2_decap_8 FILLER_9_264 ();
 sg13g2_decap_8 FILLER_9_275 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_304 ();
 sg13g2_decap_4 FILLER_9_311 ();
 sg13g2_fill_2 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_fill_2 FILLER_9_361 ();
 sg13g2_fill_1 FILLER_9_363 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_decap_4 FILLER_9_380 ();
 sg13g2_fill_1 FILLER_9_388 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_decap_8 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_9_415 ();
 sg13g2_decap_8 FILLER_9_422 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_fill_2 FILLER_10_21 ();
 sg13g2_decap_4 FILLER_10_37 ();
 sg13g2_decap_4 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_50 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_fill_2 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_72 ();
 sg13g2_decap_4 FILLER_10_87 ();
 sg13g2_decap_8 FILLER_10_101 ();
 sg13g2_fill_1 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_fill_1 FILLER_10_154 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_decap_4 FILLER_10_172 ();
 sg13g2_fill_2 FILLER_10_176 ();
 sg13g2_decap_4 FILLER_10_186 ();
 sg13g2_fill_1 FILLER_10_190 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_fill_1 FILLER_10_219 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_4 FILLER_10_252 ();
 sg13g2_fill_2 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_267 ();
 sg13g2_fill_2 FILLER_10_274 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_307 ();
 sg13g2_decap_4 FILLER_10_314 ();
 sg13g2_fill_2 FILLER_10_318 ();
 sg13g2_decap_4 FILLER_10_324 ();
 sg13g2_fill_1 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_fill_2 FILLER_10_348 ();
 sg13g2_fill_1 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_fill_2 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_10_384 ();
 sg13g2_fill_1 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_404 ();
 sg13g2_decap_8 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_4 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_32 ();
 sg13g2_decap_4 FILLER_11_40 ();
 sg13g2_fill_2 FILLER_11_44 ();
 sg13g2_fill_1 FILLER_11_50 ();
 sg13g2_decap_8 FILLER_11_61 ();
 sg13g2_decap_8 FILLER_11_68 ();
 sg13g2_decap_4 FILLER_11_75 ();
 sg13g2_fill_1 FILLER_11_104 ();
 sg13g2_fill_2 FILLER_11_113 ();
 sg13g2_fill_1 FILLER_11_115 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_128 ();
 sg13g2_decap_8 FILLER_11_139 ();
 sg13g2_decap_8 FILLER_11_146 ();
 sg13g2_decap_8 FILLER_11_153 ();
 sg13g2_decap_8 FILLER_11_160 ();
 sg13g2_decap_8 FILLER_11_167 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_fill_1 FILLER_11_181 ();
 sg13g2_decap_4 FILLER_11_200 ();
 sg13g2_fill_1 FILLER_11_204 ();
 sg13g2_fill_2 FILLER_11_226 ();
 sg13g2_fill_1 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_238 ();
 sg13g2_fill_2 FILLER_11_268 ();
 sg13g2_fill_1 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_279 ();
 sg13g2_decap_8 FILLER_11_286 ();
 sg13g2_decap_4 FILLER_11_293 ();
 sg13g2_fill_1 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_4 FILLER_11_315 ();
 sg13g2_fill_1 FILLER_11_319 ();
 sg13g2_fill_2 FILLER_11_324 ();
 sg13g2_fill_2 FILLER_11_331 ();
 sg13g2_decap_8 FILLER_11_338 ();
 sg13g2_fill_2 FILLER_11_345 ();
 sg13g2_fill_2 FILLER_11_351 ();
 sg13g2_fill_1 FILLER_11_353 ();
 sg13g2_fill_1 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_4 FILLER_11_391 ();
 sg13g2_fill_2 FILLER_11_395 ();
 sg13g2_fill_2 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_fill_2 FILLER_12_31 ();
 sg13g2_decap_8 FILLER_12_41 ();
 sg13g2_decap_4 FILLER_12_48 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_4 FILLER_12_63 ();
 sg13g2_fill_2 FILLER_12_67 ();
 sg13g2_fill_2 FILLER_12_78 ();
 sg13g2_fill_1 FILLER_12_80 ();
 sg13g2_fill_2 FILLER_12_85 ();
 sg13g2_fill_1 FILLER_12_87 ();
 sg13g2_decap_8 FILLER_12_108 ();
 sg13g2_decap_8 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_decap_8 FILLER_12_134 ();
 sg13g2_decap_8 FILLER_12_141 ();
 sg13g2_decap_4 FILLER_12_148 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_fill_2 FILLER_12_165 ();
 sg13g2_decap_4 FILLER_12_172 ();
 sg13g2_fill_2 FILLER_12_176 ();
 sg13g2_decap_8 FILLER_12_194 ();
 sg13g2_decap_8 FILLER_12_201 ();
 sg13g2_fill_1 FILLER_12_208 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_fill_2 FILLER_12_234 ();
 sg13g2_decap_8 FILLER_12_241 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_4 FILLER_12_266 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_fill_2 FILLER_12_289 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_4 FILLER_12_312 ();
 sg13g2_fill_1 FILLER_12_316 ();
 sg13g2_decap_8 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_341 ();
 sg13g2_decap_4 FILLER_12_348 ();
 sg13g2_fill_1 FILLER_12_352 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_4 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_4 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_410 ();
 sg13g2_decap_8 FILLER_12_415 ();
 sg13g2_decap_8 FILLER_12_422 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_14 ();
 sg13g2_fill_1 FILLER_13_16 ();
 sg13g2_fill_2 FILLER_13_27 ();
 sg13g2_fill_1 FILLER_13_42 ();
 sg13g2_fill_1 FILLER_13_48 ();
 sg13g2_decap_8 FILLER_13_54 ();
 sg13g2_decap_4 FILLER_13_61 ();
 sg13g2_fill_2 FILLER_13_65 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_decap_4 FILLER_13_78 ();
 sg13g2_decap_4 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_101 ();
 sg13g2_decap_4 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_125 ();
 sg13g2_fill_2 FILLER_13_132 ();
 sg13g2_decap_8 FILLER_13_144 ();
 sg13g2_decap_4 FILLER_13_151 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_decap_8 FILLER_13_167 ();
 sg13g2_decap_8 FILLER_13_187 ();
 sg13g2_fill_2 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_fill_2 FILLER_13_201 ();
 sg13g2_decap_8 FILLER_13_208 ();
 sg13g2_fill_1 FILLER_13_215 ();
 sg13g2_decap_4 FILLER_13_229 ();
 sg13g2_fill_2 FILLER_13_233 ();
 sg13g2_decap_8 FILLER_13_240 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_decap_8 FILLER_13_254 ();
 sg13g2_decap_8 FILLER_13_261 ();
 sg13g2_decap_4 FILLER_13_268 ();
 sg13g2_fill_1 FILLER_13_272 ();
 sg13g2_decap_4 FILLER_13_281 ();
 sg13g2_decap_8 FILLER_13_289 ();
 sg13g2_fill_2 FILLER_13_296 ();
 sg13g2_fill_1 FILLER_13_307 ();
 sg13g2_decap_8 FILLER_13_314 ();
 sg13g2_fill_1 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_4 FILLER_13_346 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_fill_1 FILLER_13_386 ();
 sg13g2_fill_1 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_18 ();
 sg13g2_decap_4 FILLER_14_25 ();
 sg13g2_fill_1 FILLER_14_29 ();
 sg13g2_decap_8 FILLER_14_40 ();
 sg13g2_decap_8 FILLER_14_47 ();
 sg13g2_decap_8 FILLER_14_54 ();
 sg13g2_fill_2 FILLER_14_61 ();
 sg13g2_decap_8 FILLER_14_67 ();
 sg13g2_decap_4 FILLER_14_74 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_fill_2 FILLER_14_96 ();
 sg13g2_fill_1 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_103 ();
 sg13g2_fill_2 FILLER_14_110 ();
 sg13g2_decap_8 FILLER_14_121 ();
 sg13g2_decap_8 FILLER_14_128 ();
 sg13g2_fill_2 FILLER_14_135 ();
 sg13g2_decap_8 FILLER_14_141 ();
 sg13g2_decap_8 FILLER_14_148 ();
 sg13g2_decap_4 FILLER_14_155 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_decap_4 FILLER_14_164 ();
 sg13g2_decap_8 FILLER_14_177 ();
 sg13g2_decap_8 FILLER_14_184 ();
 sg13g2_decap_8 FILLER_14_191 ();
 sg13g2_decap_4 FILLER_14_198 ();
 sg13g2_fill_2 FILLER_14_212 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_4 FILLER_14_224 ();
 sg13g2_fill_2 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_234 ();
 sg13g2_decap_4 FILLER_14_241 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_4 FILLER_14_272 ();
 sg13g2_fill_2 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_decap_4 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_fill_2 FILLER_14_327 ();
 sg13g2_fill_1 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_4 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_4 FILLER_14_382 ();
 sg13g2_fill_2 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_401 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_decap_8 FILLER_14_419 ();
 sg13g2_decap_4 FILLER_14_426 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_16 ();
 sg13g2_fill_2 FILLER_15_23 ();
 sg13g2_fill_1 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_31 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_fill_2 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_83 ();
 sg13g2_decap_8 FILLER_15_90 ();
 sg13g2_decap_8 FILLER_15_97 ();
 sg13g2_decap_8 FILLER_15_104 ();
 sg13g2_decap_8 FILLER_15_111 ();
 sg13g2_fill_1 FILLER_15_118 ();
 sg13g2_decap_4 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_127 ();
 sg13g2_decap_4 FILLER_15_159 ();
 sg13g2_fill_2 FILLER_15_163 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_decap_4 FILLER_15_176 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_fill_2 FILLER_15_225 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_4 FILLER_15_268 ();
 sg13g2_fill_1 FILLER_15_272 ();
 sg13g2_decap_4 FILLER_15_286 ();
 sg13g2_fill_2 FILLER_15_290 ();
 sg13g2_fill_2 FILLER_15_296 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_fill_2 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_305 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_4 FILLER_15_327 ();
 sg13g2_fill_2 FILLER_15_331 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_fill_1 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_4 ();
 sg13g2_fill_1 FILLER_16_62 ();
 sg13g2_decap_8 FILLER_16_93 ();
 sg13g2_decap_4 FILLER_16_100 ();
 sg13g2_fill_1 FILLER_16_104 ();
 sg13g2_decap_8 FILLER_16_131 ();
 sg13g2_decap_8 FILLER_16_138 ();
 sg13g2_fill_1 FILLER_16_145 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_decap_8 FILLER_16_184 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_197 ();
 sg13g2_decap_8 FILLER_16_204 ();
 sg13g2_decap_4 FILLER_16_211 ();
 sg13g2_fill_2 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_decap_4 FILLER_16_237 ();
 sg13g2_fill_1 FILLER_16_241 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_fill_1 FILLER_16_281 ();
 sg13g2_fill_1 FILLER_16_290 ();
 sg13g2_decap_4 FILLER_16_296 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_1 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_320 ();
 sg13g2_fill_2 FILLER_16_327 ();
 sg13g2_fill_1 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_fill_2 FILLER_16_361 ();
 sg13g2_fill_1 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_383 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_fill_1 FILLER_16_397 ();
 sg13g2_decap_4 FILLER_16_402 ();
 sg13g2_fill_1 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_419 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_2 FILLER_17_14 ();
 sg13g2_fill_1 FILLER_17_16 ();
 sg13g2_decap_8 FILLER_17_32 ();
 sg13g2_fill_1 FILLER_17_39 ();
 sg13g2_decap_8 FILLER_17_45 ();
 sg13g2_fill_2 FILLER_17_52 ();
 sg13g2_fill_2 FILLER_17_64 ();
 sg13g2_decap_8 FILLER_17_75 ();
 sg13g2_decap_8 FILLER_17_82 ();
 sg13g2_fill_1 FILLER_17_89 ();
 sg13g2_fill_2 FILLER_17_110 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_117 ();
 sg13g2_decap_8 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_135 ();
 sg13g2_decap_4 FILLER_17_151 ();
 sg13g2_fill_2 FILLER_17_155 ();
 sg13g2_decap_4 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_166 ();
 sg13g2_decap_8 FILLER_17_181 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_decap_8 FILLER_17_201 ();
 sg13g2_decap_8 FILLER_17_208 ();
 sg13g2_fill_2 FILLER_17_225 ();
 sg13g2_decap_4 FILLER_17_235 ();
 sg13g2_decap_4 FILLER_17_243 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_fill_2 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_269 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_fill_1 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_302 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_316 ();
 sg13g2_decap_4 FILLER_17_323 ();
 sg13g2_fill_2 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_4 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_4 FILLER_17_424 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_25 ();
 sg13g2_decap_4 FILLER_18_32 ();
 sg13g2_decap_8 FILLER_18_40 ();
 sg13g2_decap_8 FILLER_18_47 ();
 sg13g2_decap_8 FILLER_18_54 ();
 sg13g2_decap_8 FILLER_18_61 ();
 sg13g2_decap_4 FILLER_18_68 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_decap_4 FILLER_18_88 ();
 sg13g2_fill_1 FILLER_18_92 ();
 sg13g2_decap_8 FILLER_18_111 ();
 sg13g2_decap_8 FILLER_18_118 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_129 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_fill_1 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_145 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_fill_1 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_177 ();
 sg13g2_decap_4 FILLER_18_195 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_decap_8 FILLER_18_234 ();
 sg13g2_decap_4 FILLER_18_241 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_260 ();
 sg13g2_fill_1 FILLER_18_269 ();
 sg13g2_decap_4 FILLER_18_276 ();
 sg13g2_fill_1 FILLER_18_285 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_296 ();
 sg13g2_fill_2 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_decap_4 FILLER_18_332 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_fill_2 FILLER_18_359 ();
 sg13g2_fill_1 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_fill_1 FILLER_18_385 ();
 sg13g2_decap_4 FILLER_18_398 ();
 sg13g2_fill_2 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_27 ();
 sg13g2_decap_8 FILLER_19_55 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_decap_8 FILLER_19_131 ();
 sg13g2_decap_8 FILLER_19_138 ();
 sg13g2_decap_8 FILLER_19_145 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_169 ();
 sg13g2_decap_8 FILLER_19_176 ();
 sg13g2_decap_8 FILLER_19_183 ();
 sg13g2_decap_4 FILLER_19_190 ();
 sg13g2_fill_1 FILLER_19_194 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_decap_8 FILLER_19_268 ();
 sg13g2_fill_2 FILLER_19_279 ();
 sg13g2_fill_1 FILLER_19_281 ();
 sg13g2_fill_2 FILLER_19_305 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_4 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_decap_4 FILLER_19_363 ();
 sg13g2_decap_8 FILLER_19_423 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_11 ();
 sg13g2_fill_2 FILLER_20_18 ();
 sg13g2_fill_2 FILLER_20_35 ();
 sg13g2_fill_1 FILLER_20_37 ();
 sg13g2_fill_2 FILLER_20_43 ();
 sg13g2_fill_2 FILLER_20_49 ();
 sg13g2_fill_1 FILLER_20_51 ();
 sg13g2_fill_1 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_fill_2 FILLER_20_74 ();
 sg13g2_fill_1 FILLER_20_76 ();
 sg13g2_decap_4 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_85 ();
 sg13g2_decap_8 FILLER_20_93 ();
 sg13g2_decap_8 FILLER_20_100 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_114 ();
 sg13g2_fill_2 FILLER_20_121 ();
 sg13g2_fill_1 FILLER_20_123 ();
 sg13g2_decap_4 FILLER_20_132 ();
 sg13g2_fill_1 FILLER_20_144 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_fill_1 FILLER_20_163 ();
 sg13g2_fill_1 FILLER_20_169 ();
 sg13g2_decap_4 FILLER_20_178 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_4 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_225 ();
 sg13g2_decap_4 FILLER_20_232 ();
 sg13g2_decap_8 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_265 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_fill_1 FILLER_20_279 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_293 ();
 sg13g2_fill_1 FILLER_20_300 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_decap_4 FILLER_20_313 ();
 sg13g2_fill_2 FILLER_20_317 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_fill_2 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_349 ();
 sg13g2_decap_4 FILLER_20_366 ();
 sg13g2_fill_2 FILLER_20_370 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_fill_2 FILLER_20_400 ();
 sg13g2_fill_1 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_20_414 ();
 sg13g2_decap_8 FILLER_20_421 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_4 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_40 ();
 sg13g2_decap_8 FILLER_21_47 ();
 sg13g2_decap_4 FILLER_21_54 ();
 sg13g2_decap_4 FILLER_21_64 ();
 sg13g2_decap_4 FILLER_21_71 ();
 sg13g2_fill_2 FILLER_21_75 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_114 ();
 sg13g2_decap_4 FILLER_21_121 ();
 sg13g2_fill_2 FILLER_21_125 ();
 sg13g2_decap_8 FILLER_21_145 ();
 sg13g2_fill_2 FILLER_21_152 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_167 ();
 sg13g2_fill_2 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_181 ();
 sg13g2_decap_4 FILLER_21_186 ();
 sg13g2_fill_1 FILLER_21_190 ();
 sg13g2_decap_4 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_211 ();
 sg13g2_decap_4 FILLER_21_220 ();
 sg13g2_decap_8 FILLER_21_255 ();
 sg13g2_decap_8 FILLER_21_262 ();
 sg13g2_decap_8 FILLER_21_269 ();
 sg13g2_fill_1 FILLER_21_276 ();
 sg13g2_fill_2 FILLER_21_293 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_4 FILLER_21_320 ();
 sg13g2_fill_1 FILLER_21_328 ();
 sg13g2_fill_2 FILLER_21_334 ();
 sg13g2_fill_1 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_4 FILLER_21_369 ();
 sg13g2_fill_1 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_fill_1 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_4 FILLER_21_399 ();
 sg13g2_fill_1 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_22_26 ();
 sg13g2_fill_1 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_60 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_decap_8 FILLER_22_92 ();
 sg13g2_decap_4 FILLER_22_99 ();
 sg13g2_decap_4 FILLER_22_109 ();
 sg13g2_fill_1 FILLER_22_113 ();
 sg13g2_fill_1 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_124 ();
 sg13g2_fill_2 FILLER_22_131 ();
 sg13g2_fill_2 FILLER_22_138 ();
 sg13g2_fill_1 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_167 ();
 sg13g2_fill_1 FILLER_22_174 ();
 sg13g2_decap_4 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_215 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_decap_8 FILLER_22_229 ();
 sg13g2_fill_2 FILLER_22_236 ();
 sg13g2_fill_1 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_decap_8 FILLER_22_251 ();
 sg13g2_decap_8 FILLER_22_258 ();
 sg13g2_decap_8 FILLER_22_265 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_320 ();
 sg13g2_decap_4 FILLER_22_357 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_fill_1 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_8 FILLER_22_405 ();
 sg13g2_fill_1 FILLER_22_412 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_4 FILLER_22_424 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_12 ();
 sg13g2_fill_1 FILLER_23_26 ();
 sg13g2_decap_8 FILLER_23_59 ();
 sg13g2_decap_4 FILLER_23_66 ();
 sg13g2_fill_2 FILLER_23_75 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_90 ();
 sg13g2_fill_2 FILLER_23_95 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_fill_1 FILLER_23_114 ();
 sg13g2_fill_2 FILLER_23_132 ();
 sg13g2_fill_1 FILLER_23_134 ();
 sg13g2_fill_1 FILLER_23_153 ();
 sg13g2_fill_2 FILLER_23_171 ();
 sg13g2_fill_1 FILLER_23_173 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_fill_2 FILLER_23_186 ();
 sg13g2_fill_1 FILLER_23_188 ();
 sg13g2_fill_1 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_202 ();
 sg13g2_decap_8 FILLER_23_209 ();
 sg13g2_decap_8 FILLER_23_216 ();
 sg13g2_fill_2 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_225 ();
 sg13g2_decap_4 FILLER_23_236 ();
 sg13g2_fill_1 FILLER_23_240 ();
 sg13g2_fill_2 FILLER_23_259 ();
 sg13g2_fill_1 FILLER_23_261 ();
 sg13g2_decap_8 FILLER_23_276 ();
 sg13g2_decap_4 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_411 ();
 sg13g2_decap_8 FILLER_23_418 ();
 sg13g2_decap_4 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_51 ();
 sg13g2_fill_1 FILLER_24_57 ();
 sg13g2_decap_8 FILLER_24_83 ();
 sg13g2_decap_4 FILLER_24_90 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_fill_1 FILLER_24_106 ();
 sg13g2_decap_4 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_116 ();
 sg13g2_decap_4 FILLER_24_126 ();
 sg13g2_fill_2 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_decap_8 FILLER_24_180 ();
 sg13g2_decap_4 FILLER_24_187 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_decap_4 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_decap_8 FILLER_24_219 ();
 sg13g2_decap_8 FILLER_24_226 ();
 sg13g2_fill_2 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_267 ();
 sg13g2_fill_2 FILLER_24_274 ();
 sg13g2_fill_2 FILLER_24_309 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_1 FILLER_24_368 ();
 sg13g2_fill_1 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_384 ();
 sg13g2_fill_1 FILLER_24_397 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_11 ();
 sg13g2_decap_4 FILLER_25_18 ();
 sg13g2_fill_1 FILLER_25_22 ();
 sg13g2_decap_8 FILLER_25_33 ();
 sg13g2_decap_8 FILLER_25_40 ();
 sg13g2_decap_8 FILLER_25_47 ();
 sg13g2_fill_2 FILLER_25_54 ();
 sg13g2_fill_2 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_62 ();
 sg13g2_fill_2 FILLER_25_73 ();
 sg13g2_fill_1 FILLER_25_75 ();
 sg13g2_decap_4 FILLER_25_90 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_131 ();
 sg13g2_decap_4 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_142 ();
 sg13g2_decap_8 FILLER_25_152 ();
 sg13g2_decap_8 FILLER_25_159 ();
 sg13g2_decap_4 FILLER_25_166 ();
 sg13g2_fill_2 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_4 FILLER_25_214 ();
 sg13g2_fill_1 FILLER_25_218 ();
 sg13g2_fill_1 FILLER_25_230 ();
 sg13g2_fill_2 FILLER_25_236 ();
 sg13g2_decap_8 FILLER_25_244 ();
 sg13g2_decap_8 FILLER_25_251 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_fill_2 FILLER_25_272 ();
 sg13g2_fill_1 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_285 ();
 sg13g2_decap_4 FILLER_25_292 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_fill_2 FILLER_25_329 ();
 sg13g2_fill_1 FILLER_25_331 ();
 sg13g2_fill_1 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_4 FILLER_25_356 ();
 sg13g2_decap_4 FILLER_25_373 ();
 sg13g2_fill_2 FILLER_25_377 ();
 sg13g2_decap_4 FILLER_25_388 ();
 sg13g2_fill_1 FILLER_25_392 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_2 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_25_414 ();
 sg13g2_decap_8 FILLER_25_421 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_4 FILLER_26_31 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_40 ();
 sg13g2_fill_1 FILLER_26_44 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_decap_8 FILLER_26_76 ();
 sg13g2_decap_8 FILLER_26_83 ();
 sg13g2_decap_4 FILLER_26_90 ();
 sg13g2_fill_2 FILLER_26_99 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_107 ();
 sg13g2_decap_8 FILLER_26_114 ();
 sg13g2_decap_4 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_4 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_206 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_decap_4 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_decap_4 FILLER_26_236 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_289 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_310 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_decap_8 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_331 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_4 FILLER_26_350 ();
 sg13g2_fill_1 FILLER_26_354 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_fill_1 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_fill_2 FILLER_26_396 ();
 sg13g2_fill_1 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_26_404 ();
 sg13g2_decap_8 FILLER_26_411 ();
 sg13g2_decap_8 FILLER_26_418 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_15 ();
 sg13g2_fill_2 FILLER_27_22 ();
 sg13g2_fill_1 FILLER_27_55 ();
 sg13g2_decap_8 FILLER_27_66 ();
 sg13g2_fill_1 FILLER_27_73 ();
 sg13g2_fill_2 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_decap_4 FILLER_27_86 ();
 sg13g2_fill_2 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_104 ();
 sg13g2_decap_8 FILLER_27_111 ();
 sg13g2_decap_8 FILLER_27_118 ();
 sg13g2_decap_4 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_129 ();
 sg13g2_decap_8 FILLER_27_144 ();
 sg13g2_decap_8 FILLER_27_151 ();
 sg13g2_decap_8 FILLER_27_158 ();
 sg13g2_decap_4 FILLER_27_165 ();
 sg13g2_decap_8 FILLER_27_174 ();
 sg13g2_decap_4 FILLER_27_181 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_fill_2 FILLER_27_191 ();
 sg13g2_decap_4 FILLER_27_206 ();
 sg13g2_fill_2 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_fill_1 FILLER_27_224 ();
 sg13g2_decap_4 FILLER_27_234 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_246 ();
 sg13g2_decap_4 FILLER_27_258 ();
 sg13g2_decap_8 FILLER_27_269 ();
 sg13g2_decap_4 FILLER_27_276 ();
 sg13g2_fill_2 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_288 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_297 ();
 sg13g2_decap_8 FILLER_27_306 ();
 sg13g2_decap_8 FILLER_27_313 ();
 sg13g2_fill_2 FILLER_27_324 ();
 sg13g2_fill_1 FILLER_27_326 ();
 sg13g2_decap_4 FILLER_27_349 ();
 sg13g2_fill_1 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_365 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_fill_2 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_403 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_4 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_24 ();
 sg13g2_decap_4 FILLER_28_41 ();
 sg13g2_fill_1 FILLER_28_45 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_4 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_76 ();
 sg13g2_fill_2 FILLER_28_83 ();
 sg13g2_fill_1 FILLER_28_85 ();
 sg13g2_fill_2 FILLER_28_89 ();
 sg13g2_fill_1 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_100 ();
 sg13g2_decap_8 FILLER_28_106 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_137 ();
 sg13g2_fill_1 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_decap_4 FILLER_28_180 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_209 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_decap_4 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_220 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_decap_4 FILLER_28_234 ();
 sg13g2_fill_1 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_259 ();
 sg13g2_fill_1 FILLER_28_261 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_fill_2 FILLER_28_287 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_decap_4 FILLER_28_321 ();
 sg13g2_fill_2 FILLER_28_333 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_decap_4 FILLER_28_385 ();
 sg13g2_fill_1 FILLER_28_389 ();
 sg13g2_fill_2 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_403 ();
 sg13g2_fill_1 FILLER_28_410 ();
 sg13g2_decap_8 FILLER_28_415 ();
 sg13g2_decap_8 FILLER_28_422 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_36 ();
 sg13g2_fill_2 FILLER_29_43 ();
 sg13g2_fill_1 FILLER_29_45 ();
 sg13g2_decap_8 FILLER_29_55 ();
 sg13g2_fill_2 FILLER_29_62 ();
 sg13g2_fill_1 FILLER_29_64 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_decap_4 FILLER_29_102 ();
 sg13g2_decap_8 FILLER_29_125 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_decap_8 FILLER_29_139 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_decap_4 FILLER_29_153 ();
 sg13g2_fill_2 FILLER_29_157 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_decap_8 FILLER_29_188 ();
 sg13g2_decap_4 FILLER_29_195 ();
 sg13g2_fill_2 FILLER_29_199 ();
 sg13g2_fill_1 FILLER_29_209 ();
 sg13g2_fill_2 FILLER_29_215 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_fill_1 FILLER_29_242 ();
 sg13g2_fill_1 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_decap_8 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_decap_8 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_fill_1 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_fill_1 FILLER_29_389 ();
 sg13g2_fill_2 FILLER_29_404 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_15 ();
 sg13g2_fill_1 FILLER_30_19 ();
 sg13g2_decap_4 FILLER_30_40 ();
 sg13g2_fill_1 FILLER_30_44 ();
 sg13g2_decap_8 FILLER_30_76 ();
 sg13g2_fill_2 FILLER_30_83 ();
 sg13g2_fill_1 FILLER_30_85 ();
 sg13g2_fill_1 FILLER_30_89 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_190 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_257 ();
 sg13g2_decap_8 FILLER_30_264 ();
 sg13g2_decap_8 FILLER_30_271 ();
 sg13g2_decap_8 FILLER_30_278 ();
 sg13g2_decap_4 FILLER_30_285 ();
 sg13g2_decap_8 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_327 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_fill_2 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_fill_1 FILLER_30_385 ();
 sg13g2_fill_2 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_decap_8 FILLER_30_409 ();
 sg13g2_decap_8 FILLER_30_416 ();
 sg13g2_decap_8 FILLER_30_423 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_21 ();
 sg13g2_fill_1 FILLER_31_23 ();
 sg13g2_fill_2 FILLER_31_33 ();
 sg13g2_fill_1 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_45 ();
 sg13g2_decap_4 FILLER_31_52 ();
 sg13g2_fill_2 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_62 ();
 sg13g2_decap_8 FILLER_31_69 ();
 sg13g2_decap_8 FILLER_31_76 ();
 sg13g2_fill_1 FILLER_31_83 ();
 sg13g2_decap_8 FILLER_31_104 ();
 sg13g2_fill_2 FILLER_31_111 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_128 ();
 sg13g2_fill_2 FILLER_31_135 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_decap_4 FILLER_31_144 ();
 sg13g2_fill_2 FILLER_31_148 ();
 sg13g2_fill_2 FILLER_31_155 ();
 sg13g2_fill_2 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_decap_8 FILLER_31_188 ();
 sg13g2_fill_2 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_208 ();
 sg13g2_decap_8 FILLER_31_215 ();
 sg13g2_decap_4 FILLER_31_222 ();
 sg13g2_fill_1 FILLER_31_226 ();
 sg13g2_decap_8 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_261 ();
 sg13g2_decap_4 FILLER_31_268 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_313 ();
 sg13g2_decap_8 FILLER_31_319 ();
 sg13g2_decap_4 FILLER_31_340 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_decap_4 FILLER_31_362 ();
 sg13g2_decap_4 FILLER_31_370 ();
 sg13g2_fill_1 FILLER_31_374 ();
 sg13g2_fill_1 FILLER_31_391 ();
 sg13g2_decap_8 FILLER_31_411 ();
 sg13g2_decap_8 FILLER_31_418 ();
 sg13g2_decap_4 FILLER_31_425 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_4 FILLER_32_21 ();
 sg13g2_decap_4 FILLER_32_30 ();
 sg13g2_fill_1 FILLER_32_60 ();
 sg13g2_fill_2 FILLER_32_69 ();
 sg13g2_decap_8 FILLER_32_80 ();
 sg13g2_fill_2 FILLER_32_87 ();
 sg13g2_decap_8 FILLER_32_103 ();
 sg13g2_decap_4 FILLER_32_110 ();
 sg13g2_fill_2 FILLER_32_118 ();
 sg13g2_fill_1 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_125 ();
 sg13g2_fill_1 FILLER_32_127 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_decap_4 FILLER_32_148 ();
 sg13g2_fill_2 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_172 ();
 sg13g2_fill_2 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_decap_4 FILLER_32_216 ();
 sg13g2_fill_1 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_257 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_fill_2 FILLER_32_298 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_decap_4 FILLER_32_312 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_decap_8 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_fill_2 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_decap_4 FILLER_32_374 ();
 sg13g2_decap_4 FILLER_32_390 ();
 sg13g2_fill_1 FILLER_32_394 ();
 sg13g2_decap_4 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_417 ();
 sg13g2_decap_4 FILLER_32_424 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_61 ();
 sg13g2_fill_2 FILLER_33_68 ();
 sg13g2_fill_1 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_92 ();
 sg13g2_decap_8 FILLER_33_104 ();
 sg13g2_decap_4 FILLER_33_111 ();
 sg13g2_fill_1 FILLER_33_115 ();
 sg13g2_decap_8 FILLER_33_129 ();
 sg13g2_decap_8 FILLER_33_136 ();
 sg13g2_decap_4 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_decap_8 FILLER_33_163 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_184 ();
 sg13g2_decap_8 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_204 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_215 ();
 sg13g2_fill_2 FILLER_33_221 ();
 sg13g2_decap_4 FILLER_33_228 ();
 sg13g2_decap_4 FILLER_33_240 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_decap_8 FILLER_33_250 ();
 sg13g2_decap_8 FILLER_33_257 ();
 sg13g2_fill_2 FILLER_33_264 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_279 ();
 sg13g2_fill_2 FILLER_33_286 ();
 sg13g2_fill_1 FILLER_33_288 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_339 ();
 sg13g2_fill_2 FILLER_33_345 ();
 sg13g2_fill_2 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_decap_4 FILLER_33_364 ();
 sg13g2_fill_1 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_fill_2 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_424 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_9 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_21 ();
 sg13g2_fill_1 FILLER_34_23 ();
 sg13g2_decap_8 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_41 ();
 sg13g2_fill_2 FILLER_34_47 ();
 sg13g2_fill_1 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_55 ();
 sg13g2_decap_4 FILLER_34_62 ();
 sg13g2_fill_2 FILLER_34_66 ();
 sg13g2_decap_8 FILLER_34_73 ();
 sg13g2_decap_4 FILLER_34_80 ();
 sg13g2_fill_2 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_102 ();
 sg13g2_decap_4 FILLER_34_109 ();
 sg13g2_fill_2 FILLER_34_113 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_decap_4 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_151 ();
 sg13g2_decap_8 FILLER_34_178 ();
 sg13g2_decap_4 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_194 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_fill_2 FILLER_34_212 ();
 sg13g2_decap_4 FILLER_34_219 ();
 sg13g2_fill_2 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_230 ();
 sg13g2_fill_2 FILLER_34_238 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_decap_4 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_249 ();
 sg13g2_fill_2 FILLER_34_257 ();
 sg13g2_fill_1 FILLER_34_271 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_decap_4 FILLER_34_305 ();
 sg13g2_decap_8 FILLER_34_314 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_decap_4 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_332 ();
 sg13g2_decap_4 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_34_351 ();
 sg13g2_decap_4 FILLER_34_358 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_decap_4 FILLER_34_375 ();
 sg13g2_fill_1 FILLER_34_379 ();
 sg13g2_fill_1 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_fill_1 FILLER_34_409 ();
 sg13g2_decap_8 FILLER_34_414 ();
 sg13g2_decap_8 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_11 ();
 sg13g2_fill_2 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_23 ();
 sg13g2_decap_8 FILLER_35_29 ();
 sg13g2_decap_8 FILLER_35_36 ();
 sg13g2_fill_2 FILLER_35_78 ();
 sg13g2_fill_1 FILLER_35_80 ();
 sg13g2_decap_4 FILLER_35_86 ();
 sg13g2_fill_2 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_122 ();
 sg13g2_decap_8 FILLER_35_127 ();
 sg13g2_decap_8 FILLER_35_134 ();
 sg13g2_decap_8 FILLER_35_141 ();
 sg13g2_decap_8 FILLER_35_148 ();
 sg13g2_decap_4 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_159 ();
 sg13g2_decap_8 FILLER_35_167 ();
 sg13g2_decap_4 FILLER_35_174 ();
 sg13g2_decap_4 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_decap_8 FILLER_35_215 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_261 ();
 sg13g2_decap_8 FILLER_35_268 ();
 sg13g2_fill_2 FILLER_35_275 ();
 sg13g2_fill_1 FILLER_35_277 ();
 sg13g2_fill_2 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_decap_4 FILLER_35_337 ();
 sg13g2_fill_1 FILLER_35_341 ();
 sg13g2_decap_4 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_2 FILLER_35_357 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_fill_2 FILLER_35_370 ();
 sg13g2_fill_1 FILLER_35_372 ();
 sg13g2_decap_4 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_391 ();
 sg13g2_fill_1 FILLER_35_402 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_34 ();
 sg13g2_decap_8 FILLER_36_41 ();
 sg13g2_decap_8 FILLER_36_52 ();
 sg13g2_decap_8 FILLER_36_59 ();
 sg13g2_decap_8 FILLER_36_66 ();
 sg13g2_decap_8 FILLER_36_73 ();
 sg13g2_decap_8 FILLER_36_80 ();
 sg13g2_decap_8 FILLER_36_87 ();
 sg13g2_decap_4 FILLER_36_94 ();
 sg13g2_fill_1 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_103 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_117 ();
 sg13g2_decap_8 FILLER_36_124 ();
 sg13g2_decap_4 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_fill_2 FILLER_36_182 ();
 sg13g2_decap_4 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_decap_8 FILLER_36_204 ();
 sg13g2_decap_8 FILLER_36_211 ();
 sg13g2_decap_8 FILLER_36_218 ();
 sg13g2_fill_2 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_decap_4 FILLER_36_246 ();
 sg13g2_fill_1 FILLER_36_250 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_299 ();
 sg13g2_decap_8 FILLER_36_306 ();
 sg13g2_decap_4 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_335 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_fill_2 FILLER_36_348 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_decap_4 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_391 ();
 sg13g2_decap_8 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_fill_2 FILLER_36_409 ();
 sg13g2_decap_8 FILLER_36_416 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_fill_2 FILLER_37_36 ();
 sg13g2_fill_1 FILLER_37_38 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_4 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_88 ();
 sg13g2_decap_4 FILLER_37_97 ();
 sg13g2_decap_8 FILLER_37_131 ();
 sg13g2_decap_4 FILLER_37_138 ();
 sg13g2_fill_2 FILLER_37_142 ();
 sg13g2_decap_4 FILLER_37_178 ();
 sg13g2_fill_2 FILLER_37_182 ();
 sg13g2_decap_4 FILLER_37_210 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_decap_8 FILLER_37_261 ();
 sg13g2_decap_8 FILLER_37_268 ();
 sg13g2_decap_8 FILLER_37_275 ();
 sg13g2_decap_8 FILLER_37_282 ();
 sg13g2_decap_8 FILLER_37_289 ();
 sg13g2_decap_8 FILLER_37_296 ();
 sg13g2_decap_8 FILLER_37_303 ();
 sg13g2_decap_4 FILLER_37_310 ();
 sg13g2_fill_2 FILLER_37_314 ();
 sg13g2_fill_2 FILLER_37_320 ();
 sg13g2_decap_4 FILLER_37_327 ();
 sg13g2_fill_1 FILLER_37_331 ();
 sg13g2_fill_1 FILLER_37_341 ();
 sg13g2_decap_4 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_355 ();
 sg13g2_decap_4 FILLER_37_372 ();
 sg13g2_fill_1 FILLER_37_376 ();
 sg13g2_fill_1 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_390 ();
 sg13g2_fill_1 FILLER_37_421 ();
 sg13g2_decap_4 FILLER_37_426 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_11 ();
 sg13g2_decap_8 FILLER_38_16 ();
 sg13g2_decap_8 FILLER_38_23 ();
 sg13g2_decap_8 FILLER_38_30 ();
 sg13g2_decap_8 FILLER_38_37 ();
 sg13g2_decap_4 FILLER_38_44 ();
 sg13g2_decap_8 FILLER_38_52 ();
 sg13g2_decap_8 FILLER_38_59 ();
 sg13g2_decap_4 FILLER_38_66 ();
 sg13g2_fill_1 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_91 ();
 sg13g2_fill_2 FILLER_38_120 ();
 sg13g2_fill_1 FILLER_38_130 ();
 sg13g2_fill_1 FILLER_38_135 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_145 ();
 sg13g2_fill_1 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_38_209 ();
 sg13g2_fill_2 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_4 FILLER_38_299 ();
 sg13g2_decap_4 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_320 ();
 sg13g2_decap_4 FILLER_38_325 ();
 sg13g2_fill_2 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_fill_2 FILLER_38_427 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
