module tt_um_toivoh_retro_console (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire clknet_leaf_0_clk;
 wire active;
 wire \addr_pins_out[0] ;
 wire \addr_pins_out[1] ;
 wire \addr_pins_out[2] ;
 wire \addr_pins_out[3] ;
 wire \data_pins[0] ;
 wire \data_pins[1] ;
 wire \data_pins[2] ;
 wire \data_pins[3] ;
 wire dither_out;
 wire drive_uio_76;
 wire hsync;
 wire \ppu.b0_out[1] ;
 wire \ppu.b0_out[2] ;
 wire \ppu.b0_out[3] ;
 wire \ppu.base_addr_regs[0][0] ;
 wire \ppu.base_addr_regs[0][1] ;
 wire \ppu.base_addr_regs[0][2] ;
 wire \ppu.base_addr_regs[0][3] ;
 wire \ppu.base_addr_regs[0][4] ;
 wire \ppu.base_addr_regs[0][5] ;
 wire \ppu.base_addr_regs[0][6] ;
 wire \ppu.base_addr_regs[0][7] ;
 wire \ppu.base_addr_regs[0][8] ;
 wire \ppu.base_addr_regs[1][0] ;
 wire \ppu.base_addr_regs[1][1] ;
 wire \ppu.base_addr_regs[1][2] ;
 wire \ppu.base_addr_regs[1][3] ;
 wire \ppu.base_addr_regs[1][4] ;
 wire \ppu.base_addr_regs[1][5] ;
 wire \ppu.base_addr_regs[1][6] ;
 wire \ppu.base_addr_regs[1][7] ;
 wire \ppu.base_addr_regs[1][8] ;
 wire \ppu.base_addr_regs[2][1] ;
 wire \ppu.base_addr_regs[2][2] ;
 wire \ppu.base_addr_regs[2][3] ;
 wire \ppu.base_addr_regs[2][4] ;
 wire \ppu.base_addr_regs[2][5] ;
 wire \ppu.base_addr_regs[2][6] ;
 wire \ppu.base_addr_regs[2][7] ;
 wire \ppu.base_addr_regs[2][8] ;
 wire \ppu.base_addr_regs[3][1] ;
 wire \ppu.base_addr_regs[3][2] ;
 wire \ppu.base_addr_regs[3][3] ;
 wire \ppu.base_addr_regs[3][4] ;
 wire \ppu.copper_inst.addr[0] ;
 wire \ppu.copper_inst.addr[10] ;
 wire \ppu.copper_inst.addr[11] ;
 wire \ppu.copper_inst.addr[12] ;
 wire \ppu.copper_inst.addr[13] ;
 wire \ppu.copper_inst.addr[14] ;
 wire \ppu.copper_inst.addr[15] ;
 wire \ppu.copper_inst.addr[1] ;
 wire \ppu.copper_inst.addr[2] ;
 wire \ppu.copper_inst.addr[3] ;
 wire \ppu.copper_inst.addr[4] ;
 wire \ppu.copper_inst.addr[5] ;
 wire \ppu.copper_inst.addr[6] ;
 wire \ppu.copper_inst.addr[7] ;
 wire \ppu.copper_inst.addr[8] ;
 wire \ppu.copper_inst.addr[9] ;
 wire \ppu.copper_inst.cmp[0] ;
 wire \ppu.copper_inst.cmp[1] ;
 wire \ppu.copper_inst.cmp[2] ;
 wire \ppu.copper_inst.cmp[3] ;
 wire \ppu.copper_inst.cmp[4] ;
 wire \ppu.copper_inst.cmp[5] ;
 wire \ppu.copper_inst.cmp[6] ;
 wire \ppu.copper_inst.cmp[7] ;
 wire \ppu.copper_inst.cmp[8] ;
 wire \ppu.copper_inst.cmp_on ;
 wire \ppu.copper_inst.cmp_type ;
 wire \ppu.copper_inst.dt_out[0] ;
 wire \ppu.copper_inst.dt_out[1] ;
 wire \ppu.copper_inst.dt_out[2] ;
 wire \ppu.copper_inst.dt_sreg[10] ;
 wire \ppu.copper_inst.dt_sreg[11] ;
 wire \ppu.copper_inst.dt_sreg[3] ;
 wire \ppu.copper_inst.dt_sreg[4] ;
 wire \ppu.copper_inst.dt_sreg[5] ;
 wire \ppu.copper_inst.dt_sreg[6] ;
 wire \ppu.copper_inst.dt_sreg[7] ;
 wire \ppu.copper_inst.dt_sreg[8] ;
 wire \ppu.copper_inst.dt_sreg[9] ;
 wire \ppu.copper_inst.fast_mode ;
 wire \ppu.copper_inst.on ;
 wire \ppu.copper_inst.serial_counter[0] ;
 wire \ppu.copper_inst.serial_counter[1] ;
 wire \ppu.copper_inst.store[0] ;
 wire \ppu.copper_inst.store[10] ;
 wire \ppu.copper_inst.store[11] ;
 wire \ppu.copper_inst.store[12] ;
 wire \ppu.copper_inst.store[13] ;
 wire \ppu.copper_inst.store[14] ;
 wire \ppu.copper_inst.store[15] ;
 wire \ppu.copper_inst.store[1] ;
 wire \ppu.copper_inst.store[2] ;
 wire \ppu.copper_inst.store[3] ;
 wire \ppu.copper_inst.store[4] ;
 wire \ppu.copper_inst.store[5] ;
 wire \ppu.copper_inst.store[6] ;
 wire \ppu.copper_inst.store[7] ;
 wire \ppu.copper_inst.store[8] ;
 wire \ppu.copper_inst.store[9] ;
 wire \ppu.copper_inst.store_valid ;
 wire \ppu.copper_inst.x_cmp[0] ;
 wire \ppu.copper_inst.x_cmp[1] ;
 wire \ppu.copper_inst.x_cmp[2] ;
 wire \ppu.copper_inst.x_cmp[3] ;
 wire \ppu.copper_inst.x_cmp[4] ;
 wire \ppu.copper_inst.x_cmp[8] ;
 wire \ppu.curr_pal_addr[0] ;
 wire \ppu.curr_pal_addr[1] ;
 wire \ppu.curr_pal_addr[2] ;
 wire \ppu.curr_pal_addr[3] ;
 wire \ppu.depth_out_s[0] ;
 wire \ppu.depth_out_s[1] ;
 wire \ppu.depth_out_t[0] ;
 wire \ppu.depth_out_t[1] ;
 wire \ppu.display_mask[0] ;
 wire \ppu.display_mask[1] ;
 wire \ppu.display_mask[2] ;
 wire \ppu.display_mask[3] ;
 wire \ppu.display_mask[4] ;
 wire \ppu.display_mask[5] ;
 wire \ppu.dither_g.u[0] ;
 wire \ppu.dither_g.u[1] ;
 wire \ppu.dither_g.u[2] ;
 wire \ppu.dither_r.u[1] ;
 wire \ppu.dither_r.u[2] ;
 wire \ppu.gfxmode1[0] ;
 wire \ppu.gfxmode1[1] ;
 wire \ppu.gfxmode1[2] ;
 wire \ppu.gfxmode1[3] ;
 wire \ppu.gfxmode1[4] ;
 wire \ppu.gfxmode1[5] ;
 wire \ppu.gfxmode1[6] ;
 wire \ppu.gfxmode1[7] ;
 wire \ppu.gfxmode1[8] ;
 wire \ppu.gfxmode2[0] ;
 wire \ppu.gfxmode2[1] ;
 wire \ppu.gfxmode2[2] ;
 wire \ppu.gfxmode2[3] ;
 wire \ppu.gfxmode2[4] ;
 wire \ppu.gfxmode2[5] ;
 wire \ppu.gfxmode2[6] ;
 wire \ppu.gfxmode2[7] ;
 wire \ppu.gfxmode2[8] ;
 wire \ppu.gfxmode3[0] ;
 wire \ppu.gfxmode3[1] ;
 wire \ppu.gfxmode3[2] ;
 wire \ppu.gfxmode3[3] ;
 wire \ppu.gfxmode3[4] ;
 wire \ppu.gfxmode3[5] ;
 wire \ppu.gfxmode3[6] ;
 wire \ppu.gfxmode3[7] ;
 wire \ppu.gfxmode3[8] ;
 wire \ppu.pal[0][0] ;
 wire \ppu.pal[0][1] ;
 wire \ppu.pal[0][2] ;
 wire \ppu.pal[0][3] ;
 wire \ppu.pal[0][4] ;
 wire \ppu.pal[0][5] ;
 wire \ppu.pal[0][6] ;
 wire \ppu.pal[0][7] ;
 wire \ppu.pal[10][0] ;
 wire \ppu.pal[10][1] ;
 wire \ppu.pal[10][2] ;
 wire \ppu.pal[10][3] ;
 wire \ppu.pal[10][4] ;
 wire \ppu.pal[10][5] ;
 wire \ppu.pal[10][6] ;
 wire \ppu.pal[10][7] ;
 wire \ppu.pal[11][0] ;
 wire \ppu.pal[11][1] ;
 wire \ppu.pal[11][2] ;
 wire \ppu.pal[11][3] ;
 wire \ppu.pal[11][4] ;
 wire \ppu.pal[11][5] ;
 wire \ppu.pal[11][6] ;
 wire \ppu.pal[11][7] ;
 wire \ppu.pal[12][0] ;
 wire \ppu.pal[12][1] ;
 wire \ppu.pal[12][2] ;
 wire \ppu.pal[12][3] ;
 wire \ppu.pal[12][4] ;
 wire \ppu.pal[12][5] ;
 wire \ppu.pal[12][6] ;
 wire \ppu.pal[12][7] ;
 wire \ppu.pal[13][0] ;
 wire \ppu.pal[13][1] ;
 wire \ppu.pal[13][2] ;
 wire \ppu.pal[13][3] ;
 wire \ppu.pal[13][4] ;
 wire \ppu.pal[13][5] ;
 wire \ppu.pal[13][6] ;
 wire \ppu.pal[13][7] ;
 wire \ppu.pal[14][0] ;
 wire \ppu.pal[14][1] ;
 wire \ppu.pal[14][2] ;
 wire \ppu.pal[14][3] ;
 wire \ppu.pal[14][4] ;
 wire \ppu.pal[14][5] ;
 wire \ppu.pal[14][6] ;
 wire \ppu.pal[14][7] ;
 wire \ppu.pal[15][0] ;
 wire \ppu.pal[15][1] ;
 wire \ppu.pal[15][2] ;
 wire \ppu.pal[15][3] ;
 wire \ppu.pal[15][4] ;
 wire \ppu.pal[15][5] ;
 wire \ppu.pal[15][6] ;
 wire \ppu.pal[15][7] ;
 wire \ppu.pal[1][0] ;
 wire \ppu.pal[1][1] ;
 wire \ppu.pal[1][2] ;
 wire \ppu.pal[1][3] ;
 wire \ppu.pal[1][4] ;
 wire \ppu.pal[1][5] ;
 wire \ppu.pal[1][6] ;
 wire \ppu.pal[1][7] ;
 wire \ppu.pal[2][0] ;
 wire \ppu.pal[2][1] ;
 wire \ppu.pal[2][2] ;
 wire \ppu.pal[2][3] ;
 wire \ppu.pal[2][4] ;
 wire \ppu.pal[2][5] ;
 wire \ppu.pal[2][6] ;
 wire \ppu.pal[2][7] ;
 wire \ppu.pal[3][0] ;
 wire \ppu.pal[3][1] ;
 wire \ppu.pal[3][2] ;
 wire \ppu.pal[3][3] ;
 wire \ppu.pal[3][4] ;
 wire \ppu.pal[3][5] ;
 wire \ppu.pal[3][6] ;
 wire \ppu.pal[3][7] ;
 wire \ppu.pal[4][0] ;
 wire \ppu.pal[4][1] ;
 wire \ppu.pal[4][2] ;
 wire \ppu.pal[4][3] ;
 wire \ppu.pal[4][4] ;
 wire \ppu.pal[4][5] ;
 wire \ppu.pal[4][6] ;
 wire \ppu.pal[4][7] ;
 wire \ppu.pal[5][0] ;
 wire \ppu.pal[5][1] ;
 wire \ppu.pal[5][2] ;
 wire \ppu.pal[5][3] ;
 wire \ppu.pal[5][4] ;
 wire \ppu.pal[5][5] ;
 wire \ppu.pal[5][6] ;
 wire \ppu.pal[5][7] ;
 wire \ppu.pal[6][0] ;
 wire \ppu.pal[6][1] ;
 wire \ppu.pal[6][2] ;
 wire \ppu.pal[6][3] ;
 wire \ppu.pal[6][4] ;
 wire \ppu.pal[6][5] ;
 wire \ppu.pal[6][6] ;
 wire \ppu.pal[6][7] ;
 wire \ppu.pal[7][0] ;
 wire \ppu.pal[7][1] ;
 wire \ppu.pal[7][2] ;
 wire \ppu.pal[7][3] ;
 wire \ppu.pal[7][4] ;
 wire \ppu.pal[7][5] ;
 wire \ppu.pal[7][6] ;
 wire \ppu.pal[7][7] ;
 wire \ppu.pal[8][0] ;
 wire \ppu.pal[8][1] ;
 wire \ppu.pal[8][2] ;
 wire \ppu.pal[8][3] ;
 wire \ppu.pal[8][4] ;
 wire \ppu.pal[8][5] ;
 wire \ppu.pal[8][6] ;
 wire \ppu.pal[8][7] ;
 wire \ppu.pal[9][0] ;
 wire \ppu.pal[9][1] ;
 wire \ppu.pal[9][2] ;
 wire \ppu.pal[9][3] ;
 wire \ppu.pal[9][4] ;
 wire \ppu.pal[9][5] ;
 wire \ppu.pal[9][6] ;
 wire \ppu.pal[9][7] ;
 wire \ppu.pal_data_out[0] ;
 wire \ppu.pal_data_out[1] ;
 wire \ppu.pal_data_out[2] ;
 wire \ppu.pal_data_out[3] ;
 wire \ppu.pal_out[0] ;
 wire \ppu.pal_out[1] ;
 wire \ppu.pal_out[2] ;
 wire \ppu.pal_out[3] ;
 wire \ppu.pixel_out_s[0] ;
 wire \ppu.pixel_out_s[1] ;
 wire \ppu.pixel_out_s[2] ;
 wire \ppu.pixel_out_s[3] ;
 wire \ppu.pixel_out_t[0] ;
 wire \ppu.pixel_out_t[1] ;
 wire \ppu.pixel_out_t[2] ;
 wire \ppu.pixel_out_t[3] ;
 wire \ppu.ram_on ;
 wire \ppu.ram_running ;
 wire \ppu.rs2.phase_x ;
 wire \ppu.rs2.phase_y[0] ;
 wire \ppu.rs2.phase_y[1] ;
 wire \ppu.rs2.vsync0 ;
 wire \ppu.rs2.x0[5] ;
 wire \ppu.rs2.x0[6] ;
 wire \ppu.rs2.x0[7] ;
 wire \ppu.rs2.y_scan.counter[0] ;
 wire \ppu.rs2.y_scan.counter[1] ;
 wire \ppu.rs2.y_scan.counter[2] ;
 wire \ppu.rs2.y_scan.counter[3] ;
 wire \ppu.rs2.y_scan.counter[4] ;
 wire \ppu.rs2.y_scan.counter[5] ;
 wire \ppu.rs2.y_scan.counter[6] ;
 wire \ppu.rs2.y_scan.counter[7] ;
 wire \ppu.rs2.y_scan.counter[8] ;
 wire \ppu.scroll_regs[0][0] ;
 wire \ppu.scroll_regs[0][1] ;
 wire \ppu.scroll_regs[0][2] ;
 wire \ppu.scroll_regs[0][3] ;
 wire \ppu.scroll_regs[0][4] ;
 wire \ppu.scroll_regs[0][5] ;
 wire \ppu.scroll_regs[0][6] ;
 wire \ppu.scroll_regs[0][7] ;
 wire \ppu.scroll_regs[0][8] ;
 wire \ppu.scroll_regs[1][0] ;
 wire \ppu.scroll_regs[1][1] ;
 wire \ppu.scroll_regs[1][2] ;
 wire \ppu.scroll_regs[1][3] ;
 wire \ppu.scroll_regs[1][4] ;
 wire \ppu.scroll_regs[1][5] ;
 wire \ppu.scroll_regs[1][6] ;
 wire \ppu.scroll_regs[1][7] ;
 wire \ppu.scroll_regs[1][8] ;
 wire \ppu.scroll_regs[2][0] ;
 wire \ppu.scroll_regs[2][1] ;
 wire \ppu.scroll_regs[2][2] ;
 wire \ppu.scroll_regs[2][3] ;
 wire \ppu.scroll_regs[2][4] ;
 wire \ppu.scroll_regs[2][5] ;
 wire \ppu.scroll_regs[2][6] ;
 wire \ppu.scroll_regs[2][7] ;
 wire \ppu.scroll_regs[2][8] ;
 wire \ppu.scroll_regs[3][0] ;
 wire \ppu.scroll_regs[3][1] ;
 wire \ppu.scroll_regs[3][2] ;
 wire \ppu.scroll_regs[3][3] ;
 wire \ppu.scroll_regs[3][4] ;
 wire \ppu.scroll_regs[3][5] ;
 wire \ppu.scroll_regs[3][6] ;
 wire \ppu.scroll_regs[3][7] ;
 wire \ppu.scroll_regs[3][8] ;
 wire \ppu.sprite_buffer.attr_x[0][0] ;
 wire \ppu.sprite_buffer.attr_x[0][10] ;
 wire \ppu.sprite_buffer.attr_x[0][11] ;
 wire \ppu.sprite_buffer.attr_x[0][12] ;
 wire \ppu.sprite_buffer.attr_x[0][13] ;
 wire \ppu.sprite_buffer.attr_x[0][14] ;
 wire \ppu.sprite_buffer.attr_x[0][15] ;
 wire \ppu.sprite_buffer.attr_x[0][1] ;
 wire \ppu.sprite_buffer.attr_x[0][2] ;
 wire \ppu.sprite_buffer.attr_x[0][3] ;
 wire \ppu.sprite_buffer.attr_x[0][4] ;
 wire \ppu.sprite_buffer.attr_x[0][5] ;
 wire \ppu.sprite_buffer.attr_x[0][6] ;
 wire \ppu.sprite_buffer.attr_x[0][7] ;
 wire \ppu.sprite_buffer.attr_x[0][8] ;
 wire \ppu.sprite_buffer.attr_x[0][9] ;
 wire \ppu.sprite_buffer.attr_x[1][0] ;
 wire \ppu.sprite_buffer.attr_x[1][10] ;
 wire \ppu.sprite_buffer.attr_x[1][11] ;
 wire \ppu.sprite_buffer.attr_x[1][12] ;
 wire \ppu.sprite_buffer.attr_x[1][13] ;
 wire \ppu.sprite_buffer.attr_x[1][14] ;
 wire \ppu.sprite_buffer.attr_x[1][15] ;
 wire \ppu.sprite_buffer.attr_x[1][1] ;
 wire \ppu.sprite_buffer.attr_x[1][2] ;
 wire \ppu.sprite_buffer.attr_x[1][3] ;
 wire \ppu.sprite_buffer.attr_x[1][4] ;
 wire \ppu.sprite_buffer.attr_x[1][5] ;
 wire \ppu.sprite_buffer.attr_x[1][6] ;
 wire \ppu.sprite_buffer.attr_x[1][7] ;
 wire \ppu.sprite_buffer.attr_x[1][8] ;
 wire \ppu.sprite_buffer.attr_x[1][9] ;
 wire \ppu.sprite_buffer.attr_x[2][0] ;
 wire \ppu.sprite_buffer.attr_x[2][10] ;
 wire \ppu.sprite_buffer.attr_x[2][11] ;
 wire \ppu.sprite_buffer.attr_x[2][12] ;
 wire \ppu.sprite_buffer.attr_x[2][13] ;
 wire \ppu.sprite_buffer.attr_x[2][14] ;
 wire \ppu.sprite_buffer.attr_x[2][15] ;
 wire \ppu.sprite_buffer.attr_x[2][1] ;
 wire \ppu.sprite_buffer.attr_x[2][2] ;
 wire \ppu.sprite_buffer.attr_x[2][3] ;
 wire \ppu.sprite_buffer.attr_x[2][4] ;
 wire \ppu.sprite_buffer.attr_x[2][5] ;
 wire \ppu.sprite_buffer.attr_x[2][6] ;
 wire \ppu.sprite_buffer.attr_x[2][7] ;
 wire \ppu.sprite_buffer.attr_x[2][8] ;
 wire \ppu.sprite_buffer.attr_x[2][9] ;
 wire \ppu.sprite_buffer.attr_x[3][0] ;
 wire \ppu.sprite_buffer.attr_x[3][10] ;
 wire \ppu.sprite_buffer.attr_x[3][11] ;
 wire \ppu.sprite_buffer.attr_x[3][12] ;
 wire \ppu.sprite_buffer.attr_x[3][13] ;
 wire \ppu.sprite_buffer.attr_x[3][14] ;
 wire \ppu.sprite_buffer.attr_x[3][15] ;
 wire \ppu.sprite_buffer.attr_x[3][1] ;
 wire \ppu.sprite_buffer.attr_x[3][2] ;
 wire \ppu.sprite_buffer.attr_x[3][3] ;
 wire \ppu.sprite_buffer.attr_x[3][4] ;
 wire \ppu.sprite_buffer.attr_x[3][5] ;
 wire \ppu.sprite_buffer.attr_x[3][6] ;
 wire \ppu.sprite_buffer.attr_x[3][7] ;
 wire \ppu.sprite_buffer.attr_x[3][8] ;
 wire \ppu.sprite_buffer.attr_x[3][9] ;
 wire \ppu.sprite_buffer.attr_y[0][0] ;
 wire \ppu.sprite_buffer.attr_y[0][10] ;
 wire \ppu.sprite_buffer.attr_y[0][11] ;
 wire \ppu.sprite_buffer.attr_y[0][12] ;
 wire \ppu.sprite_buffer.attr_y[0][13] ;
 wire \ppu.sprite_buffer.attr_y[0][14] ;
 wire \ppu.sprite_buffer.attr_y[0][15] ;
 wire \ppu.sprite_buffer.attr_y[0][1] ;
 wire \ppu.sprite_buffer.attr_y[0][2] ;
 wire \ppu.sprite_buffer.attr_y[0][4] ;
 wire \ppu.sprite_buffer.attr_y[0][5] ;
 wire \ppu.sprite_buffer.attr_y[0][6] ;
 wire \ppu.sprite_buffer.attr_y[0][7] ;
 wire \ppu.sprite_buffer.attr_y[0][8] ;
 wire \ppu.sprite_buffer.attr_y[0][9] ;
 wire \ppu.sprite_buffer.attr_y[1][0] ;
 wire \ppu.sprite_buffer.attr_y[1][10] ;
 wire \ppu.sprite_buffer.attr_y[1][11] ;
 wire \ppu.sprite_buffer.attr_y[1][12] ;
 wire \ppu.sprite_buffer.attr_y[1][13] ;
 wire \ppu.sprite_buffer.attr_y[1][14] ;
 wire \ppu.sprite_buffer.attr_y[1][15] ;
 wire \ppu.sprite_buffer.attr_y[1][1] ;
 wire \ppu.sprite_buffer.attr_y[1][2] ;
 wire \ppu.sprite_buffer.attr_y[1][4] ;
 wire \ppu.sprite_buffer.attr_y[1][5] ;
 wire \ppu.sprite_buffer.attr_y[1][6] ;
 wire \ppu.sprite_buffer.attr_y[1][7] ;
 wire \ppu.sprite_buffer.attr_y[1][8] ;
 wire \ppu.sprite_buffer.attr_y[1][9] ;
 wire \ppu.sprite_buffer.data8[0] ;
 wire \ppu.sprite_buffer.data8[1] ;
 wire \ppu.sprite_buffer.data8[2] ;
 wire \ppu.sprite_buffer.data8[3] ;
 wire \ppu.sprite_buffer.extra_sorted_addr_bits[0] ;
 wire \ppu.sprite_buffer.extra_sorted_addr_bits[1] ;
 wire \ppu.sprite_buffer.extra_sorted_addr_bits[2] ;
 wire \ppu.sprite_buffer.final_pixels_in ;
 wire \ppu.sprite_buffer.id_buffer[0][0] ;
 wire \ppu.sprite_buffer.id_buffer[0][1] ;
 wire \ppu.sprite_buffer.id_buffer[0][2] ;
 wire \ppu.sprite_buffer.id_buffer[0][3] ;
 wire \ppu.sprite_buffer.id_buffer[0][4] ;
 wire \ppu.sprite_buffer.id_buffer[0][5] ;
 wire \ppu.sprite_buffer.id_buffer[1][0] ;
 wire \ppu.sprite_buffer.id_buffer[1][1] ;
 wire \ppu.sprite_buffer.id_buffer[1][2] ;
 wire \ppu.sprite_buffer.id_buffer[1][3] ;
 wire \ppu.sprite_buffer.id_buffer[1][4] ;
 wire \ppu.sprite_buffer.id_buffer[1][5] ;
 wire \ppu.sprite_buffer.id_buffer[2][0] ;
 wire \ppu.sprite_buffer.id_buffer[2][1] ;
 wire \ppu.sprite_buffer.id_buffer[2][2] ;
 wire \ppu.sprite_buffer.id_buffer[2][3] ;
 wire \ppu.sprite_buffer.id_buffer[2][4] ;
 wire \ppu.sprite_buffer.id_buffer[2][5] ;
 wire \ppu.sprite_buffer.id_buffer[3][0] ;
 wire \ppu.sprite_buffer.id_buffer[3][1] ;
 wire \ppu.sprite_buffer.id_buffer[3][2] ;
 wire \ppu.sprite_buffer.id_buffer[3][3] ;
 wire \ppu.sprite_buffer.id_buffer[3][4] ;
 wire \ppu.sprite_buffer.id_buffer[3][5] ;
 wire \ppu.sprite_buffer.in_counter_idy[0] ;
 wire \ppu.sprite_buffer.in_counter_idy[1] ;
 wire \ppu.sprite_buffer.in_counters[1][0] ;
 wire \ppu.sprite_buffer.in_counters[1][1] ;
 wire \ppu.sprite_buffer.in_counters[1][2] ;
 wire \ppu.sprite_buffer.in_counters[2][1] ;
 wire \ppu.sprite_buffer.in_counters[2][2] ;
 wire \ppu.sprite_buffer.oam_load_sprite_valid ;
 wire \ppu.sprite_buffer.oam_req_step ;
 wire \ppu.sprite_buffer.out_counter_oam[0] ;
 wire \ppu.sprite_buffer.out_counter_oam[1] ;
 wire \ppu.sprite_buffer.out_counters[0][0] ;
 wire \ppu.sprite_buffer.out_counters[0][1] ;
 wire \ppu.sprite_buffer.out_counters[0][2] ;
 wire \ppu.sprite_buffer.out_counters[2][0] ;
 wire \ppu.sprite_buffer.out_counters[2][1] ;
 wire \ppu.sprite_buffer.out_counters[2][2] ;
 wire \ppu.sprite_buffer.scan_enabled ;
 wire \ppu.sprite_buffer.scan_on ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[0][0] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[0][1] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[0][2] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[1][0] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[1][1] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[1][2] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[2][0] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[2][1] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[2][2] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[3][0] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[3][1] ;
 wire \ppu.sprite_buffer.sprite_catch_up_counters[3][2] ;
 wire \ppu.sprite_buffer.sprite_ids[0][0] ;
 wire \ppu.sprite_buffer.sprite_ids[0][1] ;
 wire \ppu.sprite_buffer.sprite_ids[0][2] ;
 wire \ppu.sprite_buffer.sprite_ids[0][3] ;
 wire \ppu.sprite_buffer.sprite_ids[0][4] ;
 wire \ppu.sprite_buffer.sprite_ids[0][5] ;
 wire \ppu.sprite_buffer.sprite_ids[1][0] ;
 wire \ppu.sprite_buffer.sprite_ids[1][1] ;
 wire \ppu.sprite_buffer.sprite_ids[1][2] ;
 wire \ppu.sprite_buffer.sprite_ids[1][3] ;
 wire \ppu.sprite_buffer.sprite_ids[1][4] ;
 wire \ppu.sprite_buffer.sprite_ids[1][5] ;
 wire \ppu.sprite_buffer.sprite_ids[2][0] ;
 wire \ppu.sprite_buffer.sprite_ids[2][1] ;
 wire \ppu.sprite_buffer.sprite_ids[2][2] ;
 wire \ppu.sprite_buffer.sprite_ids[2][3] ;
 wire \ppu.sprite_buffer.sprite_ids[2][4] ;
 wire \ppu.sprite_buffer.sprite_ids[2][5] ;
 wire \ppu.sprite_buffer.sprite_ids[3][0] ;
 wire \ppu.sprite_buffer.sprite_ids[3][1] ;
 wire \ppu.sprite_buffer.sprite_ids[3][2] ;
 wire \ppu.sprite_buffer.sprite_ids[3][3] ;
 wire \ppu.sprite_buffer.sprite_ids[3][4] ;
 wire \ppu.sprite_buffer.sprite_ids[3][5] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][0] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][10] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][11] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][12] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][13] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][14] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][15] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][16] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][17] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][18] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][19] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][1] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][20] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][21] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][22] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][23] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][24] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][25] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][26] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][27] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][28] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][29] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][2] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][30] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][31] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][3] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][4] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][5] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][6] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][7] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][8] ;
 wire \ppu.sprite_buffer.sprite_pixels[0][9] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][0] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][10] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][11] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][12] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][13] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][14] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][15] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][16] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][17] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][18] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][19] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][1] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][20] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][21] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][22] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][23] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][24] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][25] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][26] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][27] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][28] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][29] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][2] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][30] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][31] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][3] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][4] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][5] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][6] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][7] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][8] ;
 wire \ppu.sprite_buffer.sprite_pixels[1][9] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][0] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][10] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][11] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][12] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][13] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][14] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][15] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][16] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][17] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][18] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][19] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][1] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][20] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][21] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][22] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][23] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][24] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][25] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][26] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][27] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][28] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][29] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][2] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][30] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][31] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][3] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][4] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][5] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][6] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][7] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][8] ;
 wire \ppu.sprite_buffer.sprite_pixels[2][9] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][0] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][10] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][11] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][12] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][13] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][14] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][15] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][16] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][17] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][18] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][19] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][1] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][20] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][21] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][22] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][23] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][24] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][25] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][26] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][27] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][28] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][29] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][2] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][30] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][31] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][3] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][4] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][5] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][6] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][7] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][8] ;
 wire \ppu.sprite_buffer.sprite_pixels[3][9] ;
 wire \ppu.sprite_buffer.top_color[0] ;
 wire \ppu.sprite_buffer.top_color[1] ;
 wire \ppu.sprite_buffer.top_color[2] ;
 wire \ppu.sprite_buffer.top_color[3] ;
 wire \ppu.sprite_buffer.top_depth[0] ;
 wire \ppu.sprite_buffer.top_depth[1] ;
 wire \ppu.sprite_buffer.top_prio[0] ;
 wire \ppu.sprite_buffer.top_prio[1] ;
 wire \ppu.sprite_buffer.top_prio[2] ;
 wire \ppu.sprite_buffer.top_prio[3] ;
 wire \ppu.sprite_buffer.top_prio[4] ;
 wire \ppu.sprite_buffer.top_prio[5] ;
 wire \ppu.sprite_buffer.top_prio[6] ;
 wire \ppu.sprite_buffer.valid_sprites[0] ;
 wire \ppu.sprite_buffer.valid_sprites[1] ;
 wire \ppu.sprite_buffer.valid_sprites[2] ;
 wire \ppu.sprite_buffer.valid_sprites[3] ;
 wire \ppu.sprite_buffer.y_matched0 ;
 wire \ppu.sync_delay[0] ;
 wire \ppu.sync_delay[1] ;
 wire \ppu.sync_delay[2] ;
 wire \ppu.tilemap.attr[0][0] ;
 wire \ppu.tilemap.attr[0][1] ;
 wire \ppu.tilemap.attr[0][2] ;
 wire \ppu.tilemap.attr[0][3] ;
 wire \ppu.tilemap.attr[0][4] ;
 wire \ppu.tilemap.attr[1][0] ;
 wire \ppu.tilemap.attr[1][1] ;
 wire \ppu.tilemap.attr[1][2] ;
 wire \ppu.tilemap.attr[1][3] ;
 wire \ppu.tilemap.attr[1][4] ;
 wire \ppu.tilemap.map_pixels[0][0] ;
 wire \ppu.tilemap.map_pixels[0][10] ;
 wire \ppu.tilemap.map_pixels[0][11] ;
 wire \ppu.tilemap.map_pixels[0][12] ;
 wire \ppu.tilemap.map_pixels[0][13] ;
 wire \ppu.tilemap.map_pixels[0][14] ;
 wire \ppu.tilemap.map_pixels[0][15] ;
 wire \ppu.tilemap.map_pixels[0][1] ;
 wire \ppu.tilemap.map_pixels[0][2] ;
 wire \ppu.tilemap.map_pixels[0][3] ;
 wire \ppu.tilemap.map_pixels[0][4] ;
 wire \ppu.tilemap.map_pixels[0][5] ;
 wire \ppu.tilemap.map_pixels[0][6] ;
 wire \ppu.tilemap.map_pixels[0][7] ;
 wire \ppu.tilemap.map_pixels[0][8] ;
 wire \ppu.tilemap.map_pixels[0][9] ;
 wire \ppu.tilemap.map_pixels[1][0] ;
 wire \ppu.tilemap.map_pixels[1][10] ;
 wire \ppu.tilemap.map_pixels[1][11] ;
 wire \ppu.tilemap.map_pixels[1][12] ;
 wire \ppu.tilemap.map_pixels[1][13] ;
 wire \ppu.tilemap.map_pixels[1][14] ;
 wire \ppu.tilemap.map_pixels[1][15] ;
 wire \ppu.tilemap.map_pixels[1][1] ;
 wire \ppu.tilemap.map_pixels[1][2] ;
 wire \ppu.tilemap.map_pixels[1][3] ;
 wire \ppu.tilemap.map_pixels[1][4] ;
 wire \ppu.tilemap.map_pixels[1][5] ;
 wire \ppu.tilemap.map_pixels[1][6] ;
 wire \ppu.tilemap.map_pixels[1][7] ;
 wire \ppu.tilemap.map_pixels[1][8] ;
 wire \ppu.tilemap.map_pixels[1][9] ;
 wire \ppu.tilemap.next_attr[0][0] ;
 wire \ppu.tilemap.next_attr[0][1] ;
 wire \ppu.tilemap.next_attr[0][2] ;
 wire \ppu.tilemap.next_attr[0][3] ;
 wire \ppu.tilemap.next_attr[0][4] ;
 wire \ppu.tilemap.next_attr[1][0] ;
 wire \ppu.tilemap.next_attr[1][1] ;
 wire \ppu.tilemap.next_attr[1][2] ;
 wire \ppu.tilemap.next_attr[1][3] ;
 wire \ppu.tilemap.next_attr[1][4] ;
 wire \ppu.vsync ;
 wire \ppu_ctrl[0] ;
 wire \ppu_ctrl[2] ;
 wire \ppu_ctrl[4] ;
 wire reset;
 wire \rx_in_reg[0] ;
 wire \rx_in_reg[1] ;
 wire \synth.controller.counter[0] ;
 wire \synth.controller.counter[1] ;
 wire \synth.controller.counter[2] ;
 wire \synth.controller.counter[3] ;
 wire \synth.controller.curr_voice[0] ;
 wire \synth.controller.curr_voice[1] ;
 wire \synth.controller.ext_tx_request ;
 wire \synth.controller.out[0] ;
 wire \synth.controller.out[10] ;
 wire \synth.controller.out[11] ;
 wire \synth.controller.out[12] ;
 wire \synth.controller.out[13] ;
 wire \synth.controller.out[14] ;
 wire \synth.controller.out[15] ;
 wire \synth.controller.out[1] ;
 wire \synth.controller.out[2] ;
 wire \synth.controller.out[3] ;
 wire \synth.controller.out[4] ;
 wire \synth.controller.out[5] ;
 wire \synth.controller.out[6] ;
 wire \synth.controller.out[7] ;
 wire \synth.controller.out[8] ;
 wire \synth.controller.out[9] ;
 wire \synth.controller.out_reg[0] ;
 wire \synth.controller.out_reg[10] ;
 wire \synth.controller.out_reg[11] ;
 wire \synth.controller.out_reg[12] ;
 wire \synth.controller.out_reg[13] ;
 wire \synth.controller.out_reg[14] ;
 wire \synth.controller.out_reg[15] ;
 wire \synth.controller.out_reg[1] ;
 wire \synth.controller.out_reg[2] ;
 wire \synth.controller.out_reg[3] ;
 wire \synth.controller.out_reg[4] ;
 wire \synth.controller.out_reg[5] ;
 wire \synth.controller.out_reg[6] ;
 wire \synth.controller.out_reg[7] ;
 wire \synth.controller.out_reg[8] ;
 wire \synth.controller.out_reg[9] ;
 wire \synth.controller.out_reg_valid ;
 wire \synth.controller.out_valid ;
 wire \synth.controller.read_index_reg[0] ;
 wire \synth.controller.read_index_reg[1] ;
 wire \synth.controller.read_index_reg[2] ;
 wire \synth.controller.read_index_reg[3] ;
 wire \synth.controller.reg_waddr[0] ;
 wire \synth.controller.reg_waddr[1] ;
 wire \synth.controller.reg_waddr[2] ;
 wire \synth.controller.reg_waddr[3] ;
 wire \synth.controller.reg_wdata[0] ;
 wire \synth.controller.reg_wdata[1] ;
 wire \synth.controller.reg_wdata[2] ;
 wire \synth.controller.reg_wdata[3] ;
 wire \synth.controller.reg_wdata[4] ;
 wire \synth.controller.reg_wdata[5] ;
 wire \synth.controller.reg_wdata[6] ;
 wire \synth.controller.reg_wdata[7] ;
 wire \synth.controller.rx_buffer[12] ;
 wire \synth.controller.rx_buffer[13] ;
 wire \synth.controller.rx_buffer[14] ;
 wire \synth.controller.rx_buffer[15] ;
 wire \synth.controller.rx_buffer_valid ;
 wire \synth.controller.rx_counter[0] ;
 wire \synth.controller.rx_counter[1] ;
 wire \synth.controller.rx_counter[2] ;
 wire \synth.controller.rx_counter[3] ;
 wire \synth.controller.rx_sbs[0] ;
 wire \synth.controller.rx_sbs[1] ;
 wire \synth.controller.sample_counter[0] ;
 wire \synth.controller.sample_counter[1] ;
 wire \synth.controller.sample_credits[0] ;
 wire \synth.controller.sample_credits[1] ;
 wire \synth.controller.sbio_credits[0] ;
 wire \synth.controller.sbio_credits[1] ;
 wire \synth.controller.sbio_credits[2] ;
 wire \synth.controller.sbio_tx.counter[0] ;
 wire \synth.controller.sbio_tx.counter[1] ;
 wire \synth.controller.sbio_tx.counter[2] ;
 wire \synth.controller.sbio_tx.counter[3] ;
 wire \synth.controller.sbio_tx.start_present ;
 wire \synth.controller.scanning_out ;
 wire \synth.controller.step_sample ;
 wire \synth.controller.sweep_addr_index[0] ;
 wire \synth.controller.sweep_addr_index[1] ;
 wire \synth.controller.sweep_addr_index[2] ;
 wire \synth.controller.sweep_data_index[0] ;
 wire \synth.controller.sweep_data_index[1] ;
 wire \synth.controller.sweep_data_index[2] ;
 wire \synth.controller.tap_pos[0] ;
 wire \synth.controller.tap_pos[1] ;
 wire \synth.controller.tx_outstanding[0] ;
 wire \synth.controller.tx_outstanding[1] ;
 wire \synth.controller.tx_outstanding[2] ;
 wire \synth.controller.tx_source[0] ;
 wire \synth.controller.tx_source[1] ;
 wire \synth.controller.write_index_reg[0] ;
 wire \synth.controller.write_index_reg[1] ;
 wire \synth.controller.write_index_reg[2] ;
 wire \synth.controller.write_index_reg[3] ;
 wire \synth.voice.a_sel_reg[1] ;
 wire \synth.voice.a_sel_reg[2] ;
 wire \synth.voice.a_sel_reg[3] ;
 wire \synth.voice.acc[0] ;
 wire \synth.voice.acc[1] ;
 wire \synth.voice.acc[2] ;
 wire \synth.voice.acc[3] ;
 wire \synth.voice.accs[1][0] ;
 wire \synth.voice.accs[1][10] ;
 wire \synth.voice.accs[1][11] ;
 wire \synth.voice.accs[1][12] ;
 wire \synth.voice.accs[1][13] ;
 wire \synth.voice.accs[1][14] ;
 wire \synth.voice.accs[1][15] ;
 wire \synth.voice.accs[1][16] ;
 wire \synth.voice.accs[1][17] ;
 wire \synth.voice.accs[1][18] ;
 wire \synth.voice.accs[1][19] ;
 wire \synth.voice.accs[1][1] ;
 wire \synth.voice.accs[1][2] ;
 wire \synth.voice.accs[1][3] ;
 wire \synth.voice.accs[1][4] ;
 wire \synth.voice.accs[1][5] ;
 wire \synth.voice.accs[1][6] ;
 wire \synth.voice.accs[1][7] ;
 wire \synth.voice.accs[1][8] ;
 wire \synth.voice.accs[1][9] ;
 wire \synth.voice.accs[2][0] ;
 wire \synth.voice.accs[2][10] ;
 wire \synth.voice.accs[2][11] ;
 wire \synth.voice.accs[2][12] ;
 wire \synth.voice.accs[2][13] ;
 wire \synth.voice.accs[2][14] ;
 wire \synth.voice.accs[2][15] ;
 wire \synth.voice.accs[2][16] ;
 wire \synth.voice.accs[2][17] ;
 wire \synth.voice.accs[2][18] ;
 wire \synth.voice.accs[2][19] ;
 wire \synth.voice.accs[2][1] ;
 wire \synth.voice.accs[2][2] ;
 wire \synth.voice.accs[2][3] ;
 wire \synth.voice.accs[2][4] ;
 wire \synth.voice.accs[2][5] ;
 wire \synth.voice.accs[2][6] ;
 wire \synth.voice.accs[2][7] ;
 wire \synth.voice.accs[2][8] ;
 wire \synth.voice.accs[2][9] ;
 wire \synth.voice.accs[3][0] ;
 wire \synth.voice.accs[3][10] ;
 wire \synth.voice.accs[3][11] ;
 wire \synth.voice.accs[3][12] ;
 wire \synth.voice.accs[3][13] ;
 wire \synth.voice.accs[3][14] ;
 wire \synth.voice.accs[3][15] ;
 wire \synth.voice.accs[3][16] ;
 wire \synth.voice.accs[3][17] ;
 wire \synth.voice.accs[3][18] ;
 wire \synth.voice.accs[3][19] ;
 wire \synth.voice.accs[3][1] ;
 wire \synth.voice.accs[3][2] ;
 wire \synth.voice.accs[3][3] ;
 wire \synth.voice.accs[3][4] ;
 wire \synth.voice.accs[3][5] ;
 wire \synth.voice.accs[3][6] ;
 wire \synth.voice.accs[3][7] ;
 wire \synth.voice.accs[3][8] ;
 wire \synth.voice.accs[3][9] ;
 wire \synth.voice.accs[4][0] ;
 wire \synth.voice.accs[4][10] ;
 wire \synth.voice.accs[4][11] ;
 wire \synth.voice.accs[4][12] ;
 wire \synth.voice.accs[4][13] ;
 wire \synth.voice.accs[4][14] ;
 wire \synth.voice.accs[4][15] ;
 wire \synth.voice.accs[4][16] ;
 wire \synth.voice.accs[4][17] ;
 wire \synth.voice.accs[4][18] ;
 wire \synth.voice.accs[4][19] ;
 wire \synth.voice.accs[4][1] ;
 wire \synth.voice.accs[4][2] ;
 wire \synth.voice.accs[4][3] ;
 wire \synth.voice.accs[4][4] ;
 wire \synth.voice.accs[4][5] ;
 wire \synth.voice.accs[4][6] ;
 wire \synth.voice.accs[4][7] ;
 wire \synth.voice.accs[4][8] ;
 wire \synth.voice.accs[4][9] ;
 wire \synth.voice.accs[5][0] ;
 wire \synth.voice.accs[5][10] ;
 wire \synth.voice.accs[5][11] ;
 wire \synth.voice.accs[5][12] ;
 wire \synth.voice.accs[5][13] ;
 wire \synth.voice.accs[5][14] ;
 wire \synth.voice.accs[5][15] ;
 wire \synth.voice.accs[5][16] ;
 wire \synth.voice.accs[5][17] ;
 wire \synth.voice.accs[5][18] ;
 wire \synth.voice.accs[5][19] ;
 wire \synth.voice.accs[5][1] ;
 wire \synth.voice.accs[5][2] ;
 wire \synth.voice.accs[5][3] ;
 wire \synth.voice.accs[5][4] ;
 wire \synth.voice.accs[5][5] ;
 wire \synth.voice.accs[5][6] ;
 wire \synth.voice.accs[5][7] ;
 wire \synth.voice.accs[5][8] ;
 wire \synth.voice.accs[5][9] ;
 wire \synth.voice.b_sel_reg[0] ;
 wire \synth.voice.b_sel_reg[2] ;
 wire \synth.voice.bpf_en[0] ;
 wire \synth.voice.bpf_en[1] ;
 wire \synth.voice.bpf_en[2] ;
 wire \synth.voice.coeff_index[0] ;
 wire \synth.voice.coeff_index[1] ;
 wire \synth.voice.coeff_index[2] ;
 wire \synth.voice.coeff_index[3] ;
 wire \synth.voice.coeff_index[4] ;
 wire \synth.voice.delayed_p[0] ;
 wire \synth.voice.delayed_p[1] ;
 wire \synth.voice.delayed_s ;
 wire \synth.voice.fir_table.exp[0] ;
 wire \synth.voice.fir_table.exp[1] ;
 wire \synth.voice.fir_table.exp[2] ;
 wire \synth.voice.fir_table.exp[3] ;
 wire \synth.voice.fir_table.i_term[0] ;
 wire \synth.voice.fir_table.i_term[1] ;
 wire \synth.voice.fir_table.i_term[2] ;
 wire \synth.voice.fir_table.sign ;
 wire \synth.voice.flip_sign ;
 wire \synth.voice.flip_sign_fir ;
 wire \synth.voice.flip_sign_reg ;
 wire \synth.voice.float_period[0][0] ;
 wire \synth.voice.float_period[0][10] ;
 wire \synth.voice.float_period[0][11] ;
 wire \synth.voice.float_period[0][12] ;
 wire \synth.voice.float_period[0][13] ;
 wire \synth.voice.float_period[0][1] ;
 wire \synth.voice.float_period[0][2] ;
 wire \synth.voice.float_period[0][3] ;
 wire \synth.voice.float_period[0][4] ;
 wire \synth.voice.float_period[0][5] ;
 wire \synth.voice.float_period[0][6] ;
 wire \synth.voice.float_period[0][7] ;
 wire \synth.voice.float_period[0][8] ;
 wire \synth.voice.float_period[0][9] ;
 wire \synth.voice.float_period[1][0] ;
 wire \synth.voice.float_period[1][10] ;
 wire \synth.voice.float_period[1][11] ;
 wire \synth.voice.float_period[1][12] ;
 wire \synth.voice.float_period[1][13] ;
 wire \synth.voice.float_period[1][1] ;
 wire \synth.voice.float_period[1][2] ;
 wire \synth.voice.float_period[1][3] ;
 wire \synth.voice.float_period[1][4] ;
 wire \synth.voice.float_period[1][5] ;
 wire \synth.voice.float_period[1][6] ;
 wire \synth.voice.float_period[1][7] ;
 wire \synth.voice.float_period[1][8] ;
 wire \synth.voice.float_period[1][9] ;
 wire \synth.voice.genblk4[0].next_state_scan[10] ;
 wire \synth.voice.genblk4[0].next_state_scan[11] ;
 wire \synth.voice.genblk4[0].next_state_scan[12] ;
 wire \synth.voice.genblk4[0].next_state_scan[13] ;
 wire \synth.voice.genblk4[0].next_state_scan[4] ;
 wire \synth.voice.genblk4[0].next_state_scan[5] ;
 wire \synth.voice.genblk4[0].next_state_scan[6] ;
 wire \synth.voice.genblk4[0].next_state_scan[7] ;
 wire \synth.voice.genblk4[0].next_state_scan[8] ;
 wire \synth.voice.genblk4[0].next_state_scan[9] ;
 wire \synth.voice.genblk4[10].next_state_scan[0] ;
 wire \synth.voice.genblk4[10].next_state_scan[10] ;
 wire \synth.voice.genblk4[10].next_state_scan[11] ;
 wire \synth.voice.genblk4[10].next_state_scan[12] ;
 wire \synth.voice.genblk4[10].next_state_scan[13] ;
 wire \synth.voice.genblk4[10].next_state_scan[1] ;
 wire \synth.voice.genblk4[10].next_state_scan[2] ;
 wire \synth.voice.genblk4[10].next_state_scan[3] ;
 wire \synth.voice.genblk4[10].next_state_scan[4] ;
 wire \synth.voice.genblk4[10].next_state_scan[5] ;
 wire \synth.voice.genblk4[10].next_state_scan[6] ;
 wire \synth.voice.genblk4[10].next_state_scan[7] ;
 wire \synth.voice.genblk4[10].next_state_scan[8] ;
 wire \synth.voice.genblk4[10].next_state_scan[9] ;
 wire \synth.voice.genblk4[11].next_state_scan[10] ;
 wire \synth.voice.genblk4[11].next_state_scan[11] ;
 wire \synth.voice.genblk4[11].next_state_scan[12] ;
 wire \synth.voice.genblk4[11].next_state_scan[13] ;
 wire \synth.voice.genblk4[11].next_state_scan[3] ;
 wire \synth.voice.genblk4[11].next_state_scan[4] ;
 wire \synth.voice.genblk4[11].next_state_scan[5] ;
 wire \synth.voice.genblk4[11].next_state_scan[6] ;
 wire \synth.voice.genblk4[11].next_state_scan[7] ;
 wire \synth.voice.genblk4[11].next_state_scan[8] ;
 wire \synth.voice.genblk4[11].next_state_scan[9] ;
 wire \synth.voice.genblk4[1].next_state_scan[0] ;
 wire \synth.voice.genblk4[1].next_state_scan[10] ;
 wire \synth.voice.genblk4[1].next_state_scan[11] ;
 wire \synth.voice.genblk4[1].next_state_scan[12] ;
 wire \synth.voice.genblk4[1].next_state_scan[13] ;
 wire \synth.voice.genblk4[1].next_state_scan[1] ;
 wire \synth.voice.genblk4[1].next_state_scan[2] ;
 wire \synth.voice.genblk4[1].next_state_scan[3] ;
 wire \synth.voice.genblk4[1].next_state_scan[4] ;
 wire \synth.voice.genblk4[1].next_state_scan[5] ;
 wire \synth.voice.genblk4[1].next_state_scan[6] ;
 wire \synth.voice.genblk4[1].next_state_scan[7] ;
 wire \synth.voice.genblk4[1].next_state_scan[8] ;
 wire \synth.voice.genblk4[1].next_state_scan[9] ;
 wire \synth.voice.genblk4[2].next_state_scan[0] ;
 wire \synth.voice.genblk4[2].next_state_scan[10] ;
 wire \synth.voice.genblk4[2].next_state_scan[11] ;
 wire \synth.voice.genblk4[2].next_state_scan[12] ;
 wire \synth.voice.genblk4[2].next_state_scan[13] ;
 wire \synth.voice.genblk4[2].next_state_scan[1] ;
 wire \synth.voice.genblk4[2].next_state_scan[2] ;
 wire \synth.voice.genblk4[2].next_state_scan[3] ;
 wire \synth.voice.genblk4[2].next_state_scan[4] ;
 wire \synth.voice.genblk4[2].next_state_scan[5] ;
 wire \synth.voice.genblk4[2].next_state_scan[6] ;
 wire \synth.voice.genblk4[2].next_state_scan[7] ;
 wire \synth.voice.genblk4[2].next_state_scan[8] ;
 wire \synth.voice.genblk4[2].next_state_scan[9] ;
 wire \synth.voice.genblk4[3].next_state_scan[0] ;
 wire \synth.voice.genblk4[3].next_state_scan[10] ;
 wire \synth.voice.genblk4[3].next_state_scan[11] ;
 wire \synth.voice.genblk4[3].next_state_scan[12] ;
 wire \synth.voice.genblk4[3].next_state_scan[13] ;
 wire \synth.voice.genblk4[3].next_state_scan[1] ;
 wire \synth.voice.genblk4[3].next_state_scan[2] ;
 wire \synth.voice.genblk4[3].next_state_scan[3] ;
 wire \synth.voice.genblk4[3].next_state_scan[4] ;
 wire \synth.voice.genblk4[3].next_state_scan[5] ;
 wire \synth.voice.genblk4[3].next_state_scan[6] ;
 wire \synth.voice.genblk4[3].next_state_scan[7] ;
 wire \synth.voice.genblk4[3].next_state_scan[8] ;
 wire \synth.voice.genblk4[3].next_state_scan[9] ;
 wire \synth.voice.genblk4[4].next_state_scan[0] ;
 wire \synth.voice.genblk4[4].next_state_scan[1] ;
 wire \synth.voice.genblk4[4].next_state_scan[2] ;
 wire \synth.voice.genblk4[4].next_state_scan[3] ;
 wire \synth.voice.genblk4[4].next_state_scan[4] ;
 wire \synth.voice.genblk4[4].next_state_scan[5] ;
 wire \synth.voice.genblk4[6].next_state_scan[10] ;
 wire \synth.voice.genblk4[6].next_state_scan[11] ;
 wire \synth.voice.genblk4[6].next_state_scan[12] ;
 wire \synth.voice.genblk4[6].next_state_scan[13] ;
 wire \synth.voice.genblk4[6].next_state_scan[2] ;
 wire \synth.voice.genblk4[6].next_state_scan[3] ;
 wire \synth.voice.genblk4[6].next_state_scan[4] ;
 wire \synth.voice.genblk4[6].next_state_scan[5] ;
 wire \synth.voice.genblk4[6].next_state_scan[6] ;
 wire \synth.voice.genblk4[6].next_state_scan[7] ;
 wire \synth.voice.genblk4[6].next_state_scan[8] ;
 wire \synth.voice.genblk4[6].next_state_scan[9] ;
 wire \synth.voice.genblk4[7].next_state_scan[0] ;
 wire \synth.voice.genblk4[7].next_state_scan[10] ;
 wire \synth.voice.genblk4[7].next_state_scan[11] ;
 wire \synth.voice.genblk4[7].next_state_scan[12] ;
 wire \synth.voice.genblk4[7].next_state_scan[13] ;
 wire \synth.voice.genblk4[7].next_state_scan[1] ;
 wire \synth.voice.genblk4[7].next_state_scan[2] ;
 wire \synth.voice.genblk4[7].next_state_scan[3] ;
 wire \synth.voice.genblk4[7].next_state_scan[4] ;
 wire \synth.voice.genblk4[7].next_state_scan[5] ;
 wire \synth.voice.genblk4[7].next_state_scan[6] ;
 wire \synth.voice.genblk4[7].next_state_scan[7] ;
 wire \synth.voice.genblk4[7].next_state_scan[8] ;
 wire \synth.voice.genblk4[7].next_state_scan[9] ;
 wire \synth.voice.genblk4[8].next_state_scan[0] ;
 wire \synth.voice.genblk4[8].next_state_scan[10] ;
 wire \synth.voice.genblk4[8].next_state_scan[11] ;
 wire \synth.voice.genblk4[8].next_state_scan[12] ;
 wire \synth.voice.genblk4[8].next_state_scan[13] ;
 wire \synth.voice.genblk4[8].next_state_scan[1] ;
 wire \synth.voice.genblk4[8].next_state_scan[2] ;
 wire \synth.voice.genblk4[8].next_state_scan[3] ;
 wire \synth.voice.genblk4[8].next_state_scan[4] ;
 wire \synth.voice.genblk4[8].next_state_scan[5] ;
 wire \synth.voice.genblk4[8].next_state_scan[6] ;
 wire \synth.voice.genblk4[8].next_state_scan[7] ;
 wire \synth.voice.genblk4[8].next_state_scan[8] ;
 wire \synth.voice.genblk4[8].next_state_scan[9] ;
 wire \synth.voice.genblk4[9].next_state_scan[0] ;
 wire \synth.voice.genblk4[9].next_state_scan[10] ;
 wire \synth.voice.genblk4[9].next_state_scan[11] ;
 wire \synth.voice.genblk4[9].next_state_scan[12] ;
 wire \synth.voice.genblk4[9].next_state_scan[13] ;
 wire \synth.voice.genblk4[9].next_state_scan[1] ;
 wire \synth.voice.genblk4[9].next_state_scan[2] ;
 wire \synth.voice.genblk4[9].next_state_scan[3] ;
 wire \synth.voice.genblk4[9].next_state_scan[4] ;
 wire \synth.voice.genblk4[9].next_state_scan[5] ;
 wire \synth.voice.genblk4[9].next_state_scan[6] ;
 wire \synth.voice.genblk4[9].next_state_scan[7] ;
 wire \synth.voice.genblk4[9].next_state_scan[8] ;
 wire \synth.voice.genblk4[9].next_state_scan[9] ;
 wire \synth.voice.lfsr[0] ;
 wire \synth.voice.lfsr[1] ;
 wire \synth.voice.mods[1][2] ;
 wire \synth.voice.mods[1][3] ;
 wire \synth.voice.mods[2][8] ;
 wire \synth.voice.mods[2][9] ;
 wire \synth.voice.next_sweep_oct_counter[0] ;
 wire \synth.voice.oct_counter[0] ;
 wire \synth.voice.oct_counter[10] ;
 wire \synth.voice.oct_counter[1] ;
 wire \synth.voice.oct_counter[2] ;
 wire \synth.voice.oct_counter[3] ;
 wire \synth.voice.oct_counter[4] ;
 wire \synth.voice.oct_counter[5] ;
 wire \synth.voice.oct_counter[6] ;
 wire \synth.voice.oct_counter[7] ;
 wire \synth.voice.oct_counter[8] ;
 wire \synth.voice.oct_counter[9] ;
 wire \synth.voice.params[24] ;
 wire \synth.voice.params[25] ;
 wire \synth.voice.params[8] ;
 wire \synth.voice.params[9] ;
 wire \synth.voice.restart_acc ;
 wire \synth.voice.rshift[0] ;
 wire \synth.voice.rshift[1] ;
 wire \synth.voice.rshift[2] ;
 wire \synth.voice.rshift[3] ;
 wire \synth.voice.rshift_reg0[0] ;
 wire \synth.voice.rshift_reg0[1] ;
 wire \synth.voice.rshift_reg0[2] ;
 wire \synth.voice.rshift_reg0[3] ;
 wire \synth.voice.rshift_reg[0] ;
 wire \synth.voice.rshift_reg[1] ;
 wire \synth.voice.rshift_reg[2] ;
 wire \synth.voice.rshift_reg[3] ;
 wire \synth.voice.scan_accs ;
 wire \synth.voice.scan_accs_reg ;
 wire \synth.voice.scan_outs[11][0] ;
 wire \synth.voice.scan_outs[11][1] ;
 wire \synth.voice.scan_outs[2][0] ;
 wire \synth.voice.scan_outs[2][1] ;
 wire \synth.voice.scan_outs[3][0] ;
 wire \synth.voice.scan_outs[3][1] ;
 wire \synth.voice.scan_outs[4][0] ;
 wire \synth.voice.scan_outs[4][1] ;
 wire \synth.voice.sweep_oct_counter[0] ;
 wire \synth.voice.sweep_oct_counter[10] ;
 wire \synth.voice.sweep_oct_counter[11] ;
 wire \synth.voice.sweep_oct_counter[12] ;
 wire \synth.voice.sweep_oct_counter[13] ;
 wire \synth.voice.sweep_oct_counter[1] ;
 wire \synth.voice.sweep_oct_counter[2] ;
 wire \synth.voice.sweep_oct_counter[3] ;
 wire \synth.voice.sweep_oct_counter[4] ;
 wire \synth.voice.sweep_oct_counter[5] ;
 wire \synth.voice.sweep_oct_counter[6] ;
 wire \synth.voice.sweep_oct_counter[7] ;
 wire \synth.voice.sweep_oct_counter[8] ;
 wire \synth.voice.sweep_oct_counter[9] ;
 wire \synth.voice.target_reg[1] ;
 wire \synth.voice.target_reg[2] ;
 wire \synth.voice.target_reg[3] ;
 wire \synth.voice.wave_reg[0] ;
 wire \synth.voice.wave_reg[1] ;
 wire \synth.voice.wave_reg[2] ;
 wire \synth.voice.wave_reg[3] ;
 wire \synth.voice.wave_reg[4] ;
 wire \synth.voice.wave_reg[5] ;
 wire \synth.voice.wave_reg[6] ;
 wire \synth.voice.wave_reg[7] ;
 wire \synth.voice.wave_reg[8] ;
 wire \synth.voice.wave_reg[9] ;
 wire \synth.voice.zero_shifter_out ;
 wire \synth.voice.zero_shifter_out_reg ;
 wire \uio_out0[6] ;
 wire \uio_out0[7] ;
 wire \uo_out0[0] ;
 wire \uo_out0[1] ;
 wire \uo_out0[2] ;
 wire \uo_out0[4] ;
 wire \uo_out0[5] ;
 wire \uo_out0[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _09048_ (.A(\synth.voice.fir_table.i_term[0] ),
    .X(_01715_));
 sg13g2_buf_2 _09049_ (.A(\synth.voice.fir_table.i_term[1] ),
    .X(_01716_));
 sg13g2_nor2_1 _09050_ (.A(_01715_),
    .B(_01716_),
    .Y(_01717_));
 sg13g2_nand2_1 _09051_ (.Y(_01718_),
    .A(_01717_),
    .B(_00045_));
 sg13g2_inv_1 _09052_ (.Y(_01719_),
    .A(_01718_));
 sg13g2_inv_4 _09053_ (.A(\synth.controller.tap_pos[1] ),
    .Y(_01720_));
 sg13g2_nor2_1 _09054_ (.A(\synth.controller.tap_pos[0] ),
    .B(_01720_),
    .Y(_01721_));
 sg13g2_inv_1 _09055_ (.Y(_01722_),
    .A(_01721_));
 sg13g2_nand2_1 _09056_ (.Y(_01723_),
    .A(_01719_),
    .B(_01722_));
 sg13g2_buf_1 _09057_ (.A(\synth.controller.counter[3] ),
    .X(_01724_));
 sg13g2_buf_2 _09058_ (.A(\synth.controller.counter[2] ),
    .X(_01725_));
 sg13g2_nor2_2 _09059_ (.A(_01724_),
    .B(_01725_),
    .Y(_01726_));
 sg13g2_buf_8 _09060_ (.A(\synth.controller.counter[0] ),
    .X(_01727_));
 sg13g2_buf_2 _09061_ (.A(\synth.controller.counter[1] ),
    .X(_01728_));
 sg13g2_nor2_1 _09062_ (.A(_01727_),
    .B(_01728_),
    .Y(_01729_));
 sg13g2_buf_8 _09063_ (.A(_01729_),
    .X(_01730_));
 sg13g2_nand2_2 _09064_ (.Y(_01731_),
    .A(_01726_),
    .B(_01730_));
 sg13g2_inv_1 _09065_ (.Y(_01732_),
    .A(_01731_));
 sg13g2_inv_1 _09066_ (.Y(_01733_),
    .A(_01726_));
 sg13g2_inv_1 _09067_ (.Y(_01734_),
    .A(_01725_));
 sg13g2_inv_8 _09068_ (.Y(_01735_),
    .A(_01730_));
 sg13g2_nor3_2 _09069_ (.A(_01724_),
    .B(_01734_),
    .C(_01735_),
    .Y(_01736_));
 sg13g2_inv_1 _09070_ (.Y(_01737_),
    .A(_01736_));
 sg13g2_a22oi_1 _09071_ (.Y(_01738_),
    .B1(_01733_),
    .B2(_01737_),
    .A2(_01732_),
    .A1(_01723_));
 sg13g2_buf_1 _09072_ (.A(_01738_),
    .X(_01739_));
 sg13g2_inv_1 _09073_ (.Y(_01740_),
    .A(_01739_));
 sg13g2_inv_1 _09074_ (.Y(_01741_),
    .A(\synth.voice.bpf_en[1] ));
 sg13g2_inv_1 _09075_ (.Y(_01742_),
    .A(_01728_));
 sg13g2_a21oi_1 _09076_ (.A1(_01741_),
    .A2(_01727_),
    .Y(_01743_),
    .B1(_01742_));
 sg13g2_o21ai_1 _09077_ (.B1(_01743_),
    .Y(_01744_),
    .A1(_01727_),
    .A2(\synth.voice.bpf_en[0] ));
 sg13g2_buf_1 _09078_ (.A(_01730_),
    .X(_01745_));
 sg13g2_nand2_1 _09079_ (.Y(_01746_),
    .A(_01745_),
    .B(\synth.voice.bpf_en[2] ));
 sg13g2_a221oi_1 _09080_ (.B2(_01746_),
    .C1(_00046_),
    .B1(_01744_),
    .A1(_01732_),
    .Y(_01747_),
    .A2(_01719_));
 sg13g2_nor2_1 _09081_ (.A(_01718_),
    .B(_01731_),
    .Y(_01748_));
 sg13g2_buf_8 _09082_ (.A(_01748_),
    .X(_01749_));
 sg13g2_inv_1 _09083_ (.Y(_01750_),
    .A(\synth.controller.tap_pos[0] ));
 sg13g2_nor2_1 _09084_ (.A(\synth.controller.tap_pos[1] ),
    .B(_01750_),
    .Y(_01751_));
 sg13g2_nand2_1 _09085_ (.Y(_01752_),
    .A(_01749_),
    .B(_01751_));
 sg13g2_inv_1 _09086_ (.Y(_01753_),
    .A(_01752_));
 sg13g2_inv_1 _09087_ (.Y(_01754_),
    .A(_01727_));
 sg13g2_nor2_1 _09088_ (.A(_01728_),
    .B(_01754_),
    .Y(_01755_));
 sg13g2_inv_2 _09089_ (.Y(_01756_),
    .A(_01755_));
 sg13g2_nor2_1 _09090_ (.A(_01733_),
    .B(_01756_),
    .Y(_01757_));
 sg13g2_nor2_2 _09091_ (.A(_01757_),
    .B(_01749_),
    .Y(_01758_));
 sg13g2_nor2_1 _09092_ (.A(_01757_),
    .B(_01753_),
    .Y(_01759_));
 sg13g2_nor2_1 _09093_ (.A(\synth.voice.scan_outs[11][0] ),
    .B(_01759_),
    .Y(_01760_));
 sg13g2_nor3_1 _09094_ (.A(_01753_),
    .B(_01758_),
    .C(_01760_),
    .Y(_01761_));
 sg13g2_or2_1 _09095_ (.X(_01762_),
    .B(_01761_),
    .A(_01747_));
 sg13g2_buf_1 _09096_ (.A(_01762_),
    .X(_01763_));
 sg13g2_nor2_1 _09097_ (.A(net202),
    .B(_01763_),
    .Y(_00005_));
 sg13g2_buf_1 _09098_ (.A(_01739_),
    .X(_01764_));
 sg13g2_buf_1 _09099_ (.A(\synth.voice.scan_outs[11][1] ),
    .X(_01765_));
 sg13g2_inv_1 _09100_ (.Y(_01766_),
    .A(\synth.voice.scan_outs[11][0] ));
 sg13g2_nor2_1 _09101_ (.A(_01765_),
    .B(_01766_),
    .Y(_01767_));
 sg13g2_nand2_1 _09102_ (.Y(_01768_),
    .A(_01753_),
    .B(_01767_));
 sg13g2_and3_1 _09103_ (.X(_00007_),
    .A(net201),
    .B(_01749_),
    .C(_01768_));
 sg13g2_inv_1 _09104_ (.Y(_01769_),
    .A(_01763_));
 sg13g2_nor2_1 _09105_ (.A(net202),
    .B(_01769_),
    .Y(_00003_));
 sg13g2_nand3b_1 _09106_ (.B(net201),
    .C(_01768_),
    .Y(_00006_),
    .A_N(_01757_));
 sg13g2_inv_1 _09107_ (.Y(_01770_),
    .A(\synth.voice.genblk4[9].next_state_scan[12] ));
 sg13g2_nand2_2 _09108_ (.Y(_01771_),
    .A(_01727_),
    .B(_01728_));
 sg13g2_inv_2 _09109_ (.Y(_01772_),
    .A(_01771_));
 sg13g2_buf_1 _09110_ (.A(_01772_),
    .X(_01773_));
 sg13g2_nand2_1 _09111_ (.Y(_01774_),
    .A(_01735_),
    .B(_01771_));
 sg13g2_buf_8 _09112_ (.A(_01774_),
    .X(_01775_));
 sg13g2_inv_1 _09113_ (.Y(_01776_),
    .A(_01775_));
 sg13g2_nor2_1 _09114_ (.A(\synth.voice.genblk4[10].next_state_scan[9] ),
    .B(_01735_),
    .Y(_01777_));
 sg13g2_a221oi_1 _09115_ (.B2(_00081_),
    .C1(_01777_),
    .B1(_01776_),
    .A1(_01770_),
    .Y(_01778_),
    .A2(_01773_));
 sg13g2_nand2_1 _09116_ (.Y(_01779_),
    .A(_01778_),
    .B(_01758_));
 sg13g2_inv_1 _09117_ (.Y(_01780_),
    .A(_01779_));
 sg13g2_inv_1 _09118_ (.Y(_01781_),
    .A(\synth.voice.genblk4[10].next_state_scan[11] ));
 sg13g2_nor2_1 _09119_ (.A(\synth.voice.params[24] ),
    .B(_01771_),
    .Y(_01782_));
 sg13g2_a221oi_1 _09120_ (.B2(_00083_),
    .C1(_01782_),
    .B1(_01776_),
    .A1(_01781_),
    .Y(_01783_),
    .A2(net300));
 sg13g2_inv_1 _09121_ (.Y(_01784_),
    .A(\synth.voice.genblk4[10].next_state_scan[10] ));
 sg13g2_nor2_1 _09122_ (.A(\synth.voice.genblk4[9].next_state_scan[13] ),
    .B(_01771_),
    .Y(_01785_));
 sg13g2_a221oi_1 _09123_ (.B2(_00082_),
    .C1(_01785_),
    .B1(_01776_),
    .A1(_01784_),
    .Y(_01786_),
    .A2(net300));
 sg13g2_nand3_1 _09124_ (.B(_01783_),
    .C(_01786_),
    .A(_01780_),
    .Y(_01787_));
 sg13g2_nand3_1 _09125_ (.B(_00080_),
    .C(net201),
    .A(_01787_),
    .Y(_01788_));
 sg13g2_nor2_1 _09126_ (.A(_01763_),
    .B(_01788_),
    .Y(_00010_));
 sg13g2_buf_2 _09127_ (.A(reset),
    .X(_01789_));
 sg13g2_buf_1 _09128_ (.A(_01789_),
    .X(_01790_));
 sg13g2_nor3_1 _09129_ (.A(net394),
    .B(_01731_),
    .C(_01719_),
    .Y(_00009_));
 sg13g2_nor2_1 _09130_ (.A(_01769_),
    .B(_01788_),
    .Y(_00008_));
 sg13g2_nand3_1 _09131_ (.B(_01720_),
    .C(\synth.controller.step_sample ),
    .A(_01750_),
    .Y(_01791_));
 sg13g2_nand2_1 _09132_ (.Y(_01792_),
    .A(\synth.controller.sample_counter[0] ),
    .B(\synth.controller.sample_counter[1] ));
 sg13g2_inv_1 _09133_ (.Y(_01793_),
    .A(_01715_));
 sg13g2_inv_1 _09134_ (.Y(_01794_),
    .A(_00045_));
 sg13g2_nor3_1 _09135_ (.A(_01716_),
    .B(_01793_),
    .C(_01794_),
    .Y(_01795_));
 sg13g2_buf_2 _09136_ (.A(_01795_),
    .X(_01796_));
 sg13g2_inv_1 _09137_ (.Y(_01797_),
    .A(_01796_));
 sg13g2_nor3_1 _09138_ (.A(_01791_),
    .B(_01792_),
    .C(_01797_),
    .Y(\synth.voice.restart_acc ));
 sg13g2_nor2_1 _09139_ (.A(\synth.voice.restart_acc ),
    .B(net201),
    .Y(_00004_));
 sg13g2_inv_1 _09140_ (.Y(_00000_),
    .A(net1));
 sg13g2_inv_1 _09141_ (.Y(_01798_),
    .A(_01789_));
 sg13g2_nand2_1 _09142_ (.Y(_01799_),
    .A(_01798_),
    .B(\ppu_ctrl[0] ));
 sg13g2_buf_1 _09143_ (.A(_01799_),
    .X(_01800_));
 sg13g2_buf_2 _09144_ (.A(\ppu.rs2.phase_x ),
    .X(_01801_));
 sg13g2_inv_2 _09145_ (.Y(_01802_),
    .A(_01801_));
 sg13g2_buf_1 _09146_ (.A(\ppu.copper_inst.x_cmp[4] ),
    .X(_01803_));
 sg13g2_inv_1 _09147_ (.Y(_01804_),
    .A(_01803_));
 sg13g2_buf_1 _09148_ (.A(_01801_),
    .X(_01805_));
 sg13g2_nor2b_1 _09149_ (.A(_01805_),
    .B_N(\ppu.gfxmode1[7] ),
    .Y(_01806_));
 sg13g2_a21oi_1 _09150_ (.A1(net393),
    .A2(\ppu.gfxmode3[4] ),
    .Y(_01807_),
    .B1(_01806_));
 sg13g2_xnor2_1 _09151_ (.Y(_01808_),
    .A(_01804_),
    .B(_01807_));
 sg13g2_nor2_1 _09152_ (.A(\ppu.gfxmode3[7] ),
    .B(_01802_),
    .Y(_01809_));
 sg13g2_xnor2_1 _09153_ (.Y(_01810_),
    .A(_00030_),
    .B(_01809_));
 sg13g2_buf_2 _09154_ (.A(\ppu.rs2.x0[6] ),
    .X(_01811_));
 sg13g2_inv_1 _09155_ (.Y(_01812_),
    .A(_01811_));
 sg13g2_nand2_1 _09156_ (.Y(_01813_),
    .A(net393),
    .B(\ppu.gfxmode3[6] ));
 sg13g2_xnor2_1 _09157_ (.Y(_01814_),
    .A(_01812_),
    .B(_01813_));
 sg13g2_nand3_1 _09158_ (.B(_01810_),
    .C(_01814_),
    .A(_01808_),
    .Y(_01815_));
 sg13g2_buf_2 _09159_ (.A(\ppu.copper_inst.x_cmp[1] ),
    .X(_01816_));
 sg13g2_buf_1 _09160_ (.A(net393),
    .X(_01817_));
 sg13g2_nor2b_1 _09161_ (.A(net347),
    .B_N(\ppu.gfxmode1[4] ),
    .Y(_01818_));
 sg13g2_a21oi_1 _09162_ (.A1(net347),
    .A2(\ppu.gfxmode3[1] ),
    .Y(_01819_),
    .B1(_01818_));
 sg13g2_xnor2_1 _09163_ (.Y(_01820_),
    .A(_01816_),
    .B(_01819_));
 sg13g2_buf_1 _09164_ (.A(\ppu.copper_inst.x_cmp[0] ),
    .X(_01821_));
 sg13g2_buf_1 _09165_ (.A(net409),
    .X(_01822_));
 sg13g2_buf_1 _09166_ (.A(net392),
    .X(_01823_));
 sg13g2_nor2b_1 _09167_ (.A(net347),
    .B_N(\ppu.gfxmode1[3] ),
    .Y(_01824_));
 sg13g2_a21oi_1 _09168_ (.A1(net347),
    .A2(\ppu.gfxmode3[0] ),
    .Y(_01825_),
    .B1(_01824_));
 sg13g2_xnor2_1 _09169_ (.Y(_01826_),
    .A(net346),
    .B(_01825_));
 sg13g2_buf_2 _09170_ (.A(\ppu.copper_inst.x_cmp[8] ),
    .X(_01827_));
 sg13g2_nand2_1 _09171_ (.Y(_01828_),
    .A(net393),
    .B(\ppu.gfxmode3[8] ));
 sg13g2_xnor2_1 _09172_ (.Y(_01829_),
    .A(_01827_),
    .B(_01828_));
 sg13g2_buf_2 _09173_ (.A(\ppu.rs2.x0[5] ),
    .X(_01830_));
 sg13g2_inv_1 _09174_ (.Y(_01831_),
    .A(_01830_));
 sg13g2_inv_1 _09175_ (.Y(_01832_),
    .A(\ppu.gfxmode1[8] ));
 sg13g2_nand2_1 _09176_ (.Y(_01833_),
    .A(_01801_),
    .B(\ppu.gfxmode3[5] ));
 sg13g2_o21ai_1 _09177_ (.B1(_01833_),
    .Y(_01834_),
    .A1(net393),
    .A2(_01832_));
 sg13g2_nor2_1 _09178_ (.A(_01831_),
    .B(_01834_),
    .Y(_01835_));
 sg13g2_buf_2 _09179_ (.A(\ppu.copper_inst.x_cmp[3] ),
    .X(_01836_));
 sg13g2_inv_1 _09180_ (.Y(_01837_),
    .A(_01836_));
 sg13g2_inv_1 _09181_ (.Y(_01838_),
    .A(\ppu.gfxmode1[6] ));
 sg13g2_nand2_1 _09182_ (.Y(_01839_),
    .A(_01801_),
    .B(\ppu.gfxmode3[3] ));
 sg13g2_o21ai_1 _09183_ (.B1(_01839_),
    .Y(_01840_),
    .A1(net393),
    .A2(_01838_));
 sg13g2_nor2_1 _09184_ (.A(_01837_),
    .B(_01840_),
    .Y(_01841_));
 sg13g2_nor2b_1 _09185_ (.A(_01830_),
    .B_N(_01834_),
    .Y(_01842_));
 sg13g2_nor4_1 _09186_ (.A(_01829_),
    .B(_01835_),
    .C(_01841_),
    .D(_01842_),
    .Y(_01843_));
 sg13g2_inv_1 _09187_ (.Y(_01844_),
    .A(\ppu.copper_inst.x_cmp[2] ));
 sg13g2_nor2b_1 _09188_ (.A(net393),
    .B_N(\ppu.gfxmode1[5] ),
    .Y(_01845_));
 sg13g2_a21oi_1 _09189_ (.A1(\ppu.gfxmode3[2] ),
    .A2(net393),
    .Y(_01846_),
    .B1(_01845_));
 sg13g2_xnor2_1 _09190_ (.Y(_01847_),
    .A(_01844_),
    .B(_01846_));
 sg13g2_nand2_1 _09191_ (.Y(_01848_),
    .A(_01840_),
    .B(_01837_));
 sg13g2_nand3_1 _09192_ (.B(_01847_),
    .C(_01848_),
    .A(_01843_),
    .Y(_01849_));
 sg13g2_nor4_2 _09193_ (.A(_01815_),
    .B(_01820_),
    .C(_01826_),
    .Y(_01850_),
    .D(_01849_));
 sg13g2_nor2b_1 _09194_ (.A(_01802_),
    .B_N(_01850_),
    .Y(_01851_));
 sg13g2_nor2_1 _09195_ (.A(net298),
    .B(_01851_),
    .Y(_01852_));
 sg13g2_buf_1 _09196_ (.A(_01852_),
    .X(_01853_));
 sg13g2_buf_8 _09197_ (.A(\ppu.copper_inst.serial_counter[1] ),
    .X(_01854_));
 sg13g2_buf_8 _09198_ (.A(\ppu.copper_inst.serial_counter[0] ),
    .X(_01855_));
 sg13g2_nand2_1 _09199_ (.Y(_01856_),
    .A(_01854_),
    .B(_01855_));
 sg13g2_buf_8 _09200_ (.A(_01856_),
    .X(_01857_));
 sg13g2_buf_1 _09201_ (.A(\ppu.sprite_buffer.scan_on ),
    .X(_01858_));
 sg13g2_buf_1 _09202_ (.A(\ppu.copper_inst.dt_out[1] ),
    .X(_01859_));
 sg13g2_buf_1 _09203_ (.A(\ppu.copper_inst.dt_out[0] ),
    .X(_01860_));
 sg13g2_inv_1 _09204_ (.Y(_01861_),
    .A(_01860_));
 sg13g2_inv_1 _09205_ (.Y(_01862_),
    .A(_00031_));
 sg13g2_nor3_2 _09206_ (.A(_01859_),
    .B(_01861_),
    .C(_01862_),
    .Y(_01863_));
 sg13g2_nand2b_1 _09207_ (.Y(_01864_),
    .B(_01863_),
    .A_N(_01858_));
 sg13g2_buf_2 _09208_ (.A(\ppu.rs2.y_scan.counter[0] ),
    .X(_01865_));
 sg13g2_buf_1 _09209_ (.A(\data_pins[3] ),
    .X(_01866_));
 sg13g2_inv_2 _09210_ (.Y(_01867_),
    .A(net408));
 sg13g2_inv_1 _09211_ (.Y(_01868_),
    .A(\ppu.sprite_buffer.y_matched0 ));
 sg13g2_a21oi_1 _09212_ (.A1(_01865_),
    .A2(\data_pins[2] ),
    .Y(_01869_),
    .B1(_01868_));
 sg13g2_o21ai_1 _09213_ (.B1(_01869_),
    .Y(_01870_),
    .A1(_01865_),
    .A2(_01867_));
 sg13g2_buf_1 _09214_ (.A(\ppu.sprite_buffer.in_counter_idy[0] ),
    .X(_01871_));
 sg13g2_buf_1 _09215_ (.A(\ppu.sprite_buffer.in_counter_idy[1] ),
    .X(_01872_));
 sg13g2_inv_1 _09216_ (.Y(_01873_),
    .A(_01872_));
 sg13g2_nor2_1 _09217_ (.A(_01871_),
    .B(_01873_),
    .Y(_01874_));
 sg13g2_inv_1 _09218_ (.Y(_01875_),
    .A(_01871_));
 sg13g2_nor2_1 _09219_ (.A(_01872_),
    .B(_01875_),
    .Y(_01876_));
 sg13g2_nor3_1 _09220_ (.A(_00077_),
    .B(_01874_),
    .C(_01876_),
    .Y(_01877_));
 sg13g2_buf_1 _09221_ (.A(\ppu.sprite_buffer.out_counter_oam[0] ),
    .X(_01878_));
 sg13g2_xnor2_1 _09222_ (.Y(_01879_),
    .A(_01878_),
    .B(_01871_));
 sg13g2_inv_1 _09223_ (.Y(_01880_),
    .A(_01879_));
 sg13g2_o21ai_1 _09224_ (.B1(_00077_),
    .Y(_01881_),
    .A1(_01874_),
    .A2(_01876_));
 sg13g2_nand3b_1 _09225_ (.B(_01880_),
    .C(_01881_),
    .Y(_01882_),
    .A_N(_01877_));
 sg13g2_nand2_1 _09226_ (.Y(_01883_),
    .A(_01882_),
    .B(_01858_));
 sg13g2_inv_1 _09227_ (.Y(_01884_),
    .A(_01883_));
 sg13g2_a21oi_1 _09228_ (.A1(_01864_),
    .A2(_01870_),
    .Y(_01885_),
    .B1(_01884_));
 sg13g2_inv_1 _09229_ (.Y(_01886_),
    .A(_01885_));
 sg13g2_nor2_1 _09230_ (.A(net345),
    .B(_01886_),
    .Y(_01887_));
 sg13g2_inv_1 _09231_ (.Y(_01888_),
    .A(_01887_));
 sg13g2_nand2_1 _09232_ (.Y(_01889_),
    .A(_01888_),
    .B(_01858_));
 sg13g2_buf_1 _09233_ (.A(net345),
    .X(_01890_));
 sg13g2_buf_1 _09234_ (.A(net297),
    .X(_01891_));
 sg13g2_inv_1 _09235_ (.Y(_01892_),
    .A(\ppu.copper_inst.dt_sreg[6] ));
 sg13g2_nor3_1 _09236_ (.A(\ppu.copper_inst.dt_sreg[7] ),
    .B(\ppu.copper_inst.dt_sreg[8] ),
    .C(_01892_),
    .Y(_01893_));
 sg13g2_nor4_1 _09237_ (.A(_01858_),
    .B(net264),
    .C(_01893_),
    .D(_01863_),
    .Y(_01894_));
 sg13g2_inv_1 _09238_ (.Y(_01895_),
    .A(\ppu.copper_inst.dt_sreg[4] ));
 sg13g2_nand3_1 _09239_ (.B(\ppu.copper_inst.dt_sreg[3] ),
    .C(_00035_),
    .A(_01895_),
    .Y(_01896_));
 sg13g2_inv_1 _09240_ (.Y(_01897_),
    .A(\ppu.copper_inst.dt_sreg[10] ));
 sg13g2_inv_1 _09241_ (.Y(_01898_),
    .A(\ppu.copper_inst.dt_sreg[11] ));
 sg13g2_nand3_1 _09242_ (.B(_01898_),
    .C(\ppu.copper_inst.dt_sreg[9] ),
    .A(_01897_),
    .Y(_01899_));
 sg13g2_nand4_1 _09243_ (.B(_01894_),
    .C(_01896_),
    .A(_01882_),
    .Y(_01900_),
    .D(_01899_));
 sg13g2_nand3_1 _09244_ (.B(_01889_),
    .C(_01900_),
    .A(_01853_),
    .Y(_00015_));
 sg13g2_inv_1 _09245_ (.Y(_01901_),
    .A(_01859_));
 sg13g2_nor3_2 _09246_ (.A(\ppu.copper_inst.dt_out[2] ),
    .B(_01901_),
    .C(_01861_),
    .Y(_01902_));
 sg13g2_inv_4 _09247_ (.A(net345),
    .Y(_01903_));
 sg13g2_buf_1 _09248_ (.A(_01903_),
    .X(_01904_));
 sg13g2_buf_1 _09249_ (.A(_01904_),
    .X(_01905_));
 sg13g2_nand2_1 _09250_ (.Y(_01906_),
    .A(_01902_),
    .B(net254));
 sg13g2_inv_1 _09251_ (.Y(_01907_),
    .A(_01906_));
 sg13g2_inv_1 _09252_ (.Y(_01908_),
    .A(\ppu.sprite_buffer.final_pixels_in ));
 sg13g2_buf_1 _09253_ (.A(\ppu.sprite_buffer.in_counters[2][1] ),
    .X(_01909_));
 sg13g2_nand3_1 _09254_ (.B(_01909_),
    .C(\ppu.sprite_buffer.in_counters[2][2] ),
    .A(_01902_),
    .Y(_01910_));
 sg13g2_nor2_1 _09255_ (.A(_01908_),
    .B(_01910_),
    .Y(_01911_));
 sg13g2_inv_1 _09256_ (.Y(_01912_),
    .A(_01853_));
 sg13g2_buf_1 _09257_ (.A(_01912_),
    .X(_01913_));
 sg13g2_a21oi_1 _09258_ (.A1(_01907_),
    .A2(_01911_),
    .Y(_01914_),
    .B1(net146));
 sg13g2_buf_1 _09259_ (.A(_01914_),
    .X(_01915_));
 sg13g2_inv_1 _09260_ (.Y(_01916_),
    .A(_00063_));
 sg13g2_inv_2 _09261_ (.Y(_01917_),
    .A(_01854_));
 sg13g2_inv_8 _09262_ (.Y(_01918_),
    .A(_01855_));
 sg13g2_nand2_1 _09263_ (.Y(_01919_),
    .A(_01917_),
    .B(net391));
 sg13g2_buf_2 _09264_ (.A(_01919_),
    .X(_01920_));
 sg13g2_buf_1 _09265_ (.A(_01920_),
    .X(_01921_));
 sg13g2_nor2_1 _09266_ (.A(_01855_),
    .B(_01917_),
    .Y(_01922_));
 sg13g2_buf_2 _09267_ (.A(_01922_),
    .X(_01923_));
 sg13g2_a22oi_1 _09268_ (.Y(_01924_),
    .B1(\ppu.sprite_buffer.attr_x[3][7] ),
    .B2(net263),
    .A2(\ppu.sprite_buffer.attr_x[2][7] ),
    .A1(_01923_));
 sg13g2_nor2_1 _09269_ (.A(_01854_),
    .B(_01918_),
    .Y(_01925_));
 sg13g2_buf_1 _09270_ (.A(_01925_),
    .X(_01926_));
 sg13g2_buf_1 _09271_ (.A(net296),
    .X(_01927_));
 sg13g2_nand2_1 _09272_ (.Y(_01928_),
    .A(net261),
    .B(\ppu.sprite_buffer.attr_x[1][7] ));
 sg13g2_nand3_1 _09273_ (.B(_01920_),
    .C(_01928_),
    .A(_01924_),
    .Y(_01929_));
 sg13g2_o21ai_1 _09274_ (.B1(_01929_),
    .Y(_01930_),
    .A1(_01916_),
    .A2(net262));
 sg13g2_xor2_1 _09275_ (.B(_01930_),
    .A(_00030_),
    .X(_01931_));
 sg13g2_inv_1 _09276_ (.Y(_01932_),
    .A(_00071_));
 sg13g2_buf_1 _09277_ (.A(_01917_),
    .X(_01933_));
 sg13g2_o21ai_1 _09278_ (.B1(net391),
    .Y(_01934_),
    .A1(\ppu.sprite_buffer.attr_x[2][1] ),
    .A2(net344));
 sg13g2_nand2_1 _09279_ (.Y(_01935_),
    .A(_01903_),
    .B(\ppu.sprite_buffer.attr_x[3][1] ));
 sg13g2_nand2_1 _09280_ (.Y(_01936_),
    .A(net296),
    .B(\ppu.sprite_buffer.attr_x[1][1] ));
 sg13g2_nand3_1 _09281_ (.B(_01935_),
    .C(_01936_),
    .A(_01934_),
    .Y(_01937_));
 sg13g2_o21ai_1 _09282_ (.B1(_01937_),
    .Y(_01938_),
    .A1(_01932_),
    .A2(_01920_));
 sg13g2_xnor2_1 _09283_ (.Y(_01939_),
    .A(_00033_),
    .B(_01938_));
 sg13g2_a22oi_1 _09284_ (.Y(_01940_),
    .B1(\ppu.sprite_buffer.attr_x[3][0] ),
    .B2(_01903_),
    .A2(\ppu.sprite_buffer.attr_x[2][0] ),
    .A1(_01923_));
 sg13g2_nand2_1 _09285_ (.Y(_01941_),
    .A(net296),
    .B(\ppu.sprite_buffer.attr_x[1][0] ));
 sg13g2_nand3_1 _09286_ (.B(_01920_),
    .C(_01941_),
    .A(_01940_),
    .Y(_01942_));
 sg13g2_buf_2 _09287_ (.A(_00032_),
    .X(_01943_));
 sg13g2_inv_4 _09288_ (.A(_01920_),
    .Y(_01944_));
 sg13g2_nand2_1 _09289_ (.Y(_01945_),
    .A(net260),
    .B(_00072_));
 sg13g2_nand3_1 _09290_ (.B(_01943_),
    .C(_01945_),
    .A(_01942_),
    .Y(_01946_));
 sg13g2_buf_1 _09291_ (.A(_01946_),
    .X(_01947_));
 sg13g2_nand2_1 _09292_ (.Y(_01948_),
    .A(_01939_),
    .B(_01947_));
 sg13g2_inv_1 _09293_ (.Y(_01949_),
    .A(_01948_));
 sg13g2_o21ai_1 _09294_ (.B1(net391),
    .Y(_01950_),
    .A1(\ppu.sprite_buffer.attr_x[2][2] ),
    .A2(net344));
 sg13g2_nand2_1 _09295_ (.Y(_01951_),
    .A(_01903_),
    .B(\ppu.sprite_buffer.attr_x[3][2] ));
 sg13g2_nand2_1 _09296_ (.Y(_01952_),
    .A(net296),
    .B(\ppu.sprite_buffer.attr_x[1][2] ));
 sg13g2_nand3_1 _09297_ (.B(_01951_),
    .C(_01952_),
    .A(_01950_),
    .Y(_01953_));
 sg13g2_nand2_1 _09298_ (.Y(_01954_),
    .A(net260),
    .B(_00070_));
 sg13g2_nand2_1 _09299_ (.Y(_01955_),
    .A(_01953_),
    .B(_01954_));
 sg13g2_inv_1 _09300_ (.Y(_01956_),
    .A(_01955_));
 sg13g2_inv_1 _09301_ (.Y(_01957_),
    .A(_00034_));
 sg13g2_nand2_1 _09302_ (.Y(_01958_),
    .A(_01956_),
    .B(_01957_));
 sg13g2_nand2_1 _09303_ (.Y(_01959_),
    .A(_01955_),
    .B(_00034_));
 sg13g2_nand2_1 _09304_ (.Y(_01960_),
    .A(_01958_),
    .B(_01959_));
 sg13g2_nand2_1 _09305_ (.Y(_01961_),
    .A(_01949_),
    .B(_01960_));
 sg13g2_nand2_1 _09306_ (.Y(_01962_),
    .A(_01938_),
    .B(_01816_));
 sg13g2_inv_1 _09307_ (.Y(_01963_),
    .A(_01962_));
 sg13g2_nor2_1 _09308_ (.A(_01844_),
    .B(_01956_),
    .Y(_01964_));
 sg13g2_a21oi_1 _09309_ (.A1(_01960_),
    .A2(_01963_),
    .Y(_01965_),
    .B1(_01964_));
 sg13g2_nand2_1 _09310_ (.Y(_01966_),
    .A(_01961_),
    .B(_01965_));
 sg13g2_inv_1 _09311_ (.Y(_01967_),
    .A(_00064_));
 sg13g2_o21ai_1 _09312_ (.B1(net391),
    .Y(_01968_),
    .A1(\ppu.sprite_buffer.attr_x[2][6] ),
    .A2(net344));
 sg13g2_nand2_1 _09313_ (.Y(_01969_),
    .A(_01903_),
    .B(\ppu.sprite_buffer.attr_x[3][6] ));
 sg13g2_nand2_1 _09314_ (.Y(_01970_),
    .A(net261),
    .B(\ppu.sprite_buffer.attr_x[1][6] ));
 sg13g2_nand3_1 _09315_ (.B(_01969_),
    .C(_01970_),
    .A(_01968_),
    .Y(_01971_));
 sg13g2_o21ai_1 _09316_ (.B1(_01971_),
    .Y(_01972_),
    .A1(_01967_),
    .A2(net262));
 sg13g2_xnor2_1 _09317_ (.Y(_01973_),
    .A(_00065_),
    .B(_01972_));
 sg13g2_inv_1 _09318_ (.Y(_01974_),
    .A(_00066_));
 sg13g2_o21ai_1 _09319_ (.B1(net391),
    .Y(_01975_),
    .A1(\ppu.sprite_buffer.attr_x[2][5] ),
    .A2(net344));
 sg13g2_nand2_1 _09320_ (.Y(_01976_),
    .A(_01903_),
    .B(\ppu.sprite_buffer.attr_x[3][5] ));
 sg13g2_nand2_1 _09321_ (.Y(_01977_),
    .A(net296),
    .B(\ppu.sprite_buffer.attr_x[1][5] ));
 sg13g2_nand3_1 _09322_ (.B(_01976_),
    .C(_01977_),
    .A(_01975_),
    .Y(_01978_));
 sg13g2_o21ai_1 _09323_ (.B1(_01978_),
    .Y(_01979_),
    .A1(_01974_),
    .A2(_01920_));
 sg13g2_xnor2_1 _09324_ (.Y(_01980_),
    .A(_00067_),
    .B(_01979_));
 sg13g2_nand2_1 _09325_ (.Y(_01981_),
    .A(_01973_),
    .B(_01980_));
 sg13g2_o21ai_1 _09326_ (.B1(net391),
    .Y(_01982_),
    .A1(\ppu.sprite_buffer.attr_x[2][4] ),
    .A2(net344));
 sg13g2_nand2_1 _09327_ (.Y(_01983_),
    .A(_01903_),
    .B(\ppu.sprite_buffer.attr_x[3][4] ));
 sg13g2_nand2_1 _09328_ (.Y(_01984_),
    .A(net296),
    .B(\ppu.sprite_buffer.attr_x[1][4] ));
 sg13g2_nand3_1 _09329_ (.B(_01983_),
    .C(_01984_),
    .A(_01982_),
    .Y(_01985_));
 sg13g2_nand2_1 _09330_ (.Y(_01986_),
    .A(net260),
    .B(_00068_));
 sg13g2_nand2_1 _09331_ (.Y(_01987_),
    .A(_01985_),
    .B(_01986_));
 sg13g2_inv_1 _09332_ (.Y(_01988_),
    .A(_01987_));
 sg13g2_nor2_1 _09333_ (.A(_01804_),
    .B(_01988_),
    .Y(_01989_));
 sg13g2_inv_1 _09334_ (.Y(_01990_),
    .A(_01989_));
 sg13g2_nor2_1 _09335_ (.A(_01803_),
    .B(_01987_),
    .Y(_01991_));
 sg13g2_inv_1 _09336_ (.Y(_01992_),
    .A(_01991_));
 sg13g2_nand2_1 _09337_ (.Y(_01993_),
    .A(_01990_),
    .B(_01992_));
 sg13g2_inv_1 _09338_ (.Y(_01994_),
    .A(_00069_));
 sg13g2_o21ai_1 _09339_ (.B1(net391),
    .Y(_01995_),
    .A1(\ppu.sprite_buffer.attr_x[2][3] ),
    .A2(_01933_));
 sg13g2_nand2_1 _09340_ (.Y(_01996_),
    .A(_01903_),
    .B(\ppu.sprite_buffer.attr_x[3][3] ));
 sg13g2_nand2_1 _09341_ (.Y(_01997_),
    .A(net296),
    .B(\ppu.sprite_buffer.attr_x[1][3] ));
 sg13g2_nand3_1 _09342_ (.B(_01996_),
    .C(_01997_),
    .A(_01995_),
    .Y(_01998_));
 sg13g2_o21ai_1 _09343_ (.B1(_01998_),
    .Y(_01999_),
    .A1(_01994_),
    .A2(_01920_));
 sg13g2_nor2_1 _09344_ (.A(_01836_),
    .B(_01999_),
    .Y(_02000_));
 sg13g2_inv_1 _09345_ (.Y(_02001_),
    .A(_02000_));
 sg13g2_nand2_1 _09346_ (.Y(_02002_),
    .A(_01999_),
    .B(_01836_));
 sg13g2_nand2_1 _09347_ (.Y(_02003_),
    .A(_02001_),
    .B(_02002_));
 sg13g2_nor2_1 _09348_ (.A(_01993_),
    .B(_02003_),
    .Y(_02004_));
 sg13g2_inv_1 _09349_ (.Y(_02005_),
    .A(_02004_));
 sg13g2_nor2_1 _09350_ (.A(_01981_),
    .B(_02005_),
    .Y(_02006_));
 sg13g2_nand2_1 _09351_ (.Y(_02007_),
    .A(_01966_),
    .B(_02006_));
 sg13g2_inv_1 _09352_ (.Y(_02008_),
    .A(_02002_));
 sg13g2_a21oi_1 _09353_ (.A1(_02008_),
    .A2(_01992_),
    .Y(_02009_),
    .B1(_01989_));
 sg13g2_nor2_1 _09354_ (.A(_01981_),
    .B(_02009_),
    .Y(_02010_));
 sg13g2_nand2_1 _09355_ (.Y(_02011_),
    .A(_01979_),
    .B(_01830_));
 sg13g2_inv_1 _09356_ (.Y(_02012_),
    .A(_01973_));
 sg13g2_nand2_1 _09357_ (.Y(_02013_),
    .A(_01972_),
    .B(_01811_));
 sg13g2_o21ai_1 _09358_ (.B1(_02013_),
    .Y(_02014_),
    .A1(_02011_),
    .A2(_02012_));
 sg13g2_nor2_1 _09359_ (.A(_02010_),
    .B(_02014_),
    .Y(_02015_));
 sg13g2_nand2_1 _09360_ (.Y(_02016_),
    .A(_02007_),
    .B(_02015_));
 sg13g2_xnor2_1 _09361_ (.Y(_02017_),
    .A(_01931_),
    .B(_02016_));
 sg13g2_nand2_1 _09362_ (.Y(_02018_),
    .A(_01948_),
    .B(_01962_));
 sg13g2_inv_1 _09363_ (.Y(_02019_),
    .A(_01960_));
 sg13g2_nor2_1 _09364_ (.A(_02019_),
    .B(_02003_),
    .Y(_02020_));
 sg13g2_nand2_1 _09365_ (.Y(_02021_),
    .A(_02018_),
    .B(_02020_));
 sg13g2_a21oi_1 _09366_ (.A1(_02001_),
    .A2(_01964_),
    .Y(_02022_),
    .B1(_02008_));
 sg13g2_nand2_1 _09367_ (.Y(_02023_),
    .A(_02021_),
    .B(_02022_));
 sg13g2_xor2_1 _09368_ (.B(_02023_),
    .A(_01993_),
    .X(_02024_));
 sg13g2_nand2b_1 _09369_ (.Y(_02025_),
    .B(_01966_),
    .A_N(_02003_));
 sg13g2_nand3_1 _09370_ (.B(_01965_),
    .C(_02003_),
    .A(_01961_),
    .Y(_02026_));
 sg13g2_nand2_1 _09371_ (.Y(_02027_),
    .A(_01926_),
    .B(\ppu.sprite_buffer.attr_x[1][13] ));
 sg13g2_inv_2 _09372_ (.Y(_02028_),
    .A(_01923_));
 sg13g2_inv_1 _09373_ (.Y(_02029_),
    .A(\ppu.sprite_buffer.attr_x[3][13] ));
 sg13g2_o21ai_1 _09374_ (.B1(_01855_),
    .Y(_02030_),
    .A1(net344),
    .A2(_02029_));
 sg13g2_o21ai_1 _09375_ (.B1(_02030_),
    .Y(_02031_),
    .A1(\ppu.sprite_buffer.attr_x[2][13] ),
    .A2(_02028_));
 sg13g2_a22oi_1 _09376_ (.Y(_02032_),
    .B1(_02027_),
    .B2(_02031_),
    .A2(net260),
    .A1(_00073_));
 sg13g2_inv_1 _09377_ (.Y(_02033_),
    .A(_02032_));
 sg13g2_nand2_1 _09378_ (.Y(_02034_),
    .A(_01926_),
    .B(\ppu.sprite_buffer.attr_x[1][14] ));
 sg13g2_inv_1 _09379_ (.Y(_02035_),
    .A(\ppu.sprite_buffer.attr_x[3][14] ));
 sg13g2_o21ai_1 _09380_ (.B1(_01855_),
    .Y(_02036_),
    .A1(net344),
    .A2(_02035_));
 sg13g2_o21ai_1 _09381_ (.B1(_02036_),
    .Y(_02037_),
    .A1(\ppu.sprite_buffer.attr_x[2][14] ),
    .A2(_02028_));
 sg13g2_a22oi_1 _09382_ (.Y(_02038_),
    .B1(_02034_),
    .B2(_02037_),
    .A2(net260),
    .A1(_00074_));
 sg13g2_inv_1 _09383_ (.Y(_02039_),
    .A(_02038_));
 sg13g2_nor2_1 _09384_ (.A(_02033_),
    .B(_02039_),
    .Y(_02040_));
 sg13g2_inv_1 _09385_ (.Y(_02041_),
    .A(\ppu.sprite_buffer.attr_x[1][12] ));
 sg13g2_inv_1 _09386_ (.Y(_02042_),
    .A(net296));
 sg13g2_nor2_1 _09387_ (.A(_02041_),
    .B(_02042_),
    .Y(_02043_));
 sg13g2_inv_1 _09388_ (.Y(_02044_),
    .A(\ppu.sprite_buffer.attr_x[0][12] ));
 sg13g2_nor2_1 _09389_ (.A(_02044_),
    .B(_01920_),
    .Y(_02045_));
 sg13g2_inv_1 _09390_ (.Y(_02046_),
    .A(\ppu.sprite_buffer.attr_x[3][12] ));
 sg13g2_nand2_1 _09391_ (.Y(_02047_),
    .A(_01923_),
    .B(\ppu.sprite_buffer.attr_x[2][12] ));
 sg13g2_o21ai_1 _09392_ (.B1(_02047_),
    .Y(_02048_),
    .A1(_02046_),
    .A2(net345));
 sg13g2_or3_1 _09393_ (.A(_02043_),
    .B(_02045_),
    .C(_02048_),
    .X(_02049_));
 sg13g2_buf_1 _09394_ (.A(_02049_),
    .X(_02050_));
 sg13g2_buf_1 _09395_ (.A(net260),
    .X(_02051_));
 sg13g2_nand2_1 _09396_ (.Y(_02052_),
    .A(_01927_),
    .B(\ppu.sprite_buffer.attr_x[1][15] ));
 sg13g2_buf_1 _09397_ (.A(net391),
    .X(_02053_));
 sg13g2_a221oi_1 _09398_ (.B2(\ppu.sprite_buffer.attr_x[3][15] ),
    .C1(_01944_),
    .B1(net263),
    .A1(_02053_),
    .Y(_02054_),
    .A2(\ppu.sprite_buffer.attr_x[2][15] ));
 sg13g2_a22oi_1 _09399_ (.Y(_02055_),
    .B1(_02052_),
    .B2(_02054_),
    .A2(net253),
    .A1(_00075_));
 sg13g2_nand3_1 _09400_ (.B(_02050_),
    .C(_02055_),
    .A(_02040_),
    .Y(_02056_));
 sg13g2_buf_1 _09401_ (.A(_02056_),
    .X(_02057_));
 sg13g2_buf_1 _09402_ (.A(_02057_),
    .X(_02058_));
 sg13g2_inv_2 _09403_ (.Y(_02059_),
    .A(net145));
 sg13g2_nand3_1 _09404_ (.B(_02026_),
    .C(_02059_),
    .A(_02025_),
    .Y(_02060_));
 sg13g2_nand3_1 _09405_ (.B(_02060_),
    .C(_01817_),
    .A(_02024_),
    .Y(_02061_));
 sg13g2_nor2_1 _09406_ (.A(_02017_),
    .B(_02061_),
    .Y(_02062_));
 sg13g2_buf_1 _09407_ (.A(_01855_),
    .X(_02063_));
 sg13g2_inv_1 _09408_ (.Y(_02064_),
    .A(\ppu.sprite_buffer.attr_x[2][8] ));
 sg13g2_a22oi_1 _09409_ (.Y(_02065_),
    .B1(\ppu.sprite_buffer.attr_x[3][8] ),
    .B2(net263),
    .A2(\ppu.sprite_buffer.attr_x[1][8] ),
    .A1(net261));
 sg13g2_o21ai_1 _09410_ (.B1(_02065_),
    .Y(_02066_),
    .A1(_02063_),
    .A2(_02064_));
 sg13g2_nand2_1 _09411_ (.Y(_02067_),
    .A(net253),
    .B(_00062_));
 sg13g2_o21ai_1 _09412_ (.B1(_02067_),
    .Y(_02068_),
    .A1(net253),
    .A2(_02066_));
 sg13g2_xnor2_1 _09413_ (.Y(_02069_),
    .A(_00040_),
    .B(_02068_));
 sg13g2_inv_1 _09414_ (.Y(_02070_),
    .A(_01980_));
 sg13g2_nor2_1 _09415_ (.A(_01993_),
    .B(_02070_),
    .Y(_02071_));
 sg13g2_nor2_1 _09416_ (.A(_02012_),
    .B(_01931_),
    .Y(_02072_));
 sg13g2_nand3_1 _09417_ (.B(_02071_),
    .C(_02072_),
    .A(_02023_),
    .Y(_02073_));
 sg13g2_o21ai_1 _09418_ (.B1(_02011_),
    .Y(_02074_),
    .A1(_01990_),
    .A2(_02070_));
 sg13g2_buf_2 _09419_ (.A(\ppu.rs2.x0[7] ),
    .X(_02075_));
 sg13g2_nand2_1 _09420_ (.Y(_02076_),
    .A(_01930_),
    .B(_02075_));
 sg13g2_o21ai_1 _09421_ (.B1(_02076_),
    .Y(_02077_),
    .A1(_02013_),
    .A2(_01931_));
 sg13g2_a21oi_1 _09422_ (.A1(_02074_),
    .A2(_02072_),
    .Y(_02078_),
    .B1(_02077_));
 sg13g2_nand2_1 _09423_ (.Y(_02079_),
    .A(_02073_),
    .B(_02078_));
 sg13g2_xnor2_1 _09424_ (.Y(_02080_),
    .A(_02069_),
    .B(_02079_));
 sg13g2_nand4_1 _09425_ (.B(_01947_),
    .C(_01960_),
    .A(_02004_),
    .Y(_02081_),
    .D(_01939_));
 sg13g2_nor2_1 _09426_ (.A(_01965_),
    .B(_02005_),
    .Y(_02082_));
 sg13g2_nor2b_1 _09427_ (.A(_02082_),
    .B_N(_02009_),
    .Y(_02083_));
 sg13g2_nand2_1 _09428_ (.Y(_02084_),
    .A(_02081_),
    .B(_02083_));
 sg13g2_xnor2_1 _09429_ (.Y(_02085_),
    .A(_02070_),
    .B(_02084_));
 sg13g2_inv_1 _09430_ (.Y(_02086_),
    .A(_02022_));
 sg13g2_a21oi_1 _09431_ (.A1(_02086_),
    .A2(_02071_),
    .Y(_02087_),
    .B1(_02074_));
 sg13g2_nand3_1 _09432_ (.B(_02020_),
    .C(_02071_),
    .A(_02018_),
    .Y(_02088_));
 sg13g2_nand2_1 _09433_ (.Y(_02089_),
    .A(_02087_),
    .B(_02088_));
 sg13g2_xnor2_1 _09434_ (.Y(_02090_),
    .A(_02012_),
    .B(_02089_));
 sg13g2_nor2_1 _09435_ (.A(_02085_),
    .B(_02090_),
    .Y(_02091_));
 sg13g2_nand3_1 _09436_ (.B(_02080_),
    .C(_02091_),
    .A(_02062_),
    .Y(_02092_));
 sg13g2_nor2_2 _09437_ (.A(_01912_),
    .B(_02092_),
    .Y(_02093_));
 sg13g2_nand2_1 _09438_ (.Y(_02094_),
    .A(_01942_),
    .B(_01945_));
 sg13g2_inv_2 _09439_ (.Y(_02095_),
    .A(_01943_));
 sg13g2_nand2_1 _09440_ (.Y(_02096_),
    .A(_02094_),
    .B(_02095_));
 sg13g2_nand2_1 _09441_ (.Y(_02097_),
    .A(_02096_),
    .B(_01947_));
 sg13g2_buf_2 _09442_ (.A(_02097_),
    .X(_02098_));
 sg13g2_xor2_1 _09443_ (.B(_01939_),
    .A(_01947_),
    .X(_02099_));
 sg13g2_nand2_1 _09444_ (.Y(_02100_),
    .A(_02099_),
    .B(_02098_));
 sg13g2_inv_1 _09445_ (.Y(_02101_),
    .A(_02100_));
 sg13g2_a21oi_1 _09446_ (.A1(_02096_),
    .A2(_01949_),
    .Y(_02102_),
    .B1(_02101_));
 sg13g2_nor2_1 _09447_ (.A(_02059_),
    .B(_02102_),
    .Y(_02103_));
 sg13g2_a21oi_1 _09448_ (.A1(_02059_),
    .A2(_02098_),
    .Y(_02104_),
    .B1(_02103_));
 sg13g2_nand2_2 _09449_ (.Y(_02105_),
    .A(_02093_),
    .B(_02104_));
 sg13g2_inv_1 _09450_ (.Y(_02106_),
    .A(_02098_));
 sg13g2_a22oi_1 _09451_ (.Y(_02107_),
    .B1(\ppu.sprite_buffer.valid_sprites[0] ),
    .B2(_02051_),
    .A2(\ppu.sprite_buffer.valid_sprites[3] ),
    .A1(net263));
 sg13g2_buf_1 _09452_ (.A(_01927_),
    .X(_02108_));
 sg13g2_buf_1 _09453_ (.A(_01923_),
    .X(_02109_));
 sg13g2_a22oi_1 _09454_ (.Y(_02110_),
    .B1(\ppu.sprite_buffer.valid_sprites[2] ),
    .B2(net259),
    .A2(\ppu.sprite_buffer.valid_sprites[1] ),
    .A1(net252));
 sg13g2_nand2_1 _09455_ (.Y(_02111_),
    .A(_02107_),
    .B(_02110_));
 sg13g2_nand4_1 _09456_ (.B(_02080_),
    .C(_02091_),
    .A(_02062_),
    .Y(_02112_),
    .D(_02111_));
 sg13g2_a21oi_2 _09457_ (.B1(_02112_),
    .Y(_02113_),
    .A2(_02106_),
    .A1(_02058_));
 sg13g2_nand2_1 _09458_ (.Y(_02114_),
    .A(_02113_),
    .B(net254));
 sg13g2_nor3_1 _09459_ (.A(\ppu.sprite_buffer.sprite_catch_up_counters[3][0] ),
    .B(\ppu.sprite_buffer.sprite_catch_up_counters[3][1] ),
    .C(\ppu.sprite_buffer.sprite_catch_up_counters[3][2] ),
    .Y(_02115_));
 sg13g2_inv_1 _09460_ (.Y(_02116_),
    .A(_02115_));
 sg13g2_nand3_1 _09461_ (.B(_01910_),
    .C(_02116_),
    .A(_02114_),
    .Y(_02117_));
 sg13g2_nor2b_1 _09462_ (.A(_02117_),
    .B_N(_00127_),
    .Y(_02118_));
 sg13g2_nor2b_1 _09463_ (.A(_00127_),
    .B_N(_02117_),
    .Y(_02119_));
 sg13g2_o21ai_1 _09464_ (.B1(_01915_),
    .Y(_02120_),
    .A1(_02118_),
    .A2(_02119_));
 sg13g2_o21ai_1 _09465_ (.B1(_02120_),
    .Y(_00025_),
    .A1(_01915_),
    .A2(_02105_));
 sg13g2_xnor2_1 _09466_ (.Y(_02121_),
    .A(_02019_),
    .B(_02018_));
 sg13g2_inv_1 _09467_ (.Y(_02122_),
    .A(_02121_));
 sg13g2_nor2_1 _09468_ (.A(_02100_),
    .B(_02122_),
    .Y(_02123_));
 sg13g2_inv_1 _09469_ (.Y(_02124_),
    .A(_02123_));
 sg13g2_nand2_1 _09470_ (.Y(_02125_),
    .A(_02122_),
    .B(_02100_));
 sg13g2_and3_1 _09471_ (.X(_02126_),
    .A(_02124_),
    .B(net145),
    .C(_02125_));
 sg13g2_nor2b_1 _09472_ (.A(net145),
    .B_N(_02102_),
    .Y(_02127_));
 sg13g2_o21ai_1 _09473_ (.B1(_02093_),
    .Y(_02128_),
    .A1(_02126_),
    .A2(_02127_));
 sg13g2_buf_1 _09474_ (.A(_02128_),
    .X(_02129_));
 sg13g2_xor2_1 _09475_ (.B(_02118_),
    .A(\ppu.sprite_buffer.sprite_catch_up_counters[3][1] ),
    .X(_02130_));
 sg13g2_nand2_1 _09476_ (.Y(_02131_),
    .A(_02130_),
    .B(_01915_));
 sg13g2_o21ai_1 _09477_ (.B1(_02131_),
    .Y(_00026_),
    .A1(_01915_),
    .A2(_02129_));
 sg13g2_o21ai_1 _09478_ (.B1(_02124_),
    .Y(_02132_),
    .A1(net145),
    .A2(_02125_));
 sg13g2_a21o_1 _09479_ (.A2(_02026_),
    .A1(_02025_),
    .B1(_02059_),
    .X(_02133_));
 sg13g2_nor2_1 _09480_ (.A(_02123_),
    .B(_02133_),
    .Y(_02134_));
 sg13g2_a21oi_1 _09481_ (.A1(_02132_),
    .A2(_02133_),
    .Y(_02135_),
    .B1(_02134_));
 sg13g2_nand2_2 _09482_ (.Y(_02136_),
    .A(_02093_),
    .B(_02135_));
 sg13g2_nand2b_1 _09483_ (.Y(_02137_),
    .B(_02118_),
    .A_N(\ppu.sprite_buffer.sprite_catch_up_counters[3][1] ));
 sg13g2_xnor2_1 _09484_ (.Y(_02138_),
    .A(\ppu.sprite_buffer.sprite_catch_up_counters[3][2] ),
    .B(_02137_));
 sg13g2_nand2_1 _09485_ (.Y(_02139_),
    .A(_02138_),
    .B(_01915_));
 sg13g2_o21ai_1 _09486_ (.B1(_02139_),
    .Y(_00027_),
    .A1(_01915_),
    .A2(_02136_));
 sg13g2_buf_1 _09487_ (.A(net259),
    .X(_02140_));
 sg13g2_inv_1 _09488_ (.Y(_02141_),
    .A(_01909_));
 sg13g2_nand3_1 _09489_ (.B(_02141_),
    .C(\ppu.sprite_buffer.in_counters[2][2] ),
    .A(_01902_),
    .Y(_02142_));
 sg13g2_nor2_1 _09490_ (.A(_01908_),
    .B(_02142_),
    .Y(_02143_));
 sg13g2_a21oi_1 _09491_ (.A1(net251),
    .A2(_02143_),
    .Y(_02144_),
    .B1(_01912_));
 sg13g2_buf_1 _09492_ (.A(_02144_),
    .X(_02145_));
 sg13g2_nor3_1 _09493_ (.A(\ppu.sprite_buffer.sprite_catch_up_counters[2][0] ),
    .B(\ppu.sprite_buffer.sprite_catch_up_counters[2][1] ),
    .C(\ppu.sprite_buffer.sprite_catch_up_counters[2][2] ),
    .Y(_02146_));
 sg13g2_nand2_1 _09494_ (.Y(_02147_),
    .A(_02113_),
    .B(net259));
 sg13g2_nand3b_1 _09495_ (.B(_02147_),
    .C(_02142_),
    .Y(_02148_),
    .A_N(_02146_));
 sg13g2_nor2b_1 _09496_ (.A(_02148_),
    .B_N(_00128_),
    .Y(_02149_));
 sg13g2_nor2b_1 _09497_ (.A(_00128_),
    .B_N(_02148_),
    .Y(_02150_));
 sg13g2_o21ai_1 _09498_ (.B1(_02145_),
    .Y(_02151_),
    .A1(_02149_),
    .A2(_02150_));
 sg13g2_o21ai_1 _09499_ (.B1(_02151_),
    .Y(_00022_),
    .A1(_02105_),
    .A2(_02145_));
 sg13g2_xor2_1 _09500_ (.B(_02149_),
    .A(\ppu.sprite_buffer.sprite_catch_up_counters[2][1] ),
    .X(_02152_));
 sg13g2_nand2_1 _09501_ (.Y(_02153_),
    .A(_02152_),
    .B(_02145_));
 sg13g2_o21ai_1 _09502_ (.B1(_02153_),
    .Y(_00023_),
    .A1(_02129_),
    .A2(_02145_));
 sg13g2_nand2b_1 _09503_ (.Y(_02154_),
    .B(_02149_),
    .A_N(\ppu.sprite_buffer.sprite_catch_up_counters[2][1] ));
 sg13g2_xnor2_1 _09504_ (.Y(_02155_),
    .A(\ppu.sprite_buffer.sprite_catch_up_counters[2][2] ),
    .B(_02154_));
 sg13g2_nand2_1 _09505_ (.Y(_02156_),
    .A(_02155_),
    .B(_02145_));
 sg13g2_o21ai_1 _09506_ (.B1(_02156_),
    .Y(_00024_),
    .A1(_02136_),
    .A2(_02145_));
 sg13g2_inv_1 _09507_ (.Y(_02157_),
    .A(\ppu.sprite_buffer.in_counters[2][2] ));
 sg13g2_nand3_1 _09508_ (.B(_01909_),
    .C(_02157_),
    .A(_01902_),
    .Y(_02158_));
 sg13g2_nand2b_1 _09509_ (.Y(_02159_),
    .B(\ppu.sprite_buffer.final_pixels_in ),
    .A_N(_02158_));
 sg13g2_nor2_1 _09510_ (.A(_02042_),
    .B(_02159_),
    .Y(_02160_));
 sg13g2_nor2_1 _09511_ (.A(_02160_),
    .B(_01912_),
    .Y(_02161_));
 sg13g2_buf_1 _09512_ (.A(_02161_),
    .X(_02162_));
 sg13g2_nand2_1 _09513_ (.Y(_02163_),
    .A(_02113_),
    .B(net252));
 sg13g2_nor3_1 _09514_ (.A(\ppu.sprite_buffer.sprite_catch_up_counters[1][0] ),
    .B(\ppu.sprite_buffer.sprite_catch_up_counters[1][1] ),
    .C(\ppu.sprite_buffer.sprite_catch_up_counters[1][2] ),
    .Y(_02164_));
 sg13g2_inv_1 _09515_ (.Y(_02165_),
    .A(_02164_));
 sg13g2_nand3_1 _09516_ (.B(_02158_),
    .C(_02165_),
    .A(_02163_),
    .Y(_02166_));
 sg13g2_nor2b_1 _09517_ (.A(_02166_),
    .B_N(_00129_),
    .Y(_02167_));
 sg13g2_nor2b_1 _09518_ (.A(_00129_),
    .B_N(_02166_),
    .Y(_02168_));
 sg13g2_o21ai_1 _09519_ (.B1(_02162_),
    .Y(_02169_),
    .A1(_02167_),
    .A2(_02168_));
 sg13g2_o21ai_1 _09520_ (.B1(_02169_),
    .Y(_00019_),
    .A1(_02105_),
    .A2(_02162_));
 sg13g2_inv_1 _09521_ (.Y(_02170_),
    .A(\ppu.sprite_buffer.sprite_catch_up_counters[1][1] ));
 sg13g2_nor2_1 _09522_ (.A(_02170_),
    .B(_02167_),
    .Y(_02171_));
 sg13g2_nor2b_1 _09523_ (.A(\ppu.sprite_buffer.sprite_catch_up_counters[1][1] ),
    .B_N(_02167_),
    .Y(_02172_));
 sg13g2_o21ai_1 _09524_ (.B1(_02162_),
    .Y(_02173_),
    .A1(_02171_),
    .A2(_02172_));
 sg13g2_o21ai_1 _09525_ (.B1(_02173_),
    .Y(_00020_),
    .A1(_02129_),
    .A2(_02162_));
 sg13g2_a21o_1 _09526_ (.A2(_02170_),
    .A1(_02167_),
    .B1(\ppu.sprite_buffer.sprite_catch_up_counters[1][2] ),
    .X(_02174_));
 sg13g2_nand2_1 _09527_ (.Y(_02175_),
    .A(_02172_),
    .B(\ppu.sprite_buffer.sprite_catch_up_counters[1][2] ));
 sg13g2_nand3_1 _09528_ (.B(_02175_),
    .C(_02162_),
    .A(_02174_),
    .Y(_02176_));
 sg13g2_o21ai_1 _09529_ (.B1(_02176_),
    .Y(_00021_),
    .A1(_02136_),
    .A2(_02162_));
 sg13g2_nand3_1 _09530_ (.B(_02141_),
    .C(_02157_),
    .A(_01902_),
    .Y(_02177_));
 sg13g2_nand2b_1 _09531_ (.Y(_02178_),
    .B(\ppu.sprite_buffer.final_pixels_in ),
    .A_N(_02177_));
 sg13g2_nor2_1 _09532_ (.A(net262),
    .B(_02178_),
    .Y(_02179_));
 sg13g2_nor2_1 _09533_ (.A(_02179_),
    .B(_01912_),
    .Y(_02180_));
 sg13g2_buf_1 _09534_ (.A(_02180_),
    .X(_02181_));
 sg13g2_buf_1 _09535_ (.A(net253),
    .X(_02182_));
 sg13g2_nand2_1 _09536_ (.Y(_02183_),
    .A(_02113_),
    .B(net237));
 sg13g2_nor3_1 _09537_ (.A(\ppu.sprite_buffer.sprite_catch_up_counters[0][0] ),
    .B(\ppu.sprite_buffer.sprite_catch_up_counters[0][1] ),
    .C(\ppu.sprite_buffer.sprite_catch_up_counters[0][2] ),
    .Y(_02184_));
 sg13g2_inv_1 _09538_ (.Y(_02185_),
    .A(_02184_));
 sg13g2_nand3_1 _09539_ (.B(_02177_),
    .C(_02185_),
    .A(_02183_),
    .Y(_02186_));
 sg13g2_nor2b_1 _09540_ (.A(_02186_),
    .B_N(_00130_),
    .Y(_02187_));
 sg13g2_nor2b_1 _09541_ (.A(_00130_),
    .B_N(_02186_),
    .Y(_02188_));
 sg13g2_o21ai_1 _09542_ (.B1(_02181_),
    .Y(_02189_),
    .A1(_02187_),
    .A2(_02188_));
 sg13g2_o21ai_1 _09543_ (.B1(_02189_),
    .Y(_00016_),
    .A1(_02105_),
    .A2(_02181_));
 sg13g2_inv_1 _09544_ (.Y(_02190_),
    .A(\ppu.sprite_buffer.sprite_catch_up_counters[0][1] ));
 sg13g2_nor2_1 _09545_ (.A(_02190_),
    .B(_02187_),
    .Y(_02191_));
 sg13g2_nor2b_1 _09546_ (.A(\ppu.sprite_buffer.sprite_catch_up_counters[0][1] ),
    .B_N(_02187_),
    .Y(_02192_));
 sg13g2_o21ai_1 _09547_ (.B1(_02181_),
    .Y(_02193_),
    .A1(_02191_),
    .A2(_02192_));
 sg13g2_o21ai_1 _09548_ (.B1(_02193_),
    .Y(_00017_),
    .A1(_02129_),
    .A2(_02181_));
 sg13g2_a21o_1 _09549_ (.A2(_02190_),
    .A1(_02187_),
    .B1(\ppu.sprite_buffer.sprite_catch_up_counters[0][2] ),
    .X(_02194_));
 sg13g2_nand2_1 _09550_ (.Y(_02195_),
    .A(_02192_),
    .B(\ppu.sprite_buffer.sprite_catch_up_counters[0][2] ));
 sg13g2_nand3_1 _09551_ (.B(_02195_),
    .C(_02181_),
    .A(_02194_),
    .Y(_02196_));
 sg13g2_o21ai_1 _09552_ (.B1(_02196_),
    .Y(_00018_),
    .A1(_02136_),
    .A2(_02181_));
 sg13g2_buf_1 _09553_ (.A(net298),
    .X(_02197_));
 sg13g2_buf_1 _09554_ (.A(net258),
    .X(_02198_));
 sg13g2_nand2_2 _09555_ (.Y(_02199_),
    .A(_01850_),
    .B(net263));
 sg13g2_inv_1 _09556_ (.Y(_02200_),
    .A(_02199_));
 sg13g2_inv_1 _09557_ (.Y(_02201_),
    .A(\ppu.gfxmode1[0] ));
 sg13g2_nand2_1 _09558_ (.Y(_02202_),
    .A(_01802_),
    .B(\ppu.gfxmode2[0] ));
 sg13g2_o21ai_1 _09559_ (.B1(_02202_),
    .Y(_02203_),
    .A1(_01802_),
    .A2(_02201_));
 sg13g2_nor3_1 _09560_ (.A(_02095_),
    .B(net264),
    .C(_01850_),
    .Y(_02204_));
 sg13g2_a21oi_1 _09561_ (.A1(_02200_),
    .A2(_02203_),
    .Y(_02205_),
    .B1(_02204_));
 sg13g2_nor2_1 _09562_ (.A(net298),
    .B(net254),
    .Y(_02206_));
 sg13g2_buf_1 _09563_ (.A(_02206_),
    .X(_02207_));
 sg13g2_a22oi_1 _09564_ (.Y(_02208_),
    .B1(_02095_),
    .B2(_02207_),
    .A2(net258),
    .A1(\ppu.gfxmode1[0] ));
 sg13g2_o21ai_1 _09565_ (.B1(_02208_),
    .Y(_00011_),
    .A1(net250),
    .A2(_02205_));
 sg13g2_inv_2 _09566_ (.Y(_02209_),
    .A(net409));
 sg13g2_nor2_2 _09567_ (.A(_02209_),
    .B(net297),
    .Y(_02210_));
 sg13g2_xnor2_1 _09568_ (.Y(_02211_),
    .A(_01816_),
    .B(_02210_));
 sg13g2_inv_1 _09569_ (.Y(_02212_),
    .A(\ppu.gfxmode1[1] ));
 sg13g2_a21oi_1 _09570_ (.A1(net347),
    .A2(_02212_),
    .Y(_02213_),
    .B1(_01800_));
 sg13g2_o21ai_1 _09571_ (.B1(_02213_),
    .Y(_02214_),
    .A1(_01817_),
    .A2(\ppu.gfxmode2[1] ));
 sg13g2_nor2_1 _09572_ (.A(net298),
    .B(_02200_),
    .Y(_02215_));
 sg13g2_buf_2 _09573_ (.A(_02215_),
    .X(_02216_));
 sg13g2_inv_1 _09574_ (.Y(_02217_),
    .A(_02216_));
 sg13g2_a22oi_1 _09575_ (.Y(_02218_),
    .B1(_02214_),
    .B2(_02217_),
    .A2(_02211_),
    .A1(_02199_));
 sg13g2_a21o_1 _09576_ (.A2(net250),
    .A1(\ppu.gfxmode1[1] ),
    .B1(_02218_),
    .X(_00012_));
 sg13g2_inv_1 _09577_ (.Y(_02219_),
    .A(\ppu.gfxmode1[2] ));
 sg13g2_inv_1 _09578_ (.Y(_02220_),
    .A(net298));
 sg13g2_buf_1 _09579_ (.A(_02220_),
    .X(_02221_));
 sg13g2_nand2_1 _09580_ (.Y(_02222_),
    .A(_01802_),
    .B(\ppu.gfxmode2[2] ));
 sg13g2_nand2_1 _09581_ (.Y(_02223_),
    .A(net347),
    .B(\ppu.gfxmode1[2] ));
 sg13g2_a21oi_1 _09582_ (.A1(_02222_),
    .A2(_02223_),
    .Y(_02224_),
    .B1(net258));
 sg13g2_inv_1 _09583_ (.Y(_02225_),
    .A(_00033_));
 sg13g2_nand2_1 _09584_ (.Y(_02226_),
    .A(_02210_),
    .B(_02225_));
 sg13g2_xnor2_1 _09585_ (.Y(_02227_),
    .A(_01844_),
    .B(_02226_));
 sg13g2_nand2_1 _09586_ (.Y(_02228_),
    .A(_02199_),
    .B(_02227_));
 sg13g2_o21ai_1 _09587_ (.B1(_02228_),
    .Y(_02229_),
    .A1(_02224_),
    .A2(_02216_));
 sg13g2_o21ai_1 _09588_ (.B1(_02229_),
    .Y(_00013_),
    .A1(_02219_),
    .A2(net249));
 sg13g2_inv_1 _09589_ (.Y(_02230_),
    .A(\ppu.copper_inst.store[6] ));
 sg13g2_nor3_1 _09590_ (.A(_01859_),
    .B(_01860_),
    .C(_00031_),
    .Y(_02231_));
 sg13g2_nand2_1 _09591_ (.Y(_02232_),
    .A(_02231_),
    .B(\ppu.copper_inst.on ));
 sg13g2_nor2b_1 _09592_ (.A(_02232_),
    .B_N(_00076_),
    .Y(_02233_));
 sg13g2_buf_1 _09593_ (.A(net254),
    .X(_02234_));
 sg13g2_nand2_1 _09594_ (.Y(_02235_),
    .A(_02233_),
    .B(net236));
 sg13g2_buf_1 _09595_ (.A(_02235_),
    .X(_02236_));
 sg13g2_buf_1 _09596_ (.A(_00043_),
    .X(_02237_));
 sg13g2_inv_1 _09597_ (.Y(_02238_),
    .A(_02237_));
 sg13g2_buf_2 _09598_ (.A(\ppu.rs2.y_scan.counter[7] ),
    .X(_02239_));
 sg13g2_buf_2 _09599_ (.A(\ppu.rs2.y_scan.counter[6] ),
    .X(_02240_));
 sg13g2_buf_1 _09600_ (.A(\ppu.rs2.y_scan.counter[5] ),
    .X(_02241_));
 sg13g2_buf_2 _09601_ (.A(\ppu.rs2.y_scan.counter[4] ),
    .X(_02242_));
 sg13g2_buf_2 _09602_ (.A(\ppu.rs2.y_scan.counter[1] ),
    .X(_02243_));
 sg13g2_nor2_2 _09603_ (.A(_02243_),
    .B(_01865_),
    .Y(_02244_));
 sg13g2_buf_2 _09604_ (.A(\ppu.rs2.y_scan.counter[2] ),
    .X(_02245_));
 sg13g2_inv_2 _09605_ (.Y(_02246_),
    .A(_02245_));
 sg13g2_nand2_1 _09606_ (.Y(_02247_),
    .A(_02244_),
    .B(_02246_));
 sg13g2_nor2_1 _09607_ (.A(\ppu.rs2.y_scan.counter[3] ),
    .B(_02247_),
    .Y(_02248_));
 sg13g2_inv_1 _09608_ (.Y(_02249_),
    .A(_02248_));
 sg13g2_nor2_1 _09609_ (.A(_02242_),
    .B(_02249_),
    .Y(_02250_));
 sg13g2_inv_1 _09610_ (.Y(_02251_),
    .A(_02250_));
 sg13g2_nor2_1 _09611_ (.A(_02241_),
    .B(_02251_),
    .Y(_02252_));
 sg13g2_inv_1 _09612_ (.Y(_02253_),
    .A(_02252_));
 sg13g2_nor2_1 _09613_ (.A(_02240_),
    .B(_02253_),
    .Y(_02254_));
 sg13g2_inv_1 _09614_ (.Y(_02255_),
    .A(_02254_));
 sg13g2_nor2_1 _09615_ (.A(_02239_),
    .B(_02255_),
    .Y(_02256_));
 sg13g2_inv_1 _09616_ (.Y(_02257_),
    .A(_02256_));
 sg13g2_nor2_1 _09617_ (.A(_02238_),
    .B(_02257_),
    .Y(_02258_));
 sg13g2_buf_1 _09618_ (.A(_02258_),
    .X(_02259_));
 sg13g2_inv_1 _09619_ (.Y(_02260_),
    .A(net122));
 sg13g2_nor2_1 _09620_ (.A(_00180_),
    .B(_02199_),
    .Y(_02261_));
 sg13g2_inv_1 _09621_ (.Y(_02262_),
    .A(_02261_));
 sg13g2_nor2_2 _09622_ (.A(_02260_),
    .B(net184),
    .Y(_02263_));
 sg13g2_buf_1 _09623_ (.A(\ppu.rs2.phase_y[0] ),
    .X(_02264_));
 sg13g2_buf_2 _09624_ (.A(\ppu.rs2.phase_y[1] ),
    .X(_02265_));
 sg13g2_inv_1 _09625_ (.Y(_02266_),
    .A(_02265_));
 sg13g2_nor2_1 _09626_ (.A(_02264_),
    .B(_02266_),
    .Y(_02267_));
 sg13g2_nand2_1 _09627_ (.Y(_02268_),
    .A(_02263_),
    .B(_02267_));
 sg13g2_inv_1 _09628_ (.Y(_02269_),
    .A(_02268_));
 sg13g2_nor2_2 _09629_ (.A(net298),
    .B(_02269_),
    .Y(_02270_));
 sg13g2_nand3_1 _09630_ (.B(\ppu.copper_inst.fast_mode ),
    .C(_02236_),
    .A(_02270_),
    .Y(_02271_));
 sg13g2_o21ai_1 _09631_ (.B1(_02271_),
    .Y(_00014_),
    .A1(_02230_),
    .A2(_02236_));
 sg13g2_buf_1 _09632_ (.A(drive_uio_76),
    .X(_02272_));
 sg13g2_mux2_1 _09633_ (.A0(net8),
    .A1(net6),
    .S(_02272_),
    .X(_00001_));
 sg13g2_mux2_1 _09634_ (.A0(net9),
    .A1(net7),
    .S(_02272_),
    .X(_00002_));
 sg13g2_nor2_1 _09635_ (.A(\ppu.sync_delay[0] ),
    .B(\ppu.sync_delay[1] ),
    .Y(_02273_));
 sg13g2_inv_1 _09636_ (.Y(_02274_),
    .A(\ppu.sync_delay[2] ));
 sg13g2_a21oi_1 _09637_ (.A1(_02273_),
    .A2(_02274_),
    .Y(_02275_),
    .B1(net298));
 sg13g2_buf_2 _09638_ (.A(_02275_),
    .X(_02276_));
 sg13g2_inv_1 _09639_ (.Y(_02277_),
    .A(_00180_));
 sg13g2_nor2_1 _09640_ (.A(_01827_),
    .B(_02075_),
    .Y(_02278_));
 sg13g2_nor2_1 _09641_ (.A(_02277_),
    .B(_02278_),
    .Y(_02279_));
 sg13g2_xnor2_1 _09642_ (.Y(_02280_),
    .A(\ppu.gfxmode2[7] ),
    .B(_02279_));
 sg13g2_nand2_1 _09643_ (.Y(_02281_),
    .A(_02276_),
    .B(hsync));
 sg13g2_o21ai_1 _09644_ (.B1(_02281_),
    .Y(_00184_),
    .A1(_02276_),
    .A2(_02280_));
 sg13g2_xnor2_1 _09645_ (.Y(_02282_),
    .A(\ppu.gfxmode2[8] ),
    .B(\ppu.rs2.vsync0 ));
 sg13g2_nand2_1 _09646_ (.Y(_02283_),
    .A(_02276_),
    .B(\ppu.vsync ));
 sg13g2_o21ai_1 _09647_ (.B1(_02283_),
    .Y(_00185_),
    .A1(_02276_),
    .A2(_02282_));
 sg13g2_buf_1 _09648_ (.A(active),
    .X(_02284_));
 sg13g2_inv_1 _09649_ (.Y(_02285_),
    .A(_02284_));
 sg13g2_nor2_2 _09650_ (.A(_02265_),
    .B(net407),
    .Y(_02286_));
 sg13g2_inv_4 _09651_ (.A(_02286_),
    .Y(_02287_));
 sg13g2_nor3_2 _09652_ (.A(_01802_),
    .B(_02278_),
    .C(_02287_),
    .Y(_02288_));
 sg13g2_nor2_1 _09653_ (.A(_02276_),
    .B(_02288_),
    .Y(_02289_));
 sg13g2_a21oi_1 _09654_ (.A1(net389),
    .A2(_02276_),
    .Y(_00186_),
    .B1(_02289_));
 sg13g2_inv_1 _09655_ (.Y(_02290_),
    .A(\ppu.copper_inst.store[7] ));
 sg13g2_buf_1 _09656_ (.A(_02290_),
    .X(_02291_));
 sg13g2_buf_1 _09657_ (.A(\ppu.copper_inst.store[2] ),
    .X(_02292_));
 sg13g2_buf_1 _09658_ (.A(\ppu.copper_inst.store[3] ),
    .X(_02293_));
 sg13g2_inv_1 _09659_ (.Y(_02294_),
    .A(_02293_));
 sg13g2_a21oi_1 _09660_ (.A1(_01802_),
    .A2(_01830_),
    .Y(_02295_),
    .B1(_01811_));
 sg13g2_nor3_1 _09661_ (.A(_01801_),
    .B(_01831_),
    .C(_01812_),
    .Y(_02296_));
 sg13g2_buf_2 _09662_ (.A(\ppu.copper_inst.cmp_type ),
    .X(_02297_));
 sg13g2_inv_1 _09663_ (.Y(_02298_),
    .A(_02297_));
 sg13g2_buf_1 _09664_ (.A(_02298_),
    .X(_02299_));
 sg13g2_o21ai_1 _09665_ (.B1(net342),
    .Y(_02300_),
    .A1(_02295_),
    .A2(_02296_));
 sg13g2_o21ai_1 _09666_ (.B1(_02297_),
    .Y(_02301_),
    .A1(_02240_),
    .A2(_02287_));
 sg13g2_nand2_1 _09667_ (.Y(_02302_),
    .A(_02300_),
    .B(_02301_));
 sg13g2_nand2_1 _09668_ (.Y(_02303_),
    .A(_02302_),
    .B(\ppu.copper_inst.cmp[6] ));
 sg13g2_buf_1 _09669_ (.A(\ppu.copper_inst.cmp[5] ),
    .X(_02304_));
 sg13g2_xor2_1 _09670_ (.B(_01830_),
    .A(_01801_),
    .X(_02305_));
 sg13g2_buf_8 _09671_ (.A(_02286_),
    .X(_02306_));
 sg13g2_inv_1 _09672_ (.Y(_02307_),
    .A(_02241_));
 sg13g2_nand3_1 _09673_ (.B(_02297_),
    .C(_02307_),
    .A(net341),
    .Y(_02308_));
 sg13g2_o21ai_1 _09674_ (.B1(_02308_),
    .Y(_02309_),
    .A1(_02297_),
    .A2(_02305_));
 sg13g2_nor2b_1 _09675_ (.A(_02304_),
    .B_N(_02309_),
    .Y(_02310_));
 sg13g2_nand2_1 _09676_ (.Y(_02311_),
    .A(_02303_),
    .B(_02310_));
 sg13g2_inv_1 _09677_ (.Y(_02312_),
    .A(\ppu.copper_inst.cmp[6] ));
 sg13g2_nand3_1 _09678_ (.B(_02312_),
    .C(_02301_),
    .A(_02300_),
    .Y(_02313_));
 sg13g2_nand2_1 _09679_ (.Y(_02314_),
    .A(_02311_),
    .B(_02313_));
 sg13g2_buf_1 _09680_ (.A(\ppu.copper_inst.cmp[7] ),
    .X(_02315_));
 sg13g2_nor2_1 _09681_ (.A(_02239_),
    .B(net342),
    .Y(_02316_));
 sg13g2_nand2_1 _09682_ (.Y(_02317_),
    .A(_01801_),
    .B(_02075_));
 sg13g2_inv_1 _09683_ (.Y(_02318_),
    .A(_02317_));
 sg13g2_a22oi_1 _09684_ (.Y(_02319_),
    .B1(net342),
    .B2(_02318_),
    .A2(net341),
    .A1(_02316_));
 sg13g2_xnor2_1 _09685_ (.Y(_02320_),
    .A(_02315_),
    .B(_02319_));
 sg13g2_buf_2 _09686_ (.A(\ppu.rs2.y_scan.counter[8] ),
    .X(_02321_));
 sg13g2_nor2_1 _09687_ (.A(_02321_),
    .B(_02298_),
    .Y(_02322_));
 sg13g2_nand2_1 _09688_ (.Y(_02323_),
    .A(_02322_),
    .B(_02286_));
 sg13g2_o21ai_1 _09689_ (.B1(_02323_),
    .Y(_02324_),
    .A1(_02297_),
    .A2(_00040_));
 sg13g2_or2_1 _09690_ (.X(_02325_),
    .B(_02324_),
    .A(_00039_));
 sg13g2_nand2_1 _09691_ (.Y(_02326_),
    .A(_02324_),
    .B(_00039_));
 sg13g2_nand2_1 _09692_ (.Y(_02327_),
    .A(_02325_),
    .B(_02326_));
 sg13g2_nor2_1 _09693_ (.A(_02320_),
    .B(_02327_),
    .Y(_02328_));
 sg13g2_nand2_1 _09694_ (.Y(_02329_),
    .A(_02314_),
    .B(_02328_));
 sg13g2_o21ai_1 _09695_ (.B1(_02326_),
    .Y(_02330_),
    .A1(_02315_),
    .A2(_02319_));
 sg13g2_nand2_1 _09696_ (.Y(_02331_),
    .A(_02330_),
    .B(_02325_));
 sg13g2_nand2_1 _09697_ (.Y(_02332_),
    .A(_02329_),
    .B(_02331_));
 sg13g2_nand3_1 _09698_ (.B(_02297_),
    .C(_02246_),
    .A(net341),
    .Y(_02333_));
 sg13g2_nand2_1 _09699_ (.Y(_02334_),
    .A(_01957_),
    .B(net342));
 sg13g2_nand3_1 _09700_ (.B(\ppu.copper_inst.cmp[2] ),
    .C(_02334_),
    .A(_02333_),
    .Y(_02335_));
 sg13g2_nor2_1 _09701_ (.A(_02243_),
    .B(net342),
    .Y(_02336_));
 sg13g2_nand2_1 _09702_ (.Y(_02337_),
    .A(_02336_),
    .B(net341));
 sg13g2_nand2_1 _09703_ (.Y(_02338_),
    .A(_02225_),
    .B(_02299_));
 sg13g2_a21oi_1 _09704_ (.A1(_02337_),
    .A2(_02338_),
    .Y(_02339_),
    .B1(\ppu.copper_inst.cmp[1] ));
 sg13g2_a21oi_1 _09705_ (.A1(_02333_),
    .A2(_02334_),
    .Y(_02340_),
    .B1(\ppu.copper_inst.cmp[2] ));
 sg13g2_a21oi_1 _09706_ (.A1(_02335_),
    .A2(_02339_),
    .Y(_02341_),
    .B1(_02340_));
 sg13g2_inv_2 _09707_ (.Y(_02342_),
    .A(\ppu.rs2.y_scan.counter[3] ));
 sg13g2_nand3_1 _09708_ (.B(_02297_),
    .C(_02342_),
    .A(_02286_),
    .Y(_02343_));
 sg13g2_nand2b_1 _09709_ (.Y(_02344_),
    .B(net342),
    .A_N(_00037_));
 sg13g2_a21oi_1 _09710_ (.A1(_02343_),
    .A2(_02344_),
    .Y(_02345_),
    .B1(\ppu.copper_inst.cmp[3] ));
 sg13g2_nand3_1 _09711_ (.B(\ppu.copper_inst.cmp[3] ),
    .C(_02344_),
    .A(_02343_),
    .Y(_02346_));
 sg13g2_nor2b_1 _09712_ (.A(_02345_),
    .B_N(_02346_),
    .Y(_02347_));
 sg13g2_buf_1 _09713_ (.A(\ppu.copper_inst.cmp[4] ),
    .X(_02348_));
 sg13g2_inv_1 _09714_ (.Y(_02349_),
    .A(_00038_));
 sg13g2_nor2_1 _09715_ (.A(_02242_),
    .B(_02298_),
    .Y(_02350_));
 sg13g2_a22oi_1 _09716_ (.Y(_02351_),
    .B1(_02306_),
    .B2(_02350_),
    .A2(_02349_),
    .A1(_02299_));
 sg13g2_xor2_1 _09717_ (.B(_02351_),
    .A(_02348_),
    .X(_02352_));
 sg13g2_nand2_1 _09718_ (.Y(_02353_),
    .A(_02347_),
    .B(_02352_));
 sg13g2_nor2_1 _09719_ (.A(_02341_),
    .B(_02353_),
    .Y(_02354_));
 sg13g2_nand2_1 _09720_ (.Y(_02355_),
    .A(_02351_),
    .B(_02348_));
 sg13g2_nor2_1 _09721_ (.A(_02348_),
    .B(_02351_),
    .Y(_02356_));
 sg13g2_a21oi_1 _09722_ (.A1(_02345_),
    .A2(_02355_),
    .Y(_02357_),
    .B1(_02356_));
 sg13g2_nor2b_1 _09723_ (.A(_02354_),
    .B_N(_02357_),
    .Y(_02358_));
 sg13g2_xor2_1 _09724_ (.B(_02309_),
    .A(_02304_),
    .X(_02359_));
 sg13g2_nand2_1 _09725_ (.Y(_02360_),
    .A(_02303_),
    .B(_02313_));
 sg13g2_nor2_1 _09726_ (.A(_02359_),
    .B(_02360_),
    .Y(_02361_));
 sg13g2_nand2_1 _09727_ (.Y(_02362_),
    .A(_02361_),
    .B(_02328_));
 sg13g2_nor2_1 _09728_ (.A(_02358_),
    .B(_02362_),
    .Y(_02363_));
 sg13g2_nor2_1 _09729_ (.A(_02332_),
    .B(_02363_),
    .Y(_02364_));
 sg13g2_nor2b_1 _09730_ (.A(_02340_),
    .B_N(_02335_),
    .Y(_02365_));
 sg13g2_nand3_1 _09731_ (.B(\ppu.copper_inst.cmp[1] ),
    .C(_02338_),
    .A(_02337_),
    .Y(_02366_));
 sg13g2_nor2b_1 _09732_ (.A(_02339_),
    .B_N(_02366_),
    .Y(_02367_));
 sg13g2_nand2_1 _09733_ (.Y(_02368_),
    .A(_02365_),
    .B(_02367_));
 sg13g2_nor2_1 _09734_ (.A(_02368_),
    .B(_02353_),
    .Y(_02369_));
 sg13g2_nand3_1 _09735_ (.B(_00036_),
    .C(_02297_),
    .A(net341),
    .Y(_02370_));
 sg13g2_nand2_1 _09736_ (.Y(_02371_),
    .A(net342),
    .B(net409));
 sg13g2_nand3_1 _09737_ (.B(\ppu.copper_inst.cmp[0] ),
    .C(_02371_),
    .A(_02370_),
    .Y(_02372_));
 sg13g2_nand4_1 _09738_ (.B(_02369_),
    .C(_02372_),
    .A(_02361_),
    .Y(_02373_),
    .D(_02328_));
 sg13g2_nand3_1 _09739_ (.B(\ppu.copper_inst.cmp_on ),
    .C(_02373_),
    .A(_02364_),
    .Y(_02374_));
 sg13g2_nand2_1 _09740_ (.Y(_02375_),
    .A(\ppu.copper_inst.on ),
    .B(\ppu.copper_inst.store_valid ));
 sg13g2_inv_1 _09741_ (.Y(_02376_),
    .A(_02375_));
 sg13g2_nand2_1 _09742_ (.Y(_02377_),
    .A(_02374_),
    .B(_02376_));
 sg13g2_nor2_2 _09743_ (.A(net297),
    .B(_02377_),
    .Y(_02378_));
 sg13g2_inv_2 _09744_ (.Y(_02379_),
    .A(_02378_));
 sg13g2_nor3_2 _09745_ (.A(_02292_),
    .B(_02294_),
    .C(_02379_),
    .Y(_02380_));
 sg13g2_buf_1 _09746_ (.A(\ppu.copper_inst.store[1] ),
    .X(_02381_));
 sg13g2_inv_1 _09747_ (.Y(_02382_),
    .A(_02381_));
 sg13g2_buf_1 _09748_ (.A(\ppu.copper_inst.store[0] ),
    .X(_02383_));
 sg13g2_inv_1 _09749_ (.Y(_02384_),
    .A(_02383_));
 sg13g2_inv_1 _09750_ (.Y(_02385_),
    .A(\ppu.copper_inst.store[4] ));
 sg13g2_nor2_1 _09751_ (.A(\ppu.copper_inst.store[5] ),
    .B(_02385_),
    .Y(_02386_));
 sg13g2_buf_2 _09752_ (.A(_02386_),
    .X(_02387_));
 sg13g2_nand4_1 _09753_ (.B(_02382_),
    .C(_02384_),
    .A(_02380_),
    .Y(_02388_),
    .D(_02387_));
 sg13g2_buf_1 _09754_ (.A(_02388_),
    .X(_02389_));
 sg13g2_buf_1 _09755_ (.A(net108),
    .X(_02390_));
 sg13g2_nand2_1 _09756_ (.Y(_02391_),
    .A(net102),
    .B(\ppu.base_addr_regs[0][0] ));
 sg13g2_o21ai_1 _09757_ (.B1(_02391_),
    .Y(_00187_),
    .A1(_02291_),
    .A2(net102));
 sg13g2_buf_1 _09758_ (.A(\ppu.copper_inst.store[8] ),
    .X(_02392_));
 sg13g2_inv_1 _09759_ (.Y(_02393_),
    .A(_02392_));
 sg13g2_buf_1 _09760_ (.A(_02393_),
    .X(_02394_));
 sg13g2_nand2_1 _09761_ (.Y(_02395_),
    .A(net108),
    .B(\ppu.base_addr_regs[0][1] ));
 sg13g2_o21ai_1 _09762_ (.B1(_02395_),
    .Y(_00188_),
    .A1(net340),
    .A2(net102));
 sg13g2_buf_2 _09763_ (.A(\ppu.copper_inst.store[9] ),
    .X(_02396_));
 sg13g2_inv_1 _09764_ (.Y(_02397_),
    .A(_02396_));
 sg13g2_buf_1 _09765_ (.A(_02397_),
    .X(_02398_));
 sg13g2_nand2_1 _09766_ (.Y(_02399_),
    .A(net108),
    .B(\ppu.base_addr_regs[0][2] ));
 sg13g2_o21ai_1 _09767_ (.B1(_02399_),
    .Y(_00189_),
    .A1(net339),
    .A2(net102));
 sg13g2_buf_1 _09768_ (.A(\ppu.copper_inst.store[10] ),
    .X(_02400_));
 sg13g2_inv_1 _09769_ (.Y(_02401_),
    .A(_02400_));
 sg13g2_buf_1 _09770_ (.A(_02401_),
    .X(_02402_));
 sg13g2_nand2_1 _09771_ (.Y(_02403_),
    .A(net108),
    .B(\ppu.base_addr_regs[0][3] ));
 sg13g2_o21ai_1 _09772_ (.B1(_02403_),
    .Y(_00190_),
    .A1(_02402_),
    .A2(net102));
 sg13g2_buf_1 _09773_ (.A(\ppu.copper_inst.store[11] ),
    .X(_02404_));
 sg13g2_inv_1 _09774_ (.Y(_02405_),
    .A(_02404_));
 sg13g2_buf_1 _09775_ (.A(_02405_),
    .X(_02406_));
 sg13g2_nand2_1 _09776_ (.Y(_02407_),
    .A(net108),
    .B(\ppu.base_addr_regs[0][4] ));
 sg13g2_o21ai_1 _09777_ (.B1(_02407_),
    .Y(_00191_),
    .A1(net337),
    .A2(net102));
 sg13g2_buf_2 _09778_ (.A(\ppu.copper_inst.store[12] ),
    .X(_02408_));
 sg13g2_inv_1 _09779_ (.Y(_02409_),
    .A(_02408_));
 sg13g2_nand2_1 _09780_ (.Y(_02410_),
    .A(net108),
    .B(\ppu.base_addr_regs[0][5] ));
 sg13g2_o21ai_1 _09781_ (.B1(_02410_),
    .Y(_00192_),
    .A1(net387),
    .A2(net102));
 sg13g2_buf_1 _09782_ (.A(\ppu.copper_inst.store[13] ),
    .X(_02411_));
 sg13g2_inv_2 _09783_ (.Y(_02412_),
    .A(net406));
 sg13g2_nand2_1 _09784_ (.Y(_02413_),
    .A(net108),
    .B(\ppu.base_addr_regs[0][6] ));
 sg13g2_o21ai_1 _09785_ (.B1(_02413_),
    .Y(_00193_),
    .A1(_02412_),
    .A2(net102));
 sg13g2_buf_1 _09786_ (.A(\ppu.copper_inst.store[14] ),
    .X(_02414_));
 sg13g2_inv_1 _09787_ (.Y(_02415_),
    .A(_02414_));
 sg13g2_nand2_1 _09788_ (.Y(_02416_),
    .A(_02389_),
    .B(\ppu.base_addr_regs[0][7] ));
 sg13g2_o21ai_1 _09789_ (.B1(_02416_),
    .Y(_00194_),
    .A1(_02415_),
    .A2(_02390_));
 sg13g2_buf_1 _09790_ (.A(\ppu.copper_inst.store[15] ),
    .X(_02417_));
 sg13g2_inv_1 _09791_ (.Y(_02418_),
    .A(_02417_));
 sg13g2_nand2_1 _09792_ (.Y(_02419_),
    .A(net108),
    .B(\ppu.base_addr_regs[0][8] ));
 sg13g2_o21ai_1 _09793_ (.B1(_02419_),
    .Y(_00195_),
    .A1(net385),
    .A2(_02390_));
 sg13g2_inv_1 _09794_ (.Y(_02420_),
    .A(_02387_));
 sg13g2_inv_1 _09795_ (.Y(_02421_),
    .A(_02380_));
 sg13g2_nor4_1 _09796_ (.A(_02381_),
    .B(_02384_),
    .C(_02420_),
    .D(_02421_),
    .Y(_02422_));
 sg13g2_buf_1 _09797_ (.A(_02422_),
    .X(_02423_));
 sg13g2_buf_1 _09798_ (.A(net101),
    .X(_02424_));
 sg13g2_nor2_1 _09799_ (.A(\ppu.base_addr_regs[1][0] ),
    .B(net91),
    .Y(_02425_));
 sg13g2_a21oi_1 _09800_ (.A1(_02291_),
    .A2(net91),
    .Y(_00196_),
    .B1(_02425_));
 sg13g2_nor2_1 _09801_ (.A(\ppu.base_addr_regs[1][1] ),
    .B(net101),
    .Y(_02426_));
 sg13g2_a21oi_1 _09802_ (.A1(_02394_),
    .A2(net91),
    .Y(_00197_),
    .B1(_02426_));
 sg13g2_nor2_1 _09803_ (.A(\ppu.base_addr_regs[1][2] ),
    .B(net101),
    .Y(_02427_));
 sg13g2_a21oi_1 _09804_ (.A1(_02398_),
    .A2(net91),
    .Y(_00198_),
    .B1(_02427_));
 sg13g2_nor2_1 _09805_ (.A(\ppu.base_addr_regs[1][3] ),
    .B(net101),
    .Y(_02428_));
 sg13g2_a21oi_1 _09806_ (.A1(net338),
    .A2(net91),
    .Y(_00199_),
    .B1(_02428_));
 sg13g2_nor2_1 _09807_ (.A(\ppu.base_addr_regs[1][4] ),
    .B(_02423_),
    .Y(_02429_));
 sg13g2_a21oi_1 _09808_ (.A1(_02406_),
    .A2(_02424_),
    .Y(_00200_),
    .B1(_02429_));
 sg13g2_nor2_1 _09809_ (.A(\ppu.base_addr_regs[1][5] ),
    .B(net101),
    .Y(_02430_));
 sg13g2_a21oi_1 _09810_ (.A1(net387),
    .A2(net91),
    .Y(_00201_),
    .B1(_02430_));
 sg13g2_nor2_1 _09811_ (.A(\ppu.base_addr_regs[1][6] ),
    .B(net101),
    .Y(_02431_));
 sg13g2_a21oi_1 _09812_ (.A1(_02412_),
    .A2(net91),
    .Y(_00202_),
    .B1(_02431_));
 sg13g2_nor2_1 _09813_ (.A(\ppu.base_addr_regs[1][7] ),
    .B(net101),
    .Y(_02432_));
 sg13g2_a21oi_1 _09814_ (.A1(net386),
    .A2(_02424_),
    .Y(_00203_),
    .B1(_02432_));
 sg13g2_nor2_1 _09815_ (.A(\ppu.base_addr_regs[1][8] ),
    .B(net101),
    .Y(_02433_));
 sg13g2_a21oi_1 _09816_ (.A1(_02418_),
    .A2(net91),
    .Y(_00204_),
    .B1(_02433_));
 sg13g2_nor2_1 _09817_ (.A(_02383_),
    .B(_02382_),
    .Y(_02434_));
 sg13g2_nand3_1 _09818_ (.B(_02387_),
    .C(_02434_),
    .A(_02380_),
    .Y(_02435_));
 sg13g2_buf_1 _09819_ (.A(_02435_),
    .X(_02436_));
 sg13g2_buf_1 _09820_ (.A(_02436_),
    .X(_02437_));
 sg13g2_nand2_1 _09821_ (.Y(_02438_),
    .A(net100),
    .B(\ppu.base_addr_regs[2][1] ));
 sg13g2_o21ai_1 _09822_ (.B1(_02438_),
    .Y(_00205_),
    .A1(net340),
    .A2(net100));
 sg13g2_nand2_1 _09823_ (.Y(_02439_),
    .A(_02437_),
    .B(\ppu.base_addr_regs[2][2] ));
 sg13g2_o21ai_1 _09824_ (.B1(_02439_),
    .Y(_00206_),
    .A1(net339),
    .A2(_02437_));
 sg13g2_inv_1 _09825_ (.Y(_02440_),
    .A(\ppu.base_addr_regs[2][3] ));
 sg13g2_nor2_1 _09826_ (.A(_02400_),
    .B(_02436_),
    .Y(_02441_));
 sg13g2_a21oi_1 _09827_ (.A1(_02440_),
    .A2(net100),
    .Y(_00207_),
    .B1(_02441_));
 sg13g2_inv_1 _09828_ (.Y(_02442_),
    .A(\ppu.base_addr_regs[2][4] ));
 sg13g2_nor2_1 _09829_ (.A(_02404_),
    .B(_02436_),
    .Y(_02443_));
 sg13g2_a21oi_1 _09830_ (.A1(_02442_),
    .A2(net100),
    .Y(_00208_),
    .B1(_02443_));
 sg13g2_inv_1 _09831_ (.Y(_02444_),
    .A(\ppu.base_addr_regs[2][5] ));
 sg13g2_nor2_1 _09832_ (.A(_02408_),
    .B(_02436_),
    .Y(_02445_));
 sg13g2_a21oi_1 _09833_ (.A1(_02444_),
    .A2(net100),
    .Y(_00209_),
    .B1(_02445_));
 sg13g2_inv_1 _09834_ (.Y(_02446_),
    .A(\ppu.base_addr_regs[2][6] ));
 sg13g2_nor2_1 _09835_ (.A(net406),
    .B(_02436_),
    .Y(_02447_));
 sg13g2_a21oi_1 _09836_ (.A1(_02446_),
    .A2(net100),
    .Y(_00210_),
    .B1(_02447_));
 sg13g2_nand2_1 _09837_ (.Y(_02448_),
    .A(_02436_),
    .B(\ppu.base_addr_regs[2][7] ));
 sg13g2_o21ai_1 _09838_ (.B1(_02448_),
    .Y(_00211_),
    .A1(net386),
    .A2(net100));
 sg13g2_nand2_1 _09839_ (.Y(_02449_),
    .A(_02436_),
    .B(\ppu.base_addr_regs[2][8] ));
 sg13g2_o21ai_1 _09840_ (.B1(_02449_),
    .Y(_00212_),
    .A1(net385),
    .A2(net100));
 sg13g2_inv_1 _09841_ (.Y(_02450_),
    .A(\ppu.base_addr_regs[3][1] ));
 sg13g2_nand2_1 _09842_ (.Y(_02451_),
    .A(_02381_),
    .B(_02383_));
 sg13g2_inv_1 _09843_ (.Y(_02452_),
    .A(_02451_));
 sg13g2_nand3_1 _09844_ (.B(_02387_),
    .C(_02452_),
    .A(_02380_),
    .Y(_02453_));
 sg13g2_buf_2 _09845_ (.A(_02453_),
    .X(_02454_));
 sg13g2_nor2_1 _09846_ (.A(_02392_),
    .B(_02454_),
    .Y(_02455_));
 sg13g2_a21oi_1 _09847_ (.A1(_02450_),
    .A2(_02454_),
    .Y(_00213_),
    .B1(_02455_));
 sg13g2_inv_1 _09848_ (.Y(_02456_),
    .A(\ppu.base_addr_regs[3][2] ));
 sg13g2_nor2_1 _09849_ (.A(_02396_),
    .B(_02454_),
    .Y(_02457_));
 sg13g2_a21oi_1 _09850_ (.A1(_02456_),
    .A2(_02454_),
    .Y(_00214_),
    .B1(_02457_));
 sg13g2_nand2_1 _09851_ (.Y(_02458_),
    .A(_02454_),
    .B(\ppu.base_addr_regs[3][3] ));
 sg13g2_o21ai_1 _09852_ (.B1(_02458_),
    .Y(_00215_),
    .A1(_02402_),
    .A2(_02454_));
 sg13g2_nand2_1 _09853_ (.Y(_02459_),
    .A(_02454_),
    .B(\ppu.base_addr_regs[3][4] ));
 sg13g2_o21ai_1 _09854_ (.B1(_02459_),
    .Y(_00216_),
    .A1(net337),
    .A2(_02454_));
 sg13g2_inv_1 _09855_ (.Y(_02460_),
    .A(_02292_));
 sg13g2_nor4_2 _09856_ (.A(_02460_),
    .B(_02293_),
    .C(_02420_),
    .Y(_02461_),
    .D(_02379_));
 sg13g2_nand2_1 _09857_ (.Y(_02462_),
    .A(_02461_),
    .B(_02451_));
 sg13g2_buf_1 _09858_ (.A(_02462_),
    .X(_02463_));
 sg13g2_buf_1 _09859_ (.A(net107),
    .X(_02464_));
 sg13g2_nand2_1 _09860_ (.Y(_02465_),
    .A(net99),
    .B(\ppu.copper_inst.cmp[0] ));
 sg13g2_o21ai_1 _09861_ (.B1(_02465_),
    .Y(_00233_),
    .A1(net388),
    .A2(net99));
 sg13g2_nand2_1 _09862_ (.Y(_02466_),
    .A(net107),
    .B(\ppu.copper_inst.cmp[1] ));
 sg13g2_o21ai_1 _09863_ (.B1(_02466_),
    .Y(_00234_),
    .A1(net340),
    .A2(net99));
 sg13g2_nand2_1 _09864_ (.Y(_02467_),
    .A(_02463_),
    .B(\ppu.copper_inst.cmp[2] ));
 sg13g2_o21ai_1 _09865_ (.B1(_02467_),
    .Y(_00235_),
    .A1(net339),
    .A2(_02464_));
 sg13g2_nand2_1 _09866_ (.Y(_02468_),
    .A(net107),
    .B(\ppu.copper_inst.cmp[3] ));
 sg13g2_o21ai_1 _09867_ (.B1(_02468_),
    .Y(_00236_),
    .A1(net338),
    .A2(net99));
 sg13g2_nand2_1 _09868_ (.Y(_02469_),
    .A(net107),
    .B(_02348_));
 sg13g2_o21ai_1 _09869_ (.B1(_02469_),
    .Y(_00237_),
    .A1(net337),
    .A2(net99));
 sg13g2_nand2_1 _09870_ (.Y(_02470_),
    .A(net107),
    .B(_02304_));
 sg13g2_o21ai_1 _09871_ (.B1(_02470_),
    .Y(_00238_),
    .A1(_02409_),
    .A2(net99));
 sg13g2_nor2_1 _09872_ (.A(net406),
    .B(net107),
    .Y(_02471_));
 sg13g2_a21oi_1 _09873_ (.A1(_02312_),
    .A2(net99),
    .Y(_00239_),
    .B1(_02471_));
 sg13g2_nand2_1 _09874_ (.Y(_02472_),
    .A(net107),
    .B(_02315_));
 sg13g2_o21ai_1 _09875_ (.B1(_02472_),
    .Y(_00240_),
    .A1(net386),
    .A2(net99));
 sg13g2_nand2_1 _09876_ (.Y(_02473_),
    .A(net107),
    .B(\ppu.copper_inst.cmp[8] ));
 sg13g2_o21ai_1 _09877_ (.B1(_02473_),
    .Y(_00241_),
    .A1(_02418_),
    .A2(_02464_));
 sg13g2_nand2_1 _09878_ (.Y(_02474_),
    .A(_02270_),
    .B(_02378_));
 sg13g2_nor2_1 _09879_ (.A(_02383_),
    .B(_02474_),
    .Y(_02475_));
 sg13g2_a21oi_1 _09880_ (.A1(net342),
    .A2(_02474_),
    .Y(_00243_),
    .B1(_02475_));
 sg13g2_nand2_1 _09881_ (.Y(_02476_),
    .A(_02292_),
    .B(_02293_));
 sg13g2_inv_1 _09882_ (.Y(_02477_),
    .A(_02476_));
 sg13g2_nand2_1 _09883_ (.Y(_02478_),
    .A(_02452_),
    .B(_02477_));
 sg13g2_nand4_1 _09884_ (.B(\ppu.copper_inst.store_valid ),
    .C(\ppu.copper_inst.store[5] ),
    .A(net236),
    .Y(_02479_),
    .D(\ppu.copper_inst.store[4] ));
 sg13g2_o21ai_1 _09885_ (.B1(\ppu.copper_inst.on ),
    .Y(_02480_),
    .A1(_02478_),
    .A2(_02479_));
 sg13g2_nand2_1 _09886_ (.Y(_00244_),
    .A(_02270_),
    .B(_02480_));
 sg13g2_buf_1 _09887_ (.A(net237),
    .X(_02481_));
 sg13g2_nand2_1 _09888_ (.Y(_02482_),
    .A(_02233_),
    .B(net216));
 sg13g2_buf_2 _09889_ (.A(_02482_),
    .X(_02483_));
 sg13g2_buf_1 _09890_ (.A(\data_pins[0] ),
    .X(_02484_));
 sg13g2_buf_1 _09891_ (.A(_02484_),
    .X(_02485_));
 sg13g2_nor2_1 _09892_ (.A(net384),
    .B(_02483_),
    .Y(_02486_));
 sg13g2_a21oi_1 _09893_ (.A1(_02384_),
    .A2(_02483_),
    .Y(_00245_),
    .B1(_02486_));
 sg13g2_nand2_1 _09894_ (.Y(_02487_),
    .A(_02233_),
    .B(net251));
 sg13g2_buf_2 _09895_ (.A(_02487_),
    .X(_02488_));
 sg13g2_buf_1 _09896_ (.A(\data_pins[2] ),
    .X(_02489_));
 sg13g2_nor2_1 _09897_ (.A(net404),
    .B(_02488_),
    .Y(_02490_));
 sg13g2_a21oi_1 _09898_ (.A1(net338),
    .A2(_02488_),
    .Y(_00246_),
    .B1(_02490_));
 sg13g2_nor2_1 _09899_ (.A(net408),
    .B(_02488_),
    .Y(_02491_));
 sg13g2_a21oi_1 _09900_ (.A1(net337),
    .A2(_02488_),
    .Y(_00247_),
    .B1(_02491_));
 sg13g2_nor2_1 _09901_ (.A(net384),
    .B(net200),
    .Y(_02492_));
 sg13g2_a21oi_1 _09902_ (.A1(net387),
    .A2(net200),
    .Y(_00248_),
    .B1(_02492_));
 sg13g2_buf_1 _09903_ (.A(\data_pins[1] ),
    .X(_02493_));
 sg13g2_buf_1 _09904_ (.A(net403),
    .X(_02494_));
 sg13g2_nor2_1 _09905_ (.A(net383),
    .B(net200),
    .Y(_02495_));
 sg13g2_a21oi_1 _09906_ (.A1(_02412_),
    .A2(net200),
    .Y(_00249_),
    .B1(_02495_));
 sg13g2_nor2_1 _09907_ (.A(net404),
    .B(net200),
    .Y(_02496_));
 sg13g2_a21oi_1 _09908_ (.A1(_02415_),
    .A2(net200),
    .Y(_00250_),
    .B1(_02496_));
 sg13g2_nor2_1 _09909_ (.A(net408),
    .B(net200),
    .Y(_02497_));
 sg13g2_a21oi_1 _09910_ (.A1(net385),
    .A2(net200),
    .Y(_00251_),
    .B1(_02497_));
 sg13g2_nor2_1 _09911_ (.A(net383),
    .B(_02483_),
    .Y(_02498_));
 sg13g2_a21oi_1 _09912_ (.A1(_02382_),
    .A2(_02483_),
    .Y(_00252_),
    .B1(_02498_));
 sg13g2_nor2_1 _09913_ (.A(net404),
    .B(_02483_),
    .Y(_02499_));
 sg13g2_a21oi_1 _09914_ (.A1(_02460_),
    .A2(_02483_),
    .Y(_00253_),
    .B1(_02499_));
 sg13g2_nor2_1 _09915_ (.A(net408),
    .B(_02483_),
    .Y(_02500_));
 sg13g2_a21oi_1 _09916_ (.A1(_02294_),
    .A2(_02483_),
    .Y(_00254_),
    .B1(_02500_));
 sg13g2_buf_1 _09917_ (.A(net252),
    .X(_02501_));
 sg13g2_nand2_1 _09918_ (.Y(_02502_),
    .A(_02233_),
    .B(net235));
 sg13g2_buf_2 _09919_ (.A(_02502_),
    .X(_02503_));
 sg13g2_nor2_1 _09920_ (.A(net384),
    .B(_02503_),
    .Y(_02504_));
 sg13g2_a21oi_1 _09921_ (.A1(_02385_),
    .A2(_02503_),
    .Y(_00255_),
    .B1(_02504_));
 sg13g2_inv_1 _09922_ (.Y(_02505_),
    .A(net403));
 sg13g2_nand2_1 _09923_ (.Y(_02506_),
    .A(_02503_),
    .B(\ppu.copper_inst.store[5] ));
 sg13g2_o21ai_1 _09924_ (.B1(_02506_),
    .Y(_00256_),
    .A1(net382),
    .A2(_02503_));
 sg13g2_nor2_1 _09925_ (.A(net404),
    .B(_02503_),
    .Y(_02507_));
 sg13g2_a21oi_1 _09926_ (.A1(_02230_),
    .A2(_02503_),
    .Y(_00257_),
    .B1(_02507_));
 sg13g2_nor2_1 _09927_ (.A(net408),
    .B(_02503_),
    .Y(_02508_));
 sg13g2_a21oi_1 _09928_ (.A1(net388),
    .A2(_02503_),
    .Y(_00258_),
    .B1(_02508_));
 sg13g2_nor2_1 _09929_ (.A(net384),
    .B(_02488_),
    .Y(_02509_));
 sg13g2_a21oi_1 _09930_ (.A1(_02394_),
    .A2(_02488_),
    .Y(_00259_),
    .B1(_02509_));
 sg13g2_nor2_1 _09931_ (.A(net383),
    .B(_02488_),
    .Y(_02510_));
 sg13g2_a21oi_1 _09932_ (.A1(_02398_),
    .A2(_02488_),
    .Y(_00260_),
    .B1(_02510_));
 sg13g2_inv_1 _09933_ (.Y(_02511_),
    .A(\ppu.copper_inst.store_valid ));
 sg13g2_inv_1 _09934_ (.Y(_02512_),
    .A(_02207_));
 sg13g2_inv_1 _09935_ (.Y(_02513_),
    .A(_02377_));
 sg13g2_o21ai_1 _09936_ (.B1(_02232_),
    .Y(_02514_),
    .A1(_00076_),
    .A2(_02513_));
 sg13g2_nor2_1 _09937_ (.A(net264),
    .B(_01800_),
    .Y(_02515_));
 sg13g2_nand3_1 _09938_ (.B(_02268_),
    .C(_02515_),
    .A(_02514_),
    .Y(_02516_));
 sg13g2_o21ai_1 _09939_ (.B1(_02516_),
    .Y(_00261_),
    .A1(_02511_),
    .A2(_02512_));
 sg13g2_buf_1 _09940_ (.A(_02207_),
    .X(_02517_));
 sg13g2_buf_1 _09941_ (.A(_02207_),
    .X(_02518_));
 sg13g2_nor2_1 _09942_ (.A(\ppu.copper_inst.dt_sreg[3] ),
    .B(net198),
    .Y(_02519_));
 sg13g2_a21oi_1 _09943_ (.A1(_01861_),
    .A2(net199),
    .Y(_00429_),
    .B1(_02519_));
 sg13g2_inv_1 _09944_ (.Y(_02520_),
    .A(_02515_));
 sg13g2_inv_1 _09945_ (.Y(_02521_),
    .A(\ppu.copper_inst.dt_sreg[8] ));
 sg13g2_nor3_1 _09946_ (.A(\ppu.copper_inst.dt_sreg[7] ),
    .B(\ppu.copper_inst.dt_sreg[6] ),
    .C(_02521_),
    .Y(_02522_));
 sg13g2_nor3_1 _09947_ (.A(\ppu.copper_inst.dt_sreg[4] ),
    .B(\ppu.copper_inst.dt_sreg[3] ),
    .C(_00035_),
    .Y(_02523_));
 sg13g2_nor3_1 _09948_ (.A(_02231_),
    .B(_02522_),
    .C(_02523_),
    .Y(_02524_));
 sg13g2_or2_1 _09949_ (.X(_02525_),
    .B(_02524_),
    .A(\ppu.copper_inst.fast_mode ));
 sg13g2_buf_2 _09950_ (.A(\ppu.ram_running ),
    .X(_02526_));
 sg13g2_nand3_1 _09951_ (.B(\ppu.copper_inst.on ),
    .C(_02526_),
    .A(_02511_),
    .Y(_02527_));
 sg13g2_nor3_1 _09952_ (.A(\ppu.copper_inst.dt_sreg[10] ),
    .B(\ppu.copper_inst.dt_sreg[9] ),
    .C(_01898_),
    .Y(_02528_));
 sg13g2_nor2_1 _09953_ (.A(_02527_),
    .B(_02528_),
    .Y(_02529_));
 sg13g2_nand2_1 _09954_ (.Y(_02530_),
    .A(_02525_),
    .B(_02529_));
 sg13g2_buf_2 _09955_ (.A(_02530_),
    .X(_02531_));
 sg13g2_inv_1 _09956_ (.Y(_02532_),
    .A(_02531_));
 sg13g2_mux2_1 _09957_ (.A0(\ppu.scroll_regs[0][2] ),
    .A1(\ppu.scroll_regs[2][2] ),
    .S(net409),
    .X(_02533_));
 sg13g2_xnor2_1 _09958_ (.Y(_02534_),
    .A(_00034_),
    .B(_02533_));
 sg13g2_inv_1 _09959_ (.Y(_02535_),
    .A(\ppu.scroll_regs[0][1] ));
 sg13g2_nand2_1 _09960_ (.Y(_02536_),
    .A(net409),
    .B(\ppu.scroll_regs[2][1] ));
 sg13g2_o21ai_1 _09961_ (.B1(_02536_),
    .Y(_02537_),
    .A1(net409),
    .A2(_02535_));
 sg13g2_xnor2_1 _09962_ (.Y(_02538_),
    .A(_00033_),
    .B(_02537_));
 sg13g2_nand2_1 _09963_ (.Y(_02539_),
    .A(net409),
    .B(\ppu.scroll_regs[2][0] ));
 sg13g2_inv_1 _09964_ (.Y(_02540_),
    .A(_02539_));
 sg13g2_a21oi_1 _09965_ (.A1(_02209_),
    .A2(\ppu.scroll_regs[0][0] ),
    .Y(_02541_),
    .B1(_02540_));
 sg13g2_nor2_1 _09966_ (.A(_01943_),
    .B(_02541_),
    .Y(_02542_));
 sg13g2_nand2_1 _09967_ (.Y(_02543_),
    .A(_02538_),
    .B(_02542_));
 sg13g2_nand2_1 _09968_ (.Y(_02544_),
    .A(_02537_),
    .B(_01816_));
 sg13g2_nand2_1 _09969_ (.Y(_02545_),
    .A(_02543_),
    .B(_02544_));
 sg13g2_xnor2_1 _09970_ (.Y(_02546_),
    .A(_02534_),
    .B(_02545_));
 sg13g2_nand2_1 _09971_ (.Y(_02547_),
    .A(_02541_),
    .B(_01943_));
 sg13g2_xor2_1 _09972_ (.B(_02538_),
    .A(_02547_),
    .X(_02548_));
 sg13g2_nand2_1 _09973_ (.Y(_02549_),
    .A(_01803_),
    .B(_01830_));
 sg13g2_nor2_1 _09974_ (.A(_01812_),
    .B(_02549_),
    .Y(_02550_));
 sg13g2_nor2b_1 _09975_ (.A(_02550_),
    .B_N(_02278_),
    .Y(_02551_));
 sg13g2_nor2b_1 _09976_ (.A(net409),
    .B_N(\ppu.display_mask[3] ),
    .Y(_02552_));
 sg13g2_a21oi_1 _09977_ (.A1(\ppu.display_mask[4] ),
    .A2(net392),
    .Y(_02553_),
    .B1(_02552_));
 sg13g2_nor3_1 _09978_ (.A(_00180_),
    .B(_02551_),
    .C(_02553_),
    .Y(_02554_));
 sg13g2_nand3_1 _09979_ (.B(_02548_),
    .C(_02554_),
    .A(_02546_),
    .Y(_02555_));
 sg13g2_nor2_1 _09980_ (.A(_01815_),
    .B(_01849_),
    .Y(_02556_));
 sg13g2_nand2_1 _09981_ (.Y(_02557_),
    .A(_02556_),
    .B(_01805_));
 sg13g2_inv_1 _09982_ (.Y(_02558_),
    .A(_00029_));
 sg13g2_nand3_1 _09983_ (.B(_02558_),
    .C(_02306_),
    .A(_02557_),
    .Y(_02559_));
 sg13g2_buf_1 _09984_ (.A(_02559_),
    .X(_02560_));
 sg13g2_nor2_1 _09985_ (.A(_02555_),
    .B(_02560_),
    .Y(_02561_));
 sg13g2_nor2b_1 _09986_ (.A(_02560_),
    .B_N(\ppu.display_mask[5] ),
    .Y(_02562_));
 sg13g2_buf_1 _09987_ (.A(\ppu.sprite_buffer.out_counter_oam[1] ),
    .X(_02563_));
 sg13g2_xnor2_1 _09988_ (.Y(_02564_),
    .A(_01872_),
    .B(_02563_));
 sg13g2_a21oi_1 _09989_ (.A1(_01879_),
    .A2(_02564_),
    .Y(_02565_),
    .B1(\ppu.sprite_buffer.oam_load_sprite_valid ));
 sg13g2_buf_2 _09990_ (.A(\ppu.sprite_buffer.in_counters[1][1] ),
    .X(_02566_));
 sg13g2_xor2_1 _09991_ (.B(_02566_),
    .A(\ppu.sprite_buffer.out_counters[2][1] ),
    .X(_02567_));
 sg13g2_buf_1 _09992_ (.A(\ppu.sprite_buffer.in_counters[1][2] ),
    .X(_02568_));
 sg13g2_xor2_1 _09993_ (.B(_02568_),
    .A(\ppu.sprite_buffer.out_counters[2][2] ),
    .X(_02569_));
 sg13g2_xor2_1 _09994_ (.B(\ppu.sprite_buffer.in_counters[1][0] ),
    .A(\ppu.sprite_buffer.out_counters[2][0] ),
    .X(_02570_));
 sg13g2_nor3_1 _09995_ (.A(_02567_),
    .B(_02569_),
    .C(_02570_),
    .Y(_02571_));
 sg13g2_nand2b_1 _09996_ (.Y(_02572_),
    .B(_02571_),
    .A_N(_02565_));
 sg13g2_nand2_1 _09997_ (.Y(_02573_),
    .A(_02562_),
    .B(_02572_));
 sg13g2_nor3_1 _09998_ (.A(net234),
    .B(_02561_),
    .C(_02573_),
    .Y(_02574_));
 sg13g2_nor3_1 _09999_ (.A(_01859_),
    .B(_00031_),
    .C(_01861_),
    .Y(_02575_));
 sg13g2_buf_1 _10000_ (.A(_02575_),
    .X(_02576_));
 sg13g2_nand2b_1 _10001_ (.Y(_02577_),
    .B(net295),
    .A_N(_02560_));
 sg13g2_nor2b_1 _10002_ (.A(_02574_),
    .B_N(_02577_),
    .Y(_02578_));
 sg13g2_buf_2 _10003_ (.A(_02578_),
    .X(_02579_));
 sg13g2_buf_1 _10004_ (.A(_02579_),
    .X(_02580_));
 sg13g2_nand2_1 _10005_ (.Y(_02581_),
    .A(_02517_),
    .B(\ppu.copper_inst.dt_sreg[10] ));
 sg13g2_o21ai_1 _10006_ (.B1(_02581_),
    .Y(_00430_),
    .A1(_02520_),
    .A2(net121));
 sg13g2_o21ai_1 _10007_ (.B1(net249),
    .Y(_02582_),
    .A1(\ppu.copper_inst.dt_sreg[11] ),
    .A2(net236));
 sg13g2_inv_2 _10008_ (.Y(_02583_),
    .A(net295));
 sg13g2_a21oi_1 _10009_ (.A1(_02583_),
    .A2(_02555_),
    .Y(_02584_),
    .B1(_02560_));
 sg13g2_buf_2 _10010_ (.A(_02584_),
    .X(_02585_));
 sg13g2_nor2_1 _10011_ (.A(net234),
    .B(_02585_),
    .Y(_02586_));
 sg13g2_inv_1 _10012_ (.Y(_02587_),
    .A(_02586_));
 sg13g2_nor2_1 _10013_ (.A(net297),
    .B(_02587_),
    .Y(_02588_));
 sg13g2_nor2_1 _10014_ (.A(_02582_),
    .B(_02588_),
    .Y(_00431_));
 sg13g2_nor2_1 _10015_ (.A(\ppu.copper_inst.dt_sreg[4] ),
    .B(net198),
    .Y(_02589_));
 sg13g2_a21oi_1 _10016_ (.A1(_01901_),
    .A2(net199),
    .Y(_00432_),
    .B1(_02589_));
 sg13g2_inv_1 _10017_ (.Y(_02590_),
    .A(\ppu.copper_inst.dt_sreg[5] ));
 sg13g2_nand2_1 _10018_ (.Y(_02591_),
    .A(net198),
    .B(\ppu.copper_inst.dt_out[2] ));
 sg13g2_o21ai_1 _10019_ (.B1(_02591_),
    .Y(_00433_),
    .A1(_02590_),
    .A2(net199));
 sg13g2_nand2_1 _10020_ (.Y(_02592_),
    .A(net198),
    .B(\ppu.copper_inst.dt_sreg[3] ));
 sg13g2_o21ai_1 _10021_ (.B1(_02592_),
    .Y(_00434_),
    .A1(_01892_),
    .A2(net199));
 sg13g2_nor2_1 _10022_ (.A(\ppu.copper_inst.dt_sreg[7] ),
    .B(net198),
    .Y(_02593_));
 sg13g2_a21oi_1 _10023_ (.A1(_01895_),
    .A2(net199),
    .Y(_00435_),
    .B1(_02593_));
 sg13g2_nor2_1 _10024_ (.A(\ppu.copper_inst.dt_sreg[8] ),
    .B(net198),
    .Y(_02594_));
 sg13g2_a21oi_1 _10025_ (.A1(_02590_),
    .A2(net199),
    .Y(_00436_),
    .B1(_02594_));
 sg13g2_nor2_1 _10026_ (.A(\ppu.copper_inst.dt_sreg[9] ),
    .B(net198),
    .Y(_02595_));
 sg13g2_a21oi_1 _10027_ (.A1(_01892_),
    .A2(net199),
    .Y(_00437_),
    .B1(_02595_));
 sg13g2_nand2_1 _10028_ (.Y(_02596_),
    .A(net198),
    .B(\ppu.copper_inst.dt_sreg[7] ));
 sg13g2_o21ai_1 _10029_ (.B1(_02596_),
    .Y(_00438_),
    .A1(_01897_),
    .A2(_02517_));
 sg13g2_nor2_1 _10030_ (.A(\ppu.copper_inst.dt_sreg[11] ),
    .B(_02518_),
    .Y(_02597_));
 sg13g2_a21oi_1 _10031_ (.A1(_02521_),
    .A2(net199),
    .Y(_00439_),
    .B1(_02597_));
 sg13g2_nand2_1 _10032_ (.Y(_02598_),
    .A(\ppu.sprite_buffer.scan_enabled ),
    .B(_01858_));
 sg13g2_o21ai_1 _10033_ (.B1(_02571_),
    .Y(_02599_),
    .A1(_02598_),
    .A2(_02565_));
 sg13g2_nand3_1 _10034_ (.B(_02562_),
    .C(_02599_),
    .A(_02586_),
    .Y(_02600_));
 sg13g2_nand2_1 _10035_ (.Y(_02601_),
    .A(_02561_),
    .B(_02583_));
 sg13g2_nand2_1 _10036_ (.Y(_02602_),
    .A(_02600_),
    .B(_02601_));
 sg13g2_inv_1 _10037_ (.Y(_02603_),
    .A(_02602_));
 sg13g2_nand2_1 _10038_ (.Y(_02604_),
    .A(_02518_),
    .B(\ppu.copper_inst.dt_sreg[9] ));
 sg13g2_o21ai_1 _10039_ (.B1(_02604_),
    .Y(_00440_),
    .A1(_02520_),
    .A2(_02603_));
 sg13g2_nor4_1 _10040_ (.A(_02381_),
    .B(_02383_),
    .C(_02420_),
    .D(_02379_),
    .Y(_02605_));
 sg13g2_nor2_1 _10041_ (.A(_02292_),
    .B(_02293_),
    .Y(_02606_));
 sg13g2_nand2_1 _10042_ (.Y(_02607_),
    .A(_02605_),
    .B(_02606_));
 sg13g2_buf_1 _10043_ (.A(_02607_),
    .X(_02608_));
 sg13g2_buf_1 _10044_ (.A(net106),
    .X(_02609_));
 sg13g2_nand2_1 _10045_ (.Y(_02610_),
    .A(_02609_),
    .B(\ppu.scroll_regs[0][0] ));
 sg13g2_o21ai_1 _10046_ (.B1(_02610_),
    .Y(_00468_),
    .A1(net388),
    .A2(net98));
 sg13g2_nor2_1 _10047_ (.A(_02392_),
    .B(net106),
    .Y(_02611_));
 sg13g2_a21oi_1 _10048_ (.A1(_02535_),
    .A2(_02609_),
    .Y(_00469_),
    .B1(_02611_));
 sg13g2_nand2_1 _10049_ (.Y(_02612_),
    .A(_02608_),
    .B(\ppu.scroll_regs[0][2] ));
 sg13g2_o21ai_1 _10050_ (.B1(_02612_),
    .Y(_00470_),
    .A1(net339),
    .A2(net98));
 sg13g2_inv_1 _10051_ (.Y(_02613_),
    .A(\ppu.scroll_regs[0][3] ));
 sg13g2_nor2_1 _10052_ (.A(_02400_),
    .B(net106),
    .Y(_02614_));
 sg13g2_a21oi_1 _10053_ (.A1(_02613_),
    .A2(net98),
    .Y(_00471_),
    .B1(_02614_));
 sg13g2_inv_1 _10054_ (.Y(_02615_),
    .A(\ppu.scroll_regs[0][4] ));
 sg13g2_nor2_1 _10055_ (.A(_02404_),
    .B(net106),
    .Y(_02616_));
 sg13g2_a21oi_1 _10056_ (.A1(_02615_),
    .A2(net98),
    .Y(_00472_),
    .B1(_02616_));
 sg13g2_inv_1 _10057_ (.Y(_02617_),
    .A(\ppu.scroll_regs[0][5] ));
 sg13g2_nor2_1 _10058_ (.A(_02408_),
    .B(net106),
    .Y(_02618_));
 sg13g2_a21oi_1 _10059_ (.A1(_02617_),
    .A2(net98),
    .Y(_00473_),
    .B1(_02618_));
 sg13g2_inv_1 _10060_ (.Y(_02619_),
    .A(\ppu.scroll_regs[0][6] ));
 sg13g2_nor2_1 _10061_ (.A(net406),
    .B(net106),
    .Y(_02620_));
 sg13g2_a21oi_1 _10062_ (.A1(_02619_),
    .A2(net98),
    .Y(_00474_),
    .B1(_02620_));
 sg13g2_inv_1 _10063_ (.Y(_02621_),
    .A(\ppu.scroll_regs[0][7] ));
 sg13g2_nor2_1 _10064_ (.A(_02414_),
    .B(net106),
    .Y(_02622_));
 sg13g2_a21oi_1 _10065_ (.A1(_02621_),
    .A2(net98),
    .Y(_00475_),
    .B1(_02622_));
 sg13g2_inv_1 _10066_ (.Y(_02623_),
    .A(\ppu.scroll_regs[0][8] ));
 sg13g2_nor2_1 _10067_ (.A(_02417_),
    .B(net106),
    .Y(_02624_));
 sg13g2_a21oi_1 _10068_ (.A1(_02623_),
    .A2(net98),
    .Y(_00476_),
    .B1(_02624_));
 sg13g2_nor4_1 _10069_ (.A(_02381_),
    .B(_02384_),
    .C(_02420_),
    .D(_02379_),
    .Y(_02625_));
 sg13g2_nand2_1 _10070_ (.Y(_02626_),
    .A(_02625_),
    .B(_02606_));
 sg13g2_buf_1 _10071_ (.A(_02626_),
    .X(_02627_));
 sg13g2_buf_1 _10072_ (.A(net105),
    .X(_02628_));
 sg13g2_nand2_1 _10073_ (.Y(_02629_),
    .A(net97),
    .B(\ppu.scroll_regs[1][0] ));
 sg13g2_o21ai_1 _10074_ (.B1(_02629_),
    .Y(_00477_),
    .A1(net388),
    .A2(net97));
 sg13g2_inv_1 _10075_ (.Y(_02630_),
    .A(\ppu.scroll_regs[1][1] ));
 sg13g2_nor2_1 _10076_ (.A(_02392_),
    .B(net105),
    .Y(_02631_));
 sg13g2_a21oi_1 _10077_ (.A1(_02630_),
    .A2(_02628_),
    .Y(_00478_),
    .B1(_02631_));
 sg13g2_inv_1 _10078_ (.Y(_02632_),
    .A(\ppu.scroll_regs[1][2] ));
 sg13g2_nor2_1 _10079_ (.A(_02396_),
    .B(_02627_),
    .Y(_02633_));
 sg13g2_a21oi_1 _10080_ (.A1(_02632_),
    .A2(_02628_),
    .Y(_00479_),
    .B1(_02633_));
 sg13g2_inv_1 _10081_ (.Y(_02634_),
    .A(\ppu.scroll_regs[1][3] ));
 sg13g2_nor2_1 _10082_ (.A(_02400_),
    .B(net105),
    .Y(_02635_));
 sg13g2_a21oi_1 _10083_ (.A1(_02634_),
    .A2(net97),
    .Y(_00480_),
    .B1(_02635_));
 sg13g2_inv_1 _10084_ (.Y(_02636_),
    .A(\ppu.scroll_regs[1][4] ));
 sg13g2_nor2_1 _10085_ (.A(_02404_),
    .B(net105),
    .Y(_02637_));
 sg13g2_a21oi_1 _10086_ (.A1(_02636_),
    .A2(net97),
    .Y(_00481_),
    .B1(_02637_));
 sg13g2_inv_1 _10087_ (.Y(_02638_),
    .A(\ppu.scroll_regs[1][5] ));
 sg13g2_nor2_1 _10088_ (.A(_02408_),
    .B(net105),
    .Y(_02639_));
 sg13g2_a21oi_1 _10089_ (.A1(_02638_),
    .A2(net97),
    .Y(_00482_),
    .B1(_02639_));
 sg13g2_inv_1 _10090_ (.Y(_02640_),
    .A(\ppu.scroll_regs[1][6] ));
 sg13g2_nor2_1 _10091_ (.A(net406),
    .B(net105),
    .Y(_02641_));
 sg13g2_a21oi_1 _10092_ (.A1(_02640_),
    .A2(net97),
    .Y(_00483_),
    .B1(_02641_));
 sg13g2_inv_1 _10093_ (.Y(_02642_),
    .A(\ppu.scroll_regs[1][7] ));
 sg13g2_nor2_1 _10094_ (.A(_02414_),
    .B(net105),
    .Y(_02643_));
 sg13g2_a21oi_1 _10095_ (.A1(_02642_),
    .A2(net97),
    .Y(_00484_),
    .B1(_02643_));
 sg13g2_nand2_1 _10096_ (.Y(_02644_),
    .A(net105),
    .B(\ppu.scroll_regs[1][8] ));
 sg13g2_o21ai_1 _10097_ (.B1(_02644_),
    .Y(_00485_),
    .A1(net385),
    .A2(net97));
 sg13g2_nand4_1 _10098_ (.B(_02387_),
    .C(_02434_),
    .A(_02378_),
    .Y(_02645_),
    .D(_02606_));
 sg13g2_buf_1 _10099_ (.A(_02645_),
    .X(_02646_));
 sg13g2_buf_1 _10100_ (.A(net120),
    .X(_02647_));
 sg13g2_nand2_1 _10101_ (.Y(_02648_),
    .A(net117),
    .B(\ppu.scroll_regs[2][0] ));
 sg13g2_o21ai_1 _10102_ (.B1(_02648_),
    .Y(_00486_),
    .A1(net388),
    .A2(net117));
 sg13g2_nand2_1 _10103_ (.Y(_02649_),
    .A(net120),
    .B(\ppu.scroll_regs[2][1] ));
 sg13g2_o21ai_1 _10104_ (.B1(_02649_),
    .Y(_00487_),
    .A1(net340),
    .A2(_02647_));
 sg13g2_nand2_1 _10105_ (.Y(_02650_),
    .A(_02646_),
    .B(\ppu.scroll_regs[2][2] ));
 sg13g2_o21ai_1 _10106_ (.B1(_02650_),
    .Y(_00488_),
    .A1(net339),
    .A2(_02647_));
 sg13g2_nand2_1 _10107_ (.Y(_02651_),
    .A(net120),
    .B(\ppu.scroll_regs[2][3] ));
 sg13g2_o21ai_1 _10108_ (.B1(_02651_),
    .Y(_00489_),
    .A1(net338),
    .A2(net117));
 sg13g2_nand2_1 _10109_ (.Y(_02652_),
    .A(net120),
    .B(\ppu.scroll_regs[2][4] ));
 sg13g2_o21ai_1 _10110_ (.B1(_02652_),
    .Y(_00490_),
    .A1(net337),
    .A2(net117));
 sg13g2_nand2_1 _10111_ (.Y(_02653_),
    .A(net120),
    .B(\ppu.scroll_regs[2][5] ));
 sg13g2_o21ai_1 _10112_ (.B1(_02653_),
    .Y(_00491_),
    .A1(net387),
    .A2(net117));
 sg13g2_nand2_1 _10113_ (.Y(_02654_),
    .A(net120),
    .B(\ppu.scroll_regs[2][6] ));
 sg13g2_o21ai_1 _10114_ (.B1(_02654_),
    .Y(_00492_),
    .A1(_02412_),
    .A2(net117));
 sg13g2_nand2_1 _10115_ (.Y(_02655_),
    .A(net120),
    .B(\ppu.scroll_regs[2][7] ));
 sg13g2_o21ai_1 _10116_ (.B1(_02655_),
    .Y(_00493_),
    .A1(net386),
    .A2(net117));
 sg13g2_nand2_1 _10117_ (.Y(_02656_),
    .A(net120),
    .B(\ppu.scroll_regs[2][8] ));
 sg13g2_o21ai_1 _10118_ (.B1(_02656_),
    .Y(_00494_),
    .A1(net385),
    .A2(net117));
 sg13g2_nand4_1 _10119_ (.B(_02387_),
    .C(_02452_),
    .A(_02378_),
    .Y(_02657_),
    .D(_02606_));
 sg13g2_buf_1 _10120_ (.A(_02657_),
    .X(_02658_));
 sg13g2_buf_1 _10121_ (.A(net119),
    .X(_02659_));
 sg13g2_nand2_1 _10122_ (.Y(_02660_),
    .A(net116),
    .B(\ppu.scroll_regs[3][0] ));
 sg13g2_o21ai_1 _10123_ (.B1(_02660_),
    .Y(_00495_),
    .A1(net388),
    .A2(net116));
 sg13g2_nand2_1 _10124_ (.Y(_02661_),
    .A(net119),
    .B(\ppu.scroll_regs[3][1] ));
 sg13g2_o21ai_1 _10125_ (.B1(_02661_),
    .Y(_00496_),
    .A1(net340),
    .A2(_02659_));
 sg13g2_nand2_1 _10126_ (.Y(_02662_),
    .A(net119),
    .B(\ppu.scroll_regs[3][2] ));
 sg13g2_o21ai_1 _10127_ (.B1(_02662_),
    .Y(_00497_),
    .A1(net339),
    .A2(net116));
 sg13g2_nand2_1 _10128_ (.Y(_02663_),
    .A(_02658_),
    .B(\ppu.scroll_regs[3][3] ));
 sg13g2_o21ai_1 _10129_ (.B1(_02663_),
    .Y(_00498_),
    .A1(net338),
    .A2(_02659_));
 sg13g2_nand2_1 _10130_ (.Y(_02664_),
    .A(net119),
    .B(\ppu.scroll_regs[3][4] ));
 sg13g2_o21ai_1 _10131_ (.B1(_02664_),
    .Y(_00499_),
    .A1(net337),
    .A2(net116));
 sg13g2_nand2_1 _10132_ (.Y(_02665_),
    .A(net119),
    .B(\ppu.scroll_regs[3][5] ));
 sg13g2_o21ai_1 _10133_ (.B1(_02665_),
    .Y(_00500_),
    .A1(net387),
    .A2(net116));
 sg13g2_nand2_1 _10134_ (.Y(_02666_),
    .A(net119),
    .B(\ppu.scroll_regs[3][6] ));
 sg13g2_o21ai_1 _10135_ (.B1(_02666_),
    .Y(_00501_),
    .A1(_02412_),
    .A2(net116));
 sg13g2_nand2_1 _10136_ (.Y(_02667_),
    .A(net119),
    .B(\ppu.scroll_regs[3][7] ));
 sg13g2_o21ai_1 _10137_ (.B1(_02667_),
    .Y(_00502_),
    .A1(net386),
    .A2(net116));
 sg13g2_nand2_1 _10138_ (.Y(_02668_),
    .A(net119),
    .B(\ppu.scroll_regs[3][8] ));
 sg13g2_o21ai_1 _10139_ (.B1(_02668_),
    .Y(_00503_),
    .A1(net385),
    .A2(net116));
 sg13g2_nor3_1 _10140_ (.A(_01860_),
    .B(\ppu.copper_inst.dt_out[2] ),
    .C(_01901_),
    .Y(_02669_));
 sg13g2_buf_1 _10141_ (.A(_02669_),
    .X(_02670_));
 sg13g2_inv_1 _10142_ (.Y(_02671_),
    .A(_02566_));
 sg13g2_inv_1 _10143_ (.Y(_02672_),
    .A(\ppu.sprite_buffer.in_counters[1][0] ));
 sg13g2_nor2_1 _10144_ (.A(_02568_),
    .B(_02672_),
    .Y(_02673_));
 sg13g2_nand3_1 _10145_ (.B(_02671_),
    .C(_02673_),
    .A(_02670_),
    .Y(_02674_));
 sg13g2_buf_2 _10146_ (.A(_02674_),
    .X(_02675_));
 sg13g2_buf_1 _10147_ (.A(_02675_),
    .X(_02676_));
 sg13g2_mux2_1 _10148_ (.A0(\ppu.sprite_buffer.attr_x[0][4] ),
    .A1(\ppu.sprite_buffer.attr_x[0][0] ),
    .S(net233),
    .X(_00506_));
 sg13g2_inv_1 _10149_ (.Y(_02677_),
    .A(\ppu.sprite_buffer.attr_x[0][10] ));
 sg13g2_buf_1 _10150_ (.A(_02675_),
    .X(_02678_));
 sg13g2_nor2_1 _10151_ (.A(\ppu.sprite_buffer.attr_x[0][14] ),
    .B(_02675_),
    .Y(_02679_));
 sg13g2_a21oi_1 _10152_ (.A1(_02677_),
    .A2(net232),
    .Y(_00507_),
    .B1(_02679_));
 sg13g2_inv_1 _10153_ (.Y(_02680_),
    .A(\ppu.sprite_buffer.attr_x[0][11] ));
 sg13g2_nor2_1 _10154_ (.A(\ppu.sprite_buffer.attr_x[0][15] ),
    .B(_02675_),
    .Y(_02681_));
 sg13g2_a21oi_1 _10155_ (.A1(_02680_),
    .A2(_02678_),
    .Y(_00508_),
    .B1(_02681_));
 sg13g2_nor2_1 _10156_ (.A(net384),
    .B(_02675_),
    .Y(_02682_));
 sg13g2_a21oi_1 _10157_ (.A1(_02044_),
    .A2(net232),
    .Y(_00509_),
    .B1(_02682_));
 sg13g2_inv_1 _10158_ (.Y(_02683_),
    .A(\ppu.sprite_buffer.attr_x[0][13] ));
 sg13g2_nor2_1 _10159_ (.A(net383),
    .B(_02675_),
    .Y(_02684_));
 sg13g2_a21oi_1 _10160_ (.A1(_02683_),
    .A2(net232),
    .Y(_00510_),
    .B1(_02684_));
 sg13g2_inv_1 _10161_ (.Y(_02685_),
    .A(net404));
 sg13g2_buf_1 _10162_ (.A(_02685_),
    .X(_02686_));
 sg13g2_nand2_1 _10163_ (.Y(_02687_),
    .A(net233),
    .B(\ppu.sprite_buffer.attr_x[0][14] ));
 sg13g2_o21ai_1 _10164_ (.B1(_02687_),
    .Y(_00511_),
    .A1(net336),
    .A2(net232));
 sg13g2_buf_1 _10165_ (.A(_01867_),
    .X(_02688_));
 sg13g2_nand2_1 _10166_ (.Y(_02689_),
    .A(net233),
    .B(\ppu.sprite_buffer.attr_x[0][15] ));
 sg13g2_o21ai_1 _10167_ (.B1(_02689_),
    .Y(_00512_),
    .A1(net335),
    .A2(_02678_));
 sg13g2_mux2_1 _10168_ (.A0(\ppu.sprite_buffer.attr_x[0][5] ),
    .A1(\ppu.sprite_buffer.attr_x[0][1] ),
    .S(_02676_),
    .X(_00513_));
 sg13g2_mux2_1 _10169_ (.A0(\ppu.sprite_buffer.attr_x[0][6] ),
    .A1(\ppu.sprite_buffer.attr_x[0][2] ),
    .S(net233),
    .X(_00514_));
 sg13g2_mux2_1 _10170_ (.A0(\ppu.sprite_buffer.attr_x[0][7] ),
    .A1(\ppu.sprite_buffer.attr_x[0][3] ),
    .S(net233),
    .X(_00515_));
 sg13g2_mux2_1 _10171_ (.A0(\ppu.sprite_buffer.attr_x[0][8] ),
    .A1(\ppu.sprite_buffer.attr_x[0][4] ),
    .S(net233),
    .X(_00516_));
 sg13g2_mux2_1 _10172_ (.A0(\ppu.sprite_buffer.attr_x[0][9] ),
    .A1(\ppu.sprite_buffer.attr_x[0][5] ),
    .S(_02676_),
    .X(_00517_));
 sg13g2_nand2_1 _10173_ (.Y(_02690_),
    .A(net233),
    .B(\ppu.sprite_buffer.attr_x[0][6] ));
 sg13g2_o21ai_1 _10174_ (.B1(_02690_),
    .Y(_00518_),
    .A1(_02677_),
    .A2(net232));
 sg13g2_nand2_1 _10175_ (.Y(_02691_),
    .A(net233),
    .B(\ppu.sprite_buffer.attr_x[0][7] ));
 sg13g2_o21ai_1 _10176_ (.B1(_02691_),
    .Y(_00519_),
    .A1(_02680_),
    .A2(net232));
 sg13g2_nand2_1 _10177_ (.Y(_02692_),
    .A(_02675_),
    .B(\ppu.sprite_buffer.attr_x[0][8] ));
 sg13g2_o21ai_1 _10178_ (.B1(_02692_),
    .Y(_00520_),
    .A1(_02044_),
    .A2(net232));
 sg13g2_nand2_1 _10179_ (.Y(_02693_),
    .A(_02675_),
    .B(\ppu.sprite_buffer.attr_x[0][9] ));
 sg13g2_o21ai_1 _10180_ (.B1(_02693_),
    .Y(_00521_),
    .A1(_02683_),
    .A2(net232));
 sg13g2_nand3_1 _10181_ (.B(_02566_),
    .C(_02673_),
    .A(_02670_),
    .Y(_02694_));
 sg13g2_buf_2 _10182_ (.A(_02694_),
    .X(_02695_));
 sg13g2_buf_1 _10183_ (.A(_02695_),
    .X(_02696_));
 sg13g2_mux2_1 _10184_ (.A0(\ppu.sprite_buffer.attr_x[1][4] ),
    .A1(\ppu.sprite_buffer.attr_x[1][0] ),
    .S(net231),
    .X(_00522_));
 sg13g2_inv_1 _10185_ (.Y(_02697_),
    .A(\ppu.sprite_buffer.attr_x[1][10] ));
 sg13g2_buf_1 _10186_ (.A(_02695_),
    .X(_02698_));
 sg13g2_nor2_1 _10187_ (.A(\ppu.sprite_buffer.attr_x[1][14] ),
    .B(_02695_),
    .Y(_02699_));
 sg13g2_a21oi_1 _10188_ (.A1(_02697_),
    .A2(net230),
    .Y(_00523_),
    .B1(_02699_));
 sg13g2_inv_1 _10189_ (.Y(_02700_),
    .A(\ppu.sprite_buffer.attr_x[1][11] ));
 sg13g2_nor2_1 _10190_ (.A(\ppu.sprite_buffer.attr_x[1][15] ),
    .B(_02695_),
    .Y(_02701_));
 sg13g2_a21oi_1 _10191_ (.A1(_02700_),
    .A2(net230),
    .Y(_00524_),
    .B1(_02701_));
 sg13g2_nor2_1 _10192_ (.A(net384),
    .B(_02695_),
    .Y(_02702_));
 sg13g2_a21oi_1 _10193_ (.A1(_02041_),
    .A2(net230),
    .Y(_00525_),
    .B1(_02702_));
 sg13g2_inv_1 _10194_ (.Y(_02703_),
    .A(\ppu.sprite_buffer.attr_x[1][13] ));
 sg13g2_nor2_1 _10195_ (.A(net383),
    .B(_02695_),
    .Y(_02704_));
 sg13g2_a21oi_1 _10196_ (.A1(_02703_),
    .A2(net230),
    .Y(_00526_),
    .B1(_02704_));
 sg13g2_nand2_1 _10197_ (.Y(_02705_),
    .A(net231),
    .B(\ppu.sprite_buffer.attr_x[1][14] ));
 sg13g2_o21ai_1 _10198_ (.B1(_02705_),
    .Y(_00527_),
    .A1(net336),
    .A2(net230));
 sg13g2_nand2_1 _10199_ (.Y(_02706_),
    .A(_02696_),
    .B(\ppu.sprite_buffer.attr_x[1][15] ));
 sg13g2_o21ai_1 _10200_ (.B1(_02706_),
    .Y(_00528_),
    .A1(net335),
    .A2(net230));
 sg13g2_mux2_1 _10201_ (.A0(\ppu.sprite_buffer.attr_x[1][5] ),
    .A1(\ppu.sprite_buffer.attr_x[1][1] ),
    .S(net231),
    .X(_00529_));
 sg13g2_mux2_1 _10202_ (.A0(\ppu.sprite_buffer.attr_x[1][6] ),
    .A1(\ppu.sprite_buffer.attr_x[1][2] ),
    .S(net231),
    .X(_00530_));
 sg13g2_mux2_1 _10203_ (.A0(\ppu.sprite_buffer.attr_x[1][7] ),
    .A1(\ppu.sprite_buffer.attr_x[1][3] ),
    .S(net231),
    .X(_00531_));
 sg13g2_mux2_1 _10204_ (.A0(\ppu.sprite_buffer.attr_x[1][8] ),
    .A1(\ppu.sprite_buffer.attr_x[1][4] ),
    .S(net231),
    .X(_00532_));
 sg13g2_mux2_1 _10205_ (.A0(\ppu.sprite_buffer.attr_x[1][9] ),
    .A1(\ppu.sprite_buffer.attr_x[1][5] ),
    .S(net231),
    .X(_00533_));
 sg13g2_nand2_1 _10206_ (.Y(_02707_),
    .A(_02696_),
    .B(\ppu.sprite_buffer.attr_x[1][6] ));
 sg13g2_o21ai_1 _10207_ (.B1(_02707_),
    .Y(_00534_),
    .A1(_02697_),
    .A2(net230));
 sg13g2_nand2_1 _10208_ (.Y(_02708_),
    .A(net231),
    .B(\ppu.sprite_buffer.attr_x[1][7] ));
 sg13g2_o21ai_1 _10209_ (.B1(_02708_),
    .Y(_00535_),
    .A1(_02700_),
    .A2(net230));
 sg13g2_nand2_1 _10210_ (.Y(_02709_),
    .A(_02695_),
    .B(\ppu.sprite_buffer.attr_x[1][8] ));
 sg13g2_o21ai_1 _10211_ (.B1(_02709_),
    .Y(_00536_),
    .A1(_02041_),
    .A2(_02698_));
 sg13g2_nand2_1 _10212_ (.Y(_02710_),
    .A(_02695_),
    .B(\ppu.sprite_buffer.attr_x[1][9] ));
 sg13g2_o21ai_1 _10213_ (.B1(_02710_),
    .Y(_00537_),
    .A1(_02703_),
    .A2(_02698_));
 sg13g2_nand2_1 _10214_ (.Y(_02711_),
    .A(\ppu.sprite_buffer.in_counters[1][0] ),
    .B(_02568_));
 sg13g2_inv_1 _10215_ (.Y(_02712_),
    .A(_02711_));
 sg13g2_nand3_1 _10216_ (.B(_02671_),
    .C(_02712_),
    .A(_02670_),
    .Y(_02713_));
 sg13g2_buf_1 _10217_ (.A(_02713_),
    .X(_02714_));
 sg13g2_buf_1 _10218_ (.A(net248),
    .X(_02715_));
 sg13g2_mux2_1 _10219_ (.A0(\ppu.sprite_buffer.attr_x[2][4] ),
    .A1(\ppu.sprite_buffer.attr_x[2][0] ),
    .S(_02715_),
    .X(_00538_));
 sg13g2_inv_1 _10220_ (.Y(_02716_),
    .A(\ppu.sprite_buffer.attr_x[2][10] ));
 sg13g2_buf_1 _10221_ (.A(net248),
    .X(_02717_));
 sg13g2_nor2_1 _10222_ (.A(\ppu.sprite_buffer.attr_x[2][14] ),
    .B(net248),
    .Y(_02718_));
 sg13g2_a21oi_1 _10223_ (.A1(_02716_),
    .A2(net228),
    .Y(_00539_),
    .B1(_02718_));
 sg13g2_inv_1 _10224_ (.Y(_02719_),
    .A(\ppu.sprite_buffer.attr_x[2][11] ));
 sg13g2_nor2_1 _10225_ (.A(\ppu.sprite_buffer.attr_x[2][15] ),
    .B(_02714_),
    .Y(_02720_));
 sg13g2_a21oi_1 _10226_ (.A1(_02719_),
    .A2(net228),
    .Y(_00540_),
    .B1(_02720_));
 sg13g2_inv_1 _10227_ (.Y(_02721_),
    .A(net405));
 sg13g2_nand2_1 _10228_ (.Y(_02722_),
    .A(_02715_),
    .B(\ppu.sprite_buffer.attr_x[2][12] ));
 sg13g2_o21ai_1 _10229_ (.B1(_02722_),
    .Y(_00541_),
    .A1(net381),
    .A2(_02717_));
 sg13g2_nand2_1 _10230_ (.Y(_02723_),
    .A(net229),
    .B(\ppu.sprite_buffer.attr_x[2][13] ));
 sg13g2_o21ai_1 _10231_ (.B1(_02723_),
    .Y(_00542_),
    .A1(net382),
    .A2(net228));
 sg13g2_nand2_1 _10232_ (.Y(_02724_),
    .A(net229),
    .B(\ppu.sprite_buffer.attr_x[2][14] ));
 sg13g2_o21ai_1 _10233_ (.B1(_02724_),
    .Y(_00543_),
    .A1(net336),
    .A2(net228));
 sg13g2_nand2_1 _10234_ (.Y(_02725_),
    .A(net229),
    .B(\ppu.sprite_buffer.attr_x[2][15] ));
 sg13g2_o21ai_1 _10235_ (.B1(_02725_),
    .Y(_00544_),
    .A1(net335),
    .A2(net228));
 sg13g2_mux2_1 _10236_ (.A0(\ppu.sprite_buffer.attr_x[2][5] ),
    .A1(\ppu.sprite_buffer.attr_x[2][1] ),
    .S(net229),
    .X(_00545_));
 sg13g2_mux2_1 _10237_ (.A0(\ppu.sprite_buffer.attr_x[2][6] ),
    .A1(\ppu.sprite_buffer.attr_x[2][2] ),
    .S(net229),
    .X(_00546_));
 sg13g2_mux2_1 _10238_ (.A0(\ppu.sprite_buffer.attr_x[2][7] ),
    .A1(\ppu.sprite_buffer.attr_x[2][3] ),
    .S(net229),
    .X(_00547_));
 sg13g2_nand2_1 _10239_ (.Y(_02726_),
    .A(net248),
    .B(\ppu.sprite_buffer.attr_x[2][4] ));
 sg13g2_o21ai_1 _10240_ (.B1(_02726_),
    .Y(_00548_),
    .A1(_02064_),
    .A2(net228));
 sg13g2_inv_1 _10241_ (.Y(_02727_),
    .A(\ppu.sprite_buffer.attr_x[2][9] ));
 sg13g2_nand2_1 _10242_ (.Y(_02728_),
    .A(net248),
    .B(\ppu.sprite_buffer.attr_x[2][5] ));
 sg13g2_o21ai_1 _10243_ (.B1(_02728_),
    .Y(_00549_),
    .A1(_02727_),
    .A2(net228));
 sg13g2_nand2_1 _10244_ (.Y(_02729_),
    .A(net248),
    .B(\ppu.sprite_buffer.attr_x[2][6] ));
 sg13g2_o21ai_1 _10245_ (.B1(_02729_),
    .Y(_00550_),
    .A1(_02716_),
    .A2(net229));
 sg13g2_nand2_1 _10246_ (.Y(_02730_),
    .A(_02714_),
    .B(\ppu.sprite_buffer.attr_x[2][7] ));
 sg13g2_o21ai_1 _10247_ (.B1(_02730_),
    .Y(_00551_),
    .A1(_02719_),
    .A2(net229));
 sg13g2_nor2_1 _10248_ (.A(\ppu.sprite_buffer.attr_x[2][12] ),
    .B(net248),
    .Y(_02731_));
 sg13g2_a21oi_1 _10249_ (.A1(_02064_),
    .A2(_02717_),
    .Y(_00552_),
    .B1(_02731_));
 sg13g2_nor2_1 _10250_ (.A(\ppu.sprite_buffer.attr_x[2][13] ),
    .B(net248),
    .Y(_02732_));
 sg13g2_a21oi_1 _10251_ (.A1(_02727_),
    .A2(net228),
    .Y(_00553_),
    .B1(_02732_));
 sg13g2_nand3_1 _10252_ (.B(_02566_),
    .C(_02712_),
    .A(_02670_),
    .Y(_02733_));
 sg13g2_buf_2 _10253_ (.A(_02733_),
    .X(_02734_));
 sg13g2_buf_1 _10254_ (.A(_02734_),
    .X(_02735_));
 sg13g2_mux2_1 _10255_ (.A0(\ppu.sprite_buffer.attr_x[3][4] ),
    .A1(\ppu.sprite_buffer.attr_x[3][0] ),
    .S(net227),
    .X(_00554_));
 sg13g2_inv_1 _10256_ (.Y(_02736_),
    .A(\ppu.sprite_buffer.attr_x[3][10] ));
 sg13g2_buf_1 _10257_ (.A(_02734_),
    .X(_02737_));
 sg13g2_nor2_1 _10258_ (.A(\ppu.sprite_buffer.attr_x[3][14] ),
    .B(_02734_),
    .Y(_02738_));
 sg13g2_a21oi_1 _10259_ (.A1(_02736_),
    .A2(net226),
    .Y(_00555_),
    .B1(_02738_));
 sg13g2_inv_1 _10260_ (.Y(_02739_),
    .A(\ppu.sprite_buffer.attr_x[3][11] ));
 sg13g2_nor2_1 _10261_ (.A(\ppu.sprite_buffer.attr_x[3][15] ),
    .B(_02734_),
    .Y(_02740_));
 sg13g2_a21oi_1 _10262_ (.A1(_02739_),
    .A2(net226),
    .Y(_00556_),
    .B1(_02740_));
 sg13g2_nor2_1 _10263_ (.A(net384),
    .B(_02734_),
    .Y(_02741_));
 sg13g2_a21oi_1 _10264_ (.A1(_02046_),
    .A2(net226),
    .Y(_00557_),
    .B1(_02741_));
 sg13g2_nor2_1 _10265_ (.A(net383),
    .B(_02734_),
    .Y(_02742_));
 sg13g2_a21oi_1 _10266_ (.A1(_02029_),
    .A2(net226),
    .Y(_00558_),
    .B1(_02742_));
 sg13g2_nor2_1 _10267_ (.A(net404),
    .B(_02734_),
    .Y(_02743_));
 sg13g2_a21oi_1 _10268_ (.A1(_02035_),
    .A2(net226),
    .Y(_00559_),
    .B1(_02743_));
 sg13g2_nand2_1 _10269_ (.Y(_02744_),
    .A(net227),
    .B(\ppu.sprite_buffer.attr_x[3][15] ));
 sg13g2_o21ai_1 _10270_ (.B1(_02744_),
    .Y(_00560_),
    .A1(net335),
    .A2(_02737_));
 sg13g2_mux2_1 _10271_ (.A0(\ppu.sprite_buffer.attr_x[3][5] ),
    .A1(\ppu.sprite_buffer.attr_x[3][1] ),
    .S(net227),
    .X(_00561_));
 sg13g2_mux2_1 _10272_ (.A0(\ppu.sprite_buffer.attr_x[3][6] ),
    .A1(\ppu.sprite_buffer.attr_x[3][2] ),
    .S(net227),
    .X(_00562_));
 sg13g2_mux2_1 _10273_ (.A0(\ppu.sprite_buffer.attr_x[3][7] ),
    .A1(\ppu.sprite_buffer.attr_x[3][3] ),
    .S(net227),
    .X(_00563_));
 sg13g2_mux2_1 _10274_ (.A0(\ppu.sprite_buffer.attr_x[3][8] ),
    .A1(\ppu.sprite_buffer.attr_x[3][4] ),
    .S(net227),
    .X(_00564_));
 sg13g2_mux2_1 _10275_ (.A0(\ppu.sprite_buffer.attr_x[3][9] ),
    .A1(\ppu.sprite_buffer.attr_x[3][5] ),
    .S(net227),
    .X(_00565_));
 sg13g2_nand2_1 _10276_ (.Y(_02745_),
    .A(net227),
    .B(\ppu.sprite_buffer.attr_x[3][6] ));
 sg13g2_o21ai_1 _10277_ (.B1(_02745_),
    .Y(_00566_),
    .A1(_02736_),
    .A2(net226));
 sg13g2_nand2_1 _10278_ (.Y(_02746_),
    .A(_02735_),
    .B(\ppu.sprite_buffer.attr_x[3][7] ));
 sg13g2_o21ai_1 _10279_ (.B1(_02746_),
    .Y(_00567_),
    .A1(_02739_),
    .A2(_02737_));
 sg13g2_nand2_1 _10280_ (.Y(_02747_),
    .A(_02735_),
    .B(\ppu.sprite_buffer.attr_x[3][8] ));
 sg13g2_o21ai_1 _10281_ (.B1(_02747_),
    .Y(_00568_),
    .A1(_02046_),
    .A2(net226));
 sg13g2_nand2_1 _10282_ (.Y(_02748_),
    .A(_02734_),
    .B(\ppu.sprite_buffer.attr_x[3][9] ));
 sg13g2_o21ai_1 _10283_ (.B1(_02748_),
    .Y(_00569_),
    .A1(_02029_),
    .A2(net226));
 sg13g2_inv_1 _10284_ (.Y(_02749_),
    .A(\ppu.sprite_buffer.attr_y[0][0] ));
 sg13g2_nand3_1 _10285_ (.B(_02671_),
    .C(_00061_),
    .A(_02670_),
    .Y(_02750_));
 sg13g2_buf_1 _10286_ (.A(_02750_),
    .X(_02751_));
 sg13g2_buf_1 _10287_ (.A(_02751_),
    .X(_02752_));
 sg13g2_buf_1 _10288_ (.A(_02751_),
    .X(_02753_));
 sg13g2_nor2_1 _10289_ (.A(\ppu.sprite_buffer.attr_y[0][4] ),
    .B(net224),
    .Y(_02754_));
 sg13g2_a21oi_1 _10290_ (.A1(_02749_),
    .A2(net225),
    .Y(_00570_),
    .B1(_02754_));
 sg13g2_inv_1 _10291_ (.Y(_02755_),
    .A(\ppu.sprite_buffer.attr_y[0][10] ));
 sg13g2_nor2_1 _10292_ (.A(\ppu.sprite_buffer.attr_y[0][14] ),
    .B(net224),
    .Y(_02756_));
 sg13g2_a21oi_1 _10293_ (.A1(_02755_),
    .A2(net225),
    .Y(_00571_),
    .B1(_02756_));
 sg13g2_inv_1 _10294_ (.Y(_02757_),
    .A(\ppu.sprite_buffer.attr_y[0][11] ));
 sg13g2_nor2_1 _10295_ (.A(\ppu.sprite_buffer.attr_y[0][15] ),
    .B(net224),
    .Y(_02758_));
 sg13g2_a21oi_1 _10296_ (.A1(_02757_),
    .A2(net225),
    .Y(_00572_),
    .B1(_02758_));
 sg13g2_inv_1 _10297_ (.Y(_02759_),
    .A(\ppu.sprite_buffer.attr_y[0][12] ));
 sg13g2_buf_1 _10298_ (.A(_02751_),
    .X(_02760_));
 sg13g2_nor2_1 _10299_ (.A(net384),
    .B(net223),
    .Y(_02761_));
 sg13g2_a21oi_1 _10300_ (.A1(_02759_),
    .A2(net225),
    .Y(_00573_),
    .B1(_02761_));
 sg13g2_inv_1 _10301_ (.Y(_02762_),
    .A(\ppu.sprite_buffer.attr_y[0][13] ));
 sg13g2_nor2_1 _10302_ (.A(net383),
    .B(net223),
    .Y(_02763_));
 sg13g2_a21oi_1 _10303_ (.A1(_02762_),
    .A2(_02752_),
    .Y(_00574_),
    .B1(_02763_));
 sg13g2_nand2_1 _10304_ (.Y(_02764_),
    .A(net224),
    .B(\ppu.sprite_buffer.attr_y[0][14] ));
 sg13g2_o21ai_1 _10305_ (.B1(_02764_),
    .Y(_00575_),
    .A1(net336),
    .A2(net224));
 sg13g2_nand2_1 _10306_ (.Y(_02765_),
    .A(net224),
    .B(\ppu.sprite_buffer.attr_y[0][15] ));
 sg13g2_o21ai_1 _10307_ (.B1(_02765_),
    .Y(_00576_),
    .A1(_02688_),
    .A2(net224));
 sg13g2_inv_1 _10308_ (.Y(_02766_),
    .A(\ppu.sprite_buffer.attr_y[0][1] ));
 sg13g2_nor2_1 _10309_ (.A(\ppu.sprite_buffer.attr_y[0][5] ),
    .B(net223),
    .Y(_02767_));
 sg13g2_a21oi_1 _10310_ (.A1(_02766_),
    .A2(net225),
    .Y(_00577_),
    .B1(_02767_));
 sg13g2_inv_1 _10311_ (.Y(_02768_),
    .A(\ppu.sprite_buffer.attr_y[0][2] ));
 sg13g2_nor2_1 _10312_ (.A(\ppu.sprite_buffer.attr_y[0][6] ),
    .B(net223),
    .Y(_02769_));
 sg13g2_a21oi_1 _10313_ (.A1(_02768_),
    .A2(net225),
    .Y(_00578_),
    .B1(_02769_));
 sg13g2_inv_1 _10314_ (.Y(_02770_),
    .A(\ppu.sprite_buffer.attr_y[0][4] ));
 sg13g2_nor2_1 _10315_ (.A(\ppu.sprite_buffer.attr_y[0][8] ),
    .B(net223),
    .Y(_02771_));
 sg13g2_a21oi_1 _10316_ (.A1(_02770_),
    .A2(net225),
    .Y(_00579_),
    .B1(_02771_));
 sg13g2_inv_1 _10317_ (.Y(_02772_),
    .A(\ppu.sprite_buffer.attr_y[0][5] ));
 sg13g2_nor2_1 _10318_ (.A(\ppu.sprite_buffer.attr_y[0][9] ),
    .B(net223),
    .Y(_02773_));
 sg13g2_a21oi_1 _10319_ (.A1(_02772_),
    .A2(_02752_),
    .Y(_00580_),
    .B1(_02773_));
 sg13g2_inv_1 _10320_ (.Y(_02774_),
    .A(\ppu.sprite_buffer.attr_y[0][6] ));
 sg13g2_nor2_1 _10321_ (.A(\ppu.sprite_buffer.attr_y[0][10] ),
    .B(_02760_),
    .Y(_02775_));
 sg13g2_a21oi_1 _10322_ (.A1(_02774_),
    .A2(net225),
    .Y(_00581_),
    .B1(_02775_));
 sg13g2_inv_1 _10323_ (.Y(_02776_),
    .A(\ppu.sprite_buffer.attr_y[0][7] ));
 sg13g2_nor2_1 _10324_ (.A(\ppu.sprite_buffer.attr_y[0][11] ),
    .B(net223),
    .Y(_02777_));
 sg13g2_a21oi_1 _10325_ (.A1(_02776_),
    .A2(net224),
    .Y(_00582_),
    .B1(_02777_));
 sg13g2_inv_1 _10326_ (.Y(_02778_),
    .A(\ppu.sprite_buffer.attr_y[0][8] ));
 sg13g2_nor2_1 _10327_ (.A(\ppu.sprite_buffer.attr_y[0][12] ),
    .B(net223),
    .Y(_02779_));
 sg13g2_a21oi_1 _10328_ (.A1(_02778_),
    .A2(_02753_),
    .Y(_00583_),
    .B1(_02779_));
 sg13g2_inv_1 _10329_ (.Y(_02780_),
    .A(\ppu.sprite_buffer.attr_y[0][9] ));
 sg13g2_nor2_1 _10330_ (.A(\ppu.sprite_buffer.attr_y[0][13] ),
    .B(_02760_),
    .Y(_02781_));
 sg13g2_a21oi_1 _10331_ (.A1(_02780_),
    .A2(_02753_),
    .Y(_00584_),
    .B1(_02781_));
 sg13g2_nand3_1 _10332_ (.B(_02566_),
    .C(_00061_),
    .A(_02670_),
    .Y(_02782_));
 sg13g2_buf_1 _10333_ (.A(_02782_),
    .X(_02783_));
 sg13g2_buf_1 _10334_ (.A(_02783_),
    .X(_02784_));
 sg13g2_mux2_1 _10335_ (.A0(\ppu.sprite_buffer.attr_y[1][4] ),
    .A1(\ppu.sprite_buffer.attr_y[1][0] ),
    .S(net222),
    .X(_00585_));
 sg13g2_inv_1 _10336_ (.Y(_02785_),
    .A(\ppu.sprite_buffer.attr_y[1][10] ));
 sg13g2_buf_1 _10337_ (.A(_02783_),
    .X(_02786_));
 sg13g2_nor2_1 _10338_ (.A(\ppu.sprite_buffer.attr_y[1][14] ),
    .B(_02783_),
    .Y(_02787_));
 sg13g2_a21oi_1 _10339_ (.A1(_02785_),
    .A2(net221),
    .Y(_00586_),
    .B1(_02787_));
 sg13g2_inv_1 _10340_ (.Y(_02788_),
    .A(\ppu.sprite_buffer.attr_y[1][11] ));
 sg13g2_nor2_1 _10341_ (.A(\ppu.sprite_buffer.attr_y[1][15] ),
    .B(_02783_),
    .Y(_02789_));
 sg13g2_a21oi_1 _10342_ (.A1(_02788_),
    .A2(net221),
    .Y(_00587_),
    .B1(_02789_));
 sg13g2_inv_1 _10343_ (.Y(_02790_),
    .A(\ppu.sprite_buffer.attr_y[1][12] ));
 sg13g2_nor2_1 _10344_ (.A(_02485_),
    .B(_02783_),
    .Y(_02791_));
 sg13g2_a21oi_1 _10345_ (.A1(_02790_),
    .A2(net221),
    .Y(_00588_),
    .B1(_02791_));
 sg13g2_inv_1 _10346_ (.Y(_02792_),
    .A(\ppu.sprite_buffer.attr_y[1][13] ));
 sg13g2_nor2_1 _10347_ (.A(net383),
    .B(_02783_),
    .Y(_02793_));
 sg13g2_a21oi_1 _10348_ (.A1(_02792_),
    .A2(net221),
    .Y(_00589_),
    .B1(_02793_));
 sg13g2_nand2_1 _10349_ (.Y(_02794_),
    .A(net222),
    .B(\ppu.sprite_buffer.attr_y[1][14] ));
 sg13g2_o21ai_1 _10350_ (.B1(_02794_),
    .Y(_00590_),
    .A1(_02686_),
    .A2(net221));
 sg13g2_nand2_1 _10351_ (.Y(_02795_),
    .A(net222),
    .B(\ppu.sprite_buffer.attr_y[1][15] ));
 sg13g2_o21ai_1 _10352_ (.B1(_02795_),
    .Y(_00591_),
    .A1(net335),
    .A2(net221));
 sg13g2_mux2_1 _10353_ (.A0(\ppu.sprite_buffer.attr_y[1][5] ),
    .A1(\ppu.sprite_buffer.attr_y[1][1] ),
    .S(net222),
    .X(_00592_));
 sg13g2_mux2_1 _10354_ (.A0(\ppu.sprite_buffer.attr_y[1][6] ),
    .A1(\ppu.sprite_buffer.attr_y[1][2] ),
    .S(net222),
    .X(_00593_));
 sg13g2_mux2_1 _10355_ (.A0(\ppu.sprite_buffer.attr_y[1][8] ),
    .A1(\ppu.sprite_buffer.attr_y[1][4] ),
    .S(net222),
    .X(_00594_));
 sg13g2_mux2_1 _10356_ (.A0(\ppu.sprite_buffer.attr_y[1][9] ),
    .A1(\ppu.sprite_buffer.attr_y[1][5] ),
    .S(_02784_),
    .X(_00595_));
 sg13g2_nand2_1 _10357_ (.Y(_02796_),
    .A(net222),
    .B(\ppu.sprite_buffer.attr_y[1][6] ));
 sg13g2_o21ai_1 _10358_ (.B1(_02796_),
    .Y(_00596_),
    .A1(_02785_),
    .A2(_02786_));
 sg13g2_nand2_1 _10359_ (.Y(_02797_),
    .A(net222),
    .B(\ppu.sprite_buffer.attr_y[1][7] ));
 sg13g2_o21ai_1 _10360_ (.B1(_02797_),
    .Y(_00597_),
    .A1(_02788_),
    .A2(_02786_));
 sg13g2_nand2_1 _10361_ (.Y(_02798_),
    .A(_02784_),
    .B(\ppu.sprite_buffer.attr_y[1][8] ));
 sg13g2_o21ai_1 _10362_ (.B1(_02798_),
    .Y(_00598_),
    .A1(_02790_),
    .A2(net221));
 sg13g2_nand2_1 _10363_ (.Y(_02799_),
    .A(_02783_),
    .B(\ppu.sprite_buffer.attr_y[1][9] ));
 sg13g2_o21ai_1 _10364_ (.B1(_02799_),
    .Y(_00599_),
    .A1(_02792_),
    .A2(net221));
 sg13g2_inv_1 _10365_ (.Y(_02800_),
    .A(\ppu.sprite_buffer.id_buffer[0][0] ));
 sg13g2_nor2_1 _10366_ (.A(_01890_),
    .B(_01870_),
    .Y(_02801_));
 sg13g2_nand2_1 _10367_ (.Y(_02802_),
    .A(_01884_),
    .B(_02801_));
 sg13g2_inv_1 _10368_ (.Y(_02803_),
    .A(_02802_));
 sg13g2_nand3_1 _10369_ (.B(_01875_),
    .C(_01873_),
    .A(_02803_),
    .Y(_02804_));
 sg13g2_buf_1 _10370_ (.A(_02804_),
    .X(_02805_));
 sg13g2_buf_1 _10371_ (.A(_02805_),
    .X(_02806_));
 sg13g2_buf_1 _10372_ (.A(\ppu.sprite_buffer.data8[0] ),
    .X(_02807_));
 sg13g2_nor2_1 _10373_ (.A(_02807_),
    .B(net144),
    .Y(_02808_));
 sg13g2_a21oi_1 _10374_ (.A1(_02800_),
    .A2(net144),
    .Y(_00603_),
    .B1(_02808_));
 sg13g2_inv_1 _10375_ (.Y(_02809_),
    .A(\ppu.sprite_buffer.id_buffer[0][1] ));
 sg13g2_buf_2 _10376_ (.A(\ppu.sprite_buffer.data8[1] ),
    .X(_02810_));
 sg13g2_nor2_1 _10377_ (.A(_02810_),
    .B(_02806_),
    .Y(_02811_));
 sg13g2_a21oi_1 _10378_ (.A1(_02809_),
    .A2(net144),
    .Y(_00604_),
    .B1(_02811_));
 sg13g2_inv_1 _10379_ (.Y(_02812_),
    .A(\ppu.sprite_buffer.id_buffer[0][2] ));
 sg13g2_buf_2 _10380_ (.A(\ppu.sprite_buffer.data8[2] ),
    .X(_02813_));
 sg13g2_nor2_1 _10381_ (.A(_02813_),
    .B(_02806_),
    .Y(_02814_));
 sg13g2_a21oi_1 _10382_ (.A1(_02812_),
    .A2(net144),
    .Y(_00605_),
    .B1(_02814_));
 sg13g2_inv_1 _10383_ (.Y(_02815_),
    .A(\ppu.sprite_buffer.id_buffer[0][3] ));
 sg13g2_buf_2 _10384_ (.A(\ppu.sprite_buffer.data8[3] ),
    .X(_02816_));
 sg13g2_nor2_1 _10385_ (.A(_02816_),
    .B(net144),
    .Y(_02817_));
 sg13g2_a21oi_1 _10386_ (.A1(_02815_),
    .A2(net144),
    .Y(_00606_),
    .B1(_02817_));
 sg13g2_inv_1 _10387_ (.Y(_02818_),
    .A(\ppu.sprite_buffer.id_buffer[0][4] ));
 sg13g2_nor2_1 _10388_ (.A(_02485_),
    .B(_02805_),
    .Y(_02819_));
 sg13g2_a21oi_1 _10389_ (.A1(_02818_),
    .A2(net144),
    .Y(_00607_),
    .B1(_02819_));
 sg13g2_inv_1 _10390_ (.Y(_02820_),
    .A(\ppu.sprite_buffer.id_buffer[0][5] ));
 sg13g2_nor2_1 _10391_ (.A(_02494_),
    .B(_02805_),
    .Y(_02821_));
 sg13g2_a21oi_1 _10392_ (.A1(_02820_),
    .A2(net144),
    .Y(_00608_),
    .B1(_02821_));
 sg13g2_inv_1 _10393_ (.Y(_02822_),
    .A(\ppu.sprite_buffer.id_buffer[1][0] ));
 sg13g2_nand2_1 _10394_ (.Y(_02823_),
    .A(_02803_),
    .B(_01876_));
 sg13g2_buf_1 _10395_ (.A(_02823_),
    .X(_02824_));
 sg13g2_nor2_1 _10396_ (.A(_02807_),
    .B(net163),
    .Y(_02825_));
 sg13g2_a21oi_1 _10397_ (.A1(_02822_),
    .A2(net163),
    .Y(_00609_),
    .B1(_02825_));
 sg13g2_inv_1 _10398_ (.Y(_02826_),
    .A(\ppu.sprite_buffer.id_buffer[1][1] ));
 sg13g2_nor2_1 _10399_ (.A(_02810_),
    .B(net163),
    .Y(_02827_));
 sg13g2_a21oi_1 _10400_ (.A1(_02826_),
    .A2(net163),
    .Y(_00610_),
    .B1(_02827_));
 sg13g2_inv_1 _10401_ (.Y(_02828_),
    .A(\ppu.sprite_buffer.id_buffer[1][2] ));
 sg13g2_nor2_1 _10402_ (.A(_02813_),
    .B(net163),
    .Y(_02829_));
 sg13g2_a21oi_1 _10403_ (.A1(_02828_),
    .A2(net163),
    .Y(_00611_),
    .B1(_02829_));
 sg13g2_inv_1 _10404_ (.Y(_02830_),
    .A(\ppu.sprite_buffer.id_buffer[1][3] ));
 sg13g2_nor2_1 _10405_ (.A(_02816_),
    .B(net163),
    .Y(_02831_));
 sg13g2_a21oi_1 _10406_ (.A1(_02830_),
    .A2(net163),
    .Y(_00612_),
    .B1(_02831_));
 sg13g2_inv_1 _10407_ (.Y(_02832_),
    .A(\ppu.sprite_buffer.id_buffer[1][4] ));
 sg13g2_nor2_1 _10408_ (.A(net405),
    .B(_02823_),
    .Y(_02833_));
 sg13g2_a21oi_1 _10409_ (.A1(_02832_),
    .A2(_02824_),
    .Y(_00613_),
    .B1(_02833_));
 sg13g2_inv_1 _10410_ (.Y(_02834_),
    .A(\ppu.sprite_buffer.id_buffer[1][5] ));
 sg13g2_nor2_1 _10411_ (.A(_02494_),
    .B(_02823_),
    .Y(_02835_));
 sg13g2_a21oi_1 _10412_ (.A1(_02834_),
    .A2(_02824_),
    .Y(_00614_),
    .B1(_02835_));
 sg13g2_inv_1 _10413_ (.Y(_02836_),
    .A(\ppu.sprite_buffer.id_buffer[2][0] ));
 sg13g2_nand2_1 _10414_ (.Y(_02837_),
    .A(_02803_),
    .B(_01874_));
 sg13g2_buf_1 _10415_ (.A(_02837_),
    .X(_02838_));
 sg13g2_nor2_1 _10416_ (.A(_02807_),
    .B(net162),
    .Y(_02839_));
 sg13g2_a21oi_1 _10417_ (.A1(_02836_),
    .A2(net162),
    .Y(_00615_),
    .B1(_02839_));
 sg13g2_inv_1 _10418_ (.Y(_02840_),
    .A(\ppu.sprite_buffer.id_buffer[2][1] ));
 sg13g2_nor2_1 _10419_ (.A(_02810_),
    .B(_02838_),
    .Y(_02841_));
 sg13g2_a21oi_1 _10420_ (.A1(_02840_),
    .A2(net162),
    .Y(_00616_),
    .B1(_02841_));
 sg13g2_inv_1 _10421_ (.Y(_02842_),
    .A(\ppu.sprite_buffer.id_buffer[2][2] ));
 sg13g2_nor2_1 _10422_ (.A(_02813_),
    .B(_02838_),
    .Y(_02843_));
 sg13g2_a21oi_1 _10423_ (.A1(_02842_),
    .A2(net162),
    .Y(_00617_),
    .B1(_02843_));
 sg13g2_inv_1 _10424_ (.Y(_02844_),
    .A(\ppu.sprite_buffer.id_buffer[2][3] ));
 sg13g2_nor2_1 _10425_ (.A(_02816_),
    .B(net162),
    .Y(_02845_));
 sg13g2_a21oi_1 _10426_ (.A1(_02844_),
    .A2(net162),
    .Y(_00618_),
    .B1(_02845_));
 sg13g2_inv_1 _10427_ (.Y(_02846_),
    .A(\ppu.sprite_buffer.id_buffer[2][4] ));
 sg13g2_nor2_1 _10428_ (.A(net405),
    .B(_02837_),
    .Y(_02847_));
 sg13g2_a21oi_1 _10429_ (.A1(_02846_),
    .A2(net162),
    .Y(_00619_),
    .B1(_02847_));
 sg13g2_inv_1 _10430_ (.Y(_02848_),
    .A(\ppu.sprite_buffer.id_buffer[2][5] ));
 sg13g2_nor2_1 _10431_ (.A(_02493_),
    .B(_02837_),
    .Y(_02849_));
 sg13g2_a21oi_1 _10432_ (.A1(_02848_),
    .A2(net162),
    .Y(_00620_),
    .B1(_02849_));
 sg13g2_inv_1 _10433_ (.Y(_02850_),
    .A(\ppu.sprite_buffer.id_buffer[3][0] ));
 sg13g2_nor2_1 _10434_ (.A(_01875_),
    .B(_02802_),
    .Y(_02851_));
 sg13g2_nand2_1 _10435_ (.Y(_02852_),
    .A(_02851_),
    .B(_01872_));
 sg13g2_buf_1 _10436_ (.A(_02852_),
    .X(_02853_));
 sg13g2_nor2_1 _10437_ (.A(_02807_),
    .B(net161),
    .Y(_02854_));
 sg13g2_a21oi_1 _10438_ (.A1(_02850_),
    .A2(net161),
    .Y(_00621_),
    .B1(_02854_));
 sg13g2_inv_1 _10439_ (.Y(_02855_),
    .A(\ppu.sprite_buffer.id_buffer[3][1] ));
 sg13g2_nor2_1 _10440_ (.A(_02810_),
    .B(net161),
    .Y(_02856_));
 sg13g2_a21oi_1 _10441_ (.A1(_02855_),
    .A2(_02853_),
    .Y(_00622_),
    .B1(_02856_));
 sg13g2_inv_1 _10442_ (.Y(_02857_),
    .A(\ppu.sprite_buffer.id_buffer[3][2] ));
 sg13g2_nor2_1 _10443_ (.A(_02813_),
    .B(net161),
    .Y(_02858_));
 sg13g2_a21oi_1 _10444_ (.A1(_02857_),
    .A2(_02853_),
    .Y(_00623_),
    .B1(_02858_));
 sg13g2_inv_1 _10445_ (.Y(_02859_),
    .A(\ppu.sprite_buffer.id_buffer[3][3] ));
 sg13g2_nor2_1 _10446_ (.A(_02816_),
    .B(net161),
    .Y(_02860_));
 sg13g2_a21oi_1 _10447_ (.A1(_02859_),
    .A2(net161),
    .Y(_00624_),
    .B1(_02860_));
 sg13g2_inv_1 _10448_ (.Y(_02861_),
    .A(\ppu.sprite_buffer.id_buffer[3][4] ));
 sg13g2_nor2_1 _10449_ (.A(_02484_),
    .B(_02852_),
    .Y(_02862_));
 sg13g2_a21oi_1 _10450_ (.A1(_02861_),
    .A2(net161),
    .Y(_00625_),
    .B1(_02862_));
 sg13g2_inv_1 _10451_ (.Y(_02863_),
    .A(\ppu.sprite_buffer.id_buffer[3][5] ));
 sg13g2_nor2_1 _10452_ (.A(_02493_),
    .B(_02852_),
    .Y(_02864_));
 sg13g2_a21oi_1 _10453_ (.A1(_02863_),
    .A2(net161),
    .Y(_00626_),
    .B1(_02864_));
 sg13g2_nand3_1 _10454_ (.B(\ppu.sprite_buffer.extra_sorted_addr_bits[2] ),
    .C(\ppu.sprite_buffer.extra_sorted_addr_bits[1] ),
    .A(_01858_),
    .Y(_02865_));
 sg13g2_buf_1 _10455_ (.A(\ppu.sprite_buffer.extra_sorted_addr_bits[0] ),
    .X(_02866_));
 sg13g2_nand2_1 _10456_ (.Y(_02867_),
    .A(_02866_),
    .B(\ppu.sprite_buffer.out_counters[0][2] ));
 sg13g2_nor2b_1 _10457_ (.A(_02600_),
    .B_N(_02573_),
    .Y(_02868_));
 sg13g2_nor2_1 _10458_ (.A(_01888_),
    .B(_02868_),
    .Y(_02869_));
 sg13g2_nor2_1 _10459_ (.A(_01890_),
    .B(_01885_),
    .Y(_02870_));
 sg13g2_a21oi_1 _10460_ (.A1(_02868_),
    .A2(_02870_),
    .Y(_02871_),
    .B1(_02869_));
 sg13g2_nor2_1 _10461_ (.A(_00079_),
    .B(_02871_),
    .Y(_02872_));
 sg13g2_xnor2_1 _10462_ (.Y(_02873_),
    .A(_00078_),
    .B(_02869_));
 sg13g2_nand2_1 _10463_ (.Y(_02874_),
    .A(_02872_),
    .B(_02873_));
 sg13g2_inv_1 _10464_ (.Y(_02875_),
    .A(_02874_));
 sg13g2_a21oi_1 _10465_ (.A1(\ppu.sprite_buffer.out_counters[0][1] ),
    .A2(_02869_),
    .Y(_02876_),
    .B1(_02875_));
 sg13g2_nor2_1 _10466_ (.A(_02867_),
    .B(_02876_),
    .Y(_02877_));
 sg13g2_inv_1 _10467_ (.Y(_02878_),
    .A(_02877_));
 sg13g2_o21ai_1 _10468_ (.B1(\ppu.sprite_buffer.scan_enabled ),
    .Y(_02879_),
    .A1(_02865_),
    .A2(_02878_));
 sg13g2_nor2_1 _10469_ (.A(_01887_),
    .B(_01851_),
    .Y(_02880_));
 sg13g2_buf_1 _10470_ (.A(net258),
    .X(_02881_));
 sg13g2_a21oi_1 _10471_ (.A1(_02879_),
    .A2(_02880_),
    .Y(_00645_),
    .B1(net247));
 sg13g2_nor2_1 _10472_ (.A(_02579_),
    .B(_02602_),
    .Y(_02882_));
 sg13g2_buf_2 _10473_ (.A(_02882_),
    .X(_02883_));
 sg13g2_inv_1 _10474_ (.Y(_02884_),
    .A(_02883_));
 sg13g2_nor2_1 _10475_ (.A(_02587_),
    .B(_02884_),
    .Y(_02885_));
 sg13g2_nor2_1 _10476_ (.A(_01878_),
    .B(_02563_),
    .Y(_02886_));
 sg13g2_buf_2 _10477_ (.A(_02886_),
    .X(_02887_));
 sg13g2_nand2_1 _10478_ (.Y(_02888_),
    .A(_02885_),
    .B(_02887_));
 sg13g2_buf_1 _10479_ (.A(_02888_),
    .X(_02889_));
 sg13g2_nand2_1 _10480_ (.Y(_02890_),
    .A(net89),
    .B(\ppu.sprite_buffer.sprite_ids[0][0] ));
 sg13g2_o21ai_1 _10481_ (.B1(_02890_),
    .Y(_00646_),
    .A1(_02800_),
    .A2(net89));
 sg13g2_nand2_1 _10482_ (.Y(_02891_),
    .A(net89),
    .B(\ppu.sprite_buffer.sprite_ids[0][1] ));
 sg13g2_o21ai_1 _10483_ (.B1(_02891_),
    .Y(_00647_),
    .A1(_02809_),
    .A2(net89));
 sg13g2_nand2_1 _10484_ (.Y(_02892_),
    .A(net89),
    .B(\ppu.sprite_buffer.sprite_ids[0][2] ));
 sg13g2_o21ai_1 _10485_ (.B1(_02892_),
    .Y(_00648_),
    .A1(_02812_),
    .A2(net89));
 sg13g2_nand2_1 _10486_ (.Y(_02893_),
    .A(net89),
    .B(\ppu.sprite_buffer.sprite_ids[0][3] ));
 sg13g2_o21ai_1 _10487_ (.B1(_02893_),
    .Y(_00649_),
    .A1(_02815_),
    .A2(net89));
 sg13g2_nand2_1 _10488_ (.Y(_02894_),
    .A(_02888_),
    .B(\ppu.sprite_buffer.sprite_ids[0][4] ));
 sg13g2_o21ai_1 _10489_ (.B1(_02894_),
    .Y(_00650_),
    .A1(_02818_),
    .A2(_02889_));
 sg13g2_nand2_1 _10490_ (.Y(_02895_),
    .A(_02888_),
    .B(\ppu.sprite_buffer.sprite_ids[0][5] ));
 sg13g2_o21ai_1 _10491_ (.B1(_02895_),
    .Y(_00651_),
    .A1(_02820_),
    .A2(_02889_));
 sg13g2_inv_1 _10492_ (.Y(_02896_),
    .A(_02563_));
 sg13g2_nand2_1 _10493_ (.Y(_02897_),
    .A(_02896_),
    .B(_01878_));
 sg13g2_inv_2 _10494_ (.Y(_02898_),
    .A(_02897_));
 sg13g2_nand2_1 _10495_ (.Y(_02899_),
    .A(_02885_),
    .B(_02898_));
 sg13g2_buf_1 _10496_ (.A(_02899_),
    .X(_02900_));
 sg13g2_nand2_1 _10497_ (.Y(_02901_),
    .A(net88),
    .B(\ppu.sprite_buffer.sprite_ids[1][0] ));
 sg13g2_o21ai_1 _10498_ (.B1(_02901_),
    .Y(_00652_),
    .A1(_02822_),
    .A2(net88));
 sg13g2_nand2_1 _10499_ (.Y(_02902_),
    .A(_02900_),
    .B(\ppu.sprite_buffer.sprite_ids[1][1] ));
 sg13g2_o21ai_1 _10500_ (.B1(_02902_),
    .Y(_00653_),
    .A1(_02826_),
    .A2(net88));
 sg13g2_nand2_1 _10501_ (.Y(_02903_),
    .A(_02900_),
    .B(\ppu.sprite_buffer.sprite_ids[1][2] ));
 sg13g2_o21ai_1 _10502_ (.B1(_02903_),
    .Y(_00654_),
    .A1(_02828_),
    .A2(net88));
 sg13g2_nand2_1 _10503_ (.Y(_02904_),
    .A(net88),
    .B(\ppu.sprite_buffer.sprite_ids[1][3] ));
 sg13g2_o21ai_1 _10504_ (.B1(_02904_),
    .Y(_00655_),
    .A1(_02830_),
    .A2(net88));
 sg13g2_nand2_1 _10505_ (.Y(_02905_),
    .A(_02899_),
    .B(\ppu.sprite_buffer.sprite_ids[1][4] ));
 sg13g2_o21ai_1 _10506_ (.B1(_02905_),
    .Y(_00656_),
    .A1(_02832_),
    .A2(net88));
 sg13g2_nand2_1 _10507_ (.Y(_02906_),
    .A(_02899_),
    .B(\ppu.sprite_buffer.sprite_ids[1][5] ));
 sg13g2_o21ai_1 _10508_ (.B1(_02906_),
    .Y(_00657_),
    .A1(_02834_),
    .A2(net88));
 sg13g2_nor2_1 _10509_ (.A(_01878_),
    .B(_02896_),
    .Y(_02907_));
 sg13g2_buf_2 _10510_ (.A(_02907_),
    .X(_02908_));
 sg13g2_nand2_1 _10511_ (.Y(_02909_),
    .A(_02885_),
    .B(_02908_));
 sg13g2_buf_1 _10512_ (.A(_02909_),
    .X(_02910_));
 sg13g2_nand2_1 _10513_ (.Y(_02911_),
    .A(net87),
    .B(\ppu.sprite_buffer.sprite_ids[2][0] ));
 sg13g2_o21ai_1 _10514_ (.B1(_02911_),
    .Y(_00658_),
    .A1(_02836_),
    .A2(net87));
 sg13g2_nand2_1 _10515_ (.Y(_02912_),
    .A(net87),
    .B(\ppu.sprite_buffer.sprite_ids[2][1] ));
 sg13g2_o21ai_1 _10516_ (.B1(_02912_),
    .Y(_00659_),
    .A1(_02840_),
    .A2(net87));
 sg13g2_nand2_1 _10517_ (.Y(_02913_),
    .A(_02910_),
    .B(\ppu.sprite_buffer.sprite_ids[2][2] ));
 sg13g2_o21ai_1 _10518_ (.B1(_02913_),
    .Y(_00660_),
    .A1(_02842_),
    .A2(_02910_));
 sg13g2_nand2_1 _10519_ (.Y(_02914_),
    .A(net87),
    .B(\ppu.sprite_buffer.sprite_ids[2][3] ));
 sg13g2_o21ai_1 _10520_ (.B1(_02914_),
    .Y(_00661_),
    .A1(_02844_),
    .A2(net87));
 sg13g2_nand2_1 _10521_ (.Y(_02915_),
    .A(_02909_),
    .B(\ppu.sprite_buffer.sprite_ids[2][4] ));
 sg13g2_o21ai_1 _10522_ (.B1(_02915_),
    .Y(_00662_),
    .A1(_02846_),
    .A2(net87));
 sg13g2_nand2_1 _10523_ (.Y(_02916_),
    .A(_02909_),
    .B(\ppu.sprite_buffer.sprite_ids[2][5] ));
 sg13g2_o21ai_1 _10524_ (.B1(_02916_),
    .Y(_00663_),
    .A1(_02848_),
    .A2(net87));
 sg13g2_nand2_1 _10525_ (.Y(_02917_),
    .A(_01878_),
    .B(_02563_));
 sg13g2_inv_2 _10526_ (.Y(_02918_),
    .A(_02917_));
 sg13g2_nand2_1 _10527_ (.Y(_02919_),
    .A(_02885_),
    .B(_02918_));
 sg13g2_buf_1 _10528_ (.A(_02919_),
    .X(_02920_));
 sg13g2_nand2_1 _10529_ (.Y(_02921_),
    .A(net86),
    .B(\ppu.sprite_buffer.sprite_ids[3][0] ));
 sg13g2_o21ai_1 _10530_ (.B1(_02921_),
    .Y(_00664_),
    .A1(_02850_),
    .A2(net86));
 sg13g2_nand2_1 _10531_ (.Y(_02922_),
    .A(net86),
    .B(\ppu.sprite_buffer.sprite_ids[3][1] ));
 sg13g2_o21ai_1 _10532_ (.B1(_02922_),
    .Y(_00665_),
    .A1(_02855_),
    .A2(net86));
 sg13g2_nand2_1 _10533_ (.Y(_02923_),
    .A(_02920_),
    .B(\ppu.sprite_buffer.sprite_ids[3][2] ));
 sg13g2_o21ai_1 _10534_ (.B1(_02923_),
    .Y(_00666_),
    .A1(_02857_),
    .A2(_02920_));
 sg13g2_nand2_1 _10535_ (.Y(_02924_),
    .A(net86),
    .B(\ppu.sprite_buffer.sprite_ids[3][3] ));
 sg13g2_o21ai_1 _10536_ (.B1(_02924_),
    .Y(_00667_),
    .A1(_02859_),
    .A2(net86));
 sg13g2_nand2_1 _10537_ (.Y(_02925_),
    .A(_02919_),
    .B(\ppu.sprite_buffer.sprite_ids[3][4] ));
 sg13g2_o21ai_1 _10538_ (.B1(_02925_),
    .Y(_00668_),
    .A1(_02861_),
    .A2(net86));
 sg13g2_nand2_1 _10539_ (.Y(_02926_),
    .A(_02919_),
    .B(\ppu.sprite_buffer.sprite_ids[3][5] ));
 sg13g2_o21ai_1 _10540_ (.B1(_02926_),
    .Y(_00669_),
    .A1(_02863_),
    .A2(net86));
 sg13g2_buf_1 _10541_ (.A(net262),
    .X(_02927_));
 sg13g2_mux2_1 _10542_ (.A0(\ppu.sprite_buffer.top_color[0] ),
    .A1(\ppu.pixel_out_s[0] ),
    .S(net246),
    .X(_00670_));
 sg13g2_mux2_1 _10543_ (.A0(\ppu.sprite_buffer.top_color[1] ),
    .A1(\ppu.pixel_out_s[1] ),
    .S(net246),
    .X(_00671_));
 sg13g2_mux2_1 _10544_ (.A0(\ppu.sprite_buffer.top_color[2] ),
    .A1(\ppu.pixel_out_s[2] ),
    .S(net246),
    .X(_00672_));
 sg13g2_mux2_1 _10545_ (.A0(\ppu.sprite_buffer.top_color[3] ),
    .A1(\ppu.pixel_out_s[3] ),
    .S(net246),
    .X(_00673_));
 sg13g2_mux2_1 _10546_ (.A0(\ppu.sprite_buffer.top_depth[0] ),
    .A1(\ppu.depth_out_s[0] ),
    .S(net246),
    .X(_00674_));
 sg13g2_inv_1 _10547_ (.Y(_02928_),
    .A(\ppu.depth_out_s[1] ));
 sg13g2_nor2_1 _10548_ (.A(\ppu.sprite_buffer.top_depth[1] ),
    .B(net246),
    .Y(_02929_));
 sg13g2_a21oi_1 _10549_ (.A1(_02928_),
    .A2(net246),
    .Y(_00675_),
    .B1(_02929_));
 sg13g2_nand3_1 _10550_ (.B(_02177_),
    .C(_02184_),
    .A(_02183_),
    .Y(_02930_));
 sg13g2_buf_2 _10551_ (.A(_02930_),
    .X(_02931_));
 sg13g2_buf_1 _10552_ (.A(_02931_),
    .X(_02932_));
 sg13g2_mux2_1 _10553_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][0] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][4] ),
    .S(_02932_),
    .X(_00676_));
 sg13g2_mux2_1 _10554_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][10] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][14] ),
    .S(net61),
    .X(_00677_));
 sg13g2_mux2_1 _10555_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][11] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][15] ),
    .S(net61),
    .X(_00678_));
 sg13g2_mux2_1 _10556_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][12] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][16] ),
    .S(net61),
    .X(_00679_));
 sg13g2_mux2_1 _10557_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][13] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][17] ),
    .S(net61),
    .X(_00680_));
 sg13g2_mux2_1 _10558_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][14] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][18] ),
    .S(net61),
    .X(_00681_));
 sg13g2_mux2_1 _10559_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][15] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][19] ),
    .S(net61),
    .X(_00682_));
 sg13g2_mux2_1 _10560_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][16] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][20] ),
    .S(net61),
    .X(_00683_));
 sg13g2_buf_2 _10561_ (.A(_02931_),
    .X(_02933_));
 sg13g2_mux2_1 _10562_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][17] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][21] ),
    .S(net60),
    .X(_00684_));
 sg13g2_mux2_1 _10563_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][18] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][22] ),
    .S(net60),
    .X(_00685_));
 sg13g2_mux2_1 _10564_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][19] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][23] ),
    .S(net60),
    .X(_00686_));
 sg13g2_mux2_1 _10565_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][1] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][5] ),
    .S(_02933_),
    .X(_00687_));
 sg13g2_mux2_1 _10566_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][20] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][24] ),
    .S(net60),
    .X(_00688_));
 sg13g2_mux2_1 _10567_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][21] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][25] ),
    .S(net60),
    .X(_00689_));
 sg13g2_mux2_1 _10568_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][22] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][26] ),
    .S(net60),
    .X(_00690_));
 sg13g2_mux2_1 _10569_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][23] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][27] ),
    .S(_02933_),
    .X(_00691_));
 sg13g2_mux2_1 _10570_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][24] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][28] ),
    .S(net60),
    .X(_00692_));
 sg13g2_mux2_1 _10571_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][25] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][29] ),
    .S(net60),
    .X(_00693_));
 sg13g2_buf_1 _10572_ (.A(_02931_),
    .X(_02934_));
 sg13g2_mux2_1 _10573_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][26] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][30] ),
    .S(net59),
    .X(_00694_));
 sg13g2_mux2_1 _10574_ (.A0(\ppu.sprite_buffer.sprite_pixels[0][27] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[0][31] ),
    .S(net59),
    .X(_00695_));
 sg13g2_buf_1 _10575_ (.A(_02931_),
    .X(_02935_));
 sg13g2_nor2_1 _10576_ (.A(\ppu.sprite_buffer.sprite_pixels[0][28] ),
    .B(net59),
    .Y(_02936_));
 sg13g2_a21oi_1 _10577_ (.A1(net381),
    .A2(net58),
    .Y(_00696_),
    .B1(_02936_));
 sg13g2_nor2_1 _10578_ (.A(\ppu.sprite_buffer.sprite_pixels[0][29] ),
    .B(net59),
    .Y(_02937_));
 sg13g2_a21oi_1 _10579_ (.A1(net382),
    .A2(net58),
    .Y(_00697_),
    .B1(_02937_));
 sg13g2_inv_1 _10580_ (.Y(_02938_),
    .A(\ppu.sprite_buffer.sprite_pixels[0][6] ));
 sg13g2_nor2_1 _10581_ (.A(\ppu.sprite_buffer.sprite_pixels[0][2] ),
    .B(_02934_),
    .Y(_02939_));
 sg13g2_a21oi_1 _10582_ (.A1(_02938_),
    .A2(net58),
    .Y(_00698_),
    .B1(_02939_));
 sg13g2_nor2_1 _10583_ (.A(\ppu.sprite_buffer.sprite_pixels[0][30] ),
    .B(net59),
    .Y(_02940_));
 sg13g2_a21oi_1 _10584_ (.A1(net336),
    .A2(net58),
    .Y(_00699_),
    .B1(_02940_));
 sg13g2_nor2_1 _10585_ (.A(\ppu.sprite_buffer.sprite_pixels[0][31] ),
    .B(_02931_),
    .Y(_02941_));
 sg13g2_a21oi_1 _10586_ (.A1(net335),
    .A2(net58),
    .Y(_00700_),
    .B1(_02941_));
 sg13g2_inv_1 _10587_ (.Y(_02942_),
    .A(\ppu.sprite_buffer.sprite_pixels[0][7] ));
 sg13g2_nor2_1 _10588_ (.A(\ppu.sprite_buffer.sprite_pixels[0][3] ),
    .B(_02931_),
    .Y(_02943_));
 sg13g2_a21oi_1 _10589_ (.A1(_02942_),
    .A2(net58),
    .Y(_00701_),
    .B1(_02943_));
 sg13g2_inv_1 _10590_ (.Y(_02944_),
    .A(\ppu.sprite_buffer.sprite_pixels[0][8] ));
 sg13g2_nor2_1 _10591_ (.A(\ppu.sprite_buffer.sprite_pixels[0][4] ),
    .B(_02931_),
    .Y(_02945_));
 sg13g2_a21oi_1 _10592_ (.A1(_02944_),
    .A2(net58),
    .Y(_00702_),
    .B1(_02945_));
 sg13g2_inv_1 _10593_ (.Y(_02946_),
    .A(\ppu.sprite_buffer.sprite_pixels[0][9] ));
 sg13g2_nor2_1 _10594_ (.A(\ppu.sprite_buffer.sprite_pixels[0][5] ),
    .B(_02931_),
    .Y(_02947_));
 sg13g2_a21oi_1 _10595_ (.A1(_02946_),
    .A2(_02935_),
    .Y(_00703_),
    .B1(_02947_));
 sg13g2_nand2_1 _10596_ (.Y(_02948_),
    .A(net59),
    .B(\ppu.sprite_buffer.sprite_pixels[0][10] ));
 sg13g2_o21ai_1 _10597_ (.B1(_02948_),
    .Y(_00704_),
    .A1(_02938_),
    .A2(net58));
 sg13g2_nand2_1 _10598_ (.Y(_02949_),
    .A(_02934_),
    .B(\ppu.sprite_buffer.sprite_pixels[0][11] ));
 sg13g2_o21ai_1 _10599_ (.B1(_02949_),
    .Y(_00705_),
    .A1(_02942_),
    .A2(_02935_));
 sg13g2_nand2_1 _10600_ (.Y(_02950_),
    .A(net59),
    .B(\ppu.sprite_buffer.sprite_pixels[0][12] ));
 sg13g2_o21ai_1 _10601_ (.B1(_02950_),
    .Y(_00706_),
    .A1(_02944_),
    .A2(_02932_));
 sg13g2_nand2_1 _10602_ (.Y(_02951_),
    .A(net59),
    .B(\ppu.sprite_buffer.sprite_pixels[0][13] ));
 sg13g2_o21ai_1 _10603_ (.B1(_02951_),
    .Y(_00707_),
    .A1(_02946_),
    .A2(net61));
 sg13g2_nand3_1 _10604_ (.B(_02158_),
    .C(_02164_),
    .A(_02163_),
    .Y(_02952_));
 sg13g2_buf_2 _10605_ (.A(_02952_),
    .X(_02953_));
 sg13g2_buf_1 _10606_ (.A(_02953_),
    .X(_02954_));
 sg13g2_mux2_1 _10607_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][0] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][4] ),
    .S(net57),
    .X(_00708_));
 sg13g2_mux2_1 _10608_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][10] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][14] ),
    .S(net57),
    .X(_00709_));
 sg13g2_mux2_1 _10609_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][11] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][15] ),
    .S(net57),
    .X(_00710_));
 sg13g2_mux2_1 _10610_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][12] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][16] ),
    .S(net57),
    .X(_00711_));
 sg13g2_mux2_1 _10611_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][13] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][17] ),
    .S(net57),
    .X(_00712_));
 sg13g2_mux2_1 _10612_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][14] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][18] ),
    .S(_02954_),
    .X(_00713_));
 sg13g2_mux2_1 _10613_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][15] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][19] ),
    .S(_02954_),
    .X(_00714_));
 sg13g2_mux2_1 _10614_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][16] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][20] ),
    .S(net57),
    .X(_00715_));
 sg13g2_buf_2 _10615_ (.A(_02953_),
    .X(_02955_));
 sg13g2_mux2_1 _10616_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][17] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][21] ),
    .S(net56),
    .X(_00716_));
 sg13g2_mux2_1 _10617_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][18] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][22] ),
    .S(net56),
    .X(_00717_));
 sg13g2_mux2_1 _10618_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][19] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][23] ),
    .S(_02955_),
    .X(_00718_));
 sg13g2_mux2_1 _10619_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][1] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][5] ),
    .S(net56),
    .X(_00719_));
 sg13g2_mux2_1 _10620_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][20] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][24] ),
    .S(net56),
    .X(_00720_));
 sg13g2_mux2_1 _10621_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][21] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][25] ),
    .S(net56),
    .X(_00721_));
 sg13g2_mux2_1 _10622_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][22] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][26] ),
    .S(net56),
    .X(_00722_));
 sg13g2_mux2_1 _10623_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][23] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][27] ),
    .S(_02955_),
    .X(_00723_));
 sg13g2_mux2_1 _10624_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][24] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][28] ),
    .S(net56),
    .X(_00724_));
 sg13g2_mux2_1 _10625_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][25] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][29] ),
    .S(net56),
    .X(_00725_));
 sg13g2_buf_1 _10626_ (.A(_02953_),
    .X(_02956_));
 sg13g2_mux2_1 _10627_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][26] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][30] ),
    .S(net55),
    .X(_00726_));
 sg13g2_mux2_1 _10628_ (.A0(\ppu.sprite_buffer.sprite_pixels[1][27] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][31] ),
    .S(_02956_),
    .X(_00727_));
 sg13g2_buf_1 _10629_ (.A(_02953_),
    .X(_02957_));
 sg13g2_nor2_1 _10630_ (.A(\ppu.sprite_buffer.sprite_pixels[1][28] ),
    .B(net55),
    .Y(_02958_));
 sg13g2_a21oi_1 _10631_ (.A1(net381),
    .A2(net54),
    .Y(_00728_),
    .B1(_02958_));
 sg13g2_nor2_1 _10632_ (.A(\ppu.sprite_buffer.sprite_pixels[1][29] ),
    .B(net55),
    .Y(_02959_));
 sg13g2_a21oi_1 _10633_ (.A1(net382),
    .A2(net54),
    .Y(_00729_),
    .B1(_02959_));
 sg13g2_inv_1 _10634_ (.Y(_02960_),
    .A(\ppu.sprite_buffer.sprite_pixels[1][6] ));
 sg13g2_nor2_1 _10635_ (.A(\ppu.sprite_buffer.sprite_pixels[1][2] ),
    .B(net55),
    .Y(_02961_));
 sg13g2_a21oi_1 _10636_ (.A1(_02960_),
    .A2(net54),
    .Y(_00730_),
    .B1(_02961_));
 sg13g2_nor2_1 _10637_ (.A(\ppu.sprite_buffer.sprite_pixels[1][30] ),
    .B(net55),
    .Y(_02962_));
 sg13g2_a21oi_1 _10638_ (.A1(net336),
    .A2(net54),
    .Y(_00731_),
    .B1(_02962_));
 sg13g2_nor2_1 _10639_ (.A(\ppu.sprite_buffer.sprite_pixels[1][31] ),
    .B(_02953_),
    .Y(_02963_));
 sg13g2_a21oi_1 _10640_ (.A1(_02688_),
    .A2(net54),
    .Y(_00732_),
    .B1(_02963_));
 sg13g2_inv_1 _10641_ (.Y(_02964_),
    .A(\ppu.sprite_buffer.sprite_pixels[1][7] ));
 sg13g2_nor2_1 _10642_ (.A(\ppu.sprite_buffer.sprite_pixels[1][3] ),
    .B(_02953_),
    .Y(_02965_));
 sg13g2_a21oi_1 _10643_ (.A1(_02964_),
    .A2(_02957_),
    .Y(_00733_),
    .B1(_02965_));
 sg13g2_inv_1 _10644_ (.Y(_02966_),
    .A(\ppu.sprite_buffer.sprite_pixels[1][8] ));
 sg13g2_nor2_1 _10645_ (.A(\ppu.sprite_buffer.sprite_pixels[1][4] ),
    .B(_02953_),
    .Y(_02967_));
 sg13g2_a21oi_1 _10646_ (.A1(_02966_),
    .A2(net54),
    .Y(_00734_),
    .B1(_02967_));
 sg13g2_inv_1 _10647_ (.Y(_02968_),
    .A(\ppu.sprite_buffer.sprite_pixels[1][9] ));
 sg13g2_nor2_1 _10648_ (.A(\ppu.sprite_buffer.sprite_pixels[1][5] ),
    .B(_02953_),
    .Y(_02969_));
 sg13g2_a21oi_1 _10649_ (.A1(_02968_),
    .A2(net54),
    .Y(_00735_),
    .B1(_02969_));
 sg13g2_nand2_1 _10650_ (.Y(_02970_),
    .A(net55),
    .B(\ppu.sprite_buffer.sprite_pixels[1][10] ));
 sg13g2_o21ai_1 _10651_ (.B1(_02970_),
    .Y(_00736_),
    .A1(_02960_),
    .A2(net54));
 sg13g2_nand2_1 _10652_ (.Y(_02971_),
    .A(_02956_),
    .B(\ppu.sprite_buffer.sprite_pixels[1][11] ));
 sg13g2_o21ai_1 _10653_ (.B1(_02971_),
    .Y(_00737_),
    .A1(_02964_),
    .A2(_02957_));
 sg13g2_nand2_1 _10654_ (.Y(_02972_),
    .A(net55),
    .B(\ppu.sprite_buffer.sprite_pixels[1][12] ));
 sg13g2_o21ai_1 _10655_ (.B1(_02972_),
    .Y(_00738_),
    .A1(_02966_),
    .A2(net57));
 sg13g2_nand2_1 _10656_ (.Y(_02973_),
    .A(net55),
    .B(\ppu.sprite_buffer.sprite_pixels[1][13] ));
 sg13g2_o21ai_1 _10657_ (.B1(_02973_),
    .Y(_00739_),
    .A1(_02968_),
    .A2(net57));
 sg13g2_nand3_1 _10658_ (.B(_02142_),
    .C(_02146_),
    .A(_02147_),
    .Y(_02974_));
 sg13g2_buf_2 _10659_ (.A(_02974_),
    .X(_02975_));
 sg13g2_buf_1 _10660_ (.A(_02975_),
    .X(_02976_));
 sg13g2_mux2_1 _10661_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][0] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][4] ),
    .S(_02976_),
    .X(_00740_));
 sg13g2_mux2_1 _10662_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][10] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][14] ),
    .S(net53),
    .X(_00741_));
 sg13g2_mux2_1 _10663_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][11] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][15] ),
    .S(net53),
    .X(_00742_));
 sg13g2_mux2_1 _10664_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][12] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][16] ),
    .S(net53),
    .X(_00743_));
 sg13g2_mux2_1 _10665_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][13] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][17] ),
    .S(net53),
    .X(_00744_));
 sg13g2_mux2_1 _10666_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][14] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][18] ),
    .S(net53),
    .X(_00745_));
 sg13g2_mux2_1 _10667_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][15] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][19] ),
    .S(net53),
    .X(_00746_));
 sg13g2_mux2_1 _10668_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][16] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][20] ),
    .S(net53),
    .X(_00747_));
 sg13g2_buf_2 _10669_ (.A(_02975_),
    .X(_02977_));
 sg13g2_mux2_1 _10670_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][17] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][21] ),
    .S(net52),
    .X(_00748_));
 sg13g2_mux2_1 _10671_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][18] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][22] ),
    .S(net52),
    .X(_00749_));
 sg13g2_mux2_1 _10672_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][19] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][23] ),
    .S(_02977_),
    .X(_00750_));
 sg13g2_mux2_1 _10673_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][1] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][5] ),
    .S(net52),
    .X(_00751_));
 sg13g2_mux2_1 _10674_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][20] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][24] ),
    .S(_02977_),
    .X(_00752_));
 sg13g2_mux2_1 _10675_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][21] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][25] ),
    .S(net52),
    .X(_00753_));
 sg13g2_mux2_1 _10676_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][22] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][26] ),
    .S(net52),
    .X(_00754_));
 sg13g2_mux2_1 _10677_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][23] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][27] ),
    .S(net52),
    .X(_00755_));
 sg13g2_mux2_1 _10678_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][24] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][28] ),
    .S(net52),
    .X(_00756_));
 sg13g2_mux2_1 _10679_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][25] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][29] ),
    .S(net52),
    .X(_00757_));
 sg13g2_buf_1 _10680_ (.A(_02975_),
    .X(_02978_));
 sg13g2_mux2_1 _10681_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][26] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][30] ),
    .S(net51),
    .X(_00758_));
 sg13g2_mux2_1 _10682_ (.A0(\ppu.sprite_buffer.sprite_pixels[2][27] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][31] ),
    .S(net51),
    .X(_00759_));
 sg13g2_buf_1 _10683_ (.A(_02975_),
    .X(_02979_));
 sg13g2_nor2_1 _10684_ (.A(\ppu.sprite_buffer.sprite_pixels[2][28] ),
    .B(net51),
    .Y(_02980_));
 sg13g2_a21oi_1 _10685_ (.A1(net381),
    .A2(net50),
    .Y(_00760_),
    .B1(_02980_));
 sg13g2_nor2_1 _10686_ (.A(\ppu.sprite_buffer.sprite_pixels[2][29] ),
    .B(net51),
    .Y(_02981_));
 sg13g2_a21oi_1 _10687_ (.A1(net382),
    .A2(net50),
    .Y(_00761_),
    .B1(_02981_));
 sg13g2_inv_1 _10688_ (.Y(_02982_),
    .A(\ppu.sprite_buffer.sprite_pixels[2][6] ));
 sg13g2_nor2_1 _10689_ (.A(\ppu.sprite_buffer.sprite_pixels[2][2] ),
    .B(_02978_),
    .Y(_02983_));
 sg13g2_a21oi_1 _10690_ (.A1(_02982_),
    .A2(net50),
    .Y(_00762_),
    .B1(_02983_));
 sg13g2_nor2_1 _10691_ (.A(\ppu.sprite_buffer.sprite_pixels[2][30] ),
    .B(net51),
    .Y(_02984_));
 sg13g2_a21oi_1 _10692_ (.A1(net336),
    .A2(net50),
    .Y(_00763_),
    .B1(_02984_));
 sg13g2_nor2_1 _10693_ (.A(\ppu.sprite_buffer.sprite_pixels[2][31] ),
    .B(_02975_),
    .Y(_02985_));
 sg13g2_a21oi_1 _10694_ (.A1(net335),
    .A2(net50),
    .Y(_00764_),
    .B1(_02985_));
 sg13g2_inv_1 _10695_ (.Y(_02986_),
    .A(\ppu.sprite_buffer.sprite_pixels[2][7] ));
 sg13g2_nor2_1 _10696_ (.A(\ppu.sprite_buffer.sprite_pixels[2][3] ),
    .B(_02975_),
    .Y(_02987_));
 sg13g2_a21oi_1 _10697_ (.A1(_02986_),
    .A2(net50),
    .Y(_00765_),
    .B1(_02987_));
 sg13g2_inv_1 _10698_ (.Y(_02988_),
    .A(\ppu.sprite_buffer.sprite_pixels[2][8] ));
 sg13g2_nor2_1 _10699_ (.A(\ppu.sprite_buffer.sprite_pixels[2][4] ),
    .B(_02975_),
    .Y(_02989_));
 sg13g2_a21oi_1 _10700_ (.A1(_02988_),
    .A2(net50),
    .Y(_00766_),
    .B1(_02989_));
 sg13g2_inv_1 _10701_ (.Y(_02990_),
    .A(\ppu.sprite_buffer.sprite_pixels[2][9] ));
 sg13g2_nor2_1 _10702_ (.A(\ppu.sprite_buffer.sprite_pixels[2][5] ),
    .B(_02975_),
    .Y(_02991_));
 sg13g2_a21oi_1 _10703_ (.A1(_02990_),
    .A2(net50),
    .Y(_00767_),
    .B1(_02991_));
 sg13g2_nand2_1 _10704_ (.Y(_02992_),
    .A(net51),
    .B(\ppu.sprite_buffer.sprite_pixels[2][10] ));
 sg13g2_o21ai_1 _10705_ (.B1(_02992_),
    .Y(_00768_),
    .A1(_02982_),
    .A2(_02979_));
 sg13g2_nand2_1 _10706_ (.Y(_02993_),
    .A(net51),
    .B(\ppu.sprite_buffer.sprite_pixels[2][11] ));
 sg13g2_o21ai_1 _10707_ (.B1(_02993_),
    .Y(_00769_),
    .A1(_02986_),
    .A2(_02979_));
 sg13g2_nand2_1 _10708_ (.Y(_02994_),
    .A(net51),
    .B(\ppu.sprite_buffer.sprite_pixels[2][12] ));
 sg13g2_o21ai_1 _10709_ (.B1(_02994_),
    .Y(_00770_),
    .A1(_02988_),
    .A2(_02976_));
 sg13g2_nand2_1 _10710_ (.Y(_02995_),
    .A(_02978_),
    .B(\ppu.sprite_buffer.sprite_pixels[2][13] ));
 sg13g2_o21ai_1 _10711_ (.B1(_02995_),
    .Y(_00771_),
    .A1(_02990_),
    .A2(net53));
 sg13g2_nand3_1 _10712_ (.B(_01910_),
    .C(_02115_),
    .A(_02114_),
    .Y(_02996_));
 sg13g2_buf_2 _10713_ (.A(_02996_),
    .X(_02997_));
 sg13g2_buf_1 _10714_ (.A(_02997_),
    .X(_02998_));
 sg13g2_mux2_1 _10715_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][0] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][4] ),
    .S(net49),
    .X(_00772_));
 sg13g2_mux2_1 _10716_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][10] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][14] ),
    .S(net49),
    .X(_00773_));
 sg13g2_mux2_1 _10717_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][11] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][15] ),
    .S(_02998_),
    .X(_00774_));
 sg13g2_mux2_1 _10718_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][12] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][16] ),
    .S(net49),
    .X(_00775_));
 sg13g2_mux2_1 _10719_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][13] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][17] ),
    .S(net49),
    .X(_00776_));
 sg13g2_mux2_1 _10720_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][14] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][18] ),
    .S(net49),
    .X(_00777_));
 sg13g2_mux2_1 _10721_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][15] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][19] ),
    .S(net49),
    .X(_00778_));
 sg13g2_mux2_1 _10722_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][16] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][20] ),
    .S(net49),
    .X(_00779_));
 sg13g2_buf_2 _10723_ (.A(_02997_),
    .X(_02999_));
 sg13g2_mux2_1 _10724_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][17] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][21] ),
    .S(net48),
    .X(_00780_));
 sg13g2_mux2_1 _10725_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][18] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][22] ),
    .S(net48),
    .X(_00781_));
 sg13g2_mux2_1 _10726_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][19] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][23] ),
    .S(_02999_),
    .X(_00782_));
 sg13g2_mux2_1 _10727_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][1] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][5] ),
    .S(net48),
    .X(_00783_));
 sg13g2_mux2_1 _10728_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][20] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][24] ),
    .S(net48),
    .X(_00784_));
 sg13g2_mux2_1 _10729_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][21] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][25] ),
    .S(net48),
    .X(_00785_));
 sg13g2_mux2_1 _10730_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][22] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][26] ),
    .S(net48),
    .X(_00786_));
 sg13g2_mux2_1 _10731_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][23] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][27] ),
    .S(_02999_),
    .X(_00787_));
 sg13g2_mux2_1 _10732_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][24] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][28] ),
    .S(net48),
    .X(_00788_));
 sg13g2_mux2_1 _10733_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][25] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][29] ),
    .S(net48),
    .X(_00789_));
 sg13g2_buf_1 _10734_ (.A(_02997_),
    .X(_03000_));
 sg13g2_mux2_1 _10735_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][26] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][30] ),
    .S(net47),
    .X(_00790_));
 sg13g2_mux2_1 _10736_ (.A0(\ppu.sprite_buffer.sprite_pixels[3][27] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[3][31] ),
    .S(net47),
    .X(_00791_));
 sg13g2_buf_1 _10737_ (.A(_02997_),
    .X(_03001_));
 sg13g2_nor2_1 _10738_ (.A(\ppu.sprite_buffer.sprite_pixels[3][28] ),
    .B(net47),
    .Y(_03002_));
 sg13g2_a21oi_1 _10739_ (.A1(_02721_),
    .A2(net46),
    .Y(_00792_),
    .B1(_03002_));
 sg13g2_nor2_1 _10740_ (.A(\ppu.sprite_buffer.sprite_pixels[3][29] ),
    .B(net47),
    .Y(_03003_));
 sg13g2_a21oi_1 _10741_ (.A1(_02505_),
    .A2(net46),
    .Y(_00793_),
    .B1(_03003_));
 sg13g2_inv_1 _10742_ (.Y(_03004_),
    .A(\ppu.sprite_buffer.sprite_pixels[3][6] ));
 sg13g2_nor2_1 _10743_ (.A(\ppu.sprite_buffer.sprite_pixels[3][2] ),
    .B(_03000_),
    .Y(_03005_));
 sg13g2_a21oi_1 _10744_ (.A1(_03004_),
    .A2(net46),
    .Y(_00794_),
    .B1(_03005_));
 sg13g2_nor2_1 _10745_ (.A(\ppu.sprite_buffer.sprite_pixels[3][30] ),
    .B(net47),
    .Y(_03006_));
 sg13g2_a21oi_1 _10746_ (.A1(net336),
    .A2(net46),
    .Y(_00795_),
    .B1(_03006_));
 sg13g2_nor2_1 _10747_ (.A(\ppu.sprite_buffer.sprite_pixels[3][31] ),
    .B(_02997_),
    .Y(_03007_));
 sg13g2_a21oi_1 _10748_ (.A1(net335),
    .A2(_03001_),
    .Y(_00796_),
    .B1(_03007_));
 sg13g2_inv_1 _10749_ (.Y(_03008_),
    .A(\ppu.sprite_buffer.sprite_pixels[3][7] ));
 sg13g2_nor2_1 _10750_ (.A(\ppu.sprite_buffer.sprite_pixels[3][3] ),
    .B(_02997_),
    .Y(_03009_));
 sg13g2_a21oi_1 _10751_ (.A1(_03008_),
    .A2(_03001_),
    .Y(_00797_),
    .B1(_03009_));
 sg13g2_inv_1 _10752_ (.Y(_03010_),
    .A(\ppu.sprite_buffer.sprite_pixels[3][8] ));
 sg13g2_nor2_1 _10753_ (.A(\ppu.sprite_buffer.sprite_pixels[3][4] ),
    .B(_02997_),
    .Y(_03011_));
 sg13g2_a21oi_1 _10754_ (.A1(_03010_),
    .A2(net46),
    .Y(_00798_),
    .B1(_03011_));
 sg13g2_inv_1 _10755_ (.Y(_03012_),
    .A(\ppu.sprite_buffer.sprite_pixels[3][9] ));
 sg13g2_nor2_1 _10756_ (.A(\ppu.sprite_buffer.sprite_pixels[3][5] ),
    .B(_02997_),
    .Y(_03013_));
 sg13g2_a21oi_1 _10757_ (.A1(_03012_),
    .A2(net46),
    .Y(_00799_),
    .B1(_03013_));
 sg13g2_nand2_1 _10758_ (.Y(_03014_),
    .A(net47),
    .B(\ppu.sprite_buffer.sprite_pixels[3][10] ));
 sg13g2_o21ai_1 _10759_ (.B1(_03014_),
    .Y(_00800_),
    .A1(_03004_),
    .A2(net46));
 sg13g2_nand2_1 _10760_ (.Y(_03015_),
    .A(net47),
    .B(\ppu.sprite_buffer.sprite_pixels[3][11] ));
 sg13g2_o21ai_1 _10761_ (.B1(_03015_),
    .Y(_00801_),
    .A1(_03008_),
    .A2(net46));
 sg13g2_nand2_1 _10762_ (.Y(_03016_),
    .A(_03000_),
    .B(\ppu.sprite_buffer.sprite_pixels[3][12] ));
 sg13g2_o21ai_1 _10763_ (.B1(_03016_),
    .Y(_00802_),
    .A1(_03010_),
    .A2(net49));
 sg13g2_nand2_1 _10764_ (.Y(_03017_),
    .A(net47),
    .B(\ppu.sprite_buffer.sprite_pixels[3][13] ));
 sg13g2_o21ai_1 _10765_ (.B1(_03017_),
    .Y(_00803_),
    .A1(_03012_),
    .A2(_02998_));
 sg13g2_inv_1 _10766_ (.Y(_03018_),
    .A(\ppu.sprite_buffer.top_prio[2] ));
 sg13g2_nand2_1 _10767_ (.Y(_03019_),
    .A(net261),
    .B(\ppu.sprite_buffer.attr_x[1][11] ));
 sg13g2_o21ai_1 _10768_ (.B1(_01855_),
    .Y(_03020_),
    .A1(_01933_),
    .A2(_02739_));
 sg13g2_o21ai_1 _10769_ (.B1(_03020_),
    .Y(_03021_),
    .A1(\ppu.sprite_buffer.attr_x[2][11] ),
    .A2(_02028_));
 sg13g2_a22oi_1 _10770_ (.Y(_03022_),
    .B1(_03019_),
    .B2(_03021_),
    .A2(net253),
    .A1(_00123_));
 sg13g2_nand2_1 _10771_ (.Y(_03023_),
    .A(net261),
    .B(\ppu.sprite_buffer.sprite_pixels[1][3] ));
 sg13g2_a21o_1 _10772_ (.A2(\ppu.sprite_buffer.sprite_pixels[3][3] ),
    .A1(_01854_),
    .B1(_01918_),
    .X(_03024_));
 sg13g2_o21ai_1 _10773_ (.B1(_03024_),
    .Y(_03025_),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][3] ),
    .A2(_02028_));
 sg13g2_a22oi_1 _10774_ (.Y(_03026_),
    .B1(_03023_),
    .B2(_03025_),
    .A2(net260),
    .A1(_00125_));
 sg13g2_inv_1 _10775_ (.Y(_03027_),
    .A(_03026_));
 sg13g2_nand2_1 _10776_ (.Y(_03028_),
    .A(net261),
    .B(\ppu.sprite_buffer.sprite_pixels[1][1] ));
 sg13g2_a21o_1 _10777_ (.A2(\ppu.sprite_buffer.sprite_pixels[3][1] ),
    .A1(_01854_),
    .B1(_02053_),
    .X(_03029_));
 sg13g2_o21ai_1 _10778_ (.B1(_03029_),
    .Y(_03030_),
    .A1(\ppu.sprite_buffer.sprite_pixels[2][1] ),
    .A2(_02028_));
 sg13g2_a22oi_1 _10779_ (.Y(_03031_),
    .B1(_03028_),
    .B2(_03030_),
    .A2(net253),
    .A1(_00124_));
 sg13g2_nor2_1 _10780_ (.A(_03031_),
    .B(_02098_),
    .Y(_03032_));
 sg13g2_a21oi_1 _10781_ (.A1(_02098_),
    .A2(_03027_),
    .Y(_03033_),
    .B1(_03032_));
 sg13g2_inv_1 _10782_ (.Y(_03034_),
    .A(_03033_));
 sg13g2_inv_1 _10783_ (.Y(_03035_),
    .A(\ppu.sprite_buffer.sprite_pixels[3][2] ));
 sg13g2_nand2_1 _10784_ (.Y(_03036_),
    .A(_01923_),
    .B(\ppu.sprite_buffer.sprite_pixels[2][2] ));
 sg13g2_o21ai_1 _10785_ (.B1(_03036_),
    .Y(_03037_),
    .A1(_03035_),
    .A2(net345));
 sg13g2_a221oi_1 _10786_ (.B2(net253),
    .C1(_03037_),
    .B1(\ppu.sprite_buffer.sprite_pixels[0][2] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][2] ),
    .Y(_03038_),
    .A2(net261));
 sg13g2_inv_1 _10787_ (.Y(_03039_),
    .A(_03038_));
 sg13g2_inv_1 _10788_ (.Y(_03040_),
    .A(\ppu.sprite_buffer.sprite_pixels[3][0] ));
 sg13g2_nand2_1 _10789_ (.Y(_03041_),
    .A(_01923_),
    .B(\ppu.sprite_buffer.sprite_pixels[2][0] ));
 sg13g2_o21ai_1 _10790_ (.B1(_03041_),
    .Y(_03042_),
    .A1(_03040_),
    .A2(net345));
 sg13g2_a221oi_1 _10791_ (.B2(net260),
    .C1(_03042_),
    .B1(\ppu.sprite_buffer.sprite_pixels[0][0] ),
    .A1(\ppu.sprite_buffer.sprite_pixels[1][0] ),
    .Y(_03043_),
    .A2(net261));
 sg13g2_nor2_1 _10792_ (.A(_03043_),
    .B(_02098_),
    .Y(_03044_));
 sg13g2_a21oi_1 _10793_ (.A1(_02098_),
    .A2(_03039_),
    .Y(_03045_),
    .B1(_03044_));
 sg13g2_nand3b_1 _10794_ (.B(_03034_),
    .C(_03045_),
    .Y(_03046_),
    .A_N(_03022_));
 sg13g2_buf_1 _10795_ (.A(_03046_),
    .X(_03047_));
 sg13g2_nor2_1 _10796_ (.A(_03031_),
    .B(_02057_),
    .Y(_03048_));
 sg13g2_nor2_1 _10797_ (.A(_03022_),
    .B(_03026_),
    .Y(_03049_));
 sg13g2_nand4_1 _10798_ (.B(_03043_),
    .C(_03038_),
    .A(_03048_),
    .Y(_03050_),
    .D(_03049_));
 sg13g2_o21ai_1 _10799_ (.B1(_03050_),
    .Y(_03051_),
    .A1(_02059_),
    .A2(_03047_));
 sg13g2_inv_1 _10800_ (.Y(_03052_),
    .A(_03051_));
 sg13g2_nor2_1 _10801_ (.A(_02028_),
    .B(_02146_),
    .Y(_03053_));
 sg13g2_a221oi_1 _10802_ (.B2(_02185_),
    .C1(_03053_),
    .B1(_02051_),
    .A1(_02165_),
    .Y(_03054_),
    .A2(net252));
 sg13g2_nand2_1 _10803_ (.Y(_03055_),
    .A(_03052_),
    .B(_03054_));
 sg13g2_a21oi_1 _10804_ (.A1(_01904_),
    .A2(_02116_),
    .Y(_03056_),
    .B1(_03055_));
 sg13g2_nor2b_1 _10805_ (.A(_02112_),
    .B_N(_03056_),
    .Y(_03057_));
 sg13g2_buf_2 _10806_ (.A(_03057_),
    .X(_03058_));
 sg13g2_buf_8 _10807_ (.A(_03058_),
    .X(_03059_));
 sg13g2_inv_1 _10808_ (.Y(_03060_),
    .A(\ppu.sprite_buffer.sprite_ids[3][2] ));
 sg13g2_nand2_1 _10809_ (.Y(_03061_),
    .A(net259),
    .B(\ppu.sprite_buffer.sprite_ids[2][2] ));
 sg13g2_o21ai_1 _10810_ (.B1(_03061_),
    .Y(_03062_),
    .A1(_03060_),
    .A2(net345));
 sg13g2_a221oi_1 _10811_ (.B2(net237),
    .C1(_03062_),
    .B1(\ppu.sprite_buffer.sprite_ids[0][2] ),
    .A1(\ppu.sprite_buffer.sprite_ids[1][2] ),
    .Y(_03063_),
    .A2(net252));
 sg13g2_nand2_1 _10812_ (.Y(_03064_),
    .A(net72),
    .B(_03063_));
 sg13g2_nor2_1 _10813_ (.A(_03018_),
    .B(_03064_),
    .Y(_03065_));
 sg13g2_inv_1 _10814_ (.Y(_03066_),
    .A(\ppu.sprite_buffer.top_prio[1] ));
 sg13g2_inv_1 _10815_ (.Y(_03067_),
    .A(\ppu.sprite_buffer.sprite_ids[3][1] ));
 sg13g2_nand2_1 _10816_ (.Y(_03068_),
    .A(net259),
    .B(\ppu.sprite_buffer.sprite_ids[2][1] ));
 sg13g2_o21ai_1 _10817_ (.B1(_03068_),
    .Y(_03069_),
    .A1(_03067_),
    .A2(net345));
 sg13g2_a221oi_1 _10818_ (.B2(net237),
    .C1(_03069_),
    .B1(\ppu.sprite_buffer.sprite_ids[0][1] ),
    .A1(\ppu.sprite_buffer.sprite_ids[1][1] ),
    .Y(_03070_),
    .A2(net252));
 sg13g2_nand2_1 _10819_ (.Y(_03071_),
    .A(net72),
    .B(_03070_));
 sg13g2_nor2_1 _10820_ (.A(_03066_),
    .B(_03071_),
    .Y(_03072_));
 sg13g2_nor2_1 _10821_ (.A(_03065_),
    .B(_03072_),
    .Y(_03073_));
 sg13g2_inv_1 _10822_ (.Y(_03074_),
    .A(\ppu.sprite_buffer.sprite_ids[3][0] ));
 sg13g2_nand2_1 _10823_ (.Y(_03075_),
    .A(net259),
    .B(\ppu.sprite_buffer.sprite_ids[2][0] ));
 sg13g2_o21ai_1 _10824_ (.B1(_03075_),
    .Y(_03076_),
    .A1(_03074_),
    .A2(net297));
 sg13g2_a221oi_1 _10825_ (.B2(_02182_),
    .C1(_03076_),
    .B1(\ppu.sprite_buffer.sprite_ids[0][0] ),
    .A1(\ppu.sprite_buffer.sprite_ids[1][0] ),
    .Y(_03077_),
    .A2(net252));
 sg13g2_nand2_1 _10826_ (.Y(_03078_),
    .A(net72),
    .B(_03077_));
 sg13g2_nand2b_1 _10827_ (.Y(_03079_),
    .B(_03078_),
    .A_N(\ppu.sprite_buffer.top_prio[0] ));
 sg13g2_nand2_1 _10828_ (.Y(_03080_),
    .A(_03071_),
    .B(_03066_));
 sg13g2_nand2_1 _10829_ (.Y(_03081_),
    .A(_03079_),
    .B(_03080_));
 sg13g2_nand2_1 _10830_ (.Y(_03082_),
    .A(_03073_),
    .B(_03081_));
 sg13g2_nand2_1 _10831_ (.Y(_03083_),
    .A(_03064_),
    .B(_03018_));
 sg13g2_a22oi_1 _10832_ (.Y(_03084_),
    .B1(\ppu.sprite_buffer.sprite_ids[3][3] ),
    .B2(net263),
    .A2(\ppu.sprite_buffer.sprite_ids[1][3] ),
    .A1(net252));
 sg13g2_buf_1 _10833_ (.A(net344),
    .X(_03085_));
 sg13g2_o21ai_1 _10834_ (.B1(net343),
    .Y(_03086_),
    .A1(\ppu.sprite_buffer.sprite_ids[2][3] ),
    .A2(net294));
 sg13g2_nand2_1 _10835_ (.Y(_03087_),
    .A(_03084_),
    .B(_03086_));
 sg13g2_o21ai_1 _10836_ (.B1(_03087_),
    .Y(_03088_),
    .A1(\ppu.sprite_buffer.sprite_ids[0][3] ),
    .A2(net262));
 sg13g2_nand3_1 _10837_ (.B(\ppu.sprite_buffer.top_prio[3] ),
    .C(_03088_),
    .A(net72),
    .Y(_03089_));
 sg13g2_nand2_1 _10838_ (.Y(_03090_),
    .A(_03083_),
    .B(_03089_));
 sg13g2_nand2_1 _10839_ (.Y(_03091_),
    .A(net72),
    .B(_03088_));
 sg13g2_nand2b_1 _10840_ (.Y(_03092_),
    .B(_03091_),
    .A_N(\ppu.sprite_buffer.top_prio[3] ));
 sg13g2_inv_1 _10841_ (.Y(_03093_),
    .A(\ppu.sprite_buffer.sprite_ids[3][4] ));
 sg13g2_nand2_1 _10842_ (.Y(_03094_),
    .A(_02109_),
    .B(\ppu.sprite_buffer.sprite_ids[2][4] ));
 sg13g2_o21ai_1 _10843_ (.B1(_03094_),
    .Y(_03095_),
    .A1(_03093_),
    .A2(_01857_));
 sg13g2_a221oi_1 _10844_ (.B2(_02182_),
    .C1(_03095_),
    .B1(\ppu.sprite_buffer.sprite_ids[0][4] ),
    .A1(\ppu.sprite_buffer.sprite_ids[1][4] ),
    .Y(_03096_),
    .A2(_02108_));
 sg13g2_nand2_1 _10845_ (.Y(_03097_),
    .A(net72),
    .B(_03096_));
 sg13g2_nand2b_1 _10846_ (.Y(_03098_),
    .B(_03097_),
    .A_N(\ppu.sprite_buffer.top_prio[4] ));
 sg13g2_nand2_1 _10847_ (.Y(_03099_),
    .A(_03092_),
    .B(_03098_));
 sg13g2_nor2_1 _10848_ (.A(_03090_),
    .B(_03099_),
    .Y(_03100_));
 sg13g2_nand3_1 _10849_ (.B(\ppu.sprite_buffer.top_prio[4] ),
    .C(_03096_),
    .A(_03059_),
    .Y(_03101_));
 sg13g2_inv_1 _10850_ (.Y(_03102_),
    .A(\ppu.sprite_buffer.sprite_ids[3][5] ));
 sg13g2_nand2_1 _10851_ (.Y(_03103_),
    .A(_02109_),
    .B(\ppu.sprite_buffer.sprite_ids[2][5] ));
 sg13g2_o21ai_1 _10852_ (.B1(_03103_),
    .Y(_03104_),
    .A1(_03102_),
    .A2(_01857_));
 sg13g2_a221oi_1 _10853_ (.B2(net253),
    .C1(_03104_),
    .B1(\ppu.sprite_buffer.sprite_ids[0][5] ),
    .A1(\ppu.sprite_buffer.sprite_ids[1][5] ),
    .Y(_03105_),
    .A2(_02108_));
 sg13g2_inv_1 _10854_ (.Y(_03106_),
    .A(_00126_));
 sg13g2_a21oi_1 _10855_ (.A1(_03105_),
    .A2(\ppu.sprite_buffer.top_prio[5] ),
    .Y(_03107_),
    .B1(_03106_));
 sg13g2_nand2b_1 _10856_ (.Y(_03108_),
    .B(_03059_),
    .A_N(_03107_));
 sg13g2_nand2_1 _10857_ (.Y(_03109_),
    .A(_03101_),
    .B(_03108_));
 sg13g2_nand2_1 _10858_ (.Y(_03110_),
    .A(_03058_),
    .B(_03105_));
 sg13g2_nand2b_1 _10859_ (.Y(_03111_),
    .B(_03110_),
    .A_N(\ppu.sprite_buffer.top_prio[5] ));
 sg13g2_inv_1 _10860_ (.Y(_03112_),
    .A(_03058_));
 sg13g2_nand2_1 _10861_ (.Y(_03113_),
    .A(_03112_),
    .B(_00126_));
 sg13g2_nand2_1 _10862_ (.Y(_03114_),
    .A(_03111_),
    .B(_03113_));
 sg13g2_nor2_1 _10863_ (.A(_03109_),
    .B(_03114_),
    .Y(_03115_));
 sg13g2_nand3_1 _10864_ (.B(_03100_),
    .C(_03115_),
    .A(_03082_),
    .Y(_03116_));
 sg13g2_nor2b_1 _10865_ (.A(_03114_),
    .B_N(_03098_),
    .Y(_03117_));
 sg13g2_nand2_1 _10866_ (.Y(_03118_),
    .A(_03089_),
    .B(_03101_));
 sg13g2_inv_1 _10867_ (.Y(_03119_),
    .A(_03108_));
 sg13g2_a21oi_1 _10868_ (.A1(_03117_),
    .A2(_03118_),
    .Y(_03120_),
    .B1(_03119_));
 sg13g2_nand2_1 _10869_ (.Y(_03121_),
    .A(_03116_),
    .B(_03120_));
 sg13g2_nand2_1 _10870_ (.Y(_03122_),
    .A(_03121_),
    .B(_03052_));
 sg13g2_buf_1 _10871_ (.A(_03122_),
    .X(_03123_));
 sg13g2_nand2_2 _10872_ (.Y(_03124_),
    .A(_03123_),
    .B(net262));
 sg13g2_buf_8 _10873_ (.A(_03124_),
    .X(_03125_));
 sg13g2_inv_1 _10874_ (.Y(_03126_),
    .A(_02050_));
 sg13g2_nor2_1 _10875_ (.A(_02033_),
    .B(_03034_),
    .Y(_03127_));
 sg13g2_inv_1 _10876_ (.Y(_03128_),
    .A(_03127_));
 sg13g2_nor2_1 _10877_ (.A(_02039_),
    .B(_03128_),
    .Y(_03129_));
 sg13g2_o21ai_1 _10878_ (.B1(_03047_),
    .Y(_03130_),
    .A1(_02038_),
    .A2(_03127_));
 sg13g2_nor2_1 _10879_ (.A(_03129_),
    .B(_03130_),
    .Y(_03131_));
 sg13g2_nor2_1 _10880_ (.A(_03126_),
    .B(_03131_),
    .Y(_03132_));
 sg13g2_a21oi_1 _10881_ (.A1(_03126_),
    .A2(_03045_),
    .Y(_03133_),
    .B1(_03132_));
 sg13g2_nor2_1 _10882_ (.A(_03043_),
    .B(net145),
    .Y(_03134_));
 sg13g2_a21oi_1 _10883_ (.A1(_03133_),
    .A2(net145),
    .Y(_03135_),
    .B1(_03134_));
 sg13g2_nor2_1 _10884_ (.A(_03135_),
    .B(_03112_),
    .Y(_03136_));
 sg13g2_nand2_1 _10885_ (.Y(_03137_),
    .A(net28),
    .B(_03136_));
 sg13g2_buf_1 _10886_ (.A(_03123_),
    .X(_03138_));
 sg13g2_nand3_1 _10887_ (.B(\ppu.sprite_buffer.top_color[0] ),
    .C(net246),
    .A(net31),
    .Y(_03139_));
 sg13g2_nand2_1 _10888_ (.Y(_00804_),
    .A(_03137_),
    .B(_03139_));
 sg13g2_xor2_1 _10889_ (.B(_03129_),
    .A(_02055_),
    .X(_03140_));
 sg13g2_nand2_1 _10890_ (.Y(_03141_),
    .A(_03140_),
    .B(_03047_));
 sg13g2_inv_1 _10891_ (.Y(_03142_),
    .A(_03141_));
 sg13g2_nand2_1 _10892_ (.Y(_03143_),
    .A(_03034_),
    .B(_02033_));
 sg13g2_nand3_1 _10893_ (.B(_03128_),
    .C(_03143_),
    .A(_03047_),
    .Y(_03144_));
 sg13g2_o21ai_1 _10894_ (.B1(net145),
    .Y(_03145_),
    .A1(_02050_),
    .A2(_03144_));
 sg13g2_a21oi_1 _10895_ (.A1(_03142_),
    .A2(_02050_),
    .Y(_03146_),
    .B1(_03145_));
 sg13g2_nor3_1 _10896_ (.A(_03048_),
    .B(_03146_),
    .C(_03112_),
    .Y(_03147_));
 sg13g2_nand2_1 _10897_ (.Y(_03148_),
    .A(net28),
    .B(_03147_));
 sg13g2_nand3_1 _10898_ (.B(\ppu.sprite_buffer.top_color[1] ),
    .C(_02927_),
    .A(net31),
    .Y(_03149_));
 sg13g2_nand2_1 _10899_ (.Y(_00805_),
    .A(_03148_),
    .B(_03149_));
 sg13g2_o21ai_1 _10900_ (.B1(net145),
    .Y(_03150_),
    .A1(_03126_),
    .A2(_03045_));
 sg13g2_a21oi_1 _10901_ (.A1(_03131_),
    .A2(_03126_),
    .Y(_03151_),
    .B1(_03150_));
 sg13g2_nor2_1 _10902_ (.A(_03039_),
    .B(_02058_),
    .Y(_03152_));
 sg13g2_nor3_1 _10903_ (.A(_03151_),
    .B(_03152_),
    .C(_03112_),
    .Y(_03153_));
 sg13g2_nand2_1 _10904_ (.Y(_03154_),
    .A(net28),
    .B(_03153_));
 sg13g2_nand3_1 _10905_ (.B(\ppu.sprite_buffer.top_color[2] ),
    .C(_02927_),
    .A(net31),
    .Y(_03155_));
 sg13g2_nand2_1 _10906_ (.Y(_00806_),
    .A(_03154_),
    .B(_03155_));
 sg13g2_a21oi_1 _10907_ (.A1(_03144_),
    .A2(_02050_),
    .Y(_03156_),
    .B1(_02059_));
 sg13g2_nand2_1 _10908_ (.Y(_03157_),
    .A(_03141_),
    .B(_03126_));
 sg13g2_a22oi_1 _10909_ (.Y(_03158_),
    .B1(_03156_),
    .B2(_03157_),
    .A2(_03026_),
    .A1(_02059_));
 sg13g2_nor2_1 _10910_ (.A(_03158_),
    .B(_03112_),
    .Y(_03159_));
 sg13g2_nand2_1 _10911_ (.Y(_03160_),
    .A(net28),
    .B(_03159_));
 sg13g2_buf_1 _10912_ (.A(_01921_),
    .X(_03161_));
 sg13g2_nand3_1 _10913_ (.B(\ppu.sprite_buffer.top_color[3] ),
    .C(net245),
    .A(_03138_),
    .Y(_03162_));
 sg13g2_nand2_1 _10914_ (.Y(_00807_),
    .A(_03160_),
    .B(_03162_));
 sg13g2_nand2_1 _10915_ (.Y(_03163_),
    .A(_02501_),
    .B(\ppu.sprite_buffer.attr_x[1][9] ));
 sg13g2_a22oi_1 _10916_ (.Y(_03164_),
    .B1(\ppu.sprite_buffer.attr_x[3][9] ),
    .B2(net236),
    .A2(\ppu.sprite_buffer.attr_x[2][9] ),
    .A1(net251));
 sg13g2_nand2_1 _10917_ (.Y(_03165_),
    .A(net216),
    .B(\ppu.sprite_buffer.attr_x[0][9] ));
 sg13g2_nand4_1 _10918_ (.B(_03163_),
    .C(_03164_),
    .A(net72),
    .Y(_03166_),
    .D(_03165_));
 sg13g2_nand2_1 _10919_ (.Y(_03167_),
    .A(net28),
    .B(_03166_));
 sg13g2_nand3_1 _10920_ (.B(\ppu.sprite_buffer.top_depth[0] ),
    .C(net245),
    .A(net31),
    .Y(_03168_));
 sg13g2_nand2_1 _10921_ (.Y(_00808_),
    .A(_03167_),
    .B(_03168_));
 sg13g2_nand2_1 _10922_ (.Y(_03169_),
    .A(net235),
    .B(\ppu.sprite_buffer.attr_x[1][10] ));
 sg13g2_a22oi_1 _10923_ (.Y(_03170_),
    .B1(\ppu.sprite_buffer.attr_x[3][10] ),
    .B2(net236),
    .A2(\ppu.sprite_buffer.attr_x[2][10] ),
    .A1(net251));
 sg13g2_nand2_1 _10924_ (.Y(_03171_),
    .A(net216),
    .B(\ppu.sprite_buffer.attr_x[0][10] ));
 sg13g2_nand4_1 _10925_ (.B(_03169_),
    .C(_03170_),
    .A(net72),
    .Y(_03172_),
    .D(_03171_));
 sg13g2_nand2_1 _10926_ (.Y(_03173_),
    .A(net28),
    .B(_03172_));
 sg13g2_nand3_1 _10927_ (.B(\ppu.sprite_buffer.top_depth[1] ),
    .C(net245),
    .A(net31),
    .Y(_03174_));
 sg13g2_nand2_1 _10928_ (.Y(_00809_),
    .A(_03173_),
    .B(_03174_));
 sg13g2_nand2_1 _10929_ (.Y(_03175_),
    .A(net28),
    .B(_03078_));
 sg13g2_nand3_1 _10930_ (.B(\ppu.sprite_buffer.top_prio[0] ),
    .C(net245),
    .A(net31),
    .Y(_03176_));
 sg13g2_nand2_1 _10931_ (.Y(_00810_),
    .A(_03175_),
    .B(_03176_));
 sg13g2_nand2_1 _10932_ (.Y(_03177_),
    .A(net28),
    .B(_03071_));
 sg13g2_nand3_1 _10933_ (.B(\ppu.sprite_buffer.top_prio[1] ),
    .C(net245),
    .A(net31),
    .Y(_03178_));
 sg13g2_nand2_1 _10934_ (.Y(_00811_),
    .A(_03177_),
    .B(_03178_));
 sg13g2_nand2_1 _10935_ (.Y(_03179_),
    .A(_03125_),
    .B(_03064_));
 sg13g2_nand3_1 _10936_ (.B(\ppu.sprite_buffer.top_prio[2] ),
    .C(net245),
    .A(net31),
    .Y(_03180_));
 sg13g2_nand2_1 _10937_ (.Y(_00812_),
    .A(_03179_),
    .B(_03180_));
 sg13g2_nand2_1 _10938_ (.Y(_03181_),
    .A(_03125_),
    .B(_03091_));
 sg13g2_nand3_1 _10939_ (.B(\ppu.sprite_buffer.top_prio[3] ),
    .C(net245),
    .A(_03138_),
    .Y(_03182_));
 sg13g2_nand2_1 _10940_ (.Y(_00813_),
    .A(_03181_),
    .B(_03182_));
 sg13g2_nand2_1 _10941_ (.Y(_03183_),
    .A(_03124_),
    .B(_03097_));
 sg13g2_nand3_1 _10942_ (.B(\ppu.sprite_buffer.top_prio[4] ),
    .C(net245),
    .A(_03123_),
    .Y(_03184_));
 sg13g2_nand2_1 _10943_ (.Y(_00814_),
    .A(_03183_),
    .B(_03184_));
 sg13g2_nand2_1 _10944_ (.Y(_03185_),
    .A(_03124_),
    .B(_03110_));
 sg13g2_nand3_1 _10945_ (.B(\ppu.sprite_buffer.top_prio[5] ),
    .C(_03161_),
    .A(_03123_),
    .Y(_03186_));
 sg13g2_nand2_1 _10946_ (.Y(_00815_),
    .A(_03185_),
    .B(_03186_));
 sg13g2_nand2_1 _10947_ (.Y(_03187_),
    .A(_03124_),
    .B(_03112_));
 sg13g2_nand3_1 _10948_ (.B(\ppu.sprite_buffer.top_prio[6] ),
    .C(_03161_),
    .A(_03123_),
    .Y(_03188_));
 sg13g2_nand2_1 _10949_ (.Y(_00816_),
    .A(_03187_),
    .B(_03188_));
 sg13g2_xnor2_1 _10950_ (.Y(_03189_),
    .A(net392),
    .B(\ppu.scroll_regs[0][0] ));
 sg13g2_nor3_1 _10951_ (.A(_01860_),
    .B(_00031_),
    .C(_01901_),
    .Y(_03190_));
 sg13g2_inv_1 _10952_ (.Y(_03191_),
    .A(_03190_));
 sg13g2_nor2_1 _10953_ (.A(_02095_),
    .B(_03191_),
    .Y(_03192_));
 sg13g2_buf_1 _10954_ (.A(_03192_),
    .X(_03193_));
 sg13g2_o21ai_1 _10955_ (.B1(net244),
    .Y(_03194_),
    .A1(net254),
    .A2(_03189_));
 sg13g2_buf_1 _10956_ (.A(_03194_),
    .X(_03195_));
 sg13g2_mux2_1 _10957_ (.A0(\ppu.tilemap.next_attr[0][0] ),
    .A1(\ppu.tilemap.attr[0][0] ),
    .S(net215),
    .X(_00825_));
 sg13g2_inv_1 _10958_ (.Y(_03196_),
    .A(\ppu.tilemap.attr[0][1] ));
 sg13g2_nor2_1 _10959_ (.A(\ppu.tilemap.next_attr[0][1] ),
    .B(net215),
    .Y(_03197_));
 sg13g2_a21oi_1 _10960_ (.A1(_03196_),
    .A2(net215),
    .Y(_00826_),
    .B1(_03197_));
 sg13g2_inv_1 _10961_ (.Y(_03198_),
    .A(\ppu.tilemap.attr[0][2] ));
 sg13g2_nor2_1 _10962_ (.A(\ppu.tilemap.next_attr[0][2] ),
    .B(net215),
    .Y(_03199_));
 sg13g2_a21oi_1 _10963_ (.A1(_03198_),
    .A2(net215),
    .Y(_00827_),
    .B1(_03199_));
 sg13g2_inv_1 _10964_ (.Y(_03200_),
    .A(\ppu.tilemap.attr[0][3] ));
 sg13g2_nor2_1 _10965_ (.A(\ppu.tilemap.next_attr[0][3] ),
    .B(net215),
    .Y(_03201_));
 sg13g2_a21oi_1 _10966_ (.A1(_03200_),
    .A2(net215),
    .Y(_00828_),
    .B1(_03201_));
 sg13g2_inv_1 _10967_ (.Y(_03202_),
    .A(\ppu.tilemap.attr[0][4] ));
 sg13g2_nor2_1 _10968_ (.A(\ppu.tilemap.next_attr[0][4] ),
    .B(_03195_),
    .Y(_03203_));
 sg13g2_a21oi_1 _10969_ (.A1(_03202_),
    .A2(net215),
    .Y(_00829_),
    .B1(_03203_));
 sg13g2_o21ai_1 _10970_ (.B1(_03190_),
    .Y(_03204_),
    .A1(_02540_),
    .A2(_02210_));
 sg13g2_buf_2 _10971_ (.A(_03204_),
    .X(_03205_));
 sg13g2_mux2_1 _10972_ (.A0(\ppu.tilemap.next_attr[1][0] ),
    .A1(\ppu.tilemap.attr[1][0] ),
    .S(_03205_),
    .X(_00830_));
 sg13g2_mux2_1 _10973_ (.A0(\ppu.tilemap.next_attr[1][1] ),
    .A1(\ppu.tilemap.attr[1][1] ),
    .S(_03205_),
    .X(_00831_));
 sg13g2_mux2_1 _10974_ (.A0(\ppu.tilemap.next_attr[1][2] ),
    .A1(\ppu.tilemap.attr[1][2] ),
    .S(_03205_),
    .X(_00832_));
 sg13g2_mux2_1 _10975_ (.A0(\ppu.tilemap.next_attr[1][3] ),
    .A1(\ppu.tilemap.attr[1][3] ),
    .S(_03205_),
    .X(_00833_));
 sg13g2_mux2_1 _10976_ (.A0(\ppu.tilemap.next_attr[1][4] ),
    .A1(\ppu.tilemap.attr[1][4] ),
    .S(_03205_),
    .X(_00834_));
 sg13g2_nand3_1 _10977_ (.B(net237),
    .C(_03189_),
    .A(_03193_),
    .Y(_03206_));
 sg13g2_buf_1 _10978_ (.A(_03206_),
    .X(_03207_));
 sg13g2_nor2_1 _10979_ (.A(net381),
    .B(net197),
    .Y(_03208_));
 sg13g2_a21oi_1 _10980_ (.A1(\ppu.tilemap.map_pixels[0][4] ),
    .A2(net197),
    .Y(_03209_),
    .B1(_03208_));
 sg13g2_inv_1 _10981_ (.Y(_03210_),
    .A(_03189_));
 sg13g2_a21oi_1 _10982_ (.A1(net263),
    .A2(_03210_),
    .Y(_03211_),
    .B1(net244));
 sg13g2_buf_1 _10983_ (.A(_03211_),
    .X(_03212_));
 sg13g2_o21ai_1 _10984_ (.B1(net197),
    .Y(_03213_),
    .A1(net264),
    .A2(_03212_));
 sg13g2_buf_2 _10985_ (.A(_03213_),
    .X(_03214_));
 sg13g2_nor2_1 _10986_ (.A(\ppu.tilemap.map_pixels[0][0] ),
    .B(_03214_),
    .Y(_03215_));
 sg13g2_a21oi_1 _10987_ (.A1(_03209_),
    .A2(_03214_),
    .Y(_00837_),
    .B1(_03215_));
 sg13g2_inv_1 _10988_ (.Y(_03216_),
    .A(\ppu.tilemap.map_pixels[0][14] ));
 sg13g2_buf_1 _10989_ (.A(_03212_),
    .X(_03217_));
 sg13g2_buf_1 _10990_ (.A(_03212_),
    .X(_03218_));
 sg13g2_nand2_1 _10991_ (.Y(_03219_),
    .A(net195),
    .B(\ppu.tilemap.map_pixels[0][10] ));
 sg13g2_o21ai_1 _10992_ (.B1(_03219_),
    .Y(_00838_),
    .A1(_03216_),
    .A2(net196));
 sg13g2_inv_1 _10993_ (.Y(_03220_),
    .A(\ppu.tilemap.map_pixels[0][15] ));
 sg13g2_nand2_1 _10994_ (.Y(_03221_),
    .A(net195),
    .B(\ppu.tilemap.map_pixels[0][11] ));
 sg13g2_o21ai_1 _10995_ (.B1(_03221_),
    .Y(_00839_),
    .A1(_03220_),
    .A2(net196));
 sg13g2_inv_1 _10996_ (.Y(_03222_),
    .A(\ppu.tilemap.map_pixels[0][12] ));
 sg13g2_inv_1 _10997_ (.Y(_03223_),
    .A(net244));
 sg13g2_nand2_1 _10998_ (.Y(_03224_),
    .A(_03223_),
    .B(\ppu.tilemap.map_pixels[0][0] ));
 sg13g2_a21oi_1 _10999_ (.A1(net405),
    .A2(net244),
    .Y(_03225_),
    .B1(net195));
 sg13g2_a22oi_1 _11000_ (.Y(_00840_),
    .B1(_03224_),
    .B2(_03225_),
    .A2(_03217_),
    .A1(_03222_));
 sg13g2_inv_1 _11001_ (.Y(_03226_),
    .A(\ppu.tilemap.map_pixels[0][1] ));
 sg13g2_nor2_1 _11002_ (.A(_03226_),
    .B(net244),
    .Y(_03227_));
 sg13g2_a21oi_1 _11003_ (.A1(net403),
    .A2(net244),
    .Y(_03228_),
    .B1(_03227_));
 sg13g2_nand2_1 _11004_ (.Y(_03229_),
    .A(net195),
    .B(\ppu.tilemap.map_pixels[0][13] ));
 sg13g2_o21ai_1 _11005_ (.B1(_03229_),
    .Y(_00841_),
    .A1(net196),
    .A2(_03228_));
 sg13g2_nand2_1 _11006_ (.Y(_03230_),
    .A(_03223_),
    .B(\ppu.tilemap.map_pixels[0][2] ));
 sg13g2_a21oi_1 _11007_ (.A1(net404),
    .A2(net244),
    .Y(_03231_),
    .B1(_03218_));
 sg13g2_a22oi_1 _11008_ (.Y(_00842_),
    .B1(_03230_),
    .B2(_03231_),
    .A2(net196),
    .A1(_03216_));
 sg13g2_nand2_1 _11009_ (.Y(_03232_),
    .A(_03223_),
    .B(\ppu.tilemap.map_pixels[0][3] ));
 sg13g2_a21oi_1 _11010_ (.A1(net408),
    .A2(net244),
    .Y(_03233_),
    .B1(net195));
 sg13g2_a22oi_1 _11011_ (.Y(_00843_),
    .B1(_03232_),
    .B2(_03233_),
    .A2(net196),
    .A1(_03220_));
 sg13g2_inv_1 _11012_ (.Y(_03234_),
    .A(\ppu.tilemap.map_pixels[0][5] ));
 sg13g2_o21ai_1 _11013_ (.B1(_03214_),
    .Y(_03235_),
    .A1(net403),
    .A2(net197));
 sg13g2_a21o_1 _11014_ (.A2(net197),
    .A1(_03234_),
    .B1(_03235_),
    .X(_03236_));
 sg13g2_o21ai_1 _11015_ (.B1(_03236_),
    .Y(_00844_),
    .A1(_03226_),
    .A2(_03214_));
 sg13g2_nor2_1 _11016_ (.A(_02685_),
    .B(net197),
    .Y(_03237_));
 sg13g2_a21oi_1 _11017_ (.A1(\ppu.tilemap.map_pixels[0][6] ),
    .A2(_03207_),
    .Y(_03238_),
    .B1(_03237_));
 sg13g2_nor2_1 _11018_ (.A(\ppu.tilemap.map_pixels[0][2] ),
    .B(_03214_),
    .Y(_03239_));
 sg13g2_a21oi_1 _11019_ (.A1(_03238_),
    .A2(_03214_),
    .Y(_00845_),
    .B1(_03239_));
 sg13g2_nor2_1 _11020_ (.A(_01867_),
    .B(net197),
    .Y(_03240_));
 sg13g2_a21oi_1 _11021_ (.A1(\ppu.tilemap.map_pixels[0][7] ),
    .A2(net197),
    .Y(_03241_),
    .B1(_03240_));
 sg13g2_nor2_1 _11022_ (.A(\ppu.tilemap.map_pixels[0][3] ),
    .B(_03214_),
    .Y(_03242_));
 sg13g2_a21oi_1 _11023_ (.A1(_03241_),
    .A2(_03214_),
    .Y(_00846_),
    .B1(_03242_));
 sg13g2_mux2_1 _11024_ (.A0(\ppu.tilemap.map_pixels[0][8] ),
    .A1(\ppu.tilemap.map_pixels[0][4] ),
    .S(net196),
    .X(_00847_));
 sg13g2_nor2_1 _11025_ (.A(\ppu.tilemap.map_pixels[0][9] ),
    .B(net195),
    .Y(_03243_));
 sg13g2_a21oi_1 _11026_ (.A1(_03234_),
    .A2(net196),
    .Y(_00848_),
    .B1(_03243_));
 sg13g2_mux2_1 _11027_ (.A0(\ppu.tilemap.map_pixels[0][10] ),
    .A1(\ppu.tilemap.map_pixels[0][6] ),
    .S(net196),
    .X(_00849_));
 sg13g2_mux2_1 _11028_ (.A0(\ppu.tilemap.map_pixels[0][11] ),
    .A1(\ppu.tilemap.map_pixels[0][7] ),
    .S(_03218_),
    .X(_00850_));
 sg13g2_nand2_1 _11029_ (.Y(_03244_),
    .A(net195),
    .B(\ppu.tilemap.map_pixels[0][8] ));
 sg13g2_o21ai_1 _11030_ (.B1(_03244_),
    .Y(_00851_),
    .A1(_03222_),
    .A2(_03217_));
 sg13g2_mux2_1 _11031_ (.A0(\ppu.tilemap.map_pixels[0][13] ),
    .A1(\ppu.tilemap.map_pixels[0][9] ),
    .S(net195),
    .X(_00852_));
 sg13g2_nor2_2 _11032_ (.A(_02209_),
    .B(_03191_),
    .Y(_03245_));
 sg13g2_inv_1 _11033_ (.Y(_03246_),
    .A(_03245_));
 sg13g2_buf_1 _11034_ (.A(net346),
    .X(_03247_));
 sg13g2_xor2_1 _11035_ (.B(\ppu.scroll_regs[2][0] ),
    .A(net293),
    .X(_03248_));
 sg13g2_nand2_1 _11036_ (.Y(_03249_),
    .A(_03248_),
    .B(net263));
 sg13g2_nand2_1 _11037_ (.Y(_03250_),
    .A(_03246_),
    .B(_03249_));
 sg13g2_inv_2 _11038_ (.Y(_03251_),
    .A(_03250_));
 sg13g2_nand3_1 _11039_ (.B(net237),
    .C(_02540_),
    .A(_03190_),
    .Y(_03252_));
 sg13g2_buf_1 _11040_ (.A(_03252_),
    .X(_03253_));
 sg13g2_o21ai_1 _11041_ (.B1(_03253_),
    .Y(_03254_),
    .A1(net264),
    .A2(_03251_));
 sg13g2_buf_2 _11042_ (.A(_03254_),
    .X(_03255_));
 sg13g2_nor2_1 _11043_ (.A(net381),
    .B(net194),
    .Y(_03256_));
 sg13g2_a21oi_1 _11044_ (.A1(\ppu.tilemap.map_pixels[1][4] ),
    .A2(net194),
    .Y(_03257_),
    .B1(_03256_));
 sg13g2_nor2_1 _11045_ (.A(\ppu.tilemap.map_pixels[1][0] ),
    .B(_03255_),
    .Y(_03258_));
 sg13g2_a21oi_1 _11046_ (.A1(_03255_),
    .A2(_03257_),
    .Y(_00853_),
    .B1(_03258_));
 sg13g2_inv_1 _11047_ (.Y(_03259_),
    .A(\ppu.tilemap.map_pixels[1][14] ));
 sg13g2_buf_1 _11048_ (.A(_03250_),
    .X(_03260_));
 sg13g2_nor2_1 _11049_ (.A(\ppu.tilemap.map_pixels[1][10] ),
    .B(net214),
    .Y(_03261_));
 sg13g2_a21oi_1 _11050_ (.A1(_03259_),
    .A2(net214),
    .Y(_00854_),
    .B1(_03261_));
 sg13g2_inv_1 _11051_ (.Y(_03262_),
    .A(\ppu.tilemap.map_pixels[1][15] ));
 sg13g2_nor2_1 _11052_ (.A(\ppu.tilemap.map_pixels[1][11] ),
    .B(net214),
    .Y(_03263_));
 sg13g2_a21oi_1 _11053_ (.A1(_03262_),
    .A2(net214),
    .Y(_00855_),
    .B1(_03263_));
 sg13g2_inv_1 _11054_ (.Y(_03264_),
    .A(\ppu.tilemap.map_pixels[1][12] ));
 sg13g2_nand2_1 _11055_ (.Y(_03265_),
    .A(_03245_),
    .B(net405));
 sg13g2_o21ai_1 _11056_ (.B1(_03246_),
    .Y(_03266_),
    .A1(\ppu.tilemap.map_pixels[1][0] ),
    .A2(_03249_));
 sg13g2_a22oi_1 _11057_ (.Y(_00856_),
    .B1(_03265_),
    .B2(_03266_),
    .A2(_03264_),
    .A1(_03251_));
 sg13g2_nand2_1 _11058_ (.Y(_03267_),
    .A(_03246_),
    .B(\ppu.tilemap.map_pixels[1][1] ));
 sg13g2_a22oi_1 _11059_ (.Y(_03268_),
    .B1(\ppu.tilemap.map_pixels[1][13] ),
    .B2(_03251_),
    .A2(_03245_),
    .A1(net403));
 sg13g2_o21ai_1 _11060_ (.B1(_03268_),
    .Y(_00857_),
    .A1(_03249_),
    .A2(_03267_));
 sg13g2_nand2_1 _11061_ (.Y(_03269_),
    .A(_03245_),
    .B(net404));
 sg13g2_o21ai_1 _11062_ (.B1(_03246_),
    .Y(_03270_),
    .A1(\ppu.tilemap.map_pixels[1][2] ),
    .A2(_03249_));
 sg13g2_a22oi_1 _11063_ (.Y(_00858_),
    .B1(_03269_),
    .B2(_03270_),
    .A2(_03259_),
    .A1(_03251_));
 sg13g2_nand2_1 _11064_ (.Y(_03271_),
    .A(_03246_),
    .B(\ppu.tilemap.map_pixels[1][3] ));
 sg13g2_a21oi_1 _11065_ (.A1(net408),
    .A2(_03245_),
    .Y(_03272_),
    .B1(_03251_));
 sg13g2_a22oi_1 _11066_ (.Y(_00859_),
    .B1(_03271_),
    .B2(_03272_),
    .A2(_03251_),
    .A1(_03262_));
 sg13g2_nor2_1 _11067_ (.A(net382),
    .B(net194),
    .Y(_03273_));
 sg13g2_a21oi_1 _11068_ (.A1(\ppu.tilemap.map_pixels[1][5] ),
    .A2(net194),
    .Y(_03274_),
    .B1(_03273_));
 sg13g2_nor2_1 _11069_ (.A(\ppu.tilemap.map_pixels[1][1] ),
    .B(_03255_),
    .Y(_03275_));
 sg13g2_a21oi_1 _11070_ (.A1(_03255_),
    .A2(_03274_),
    .Y(_00860_),
    .B1(_03275_));
 sg13g2_nor2_1 _11071_ (.A(_02685_),
    .B(net194),
    .Y(_03276_));
 sg13g2_a21oi_1 _11072_ (.A1(\ppu.tilemap.map_pixels[1][6] ),
    .A2(net194),
    .Y(_03277_),
    .B1(_03276_));
 sg13g2_nor2_1 _11073_ (.A(\ppu.tilemap.map_pixels[1][2] ),
    .B(_03255_),
    .Y(_03278_));
 sg13g2_a21oi_1 _11074_ (.A1(_03255_),
    .A2(_03277_),
    .Y(_00861_),
    .B1(_03278_));
 sg13g2_nor2_1 _11075_ (.A(_01867_),
    .B(net194),
    .Y(_03279_));
 sg13g2_a21oi_1 _11076_ (.A1(\ppu.tilemap.map_pixels[1][7] ),
    .A2(net194),
    .Y(_03280_),
    .B1(_03279_));
 sg13g2_nor2_1 _11077_ (.A(\ppu.tilemap.map_pixels[1][3] ),
    .B(_03255_),
    .Y(_03281_));
 sg13g2_a21oi_1 _11078_ (.A1(_03255_),
    .A2(_03280_),
    .Y(_00862_),
    .B1(_03281_));
 sg13g2_mux2_1 _11079_ (.A0(\ppu.tilemap.map_pixels[1][4] ),
    .A1(\ppu.tilemap.map_pixels[1][8] ),
    .S(_03260_),
    .X(_00863_));
 sg13g2_mux2_1 _11080_ (.A0(\ppu.tilemap.map_pixels[1][5] ),
    .A1(\ppu.tilemap.map_pixels[1][9] ),
    .S(_03260_),
    .X(_00864_));
 sg13g2_mux2_1 _11081_ (.A0(\ppu.tilemap.map_pixels[1][6] ),
    .A1(\ppu.tilemap.map_pixels[1][10] ),
    .S(net214),
    .X(_00865_));
 sg13g2_mux2_1 _11082_ (.A0(\ppu.tilemap.map_pixels[1][7] ),
    .A1(\ppu.tilemap.map_pixels[1][11] ),
    .S(net214),
    .X(_00866_));
 sg13g2_nor2_1 _11083_ (.A(\ppu.tilemap.map_pixels[1][8] ),
    .B(_03250_),
    .Y(_03282_));
 sg13g2_a21oi_1 _11084_ (.A1(_03264_),
    .A2(net214),
    .Y(_00867_),
    .B1(_03282_));
 sg13g2_mux2_1 _11085_ (.A0(\ppu.tilemap.map_pixels[1][9] ),
    .A1(\ppu.tilemap.map_pixels[1][13] ),
    .S(net214),
    .X(_00868_));
 sg13g2_nand3_1 _11086_ (.B(_01943_),
    .C(net251),
    .A(net295),
    .Y(_03283_));
 sg13g2_nand2_1 _11087_ (.Y(_03284_),
    .A(_03283_),
    .B(\ppu.tilemap.next_attr[0][0] ));
 sg13g2_o21ai_1 _11088_ (.B1(_03284_),
    .Y(_00869_),
    .A1(_01867_),
    .A2(_03283_));
 sg13g2_nand3_1 _11089_ (.B(_01943_),
    .C(net236),
    .A(net295),
    .Y(_03285_));
 sg13g2_buf_2 _11090_ (.A(_03285_),
    .X(_03286_));
 sg13g2_nand2_1 _11091_ (.Y(_03287_),
    .A(_03286_),
    .B(\ppu.tilemap.next_attr[0][1] ));
 sg13g2_o21ai_1 _11092_ (.B1(_03287_),
    .Y(_00870_),
    .A1(net381),
    .A2(_03286_));
 sg13g2_nand2_1 _11093_ (.Y(_03288_),
    .A(_03286_),
    .B(\ppu.tilemap.next_attr[0][2] ));
 sg13g2_o21ai_1 _11094_ (.B1(_03288_),
    .Y(_00871_),
    .A1(net382),
    .A2(_03286_));
 sg13g2_nand2_1 _11095_ (.Y(_03289_),
    .A(_03286_),
    .B(\ppu.tilemap.next_attr[0][3] ));
 sg13g2_o21ai_1 _11096_ (.B1(_03289_),
    .Y(_00872_),
    .A1(_02685_),
    .A2(_03286_));
 sg13g2_nand2_1 _11097_ (.Y(_03290_),
    .A(_03286_),
    .B(\ppu.tilemap.next_attr[0][4] ));
 sg13g2_o21ai_1 _11098_ (.B1(_03290_),
    .Y(_00873_),
    .A1(_01867_),
    .A2(_03286_));
 sg13g2_nand3_1 _11099_ (.B(_02095_),
    .C(net251),
    .A(net295),
    .Y(_03291_));
 sg13g2_nand2_1 _11100_ (.Y(_03292_),
    .A(_03291_),
    .B(\ppu.tilemap.next_attr[1][0] ));
 sg13g2_o21ai_1 _11101_ (.B1(_03292_),
    .Y(_00874_),
    .A1(_01867_),
    .A2(_03291_));
 sg13g2_nand3_1 _11102_ (.B(_02095_),
    .C(net236),
    .A(net295),
    .Y(_03293_));
 sg13g2_buf_2 _11103_ (.A(_03293_),
    .X(_03294_));
 sg13g2_nand2_1 _11104_ (.Y(_03295_),
    .A(_03294_),
    .B(\ppu.tilemap.next_attr[1][1] ));
 sg13g2_o21ai_1 _11105_ (.B1(_03295_),
    .Y(_00875_),
    .A1(net381),
    .A2(_03294_));
 sg13g2_nand2_1 _11106_ (.Y(_03296_),
    .A(_03294_),
    .B(\ppu.tilemap.next_attr[1][2] ));
 sg13g2_o21ai_1 _11107_ (.B1(_03296_),
    .Y(_00876_),
    .A1(net382),
    .A2(_03294_));
 sg13g2_nand2_1 _11108_ (.Y(_03297_),
    .A(_03294_),
    .B(\ppu.tilemap.next_attr[1][3] ));
 sg13g2_o21ai_1 _11109_ (.B1(_03297_),
    .Y(_00877_),
    .A1(_02685_),
    .A2(_03294_));
 sg13g2_nand2_1 _11110_ (.Y(_03298_),
    .A(_03294_),
    .B(\ppu.tilemap.next_attr[1][4] ));
 sg13g2_o21ai_1 _11111_ (.B1(_03298_),
    .Y(_00878_),
    .A1(_01867_),
    .A2(_03294_));
 sg13g2_buf_1 _11112_ (.A(\synth.controller.out_valid ),
    .X(_03299_));
 sg13g2_buf_1 _11113_ (.A(_03299_),
    .X(_03300_));
 sg13g2_inv_1 _11114_ (.Y(_03301_),
    .A(\synth.controller.out_reg[2] ));
 sg13g2_nand2_1 _11115_ (.Y(_03302_),
    .A(net380),
    .B(\synth.controller.out[0] ));
 sg13g2_o21ai_1 _11116_ (.B1(_03302_),
    .Y(_03303_),
    .A1(net380),
    .A2(_03301_));
 sg13g2_buf_1 _11117_ (.A(\synth.controller.sbio_tx.counter[3] ),
    .X(_03304_));
 sg13g2_buf_1 _11118_ (.A(\synth.controller.tx_source[1] ),
    .X(_03305_));
 sg13g2_buf_1 _11119_ (.A(\synth.controller.tx_source[0] ),
    .X(_03306_));
 sg13g2_inv_1 _11120_ (.Y(_03307_),
    .A(_03306_));
 sg13g2_nor2_1 _11121_ (.A(_03305_),
    .B(_03307_),
    .Y(_03308_));
 sg13g2_inv_1 _11122_ (.Y(_03309_),
    .A(_03308_));
 sg13g2_nor2_2 _11123_ (.A(_03304_),
    .B(_03309_),
    .Y(_03310_));
 sg13g2_nor2_1 _11124_ (.A(_03299_),
    .B(_03310_),
    .Y(_03311_));
 sg13g2_buf_1 _11125_ (.A(_03311_),
    .X(_03312_));
 sg13g2_buf_1 _11126_ (.A(_03312_),
    .X(_03313_));
 sg13g2_mux2_1 _11127_ (.A0(_03303_),
    .A1(\synth.controller.out_reg[0] ),
    .S(net213),
    .X(_00889_));
 sg13g2_nor2_1 _11128_ (.A(net380),
    .B(\synth.controller.out_reg[10] ),
    .Y(_03314_));
 sg13g2_buf_1 _11129_ (.A(_03299_),
    .X(_03315_));
 sg13g2_buf_1 _11130_ (.A(\synth.controller.out[10] ),
    .X(_03316_));
 sg13g2_nand2_1 _11131_ (.Y(_03317_),
    .A(net379),
    .B(_03316_));
 sg13g2_nor2b_1 _11132_ (.A(_03312_),
    .B_N(_03317_),
    .Y(_03318_));
 sg13g2_inv_1 _11133_ (.Y(_03319_),
    .A(_03299_));
 sg13g2_nand3_1 _11134_ (.B(net378),
    .C(\synth.controller.out_reg[12] ),
    .A(_03310_),
    .Y(_03320_));
 sg13g2_o21ai_1 _11135_ (.B1(_03320_),
    .Y(_00890_),
    .A1(_03314_),
    .A2(_03318_));
 sg13g2_inv_1 _11136_ (.Y(_03321_),
    .A(\synth.controller.out_reg[11] ));
 sg13g2_inv_1 _11137_ (.Y(_03322_),
    .A(\synth.controller.out[11] ));
 sg13g2_nand2_1 _11138_ (.Y(_03323_),
    .A(net378),
    .B(\synth.controller.out_reg[13] ));
 sg13g2_o21ai_1 _11139_ (.B1(_03323_),
    .Y(_03324_),
    .A1(net378),
    .A2(_03322_));
 sg13g2_buf_1 _11140_ (.A(_03312_),
    .X(_03325_));
 sg13g2_nor2_1 _11141_ (.A(_03324_),
    .B(net212),
    .Y(_03326_));
 sg13g2_a21oi_1 _11142_ (.A1(_03321_),
    .A2(net213),
    .Y(_00891_),
    .B1(_03326_));
 sg13g2_buf_1 _11143_ (.A(\synth.controller.out[12] ),
    .X(_03327_));
 sg13g2_a22oi_1 _11144_ (.Y(_03328_),
    .B1(\synth.controller.out_reg[12] ),
    .B2(net212),
    .A2(_03327_),
    .A1(net380));
 sg13g2_nand3_1 _11145_ (.B(net378),
    .C(\synth.controller.out_reg[14] ),
    .A(_03310_),
    .Y(_03329_));
 sg13g2_nand2_1 _11146_ (.Y(_00892_),
    .A(_03328_),
    .B(_03329_));
 sg13g2_buf_1 _11147_ (.A(\synth.controller.out[13] ),
    .X(_03330_));
 sg13g2_a22oi_1 _11148_ (.Y(_03331_),
    .B1(\synth.controller.out_reg[13] ),
    .B2(net212),
    .A2(_03330_),
    .A1(net380));
 sg13g2_nand3_1 _11149_ (.B(net378),
    .C(\synth.controller.out_reg[15] ),
    .A(_03310_),
    .Y(_03332_));
 sg13g2_nand2_1 _11150_ (.Y(_00893_),
    .A(_03331_),
    .B(_03332_));
 sg13g2_inv_1 _11151_ (.Y(_03333_),
    .A(\synth.controller.out[14] ));
 sg13g2_nand2_1 _11152_ (.Y(_03334_),
    .A(net212),
    .B(\synth.controller.out_reg[14] ));
 sg13g2_o21ai_1 _11153_ (.B1(_03334_),
    .Y(_00894_),
    .A1(net378),
    .A2(_03333_));
 sg13g2_inv_1 _11154_ (.Y(_03335_),
    .A(\synth.controller.out[15] ));
 sg13g2_nand2_1 _11155_ (.Y(_03336_),
    .A(net212),
    .B(\synth.controller.out_reg[15] ));
 sg13g2_o21ai_1 _11156_ (.B1(_03336_),
    .Y(_00895_),
    .A1(net378),
    .A2(_03335_));
 sg13g2_inv_1 _11157_ (.Y(_03337_),
    .A(\synth.controller.out_reg[3] ));
 sg13g2_nand2_1 _11158_ (.Y(_03338_),
    .A(net380),
    .B(\synth.controller.out[1] ));
 sg13g2_o21ai_1 _11159_ (.B1(_03338_),
    .Y(_03339_),
    .A1(net380),
    .A2(_03337_));
 sg13g2_mux2_1 _11160_ (.A0(_03339_),
    .A1(\synth.controller.out_reg[1] ),
    .S(net212),
    .X(_00896_));
 sg13g2_inv_1 _11161_ (.Y(_03340_),
    .A(\synth.controller.out_reg[4] ));
 sg13g2_nand2_1 _11162_ (.Y(_03341_),
    .A(net379),
    .B(\synth.controller.out[2] ));
 sg13g2_o21ai_1 _11163_ (.B1(_03341_),
    .Y(_03342_),
    .A1(net380),
    .A2(_03340_));
 sg13g2_nor2_1 _11164_ (.A(_03342_),
    .B(net212),
    .Y(_03343_));
 sg13g2_a21oi_1 _11165_ (.A1(_03301_),
    .A2(net213),
    .Y(_00897_),
    .B1(_03343_));
 sg13g2_inv_1 _11166_ (.Y(_03344_),
    .A(\synth.controller.out_reg[5] ));
 sg13g2_nand2_1 _11167_ (.Y(_03345_),
    .A(net379),
    .B(\synth.controller.out[3] ));
 sg13g2_o21ai_1 _11168_ (.B1(_03345_),
    .Y(_03346_),
    .A1(_03300_),
    .A2(_03344_));
 sg13g2_nor2_1 _11169_ (.A(_03346_),
    .B(net212),
    .Y(_03347_));
 sg13g2_a21oi_1 _11170_ (.A1(_03337_),
    .A2(net213),
    .Y(_00898_),
    .B1(_03347_));
 sg13g2_inv_1 _11171_ (.Y(_03348_),
    .A(\synth.controller.out_reg[6] ));
 sg13g2_nand2_1 _11172_ (.Y(_03349_),
    .A(net379),
    .B(\synth.controller.out[4] ));
 sg13g2_o21ai_1 _11173_ (.B1(_03349_),
    .Y(_03350_),
    .A1(_03315_),
    .A2(_03348_));
 sg13g2_nor2_1 _11174_ (.A(_03350_),
    .B(_03325_),
    .Y(_03351_));
 sg13g2_a21oi_1 _11175_ (.A1(_03340_),
    .A2(net213),
    .Y(_00899_),
    .B1(_03351_));
 sg13g2_inv_1 _11176_ (.Y(_03352_),
    .A(\synth.controller.out_reg[7] ));
 sg13g2_nand2_1 _11177_ (.Y(_03353_),
    .A(net379),
    .B(\synth.controller.out[5] ));
 sg13g2_o21ai_1 _11178_ (.B1(_03353_),
    .Y(_03354_),
    .A1(_03315_),
    .A2(_03352_));
 sg13g2_nor2_1 _11179_ (.A(_03354_),
    .B(_03325_),
    .Y(_03355_));
 sg13g2_a21oi_1 _11180_ (.A1(_03344_),
    .A2(net213),
    .Y(_00900_),
    .B1(_03355_));
 sg13g2_inv_1 _11181_ (.Y(_03356_),
    .A(\synth.controller.out_reg[8] ));
 sg13g2_nand2_1 _11182_ (.Y(_03357_),
    .A(_03299_),
    .B(\synth.controller.out[6] ));
 sg13g2_o21ai_1 _11183_ (.B1(_03357_),
    .Y(_03358_),
    .A1(net379),
    .A2(_03356_));
 sg13g2_nor2_1 _11184_ (.A(_03358_),
    .B(_03312_),
    .Y(_03359_));
 sg13g2_a21oi_1 _11185_ (.A1(_03348_),
    .A2(_03313_),
    .Y(_00901_),
    .B1(_03359_));
 sg13g2_inv_1 _11186_ (.Y(_03360_),
    .A(\synth.controller.out_reg[9] ));
 sg13g2_nand2_1 _11187_ (.Y(_03361_),
    .A(_03299_),
    .B(\synth.controller.out[7] ));
 sg13g2_o21ai_1 _11188_ (.B1(_03361_),
    .Y(_03362_),
    .A1(net379),
    .A2(_03360_));
 sg13g2_nor2_1 _11189_ (.A(_03362_),
    .B(_03312_),
    .Y(_03363_));
 sg13g2_a21oi_1 _11190_ (.A1(_03352_),
    .A2(_03313_),
    .Y(_00902_),
    .B1(_03363_));
 sg13g2_buf_1 _11191_ (.A(\synth.controller.out[8] ),
    .X(_03364_));
 sg13g2_nor2_1 _11192_ (.A(_03364_),
    .B(net378),
    .Y(_03365_));
 sg13g2_a221oi_1 _11193_ (.B2(_03356_),
    .C1(_03365_),
    .B1(net213),
    .A1(_03310_),
    .Y(_00903_),
    .A2(_03314_));
 sg13g2_buf_1 _11194_ (.A(\synth.controller.out[9] ),
    .X(_03366_));
 sg13g2_nand2_1 _11195_ (.Y(_03367_),
    .A(_03299_),
    .B(_03366_));
 sg13g2_o21ai_1 _11196_ (.B1(_03367_),
    .Y(_03368_),
    .A1(net379),
    .A2(_03321_));
 sg13g2_nor2_1 _11197_ (.A(_03368_),
    .B(_03312_),
    .Y(_03369_));
 sg13g2_a21oi_1 _11198_ (.A1(_03360_),
    .A2(net213),
    .Y(_00904_),
    .B1(_03369_));
 sg13g2_buf_2 _11199_ (.A(\rx_in_reg[0] ),
    .X(_03370_));
 sg13g2_inv_1 _11200_ (.Y(_03371_),
    .A(_03370_));
 sg13g2_buf_1 _11201_ (.A(\synth.controller.rx_counter[3] ),
    .X(_03372_));
 sg13g2_inv_1 _11202_ (.Y(_03373_),
    .A(net402));
 sg13g2_nand2_1 _11203_ (.Y(_03374_),
    .A(\synth.controller.rx_counter[1] ),
    .B(\synth.controller.rx_counter[0] ));
 sg13g2_inv_1 _11204_ (.Y(_03375_),
    .A(_03374_));
 sg13g2_nand2_1 _11205_ (.Y(_03376_),
    .A(_03375_),
    .B(\synth.controller.rx_counter[2] ));
 sg13g2_nor2_1 _11206_ (.A(_03373_),
    .B(_03376_),
    .Y(_03377_));
 sg13g2_inv_1 _11207_ (.Y(_03378_),
    .A(_03377_));
 sg13g2_buf_1 _11208_ (.A(\rx_in_reg[1] ),
    .X(_03379_));
 sg13g2_nand2_1 _11209_ (.Y(_03380_),
    .A(_03377_),
    .B(net401));
 sg13g2_nand2_1 _11210_ (.Y(_03381_),
    .A(_03380_),
    .B(\synth.controller.rx_sbs[0] ));
 sg13g2_o21ai_1 _11211_ (.B1(_03381_),
    .Y(_00931_),
    .A1(net377),
    .A2(_03378_));
 sg13g2_inv_1 _11212_ (.Y(_03382_),
    .A(\synth.controller.rx_sbs[1] ));
 sg13g2_inv_2 _11213_ (.Y(_03383_),
    .A(_03379_));
 sg13g2_a21oi_1 _11214_ (.A1(net377),
    .A2(_03383_),
    .Y(_03384_),
    .B1(_03378_));
 sg13g2_o21ai_1 _11215_ (.B1(_03380_),
    .Y(_00932_),
    .A1(_03382_),
    .A2(_03384_));
 sg13g2_buf_1 _11216_ (.A(\synth.controller.out_reg_valid ),
    .X(_03385_));
 sg13g2_inv_1 _11217_ (.Y(_03386_),
    .A(\synth.controller.tx_outstanding[1] ));
 sg13g2_nor2_1 _11218_ (.A(\synth.controller.sbio_credits[1] ),
    .B(_03386_),
    .Y(_03387_));
 sg13g2_inv_1 _11219_ (.Y(_03388_),
    .A(\synth.controller.tx_outstanding[0] ));
 sg13g2_nand2_1 _11220_ (.Y(_03389_),
    .A(_03388_),
    .B(\synth.controller.sbio_credits[0] ));
 sg13g2_inv_1 _11221_ (.Y(_03390_),
    .A(\synth.controller.tx_outstanding[2] ));
 sg13g2_a22oi_1 _11222_ (.Y(_03391_),
    .B1(\synth.controller.sbio_credits[1] ),
    .B2(_03386_),
    .A2(\synth.controller.sbio_credits[2] ),
    .A1(_03390_));
 sg13g2_o21ai_1 _11223_ (.B1(_03391_),
    .Y(_03392_),
    .A1(_03387_),
    .A2(_03389_));
 sg13g2_inv_1 _11224_ (.Y(_03393_),
    .A(\synth.controller.sweep_addr_index[1] ));
 sg13g2_and3_1 _11225_ (.X(_03394_),
    .A(_03393_),
    .B(\synth.controller.sweep_addr_index[0] ),
    .C(\synth.controller.sweep_addr_index[2] ));
 sg13g2_nand2b_1 _11226_ (.Y(_03395_),
    .B(_03394_),
    .A_N(\synth.controller.scanning_out ));
 sg13g2_nand2b_1 _11227_ (.Y(_03396_),
    .B(\synth.controller.tx_outstanding[2] ),
    .A_N(\synth.controller.sbio_credits[2] ));
 sg13g2_nand3_1 _11228_ (.B(_03395_),
    .C(_03396_),
    .A(_03392_),
    .Y(_03397_));
 sg13g2_inv_1 _11229_ (.Y(_03398_),
    .A(\synth.controller.ext_tx_request ));
 sg13g2_nand3b_1 _11230_ (.B(_03397_),
    .C(_03398_),
    .Y(_03399_),
    .A_N(_03385_));
 sg13g2_buf_1 _11231_ (.A(\synth.controller.sbio_tx.counter[0] ),
    .X(_03400_));
 sg13g2_buf_1 _11232_ (.A(\synth.controller.sbio_tx.counter[1] ),
    .X(_03401_));
 sg13g2_inv_1 _11233_ (.Y(_03402_),
    .A(_03401_));
 sg13g2_inv_1 _11234_ (.Y(_03403_),
    .A(\synth.controller.sbio_tx.counter[2] ));
 sg13g2_inv_2 _11235_ (.Y(_03404_),
    .A(_03304_));
 sg13g2_nor4_2 _11236_ (.A(_03400_),
    .B(_03402_),
    .C(_03403_),
    .Y(_03405_),
    .D(_03404_));
 sg13g2_nand2_2 _11237_ (.Y(_03406_),
    .A(_03399_),
    .B(_03405_));
 sg13g2_nor3_2 _11238_ (.A(_03385_),
    .B(\synth.controller.ext_tx_request ),
    .C(_03406_),
    .Y(_03407_));
 sg13g2_a21oi_1 _11239_ (.A1(_03307_),
    .A2(_03406_),
    .Y(_00959_),
    .B1(_03407_));
 sg13g2_inv_1 _11240_ (.Y(_03408_),
    .A(_03305_));
 sg13g2_o21ai_1 _11241_ (.B1(_03398_),
    .Y(_03409_),
    .A1(_03385_),
    .A2(_03394_));
 sg13g2_nor2_1 _11242_ (.A(_03409_),
    .B(_03406_),
    .Y(_03410_));
 sg13g2_a21oi_1 _11243_ (.A1(_03408_),
    .A2(_03406_),
    .Y(_00960_),
    .B1(_03410_));
 sg13g2_buf_2 _11244_ (.A(\synth.voice.delayed_s ),
    .X(_03411_));
 sg13g2_inv_1 _11245_ (.Y(_03412_),
    .A(_03411_));
 sg13g2_inv_1 _11246_ (.Y(_03413_),
    .A(\synth.voice.delayed_p[0] ));
 sg13g2_nand2_1 _11247_ (.Y(_03414_),
    .A(_01772_),
    .B(_01726_));
 sg13g2_buf_2 _11248_ (.A(_03414_),
    .X(_03415_));
 sg13g2_buf_1 _11249_ (.A(_03415_),
    .X(_03416_));
 sg13g2_buf_1 _11250_ (.A(net243),
    .X(_03417_));
 sg13g2_buf_1 _11251_ (.A(_03417_),
    .X(_03418_));
 sg13g2_buf_1 _11252_ (.A(net211),
    .X(_03419_));
 sg13g2_nor2_1 _11253_ (.A(\synth.voice.delayed_p[1] ),
    .B(net193),
    .Y(_03420_));
 sg13g2_a21o_1 _11254_ (.A2(net193),
    .A1(_03413_),
    .B1(_03420_),
    .X(_03421_));
 sg13g2_buf_1 _11255_ (.A(_03421_),
    .X(_03422_));
 sg13g2_buf_1 _11256_ (.A(\synth.controller.sweep_data_index[1] ),
    .X(_03423_));
 sg13g2_inv_2 _11257_ (.Y(_03424_),
    .A(net400));
 sg13g2_buf_2 _11258_ (.A(\synth.controller.sweep_data_index[0] ),
    .X(_03425_));
 sg13g2_nand2_1 _11259_ (.Y(_03426_),
    .A(_03424_),
    .B(_03425_));
 sg13g2_nor2_1 _11260_ (.A(\synth.controller.sample_credits[0] ),
    .B(\synth.controller.sample_credits[1] ),
    .Y(_03427_));
 sg13g2_nor2_1 _11261_ (.A(_00051_),
    .B(_03427_),
    .Y(_03428_));
 sg13g2_nand2b_1 _11262_ (.Y(_03429_),
    .B(_03428_),
    .A_N(_03426_));
 sg13g2_inv_1 _11263_ (.Y(_03430_),
    .A(_01724_));
 sg13g2_nand2_1 _11264_ (.Y(_03431_),
    .A(_03430_),
    .B(_00047_));
 sg13g2_o21ai_1 _11265_ (.B1(_01733_),
    .Y(_03432_),
    .A1(_03431_),
    .A2(_01755_));
 sg13g2_nor2_1 _11266_ (.A(_03429_),
    .B(_03432_),
    .Y(_03433_));
 sg13g2_buf_1 _11267_ (.A(_03433_),
    .X(_03434_));
 sg13g2_nor2_1 _11268_ (.A(_01737_),
    .B(net242),
    .Y(_03435_));
 sg13g2_o21ai_1 _11269_ (.B1(_03435_),
    .Y(_03436_),
    .A1(_03411_),
    .A2(net143));
 sg13g2_inv_1 _11270_ (.Y(_03437_),
    .A(_00115_));
 sg13g2_nor2_1 _11271_ (.A(_03437_),
    .B(_03415_),
    .Y(_03438_));
 sg13g2_a21oi_2 _11272_ (.B1(_03438_),
    .Y(_03439_),
    .A2(_03415_),
    .A1(_00114_));
 sg13g2_inv_1 _11273_ (.Y(_03440_),
    .A(_03439_));
 sg13g2_buf_1 _11274_ (.A(_00112_),
    .X(_03441_));
 sg13g2_a21oi_1 _11275_ (.A1(_01730_),
    .A2(_01734_),
    .Y(_03442_),
    .B1(_03430_));
 sg13g2_nor3_1 _11276_ (.A(_01724_),
    .B(_01734_),
    .C(_01756_),
    .Y(_03443_));
 sg13g2_nor2_1 _11277_ (.A(_03442_),
    .B(_03443_),
    .Y(_03444_));
 sg13g2_nand2_1 _11278_ (.Y(_03445_),
    .A(net242),
    .B(_03444_));
 sg13g2_buf_2 _11279_ (.A(_03445_),
    .X(_03446_));
 sg13g2_inv_4 _11280_ (.A(_03446_),
    .Y(_03447_));
 sg13g2_buf_8 _11281_ (.A(_03447_),
    .X(_03448_));
 sg13g2_nor2_2 _11282_ (.A(_03441_),
    .B(net183),
    .Y(_03449_));
 sg13g2_inv_1 _11283_ (.Y(_03450_),
    .A(\synth.voice.float_period[0][10] ));
 sg13g2_buf_1 _11284_ (.A(\synth.voice.float_period[1][10] ),
    .X(_03451_));
 sg13g2_nor2_1 _11285_ (.A(_03451_),
    .B(_03415_),
    .Y(_03452_));
 sg13g2_a21oi_1 _11286_ (.A1(_03450_),
    .A2(_03416_),
    .Y(_03453_),
    .B1(_03452_));
 sg13g2_buf_2 _11287_ (.A(_03453_),
    .X(_03454_));
 sg13g2_nand3_1 _11288_ (.B(_00113_),
    .C(_03454_),
    .A(_03449_),
    .Y(_03455_));
 sg13g2_buf_8 _11289_ (.A(_03446_),
    .X(_03456_));
 sg13g2_inv_2 _11290_ (.Y(_03457_),
    .A(_03454_));
 sg13g2_nand3_1 _11291_ (.B(_03441_),
    .C(_03457_),
    .A(net192),
    .Y(_03458_));
 sg13g2_nand2_1 _11292_ (.Y(_03459_),
    .A(_03455_),
    .B(_03458_));
 sg13g2_inv_1 _11293_ (.Y(_03460_),
    .A(_00113_));
 sg13g2_nand2b_1 _11294_ (.Y(_03461_),
    .B(_03460_),
    .A_N(_03441_));
 sg13g2_a21oi_1 _11295_ (.A1(_03456_),
    .A2(_03461_),
    .Y(_03462_),
    .B1(_00116_));
 sg13g2_xor2_1 _11296_ (.B(_03446_),
    .A(_00117_),
    .X(_03463_));
 sg13g2_xor2_1 _11297_ (.B(_03463_),
    .A(_03462_),
    .X(_03464_));
 sg13g2_a21o_1 _11298_ (.A2(_00117_),
    .A1(_03464_),
    .B1(_03457_),
    .X(_03465_));
 sg13g2_inv_1 _11299_ (.Y(_03466_),
    .A(_00116_));
 sg13g2_xnor2_1 _11300_ (.Y(_03467_),
    .A(_03466_),
    .B(net192));
 sg13g2_nand2_1 _11301_ (.Y(_03468_),
    .A(_03449_),
    .B(\synth.voice.oct_counter[1] ));
 sg13g2_xor2_1 _11302_ (.B(_03468_),
    .A(_03467_),
    .X(_03469_));
 sg13g2_o21ai_1 _11303_ (.B1(_03457_),
    .Y(_03470_),
    .A1(_03466_),
    .A2(_03469_));
 sg13g2_nor2b_1 _11304_ (.A(_03440_),
    .B_N(_03470_),
    .Y(_03471_));
 sg13g2_a22oi_1 _11305_ (.Y(_03472_),
    .B1(_03465_),
    .B2(_03471_),
    .A2(_03459_),
    .A1(_03440_));
 sg13g2_nor2_1 _11306_ (.A(\synth.voice.float_period[1][13] ),
    .B(_03415_),
    .Y(_03473_));
 sg13g2_nand2b_1 _11307_ (.Y(_03474_),
    .B(_03415_),
    .A_N(\synth.voice.float_period[0][13] ));
 sg13g2_nand2b_1 _11308_ (.Y(_03475_),
    .B(_03474_),
    .A_N(_03473_));
 sg13g2_nor2_1 _11309_ (.A(\synth.voice.float_period[1][12] ),
    .B(_03415_),
    .Y(_03476_));
 sg13g2_nand2b_1 _11310_ (.Y(_03477_),
    .B(_03415_),
    .A_N(\synth.voice.float_period[0][12] ));
 sg13g2_nand2b_2 _11311_ (.Y(_03478_),
    .B(_03477_),
    .A_N(_03476_));
 sg13g2_inv_2 _11312_ (.Y(_03479_),
    .A(_03478_));
 sg13g2_nand3_1 _11313_ (.B(_03475_),
    .C(_03479_),
    .A(_03472_),
    .Y(_03480_));
 sg13g2_inv_1 _11314_ (.Y(_03481_),
    .A(_03480_));
 sg13g2_buf_1 _11315_ (.A(\synth.voice.oct_counter[7] ),
    .X(_03482_));
 sg13g2_inv_1 _11316_ (.Y(_03483_),
    .A(_03482_));
 sg13g2_nor2_1 _11317_ (.A(_03483_),
    .B(net192),
    .Y(_03484_));
 sg13g2_nor2_1 _11318_ (.A(_03482_),
    .B(_03447_),
    .Y(_03485_));
 sg13g2_nor2_1 _11319_ (.A(_03484_),
    .B(_03485_),
    .Y(_03486_));
 sg13g2_inv_1 _11320_ (.Y(_03487_),
    .A(_03486_));
 sg13g2_nor2_1 _11321_ (.A(\synth.voice.oct_counter[6] ),
    .B(_03447_),
    .Y(_03488_));
 sg13g2_buf_2 _11322_ (.A(\synth.voice.oct_counter[4] ),
    .X(_03489_));
 sg13g2_xnor2_1 _11323_ (.Y(_03490_),
    .A(_03489_),
    .B(net192));
 sg13g2_nand3_1 _11324_ (.B(_03490_),
    .C(_03462_),
    .A(_03463_),
    .Y(_03491_));
 sg13g2_buf_1 _11325_ (.A(\synth.voice.oct_counter[3] ),
    .X(_03492_));
 sg13g2_o21ai_1 _11326_ (.B1(net183),
    .Y(_03493_),
    .A1(_03489_),
    .A2(_03492_));
 sg13g2_nand2_1 _11327_ (.Y(_03494_),
    .A(_03491_),
    .B(_03493_));
 sg13g2_inv_1 _11328_ (.Y(_03495_),
    .A(\synth.voice.oct_counter[5] ));
 sg13g2_nor2_1 _11329_ (.A(_03495_),
    .B(_03446_),
    .Y(_03496_));
 sg13g2_nor2_1 _11330_ (.A(\synth.voice.oct_counter[5] ),
    .B(_03447_),
    .Y(_03497_));
 sg13g2_nor2_1 _11331_ (.A(_03496_),
    .B(_03497_),
    .Y(_03498_));
 sg13g2_nand2_1 _11332_ (.Y(_03499_),
    .A(_03494_),
    .B(_03498_));
 sg13g2_inv_1 _11333_ (.Y(_03500_),
    .A(\synth.voice.oct_counter[6] ));
 sg13g2_nor2_1 _11334_ (.A(_03500_),
    .B(_03446_),
    .Y(_03501_));
 sg13g2_nor2_1 _11335_ (.A(_03496_),
    .B(_03501_),
    .Y(_03502_));
 sg13g2_o21ai_1 _11336_ (.B1(_03502_),
    .Y(_03503_),
    .A1(_03488_),
    .A2(_03499_));
 sg13g2_xnor2_1 _11337_ (.Y(_03504_),
    .A(_03487_),
    .B(_03503_));
 sg13g2_nand3_1 _11338_ (.B(_03483_),
    .C(_03454_),
    .A(_03504_),
    .Y(_03505_));
 sg13g2_nand2_1 _11339_ (.Y(_03506_),
    .A(_03498_),
    .B(_03490_));
 sg13g2_nor2_1 _11340_ (.A(_00116_),
    .B(_03456_),
    .Y(_03507_));
 sg13g2_a22oi_1 _11341_ (.Y(_03508_),
    .B1(_03507_),
    .B2(_03463_),
    .A2(net183),
    .A1(_03492_));
 sg13g2_o21ai_1 _11342_ (.B1(_03448_),
    .Y(_03509_),
    .A1(_03489_),
    .A2(\synth.voice.oct_counter[5] ));
 sg13g2_o21ai_1 _11343_ (.B1(_03509_),
    .Y(_03510_),
    .A1(_03506_),
    .A2(_03508_));
 sg13g2_inv_1 _11344_ (.Y(_03511_),
    .A(_03510_));
 sg13g2_nand2_1 _11345_ (.Y(_03512_),
    .A(_03463_),
    .B(_03467_));
 sg13g2_nor2_1 _11346_ (.A(_03512_),
    .B(_03506_),
    .Y(_03513_));
 sg13g2_inv_1 _11347_ (.Y(_03514_),
    .A(_03468_));
 sg13g2_nand2_1 _11348_ (.Y(_03515_),
    .A(_03513_),
    .B(_03514_));
 sg13g2_nand2_1 _11349_ (.Y(_03516_),
    .A(_03511_),
    .B(_03515_));
 sg13g2_nor2_1 _11350_ (.A(_03501_),
    .B(_03488_),
    .Y(_03517_));
 sg13g2_nand2_1 _11351_ (.Y(_03518_),
    .A(_03516_),
    .B(_03517_));
 sg13g2_inv_1 _11352_ (.Y(_03519_),
    .A(_03517_));
 sg13g2_nand3_1 _11353_ (.B(_03515_),
    .C(_03519_),
    .A(_03511_),
    .Y(_03520_));
 sg13g2_nand4_1 _11354_ (.B(_03520_),
    .C(_03500_),
    .A(_03518_),
    .Y(_03521_),
    .D(_03457_));
 sg13g2_nand3_1 _11355_ (.B(_03521_),
    .C(_03439_),
    .A(_03505_),
    .Y(_03522_));
 sg13g2_o21ai_1 _11356_ (.B1(_03508_),
    .Y(_03523_),
    .A1(_03468_),
    .A2(_03512_));
 sg13g2_xnor2_1 _11357_ (.Y(_03524_),
    .A(_03490_),
    .B(_03523_));
 sg13g2_nor3_1 _11358_ (.A(_03489_),
    .B(_03454_),
    .C(_03524_),
    .Y(_03525_));
 sg13g2_inv_1 _11359_ (.Y(_03526_),
    .A(_03498_));
 sg13g2_xnor2_1 _11360_ (.Y(_03527_),
    .A(_03526_),
    .B(_03494_));
 sg13g2_nand3_1 _11361_ (.B(_03495_),
    .C(_03454_),
    .A(_03527_),
    .Y(_03528_));
 sg13g2_nand3b_1 _11362_ (.B(_03440_),
    .C(_03528_),
    .Y(_03529_),
    .A_N(_03525_));
 sg13g2_nand3_1 _11363_ (.B(_03478_),
    .C(_03529_),
    .A(_03522_),
    .Y(_03530_));
 sg13g2_inv_1 _11364_ (.Y(_03531_),
    .A(_03475_));
 sg13g2_nand2_1 _11365_ (.Y(_03532_),
    .A(_03530_),
    .B(_03531_));
 sg13g2_xor2_1 _11366_ (.B(net192),
    .A(\synth.voice.oct_counter[10] ),
    .X(_03533_));
 sg13g2_a21oi_1 _11367_ (.A1(_03500_),
    .A2(_03483_),
    .Y(_03534_),
    .B1(net192));
 sg13g2_buf_1 _11368_ (.A(\synth.voice.oct_counter[9] ),
    .X(_03535_));
 sg13g2_nor2_1 _11369_ (.A(_03535_),
    .B(net183),
    .Y(_03536_));
 sg13g2_inv_1 _11370_ (.Y(_03537_),
    .A(_03536_));
 sg13g2_nand2_1 _11371_ (.Y(_03538_),
    .A(net183),
    .B(_03535_));
 sg13g2_nand2_1 _11372_ (.Y(_03539_),
    .A(_03537_),
    .B(_03538_));
 sg13g2_buf_1 _11373_ (.A(\synth.voice.oct_counter[8] ),
    .X(_03540_));
 sg13g2_inv_1 _11374_ (.Y(_03541_),
    .A(_03540_));
 sg13g2_nor2_1 _11375_ (.A(_03541_),
    .B(net192),
    .Y(_03542_));
 sg13g2_nor2_1 _11376_ (.A(_03540_),
    .B(_03447_),
    .Y(_03543_));
 sg13g2_nor2_1 _11377_ (.A(_03542_),
    .B(_03543_),
    .Y(_03544_));
 sg13g2_inv_1 _11378_ (.Y(_03545_),
    .A(_03544_));
 sg13g2_nor2_1 _11379_ (.A(_03539_),
    .B(_03545_),
    .Y(_03546_));
 sg13g2_nor2_1 _11380_ (.A(_03519_),
    .B(_03487_),
    .Y(_03547_));
 sg13g2_and2_1 _11381_ (.A(_03547_),
    .B(_03546_),
    .X(_03548_));
 sg13g2_nand2b_1 _11382_ (.Y(_03549_),
    .B(_03538_),
    .A_N(_03542_));
 sg13g2_a221oi_1 _11383_ (.B2(_03548_),
    .C1(_03549_),
    .B1(_03510_),
    .A1(_03534_),
    .Y(_03550_),
    .A2(_03546_));
 sg13g2_nand3_1 _11384_ (.B(_03513_),
    .C(_03514_),
    .A(_03548_),
    .Y(_03551_));
 sg13g2_nand2_1 _11385_ (.Y(_03552_),
    .A(_03550_),
    .B(_03551_));
 sg13g2_nand2b_1 _11386_ (.Y(_03553_),
    .B(_03552_),
    .A_N(_03533_));
 sg13g2_nand3_1 _11387_ (.B(_03551_),
    .C(_03533_),
    .A(_03550_),
    .Y(_03554_));
 sg13g2_nor3_1 _11388_ (.A(\synth.voice.oct_counter[10] ),
    .B(_03454_),
    .C(_03440_),
    .Y(_03555_));
 sg13g2_nand3_1 _11389_ (.B(_03554_),
    .C(_03555_),
    .A(_03553_),
    .Y(_03556_));
 sg13g2_inv_1 _11390_ (.Y(_03557_),
    .A(_03539_));
 sg13g2_inv_1 _11391_ (.Y(_03558_),
    .A(_03507_));
 sg13g2_nand2_1 _11392_ (.Y(_03559_),
    .A(_03463_),
    .B(_03490_));
 sg13g2_o21ai_1 _11393_ (.B1(net183),
    .Y(_03560_),
    .A1(_03489_),
    .A2(_03492_));
 sg13g2_o21ai_1 _11394_ (.B1(_03560_),
    .Y(_03561_),
    .A1(_03558_),
    .A2(_03559_));
 sg13g2_nand2_1 _11395_ (.Y(_03562_),
    .A(_03486_),
    .B(_03544_));
 sg13g2_nor3_1 _11396_ (.A(_03526_),
    .B(_03519_),
    .C(_03562_),
    .Y(_03563_));
 sg13g2_o21ai_1 _11397_ (.B1(_03448_),
    .Y(_03564_),
    .A1(_03482_),
    .A2(_03540_));
 sg13g2_o21ai_1 _11398_ (.B1(_03564_),
    .Y(_03565_),
    .A1(_03502_),
    .A2(_03562_));
 sg13g2_a21oi_1 _11399_ (.A1(_03561_),
    .A2(_03563_),
    .Y(_03566_),
    .B1(_03565_));
 sg13g2_inv_1 _11400_ (.Y(_03567_),
    .A(_03467_));
 sg13g2_nor3_1 _11401_ (.A(_00113_),
    .B(_03567_),
    .C(_03559_),
    .Y(_03568_));
 sg13g2_nand3_1 _11402_ (.B(_03568_),
    .C(_03449_),
    .A(_03563_),
    .Y(_03569_));
 sg13g2_nand2_1 _11403_ (.Y(_03570_),
    .A(_03566_),
    .B(_03569_));
 sg13g2_xnor2_1 _11404_ (.Y(_03571_),
    .A(_03557_),
    .B(_03570_));
 sg13g2_o21ai_1 _11405_ (.B1(_03454_),
    .Y(_03572_),
    .A1(_03535_),
    .A2(_03571_));
 sg13g2_nand3b_1 _11406_ (.B(_03523_),
    .C(_03547_),
    .Y(_03573_),
    .A_N(_03506_));
 sg13g2_inv_1 _11407_ (.Y(_03574_),
    .A(_03509_));
 sg13g2_a21oi_1 _11408_ (.A1(_03547_),
    .A2(_03574_),
    .Y(_03575_),
    .B1(_03534_));
 sg13g2_nand2_1 _11409_ (.Y(_03576_),
    .A(_03573_),
    .B(_03575_));
 sg13g2_nand2_1 _11410_ (.Y(_03577_),
    .A(_03576_),
    .B(_03544_));
 sg13g2_nand3_1 _11411_ (.B(_03545_),
    .C(_03575_),
    .A(_03573_),
    .Y(_03578_));
 sg13g2_nand3_1 _11412_ (.B(_03578_),
    .C(_03541_),
    .A(_03577_),
    .Y(_03579_));
 sg13g2_nand2_1 _11413_ (.Y(_03580_),
    .A(_03579_),
    .B(_03457_));
 sg13g2_nand3_1 _11414_ (.B(_03580_),
    .C(_03440_),
    .A(_03572_),
    .Y(_03581_));
 sg13g2_a21oi_1 _11415_ (.A1(_03556_),
    .A2(_03581_),
    .Y(_03582_),
    .B1(_03478_));
 sg13g2_nor2_1 _11416_ (.A(_03532_),
    .B(_03582_),
    .Y(_03583_));
 sg13g2_nor2_1 _11417_ (.A(_03481_),
    .B(_03583_),
    .Y(_03584_));
 sg13g2_nand2b_1 _11418_ (.Y(_03585_),
    .B(_03584_),
    .A_N(_03436_));
 sg13g2_nor3_1 _11419_ (.A(_03304_),
    .B(_03306_),
    .C(_03305_),
    .Y(_03586_));
 sg13g2_inv_1 _11420_ (.Y(_03587_),
    .A(_03586_));
 sg13g2_nor2_1 _11421_ (.A(\synth.controller.read_index_reg[3] ),
    .B(_03587_),
    .Y(_03588_));
 sg13g2_inv_1 _11422_ (.Y(_03589_),
    .A(_03588_));
 sg13g2_nor2_1 _11423_ (.A(\synth.controller.read_index_reg[2] ),
    .B(_03589_),
    .Y(_03590_));
 sg13g2_buf_1 _11424_ (.A(\synth.controller.read_index_reg[1] ),
    .X(_03591_));
 sg13g2_inv_1 _11425_ (.Y(_03592_),
    .A(_00057_));
 sg13g2_nor2_1 _11426_ (.A(_03592_),
    .B(_03587_),
    .Y(_03593_));
 sg13g2_inv_1 _11427_ (.Y(_03594_),
    .A(_03593_));
 sg13g2_nor2_1 _11428_ (.A(_03591_),
    .B(_03594_),
    .Y(_03595_));
 sg13g2_buf_1 _11429_ (.A(\synth.controller.write_index_reg[1] ),
    .X(_03596_));
 sg13g2_inv_1 _11430_ (.Y(_03597_),
    .A(_00111_));
 sg13g2_inv_1 _11431_ (.Y(_03598_),
    .A(\synth.controller.rx_sbs[0] ));
 sg13g2_nor3_1 _11432_ (.A(net402),
    .B(\synth.controller.rx_sbs[1] ),
    .C(_03598_),
    .Y(_03599_));
 sg13g2_inv_1 _11433_ (.Y(_03600_),
    .A(_03599_));
 sg13g2_nor2_1 _11434_ (.A(_03597_),
    .B(_03600_),
    .Y(_03601_));
 sg13g2_inv_1 _11435_ (.Y(_03602_),
    .A(_03601_));
 sg13g2_nor2_1 _11436_ (.A(_03596_),
    .B(_03602_),
    .Y(_03603_));
 sg13g2_buf_1 _11437_ (.A(\synth.controller.write_index_reg[2] ),
    .X(_03604_));
 sg13g2_nor2_1 _11438_ (.A(\synth.controller.write_index_reg[3] ),
    .B(_03600_),
    .Y(_03605_));
 sg13g2_inv_1 _11439_ (.Y(_03606_),
    .A(_03605_));
 sg13g2_nor2_1 _11440_ (.A(_03604_),
    .B(_03606_),
    .Y(_03607_));
 sg13g2_a22oi_1 _11441_ (.Y(_03608_),
    .B1(_03603_),
    .B2(_03607_),
    .A2(_03595_),
    .A1(_03590_));
 sg13g2_buf_1 _11442_ (.A(_03608_),
    .X(_03609_));
 sg13g2_nand2_1 _11443_ (.Y(_03610_),
    .A(_03585_),
    .B(_03609_));
 sg13g2_inv_1 _11444_ (.Y(_03611_),
    .A(_03609_));
 sg13g2_buf_1 _11445_ (.A(_03611_),
    .X(_03612_));
 sg13g2_nor3_1 _11446_ (.A(_03454_),
    .B(_03531_),
    .C(_03479_),
    .Y(_03613_));
 sg13g2_buf_2 _11447_ (.A(_03613_),
    .X(_03614_));
 sg13g2_buf_1 _11448_ (.A(_03614_),
    .X(_03615_));
 sg13g2_inv_1 _11449_ (.Y(_03616_),
    .A(_00098_));
 sg13g2_nor2_1 _11450_ (.A(_00097_),
    .B(net220),
    .Y(_03617_));
 sg13g2_a21o_1 _11451_ (.A2(_03417_),
    .A1(_03616_),
    .B1(_03617_),
    .X(_03618_));
 sg13g2_inv_1 _11452_ (.Y(_03619_),
    .A(_03618_));
 sg13g2_inv_1 _11453_ (.Y(_03620_),
    .A(_00100_));
 sg13g2_nor2_1 _11454_ (.A(_00099_),
    .B(net220),
    .Y(_03621_));
 sg13g2_a21o_1 _11455_ (.A2(net220),
    .A1(_03620_),
    .B1(_03621_),
    .X(_03622_));
 sg13g2_buf_1 _11456_ (.A(_03622_),
    .X(_03623_));
 sg13g2_nor2_1 _11457_ (.A(_03623_),
    .B(net160),
    .Y(_03624_));
 sg13g2_a21oi_1 _11458_ (.A1(_03615_),
    .A2(_03619_),
    .Y(_03625_),
    .B1(_03624_));
 sg13g2_nor2_1 _11459_ (.A(_03531_),
    .B(_03479_),
    .Y(_03626_));
 sg13g2_nand2_1 _11460_ (.Y(_03627_),
    .A(_03626_),
    .B(_03440_));
 sg13g2_buf_8 _11461_ (.A(_03627_),
    .X(_03628_));
 sg13g2_inv_8 _11462_ (.Y(_03629_),
    .A(_03628_));
 sg13g2_inv_1 _11463_ (.Y(_03630_),
    .A(_00103_));
 sg13g2_nor2_1 _11464_ (.A(_03630_),
    .B(net243),
    .Y(_03631_));
 sg13g2_a21oi_2 _11465_ (.B1(_03631_),
    .Y(_03632_),
    .A2(net243),
    .A1(_00104_));
 sg13g2_inv_1 _11466_ (.Y(_03633_),
    .A(_00102_));
 sg13g2_nor2_1 _11467_ (.A(_00101_),
    .B(net243),
    .Y(_03634_));
 sg13g2_a21o_1 _11468_ (.A2(net243),
    .A1(_03633_),
    .B1(_03634_),
    .X(_03635_));
 sg13g2_inv_1 _11469_ (.Y(_03636_),
    .A(_03635_));
 sg13g2_nand2_1 _11470_ (.Y(_03637_),
    .A(net160),
    .B(_03636_));
 sg13g2_o21ai_1 _11471_ (.B1(_03637_),
    .Y(_03638_),
    .A1(net160),
    .A2(_03632_));
 sg13g2_nor2_1 _11472_ (.A(net142),
    .B(_03638_),
    .Y(_03639_));
 sg13g2_a21o_1 _11473_ (.A2(net142),
    .A1(_03625_),
    .B1(_03639_),
    .X(_03640_));
 sg13g2_inv_1 _11474_ (.Y(_03641_),
    .A(_03640_));
 sg13g2_inv_1 _11475_ (.Y(_03642_),
    .A(_03623_));
 sg13g2_nor2_1 _11476_ (.A(_03635_),
    .B(net160),
    .Y(_03643_));
 sg13g2_a21oi_1 _11477_ (.A1(net160),
    .A2(_03642_),
    .Y(_03644_),
    .B1(_03643_));
 sg13g2_inv_1 _11478_ (.Y(_03645_),
    .A(_00096_));
 sg13g2_nor2_1 _11479_ (.A(_00090_),
    .B(net220),
    .Y(_03646_));
 sg13g2_a21o_1 _11480_ (.A2(net220),
    .A1(_03645_),
    .B1(_03646_),
    .X(_03647_));
 sg13g2_nor2_1 _11481_ (.A(_03619_),
    .B(_03614_),
    .Y(_03648_));
 sg13g2_a21oi_1 _11482_ (.A1(net160),
    .A2(_03647_),
    .Y(_03649_),
    .B1(_03648_));
 sg13g2_nor2_1 _11483_ (.A(_03628_),
    .B(_03649_),
    .Y(_03650_));
 sg13g2_a21oi_1 _11484_ (.A1(_03644_),
    .A2(net159),
    .Y(_03651_),
    .B1(_03650_));
 sg13g2_nand2_1 _11485_ (.Y(_03652_),
    .A(_03614_),
    .B(_03439_));
 sg13g2_inv_1 _11486_ (.Y(_03653_),
    .A(_03652_));
 sg13g2_inv_1 _11487_ (.Y(_03654_),
    .A(_00106_));
 sg13g2_nor2_1 _11488_ (.A(_00105_),
    .B(net243),
    .Y(_03655_));
 sg13g2_a21o_1 _11489_ (.A2(net243),
    .A1(_03654_),
    .B1(_03655_),
    .X(_03656_));
 sg13g2_buf_1 _11490_ (.A(_03656_),
    .X(_03657_));
 sg13g2_inv_1 _11491_ (.Y(_03658_),
    .A(_03657_));
 sg13g2_nor2_2 _11492_ (.A(_03614_),
    .B(net142),
    .Y(_03659_));
 sg13g2_inv_1 _11493_ (.Y(_03660_),
    .A(_00060_));
 sg13g2_nor2_1 _11494_ (.A(_03660_),
    .B(_03416_),
    .Y(_03661_));
 sg13g2_a21oi_1 _11495_ (.A1(_00107_),
    .A2(net243),
    .Y(_03662_),
    .B1(_03661_));
 sg13g2_inv_1 _11496_ (.Y(_03663_),
    .A(_03662_));
 sg13g2_a22oi_1 _11497_ (.Y(_03664_),
    .B1(_03659_),
    .B2(_03663_),
    .A2(_03658_),
    .A1(_03653_));
 sg13g2_nand2_1 _11498_ (.Y(_03665_),
    .A(_03638_),
    .B(net142));
 sg13g2_nand2_1 _11499_ (.Y(_03666_),
    .A(_03664_),
    .B(_03665_));
 sg13g2_nand3_1 _11500_ (.B(_03651_),
    .C(_03666_),
    .A(_03641_),
    .Y(_03667_));
 sg13g2_buf_1 _11501_ (.A(_00054_),
    .X(_03668_));
 sg13g2_inv_1 _11502_ (.Y(_03669_),
    .A(_03668_));
 sg13g2_nor2_1 _11503_ (.A(_03632_),
    .B(_03652_),
    .Y(_03670_));
 sg13g2_inv_2 _11504_ (.Y(_03671_),
    .A(_03659_));
 sg13g2_nor2_1 _11505_ (.A(_03657_),
    .B(_03671_),
    .Y(_03672_));
 sg13g2_nor2_1 _11506_ (.A(net159),
    .B(_03644_),
    .Y(_03673_));
 sg13g2_nor3_1 _11507_ (.A(_03670_),
    .B(_03672_),
    .C(_03673_),
    .Y(_03674_));
 sg13g2_nor3_1 _11508_ (.A(_03669_),
    .B(_03611_),
    .C(_03674_),
    .Y(_03675_));
 sg13g2_inv_1 _11509_ (.Y(_03676_),
    .A(_00095_));
 sg13g2_nor2_1 _11510_ (.A(_00089_),
    .B(net220),
    .Y(_03677_));
 sg13g2_a21o_1 _11511_ (.A2(net220),
    .A1(_03676_),
    .B1(_03677_),
    .X(_03678_));
 sg13g2_buf_1 _11512_ (.A(_03678_),
    .X(_03679_));
 sg13g2_inv_1 _11513_ (.Y(_03680_),
    .A(_03647_));
 sg13g2_nor2_1 _11514_ (.A(_03680_),
    .B(_03614_),
    .Y(_03681_));
 sg13g2_a21o_1 _11515_ (.A2(_03679_),
    .A1(_03615_),
    .B1(_03681_),
    .X(_03682_));
 sg13g2_inv_1 _11516_ (.Y(_03683_),
    .A(_03682_));
 sg13g2_nor2_1 _11517_ (.A(net142),
    .B(_03625_),
    .Y(_03684_));
 sg13g2_a21oi_2 _11518_ (.B1(_03684_),
    .Y(_03685_),
    .A2(_03683_),
    .A1(_03629_));
 sg13g2_nor2b_2 _11519_ (.A(net159),
    .B_N(_03614_),
    .Y(_03686_));
 sg13g2_nor2b_1 _11520_ (.A(net211),
    .B_N(_00134_),
    .Y(_03687_));
 sg13g2_a21oi_1 _11521_ (.A1(_00133_),
    .A2(net211),
    .Y(_03688_),
    .B1(_03687_));
 sg13g2_nand2_1 _11522_ (.Y(_03689_),
    .A(_03686_),
    .B(_03688_));
 sg13g2_nand2_1 _11523_ (.Y(_03690_),
    .A(_03685_),
    .B(_03689_));
 sg13g2_nand2_1 _11524_ (.Y(_03691_),
    .A(_03675_),
    .B(_03690_));
 sg13g2_nor2b_1 _11525_ (.A(net211),
    .B_N(_00136_),
    .Y(_03692_));
 sg13g2_a21oi_1 _11526_ (.A1(_00135_),
    .A2(net211),
    .Y(_03693_),
    .B1(_03692_));
 sg13g2_nand2_1 _11527_ (.Y(_03694_),
    .A(net142),
    .B(_03693_));
 sg13g2_inv_1 _11528_ (.Y(_03695_),
    .A(_03679_));
 sg13g2_inv_1 _11529_ (.Y(_03696_),
    .A(_00093_));
 sg13g2_nor2_1 _11530_ (.A(_00087_),
    .B(net220),
    .Y(_03697_));
 sg13g2_a21o_1 _11531_ (.A2(net211),
    .A1(_03696_),
    .B1(_03697_),
    .X(_03698_));
 sg13g2_buf_1 _11532_ (.A(_03698_),
    .X(_03699_));
 sg13g2_nand2_1 _11533_ (.Y(_03700_),
    .A(_03614_),
    .B(_03699_));
 sg13g2_o21ai_1 _11534_ (.B1(_03700_),
    .Y(_03701_),
    .A1(net160),
    .A2(_03695_));
 sg13g2_inv_1 _11535_ (.Y(_03702_),
    .A(_00091_));
 sg13g2_nor2_1 _11536_ (.A(_00084_),
    .B(net211),
    .Y(_03703_));
 sg13g2_a21o_1 _11537_ (.A2(net211),
    .A1(_03702_),
    .B1(_03703_),
    .X(_03704_));
 sg13g2_nor2b_1 _11538_ (.A(_03614_),
    .B_N(_03699_),
    .Y(_03705_));
 sg13g2_a21o_1 _11539_ (.A2(_03704_),
    .A1(net160),
    .B1(_03705_),
    .X(_03706_));
 sg13g2_nor2_1 _11540_ (.A(net159),
    .B(_03706_),
    .Y(_03707_));
 sg13g2_a21oi_1 _11541_ (.A1(net159),
    .A2(_03683_),
    .Y(_03708_),
    .B1(_03707_));
 sg13g2_nor2_1 _11542_ (.A(_00138_),
    .B(_03418_),
    .Y(_03709_));
 sg13g2_nand2b_1 _11543_ (.Y(_03710_),
    .B(_03418_),
    .A_N(_00137_));
 sg13g2_nand2b_1 _11544_ (.Y(_03711_),
    .B(_03710_),
    .A_N(_03709_));
 sg13g2_nand3b_1 _11545_ (.B(_03711_),
    .C(_03671_),
    .Y(_03712_),
    .A_N(_03708_));
 sg13g2_o21ai_1 _11546_ (.B1(_03712_),
    .Y(_03713_),
    .A1(_03694_),
    .A2(_03701_));
 sg13g2_nor2_1 _11547_ (.A(net142),
    .B(_03649_),
    .Y(_03714_));
 sg13g2_a21o_1 _11548_ (.A2(net142),
    .A1(_03701_),
    .B1(_03714_),
    .X(_03715_));
 sg13g2_nand2_1 _11549_ (.Y(_03716_),
    .A(_03715_),
    .B(_03694_));
 sg13g2_nor2_1 _11550_ (.A(_03689_),
    .B(_03685_),
    .Y(_03717_));
 sg13g2_a21oi_1 _11551_ (.A1(_03713_),
    .A2(_03716_),
    .Y(_03718_),
    .B1(_03717_));
 sg13g2_nor3_1 _11552_ (.A(_03667_),
    .B(_03691_),
    .C(_03718_),
    .Y(_03719_));
 sg13g2_a22oi_1 _11553_ (.Y(_03720_),
    .B1(_03719_),
    .B2(_03610_),
    .A2(net182),
    .A1(\synth.voice.delayed_p[1] ));
 sg13g2_o21ai_1 _11554_ (.B1(_03720_),
    .Y(_01098_),
    .A1(_03412_),
    .A2(_03610_));
 sg13g2_inv_2 _11555_ (.Y(_03721_),
    .A(_03425_));
 sg13g2_nand3_1 _11556_ (.B(net400),
    .C(\synth.voice.genblk4[6].next_state_scan[7] ),
    .A(_03721_),
    .Y(_03722_));
 sg13g2_buf_1 _11557_ (.A(_03425_),
    .X(_03723_));
 sg13g2_nand3_1 _11558_ (.B(net376),
    .C(\synth.voice.genblk4[7].next_state_scan[1] ),
    .A(net400),
    .Y(_03724_));
 sg13g2_nand2_1 _11559_ (.Y(_03725_),
    .A(_03424_),
    .B(\synth.voice.genblk4[7].next_state_scan[11] ));
 sg13g2_nand3_1 _11560_ (.B(_03724_),
    .C(_03725_),
    .A(_03722_),
    .Y(_03726_));
 sg13g2_buf_2 _11561_ (.A(\synth.controller.sweep_data_index[2] ),
    .X(_03727_));
 sg13g2_nor2_1 _11562_ (.A(net400),
    .B(_03727_),
    .Y(_03728_));
 sg13g2_inv_2 _11563_ (.Y(_03729_),
    .A(_03728_));
 sg13g2_nand2_1 _11564_ (.Y(_03730_),
    .A(_03726_),
    .B(net334));
 sg13g2_inv_1 _11565_ (.Y(_03731_),
    .A(\synth.voice.float_period[0][5] ));
 sg13g2_buf_1 _11566_ (.A(\synth.voice.float_period[1][5] ),
    .X(_03732_));
 sg13g2_nand2_1 _11567_ (.Y(_03733_),
    .A(net376),
    .B(_03732_));
 sg13g2_o21ai_1 _11568_ (.B1(_03733_),
    .Y(_03734_),
    .A1(net376),
    .A2(_03731_));
 sg13g2_buf_1 _11569_ (.A(_03728_),
    .X(_03735_));
 sg13g2_nand2_1 _11570_ (.Y(_03736_),
    .A(_03734_),
    .B(net333));
 sg13g2_a21oi_1 _11571_ (.A1(_03730_),
    .A2(_03736_),
    .Y(_03737_),
    .B1(\synth.controller.reg_wdata[1] ));
 sg13g2_nor2_1 _11572_ (.A(_03425_),
    .B(_03424_),
    .Y(_03738_));
 sg13g2_buf_1 _11573_ (.A(_03738_),
    .X(_03739_));
 sg13g2_nand2_1 _11574_ (.Y(_03740_),
    .A(net292),
    .B(\synth.voice.genblk4[6].next_state_scan[6] ));
 sg13g2_nand3_1 _11575_ (.B(net376),
    .C(\synth.voice.genblk4[7].next_state_scan[0] ),
    .A(net400),
    .Y(_03741_));
 sg13g2_buf_1 _11576_ (.A(_03424_),
    .X(_03742_));
 sg13g2_nand2_1 _11577_ (.Y(_03743_),
    .A(net332),
    .B(\synth.voice.genblk4[7].next_state_scan[10] ));
 sg13g2_nand3_1 _11578_ (.B(_03741_),
    .C(_03743_),
    .A(_03740_),
    .Y(_03744_));
 sg13g2_nand2_1 _11579_ (.Y(_03745_),
    .A(_03744_),
    .B(net334));
 sg13g2_buf_1 _11580_ (.A(\synth.voice.float_period[0][4] ),
    .X(_03746_));
 sg13g2_inv_1 _11581_ (.Y(_03747_),
    .A(\synth.voice.float_period[1][4] ));
 sg13g2_a21oi_1 _11582_ (.A1(net376),
    .A2(_03747_),
    .Y(_03748_),
    .B1(net334));
 sg13g2_o21ai_1 _11583_ (.B1(_03748_),
    .Y(_03749_),
    .A1(net376),
    .A2(_03746_));
 sg13g2_buf_1 _11584_ (.A(\synth.controller.reg_wdata[2] ),
    .X(_03750_));
 sg13g2_a21oi_1 _11585_ (.A1(_03745_),
    .A2(_03749_),
    .Y(_03751_),
    .B1(_03750_));
 sg13g2_nor2_1 _11586_ (.A(_03737_),
    .B(_03751_),
    .Y(_03752_));
 sg13g2_nand3_1 _11587_ (.B(\synth.controller.reg_wdata[1] ),
    .C(_03736_),
    .A(_03730_),
    .Y(_03753_));
 sg13g2_a22oi_1 _11588_ (.Y(_03754_),
    .B1(\synth.voice.genblk4[6].next_state_scan[8] ),
    .B2(net292),
    .A2(\synth.voice.genblk4[7].next_state_scan[12] ),
    .A1(net332));
 sg13g2_nand2_1 _11589_ (.Y(_03755_),
    .A(net400),
    .B(_03425_));
 sg13g2_inv_1 _11590_ (.Y(_03756_),
    .A(_03755_));
 sg13g2_buf_1 _11591_ (.A(\synth.voice.genblk4[7].next_state_scan[2] ),
    .X(_03757_));
 sg13g2_nand2_1 _11592_ (.Y(_03758_),
    .A(_03756_),
    .B(_03757_));
 sg13g2_nand2_1 _11593_ (.Y(_03759_),
    .A(_03754_),
    .B(_03758_));
 sg13g2_nand2_1 _11594_ (.Y(_03760_),
    .A(_03759_),
    .B(net334));
 sg13g2_inv_1 _11595_ (.Y(_03761_),
    .A(\synth.voice.float_period[0][6] ));
 sg13g2_buf_1 _11596_ (.A(\synth.voice.float_period[1][6] ),
    .X(_03762_));
 sg13g2_o21ai_1 _11597_ (.B1(_03728_),
    .Y(_03763_),
    .A1(_03721_),
    .A2(_03762_));
 sg13g2_a21oi_1 _11598_ (.A1(_03721_),
    .A2(_03761_),
    .Y(_03764_),
    .B1(_03763_));
 sg13g2_buf_1 _11599_ (.A(\synth.controller.reg_wdata[0] ),
    .X(_03765_));
 sg13g2_nor2b_1 _11600_ (.A(_03764_),
    .B_N(_03765_),
    .Y(_03766_));
 sg13g2_nand2_1 _11601_ (.Y(_03767_),
    .A(_03760_),
    .B(_03766_));
 sg13g2_nand2_1 _11602_ (.Y(_03768_),
    .A(_03753_),
    .B(_03767_));
 sg13g2_nand2_1 _11603_ (.Y(_03769_),
    .A(_03752_),
    .B(_03768_));
 sg13g2_nand3_1 _11604_ (.B(_03749_),
    .C(_03750_),
    .A(_03745_),
    .Y(_03770_));
 sg13g2_nand2_1 _11605_ (.Y(_03771_),
    .A(_03769_),
    .B(_03770_));
 sg13g2_inv_1 _11606_ (.Y(_03772_),
    .A(\synth.voice.mods[1][3] ));
 sg13g2_buf_1 _11607_ (.A(\synth.voice.genblk4[7].next_state_scan[9] ),
    .X(_03773_));
 sg13g2_a22oi_1 _11608_ (.Y(_03774_),
    .B1(\synth.voice.genblk4[6].next_state_scan[5] ),
    .B2(net292),
    .A2(_03773_),
    .A1(net332));
 sg13g2_o21ai_1 _11609_ (.B1(_03774_),
    .Y(_03775_),
    .A1(_03772_),
    .A2(_03755_));
 sg13g2_nand2_1 _11610_ (.Y(_03776_),
    .A(_03775_),
    .B(net334));
 sg13g2_nor2_1 _11611_ (.A(net376),
    .B(\synth.voice.float_period[0][3] ),
    .Y(_03777_));
 sg13g2_nor2_1 _11612_ (.A(\synth.voice.float_period[1][3] ),
    .B(_03721_),
    .Y(_03778_));
 sg13g2_nor3_1 _11613_ (.A(_03777_),
    .B(_03778_),
    .C(net334),
    .Y(_03779_));
 sg13g2_inv_1 _11614_ (.Y(_03780_),
    .A(_03779_));
 sg13g2_nand2_1 _11615_ (.Y(_03781_),
    .A(_03776_),
    .B(_03780_));
 sg13g2_inv_1 _11616_ (.Y(_03782_),
    .A(\synth.controller.reg_wdata[3] ));
 sg13g2_nand2_1 _11617_ (.Y(_03783_),
    .A(_03781_),
    .B(_03782_));
 sg13g2_nand2_1 _11618_ (.Y(_03784_),
    .A(_03771_),
    .B(_03783_));
 sg13g2_a22oi_1 _11619_ (.Y(_03785_),
    .B1(\synth.voice.genblk4[6].next_state_scan[4] ),
    .B2(net292),
    .A2(\synth.voice.genblk4[7].next_state_scan[8] ),
    .A1(net332));
 sg13g2_nand2_1 _11620_ (.Y(_03786_),
    .A(_03756_),
    .B(\synth.voice.mods[1][2] ));
 sg13g2_a21o_1 _11621_ (.A2(_03786_),
    .A1(_03785_),
    .B1(net333),
    .X(_03787_));
 sg13g2_nor2_1 _11622_ (.A(net376),
    .B(\synth.voice.float_period[0][2] ),
    .Y(_03788_));
 sg13g2_nor2_1 _11623_ (.A(\synth.voice.float_period[1][2] ),
    .B(_03721_),
    .Y(_03789_));
 sg13g2_nor3_1 _11624_ (.A(_03788_),
    .B(_03789_),
    .C(net334),
    .Y(_03790_));
 sg13g2_inv_1 _11625_ (.Y(_03791_),
    .A(_03790_));
 sg13g2_nand2_1 _11626_ (.Y(_03792_),
    .A(_03787_),
    .B(_03791_));
 sg13g2_inv_1 _11627_ (.Y(_03793_),
    .A(_03792_));
 sg13g2_nor2_1 _11628_ (.A(_03782_),
    .B(_03781_),
    .Y(_03794_));
 sg13g2_a21oi_1 _11629_ (.A1(_03793_),
    .A2(\synth.controller.reg_wdata[4] ),
    .Y(_03795_),
    .B1(_03794_));
 sg13g2_nand2_1 _11630_ (.Y(_03796_),
    .A(_03784_),
    .B(_03795_));
 sg13g2_a22oi_1 _11631_ (.Y(_03797_),
    .B1(\synth.voice.genblk4[6].next_state_scan[3] ),
    .B2(_03739_),
    .A2(\synth.voice.genblk4[7].next_state_scan[7] ),
    .A1(net332));
 sg13g2_nand2_1 _11632_ (.Y(_03798_),
    .A(_03756_),
    .B(\synth.voice.genblk4[6].next_state_scan[13] ));
 sg13g2_a21o_1 _11633_ (.A2(_03798_),
    .A1(_03797_),
    .B1(net333),
    .X(_03799_));
 sg13g2_nor2_1 _11634_ (.A(_03723_),
    .B(\synth.voice.float_period[0][1] ),
    .Y(_03800_));
 sg13g2_buf_1 _11635_ (.A(_03721_),
    .X(_03801_));
 sg13g2_nor2_1 _11636_ (.A(\synth.voice.float_period[1][1] ),
    .B(_03801_),
    .Y(_03802_));
 sg13g2_nor3_1 _11637_ (.A(_03800_),
    .B(_03802_),
    .C(_03729_),
    .Y(_03803_));
 sg13g2_inv_1 _11638_ (.Y(_03804_),
    .A(_03803_));
 sg13g2_nand2_1 _11639_ (.Y(_03805_),
    .A(_03799_),
    .B(_03804_));
 sg13g2_inv_1 _11640_ (.Y(_03806_),
    .A(\synth.controller.reg_wdata[4] ));
 sg13g2_a22oi_1 _11641_ (.Y(_03807_),
    .B1(_03806_),
    .B2(_03792_),
    .A2(_00121_),
    .A1(_03805_));
 sg13g2_nand2_1 _11642_ (.Y(_03808_),
    .A(_03796_),
    .B(_03807_));
 sg13g2_buf_1 _11643_ (.A(net334),
    .X(_03809_));
 sg13g2_buf_1 _11644_ (.A(_03723_),
    .X(_03810_));
 sg13g2_nor2_1 _11645_ (.A(net330),
    .B(\synth.voice.float_period[0][0] ),
    .Y(_03811_));
 sg13g2_nor2_1 _11646_ (.A(\synth.voice.float_period[1][0] ),
    .B(_03801_),
    .Y(_03812_));
 sg13g2_nor3_2 _11647_ (.A(_03811_),
    .B(_03812_),
    .C(_03809_),
    .Y(_03813_));
 sg13g2_inv_1 _11648_ (.Y(_03814_),
    .A(_03813_));
 sg13g2_o21ai_1 _11649_ (.B1(_03814_),
    .Y(_03815_),
    .A1(_00121_),
    .A2(_03805_));
 sg13g2_inv_1 _11650_ (.Y(_03816_),
    .A(\synth.voice.genblk4[6].next_state_scan[12] ));
 sg13g2_buf_1 _11651_ (.A(\synth.voice.genblk4[7].next_state_scan[6] ),
    .X(_03817_));
 sg13g2_buf_1 _11652_ (.A(\synth.voice.genblk4[6].next_state_scan[2] ),
    .X(_03818_));
 sg13g2_a22oi_1 _11653_ (.Y(_03819_),
    .B1(_03818_),
    .B2(net292),
    .A2(_03817_),
    .A1(net332));
 sg13g2_o21ai_1 _11654_ (.B1(_03819_),
    .Y(_03820_),
    .A1(_03816_),
    .A2(_03755_));
 sg13g2_nand2_1 _11655_ (.Y(_03821_),
    .A(_03820_),
    .B(net291));
 sg13g2_nor2b_1 _11656_ (.A(_03815_),
    .B_N(_03821_),
    .Y(_03822_));
 sg13g2_nand3_1 _11657_ (.B(net291),
    .C(_03822_),
    .A(_03808_),
    .Y(_03823_));
 sg13g2_buf_1 _11658_ (.A(_00119_),
    .X(_03824_));
 sg13g2_nand2_2 _11659_ (.Y(_03825_),
    .A(net333),
    .B(_03824_));
 sg13g2_nand2_1 _11660_ (.Y(_03826_),
    .A(_03823_),
    .B(_03825_));
 sg13g2_nand2_1 _11661_ (.Y(_03827_),
    .A(_03821_),
    .B(_03749_));
 sg13g2_inv_1 _11662_ (.Y(_03828_),
    .A(_03827_));
 sg13g2_nand2_1 _11663_ (.Y(_03829_),
    .A(_03826_),
    .B(_03828_));
 sg13g2_nand3_1 _11664_ (.B(_03825_),
    .C(_03827_),
    .A(_03823_),
    .Y(_03830_));
 sg13g2_buf_1 _11665_ (.A(_03830_),
    .X(_03831_));
 sg13g2_nand2_2 _11666_ (.Y(_03832_),
    .A(_03829_),
    .B(_03831_));
 sg13g2_nand2_1 _11667_ (.Y(_03833_),
    .A(_03799_),
    .B(_03736_));
 sg13g2_nand2_1 _11668_ (.Y(_03834_),
    .A(_03808_),
    .B(_03822_));
 sg13g2_buf_1 _11669_ (.A(_03824_),
    .X(_03835_));
 sg13g2_nand2_1 _11670_ (.Y(_03836_),
    .A(_03834_),
    .B(net375));
 sg13g2_nand2_1 _11671_ (.Y(_03837_),
    .A(_03836_),
    .B(_03825_));
 sg13g2_nand2b_1 _11672_ (.Y(_03838_),
    .B(_03837_),
    .A_N(_03833_));
 sg13g2_nand3_1 _11673_ (.B(_03833_),
    .C(_03825_),
    .A(_03836_),
    .Y(_03839_));
 sg13g2_buf_1 _11674_ (.A(_03839_),
    .X(_03840_));
 sg13g2_nand2_1 _11675_ (.Y(_03841_),
    .A(_03838_),
    .B(_03840_));
 sg13g2_nor2_1 _11676_ (.A(_03832_),
    .B(_03841_),
    .Y(_03842_));
 sg13g2_nor2_1 _11677_ (.A(net375),
    .B(_03780_),
    .Y(_03843_));
 sg13g2_nor2_1 _11678_ (.A(_03835_),
    .B(_03791_),
    .Y(_03844_));
 sg13g2_nor2_1 _11679_ (.A(_03843_),
    .B(_03844_),
    .Y(_03845_));
 sg13g2_inv_1 _11680_ (.Y(_03846_),
    .A(_03845_));
 sg13g2_a21oi_1 _11681_ (.A1(_03836_),
    .A2(_03825_),
    .Y(_03847_),
    .B1(_03833_));
 sg13g2_a21oi_1 _11682_ (.A1(_03840_),
    .A2(_03831_),
    .Y(_03848_),
    .B1(_03847_));
 sg13g2_a21oi_1 _11683_ (.A1(_03842_),
    .A2(_03846_),
    .Y(_03849_),
    .B1(_03848_));
 sg13g2_nor2_1 _11684_ (.A(_03824_),
    .B(_03809_),
    .Y(_03850_));
 sg13g2_nor2_1 _11685_ (.A(_03850_),
    .B(_03779_),
    .Y(_03851_));
 sg13g2_nor2_1 _11686_ (.A(_03851_),
    .B(_03843_),
    .Y(_03852_));
 sg13g2_xor2_1 _11687_ (.B(_03790_),
    .A(_03850_),
    .X(_03853_));
 sg13g2_nand2_1 _11688_ (.Y(_03854_),
    .A(_03852_),
    .B(_03853_));
 sg13g2_nor3_1 _11689_ (.A(_03854_),
    .B(_03832_),
    .C(_03841_),
    .Y(_03855_));
 sg13g2_nand2_1 _11690_ (.Y(_03856_),
    .A(_03836_),
    .B(_03735_));
 sg13g2_nand2_1 _11691_ (.Y(_03857_),
    .A(_03856_),
    .B(_03804_));
 sg13g2_nor2_1 _11692_ (.A(_03804_),
    .B(_03856_),
    .Y(_03858_));
 sg13g2_a21oi_2 _11693_ (.B1(_03858_),
    .Y(_03859_),
    .A2(_03813_),
    .A1(_03857_));
 sg13g2_inv_1 _11694_ (.Y(_03860_),
    .A(_03859_));
 sg13g2_nand2_1 _11695_ (.Y(_03861_),
    .A(_03855_),
    .B(_03860_));
 sg13g2_nand2_1 _11696_ (.Y(_03862_),
    .A(_03849_),
    .B(_03861_));
 sg13g2_buf_1 _11697_ (.A(\synth.voice.float_period[1][7] ),
    .X(_03863_));
 sg13g2_inv_1 _11698_ (.Y(_03864_),
    .A(\synth.voice.float_period[0][7] ));
 sg13g2_a21oi_1 _11699_ (.A1(net331),
    .A2(_03864_),
    .Y(_03865_),
    .B1(net291));
 sg13g2_o21ai_1 _11700_ (.B1(_03865_),
    .Y(_03866_),
    .A1(net331),
    .A2(_03863_));
 sg13g2_nand2_1 _11701_ (.Y(_03867_),
    .A(_03776_),
    .B(_03866_));
 sg13g2_xnor2_1 _11702_ (.Y(_03868_),
    .A(net375),
    .B(_03867_));
 sg13g2_inv_1 _11703_ (.Y(_03869_),
    .A(_03868_));
 sg13g2_nand2b_1 _11704_ (.Y(_03870_),
    .B(_03787_),
    .A_N(_03764_));
 sg13g2_xnor2_1 _11705_ (.Y(_03871_),
    .A(_03835_),
    .B(_03870_));
 sg13g2_inv_1 _11706_ (.Y(_03872_),
    .A(_03871_));
 sg13g2_nor2_1 _11707_ (.A(_03869_),
    .B(_03872_),
    .Y(_03873_));
 sg13g2_buf_1 _11708_ (.A(\synth.voice.float_period[1][9] ),
    .X(_03874_));
 sg13g2_inv_1 _11709_ (.Y(_03875_),
    .A(\synth.voice.float_period[0][9] ));
 sg13g2_a21oi_1 _11710_ (.A1(net331),
    .A2(_03875_),
    .Y(_03876_),
    .B1(net291));
 sg13g2_o21ai_1 _11711_ (.B1(_03876_),
    .Y(_03877_),
    .A1(net331),
    .A2(_03874_));
 sg13g2_nand2_1 _11712_ (.Y(_03878_),
    .A(_03730_),
    .B(_03877_));
 sg13g2_xnor2_1 _11713_ (.Y(_03879_),
    .A(net375),
    .B(_03878_));
 sg13g2_inv_1 _11714_ (.Y(_03880_),
    .A(_03879_));
 sg13g2_inv_1 _11715_ (.Y(_03881_),
    .A(\synth.voice.float_period[0][8] ));
 sg13g2_a21oi_1 _11716_ (.A1(net331),
    .A2(_03881_),
    .Y(_03882_),
    .B1(net291));
 sg13g2_o21ai_1 _11717_ (.B1(_03882_),
    .Y(_03883_),
    .A1(net331),
    .A2(\synth.voice.float_period[1][8] ));
 sg13g2_nand2_1 _11718_ (.Y(_03884_),
    .A(_03745_),
    .B(_03883_));
 sg13g2_xnor2_1 _11719_ (.Y(_03885_),
    .A(net375),
    .B(_03884_));
 sg13g2_inv_1 _11720_ (.Y(_03886_),
    .A(_03885_));
 sg13g2_nor2_1 _11721_ (.A(_03880_),
    .B(_03886_),
    .Y(_03887_));
 sg13g2_nand2_1 _11722_ (.Y(_03888_),
    .A(_03873_),
    .B(_03887_));
 sg13g2_inv_1 _11723_ (.Y(_03889_),
    .A(net375));
 sg13g2_a22oi_1 _11724_ (.Y(_03890_),
    .B1(\synth.voice.genblk4[6].next_state_scan[11] ),
    .B2(net292),
    .A2(\synth.voice.mods[2][9] ),
    .A1(_03742_));
 sg13g2_nand2_1 _11725_ (.Y(_03891_),
    .A(_03756_),
    .B(\synth.voice.genblk4[7].next_state_scan[5] ));
 sg13g2_nand2_1 _11726_ (.Y(_03892_),
    .A(_03890_),
    .B(_03891_));
 sg13g2_inv_1 _11727_ (.Y(_03893_),
    .A(\synth.voice.float_period[1][13] ));
 sg13g2_o21ai_1 _11728_ (.B1(net333),
    .Y(_03894_),
    .A1(net330),
    .A2(\synth.voice.float_period[0][13] ));
 sg13g2_a21oi_1 _11729_ (.A1(net330),
    .A2(_03893_),
    .Y(_03895_),
    .B1(_03894_));
 sg13g2_a21oi_1 _11730_ (.A1(_03892_),
    .A2(net291),
    .Y(_03896_),
    .B1(_03895_));
 sg13g2_xnor2_1 _11731_ (.Y(_03897_),
    .A(net329),
    .B(_03896_));
 sg13g2_inv_1 _11732_ (.Y(_03898_),
    .A(_03897_));
 sg13g2_inv_1 _11733_ (.Y(_03899_),
    .A(\synth.voice.float_period[1][12] ));
 sg13g2_o21ai_1 _11734_ (.B1(net333),
    .Y(_03900_),
    .A1(net330),
    .A2(\synth.voice.float_period[0][12] ));
 sg13g2_a21oi_1 _11735_ (.A1(net330),
    .A2(_03899_),
    .Y(_03901_),
    .B1(_03900_));
 sg13g2_buf_1 _11736_ (.A(\synth.voice.genblk4[7].next_state_scan[4] ),
    .X(_03902_));
 sg13g2_a22oi_1 _11737_ (.Y(_03903_),
    .B1(_03902_),
    .B2(_03756_),
    .A2(\synth.voice.mods[2][8] ),
    .A1(net332));
 sg13g2_nand2_1 _11738_ (.Y(_03904_),
    .A(net292),
    .B(\synth.voice.genblk4[6].next_state_scan[10] ));
 sg13g2_a21oi_1 _11739_ (.A1(_03903_),
    .A2(_03904_),
    .Y(_03905_),
    .B1(net333));
 sg13g2_nor3_1 _11740_ (.A(net329),
    .B(_03901_),
    .C(_03905_),
    .Y(_03906_));
 sg13g2_o21ai_1 _11741_ (.B1(net329),
    .Y(_03907_),
    .A1(_03901_),
    .A2(_03905_));
 sg13g2_nor2b_1 _11742_ (.A(_03906_),
    .B_N(_03907_),
    .Y(_03908_));
 sg13g2_inv_1 _11743_ (.Y(_03909_),
    .A(_03908_));
 sg13g2_nor2_1 _11744_ (.A(_03898_),
    .B(_03909_),
    .Y(_03910_));
 sg13g2_a21oi_1 _11745_ (.A1(net331),
    .A2(_03450_),
    .Y(_03911_),
    .B1(net291));
 sg13g2_o21ai_1 _11746_ (.B1(_03911_),
    .Y(_03912_),
    .A1(net331),
    .A2(_03451_));
 sg13g2_nand2_1 _11747_ (.Y(_03913_),
    .A(_03760_),
    .B(_03912_));
 sg13g2_xnor2_1 _11748_ (.Y(_03914_),
    .A(net375),
    .B(_03913_));
 sg13g2_inv_1 _11749_ (.Y(_03915_),
    .A(_03914_));
 sg13g2_a22oi_1 _11750_ (.Y(_03916_),
    .B1(\synth.voice.genblk4[6].next_state_scan[9] ),
    .B2(net292),
    .A2(\synth.voice.genblk4[7].next_state_scan[13] ),
    .A1(_03742_));
 sg13g2_buf_1 _11751_ (.A(\synth.voice.genblk4[7].next_state_scan[3] ),
    .X(_03917_));
 sg13g2_nand2_1 _11752_ (.Y(_03918_),
    .A(_03756_),
    .B(_03917_));
 sg13g2_nand2_1 _11753_ (.Y(_03919_),
    .A(_03916_),
    .B(_03918_));
 sg13g2_inv_1 _11754_ (.Y(_03920_),
    .A(\synth.voice.float_period[1][11] ));
 sg13g2_o21ai_1 _11755_ (.B1(net333),
    .Y(_03921_),
    .A1(net330),
    .A2(\synth.voice.float_period[0][11] ));
 sg13g2_a21oi_1 _11756_ (.A1(net330),
    .A2(_03920_),
    .Y(_03922_),
    .B1(_03921_));
 sg13g2_a21oi_1 _11757_ (.A1(_03919_),
    .A2(net291),
    .Y(_03923_),
    .B1(_03922_));
 sg13g2_xnor2_1 _11758_ (.Y(_03924_),
    .A(net329),
    .B(_03923_));
 sg13g2_inv_1 _11759_ (.Y(_03925_),
    .A(_03924_));
 sg13g2_nor2_1 _11760_ (.A(_03915_),
    .B(_03925_),
    .Y(_03926_));
 sg13g2_nand2_1 _11761_ (.Y(_03927_),
    .A(_03910_),
    .B(_03926_));
 sg13g2_nor2_1 _11762_ (.A(_03888_),
    .B(_03927_),
    .Y(_03928_));
 sg13g2_nand2_1 _11763_ (.Y(_03929_),
    .A(_03862_),
    .B(_03928_));
 sg13g2_buf_1 _11764_ (.A(\synth.controller.reg_waddr[2] ),
    .X(_03930_));
 sg13g2_nand2_1 _11765_ (.Y(_03931_),
    .A(_03907_),
    .B(_03896_));
 sg13g2_nand2_1 _11766_ (.Y(_03932_),
    .A(_03913_),
    .B(net329));
 sg13g2_inv_2 _11767_ (.Y(_03933_),
    .A(_03930_));
 sg13g2_a21oi_1 _11768_ (.A1(_03932_),
    .A2(_03923_),
    .Y(_03934_),
    .B1(_03933_));
 sg13g2_a21oi_1 _11769_ (.A1(_03870_),
    .A2(net329),
    .Y(_03935_),
    .B1(_03867_));
 sg13g2_nor2_1 _11770_ (.A(_03933_),
    .B(_03935_),
    .Y(_03936_));
 sg13g2_a21oi_1 _11771_ (.A1(_03884_),
    .A2(net329),
    .Y(_03937_),
    .B1(_03878_));
 sg13g2_nor2_1 _11772_ (.A(_03933_),
    .B(_03937_),
    .Y(_03938_));
 sg13g2_a21oi_1 _11773_ (.A1(_03936_),
    .A2(_03887_),
    .Y(_03939_),
    .B1(_03938_));
 sg13g2_nor2_1 _11774_ (.A(_03927_),
    .B(_03939_),
    .Y(_03940_));
 sg13g2_a221oi_1 _11775_ (.B2(_03934_),
    .C1(_03940_),
    .B1(_03910_),
    .A1(_03930_),
    .Y(_03941_),
    .A2(_03931_));
 sg13g2_nand2_1 _11776_ (.Y(_03942_),
    .A(_03929_),
    .B(_03941_));
 sg13g2_nand2_1 _11777_ (.Y(_03943_),
    .A(_03942_),
    .B(net375));
 sg13g2_nand3_1 _11778_ (.B(_03889_),
    .C(_03941_),
    .A(_03929_),
    .Y(_03944_));
 sg13g2_buf_1 _11779_ (.A(\synth.controller.reg_waddr[1] ),
    .X(_03945_));
 sg13g2_buf_1 _11780_ (.A(\synth.controller.reg_wdata[6] ),
    .X(_03946_));
 sg13g2_inv_1 _11781_ (.Y(_03947_),
    .A(_03946_));
 sg13g2_buf_2 _11782_ (.A(\synth.voice.sweep_oct_counter[0] ),
    .X(_03948_));
 sg13g2_nand2_1 _11783_ (.Y(_03949_),
    .A(_03947_),
    .B(_03948_));
 sg13g2_nand2_1 _11784_ (.Y(_03950_),
    .A(_03948_),
    .B(\synth.voice.sweep_oct_counter[1] ));
 sg13g2_inv_1 _11785_ (.Y(_03951_),
    .A(_03950_));
 sg13g2_buf_1 _11786_ (.A(_03946_),
    .X(_03952_));
 sg13g2_inv_1 _11787_ (.Y(_03953_),
    .A(\synth.voice.sweep_oct_counter[2] ));
 sg13g2_nand3_1 _11788_ (.B(net374),
    .C(_03953_),
    .A(_03951_),
    .Y(_03954_));
 sg13g2_o21ai_1 _11789_ (.B1(_03954_),
    .Y(_03955_),
    .A1(\synth.voice.sweep_oct_counter[1] ),
    .A2(_03949_));
 sg13g2_buf_1 _11790_ (.A(\synth.controller.reg_wdata[7] ),
    .X(_03956_));
 sg13g2_a21oi_1 _11791_ (.A1(net374),
    .A2(_03948_),
    .Y(_03957_),
    .B1(_03956_));
 sg13g2_a21o_1 _11792_ (.A2(_03956_),
    .A1(_03955_),
    .B1(_03957_),
    .X(_03958_));
 sg13g2_buf_2 _11793_ (.A(\synth.controller.reg_waddr[0] ),
    .X(_03959_));
 sg13g2_inv_1 _11794_ (.Y(_03960_),
    .A(_03959_));
 sg13g2_buf_2 _11795_ (.A(\synth.voice.sweep_oct_counter[6] ),
    .X(_03961_));
 sg13g2_inv_1 _11796_ (.Y(_03962_),
    .A(\synth.voice.sweep_oct_counter[5] ));
 sg13g2_inv_1 _11797_ (.Y(_03963_),
    .A(\synth.voice.sweep_oct_counter[4] ));
 sg13g2_inv_1 _11798_ (.Y(_03964_),
    .A(\synth.voice.sweep_oct_counter[3] ));
 sg13g2_nor2_1 _11799_ (.A(_03953_),
    .B(_03950_),
    .Y(_03965_));
 sg13g2_inv_1 _11800_ (.Y(_03966_),
    .A(_03965_));
 sg13g2_nor2_1 _11801_ (.A(_03964_),
    .B(_03966_),
    .Y(_03967_));
 sg13g2_inv_1 _11802_ (.Y(_03968_),
    .A(_03967_));
 sg13g2_nor2_1 _11803_ (.A(_03963_),
    .B(_03968_),
    .Y(_03969_));
 sg13g2_inv_1 _11804_ (.Y(_03970_),
    .A(_03969_));
 sg13g2_nor2_1 _11805_ (.A(_03962_),
    .B(_03970_),
    .Y(_03971_));
 sg13g2_inv_1 _11806_ (.Y(_03972_),
    .A(_03971_));
 sg13g2_o21ai_1 _11807_ (.B1(net374),
    .Y(_03973_),
    .A1(_03961_),
    .A2(_03972_));
 sg13g2_o21ai_1 _11808_ (.B1(_03947_),
    .Y(_03974_),
    .A1(\synth.voice.sweep_oct_counter[5] ),
    .A2(_03970_));
 sg13g2_nand3_1 _11809_ (.B(_03956_),
    .C(_03974_),
    .A(_03973_),
    .Y(_03975_));
 sg13g2_nand3_1 _11810_ (.B(net374),
    .C(\synth.voice.sweep_oct_counter[3] ),
    .A(_03963_),
    .Y(_03976_));
 sg13g2_o21ai_1 _11811_ (.B1(_03976_),
    .Y(_03977_),
    .A1(net374),
    .A2(\synth.voice.sweep_oct_counter[3] ));
 sg13g2_inv_2 _11812_ (.Y(_03978_),
    .A(_03956_));
 sg13g2_nand3_1 _11813_ (.B(_03978_),
    .C(_03965_),
    .A(_03977_),
    .Y(_03979_));
 sg13g2_a21oi_1 _11814_ (.A1(_03975_),
    .A2(_03979_),
    .Y(_03980_),
    .B1(_03960_));
 sg13g2_a21oi_1 _11815_ (.A1(_03958_),
    .A2(_03960_),
    .Y(_03981_),
    .B1(_03980_));
 sg13g2_buf_1 _11816_ (.A(\synth.voice.sweep_oct_counter[11] ),
    .X(_03982_));
 sg13g2_inv_1 _11817_ (.Y(_03983_),
    .A(\synth.voice.sweep_oct_counter[12] ));
 sg13g2_nand3_1 _11818_ (.B(net374),
    .C(_03982_),
    .A(_03983_),
    .Y(_03984_));
 sg13g2_o21ai_1 _11819_ (.B1(_03984_),
    .Y(_03985_),
    .A1(net374),
    .A2(_03982_));
 sg13g2_nand2_1 _11820_ (.Y(_03986_),
    .A(_03985_),
    .B(_03978_));
 sg13g2_inv_1 _11821_ (.Y(_03987_),
    .A(\synth.voice.sweep_oct_counter[8] ));
 sg13g2_buf_1 _11822_ (.A(\synth.voice.sweep_oct_counter[7] ),
    .X(_03988_));
 sg13g2_nand3_1 _11823_ (.B(_03961_),
    .C(_03988_),
    .A(_03971_),
    .Y(_03989_));
 sg13g2_nor2_1 _11824_ (.A(_03987_),
    .B(_03989_),
    .Y(_03990_));
 sg13g2_nand3_1 _11825_ (.B(\synth.voice.sweep_oct_counter[9] ),
    .C(\synth.voice.sweep_oct_counter[10] ),
    .A(_03990_),
    .Y(_03991_));
 sg13g2_buf_1 _11826_ (.A(_03991_),
    .X(_03992_));
 sg13g2_o21ai_1 _11827_ (.B1(_03959_),
    .Y(_03993_),
    .A1(_03986_),
    .A2(_03992_));
 sg13g2_inv_1 _11828_ (.Y(_03994_),
    .A(\synth.voice.sweep_oct_counter[13] ));
 sg13g2_nand4_1 _11829_ (.B(_03956_),
    .C(\synth.voice.sweep_oct_counter[12] ),
    .A(_03994_),
    .Y(_03995_),
    .D(_00118_));
 sg13g2_nor2b_1 _11830_ (.A(_03992_),
    .B_N(_03982_),
    .Y(_03996_));
 sg13g2_nor2b_1 _11831_ (.A(_03995_),
    .B_N(_03996_),
    .Y(_03997_));
 sg13g2_nand3_1 _11832_ (.B(_03946_),
    .C(_03988_),
    .A(_03987_),
    .Y(_03998_));
 sg13g2_o21ai_1 _11833_ (.B1(_03998_),
    .Y(_03999_),
    .A1(_03952_),
    .A2(_03988_));
 sg13g2_nand4_1 _11834_ (.B(_03978_),
    .C(_03961_),
    .A(_03971_),
    .Y(_04000_),
    .D(_03999_));
 sg13g2_nor2b_1 _11835_ (.A(_03959_),
    .B_N(_04000_),
    .Y(_04001_));
 sg13g2_nand3b_1 _11836_ (.B(_03952_),
    .C(\synth.voice.sweep_oct_counter[9] ),
    .Y(_04002_),
    .A_N(\synth.voice.sweep_oct_counter[10] ));
 sg13g2_inv_1 _11837_ (.Y(_04003_),
    .A(\synth.voice.sweep_oct_counter[9] ));
 sg13g2_nand2_1 _11838_ (.Y(_04004_),
    .A(_03947_),
    .B(_04003_));
 sg13g2_a21oi_1 _11839_ (.A1(_04002_),
    .A2(_04004_),
    .Y(_04005_),
    .B1(_03978_));
 sg13g2_nand2_1 _11840_ (.Y(_04006_),
    .A(_03990_),
    .B(_04005_));
 sg13g2_inv_1 _11841_ (.Y(_04007_),
    .A(_03945_));
 sg13g2_a21oi_1 _11842_ (.A1(_04001_),
    .A2(_04006_),
    .Y(_04008_),
    .B1(_04007_));
 sg13g2_o21ai_1 _11843_ (.B1(_04008_),
    .Y(_04009_),
    .A1(_03993_),
    .A2(_03997_));
 sg13g2_o21ai_1 _11844_ (.B1(_04009_),
    .Y(_04010_),
    .A1(_03945_),
    .A2(_03981_));
 sg13g2_nand3_1 _11845_ (.B(_03944_),
    .C(_04010_),
    .A(_03943_),
    .Y(_04011_));
 sg13g2_buf_2 _11846_ (.A(\synth.controller.rx_buffer[14] ),
    .X(_04012_));
 sg13g2_nand2_2 _11847_ (.Y(_04013_),
    .A(_04011_),
    .B(_04012_));
 sg13g2_inv_1 _11848_ (.Y(_04014_),
    .A(\synth.controller.rx_buffer_valid ));
 sg13g2_nor3_1 _11849_ (.A(\synth.controller.rx_sbs[0] ),
    .B(_03382_),
    .C(_04014_),
    .Y(_04015_));
 sg13g2_buf_2 _11850_ (.A(_04015_),
    .X(_04016_));
 sg13g2_nor3_1 _11851_ (.A(net330),
    .B(_03727_),
    .C(net332),
    .Y(_04017_));
 sg13g2_nand3_1 _11852_ (.B(_04016_),
    .C(_04017_),
    .A(_04013_),
    .Y(_04018_));
 sg13g2_buf_1 _11853_ (.A(_04018_),
    .X(_04019_));
 sg13g2_inv_1 _11854_ (.Y(_04020_),
    .A(_03596_));
 sg13g2_nor2_1 _11855_ (.A(_04020_),
    .B(_03602_),
    .Y(_04021_));
 sg13g2_inv_1 _11856_ (.Y(_04022_),
    .A(_03604_));
 sg13g2_nor2_1 _11857_ (.A(_04022_),
    .B(_03606_),
    .Y(_04023_));
 sg13g2_inv_1 _11858_ (.Y(_04024_),
    .A(\synth.controller.read_index_reg[2] ));
 sg13g2_nor2_1 _11859_ (.A(_04024_),
    .B(_03589_),
    .Y(_04025_));
 sg13g2_inv_1 _11860_ (.Y(_04026_),
    .A(_04025_));
 sg13g2_inv_1 _11861_ (.Y(_04027_),
    .A(_03591_));
 sg13g2_nor2_1 _11862_ (.A(_04027_),
    .B(_03594_),
    .Y(_04028_));
 sg13g2_inv_1 _11863_ (.Y(_04029_),
    .A(_04028_));
 sg13g2_nor2_1 _11864_ (.A(_04026_),
    .B(_04029_),
    .Y(_04030_));
 sg13g2_a21oi_1 _11865_ (.A1(_04021_),
    .A2(_04023_),
    .Y(_04031_),
    .B1(_04030_));
 sg13g2_buf_2 _11866_ (.A(_04031_),
    .X(_04032_));
 sg13g2_nand2_1 _11867_ (.Y(_04033_),
    .A(_04019_),
    .B(_04032_));
 sg13g2_buf_1 _11868_ (.A(_04033_),
    .X(_04034_));
 sg13g2_inv_1 _11869_ (.Y(_04035_),
    .A(\synth.voice.genblk4[6].next_state_scan[4] ));
 sg13g2_buf_1 _11870_ (.A(_04032_),
    .X(_04036_));
 sg13g2_o21ai_1 _11871_ (.B1(_03845_),
    .Y(_04037_),
    .A1(_03854_),
    .A2(_03859_));
 sg13g2_xnor2_1 _11872_ (.Y(_04038_),
    .A(_03832_),
    .B(_04037_));
 sg13g2_buf_1 _11873_ (.A(_04012_),
    .X(_04039_));
 sg13g2_nor2_1 _11874_ (.A(net373),
    .B(_03806_),
    .Y(_04040_));
 sg13g2_a21oi_2 _11875_ (.B1(_04040_),
    .Y(_04041_),
    .A2(net373),
    .A1(_04038_));
 sg13g2_buf_1 _11876_ (.A(_04032_),
    .X(_04042_));
 sg13g2_nand2b_1 _11877_ (.Y(_04043_),
    .B(net157),
    .A_N(_04041_));
 sg13g2_o21ai_1 _11878_ (.B1(_04043_),
    .Y(_04044_),
    .A1(_04035_),
    .A2(net158));
 sg13g2_nand2_1 _11879_ (.Y(_04045_),
    .A(net30),
    .B(_04044_));
 sg13g2_buf_1 _11880_ (.A(_04019_),
    .X(_04046_));
 sg13g2_buf_1 _11881_ (.A(net157),
    .X(_04047_));
 sg13g2_nand3_1 _11882_ (.B(_03818_),
    .C(net141),
    .A(net37),
    .Y(_04048_));
 sg13g2_nand2_1 _11883_ (.Y(_01099_),
    .A(_04045_),
    .B(_04048_));
 sg13g2_inv_1 _11884_ (.Y(_04049_),
    .A(\synth.voice.genblk4[6].next_state_scan[5] ));
 sg13g2_xnor2_1 _11885_ (.Y(_04050_),
    .A(_03803_),
    .B(_03856_));
 sg13g2_nand2_1 _11886_ (.Y(_04051_),
    .A(_04050_),
    .B(_03853_));
 sg13g2_nor2b_1 _11887_ (.A(_03832_),
    .B_N(_03852_),
    .Y(_04052_));
 sg13g2_inv_1 _11888_ (.Y(_04053_),
    .A(_04052_));
 sg13g2_nor2_1 _11889_ (.A(_04051_),
    .B(_04053_),
    .Y(_04054_));
 sg13g2_nand2_1 _11890_ (.Y(_04055_),
    .A(_04054_),
    .B(_03813_));
 sg13g2_nand2_1 _11891_ (.Y(_04056_),
    .A(_03858_),
    .B(_03853_));
 sg13g2_nand2b_1 _11892_ (.Y(_04057_),
    .B(_04056_),
    .A_N(_03844_));
 sg13g2_nand2b_1 _11893_ (.Y(_04058_),
    .B(_03831_),
    .A_N(_03843_));
 sg13g2_a21oi_1 _11894_ (.A1(_04057_),
    .A2(_04052_),
    .Y(_04059_),
    .B1(_04058_));
 sg13g2_nand2_1 _11895_ (.Y(_04060_),
    .A(_04055_),
    .B(_04059_));
 sg13g2_xnor2_1 _11896_ (.Y(_04061_),
    .A(_03841_),
    .B(_04060_));
 sg13g2_inv_1 _11897_ (.Y(_04062_),
    .A(\synth.controller.reg_wdata[5] ));
 sg13g2_nor2_1 _11898_ (.A(_04012_),
    .B(_04062_),
    .Y(_04063_));
 sg13g2_a21oi_2 _11899_ (.B1(_04063_),
    .Y(_04064_),
    .A2(_04039_),
    .A1(_04061_));
 sg13g2_nand2b_1 _11900_ (.Y(_04065_),
    .B(net157),
    .A_N(_04064_));
 sg13g2_o21ai_1 _11901_ (.B1(_04065_),
    .Y(_04066_),
    .A1(_04049_),
    .A2(net158));
 sg13g2_nand2_1 _11902_ (.Y(_04067_),
    .A(net30),
    .B(_04066_));
 sg13g2_nand3_1 _11903_ (.B(\synth.voice.genblk4[6].next_state_scan[3] ),
    .C(net141),
    .A(net37),
    .Y(_04068_));
 sg13g2_nand2_1 _11904_ (.Y(_01100_),
    .A(_04067_),
    .B(_04068_));
 sg13g2_inv_1 _11905_ (.Y(_04069_),
    .A(\synth.voice.genblk4[6].next_state_scan[6] ));
 sg13g2_nand2_1 _11906_ (.Y(_04070_),
    .A(_03862_),
    .B(_03872_));
 sg13g2_nand3_1 _11907_ (.B(_03861_),
    .C(_03871_),
    .A(_03849_),
    .Y(_04071_));
 sg13g2_nand3_1 _11908_ (.B(_04071_),
    .C(_04012_),
    .A(_04070_),
    .Y(_04072_));
 sg13g2_buf_1 _11909_ (.A(_04072_),
    .X(_04073_));
 sg13g2_inv_1 _11910_ (.Y(_04074_),
    .A(_04012_));
 sg13g2_nand2_2 _11911_ (.Y(_04075_),
    .A(_03947_),
    .B(net372));
 sg13g2_nand3_1 _11912_ (.B(net157),
    .C(_04075_),
    .A(_04073_),
    .Y(_04076_));
 sg13g2_o21ai_1 _11913_ (.B1(_04076_),
    .Y(_04077_),
    .A1(_04069_),
    .A2(net158));
 sg13g2_nand2_1 _11914_ (.Y(_04078_),
    .A(net30),
    .B(_04077_));
 sg13g2_nand3_1 _11915_ (.B(\synth.voice.genblk4[6].next_state_scan[4] ),
    .C(net141),
    .A(net37),
    .Y(_04079_));
 sg13g2_nand2_1 _11916_ (.Y(_01101_),
    .A(_04078_),
    .B(_04079_));
 sg13g2_nand3_1 _11917_ (.B(_03840_),
    .C(_03871_),
    .A(_03838_),
    .Y(_04080_));
 sg13g2_buf_1 _11918_ (.A(_04080_),
    .X(_04081_));
 sg13g2_inv_1 _11919_ (.Y(_04082_),
    .A(_04081_));
 sg13g2_nand2_1 _11920_ (.Y(_04083_),
    .A(_03870_),
    .B(_03930_));
 sg13g2_o21ai_1 _11921_ (.B1(_04083_),
    .Y(_04084_),
    .A1(_03872_),
    .A2(_03840_));
 sg13g2_a21oi_1 _11922_ (.A1(_04060_),
    .A2(_04082_),
    .Y(_04085_),
    .B1(_04084_));
 sg13g2_xnor2_1 _11923_ (.Y(_04086_),
    .A(_03869_),
    .B(_04085_));
 sg13g2_buf_1 _11924_ (.A(_04039_),
    .X(_04087_));
 sg13g2_nand2_2 _11925_ (.Y(_04088_),
    .A(_04086_),
    .B(_04087_));
 sg13g2_nand2_2 _11926_ (.Y(_04089_),
    .A(_03978_),
    .B(net372));
 sg13g2_nand3_1 _11927_ (.B(net157),
    .C(_04089_),
    .A(_04088_),
    .Y(_04090_));
 sg13g2_inv_1 _11928_ (.Y(_04091_),
    .A(_04032_));
 sg13g2_buf_1 _11929_ (.A(_04091_),
    .X(_04092_));
 sg13g2_nand2_1 _11930_ (.Y(_04093_),
    .A(net140),
    .B(\synth.voice.genblk4[6].next_state_scan[7] ));
 sg13g2_nand2_1 _11931_ (.Y(_04094_),
    .A(_04090_),
    .B(_04093_));
 sg13g2_nand2_1 _11932_ (.Y(_04095_),
    .A(net30),
    .B(_04094_));
 sg13g2_nand3_1 _11933_ (.B(\synth.voice.genblk4[6].next_state_scan[5] ),
    .C(net141),
    .A(net37),
    .Y(_04096_));
 sg13g2_nand2_1 _11934_ (.Y(_01102_),
    .A(_04095_),
    .B(_04096_));
 sg13g2_a21oi_1 _11935_ (.A1(_03862_),
    .A2(_03873_),
    .Y(_04097_),
    .B1(_03936_));
 sg13g2_xnor2_1 _11936_ (.Y(_04098_),
    .A(_03886_),
    .B(_04097_));
 sg13g2_nand2_1 _11937_ (.Y(_04099_),
    .A(_04098_),
    .B(net373));
 sg13g2_nand2_1 _11938_ (.Y(_04100_),
    .A(_03960_),
    .B(net372));
 sg13g2_nand3_1 _11939_ (.B(_04042_),
    .C(_04100_),
    .A(_04099_),
    .Y(_04101_));
 sg13g2_nand2_1 _11940_ (.Y(_04102_),
    .A(net140),
    .B(\synth.voice.genblk4[6].next_state_scan[8] ));
 sg13g2_nand2_1 _11941_ (.Y(_04103_),
    .A(_04101_),
    .B(_04102_));
 sg13g2_nand2_1 _11942_ (.Y(_04104_),
    .A(net30),
    .B(_04103_));
 sg13g2_nand3_1 _11943_ (.B(\synth.voice.genblk4[6].next_state_scan[6] ),
    .C(net141),
    .A(net37),
    .Y(_04105_));
 sg13g2_nand2_1 _11944_ (.Y(_01103_),
    .A(_04104_),
    .B(_04105_));
 sg13g2_nor2_1 _11945_ (.A(_03886_),
    .B(_03869_),
    .Y(_04106_));
 sg13g2_inv_1 _11946_ (.Y(_04107_),
    .A(_04106_));
 sg13g2_nor2_1 _11947_ (.A(_04107_),
    .B(_04081_),
    .Y(_04108_));
 sg13g2_nand2b_1 _11948_ (.Y(_04109_),
    .B(_04108_),
    .A_N(_04059_));
 sg13g2_nand3_1 _11949_ (.B(_03813_),
    .C(_04108_),
    .A(_04054_),
    .Y(_04110_));
 sg13g2_a21oi_1 _11950_ (.A1(_03867_),
    .A2(_03889_),
    .Y(_04111_),
    .B1(_03884_));
 sg13g2_nor2_1 _11951_ (.A(_03933_),
    .B(_04111_),
    .Y(_04112_));
 sg13g2_a21oi_1 _11952_ (.A1(_04084_),
    .A2(_04106_),
    .Y(_04113_),
    .B1(_04112_));
 sg13g2_nand3_1 _11953_ (.B(_04110_),
    .C(_04113_),
    .A(_04109_),
    .Y(_04114_));
 sg13g2_nand2_1 _11954_ (.Y(_04115_),
    .A(_04114_),
    .B(_03880_));
 sg13g2_nand4_1 _11955_ (.B(_04110_),
    .C(_03879_),
    .A(_04109_),
    .Y(_04116_),
    .D(_04113_));
 sg13g2_nand3_1 _11956_ (.B(_04116_),
    .C(net373),
    .A(_04115_),
    .Y(_04117_));
 sg13g2_nand2_1 _11957_ (.Y(_04118_),
    .A(_04007_),
    .B(net372));
 sg13g2_nand3_1 _11958_ (.B(_04042_),
    .C(_04118_),
    .A(_04117_),
    .Y(_04119_));
 sg13g2_nand2_1 _11959_ (.Y(_04120_),
    .A(net140),
    .B(\synth.voice.genblk4[6].next_state_scan[9] ));
 sg13g2_nand2_1 _11960_ (.Y(_04121_),
    .A(_04119_),
    .B(_04120_));
 sg13g2_nand2_1 _11961_ (.Y(_04122_),
    .A(_04034_),
    .B(_04121_));
 sg13g2_nand3_1 _11962_ (.B(\synth.voice.genblk4[6].next_state_scan[7] ),
    .C(_04047_),
    .A(_04046_),
    .Y(_04123_));
 sg13g2_nand2_1 _11963_ (.Y(_01104_),
    .A(_04122_),
    .B(_04123_));
 sg13g2_nand2b_1 _11964_ (.Y(_04124_),
    .B(_03862_),
    .A_N(_03888_));
 sg13g2_nand2_1 _11965_ (.Y(_04125_),
    .A(_04124_),
    .B(_03939_));
 sg13g2_xnor2_1 _11966_ (.Y(_04126_),
    .A(_03914_),
    .B(_04125_));
 sg13g2_nand2_1 _11967_ (.Y(_04127_),
    .A(_04126_),
    .B(net373));
 sg13g2_nand2_1 _11968_ (.Y(_04128_),
    .A(_03933_),
    .B(net372));
 sg13g2_nand3_1 _11969_ (.B(_04032_),
    .C(_04128_),
    .A(_04127_),
    .Y(_04129_));
 sg13g2_nand2_1 _11970_ (.Y(_04130_),
    .A(net140),
    .B(\synth.voice.genblk4[6].next_state_scan[10] ));
 sg13g2_nand2_1 _11971_ (.Y(_04131_),
    .A(_04129_),
    .B(_04130_));
 sg13g2_nand2_1 _11972_ (.Y(_04132_),
    .A(net30),
    .B(_04131_));
 sg13g2_nand3_1 _11973_ (.B(\synth.voice.genblk4[6].next_state_scan[8] ),
    .C(net141),
    .A(net37),
    .Y(_04133_));
 sg13g2_nand2_1 _11974_ (.Y(_01105_),
    .A(_04132_),
    .B(_04133_));
 sg13g2_nor2_1 _11975_ (.A(_03880_),
    .B(_03915_),
    .Y(_04134_));
 sg13g2_nor2b_1 _11976_ (.A(_04107_),
    .B_N(_04134_),
    .Y(_04135_));
 sg13g2_nand3_1 _11977_ (.B(_04052_),
    .C(_04135_),
    .A(_04082_),
    .Y(_04136_));
 sg13g2_inv_1 _11978_ (.Y(_04137_),
    .A(_04057_));
 sg13g2_o21ai_1 _11979_ (.B1(_04137_),
    .Y(_04138_),
    .A1(_03814_),
    .A2(_04051_));
 sg13g2_nand2b_1 _11980_ (.Y(_04139_),
    .B(_04138_),
    .A_N(_04136_));
 sg13g2_a21oi_1 _11981_ (.A1(net329),
    .A2(_03878_),
    .Y(_04140_),
    .B1(_03913_));
 sg13g2_nor2_1 _11982_ (.A(_03933_),
    .B(_04140_),
    .Y(_04141_));
 sg13g2_a21oi_1 _11983_ (.A1(_04112_),
    .A2(_04134_),
    .Y(_04142_),
    .B1(_04141_));
 sg13g2_nor2b_1 _11984_ (.A(_04081_),
    .B_N(_04058_),
    .Y(_04143_));
 sg13g2_o21ai_1 _11985_ (.B1(_04135_),
    .Y(_04144_),
    .A1(_04084_),
    .A2(_04143_));
 sg13g2_nand3_1 _11986_ (.B(_04142_),
    .C(_04144_),
    .A(_04139_),
    .Y(_04145_));
 sg13g2_nand2_1 _11987_ (.Y(_04146_),
    .A(_04145_),
    .B(_03925_));
 sg13g2_nand4_1 _11988_ (.B(_04144_),
    .C(_03924_),
    .A(_04139_),
    .Y(_04147_),
    .D(_04142_));
 sg13g2_nand3_1 _11989_ (.B(_04147_),
    .C(net373),
    .A(_04146_),
    .Y(_04148_));
 sg13g2_inv_1 _11990_ (.Y(_04149_),
    .A(\synth.controller.reg_waddr[3] ));
 sg13g2_nand2_1 _11991_ (.Y(_04150_),
    .A(net372),
    .B(_04149_));
 sg13g2_nand3_1 _11992_ (.B(_04032_),
    .C(_04150_),
    .A(_04148_),
    .Y(_04151_));
 sg13g2_nand2_1 _11993_ (.Y(_04152_),
    .A(net140),
    .B(\synth.voice.genblk4[6].next_state_scan[11] ));
 sg13g2_nand2_1 _11994_ (.Y(_04153_),
    .A(_04151_),
    .B(_04152_));
 sg13g2_nand2_1 _11995_ (.Y(_04154_),
    .A(net30),
    .B(_04153_));
 sg13g2_nand3_1 _11996_ (.B(\synth.voice.genblk4[6].next_state_scan[9] ),
    .C(net141),
    .A(net37),
    .Y(_04155_));
 sg13g2_nand2_1 _11997_ (.Y(_01106_),
    .A(_04154_),
    .B(_04155_));
 sg13g2_nand2_1 _11998_ (.Y(_04156_),
    .A(_03848_),
    .B(_03873_));
 sg13g2_nand2b_1 _11999_ (.Y(_04157_),
    .B(_04156_),
    .A_N(_03936_));
 sg13g2_nand2_1 _12000_ (.Y(_04158_),
    .A(_03926_),
    .B(_03887_));
 sg13g2_inv_1 _12001_ (.Y(_04159_),
    .A(_04158_));
 sg13g2_a21o_1 _12002_ (.A2(_03938_),
    .A1(_03926_),
    .B1(_03934_),
    .X(_04160_));
 sg13g2_a21oi_1 _12003_ (.A1(_04157_),
    .A2(_04159_),
    .Y(_04161_),
    .B1(_04160_));
 sg13g2_nand3_1 _12004_ (.B(_03873_),
    .C(_04159_),
    .A(_03842_),
    .Y(_04162_));
 sg13g2_nand2b_1 _12005_ (.Y(_04163_),
    .B(_04037_),
    .A_N(_04162_));
 sg13g2_a21oi_1 _12006_ (.A1(_04161_),
    .A2(_04163_),
    .Y(_04164_),
    .B1(_03908_));
 sg13g2_nand3_1 _12007_ (.B(_03908_),
    .C(_04163_),
    .A(_04161_),
    .Y(_04165_));
 sg13g2_nand3b_1 _12008_ (.B(net373),
    .C(_04165_),
    .Y(_04166_),
    .A_N(_04164_));
 sg13g2_buf_1 _12009_ (.A(_04166_),
    .X(_04167_));
 sg13g2_inv_1 _12010_ (.Y(_04168_),
    .A(\synth.controller.rx_buffer[12] ));
 sg13g2_nand2_2 _12011_ (.Y(_04169_),
    .A(net372),
    .B(_04168_));
 sg13g2_nand3_1 _12012_ (.B(_04032_),
    .C(_04169_),
    .A(_04167_),
    .Y(_04170_));
 sg13g2_nand2_1 _12013_ (.Y(_04171_),
    .A(net140),
    .B(\synth.voice.genblk4[6].next_state_scan[12] ));
 sg13g2_nand2_1 _12014_ (.Y(_04172_),
    .A(_04170_),
    .B(_04171_));
 sg13g2_nand2_1 _12015_ (.Y(_04173_),
    .A(_04034_),
    .B(_04172_));
 sg13g2_nand3_1 _12016_ (.B(\synth.voice.genblk4[6].next_state_scan[10] ),
    .C(_04047_),
    .A(_04046_),
    .Y(_04174_));
 sg13g2_nand2_1 _12017_ (.Y(_01107_),
    .A(_04173_),
    .B(_04174_));
 sg13g2_nor2_1 _12018_ (.A(_03901_),
    .B(_03905_),
    .Y(_04175_));
 sg13g2_nand3_1 _12019_ (.B(_04175_),
    .C(_03923_),
    .A(_04140_),
    .Y(_04176_));
 sg13g2_nor2_1 _12020_ (.A(_03933_),
    .B(_03906_),
    .Y(_04177_));
 sg13g2_nand3_1 _12021_ (.B(_03908_),
    .C(_03924_),
    .A(_04134_),
    .Y(_04178_));
 sg13g2_nor2_1 _12022_ (.A(_04178_),
    .B(_04113_),
    .Y(_04179_));
 sg13g2_a21oi_1 _12023_ (.A1(_04176_),
    .A2(_04177_),
    .Y(_04180_),
    .B1(_04179_));
 sg13g2_nor3_1 _12024_ (.A(_04107_),
    .B(_04178_),
    .C(_04081_),
    .Y(_04181_));
 sg13g2_nand2_1 _12025_ (.Y(_04182_),
    .A(_04060_),
    .B(_04181_));
 sg13g2_nand2_1 _12026_ (.Y(_04183_),
    .A(_04180_),
    .B(_04182_));
 sg13g2_nand2_1 _12027_ (.Y(_04184_),
    .A(_04183_),
    .B(_03898_));
 sg13g2_nand3_1 _12028_ (.B(_04182_),
    .C(_03897_),
    .A(_04180_),
    .Y(_04185_));
 sg13g2_nand3_1 _12029_ (.B(_04185_),
    .C(net373),
    .A(_04184_),
    .Y(_04186_));
 sg13g2_buf_1 _12030_ (.A(_04186_),
    .X(_04187_));
 sg13g2_inv_1 _12031_ (.Y(_04188_),
    .A(\synth.controller.rx_buffer[13] ));
 sg13g2_nand2_2 _12032_ (.Y(_04189_),
    .A(net372),
    .B(_04188_));
 sg13g2_nand3_1 _12033_ (.B(_04032_),
    .C(_04189_),
    .A(_04187_),
    .Y(_04190_));
 sg13g2_nand2_1 _12034_ (.Y(_04191_),
    .A(net140),
    .B(\synth.voice.genblk4[6].next_state_scan[13] ));
 sg13g2_nand2_1 _12035_ (.Y(_04192_),
    .A(_04190_),
    .B(_04191_));
 sg13g2_nand2_1 _12036_ (.Y(_04193_),
    .A(net30),
    .B(_04192_));
 sg13g2_nand3_1 _12037_ (.B(\synth.voice.genblk4[6].next_state_scan[11] ),
    .C(net141),
    .A(net37),
    .Y(_04194_));
 sg13g2_nand2_1 _12038_ (.Y(_01108_),
    .A(_04193_),
    .B(_04194_));
 sg13g2_inv_1 _12039_ (.Y(_04195_),
    .A(\synth.voice.genblk4[0].next_state_scan[8] ));
 sg13g2_inv_1 _12040_ (.Y(_04196_),
    .A(net193));
 sg13g2_nor2_1 _12041_ (.A(_04196_),
    .B(_01736_),
    .Y(_04197_));
 sg13g2_nor3_1 _12042_ (.A(_03481_),
    .B(_04197_),
    .C(_03583_),
    .Y(_04198_));
 sg13g2_buf_2 _12043_ (.A(_04198_),
    .X(_04199_));
 sg13g2_inv_1 _12044_ (.Y(_04200_),
    .A(net242));
 sg13g2_nand2_1 _12045_ (.Y(_04201_),
    .A(_04200_),
    .B(_03412_));
 sg13g2_nor2_2 _12046_ (.A(_01737_),
    .B(_04201_),
    .Y(_04202_));
 sg13g2_nand3_1 _12047_ (.B(net143),
    .C(_04202_),
    .A(_04199_),
    .Y(_04203_));
 sg13g2_buf_2 _12048_ (.A(_04203_),
    .X(_04204_));
 sg13g2_nand2_1 _12049_ (.Y(_04205_),
    .A(_04204_),
    .B(_03609_));
 sg13g2_buf_1 _12050_ (.A(_04205_),
    .X(_04206_));
 sg13g2_buf_8 _12051_ (.A(_04205_),
    .X(_04207_));
 sg13g2_inv_1 _12052_ (.Y(_04208_),
    .A(_00101_));
 sg13g2_inv_1 _12053_ (.Y(_04209_),
    .A(\synth.voice.genblk4[10].next_state_scan[13] ));
 sg13g2_buf_1 _12054_ (.A(net193),
    .X(_04210_));
 sg13g2_nor2_1 _12055_ (.A(_04209_),
    .B(net181),
    .Y(_04211_));
 sg13g2_buf_1 _12056_ (.A(_04211_),
    .X(_04212_));
 sg13g2_xnor2_1 _12057_ (.Y(_04213_),
    .A(_03657_),
    .B(_03652_));
 sg13g2_nor2_1 _12058_ (.A(_03663_),
    .B(_03671_),
    .Y(_04214_));
 sg13g2_nand2_1 _12059_ (.Y(_04215_),
    .A(_04213_),
    .B(_04214_));
 sg13g2_o21ai_1 _12060_ (.B1(_04215_),
    .Y(_04216_),
    .A1(_03652_),
    .A2(_03658_));
 sg13g2_nor2_1 _12061_ (.A(_03457_),
    .B(net159),
    .Y(_04217_));
 sg13g2_xor2_1 _12062_ (.B(_04217_),
    .A(_03632_),
    .X(_04218_));
 sg13g2_nand2_1 _12063_ (.Y(_04219_),
    .A(_04216_),
    .B(_04218_));
 sg13g2_nand2_1 _12064_ (.Y(_04220_),
    .A(_04217_),
    .B(_03632_));
 sg13g2_nand2_1 _12065_ (.Y(_04221_),
    .A(_04219_),
    .B(_04220_));
 sg13g2_xnor2_1 _12066_ (.Y(_04222_),
    .A(_03636_),
    .B(_03686_));
 sg13g2_nand2_1 _12067_ (.Y(_04223_),
    .A(_04221_),
    .B(_04222_));
 sg13g2_nand2_1 _12068_ (.Y(_04224_),
    .A(_03686_),
    .B(_03635_));
 sg13g2_nand2_1 _12069_ (.Y(_04225_),
    .A(_04223_),
    .B(_04224_));
 sg13g2_nand2_1 _12070_ (.Y(_04226_),
    .A(_04225_),
    .B(_03623_));
 sg13g2_nor2_1 _12071_ (.A(_03623_),
    .B(_04225_),
    .Y(_04227_));
 sg13g2_nor2_1 _12072_ (.A(net139),
    .B(_04227_),
    .Y(_04228_));
 sg13g2_a22oi_1 _12073_ (.Y(_04229_),
    .B1(_04226_),
    .B2(_04228_),
    .A2(net139),
    .A1(_04208_));
 sg13g2_buf_1 _12074_ (.A(_03611_),
    .X(_04230_));
 sg13g2_nand2_1 _12075_ (.Y(_04231_),
    .A(net180),
    .B(\synth.voice.genblk4[0].next_state_scan[10] ));
 sg13g2_o21ai_1 _12076_ (.B1(_04231_),
    .Y(_04232_),
    .A1(net182),
    .A2(_04229_));
 sg13g2_nand2_1 _12077_ (.Y(_04233_),
    .A(net43),
    .B(_04232_));
 sg13g2_o21ai_1 _12078_ (.B1(_04233_),
    .Y(_01109_),
    .A1(_04195_),
    .A2(net44));
 sg13g2_nor2_1 _12079_ (.A(_03727_),
    .B(_03755_),
    .Y(_04234_));
 sg13g2_nand3_1 _12080_ (.B(_04016_),
    .C(_04234_),
    .A(_04013_),
    .Y(_04235_));
 sg13g2_buf_1 _12081_ (.A(_04235_),
    .X(_04236_));
 sg13g2_nand2_1 _12082_ (.Y(_04237_),
    .A(_04236_),
    .B(net157));
 sg13g2_o21ai_1 _12083_ (.B1(_04043_),
    .Y(_04238_),
    .A1(net377),
    .A2(net158));
 sg13g2_nand2_1 _12084_ (.Y(_04239_),
    .A(_04237_),
    .B(_04238_));
 sg13g2_buf_1 _12085_ (.A(_04236_),
    .X(_04240_));
 sg13g2_nand3_1 _12086_ (.B(\synth.voice.genblk4[6].next_state_scan[12] ),
    .C(net158),
    .A(net36),
    .Y(_04241_));
 sg13g2_nand2_1 _12087_ (.Y(_01110_),
    .A(_04239_),
    .B(_04241_));
 sg13g2_o21ai_1 _12088_ (.B1(_04065_),
    .Y(_04242_),
    .A1(_03383_),
    .A2(net157));
 sg13g2_nand2_1 _12089_ (.Y(_04243_),
    .A(_04237_),
    .B(_04242_));
 sg13g2_nand3_1 _12090_ (.B(\synth.voice.genblk4[6].next_state_scan[13] ),
    .C(net158),
    .A(net36),
    .Y(_04244_));
 sg13g2_nand2_1 _12091_ (.Y(_01111_),
    .A(_04243_),
    .B(_04244_));
 sg13g2_nor2_1 _12092_ (.A(_03596_),
    .B(_03600_),
    .Y(_04245_));
 sg13g2_nor2_1 _12093_ (.A(_03601_),
    .B(_04245_),
    .Y(_04246_));
 sg13g2_inv_1 _12094_ (.Y(_04247_),
    .A(_04246_));
 sg13g2_inv_1 _12095_ (.Y(_04248_),
    .A(_04023_));
 sg13g2_nor2_1 _12096_ (.A(_03591_),
    .B(_03587_),
    .Y(_04249_));
 sg13g2_nor2_1 _12097_ (.A(_03593_),
    .B(_04249_),
    .Y(_04250_));
 sg13g2_nand2_1 _12098_ (.Y(_04251_),
    .A(_04025_),
    .B(_04250_));
 sg13g2_o21ai_1 _12099_ (.B1(_04251_),
    .Y(_04252_),
    .A1(_04247_),
    .A2(_04248_));
 sg13g2_buf_2 _12100_ (.A(_04252_),
    .X(_04253_));
 sg13g2_inv_1 _12101_ (.Y(_04254_),
    .A(_04253_));
 sg13g2_nand2_1 _12102_ (.Y(_04255_),
    .A(_04236_),
    .B(net179));
 sg13g2_buf_2 _12103_ (.A(_04255_),
    .X(_04256_));
 sg13g2_inv_1 _12104_ (.Y(_04257_),
    .A(\synth.voice.genblk4[7].next_state_scan[0] ));
 sg13g2_buf_1 _12105_ (.A(net179),
    .X(_04258_));
 sg13g2_nand3_1 _12106_ (.B(_04075_),
    .C(net179),
    .A(_04073_),
    .Y(_04259_));
 sg13g2_o21ai_1 _12107_ (.B1(_04259_),
    .Y(_04260_),
    .A1(_04257_),
    .A2(net156));
 sg13g2_nand2_1 _12108_ (.Y(_04261_),
    .A(_04256_),
    .B(_04260_));
 sg13g2_buf_1 _12109_ (.A(net156),
    .X(_04262_));
 sg13g2_nand3_1 _12110_ (.B(\synth.voice.mods[1][2] ),
    .C(net138),
    .A(net36),
    .Y(_04263_));
 sg13g2_nand2_1 _12111_ (.Y(_01112_),
    .A(_04261_),
    .B(_04263_));
 sg13g2_nand3_1 _12112_ (.B(_04089_),
    .C(net179),
    .A(_04088_),
    .Y(_04264_));
 sg13g2_buf_1 _12113_ (.A(_04253_),
    .X(_04265_));
 sg13g2_nand2_1 _12114_ (.Y(_04266_),
    .A(_04265_),
    .B(\synth.voice.genblk4[7].next_state_scan[1] ));
 sg13g2_nand2_1 _12115_ (.Y(_04267_),
    .A(_04264_),
    .B(_04266_));
 sg13g2_nand2_1 _12116_ (.Y(_04268_),
    .A(_04256_),
    .B(_04267_));
 sg13g2_nand3_1 _12117_ (.B(\synth.voice.mods[1][3] ),
    .C(_04262_),
    .A(_04240_),
    .Y(_04269_));
 sg13g2_nand2_1 _12118_ (.Y(_01113_),
    .A(_04268_),
    .B(_04269_));
 sg13g2_nand3_1 _12119_ (.B(_04100_),
    .C(net179),
    .A(_04099_),
    .Y(_04270_));
 sg13g2_nand2_1 _12120_ (.Y(_04271_),
    .A(net178),
    .B(_03757_));
 sg13g2_nand2_1 _12121_ (.Y(_04272_),
    .A(_04270_),
    .B(_04271_));
 sg13g2_nand2_1 _12122_ (.Y(_04273_),
    .A(_04256_),
    .B(_04272_));
 sg13g2_nand3_1 _12123_ (.B(\synth.voice.genblk4[7].next_state_scan[0] ),
    .C(net138),
    .A(net36),
    .Y(_04274_));
 sg13g2_nand2_1 _12124_ (.Y(_01114_),
    .A(_04273_),
    .B(_04274_));
 sg13g2_nand3_1 _12125_ (.B(_04118_),
    .C(net179),
    .A(_04117_),
    .Y(_04275_));
 sg13g2_nand2_1 _12126_ (.Y(_04276_),
    .A(_04265_),
    .B(_03917_));
 sg13g2_nand2_1 _12127_ (.Y(_04277_),
    .A(_04275_),
    .B(_04276_));
 sg13g2_nand2_1 _12128_ (.Y(_04278_),
    .A(_04256_),
    .B(_04277_));
 sg13g2_nand3_1 _12129_ (.B(\synth.voice.genblk4[7].next_state_scan[1] ),
    .C(net138),
    .A(_04240_),
    .Y(_04279_));
 sg13g2_nand2_1 _12130_ (.Y(_01115_),
    .A(_04278_),
    .B(_04279_));
 sg13g2_nand3_1 _12131_ (.B(_04128_),
    .C(_04254_),
    .A(_04127_),
    .Y(_04280_));
 sg13g2_nand2_1 _12132_ (.Y(_04281_),
    .A(net178),
    .B(_03902_));
 sg13g2_nand2_1 _12133_ (.Y(_04282_),
    .A(_04280_),
    .B(_04281_));
 sg13g2_nand2_1 _12134_ (.Y(_04283_),
    .A(_04256_),
    .B(_04282_));
 sg13g2_nand3_1 _12135_ (.B(_03757_),
    .C(net138),
    .A(net36),
    .Y(_04284_));
 sg13g2_nand2_1 _12136_ (.Y(_01116_),
    .A(_04283_),
    .B(_04284_));
 sg13g2_nand3_1 _12137_ (.B(_04150_),
    .C(_04254_),
    .A(_04148_),
    .Y(_04285_));
 sg13g2_nand2_1 _12138_ (.Y(_04286_),
    .A(net178),
    .B(\synth.voice.genblk4[7].next_state_scan[5] ));
 sg13g2_nand2_1 _12139_ (.Y(_04287_),
    .A(_04285_),
    .B(_04286_));
 sg13g2_nand2_1 _12140_ (.Y(_04288_),
    .A(_04256_),
    .B(_04287_));
 sg13g2_nand3_1 _12141_ (.B(_03917_),
    .C(net138),
    .A(net36),
    .Y(_04289_));
 sg13g2_nand2_1 _12142_ (.Y(_01117_),
    .A(_04288_),
    .B(_04289_));
 sg13g2_nand3_1 _12143_ (.B(_04169_),
    .C(net156),
    .A(_04167_),
    .Y(_04290_));
 sg13g2_nand2_1 _12144_ (.Y(_04291_),
    .A(net178),
    .B(_03817_));
 sg13g2_nand2_1 _12145_ (.Y(_04292_),
    .A(_04290_),
    .B(_04291_));
 sg13g2_nand2_1 _12146_ (.Y(_04293_),
    .A(_04256_),
    .B(_04292_));
 sg13g2_nand3_1 _12147_ (.B(_03902_),
    .C(_04262_),
    .A(net36),
    .Y(_04294_));
 sg13g2_nand2_1 _12148_ (.Y(_01118_),
    .A(_04293_),
    .B(_04294_));
 sg13g2_nand3_1 _12149_ (.B(_04189_),
    .C(net179),
    .A(_04187_),
    .Y(_04295_));
 sg13g2_nand2_1 _12150_ (.Y(_04296_),
    .A(net178),
    .B(\synth.voice.genblk4[7].next_state_scan[7] ));
 sg13g2_nand2_1 _12151_ (.Y(_04297_),
    .A(_04295_),
    .B(_04296_));
 sg13g2_nand2_1 _12152_ (.Y(_04298_),
    .A(_04256_),
    .B(_04297_));
 sg13g2_nand3_1 _12153_ (.B(\synth.voice.genblk4[7].next_state_scan[5] ),
    .C(net138),
    .A(net36),
    .Y(_04299_));
 sg13g2_nand2_1 _12154_ (.Y(_01119_),
    .A(_04298_),
    .B(_04299_));
 sg13g2_inv_1 _12155_ (.Y(_04300_),
    .A(\synth.voice.genblk4[0].next_state_scan[9] ));
 sg13g2_inv_1 _12156_ (.Y(_04301_),
    .A(_00099_));
 sg13g2_nand2_1 _12157_ (.Y(_04302_),
    .A(_04226_),
    .B(_03619_));
 sg13g2_nor2_1 _12158_ (.A(_03619_),
    .B(_04226_),
    .Y(_04303_));
 sg13g2_nor2_1 _12159_ (.A(net139),
    .B(_04303_),
    .Y(_04304_));
 sg13g2_a22oi_1 _12160_ (.Y(_04305_),
    .B1(_04302_),
    .B2(_04304_),
    .A2(net139),
    .A1(_04301_));
 sg13g2_nand2_1 _12161_ (.Y(_04306_),
    .A(net180),
    .B(\synth.voice.genblk4[0].next_state_scan[11] ));
 sg13g2_o21ai_1 _12162_ (.B1(_04306_),
    .Y(_04307_),
    .A1(net182),
    .A2(_04305_));
 sg13g2_nand2_1 _12163_ (.Y(_04308_),
    .A(net43),
    .B(_04307_));
 sg13g2_o21ai_1 _12164_ (.B1(_04308_),
    .Y(_01120_),
    .A1(_04300_),
    .A2(net44));
 sg13g2_nor3_1 _12165_ (.A(net400),
    .B(_03810_),
    .C(_00051_),
    .Y(_04309_));
 sg13g2_nand3_1 _12166_ (.B(_04016_),
    .C(_04309_),
    .A(_04013_),
    .Y(_04310_));
 sg13g2_buf_1 _12167_ (.A(_04310_),
    .X(_04311_));
 sg13g2_nand2_1 _12168_ (.Y(_04312_),
    .A(_04311_),
    .B(net179));
 sg13g2_buf_2 _12169_ (.A(_04312_),
    .X(_04313_));
 sg13g2_nand2_1 _12170_ (.Y(_04314_),
    .A(_04253_),
    .B(\synth.voice.genblk4[7].next_state_scan[8] ));
 sg13g2_o21ai_1 _12171_ (.B1(_04314_),
    .Y(_04315_),
    .A1(net178),
    .A2(_04041_));
 sg13g2_nand2_1 _12172_ (.Y(_04316_),
    .A(_04313_),
    .B(_04315_));
 sg13g2_buf_1 _12173_ (.A(_04311_),
    .X(_04317_));
 sg13g2_nand3_1 _12174_ (.B(_03817_),
    .C(net138),
    .A(net35),
    .Y(_04318_));
 sg13g2_nand2_1 _12175_ (.Y(_01121_),
    .A(_04316_),
    .B(_04318_));
 sg13g2_nand2_1 _12176_ (.Y(_04319_),
    .A(_04253_),
    .B(_03773_));
 sg13g2_o21ai_1 _12177_ (.B1(_04319_),
    .Y(_04320_),
    .A1(net178),
    .A2(_04064_));
 sg13g2_nand2_1 _12178_ (.Y(_04321_),
    .A(_04313_),
    .B(_04320_));
 sg13g2_nand3_1 _12179_ (.B(\synth.voice.genblk4[7].next_state_scan[7] ),
    .C(net138),
    .A(net35),
    .Y(_04322_));
 sg13g2_nand2_1 _12180_ (.Y(_01122_),
    .A(_04321_),
    .B(_04322_));
 sg13g2_inv_1 _12181_ (.Y(_04323_),
    .A(\synth.voice.genblk4[7].next_state_scan[10] ));
 sg13g2_o21ai_1 _12182_ (.B1(_04259_),
    .Y(_04324_),
    .A1(_04323_),
    .A2(net156));
 sg13g2_nand2_1 _12183_ (.Y(_04325_),
    .A(_04313_),
    .B(_04324_));
 sg13g2_nand3_1 _12184_ (.B(\synth.voice.genblk4[7].next_state_scan[8] ),
    .C(net156),
    .A(net35),
    .Y(_04326_));
 sg13g2_nand2_1 _12185_ (.Y(_01123_),
    .A(_04325_),
    .B(_04326_));
 sg13g2_nand2_1 _12186_ (.Y(_04327_),
    .A(net178),
    .B(\synth.voice.genblk4[7].next_state_scan[11] ));
 sg13g2_nand2_1 _12187_ (.Y(_04328_),
    .A(_04264_),
    .B(_04327_));
 sg13g2_nand2_1 _12188_ (.Y(_04329_),
    .A(_04313_),
    .B(_04328_));
 sg13g2_nand3_1 _12189_ (.B(_03773_),
    .C(net156),
    .A(net35),
    .Y(_04330_));
 sg13g2_nand2_1 _12190_ (.Y(_01124_),
    .A(_04329_),
    .B(_04330_));
 sg13g2_nand2_1 _12191_ (.Y(_04331_),
    .A(_04253_),
    .B(\synth.voice.genblk4[7].next_state_scan[12] ));
 sg13g2_nand2_1 _12192_ (.Y(_04332_),
    .A(_04270_),
    .B(_04331_));
 sg13g2_nand2_1 _12193_ (.Y(_04333_),
    .A(_04313_),
    .B(_04332_));
 sg13g2_nand3_1 _12194_ (.B(\synth.voice.genblk4[7].next_state_scan[10] ),
    .C(net156),
    .A(net35),
    .Y(_04334_));
 sg13g2_nand2_1 _12195_ (.Y(_01125_),
    .A(_04333_),
    .B(_04334_));
 sg13g2_nand2_1 _12196_ (.Y(_04335_),
    .A(_04253_),
    .B(\synth.voice.genblk4[7].next_state_scan[13] ));
 sg13g2_nand2_1 _12197_ (.Y(_04336_),
    .A(_04275_),
    .B(_04335_));
 sg13g2_nand2_1 _12198_ (.Y(_04337_),
    .A(_04313_),
    .B(_04336_));
 sg13g2_nand3_1 _12199_ (.B(\synth.voice.genblk4[7].next_state_scan[11] ),
    .C(_04258_),
    .A(net35),
    .Y(_04338_));
 sg13g2_nand2_1 _12200_ (.Y(_01126_),
    .A(_04337_),
    .B(_04338_));
 sg13g2_nand2_1 _12201_ (.Y(_04339_),
    .A(_04253_),
    .B(_03370_));
 sg13g2_nand2_1 _12202_ (.Y(_04340_),
    .A(_04280_),
    .B(_04339_));
 sg13g2_nand2_1 _12203_ (.Y(_04341_),
    .A(_04313_),
    .B(_04340_));
 sg13g2_nand3_1 _12204_ (.B(\synth.voice.genblk4[7].next_state_scan[12] ),
    .C(net156),
    .A(_04317_),
    .Y(_04342_));
 sg13g2_nand2_1 _12205_ (.Y(_01127_),
    .A(_04341_),
    .B(_04342_));
 sg13g2_nand2_1 _12206_ (.Y(_04343_),
    .A(_04253_),
    .B(net401));
 sg13g2_nand2_1 _12207_ (.Y(_04344_),
    .A(_04285_),
    .B(_04343_));
 sg13g2_nand2_1 _12208_ (.Y(_04345_),
    .A(_04313_),
    .B(_04344_));
 sg13g2_nand3_1 _12209_ (.B(\synth.voice.genblk4[7].next_state_scan[13] ),
    .C(_04258_),
    .A(_04317_),
    .Y(_04346_));
 sg13g2_nand2_1 _12210_ (.Y(_01128_),
    .A(_04345_),
    .B(_04346_));
 sg13g2_inv_1 _12211_ (.Y(_04347_),
    .A(\synth.controller.write_index_reg[3] ));
 sg13g2_nor2_1 _12212_ (.A(_03604_),
    .B(_04347_),
    .Y(_04348_));
 sg13g2_nand2_1 _12213_ (.Y(_04349_),
    .A(_03603_),
    .B(_04348_));
 sg13g2_nand2_1 _12214_ (.Y(_04350_),
    .A(_04024_),
    .B(\synth.controller.read_index_reg[3] ));
 sg13g2_inv_1 _12215_ (.Y(_04351_),
    .A(_04350_));
 sg13g2_nand2_1 _12216_ (.Y(_04352_),
    .A(_03595_),
    .B(_04351_));
 sg13g2_nand2_1 _12217_ (.Y(_04353_),
    .A(_04349_),
    .B(_04352_));
 sg13g2_buf_2 _12218_ (.A(_04353_),
    .X(_04354_));
 sg13g2_inv_1 _12219_ (.Y(_04355_),
    .A(_04354_));
 sg13g2_nand2_1 _12220_ (.Y(_04356_),
    .A(_04311_),
    .B(net177));
 sg13g2_nand3_1 _12221_ (.B(_04169_),
    .C(net177),
    .A(_04167_),
    .Y(_04357_));
 sg13g2_buf_1 _12222_ (.A(_04354_),
    .X(_04358_));
 sg13g2_nand2_1 _12223_ (.Y(_04359_),
    .A(net176),
    .B(\synth.voice.genblk4[8].next_state_scan[0] ));
 sg13g2_nand2_1 _12224_ (.Y(_04360_),
    .A(_04357_),
    .B(_04359_));
 sg13g2_nand2_1 _12225_ (.Y(_04361_),
    .A(_04356_),
    .B(_04360_));
 sg13g2_nand3_1 _12226_ (.B(\synth.voice.mods[2][8] ),
    .C(net177),
    .A(net35),
    .Y(_04362_));
 sg13g2_nand2_1 _12227_ (.Y(_01129_),
    .A(_04361_),
    .B(_04362_));
 sg13g2_nand3_1 _12228_ (.B(_04189_),
    .C(_04355_),
    .A(_04187_),
    .Y(_04363_));
 sg13g2_nand2_1 _12229_ (.Y(_04364_),
    .A(_04354_),
    .B(\synth.voice.genblk4[8].next_state_scan[1] ));
 sg13g2_nand2_1 _12230_ (.Y(_04365_),
    .A(_04363_),
    .B(_04364_));
 sg13g2_nand2_1 _12231_ (.Y(_04366_),
    .A(_04356_),
    .B(_04365_));
 sg13g2_nand3_1 _12232_ (.B(\synth.voice.mods[2][9] ),
    .C(net177),
    .A(net35),
    .Y(_04367_));
 sg13g2_nand2_1 _12233_ (.Y(_01130_),
    .A(_04366_),
    .B(_04367_));
 sg13g2_inv_1 _12234_ (.Y(_04368_),
    .A(\synth.voice.genblk4[0].next_state_scan[10] ));
 sg13g2_nor3_1 _12235_ (.A(_03680_),
    .B(_03619_),
    .C(_04226_),
    .Y(_04369_));
 sg13g2_nor2_1 _12236_ (.A(_03647_),
    .B(_04303_),
    .Y(_04370_));
 sg13g2_nor3_1 _12237_ (.A(net139),
    .B(_04369_),
    .C(_04370_),
    .Y(_04371_));
 sg13g2_a21oi_1 _12238_ (.A1(\synth.voice.genblk4[1].next_state_scan[3] ),
    .A2(net139),
    .Y(_04372_),
    .B1(_04371_));
 sg13g2_nand2_1 _12239_ (.Y(_04373_),
    .A(_04230_),
    .B(\synth.voice.genblk4[0].next_state_scan[12] ));
 sg13g2_o21ai_1 _12240_ (.B1(_04373_),
    .Y(_04374_),
    .A1(net182),
    .A2(_04372_));
 sg13g2_nand2_1 _12241_ (.Y(_04375_),
    .A(net43),
    .B(_04374_));
 sg13g2_o21ai_1 _12242_ (.B1(_04375_),
    .Y(_01131_),
    .A1(_04368_),
    .A2(net44));
 sg13g2_nand4_1 _12243_ (.B(_03412_),
    .C(net143),
    .A(_04199_),
    .Y(_04376_),
    .D(_04211_));
 sg13g2_buf_1 _12244_ (.A(_04376_),
    .X(_04377_));
 sg13g2_nand2_1 _12245_ (.Y(_04378_),
    .A(_04377_),
    .B(net177));
 sg13g2_buf_2 _12246_ (.A(_04378_),
    .X(_04379_));
 sg13g2_inv_1 _12247_ (.Y(_04380_),
    .A(\synth.voice.genblk4[1].next_state_scan[7] ));
 sg13g2_nand2_1 _12248_ (.Y(_04381_),
    .A(_04354_),
    .B(\synth.voice.genblk4[8].next_state_scan[2] ));
 sg13g2_o21ai_1 _12249_ (.B1(_04381_),
    .Y(_04382_),
    .A1(_04380_),
    .A2(net176));
 sg13g2_nand2_1 _12250_ (.Y(_04383_),
    .A(_04379_),
    .B(_04382_));
 sg13g2_nand3_1 _12251_ (.B(\synth.voice.genblk4[8].next_state_scan[0] ),
    .C(net177),
    .A(_04377_),
    .Y(_04384_));
 sg13g2_nand2_1 _12252_ (.Y(_01132_),
    .A(_04383_),
    .B(_04384_));
 sg13g2_mux2_1 _12253_ (.A0(\synth.voice.genblk4[8].next_state_scan[0] ),
    .A1(\synth.voice.genblk4[8].next_state_scan[3] ),
    .S(_04354_),
    .X(_04385_));
 sg13g2_nand2_1 _12254_ (.Y(_04386_),
    .A(_04379_),
    .B(_04385_));
 sg13g2_nand3_1 _12255_ (.B(\synth.voice.genblk4[8].next_state_scan[1] ),
    .C(net177),
    .A(_04377_),
    .Y(_04387_));
 sg13g2_nand2_1 _12256_ (.Y(_01133_),
    .A(_04386_),
    .B(_04387_));
 sg13g2_nor2b_1 _12257_ (.A(net176),
    .B_N(\synth.voice.genblk4[8].next_state_scan[1] ),
    .Y(_04388_));
 sg13g2_a21oi_1 _12258_ (.A1(\synth.voice.genblk4[8].next_state_scan[4] ),
    .A2(net176),
    .Y(_04389_),
    .B1(_04388_));
 sg13g2_nor2_1 _12259_ (.A(\synth.voice.genblk4[8].next_state_scan[2] ),
    .B(_04379_),
    .Y(_04390_));
 sg13g2_a21oi_1 _12260_ (.A1(_04379_),
    .A2(_04389_),
    .Y(_01134_),
    .B1(_04390_));
 sg13g2_inv_1 _12261_ (.Y(_04391_),
    .A(\synth.voice.genblk4[8].next_state_scan[5] ));
 sg13g2_nor2_1 _12262_ (.A(\synth.voice.genblk4[8].next_state_scan[2] ),
    .B(net176),
    .Y(_04392_));
 sg13g2_a21o_1 _12263_ (.A2(net176),
    .A1(_04391_),
    .B1(_04392_),
    .X(_04393_));
 sg13g2_nor2_1 _12264_ (.A(\synth.voice.genblk4[8].next_state_scan[3] ),
    .B(_04379_),
    .Y(_04394_));
 sg13g2_a21oi_1 _12265_ (.A1(_04379_),
    .A2(_04393_),
    .Y(_01135_),
    .B1(_04394_));
 sg13g2_mux2_1 _12266_ (.A0(\synth.voice.genblk4[8].next_state_scan[3] ),
    .A1(\synth.voice.genblk4[8].next_state_scan[6] ),
    .S(_04354_),
    .X(_04395_));
 sg13g2_nand2_1 _12267_ (.Y(_04396_),
    .A(_04379_),
    .B(_04395_));
 sg13g2_nand3_1 _12268_ (.B(\synth.voice.genblk4[8].next_state_scan[4] ),
    .C(net177),
    .A(_04377_),
    .Y(_04397_));
 sg13g2_nand2_1 _12269_ (.Y(_01136_),
    .A(_04396_),
    .B(_04397_));
 sg13g2_inv_1 _12270_ (.Y(_04398_),
    .A(_00058_));
 sg13g2_inv_1 _12271_ (.Y(_04399_),
    .A(\synth.voice.genblk4[10].next_state_scan[8] ));
 sg13g2_inv_1 _12272_ (.Y(_04400_),
    .A(\synth.voice.genblk4[9].next_state_scan[11] ));
 sg13g2_a22oi_1 _12273_ (.Y(_04401_),
    .B1(_04400_),
    .B2(_01772_),
    .A2(_04399_),
    .A1(_01730_));
 sg13g2_o21ai_1 _12274_ (.B1(_04401_),
    .Y(_04402_),
    .A1(_04398_),
    .A2(net255));
 sg13g2_buf_1 _12275_ (.A(_04402_),
    .X(_04403_));
 sg13g2_nor2b_1 _12276_ (.A(net255),
    .B_N(_00085_),
    .Y(_04404_));
 sg13g2_inv_1 _12277_ (.Y(_04405_),
    .A(\synth.voice.genblk4[10].next_state_scan[7] ));
 sg13g2_inv_1 _12278_ (.Y(_04406_),
    .A(\synth.voice.genblk4[9].next_state_scan[10] ));
 sg13g2_a22oi_1 _12279_ (.Y(_04407_),
    .B1(_04406_),
    .B2(_01772_),
    .A2(_04405_),
    .A1(_01730_));
 sg13g2_nand2b_1 _12280_ (.Y(_04408_),
    .B(_04407_),
    .A_N(_04404_));
 sg13g2_inv_2 _12281_ (.Y(_04409_),
    .A(_04408_));
 sg13g2_nand2b_1 _12282_ (.Y(_04410_),
    .B(_04409_),
    .A_N(_04403_));
 sg13g2_buf_2 _12283_ (.A(_04410_),
    .X(_04411_));
 sg13g2_buf_8 _12284_ (.A(_04411_),
    .X(_04412_));
 sg13g2_inv_1 _12285_ (.Y(_04413_),
    .A(_00092_));
 sg13g2_inv_1 _12286_ (.Y(_04414_),
    .A(\synth.voice.genblk4[10].next_state_scan[3] ));
 sg13g2_inv_1 _12287_ (.Y(_04415_),
    .A(\synth.voice.genblk4[9].next_state_scan[6] ));
 sg13g2_a22oi_1 _12288_ (.Y(_04416_),
    .B1(_04415_),
    .B2(_01772_),
    .A2(_04414_),
    .A1(_01730_));
 sg13g2_o21ai_1 _12289_ (.B1(_04416_),
    .Y(_04417_),
    .A1(_04413_),
    .A2(net255));
 sg13g2_buf_1 _12290_ (.A(_04417_),
    .X(_04418_));
 sg13g2_inv_1 _12291_ (.Y(_04419_),
    .A(_04418_));
 sg13g2_nand3_1 _12292_ (.B(_03616_),
    .C(_04419_),
    .A(net137),
    .Y(_04420_));
 sg13g2_buf_1 _12293_ (.A(_04418_),
    .X(_04421_));
 sg13g2_nand3_1 _12294_ (.B(_03645_),
    .C(net191),
    .A(net137),
    .Y(_04422_));
 sg13g2_inv_1 _12295_ (.Y(_04423_),
    .A(\synth.voice.genblk4[10].next_state_scan[4] ));
 sg13g2_inv_1 _12296_ (.Y(_04424_),
    .A(\synth.voice.genblk4[9].next_state_scan[7] ));
 sg13g2_nor2b_1 _12297_ (.A(net255),
    .B_N(_00094_),
    .Y(_04425_));
 sg13g2_a221oi_1 _12298_ (.B2(net299),
    .C1(_04425_),
    .B1(_04424_),
    .A1(_04423_),
    .Y(_04426_),
    .A2(net300));
 sg13g2_buf_2 _12299_ (.A(_04426_),
    .X(_04427_));
 sg13g2_and3_1 _12300_ (.X(_04428_),
    .A(_04420_),
    .B(_04422_),
    .C(_04427_));
 sg13g2_inv_1 _12301_ (.Y(_04429_),
    .A(net137));
 sg13g2_nor2_1 _12302_ (.A(_00095_),
    .B(net191),
    .Y(_04430_));
 sg13g2_a21oi_1 _12303_ (.A1(_03696_),
    .A2(net191),
    .Y(_04431_),
    .B1(_04430_));
 sg13g2_inv_1 _12304_ (.Y(_04432_),
    .A(_04427_));
 sg13g2_buf_1 _12305_ (.A(_04432_),
    .X(_04433_));
 sg13g2_o21ai_1 _12306_ (.B1(net155),
    .Y(_04434_),
    .A1(_04429_),
    .A2(_04431_));
 sg13g2_nor2b_1 _12307_ (.A(_04428_),
    .B_N(_04434_),
    .Y(_04435_));
 sg13g2_nand2b_1 _12308_ (.Y(_04436_),
    .B(_04408_),
    .A_N(_04403_));
 sg13g2_nand2_1 _12309_ (.Y(_04437_),
    .A(_04403_),
    .B(_04409_));
 sg13g2_buf_8 _12310_ (.A(_04437_),
    .X(_04438_));
 sg13g2_nand2_1 _12311_ (.Y(_04439_),
    .A(_04436_),
    .B(_04438_));
 sg13g2_buf_8 _12312_ (.A(_04439_),
    .X(_04440_));
 sg13g2_nand2b_1 _12313_ (.Y(_04441_),
    .B(net128),
    .A_N(_00097_));
 sg13g2_nand2_1 _12314_ (.Y(_04442_),
    .A(net154),
    .B(_00097_));
 sg13g2_nand2_1 _12315_ (.Y(_04443_),
    .A(_04441_),
    .B(_04442_));
 sg13g2_inv_1 _12316_ (.Y(_04444_),
    .A(_04443_));
 sg13g2_inv_1 _12317_ (.Y(_04445_),
    .A(\synth.voice.genblk4[10].next_state_scan[5] ));
 sg13g2_inv_1 _12318_ (.Y(_04446_),
    .A(\synth.voice.genblk4[9].next_state_scan[8] ));
 sg13g2_nor2b_1 _12319_ (.A(net255),
    .B_N(_00086_),
    .Y(_04447_));
 sg13g2_a221oi_1 _12320_ (.B2(net299),
    .C1(_04447_),
    .B1(_04446_),
    .A1(_04445_),
    .Y(_04448_),
    .A2(net300));
 sg13g2_buf_1 _12321_ (.A(_04448_),
    .X(_04449_));
 sg13g2_buf_1 _12322_ (.A(_04449_),
    .X(_04450_));
 sg13g2_nand2_1 _12323_ (.Y(_04451_),
    .A(_04444_),
    .B(net175));
 sg13g2_nand2b_1 _12324_ (.Y(_04452_),
    .B(net128),
    .A_N(_00090_));
 sg13g2_nand2_1 _12325_ (.Y(_04453_),
    .A(net154),
    .B(_00090_));
 sg13g2_nand2_1 _12326_ (.Y(_04454_),
    .A(_04452_),
    .B(_04453_));
 sg13g2_inv_1 _12327_ (.Y(_04455_),
    .A(_04454_));
 sg13g2_inv_1 _12328_ (.Y(_04456_),
    .A(_04449_));
 sg13g2_nand2_1 _12329_ (.Y(_04457_),
    .A(_04455_),
    .B(net174));
 sg13g2_inv_1 _12330_ (.Y(_04458_),
    .A(\synth.voice.genblk4[10].next_state_scan[6] ));
 sg13g2_inv_1 _12331_ (.Y(_04459_),
    .A(\synth.voice.genblk4[9].next_state_scan[9] ));
 sg13g2_nor2b_1 _12332_ (.A(net255),
    .B_N(_00088_),
    .Y(_04460_));
 sg13g2_a221oi_1 _12333_ (.B2(net299),
    .C1(_04460_),
    .B1(_04459_),
    .A1(_04458_),
    .Y(_04461_),
    .A2(net300));
 sg13g2_buf_1 _12334_ (.A(_04461_),
    .X(_04462_));
 sg13g2_nand3_1 _12335_ (.B(_04457_),
    .C(net190),
    .A(_04451_),
    .Y(_04463_));
 sg13g2_nand2b_1 _12336_ (.Y(_04464_),
    .B(net128),
    .A_N(_00089_));
 sg13g2_nand2_1 _12337_ (.Y(_04465_),
    .A(net154),
    .B(_00089_));
 sg13g2_nand2_1 _12338_ (.Y(_04466_),
    .A(_04464_),
    .B(_04465_));
 sg13g2_inv_1 _12339_ (.Y(_04467_),
    .A(_04466_));
 sg13g2_nand2_1 _12340_ (.Y(_04468_),
    .A(_04467_),
    .B(net175));
 sg13g2_nand2b_1 _12341_ (.Y(_04469_),
    .B(net128),
    .A_N(_00087_));
 sg13g2_nand2_1 _12342_ (.Y(_04470_),
    .A(net154),
    .B(_00087_));
 sg13g2_nand2_1 _12343_ (.Y(_04471_),
    .A(_04469_),
    .B(_04470_));
 sg13g2_inv_1 _12344_ (.Y(_04472_),
    .A(_04471_));
 sg13g2_nand2_1 _12345_ (.Y(_04473_),
    .A(_04472_),
    .B(net174));
 sg13g2_inv_2 _12346_ (.Y(_04474_),
    .A(net190));
 sg13g2_nand3_1 _12347_ (.B(_04473_),
    .C(net173),
    .A(_04468_),
    .Y(_04475_));
 sg13g2_nand2_1 _12348_ (.Y(_04476_),
    .A(_04463_),
    .B(_04475_));
 sg13g2_nand2b_1 _12349_ (.Y(_04477_),
    .B(_04476_),
    .A_N(_04435_));
 sg13g2_nand3_1 _12350_ (.B(_04475_),
    .C(_04435_),
    .A(_04463_),
    .Y(_04478_));
 sg13g2_nand2_1 _12351_ (.Y(_04479_),
    .A(_04477_),
    .B(_04478_));
 sg13g2_nand2_1 _12352_ (.Y(_04480_),
    .A(_04411_),
    .B(_03654_));
 sg13g2_inv_1 _12353_ (.Y(_04481_),
    .A(_00104_));
 sg13g2_nand3_1 _12354_ (.B(_04481_),
    .C(_04418_),
    .A(_04411_),
    .Y(_04482_));
 sg13g2_o21ai_1 _12355_ (.B1(_04482_),
    .Y(_04483_),
    .A1(_04421_),
    .A2(_04480_));
 sg13g2_inv_1 _12356_ (.Y(_04484_),
    .A(_00107_));
 sg13g2_nand3_1 _12357_ (.B(_04484_),
    .C(_04418_),
    .A(_04411_),
    .Y(_04485_));
 sg13g2_nor2_1 _12358_ (.A(_04432_),
    .B(_04485_),
    .Y(_04486_));
 sg13g2_a21oi_1 _12359_ (.A1(_04483_),
    .A2(_04433_),
    .Y(_04487_),
    .B1(_04486_));
 sg13g2_a21oi_1 _12360_ (.A1(_04403_),
    .A2(_04409_),
    .Y(_04488_),
    .B1(_03630_));
 sg13g2_a21oi_1 _12361_ (.A1(net128),
    .A2(_03630_),
    .Y(_04489_),
    .B1(_04488_));
 sg13g2_nand2_1 _12362_ (.Y(_04490_),
    .A(_04489_),
    .B(net174));
 sg13g2_inv_1 _12363_ (.Y(_04491_),
    .A(_00105_));
 sg13g2_nand2_1 _12364_ (.Y(_04492_),
    .A(_04440_),
    .B(_04491_));
 sg13g2_nand2_1 _12365_ (.Y(_04493_),
    .A(_04438_),
    .B(_00105_));
 sg13g2_nand3_1 _12366_ (.B(net175),
    .C(_04493_),
    .A(_04492_),
    .Y(_04494_));
 sg13g2_nand3_1 _12367_ (.B(_04494_),
    .C(net173),
    .A(_04490_),
    .Y(_04495_));
 sg13g2_nand2_1 _12368_ (.Y(_04496_),
    .A(_04440_),
    .B(_03660_));
 sg13g2_nand2_1 _12369_ (.Y(_04497_),
    .A(net154),
    .B(_00060_));
 sg13g2_nand3_1 _12370_ (.B(_04456_),
    .C(_04497_),
    .A(_04496_),
    .Y(_04498_));
 sg13g2_nand2_1 _12371_ (.Y(_04499_),
    .A(_04498_),
    .B(net190));
 sg13g2_nand3b_1 _12372_ (.B(_04495_),
    .C(_04499_),
    .Y(_04500_),
    .A_N(_04487_));
 sg13g2_buf_1 _12373_ (.A(_04500_),
    .X(_04501_));
 sg13g2_nand2_1 _12374_ (.Y(_04502_),
    .A(_04495_),
    .B(_04499_));
 sg13g2_nand2_1 _12375_ (.Y(_04503_),
    .A(_04502_),
    .B(_04487_));
 sg13g2_nand2_1 _12376_ (.Y(_04504_),
    .A(_04501_),
    .B(_04503_));
 sg13g2_nand3_1 _12377_ (.B(_04484_),
    .C(_04419_),
    .A(_04412_),
    .Y(_04505_));
 sg13g2_o21ai_1 _12378_ (.B1(_04505_),
    .Y(_04506_),
    .A1(_04419_),
    .A2(_04480_));
 sg13g2_nand3_1 _12379_ (.B(_04481_),
    .C(_04419_),
    .A(net137),
    .Y(_04507_));
 sg13g2_nand3_1 _12380_ (.B(_03633_),
    .C(_04421_),
    .A(_04412_),
    .Y(_04508_));
 sg13g2_a21oi_1 _12381_ (.A1(_04507_),
    .A2(_04508_),
    .Y(_04509_),
    .B1(_04427_));
 sg13g2_a21oi_2 _12382_ (.B1(_04509_),
    .Y(_04510_),
    .A2(_04427_),
    .A1(_04506_));
 sg13g2_nand2_1 _12383_ (.Y(_04511_),
    .A(_04492_),
    .B(_04493_));
 sg13g2_nand2_1 _12384_ (.Y(_04512_),
    .A(_04511_),
    .B(net174));
 sg13g2_nand2_1 _12385_ (.Y(_04513_),
    .A(_04496_),
    .B(_04497_));
 sg13g2_nand2_1 _12386_ (.Y(_04514_),
    .A(_04513_),
    .B(_04450_));
 sg13g2_nand2_1 _12387_ (.Y(_04515_),
    .A(_04512_),
    .B(_04514_));
 sg13g2_nand2_1 _12388_ (.Y(_04516_),
    .A(_04515_),
    .B(net190));
 sg13g2_nand2_1 _12389_ (.Y(_04517_),
    .A(_04489_),
    .B(_04450_));
 sg13g2_nand2_1 _12390_ (.Y(_04518_),
    .A(net128),
    .B(_04208_));
 sg13g2_nand2_1 _12391_ (.Y(_04519_),
    .A(net154),
    .B(_00101_));
 sg13g2_nand3_1 _12392_ (.B(net174),
    .C(_04519_),
    .A(_04518_),
    .Y(_04520_));
 sg13g2_nand3_1 _12393_ (.B(_04520_),
    .C(_04474_),
    .A(_04517_),
    .Y(_04521_));
 sg13g2_nand2_1 _12394_ (.Y(_04522_),
    .A(_04516_),
    .B(_04521_));
 sg13g2_xnor2_1 _12395_ (.Y(_04523_),
    .A(_04510_),
    .B(_04522_));
 sg13g2_nor2_1 _12396_ (.A(_04504_),
    .B(_04523_),
    .Y(_04524_));
 sg13g2_nand3_1 _12397_ (.B(_04514_),
    .C(net173),
    .A(_04512_),
    .Y(_04525_));
 sg13g2_nand2_1 _12398_ (.Y(_04526_),
    .A(_04506_),
    .B(net155));
 sg13g2_nand2_1 _12399_ (.Y(_04527_),
    .A(_04525_),
    .B(_04526_));
 sg13g2_nand2b_1 _12400_ (.Y(_04528_),
    .B(_04474_),
    .A_N(_04498_));
 sg13g2_nor2_1 _12401_ (.A(_04427_),
    .B(_04485_),
    .Y(_04529_));
 sg13g2_nor2b_1 _12402_ (.A(_04528_),
    .B_N(_04529_),
    .Y(_04530_));
 sg13g2_buf_1 _12403_ (.A(_04530_),
    .X(_04531_));
 sg13g2_nor2_1 _12404_ (.A(_04526_),
    .B(_04525_),
    .Y(_04532_));
 sg13g2_a21oi_2 _12405_ (.B1(_04532_),
    .Y(_04533_),
    .A2(_04531_),
    .A1(_04527_));
 sg13g2_inv_1 _12406_ (.Y(_04534_),
    .A(_04533_));
 sg13g2_nand2_1 _12407_ (.Y(_04535_),
    .A(_04524_),
    .B(_04534_));
 sg13g2_inv_1 _12408_ (.Y(_04536_),
    .A(_04501_));
 sg13g2_nand2_1 _12409_ (.Y(_04537_),
    .A(_04522_),
    .B(_04510_));
 sg13g2_nor2_1 _12410_ (.A(_04510_),
    .B(_04522_),
    .Y(_04538_));
 sg13g2_a21oi_1 _12411_ (.A1(_04536_),
    .A2(_04537_),
    .Y(_04539_),
    .B1(_04538_));
 sg13g2_nand2_1 _12412_ (.Y(_04540_),
    .A(_04535_),
    .B(_04539_));
 sg13g2_nand3_1 _12413_ (.B(_03620_),
    .C(_04419_),
    .A(net137),
    .Y(_04541_));
 sg13g2_nand3_1 _12414_ (.B(_03616_),
    .C(net191),
    .A(net137),
    .Y(_04542_));
 sg13g2_nand2_1 _12415_ (.Y(_04543_),
    .A(_04541_),
    .B(_04542_));
 sg13g2_a21oi_1 _12416_ (.A1(_04507_),
    .A2(_04508_),
    .Y(_04544_),
    .B1(net155));
 sg13g2_a21o_1 _12417_ (.A2(_04543_),
    .A1(net155),
    .B1(_04544_),
    .X(_04545_));
 sg13g2_buf_1 _12418_ (.A(_04545_),
    .X(_04546_));
 sg13g2_nand2_1 _12419_ (.Y(_04547_),
    .A(_04444_),
    .B(net174));
 sg13g2_nand2_1 _12420_ (.Y(_04548_),
    .A(net128),
    .B(_04301_));
 sg13g2_nand2_1 _12421_ (.Y(_04549_),
    .A(net154),
    .B(_00099_));
 sg13g2_nand3_1 _12422_ (.B(net175),
    .C(_04549_),
    .A(_04548_),
    .Y(_04550_));
 sg13g2_nand3_1 _12423_ (.B(net173),
    .C(_04550_),
    .A(_04547_),
    .Y(_04551_));
 sg13g2_nand3_1 _12424_ (.B(_04520_),
    .C(_04462_),
    .A(_04517_),
    .Y(_04552_));
 sg13g2_nand2_1 _12425_ (.Y(_04553_),
    .A(_04551_),
    .B(_04552_));
 sg13g2_xnor2_1 _12426_ (.Y(_04554_),
    .A(_04546_),
    .B(_04553_));
 sg13g2_nand2_1 _12427_ (.Y(_04555_),
    .A(_04483_),
    .B(_04427_));
 sg13g2_a21oi_1 _12428_ (.A1(_04411_),
    .A2(_03620_),
    .Y(_04556_),
    .B1(_04419_));
 sg13g2_a21oi_1 _12429_ (.A1(_04411_),
    .A2(_03633_),
    .Y(_04557_),
    .B1(_04418_));
 sg13g2_nor2_1 _12430_ (.A(_04556_),
    .B(_04557_),
    .Y(_04558_));
 sg13g2_nand2_1 _12431_ (.Y(_04559_),
    .A(_04558_),
    .B(_04433_));
 sg13g2_nand2_1 _12432_ (.Y(_04560_),
    .A(_04555_),
    .B(_04559_));
 sg13g2_nand3_1 _12433_ (.B(_04494_),
    .C(net190),
    .A(_04490_),
    .Y(_04561_));
 sg13g2_nand3_1 _12434_ (.B(net175),
    .C(_04519_),
    .A(_04518_),
    .Y(_04562_));
 sg13g2_nand3_1 _12435_ (.B(net174),
    .C(_04549_),
    .A(_04548_),
    .Y(_04563_));
 sg13g2_nand3_1 _12436_ (.B(_04563_),
    .C(net173),
    .A(_04562_),
    .Y(_04564_));
 sg13g2_nand2_1 _12437_ (.Y(_04565_),
    .A(_04561_),
    .B(_04564_));
 sg13g2_nand2b_1 _12438_ (.Y(_04566_),
    .B(_04565_),
    .A_N(_04560_));
 sg13g2_nand3_1 _12439_ (.B(_04564_),
    .C(_04560_),
    .A(_04561_),
    .Y(_04567_));
 sg13g2_nand2_1 _12440_ (.Y(_04568_),
    .A(_04566_),
    .B(_04567_));
 sg13g2_inv_1 _12441_ (.Y(_04569_),
    .A(_04568_));
 sg13g2_nand2_1 _12442_ (.Y(_04570_),
    .A(_04554_),
    .B(_04569_));
 sg13g2_nand2_1 _12443_ (.Y(_04571_),
    .A(net191),
    .B(_03676_));
 sg13g2_o21ai_1 _12444_ (.B1(_04571_),
    .Y(_04572_),
    .A1(_00096_),
    .A2(net191));
 sg13g2_nand2_1 _12445_ (.Y(_04573_),
    .A(_04572_),
    .B(net137));
 sg13g2_nor2_1 _12446_ (.A(net155),
    .B(_04543_),
    .Y(_04574_));
 sg13g2_a21oi_1 _12447_ (.A1(net155),
    .A2(_04573_),
    .Y(_04575_),
    .B1(_04574_));
 sg13g2_nand2_1 _12448_ (.Y(_04576_),
    .A(_04455_),
    .B(net175));
 sg13g2_nand2_1 _12449_ (.Y(_04577_),
    .A(_04467_),
    .B(net174));
 sg13g2_nand3_1 _12450_ (.B(_04577_),
    .C(net173),
    .A(_04576_),
    .Y(_04578_));
 sg13g2_nand3_1 _12451_ (.B(net190),
    .C(_04550_),
    .A(_04547_),
    .Y(_04579_));
 sg13g2_nand2_1 _12452_ (.Y(_04580_),
    .A(_04578_),
    .B(_04579_));
 sg13g2_nand2b_1 _12453_ (.Y(_04581_),
    .B(_04580_),
    .A_N(_04575_));
 sg13g2_nand3_1 _12454_ (.B(_04579_),
    .C(_04575_),
    .A(_04578_),
    .Y(_04582_));
 sg13g2_nand2_1 _12455_ (.Y(_04583_),
    .A(_04581_),
    .B(_04582_));
 sg13g2_inv_1 _12456_ (.Y(_04584_),
    .A(_04583_));
 sg13g2_nand3_1 _12457_ (.B(_04422_),
    .C(net155),
    .A(_04420_),
    .Y(_04585_));
 sg13g2_o21ai_1 _12458_ (.B1(_04585_),
    .Y(_04586_),
    .A1(net155),
    .A2(_04558_));
 sg13g2_nand3_1 _12459_ (.B(_04457_),
    .C(net173),
    .A(_04451_),
    .Y(_04587_));
 sg13g2_nand3_1 _12460_ (.B(_04563_),
    .C(net190),
    .A(_04562_),
    .Y(_04588_));
 sg13g2_nand2_1 _12461_ (.Y(_04589_),
    .A(_04587_),
    .B(_04588_));
 sg13g2_xor2_1 _12462_ (.B(_04589_),
    .A(_04586_),
    .X(_04590_));
 sg13g2_nand2_1 _12463_ (.Y(_04591_),
    .A(_04584_),
    .B(_04590_));
 sg13g2_nor2_1 _12464_ (.A(_04570_),
    .B(_04591_),
    .Y(_04592_));
 sg13g2_nand2_1 _12465_ (.Y(_04593_),
    .A(_04540_),
    .B(_04592_));
 sg13g2_nand2b_1 _12466_ (.Y(_04594_),
    .B(_04553_),
    .A_N(_04546_));
 sg13g2_inv_1 _12467_ (.Y(_04595_),
    .A(_04567_));
 sg13g2_nor2b_1 _12468_ (.A(_04553_),
    .B_N(_04546_),
    .Y(_04596_));
 sg13g2_a21oi_1 _12469_ (.A1(_04594_),
    .A2(_04595_),
    .Y(_04597_),
    .B1(_04596_));
 sg13g2_nor2_1 _12470_ (.A(_04597_),
    .B(_04591_),
    .Y(_04598_));
 sg13g2_nor2_1 _12471_ (.A(_04586_),
    .B(_04589_),
    .Y(_04599_));
 sg13g2_inv_1 _12472_ (.Y(_04600_),
    .A(_04582_));
 sg13g2_o21ai_1 _12473_ (.B1(_04581_),
    .Y(_04601_),
    .A1(_04599_),
    .A2(_04600_));
 sg13g2_nor2b_1 _12474_ (.A(_04598_),
    .B_N(_04601_),
    .Y(_04602_));
 sg13g2_nand2_1 _12475_ (.Y(_04603_),
    .A(_04593_),
    .B(_04602_));
 sg13g2_nand2b_1 _12476_ (.Y(_04604_),
    .B(_04603_),
    .A_N(_04479_));
 sg13g2_nand3_1 _12477_ (.B(_04479_),
    .C(_04602_),
    .A(_04593_),
    .Y(_04605_));
 sg13g2_nand2_1 _12478_ (.Y(_04606_),
    .A(_04604_),
    .B(_04605_));
 sg13g2_a21oi_1 _12479_ (.A1(_04503_),
    .A2(_04532_),
    .Y(_04607_),
    .B1(_04536_));
 sg13g2_inv_1 _12480_ (.Y(_04608_),
    .A(_04607_));
 sg13g2_nor2_1 _12481_ (.A(_04568_),
    .B(_04523_),
    .Y(_04609_));
 sg13g2_nand2_1 _12482_ (.Y(_04610_),
    .A(_04608_),
    .B(_04609_));
 sg13g2_a21oi_1 _12483_ (.A1(_04538_),
    .A2(_04566_),
    .Y(_04611_),
    .B1(_04595_));
 sg13g2_nand2_1 _12484_ (.Y(_04612_),
    .A(_04610_),
    .B(_04611_));
 sg13g2_nand2_1 _12485_ (.Y(_04613_),
    .A(_04590_),
    .B(_04554_));
 sg13g2_nor2_1 _12486_ (.A(_04583_),
    .B(_04479_),
    .Y(_04614_));
 sg13g2_inv_1 _12487_ (.Y(_04615_),
    .A(_04614_));
 sg13g2_nor2_1 _12488_ (.A(_04613_),
    .B(_04615_),
    .Y(_04616_));
 sg13g2_nor2_1 _12489_ (.A(_04596_),
    .B(_04599_),
    .Y(_04617_));
 sg13g2_nand2_1 _12490_ (.Y(_04618_),
    .A(_04589_),
    .B(_04586_));
 sg13g2_nor2b_1 _12491_ (.A(_04617_),
    .B_N(_04618_),
    .Y(_04619_));
 sg13g2_nand2_1 _12492_ (.Y(_04620_),
    .A(_04619_),
    .B(_04614_));
 sg13g2_inv_1 _12493_ (.Y(_04621_),
    .A(_04478_));
 sg13g2_o21ai_1 _12494_ (.B1(_04477_),
    .Y(_04622_),
    .A1(_04600_),
    .A2(_04621_));
 sg13g2_nand2_1 _12495_ (.Y(_04623_),
    .A(_04620_),
    .B(_04622_));
 sg13g2_a21oi_1 _12496_ (.A1(_04612_),
    .A2(_04616_),
    .Y(_04624_),
    .B1(_04623_));
 sg13g2_nor2b_1 _12497_ (.A(_04532_),
    .B_N(_04527_),
    .Y(_04625_));
 sg13g2_nand3_1 _12498_ (.B(_04501_),
    .C(_04503_),
    .A(_04625_),
    .Y(_04626_));
 sg13g2_inv_1 _12499_ (.Y(_04627_),
    .A(_04609_));
 sg13g2_nor2_1 _12500_ (.A(_04626_),
    .B(_04627_),
    .Y(_04628_));
 sg13g2_nand3_1 _12501_ (.B(_04628_),
    .C(_04531_),
    .A(_04616_),
    .Y(_04629_));
 sg13g2_nand2_1 _12502_ (.Y(_04630_),
    .A(_04624_),
    .B(_04629_));
 sg13g2_nor2_1 _12503_ (.A(_03696_),
    .B(net191),
    .Y(_04631_));
 sg13g2_a21oi_1 _12504_ (.A1(_00091_),
    .A2(net191),
    .Y(_04632_),
    .B1(_04631_));
 sg13g2_a21oi_1 _12505_ (.A1(_04632_),
    .A2(net137),
    .Y(_04633_),
    .B1(_04427_));
 sg13g2_a21o_1 _12506_ (.A2(_04573_),
    .A1(_04427_),
    .B1(_04633_),
    .X(_04634_));
 sg13g2_nand2b_1 _12507_ (.Y(_04635_),
    .B(net128),
    .A_N(_00084_));
 sg13g2_a21oi_1 _12508_ (.A1(net154),
    .A2(_00084_),
    .Y(_04636_),
    .B1(net175));
 sg13g2_a22oi_1 _12509_ (.Y(_04637_),
    .B1(net175),
    .B2(_04472_),
    .A2(_04636_),
    .A1(_04635_));
 sg13g2_nand2_1 _12510_ (.Y(_04638_),
    .A(_04637_),
    .B(net173));
 sg13g2_nand3_1 _12511_ (.B(_04577_),
    .C(net190),
    .A(_04576_),
    .Y(_04639_));
 sg13g2_nand2_1 _12512_ (.Y(_04640_),
    .A(_04638_),
    .B(_04639_));
 sg13g2_xnor2_1 _12513_ (.Y(_04641_),
    .A(_04634_),
    .B(_04640_));
 sg13g2_nand2_1 _12514_ (.Y(_04642_),
    .A(_04630_),
    .B(_04641_));
 sg13g2_inv_1 _12515_ (.Y(_04643_),
    .A(_04641_));
 sg13g2_nand3_1 _12516_ (.B(_04629_),
    .C(_04643_),
    .A(_04624_),
    .Y(_04644_));
 sg13g2_nand2_1 _12517_ (.Y(_04645_),
    .A(_04642_),
    .B(_04644_));
 sg13g2_buf_2 _12518_ (.A(_04645_),
    .X(_04646_));
 sg13g2_nand2b_1 _12519_ (.Y(_04647_),
    .B(_04646_),
    .A_N(_04606_));
 sg13g2_nand2_1 _12520_ (.Y(_04648_),
    .A(_04630_),
    .B(_04643_));
 sg13g2_nand3_1 _12521_ (.B(_04629_),
    .C(_04641_),
    .A(_04624_),
    .Y(_04649_));
 sg13g2_nand2_1 _12522_ (.Y(_04650_),
    .A(_04648_),
    .B(_04649_));
 sg13g2_buf_2 _12523_ (.A(_04650_),
    .X(_04651_));
 sg13g2_nand2_1 _12524_ (.Y(_04652_),
    .A(_04651_),
    .B(_04606_));
 sg13g2_nand2_1 _12525_ (.Y(_04653_),
    .A(_04647_),
    .B(_04652_));
 sg13g2_inv_1 _12526_ (.Y(_04654_),
    .A(\synth.voice.genblk4[10].next_state_scan[2] ));
 sg13g2_inv_1 _12527_ (.Y(_04655_),
    .A(\synth.voice.genblk4[9].next_state_scan[5] ));
 sg13g2_nor2b_1 _12528_ (.A(net255),
    .B_N(_00110_),
    .Y(_04656_));
 sg13g2_a221oi_1 _12529_ (.B2(net299),
    .C1(_04656_),
    .B1(_04655_),
    .A1(_04654_),
    .Y(_04657_),
    .A2(net300));
 sg13g2_buf_1 _12530_ (.A(_04657_),
    .X(_04658_));
 sg13g2_inv_1 _12531_ (.Y(_04659_),
    .A(\synth.voice.genblk4[10].next_state_scan[1] ));
 sg13g2_inv_1 _12532_ (.Y(_04660_),
    .A(\synth.voice.genblk4[9].next_state_scan[4] ));
 sg13g2_nor2b_1 _12533_ (.A(net255),
    .B_N(_00109_),
    .Y(_04661_));
 sg13g2_a221oi_1 _12534_ (.B2(net299),
    .C1(_04661_),
    .B1(_04660_),
    .A1(_04659_),
    .Y(_04662_),
    .A2(net300));
 sg13g2_inv_1 _12535_ (.Y(_04663_),
    .A(_04662_));
 sg13g2_nor2_1 _12536_ (.A(_04658_),
    .B(_04663_),
    .Y(_04664_));
 sg13g2_buf_2 _12537_ (.A(_04664_),
    .X(_04665_));
 sg13g2_nor2_1 _12538_ (.A(_04658_),
    .B(_04662_),
    .Y(_04666_));
 sg13g2_buf_2 _12539_ (.A(_04666_),
    .X(_04667_));
 sg13g2_inv_1 _12540_ (.Y(_04668_),
    .A(_04658_));
 sg13g2_nor2_1 _12541_ (.A(_04668_),
    .B(_04663_),
    .Y(_04669_));
 sg13g2_inv_1 _12542_ (.Y(_04670_),
    .A(\synth.voice.genblk4[10].next_state_scan[0] ));
 sg13g2_inv_1 _12543_ (.Y(_04671_),
    .A(\synth.voice.genblk4[9].next_state_scan[3] ));
 sg13g2_nor2b_1 _12544_ (.A(_01775_),
    .B_N(_00108_),
    .Y(_04672_));
 sg13g2_a221oi_1 _12545_ (.B2(net299),
    .C1(_04672_),
    .B1(_04671_),
    .A1(_04670_),
    .Y(_04673_),
    .A2(net300));
 sg13g2_buf_1 _12546_ (.A(_04673_),
    .X(_04674_));
 sg13g2_nand2_1 _12547_ (.Y(_04675_),
    .A(_04669_),
    .B(_04674_));
 sg13g2_o21ai_1 _12548_ (.B1(_04501_),
    .Y(_04676_),
    .A1(_04533_),
    .A2(_04504_));
 sg13g2_nand3b_1 _12549_ (.B(_04676_),
    .C(_04609_),
    .Y(_04677_),
    .A_N(_04613_));
 sg13g2_nor2_1 _12550_ (.A(_04611_),
    .B(_04613_),
    .Y(_04678_));
 sg13g2_nor2_1 _12551_ (.A(_04619_),
    .B(_04678_),
    .Y(_04679_));
 sg13g2_nand2_1 _12552_ (.Y(_04680_),
    .A(_04677_),
    .B(_04679_));
 sg13g2_xnor2_1 _12553_ (.Y(_04681_),
    .A(_04583_),
    .B(_04680_));
 sg13g2_nor2_1 _12554_ (.A(_04675_),
    .B(_04681_),
    .Y(_04682_));
 sg13g2_nor2_1 _12555_ (.A(_04667_),
    .B(_04682_),
    .Y(_04683_));
 sg13g2_nor3_1 _12556_ (.A(_04662_),
    .B(_04674_),
    .C(_04668_),
    .Y(_04684_));
 sg13g2_nand2_1 _12557_ (.Y(_04685_),
    .A(_04651_),
    .B(_04684_));
 sg13g2_nand2_1 _12558_ (.Y(_04686_),
    .A(_04683_),
    .B(_04685_));
 sg13g2_a21oi_1 _12559_ (.A1(_04653_),
    .A2(_04665_),
    .Y(_04687_),
    .B1(_04686_));
 sg13g2_nand3_1 _12560_ (.B(_04658_),
    .C(_04674_),
    .A(_04663_),
    .Y(_04688_));
 sg13g2_nand2_1 _12561_ (.Y(_04689_),
    .A(_04646_),
    .B(_04681_));
 sg13g2_nand2b_1 _12562_ (.Y(_04690_),
    .B(_04689_),
    .A_N(_04688_));
 sg13g2_inv_1 _12563_ (.Y(_04691_),
    .A(_04669_));
 sg13g2_nand2_1 _12564_ (.Y(_04692_),
    .A(_04690_),
    .B(_04691_));
 sg13g2_nand2_1 _12565_ (.Y(_04693_),
    .A(_04692_),
    .B(_04647_));
 sg13g2_nand2_1 _12566_ (.Y(_04694_),
    .A(_04687_),
    .B(_04693_));
 sg13g2_nand2_1 _12567_ (.Y(_04695_),
    .A(_01776_),
    .B(\synth.voice.genblk4[9].next_state_scan[2] ));
 sg13g2_a22oi_1 _12568_ (.Y(_04696_),
    .B1(\synth.voice.params[25] ),
    .B2(net299),
    .A2(\synth.voice.genblk4[10].next_state_scan[12] ),
    .A1(_01745_));
 sg13g2_a21oi_1 _12569_ (.A1(_04695_),
    .A2(_04696_),
    .Y(_04697_),
    .B1(net176));
 sg13g2_buf_8 _12570_ (.A(_04646_),
    .X(_04698_));
 sg13g2_inv_1 _12571_ (.Y(_04699_),
    .A(_01758_));
 sg13g2_nor2_2 _12572_ (.A(_04699_),
    .B(_01740_),
    .Y(_04700_));
 sg13g2_inv_1 _12573_ (.Y(_04701_),
    .A(_04700_));
 sg13g2_buf_1 _12574_ (.A(_04701_),
    .X(_04702_));
 sg13g2_a21oi_1 _12575_ (.A1(net34),
    .A2(_04667_),
    .Y(_04703_),
    .B1(net136));
 sg13g2_nand3_1 _12576_ (.B(_04697_),
    .C(_04703_),
    .A(_04694_),
    .Y(_04704_));
 sg13g2_nor2_1 _12577_ (.A(_04391_),
    .B(net176),
    .Y(_04705_));
 sg13g2_a22oi_1 _12578_ (.Y(_04706_),
    .B1(net136),
    .B2(_04705_),
    .A2(_04358_),
    .A1(\synth.voice.genblk4[8].next_state_scan[7] ));
 sg13g2_nand2_1 _12579_ (.Y(_01137_),
    .A(_04704_),
    .B(_04706_));
 sg13g2_xnor2_1 _12580_ (.Y(_04707_),
    .A(_03679_),
    .B(_04369_));
 sg13g2_inv_1 _12581_ (.Y(_04708_),
    .A(_04211_));
 sg13g2_nor2_1 _12582_ (.A(\synth.voice.genblk4[1].next_state_scan[4] ),
    .B(net135),
    .Y(_04709_));
 sg13g2_a21oi_1 _12583_ (.A1(_04707_),
    .A2(net135),
    .Y(_04710_),
    .B1(_04709_));
 sg13g2_buf_1 _12584_ (.A(_03609_),
    .X(_04711_));
 sg13g2_inv_1 _12585_ (.Y(_04712_),
    .A(\synth.voice.genblk4[0].next_state_scan[13] ));
 sg13g2_nor2_1 _12586_ (.A(_04712_),
    .B(net189),
    .Y(_04713_));
 sg13g2_a21oi_1 _12587_ (.A1(_04710_),
    .A2(net189),
    .Y(_04714_),
    .B1(_04713_));
 sg13g2_nor2_1 _12588_ (.A(\synth.voice.genblk4[0].next_state_scan[11] ),
    .B(net43),
    .Y(_04715_));
 sg13g2_a21oi_1 _12589_ (.A1(net44),
    .A2(_04714_),
    .Y(_01142_),
    .B1(_04715_));
 sg13g2_inv_1 _12590_ (.Y(_04716_),
    .A(_04348_));
 sg13g2_nand2_1 _12591_ (.Y(_04717_),
    .A(_04245_),
    .B(_03597_));
 sg13g2_nand3_1 _12592_ (.B(_03592_),
    .C(_04351_),
    .A(_04249_),
    .Y(_04718_));
 sg13g2_o21ai_1 _12593_ (.B1(_04718_),
    .Y(_04719_),
    .A1(_04716_),
    .A2(_04717_));
 sg13g2_buf_1 _12594_ (.A(_04719_),
    .X(_04720_));
 sg13g2_buf_1 _12595_ (.A(_04720_),
    .X(_04721_));
 sg13g2_mux2_1 _12596_ (.A0(\synth.voice.params[8] ),
    .A1(\synth.voice.genblk4[9].next_state_scan[0] ),
    .S(net210),
    .X(_01147_));
 sg13g2_mux2_1 _12597_ (.A0(\synth.voice.params[9] ),
    .A1(\synth.voice.genblk4[9].next_state_scan[1] ),
    .S(net210),
    .X(_01148_));
 sg13g2_mux2_1 _12598_ (.A0(\synth.voice.genblk4[9].next_state_scan[0] ),
    .A1(\synth.voice.genblk4[9].next_state_scan[2] ),
    .S(net210),
    .X(_01149_));
 sg13g2_buf_1 _12599_ (.A(_04720_),
    .X(_04722_));
 sg13g2_buf_1 _12600_ (.A(net209),
    .X(_04723_));
 sg13g2_nor2_1 _12601_ (.A(\synth.voice.genblk4[9].next_state_scan[1] ),
    .B(net210),
    .Y(_04724_));
 sg13g2_a21oi_1 _12602_ (.A1(_04671_),
    .A2(net188),
    .Y(_01150_),
    .B1(_04724_));
 sg13g2_nor2_1 _12603_ (.A(\synth.voice.genblk4[9].next_state_scan[2] ),
    .B(net210),
    .Y(_04725_));
 sg13g2_a21oi_1 _12604_ (.A1(_04660_),
    .A2(_04723_),
    .Y(_01151_),
    .B1(_04725_));
 sg13g2_nor2_1 _12605_ (.A(\synth.voice.genblk4[9].next_state_scan[3] ),
    .B(net210),
    .Y(_04726_));
 sg13g2_a21oi_1 _12606_ (.A1(_04655_),
    .A2(net188),
    .Y(_01152_),
    .B1(_04726_));
 sg13g2_inv_1 _12607_ (.Y(_04727_),
    .A(\synth.voice.genblk4[0].next_state_scan[12] ));
 sg13g2_nor4_1 _12608_ (.A(_03695_),
    .B(_03680_),
    .C(_03619_),
    .D(_03642_),
    .Y(_04728_));
 sg13g2_a21oi_1 _12609_ (.A1(_04225_),
    .A2(_04728_),
    .Y(_04729_),
    .B1(_03699_));
 sg13g2_nand3_1 _12610_ (.B(_03699_),
    .C(_04728_),
    .A(_04225_),
    .Y(_04730_));
 sg13g2_nor2b_1 _12611_ (.A(_04729_),
    .B_N(_04730_),
    .Y(_04731_));
 sg13g2_inv_1 _12612_ (.Y(_04732_),
    .A(\synth.voice.genblk4[1].next_state_scan[5] ));
 sg13g2_nor2_1 _12613_ (.A(_04732_),
    .B(net135),
    .Y(_04733_));
 sg13g2_a21oi_1 _12614_ (.A1(_04731_),
    .A2(net135),
    .Y(_04734_),
    .B1(_04733_));
 sg13g2_nand2_1 _12615_ (.Y(_04735_),
    .A(_04230_),
    .B(_03370_));
 sg13g2_o21ai_1 _12616_ (.B1(_04735_),
    .Y(_04736_),
    .A1(net182),
    .A2(_04734_));
 sg13g2_nand2_1 _12617_ (.Y(_04737_),
    .A(net43),
    .B(_04736_));
 sg13g2_o21ai_1 _12618_ (.B1(_04737_),
    .Y(_01153_),
    .A1(_04727_),
    .A2(net44));
 sg13g2_nor2_1 _12619_ (.A(\synth.voice.genblk4[9].next_state_scan[4] ),
    .B(net209),
    .Y(_04738_));
 sg13g2_a21oi_1 _12620_ (.A1(_04415_),
    .A2(net188),
    .Y(_01154_),
    .B1(_04738_));
 sg13g2_nor2_1 _12621_ (.A(\synth.voice.genblk4[9].next_state_scan[5] ),
    .B(net209),
    .Y(_04739_));
 sg13g2_a21oi_1 _12622_ (.A1(_04424_),
    .A2(net188),
    .Y(_01155_),
    .B1(_04739_));
 sg13g2_nor2_1 _12623_ (.A(\synth.voice.genblk4[9].next_state_scan[6] ),
    .B(net209),
    .Y(_04740_));
 sg13g2_a21oi_1 _12624_ (.A1(_04446_),
    .A2(net188),
    .Y(_01156_),
    .B1(_04740_));
 sg13g2_nor2_1 _12625_ (.A(\synth.voice.genblk4[9].next_state_scan[7] ),
    .B(net209),
    .Y(_04741_));
 sg13g2_a21oi_1 _12626_ (.A1(_04459_),
    .A2(net188),
    .Y(_01157_),
    .B1(_04741_));
 sg13g2_nor2_1 _12627_ (.A(\synth.voice.genblk4[9].next_state_scan[8] ),
    .B(net209),
    .Y(_04742_));
 sg13g2_a21oi_1 _12628_ (.A1(_04406_),
    .A2(net188),
    .Y(_01158_),
    .B1(_04742_));
 sg13g2_nor2_1 _12629_ (.A(\synth.voice.genblk4[9].next_state_scan[9] ),
    .B(net209),
    .Y(_04743_));
 sg13g2_a21oi_1 _12630_ (.A1(_04400_),
    .A2(net188),
    .Y(_01159_),
    .B1(_04743_));
 sg13g2_nor2_1 _12631_ (.A(\synth.voice.genblk4[9].next_state_scan[10] ),
    .B(net209),
    .Y(_04744_));
 sg13g2_a21oi_1 _12632_ (.A1(_01770_),
    .A2(_04723_),
    .Y(_01160_),
    .B1(_04744_));
 sg13g2_nand2_1 _12633_ (.Y(_04745_),
    .A(net210),
    .B(\synth.voice.genblk4[9].next_state_scan[13] ));
 sg13g2_o21ai_1 _12634_ (.B1(_04745_),
    .Y(_01161_),
    .A1(_04400_),
    .A2(_04721_));
 sg13g2_nor2_1 _12635_ (.A(\synth.voice.genblk4[9].next_state_scan[12] ),
    .B(_04722_),
    .Y(_04746_));
 sg13g2_a21oi_1 _12636_ (.A1(net377),
    .A2(net210),
    .Y(_01162_),
    .B1(_04746_));
 sg13g2_nor2_1 _12637_ (.A(\synth.voice.genblk4[9].next_state_scan[13] ),
    .B(_04722_),
    .Y(_04747_));
 sg13g2_a21oi_1 _12638_ (.A1(_03383_),
    .A2(_04721_),
    .Y(_01163_),
    .B1(_04747_));
 sg13g2_inv_1 _12639_ (.Y(_04748_),
    .A(_03704_));
 sg13g2_xnor2_1 _12640_ (.Y(_04749_),
    .A(_04748_),
    .B(_04730_));
 sg13g2_nor2_1 _12641_ (.A(net139),
    .B(_04749_),
    .Y(_04750_));
 sg13g2_a21oi_1 _12642_ (.A1(\synth.voice.genblk4[1].next_state_scan[6] ),
    .A2(net139),
    .Y(_04751_),
    .B1(_04750_));
 sg13g2_nand2_1 _12643_ (.Y(_04752_),
    .A(net180),
    .B(net401));
 sg13g2_o21ai_1 _12644_ (.B1(_04752_),
    .Y(_04753_),
    .A1(net180),
    .A2(_04751_));
 sg13g2_nand2_1 _12645_ (.Y(_04754_),
    .A(net43),
    .B(_04753_));
 sg13g2_o21ai_1 _12646_ (.B1(_04754_),
    .Y(_01164_),
    .A1(_04712_),
    .A2(net44));
 sg13g2_inv_1 _12647_ (.Y(_04755_),
    .A(_04021_));
 sg13g2_nand3_1 _12648_ (.B(_03591_),
    .C(_04351_),
    .A(_03593_),
    .Y(_04756_));
 sg13g2_o21ai_1 _12649_ (.B1(_04756_),
    .Y(_04757_),
    .A1(_04716_),
    .A2(_04755_));
 sg13g2_buf_1 _12650_ (.A(_04757_),
    .X(_04758_));
 sg13g2_buf_1 _12651_ (.A(_04758_),
    .X(_04759_));
 sg13g2_buf_1 _12652_ (.A(_04758_),
    .X(_04760_));
 sg13g2_nor2_1 _12653_ (.A(\synth.voice.params[24] ),
    .B(net171),
    .Y(_04761_));
 sg13g2_a21oi_1 _12654_ (.A1(_04670_),
    .A2(_04759_),
    .Y(_01165_),
    .B1(_04761_));
 sg13g2_nor2_1 _12655_ (.A(\synth.voice.params[25] ),
    .B(net171),
    .Y(_04762_));
 sg13g2_a21oi_1 _12656_ (.A1(_04659_),
    .A2(net172),
    .Y(_01166_),
    .B1(_04762_));
 sg13g2_buf_1 _12657_ (.A(_04758_),
    .X(_04763_));
 sg13g2_nor2_1 _12658_ (.A(\synth.voice.genblk4[10].next_state_scan[0] ),
    .B(net170),
    .Y(_04764_));
 sg13g2_a21oi_1 _12659_ (.A1(_04654_),
    .A2(net172),
    .Y(_01167_),
    .B1(_04764_));
 sg13g2_nor2_1 _12660_ (.A(\synth.voice.genblk4[10].next_state_scan[1] ),
    .B(net170),
    .Y(_04765_));
 sg13g2_a21oi_1 _12661_ (.A1(_04414_),
    .A2(net172),
    .Y(_01168_),
    .B1(_04765_));
 sg13g2_nor2_1 _12662_ (.A(\synth.voice.genblk4[10].next_state_scan[2] ),
    .B(net170),
    .Y(_04766_));
 sg13g2_a21oi_1 _12663_ (.A1(_04423_),
    .A2(net172),
    .Y(_01169_),
    .B1(_04766_));
 sg13g2_nor2_1 _12664_ (.A(\synth.voice.genblk4[10].next_state_scan[3] ),
    .B(net170),
    .Y(_04767_));
 sg13g2_a21oi_1 _12665_ (.A1(_04445_),
    .A2(net172),
    .Y(_01170_),
    .B1(_04767_));
 sg13g2_nor2_1 _12666_ (.A(\synth.voice.genblk4[10].next_state_scan[4] ),
    .B(net170),
    .Y(_04768_));
 sg13g2_a21oi_1 _12667_ (.A1(_04458_),
    .A2(net172),
    .Y(_01171_),
    .B1(_04768_));
 sg13g2_nor2_1 _12668_ (.A(\synth.voice.genblk4[10].next_state_scan[5] ),
    .B(net170),
    .Y(_04769_));
 sg13g2_a21oi_1 _12669_ (.A1(_04405_),
    .A2(net172),
    .Y(_01172_),
    .B1(_04769_));
 sg13g2_nor2_1 _12670_ (.A(\synth.voice.genblk4[10].next_state_scan[6] ),
    .B(net170),
    .Y(_04770_));
 sg13g2_a21oi_1 _12671_ (.A1(_04399_),
    .A2(net172),
    .Y(_01173_),
    .B1(_04770_));
 sg13g2_nand2_1 _12672_ (.Y(_04771_),
    .A(net171),
    .B(\synth.voice.genblk4[10].next_state_scan[9] ));
 sg13g2_o21ai_1 _12673_ (.B1(_04771_),
    .Y(_01174_),
    .A1(_04405_),
    .A2(net171));
 sg13g2_nor4_1 _12674_ (.A(\synth.voice.genblk4[1].next_state_scan[0] ),
    .B(\synth.voice.genblk4[1].next_state_scan[3] ),
    .C(\synth.voice.genblk4[1].next_state_scan[2] ),
    .D(\synth.voice.genblk4[1].next_state_scan[5] ),
    .Y(_04772_));
 sg13g2_nor4_1 _12675_ (.A(\synth.voice.genblk4[1].next_state_scan[4] ),
    .B(\synth.voice.genblk4[1].next_state_scan[7] ),
    .C(\synth.voice.genblk4[1].next_state_scan[6] ),
    .D(\synth.voice.genblk4[8].next_state_scan[1] ),
    .Y(_04773_));
 sg13g2_nor2_1 _12676_ (.A(\synth.voice.lfsr[1] ),
    .B(\synth.voice.genblk4[1].next_state_scan[1] ),
    .Y(_04774_));
 sg13g2_nor3_1 _12677_ (.A(\synth.voice.genblk4[8].next_state_scan[0] ),
    .B(\synth.voice.genblk4[8].next_state_scan[3] ),
    .C(\synth.voice.genblk4[8].next_state_scan[2] ),
    .Y(_04775_));
 sg13g2_nand4_1 _12678_ (.B(_04773_),
    .C(_04774_),
    .A(_04772_),
    .Y(_04776_),
    .D(_04775_));
 sg13g2_inv_1 _12679_ (.Y(_04777_),
    .A(\synth.voice.lfsr[0] ));
 sg13g2_nand3b_1 _12680_ (.B(_04776_),
    .C(_04777_),
    .Y(_04778_),
    .A_N(\synth.voice.genblk4[8].next_state_scan[4] ));
 sg13g2_a21oi_1 _12681_ (.A1(\synth.voice.genblk4[8].next_state_scan[4] ),
    .A2(\synth.voice.lfsr[0] ),
    .Y(_04779_),
    .B1(_04708_));
 sg13g2_xnor2_1 _12682_ (.Y(_04780_),
    .A(_03663_),
    .B(_03659_));
 sg13g2_a22oi_1 _12683_ (.Y(_04781_),
    .B1(_04708_),
    .B2(_04780_),
    .A2(_04779_),
    .A1(_04778_));
 sg13g2_inv_1 _12684_ (.Y(_04782_),
    .A(_04781_));
 sg13g2_inv_1 _12685_ (.Y(_04783_),
    .A(_04717_));
 sg13g2_nand2_1 _12686_ (.Y(_04784_),
    .A(_04249_),
    .B(_03592_));
 sg13g2_inv_1 _12687_ (.Y(_04785_),
    .A(_03590_));
 sg13g2_nor2_1 _12688_ (.A(_04784_),
    .B(_04785_),
    .Y(_04786_));
 sg13g2_a21oi_1 _12689_ (.A1(_03607_),
    .A2(_04783_),
    .Y(_04787_),
    .B1(_04786_));
 sg13g2_buf_1 _12690_ (.A(_04787_),
    .X(_04788_));
 sg13g2_nand2_1 _12691_ (.Y(_04789_),
    .A(_04782_),
    .B(_04788_));
 sg13g2_inv_1 _12692_ (.Y(_04790_),
    .A(_04204_));
 sg13g2_nor2_1 _12693_ (.A(_04789_),
    .B(_04790_),
    .Y(_04791_));
 sg13g2_nand4_1 _12694_ (.B(_03702_),
    .C(\synth.voice.genblk4[11].next_state_scan[3] ),
    .A(_04749_),
    .Y(_04792_),
    .D(_01736_));
 sg13g2_a21oi_1 _12695_ (.A1(_04792_),
    .A2(net181),
    .Y(_04793_),
    .B1(_04201_));
 sg13g2_nand3_1 _12696_ (.B(_04793_),
    .C(net143),
    .A(_04199_),
    .Y(_04794_));
 sg13g2_buf_2 _12697_ (.A(_04794_),
    .X(_04795_));
 sg13g2_nand2_1 _12698_ (.Y(_04796_),
    .A(_04795_),
    .B(_04788_));
 sg13g2_buf_8 _12699_ (.A(_04796_),
    .X(_04797_));
 sg13g2_nand2_1 _12700_ (.Y(_04798_),
    .A(_04791_),
    .B(_04797_));
 sg13g2_buf_1 _12701_ (.A(_04788_),
    .X(_04799_));
 sg13g2_nand3_1 _12702_ (.B(\synth.voice.lfsr[0] ),
    .C(net153),
    .A(_04795_),
    .Y(_04800_));
 sg13g2_inv_1 _12703_ (.Y(_04801_),
    .A(_04788_));
 sg13g2_buf_1 _12704_ (.A(_04801_),
    .X(_04802_));
 sg13g2_buf_1 _12705_ (.A(net134),
    .X(_04803_));
 sg13g2_nand2_1 _12706_ (.Y(_04804_),
    .A(net127),
    .B(\synth.voice.genblk4[1].next_state_scan[0] ));
 sg13g2_nand3_1 _12707_ (.B(_04800_),
    .C(_04804_),
    .A(_04798_),
    .Y(_01175_));
 sg13g2_nor2_1 _12708_ (.A(\synth.voice.genblk4[10].next_state_scan[8] ),
    .B(net170),
    .Y(_04805_));
 sg13g2_a21oi_1 _12709_ (.A1(_01784_),
    .A2(_04759_),
    .Y(_01176_),
    .B1(_04805_));
 sg13g2_nor2_1 _12710_ (.A(\synth.voice.genblk4[10].next_state_scan[9] ),
    .B(_04763_),
    .Y(_04806_));
 sg13g2_a21oi_1 _12711_ (.A1(_01781_),
    .A2(_04760_),
    .Y(_01177_),
    .B1(_04806_));
 sg13g2_nand2_1 _12712_ (.Y(_04807_),
    .A(net171),
    .B(\synth.voice.genblk4[10].next_state_scan[12] ));
 sg13g2_o21ai_1 _12713_ (.B1(_04807_),
    .Y(_01178_),
    .A1(_01784_),
    .A2(net171));
 sg13g2_nor2_1 _12714_ (.A(\synth.voice.genblk4[10].next_state_scan[11] ),
    .B(_04763_),
    .Y(_04808_));
 sg13g2_a21oi_1 _12715_ (.A1(_04209_),
    .A2(_04760_),
    .Y(_01179_),
    .B1(_04808_));
 sg13g2_nor2_1 _12716_ (.A(\synth.voice.genblk4[10].next_state_scan[12] ),
    .B(_04758_),
    .Y(_04809_));
 sg13g2_a21oi_1 _12717_ (.A1(net377),
    .A2(net171),
    .Y(_01180_),
    .B1(_04809_));
 sg13g2_nor2_1 _12718_ (.A(\synth.voice.genblk4[10].next_state_scan[13] ),
    .B(_04758_),
    .Y(_04810_));
 sg13g2_a21oi_1 _12719_ (.A1(_03383_),
    .A2(net171),
    .Y(_01181_),
    .B1(_04810_));
 sg13g2_nand2_1 _12720_ (.Y(_04811_),
    .A(_03599_),
    .B(_04348_));
 sg13g2_nor2_1 _12721_ (.A(_04350_),
    .B(_03587_),
    .Y(_04812_));
 sg13g2_nand2_1 _12722_ (.Y(_04813_),
    .A(_04250_),
    .B(_04812_));
 sg13g2_o21ai_1 _12723_ (.B1(_04813_),
    .Y(_04814_),
    .A1(_04811_),
    .A2(_04247_));
 sg13g2_buf_1 _12724_ (.A(_04814_),
    .X(_04815_));
 sg13g2_buf_1 _12725_ (.A(net208),
    .X(_04816_));
 sg13g2_buf_1 _12726_ (.A(_04815_),
    .X(_04817_));
 sg13g2_nand2_1 _12727_ (.Y(_04818_),
    .A(net186),
    .B(\synth.voice.bpf_en[0] ));
 sg13g2_o21ai_1 _12728_ (.B1(_04818_),
    .Y(_01182_),
    .A1(_01766_),
    .A2(_04816_));
 sg13g2_nor2_1 _12729_ (.A(_01765_),
    .B(net208),
    .Y(_04819_));
 sg13g2_a21oi_1 _12730_ (.A1(_01741_),
    .A2(net187),
    .Y(_01183_),
    .B1(_04819_));
 sg13g2_mux2_1 _12731_ (.A0(\synth.voice.bpf_en[0] ),
    .A1(\synth.voice.bpf_en[2] ),
    .S(_04817_),
    .X(_01184_));
 sg13g2_nand2_1 _12732_ (.Y(_04820_),
    .A(_04817_),
    .B(\synth.voice.genblk4[11].next_state_scan[3] ));
 sg13g2_o21ai_1 _12733_ (.B1(_04820_),
    .Y(_01185_),
    .A1(_01741_),
    .A2(_04816_));
 sg13g2_nor2_1 _12734_ (.A(_04214_),
    .B(_04213_),
    .Y(_04821_));
 sg13g2_inv_1 _12735_ (.Y(_04822_),
    .A(_04215_));
 sg13g2_nor3_1 _12736_ (.A(_04212_),
    .B(_04821_),
    .C(_04822_),
    .Y(_04823_));
 sg13g2_a21oi_1 _12737_ (.A1(_03660_),
    .A2(_04212_),
    .Y(_04824_),
    .B1(_04823_));
 sg13g2_inv_1 _12738_ (.Y(_04825_),
    .A(_04824_));
 sg13g2_nand2_1 _12739_ (.Y(_04826_),
    .A(_04825_),
    .B(_04788_));
 sg13g2_nor2_1 _12740_ (.A(_04826_),
    .B(_04790_),
    .Y(_04827_));
 sg13g2_nand2_1 _12741_ (.Y(_04828_),
    .A(_04827_),
    .B(net42));
 sg13g2_nand3_1 _12742_ (.B(\synth.voice.lfsr[1] ),
    .C(net153),
    .A(_04795_),
    .Y(_04829_));
 sg13g2_nand2_1 _12743_ (.Y(_04830_),
    .A(net127),
    .B(\synth.voice.genblk4[1].next_state_scan[1] ));
 sg13g2_nand3_1 _12744_ (.B(_04829_),
    .C(_04830_),
    .A(_04828_),
    .Y(_01186_));
 sg13g2_inv_1 _12745_ (.Y(_04831_),
    .A(\synth.voice.genblk4[11].next_state_scan[4] ));
 sg13g2_nor2_1 _12746_ (.A(\synth.voice.bpf_en[2] ),
    .B(net208),
    .Y(_04832_));
 sg13g2_a21oi_1 _12747_ (.A1(_04831_),
    .A2(net187),
    .Y(_01187_),
    .B1(_04832_));
 sg13g2_inv_1 _12748_ (.Y(_04833_),
    .A(\synth.voice.genblk4[11].next_state_scan[5] ));
 sg13g2_nor2_1 _12749_ (.A(\synth.voice.genblk4[11].next_state_scan[3] ),
    .B(net208),
    .Y(_04834_));
 sg13g2_a21oi_1 _12750_ (.A1(_04833_),
    .A2(net187),
    .Y(_01188_),
    .B1(_04834_));
 sg13g2_inv_1 _12751_ (.Y(_04835_),
    .A(\synth.voice.genblk4[11].next_state_scan[6] ));
 sg13g2_nor2_1 _12752_ (.A(\synth.voice.genblk4[11].next_state_scan[4] ),
    .B(net208),
    .Y(_04836_));
 sg13g2_a21oi_1 _12753_ (.A1(_04835_),
    .A2(net187),
    .Y(_01189_),
    .B1(_04836_));
 sg13g2_inv_1 _12754_ (.Y(_04837_),
    .A(\synth.voice.genblk4[11].next_state_scan[7] ));
 sg13g2_nor2_1 _12755_ (.A(\synth.voice.genblk4[11].next_state_scan[5] ),
    .B(net208),
    .Y(_04838_));
 sg13g2_a21oi_1 _12756_ (.A1(_04837_),
    .A2(net187),
    .Y(_01190_),
    .B1(_04838_));
 sg13g2_nand2_1 _12757_ (.Y(_04839_),
    .A(net186),
    .B(\synth.voice.genblk4[11].next_state_scan[8] ));
 sg13g2_o21ai_1 _12758_ (.B1(_04839_),
    .Y(_01191_),
    .A1(_04835_),
    .A2(net187));
 sg13g2_nand2_1 _12759_ (.Y(_04840_),
    .A(net186),
    .B(\synth.voice.genblk4[11].next_state_scan[9] ));
 sg13g2_o21ai_1 _12760_ (.B1(_04840_),
    .Y(_01192_),
    .A1(_04837_),
    .A2(net186));
 sg13g2_mux2_1 _12761_ (.A0(\synth.voice.genblk4[11].next_state_scan[8] ),
    .A1(\synth.voice.genblk4[11].next_state_scan[10] ),
    .S(net186),
    .X(_01193_));
 sg13g2_mux2_1 _12762_ (.A0(\synth.voice.genblk4[11].next_state_scan[9] ),
    .A1(\synth.voice.genblk4[11].next_state_scan[11] ),
    .S(net186),
    .X(_01194_));
 sg13g2_mux2_1 _12763_ (.A0(\synth.voice.genblk4[11].next_state_scan[10] ),
    .A1(\synth.voice.genblk4[11].next_state_scan[12] ),
    .S(net186),
    .X(_01195_));
 sg13g2_mux2_1 _12764_ (.A0(\synth.voice.genblk4[11].next_state_scan[11] ),
    .A1(\synth.voice.genblk4[11].next_state_scan[13] ),
    .S(net186),
    .X(_01196_));
 sg13g2_xnor2_1 _12765_ (.Y(_04841_),
    .A(_04218_),
    .B(_04216_));
 sg13g2_nor2_1 _12766_ (.A(_04491_),
    .B(net135),
    .Y(_04842_));
 sg13g2_a21o_1 _12767_ (.A2(net135),
    .A1(_04841_),
    .B1(_04842_),
    .X(_04843_));
 sg13g2_nor2_1 _12768_ (.A(net134),
    .B(_04843_),
    .Y(_04844_));
 sg13g2_nor2b_1 _12769_ (.A(_04790_),
    .B_N(_04844_),
    .Y(_04845_));
 sg13g2_nand2_1 _12770_ (.Y(_04846_),
    .A(_04845_),
    .B(net42));
 sg13g2_nand3_1 _12771_ (.B(\synth.voice.genblk4[1].next_state_scan[0] ),
    .C(_04799_),
    .A(_04795_),
    .Y(_04847_));
 sg13g2_nand2_1 _12772_ (.Y(_04848_),
    .A(net127),
    .B(\synth.voice.genblk4[1].next_state_scan[2] ));
 sg13g2_nand3_1 _12773_ (.B(_04847_),
    .C(_04848_),
    .A(_04846_),
    .Y(_01197_));
 sg13g2_nor2_1 _12774_ (.A(\synth.voice.genblk4[11].next_state_scan[12] ),
    .B(net208),
    .Y(_04849_));
 sg13g2_a21oi_1 _12775_ (.A1(net377),
    .A2(net187),
    .Y(_01198_),
    .B1(_04849_));
 sg13g2_nor2_1 _12776_ (.A(\synth.voice.genblk4[11].next_state_scan[13] ),
    .B(net208),
    .Y(_04850_));
 sg13g2_a21oi_1 _12777_ (.A1(_03383_),
    .A2(net187),
    .Y(_01199_),
    .B1(_04850_));
 sg13g2_xnor2_1 _12778_ (.Y(_04851_),
    .A(_04222_),
    .B(_04221_));
 sg13g2_nor2_1 _12779_ (.A(_03630_),
    .B(net135),
    .Y(_04852_));
 sg13g2_a21o_1 _12780_ (.A2(net135),
    .A1(_04851_),
    .B1(_04852_),
    .X(_04853_));
 sg13g2_nor2_1 _12781_ (.A(net134),
    .B(_04853_),
    .Y(_04854_));
 sg13g2_nor2b_1 _12782_ (.A(_04790_),
    .B_N(_04854_),
    .Y(_04855_));
 sg13g2_nand2_1 _12783_ (.Y(_04856_),
    .A(_04855_),
    .B(_04797_));
 sg13g2_nand3_1 _12784_ (.B(\synth.voice.genblk4[1].next_state_scan[1] ),
    .C(_04799_),
    .A(_04795_),
    .Y(_04857_));
 sg13g2_nand2_1 _12785_ (.Y(_04858_),
    .A(net127),
    .B(\synth.voice.genblk4[1].next_state_scan[3] ));
 sg13g2_nand3_1 _12786_ (.B(_04857_),
    .C(_04858_),
    .A(_04856_),
    .Y(_01200_));
 sg13g2_nand2_1 _12787_ (.Y(_04859_),
    .A(net181),
    .B(_03875_));
 sg13g2_o21ai_1 _12788_ (.B1(_04859_),
    .Y(_04860_),
    .A1(_03874_),
    .A2(net181));
 sg13g2_nand3_1 _12789_ (.B(_03665_),
    .C(_04860_),
    .A(_03664_),
    .Y(_04861_));
 sg13g2_nand3_1 _12790_ (.B(_03609_),
    .C(_03422_),
    .A(_04861_),
    .Y(_04862_));
 sg13g2_nor2b_1 _12791_ (.A(net193),
    .B_N(\synth.voice.float_period[1][3] ),
    .Y(_04863_));
 sg13g2_a21oi_1 _12792_ (.A1(\synth.voice.float_period[0][3] ),
    .A2(net193),
    .Y(_04864_),
    .B1(_04863_));
 sg13g2_inv_1 _12793_ (.Y(_04865_),
    .A(_03715_));
 sg13g2_nand2_1 _12794_ (.Y(_04866_),
    .A(net193),
    .B(_03746_));
 sg13g2_o21ai_1 _12795_ (.B1(_04866_),
    .Y(_04867_),
    .A1(_03747_),
    .A2(net193));
 sg13g2_nand2_1 _12796_ (.Y(_04868_),
    .A(_04865_),
    .B(_04867_));
 sg13g2_o21ai_1 _12797_ (.B1(_04868_),
    .Y(_04869_),
    .A1(_03708_),
    .A2(_04864_));
 sg13g2_nand3_1 _12798_ (.B(_04748_),
    .C(_03711_),
    .A(_03659_),
    .Y(_04870_));
 sg13g2_nor2_1 _12799_ (.A(_04870_),
    .B(_03706_),
    .Y(_04871_));
 sg13g2_a21oi_1 _12800_ (.A1(net159),
    .A2(_03693_),
    .Y(_04872_),
    .B1(_04871_));
 sg13g2_a21o_1 _12801_ (.A2(_04870_),
    .A1(_03706_),
    .B1(_04872_),
    .X(_04873_));
 sg13g2_a22oi_1 _12802_ (.Y(_04874_),
    .B1(net159),
    .B2(_03701_),
    .A2(_04217_),
    .A1(_03704_));
 sg13g2_nor2b_1 _12803_ (.A(_03686_),
    .B_N(_03688_),
    .Y(_04875_));
 sg13g2_nand2_1 _12804_ (.Y(_04876_),
    .A(_04874_),
    .B(_04875_));
 sg13g2_nor2_1 _12805_ (.A(_04875_),
    .B(_04874_),
    .Y(_04877_));
 sg13g2_a221oi_1 _12806_ (.B2(_04876_),
    .C1(_04877_),
    .B1(_04873_),
    .A1(_03708_),
    .Y(_04878_),
    .A2(_04864_));
 sg13g2_nand2_1 _12807_ (.Y(_04879_),
    .A(_03419_),
    .B(_03731_));
 sg13g2_o21ai_1 _12808_ (.B1(_04879_),
    .Y(_04880_),
    .A1(_03732_),
    .A2(net181));
 sg13g2_nor2_1 _12809_ (.A(_04867_),
    .B(_04865_),
    .Y(_04881_));
 sg13g2_a21oi_1 _12810_ (.A1(_03685_),
    .A2(_04880_),
    .Y(_04882_),
    .B1(_04881_));
 sg13g2_o21ai_1 _12811_ (.B1(_04882_),
    .Y(_04883_),
    .A1(_04869_),
    .A2(_04878_));
 sg13g2_nand2_1 _12812_ (.Y(_04884_),
    .A(_03419_),
    .B(_03761_));
 sg13g2_o21ai_1 _12813_ (.B1(_04884_),
    .Y(_04885_),
    .A1(_03762_),
    .A2(net181));
 sg13g2_inv_1 _12814_ (.Y(_04886_),
    .A(_04885_));
 sg13g2_nor2_1 _12815_ (.A(_04880_),
    .B(_03685_),
    .Y(_04887_));
 sg13g2_a21oi_1 _12816_ (.A1(_03651_),
    .A2(_04886_),
    .Y(_04888_),
    .B1(_04887_));
 sg13g2_nand2_1 _12817_ (.Y(_04889_),
    .A(_04883_),
    .B(_04888_));
 sg13g2_nand2_1 _12818_ (.Y(_04890_),
    .A(net181),
    .B(_03864_));
 sg13g2_o21ai_1 _12819_ (.B1(_04890_),
    .Y(_04891_),
    .A1(_03863_),
    .A2(net181));
 sg13g2_nor2_1 _12820_ (.A(_04886_),
    .B(_03651_),
    .Y(_04892_));
 sg13g2_a21oi_1 _12821_ (.A1(_03640_),
    .A2(_04891_),
    .Y(_04893_),
    .B1(_04892_));
 sg13g2_nand2_1 _12822_ (.Y(_04894_),
    .A(_04889_),
    .B(_04893_));
 sg13g2_nand2b_1 _12823_ (.Y(_04895_),
    .B(_03641_),
    .A_N(_04891_));
 sg13g2_nand2_1 _12824_ (.Y(_04896_),
    .A(_04894_),
    .B(_04895_));
 sg13g2_inv_1 _12825_ (.Y(_04897_),
    .A(\synth.voice.float_period[1][8] ));
 sg13g2_nor2_1 _12826_ (.A(_04897_),
    .B(_04210_),
    .Y(_04898_));
 sg13g2_a21oi_1 _12827_ (.A1(\synth.voice.float_period[0][8] ),
    .A2(_04210_),
    .Y(_04899_),
    .B1(_04898_));
 sg13g2_nand2_1 _12828_ (.Y(_04900_),
    .A(_03674_),
    .B(_04899_));
 sg13g2_nand2b_1 _12829_ (.Y(_04901_),
    .B(_03666_),
    .A_N(_04860_));
 sg13g2_o21ai_1 _12830_ (.B1(_04901_),
    .Y(_04902_),
    .A1(_04899_),
    .A2(_03674_));
 sg13g2_a21oi_1 _12831_ (.A1(_04896_),
    .A2(_04900_),
    .Y(_04903_),
    .B1(_04902_));
 sg13g2_nor2_1 _12832_ (.A(_04862_),
    .B(_04903_),
    .Y(_04904_));
 sg13g2_and2_1 _12833_ (.A(_04199_),
    .B(_04202_),
    .X(_04905_));
 sg13g2_nor3_1 _12834_ (.A(_03413_),
    .B(net182),
    .C(_04905_),
    .Y(_04906_));
 sg13g2_a21oi_1 _12835_ (.A1(_04904_),
    .A2(_04905_),
    .Y(_04907_),
    .B1(_04906_));
 sg13g2_buf_2 _12836_ (.A(\synth.voice.coeff_index[0] ),
    .X(_04908_));
 sg13g2_nand2_1 _12837_ (.Y(_04909_),
    .A(net182),
    .B(_04908_));
 sg13g2_nand2_1 _12838_ (.Y(_01201_),
    .A(_04907_),
    .B(_04909_));
 sg13g2_nor2_1 _12839_ (.A(net134),
    .B(_04229_),
    .Y(_04910_));
 sg13g2_nor2b_1 _12840_ (.A(_04790_),
    .B_N(_04910_),
    .Y(_04911_));
 sg13g2_nand2_1 _12841_ (.Y(_04912_),
    .A(_04911_),
    .B(net42));
 sg13g2_nand3_1 _12842_ (.B(\synth.voice.genblk4[1].next_state_scan[2] ),
    .C(net153),
    .A(_04795_),
    .Y(_04913_));
 sg13g2_nand2_1 _12843_ (.Y(_04914_),
    .A(net127),
    .B(\synth.voice.genblk4[1].next_state_scan[4] ));
 sg13g2_nand3_1 _12844_ (.B(_04913_),
    .C(_04914_),
    .A(_04912_),
    .Y(_01202_));
 sg13g2_nor2_1 _12845_ (.A(net134),
    .B(_04305_),
    .Y(_04915_));
 sg13g2_nor2b_1 _12846_ (.A(_04790_),
    .B_N(_04915_),
    .Y(_04916_));
 sg13g2_nand2_1 _12847_ (.Y(_04917_),
    .A(_04916_),
    .B(net42));
 sg13g2_nand3_1 _12848_ (.B(\synth.voice.genblk4[1].next_state_scan[3] ),
    .C(net153),
    .A(_04795_),
    .Y(_04918_));
 sg13g2_nand2_1 _12849_ (.Y(_04919_),
    .A(net127),
    .B(\synth.voice.genblk4[1].next_state_scan[5] ));
 sg13g2_nand3_1 _12850_ (.B(_04918_),
    .C(_04919_),
    .A(_04917_),
    .Y(_01203_));
 sg13g2_inv_1 _12851_ (.Y(_04920_),
    .A(\synth.voice.genblk4[1].next_state_scan[6] ));
 sg13g2_nor2_1 _12852_ (.A(_04920_),
    .B(net153),
    .Y(_04921_));
 sg13g2_nor2b_1 _12853_ (.A(net42),
    .B_N(\synth.voice.genblk4[1].next_state_scan[4] ),
    .Y(_04922_));
 sg13g2_nor2_1 _12854_ (.A(_04921_),
    .B(_04922_),
    .Y(_04923_));
 sg13g2_nor2_1 _12855_ (.A(net134),
    .B(_04795_),
    .Y(_04924_));
 sg13g2_nand2_1 _12856_ (.Y(_04925_),
    .A(_04204_),
    .B(_04372_));
 sg13g2_nand4_1 _12857_ (.B(_04831_),
    .C(net143),
    .A(_04199_),
    .Y(_04926_),
    .D(_04202_));
 sg13g2_nand3_1 _12858_ (.B(_04925_),
    .C(_04926_),
    .A(_04924_),
    .Y(_04927_));
 sg13g2_nand2_1 _12859_ (.Y(_01204_),
    .A(_04923_),
    .B(_04927_));
 sg13g2_nor2_1 _12860_ (.A(_04380_),
    .B(net153),
    .Y(_04928_));
 sg13g2_nor2_1 _12861_ (.A(_04732_),
    .B(net42),
    .Y(_04929_));
 sg13g2_nor2_1 _12862_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sg13g2_nand2b_1 _12863_ (.Y(_04931_),
    .B(_04204_),
    .A_N(_04710_));
 sg13g2_nand4_1 _12864_ (.B(_04833_),
    .C(net143),
    .A(_04199_),
    .Y(_04932_),
    .D(_04202_));
 sg13g2_nand3_1 _12865_ (.B(_04931_),
    .C(_04932_),
    .A(_04924_),
    .Y(_04933_));
 sg13g2_nand2_1 _12866_ (.Y(_01205_),
    .A(_04930_),
    .B(_04933_));
 sg13g2_inv_1 _12867_ (.Y(_04934_),
    .A(\synth.voice.genblk4[1].next_state_scan[8] ));
 sg13g2_nor2_1 _12868_ (.A(_04934_),
    .B(net153),
    .Y(_04935_));
 sg13g2_nor2_1 _12869_ (.A(_04920_),
    .B(net42),
    .Y(_04936_));
 sg13g2_nor2_1 _12870_ (.A(_04935_),
    .B(_04936_),
    .Y(_04937_));
 sg13g2_nand2_1 _12871_ (.Y(_04938_),
    .A(_04204_),
    .B(_04734_));
 sg13g2_nand4_1 _12872_ (.B(_04835_),
    .C(net143),
    .A(_04199_),
    .Y(_04939_),
    .D(_04202_));
 sg13g2_nand3_1 _12873_ (.B(_04938_),
    .C(_04939_),
    .A(_04924_),
    .Y(_04940_));
 sg13g2_nand2_1 _12874_ (.Y(_01206_),
    .A(_04937_),
    .B(_04940_));
 sg13g2_inv_1 _12875_ (.Y(_04941_),
    .A(\synth.voice.genblk4[1].next_state_scan[9] ));
 sg13g2_nor2_1 _12876_ (.A(_04941_),
    .B(net153),
    .Y(_04942_));
 sg13g2_nor2_1 _12877_ (.A(_04380_),
    .B(net42),
    .Y(_04943_));
 sg13g2_nor2_1 _12878_ (.A(_04942_),
    .B(_04943_),
    .Y(_04944_));
 sg13g2_nand2_1 _12879_ (.Y(_04945_),
    .A(_04204_),
    .B(_04751_));
 sg13g2_nand4_1 _12880_ (.B(_04837_),
    .C(net143),
    .A(_04199_),
    .Y(_04946_),
    .D(_04202_));
 sg13g2_nand3_1 _12881_ (.B(_04945_),
    .C(_04946_),
    .A(_04924_),
    .Y(_04947_));
 sg13g2_nand2_1 _12882_ (.Y(_01207_),
    .A(_04944_),
    .B(_04947_));
 sg13g2_inv_1 _12883_ (.Y(_04948_),
    .A(_03435_));
 sg13g2_nor2_2 _12884_ (.A(_04948_),
    .B(net134),
    .Y(_04949_));
 sg13g2_inv_1 _12885_ (.Y(_04950_),
    .A(_04949_));
 sg13g2_nand2_2 _12886_ (.Y(_04951_),
    .A(_04749_),
    .B(_03702_));
 sg13g2_nor2_2 _12887_ (.A(_03411_),
    .B(_04934_),
    .Y(_04952_));
 sg13g2_inv_1 _12888_ (.Y(_04953_),
    .A(_04952_));
 sg13g2_nand2_1 _12889_ (.Y(_04954_),
    .A(_04934_),
    .B(_03411_));
 sg13g2_nand3_1 _12890_ (.B(_04953_),
    .C(_04954_),
    .A(_04951_),
    .Y(_04955_));
 sg13g2_buf_1 _12891_ (.A(\synth.voice.genblk4[1].next_state_scan[10] ),
    .X(_04956_));
 sg13g2_nor2_1 _12892_ (.A(_03435_),
    .B(_04802_),
    .Y(_04957_));
 sg13g2_buf_2 _12893_ (.A(_04957_),
    .X(_04958_));
 sg13g2_a22oi_1 _12894_ (.Y(_04959_),
    .B1(\synth.voice.genblk4[1].next_state_scan[8] ),
    .B2(_04958_),
    .A2(_04802_),
    .A1(_04956_));
 sg13g2_o21ai_1 _12895_ (.B1(_04959_),
    .Y(_01208_),
    .A1(_04950_),
    .A2(_04955_));
 sg13g2_buf_1 _12896_ (.A(_00139_),
    .X(_04960_));
 sg13g2_xnor2_1 _12897_ (.Y(_04961_),
    .A(_04960_),
    .B(_04952_));
 sg13g2_nand3_1 _12898_ (.B(_04949_),
    .C(_04961_),
    .A(_04951_),
    .Y(_04962_));
 sg13g2_a22oi_1 _12899_ (.Y(_04963_),
    .B1(\synth.voice.genblk4[1].next_state_scan[9] ),
    .B2(_04958_),
    .A2(net127),
    .A1(\synth.voice.genblk4[1].next_state_scan[11] ));
 sg13g2_nand2_1 _12900_ (.Y(_01209_),
    .A(_04962_),
    .B(_04963_));
 sg13g2_nor2_1 _12901_ (.A(_04960_),
    .B(_04953_),
    .Y(_04964_));
 sg13g2_xnor2_1 _12902_ (.Y(_04965_),
    .A(_00140_),
    .B(_04964_));
 sg13g2_nand3_1 _12903_ (.B(_04949_),
    .C(_04965_),
    .A(_04951_),
    .Y(_04966_));
 sg13g2_a22oi_1 _12904_ (.Y(_04967_),
    .B1(_04956_),
    .B2(_04958_),
    .A2(net127),
    .A1(\synth.voice.genblk4[1].next_state_scan[12] ));
 sg13g2_nand2_1 _12905_ (.Y(_01210_),
    .A(_04966_),
    .B(_04967_));
 sg13g2_inv_1 _12906_ (.Y(_04968_),
    .A(_00141_));
 sg13g2_nand2_1 _12907_ (.Y(_04969_),
    .A(\synth.voice.genblk4[1].next_state_scan[9] ),
    .B(_04956_));
 sg13g2_inv_1 _12908_ (.Y(_04970_),
    .A(_04969_));
 sg13g2_nand2_1 _12909_ (.Y(_04971_),
    .A(_04970_),
    .B(_04952_));
 sg13g2_xnor2_1 _12910_ (.Y(_04972_),
    .A(_04968_),
    .B(_04971_));
 sg13g2_nand3_1 _12911_ (.B(_04949_),
    .C(_04972_),
    .A(_04951_),
    .Y(_04973_));
 sg13g2_a22oi_1 _12912_ (.Y(_04974_),
    .B1(\synth.voice.genblk4[1].next_state_scan[11] ),
    .B2(_04958_),
    .A2(_04803_),
    .A1(\synth.voice.genblk4[1].next_state_scan[13] ));
 sg13g2_nand2_1 _12913_ (.Y(_01211_),
    .A(_04973_),
    .B(_04974_));
 sg13g2_nand3_1 _12914_ (.B(_03668_),
    .C(_04196_),
    .A(_03584_),
    .Y(_04975_));
 sg13g2_nand2b_1 _12915_ (.Y(_04976_),
    .B(_04904_),
    .A_N(_04975_));
 sg13g2_nand3_1 _12916_ (.B(\synth.voice.delayed_p[1] ),
    .C(net189),
    .A(_04975_),
    .Y(_04977_));
 sg13g2_nand2_1 _12917_ (.Y(_04978_),
    .A(net182),
    .B(\synth.voice.coeff_index[1] ));
 sg13g2_nand3_1 _12918_ (.B(_04977_),
    .C(_04978_),
    .A(_04976_),
    .Y(_01212_));
 sg13g2_inv_1 _12919_ (.Y(_04979_),
    .A(_00142_));
 sg13g2_nand3_1 _12920_ (.B(_04956_),
    .C(\synth.voice.genblk4[1].next_state_scan[11] ),
    .A(_04964_),
    .Y(_04980_));
 sg13g2_xnor2_1 _12921_ (.Y(_04981_),
    .A(_04979_),
    .B(_04980_));
 sg13g2_nand3_1 _12922_ (.B(_04949_),
    .C(_04981_),
    .A(_04951_),
    .Y(_04982_));
 sg13g2_a22oi_1 _12923_ (.Y(_04983_),
    .B1(\synth.voice.genblk4[1].next_state_scan[12] ),
    .B2(_04958_),
    .A2(_04803_),
    .A1(_03370_));
 sg13g2_nand2_1 _12924_ (.Y(_01213_),
    .A(_04982_),
    .B(_04983_));
 sg13g2_nand4_1 _12925_ (.B(_04952_),
    .C(\synth.voice.genblk4[1].next_state_scan[11] ),
    .A(_04970_),
    .Y(_04984_),
    .D(\synth.voice.genblk4[1].next_state_scan[12] ));
 sg13g2_xor2_1 _12926_ (.B(_04984_),
    .A(_00143_),
    .X(_04985_));
 sg13g2_nand3_1 _12927_ (.B(_04949_),
    .C(_04985_),
    .A(_04951_),
    .Y(_04986_));
 sg13g2_a22oi_1 _12928_ (.Y(_04987_),
    .B1(\synth.voice.genblk4[1].next_state_scan[13] ),
    .B2(_04958_),
    .A2(net134),
    .A1(net401));
 sg13g2_nand2_1 _12929_ (.Y(_01214_),
    .A(_04986_),
    .B(_04987_));
 sg13g2_buf_1 _12930_ (.A(\synth.voice.a_sel_reg[3] ),
    .X(_04988_));
 sg13g2_buf_1 _12931_ (.A(_04988_),
    .X(_04989_));
 sg13g2_buf_1 _12932_ (.A(\synth.voice.a_sel_reg[2] ),
    .X(_04990_));
 sg13g2_buf_1 _12933_ (.A(_04990_),
    .X(_04991_));
 sg13g2_buf_1 _12934_ (.A(\synth.voice.a_sel_reg[1] ),
    .X(_04992_));
 sg13g2_nand2_1 _12935_ (.Y(_04993_),
    .A(\synth.voice.genblk4[2].next_state_scan[8] ),
    .B(net399));
 sg13g2_inv_1 _12936_ (.Y(_04994_),
    .A(_04993_));
 sg13g2_a221oi_1 _12937_ (.B2(\synth.controller.out[6] ),
    .C1(_04994_),
    .B1(net370),
    .A1(\synth.voice.genblk4[3].next_state_scan[12] ),
    .Y(_04995_),
    .A2(net371));
 sg13g2_buf_1 _12938_ (.A(_04995_),
    .X(_04996_));
 sg13g2_buf_2 _12939_ (.A(_00145_),
    .X(_04997_));
 sg13g2_inv_1 _12940_ (.Y(_04998_),
    .A(_04997_));
 sg13g2_buf_2 _12941_ (.A(\synth.voice.b_sel_reg[2] ),
    .X(_04999_));
 sg13g2_buf_2 _12942_ (.A(\synth.voice.b_sel_reg[0] ),
    .X(_05000_));
 sg13g2_nor2_1 _12943_ (.A(_04999_),
    .B(_05000_),
    .Y(_05001_));
 sg13g2_buf_1 _12944_ (.A(_05001_),
    .X(_05002_));
 sg13g2_inv_2 _12945_ (.Y(_05003_),
    .A(_05000_));
 sg13g2_inv_1 _12946_ (.Y(_05004_),
    .A(\synth.voice.genblk4[3].next_state_scan[1] ));
 sg13g2_buf_1 _12947_ (.A(\synth.voice.genblk4[4].next_state_scan[5] ),
    .X(_05005_));
 sg13g2_nand2_1 _12948_ (.Y(_05006_),
    .A(_04999_),
    .B(_05005_));
 sg13g2_o21ai_1 _12949_ (.B1(_05006_),
    .Y(_05007_),
    .A1(_05003_),
    .A2(_05004_));
 sg13g2_a21oi_1 _12950_ (.A1(\synth.voice.wave_reg[9] ),
    .A2(_05002_),
    .Y(_05008_),
    .B1(_05007_));
 sg13g2_xnor2_1 _12951_ (.Y(_05009_),
    .A(_04998_),
    .B(_05008_));
 sg13g2_buf_1 _12952_ (.A(\synth.voice.rshift_reg[0] ),
    .X(_05010_));
 sg13g2_buf_1 _12953_ (.A(_05010_),
    .X(_05011_));
 sg13g2_nand2_1 _12954_ (.Y(_05012_),
    .A(_05009_),
    .B(net369));
 sg13g2_buf_1 _12955_ (.A(_04998_),
    .X(_05013_));
 sg13g2_inv_1 _12956_ (.Y(_05014_),
    .A(\synth.voice.genblk4[3].next_state_scan[0] ));
 sg13g2_buf_1 _12957_ (.A(\synth.voice.genblk4[4].next_state_scan[4] ),
    .X(_05015_));
 sg13g2_nand2_1 _12958_ (.Y(_05016_),
    .A(_04999_),
    .B(_05015_));
 sg13g2_o21ai_1 _12959_ (.B1(_05016_),
    .Y(_05017_),
    .A1(_05003_),
    .A2(_05014_));
 sg13g2_a21oi_1 _12960_ (.A1(\synth.voice.wave_reg[8] ),
    .A2(_05002_),
    .Y(_05018_),
    .B1(_05017_));
 sg13g2_xnor2_1 _12961_ (.Y(_05019_),
    .A(net326),
    .B(_05018_));
 sg13g2_inv_1 _12962_ (.Y(_05020_),
    .A(_05010_));
 sg13g2_nand2_1 _12963_ (.Y(_05021_),
    .A(_05019_),
    .B(net368));
 sg13g2_buf_1 _12964_ (.A(\synth.voice.rshift_reg[1] ),
    .X(_05022_));
 sg13g2_inv_1 _12965_ (.Y(_05023_),
    .A(_05022_));
 sg13g2_nand3_1 _12966_ (.B(_05021_),
    .C(net367),
    .A(_05012_),
    .Y(_05024_));
 sg13g2_nor2_1 _12967_ (.A(_05023_),
    .B(_05009_),
    .Y(_05025_));
 sg13g2_inv_1 _12968_ (.Y(_05026_),
    .A(_05025_));
 sg13g2_nand2_1 _12969_ (.Y(_05027_),
    .A(_05024_),
    .B(_05026_));
 sg13g2_buf_1 _12970_ (.A(\synth.voice.rshift_reg[2] ),
    .X(_05028_));
 sg13g2_inv_1 _12971_ (.Y(_05029_),
    .A(net398));
 sg13g2_nand2_1 _12972_ (.Y(_05030_),
    .A(_05027_),
    .B(net366));
 sg13g2_inv_1 _12973_ (.Y(_05031_),
    .A(_05009_));
 sg13g2_nand2_2 _12974_ (.Y(_05032_),
    .A(_05031_),
    .B(net398));
 sg13g2_nand2_1 _12975_ (.Y(_05033_),
    .A(_05030_),
    .B(_05032_));
 sg13g2_buf_1 _12976_ (.A(\synth.voice.rshift_reg[3] ),
    .X(_05034_));
 sg13g2_buf_1 _12977_ (.A(_05034_),
    .X(_05035_));
 sg13g2_buf_1 _12978_ (.A(\synth.voice.zero_shifter_out_reg ),
    .X(_05036_));
 sg13g2_a21oi_1 _12979_ (.A1(_05033_),
    .A2(net365),
    .Y(_05037_),
    .B1(net397));
 sg13g2_buf_1 _12980_ (.A(_05010_),
    .X(_05038_));
 sg13g2_inv_2 _12981_ (.Y(_05039_),
    .A(_04999_));
 sg13g2_buf_1 _12982_ (.A(\synth.voice.scan_outs[4][1] ),
    .X(_05040_));
 sg13g2_inv_1 _12983_ (.Y(_05041_),
    .A(_05040_));
 sg13g2_nand2_1 _12984_ (.Y(_05042_),
    .A(_05000_),
    .B(\synth.voice.genblk4[2].next_state_scan[11] ));
 sg13g2_o21ai_1 _12985_ (.B1(_05042_),
    .Y(_05043_),
    .A1(_05039_),
    .A2(_05041_));
 sg13g2_a21oi_1 _12986_ (.A1(\synth.voice.wave_reg[3] ),
    .A2(net327),
    .Y(_05044_),
    .B1(_05043_));
 sg13g2_xnor2_1 _12987_ (.Y(_05045_),
    .A(net326),
    .B(_05044_));
 sg13g2_buf_2 _12988_ (.A(_04997_),
    .X(_05046_));
 sg13g2_buf_1 _12989_ (.A(\synth.voice.scan_outs[4][0] ),
    .X(_05047_));
 sg13g2_inv_1 _12990_ (.Y(_05048_),
    .A(_05047_));
 sg13g2_nand2_1 _12991_ (.Y(_05049_),
    .A(_05000_),
    .B(\synth.voice.genblk4[2].next_state_scan[10] ));
 sg13g2_o21ai_1 _12992_ (.B1(_05049_),
    .Y(_05050_),
    .A1(_05048_),
    .A2(_05039_));
 sg13g2_a21oi_1 _12993_ (.A1(\synth.voice.wave_reg[2] ),
    .A2(net327),
    .Y(_05051_),
    .B1(_05050_));
 sg13g2_xnor2_1 _12994_ (.Y(_05052_),
    .A(net363),
    .B(_05051_));
 sg13g2_nor2_1 _12995_ (.A(net369),
    .B(_05052_),
    .Y(_05053_));
 sg13g2_a21oi_1 _12996_ (.A1(net364),
    .A2(_05045_),
    .Y(_05054_),
    .B1(_05053_));
 sg13g2_buf_1 _12997_ (.A(_05022_),
    .X(_05055_));
 sg13g2_nand2_1 _12998_ (.Y(_05056_),
    .A(_05054_),
    .B(_05055_));
 sg13g2_inv_1 _12999_ (.Y(_05057_),
    .A(\synth.voice.genblk4[3].next_state_scan[13] ));
 sg13g2_nand2_1 _13000_ (.Y(_05058_),
    .A(_05000_),
    .B(\synth.voice.genblk4[2].next_state_scan[9] ));
 sg13g2_o21ai_1 _13001_ (.B1(_05058_),
    .Y(_05059_),
    .A1(_05039_),
    .A2(_05057_));
 sg13g2_a21oi_1 _13002_ (.A1(\synth.voice.wave_reg[1] ),
    .A2(net327),
    .Y(_05060_),
    .B1(_05059_));
 sg13g2_xnor2_1 _13003_ (.Y(_05061_),
    .A(_05046_),
    .B(_05060_));
 sg13g2_nand2_1 _13004_ (.Y(_05062_),
    .A(_05061_),
    .B(net369));
 sg13g2_inv_1 _13005_ (.Y(_05063_),
    .A(\synth.voice.genblk4[3].next_state_scan[12] ));
 sg13g2_nand2_1 _13006_ (.Y(_05064_),
    .A(_05000_),
    .B(\synth.voice.genblk4[2].next_state_scan[8] ));
 sg13g2_o21ai_1 _13007_ (.B1(_05064_),
    .Y(_05065_),
    .A1(_05039_),
    .A2(_05063_));
 sg13g2_a21oi_1 _13008_ (.A1(\synth.voice.wave_reg[0] ),
    .A2(net327),
    .Y(_05066_),
    .B1(_05065_));
 sg13g2_xnor2_1 _13009_ (.Y(_05067_),
    .A(_05046_),
    .B(_05066_));
 sg13g2_buf_1 _13010_ (.A(net368),
    .X(_05068_));
 sg13g2_nand2_1 _13011_ (.Y(_05069_),
    .A(_05067_),
    .B(net325));
 sg13g2_nand2_1 _13012_ (.Y(_05070_),
    .A(_05062_),
    .B(_05069_));
 sg13g2_buf_1 _13013_ (.A(net367),
    .X(_05071_));
 sg13g2_nand2_1 _13014_ (.Y(_05072_),
    .A(_05070_),
    .B(_05071_));
 sg13g2_buf_1 _13015_ (.A(net366),
    .X(_05073_));
 sg13g2_nand3_1 _13016_ (.B(_05072_),
    .C(net323),
    .A(_05056_),
    .Y(_05074_));
 sg13g2_inv_1 _13017_ (.Y(_05075_),
    .A(\synth.voice.genblk4[4].next_state_scan[1] ));
 sg13g2_nand2_1 _13018_ (.Y(_05076_),
    .A(_05000_),
    .B(\synth.voice.genblk4[2].next_state_scan[13] ));
 sg13g2_o21ai_1 _13019_ (.B1(_05076_),
    .Y(_05077_),
    .A1(_05039_),
    .A2(_05075_));
 sg13g2_a21oi_1 _13020_ (.A1(\synth.voice.wave_reg[5] ),
    .A2(net327),
    .Y(_05078_),
    .B1(_05077_));
 sg13g2_xnor2_1 _13021_ (.Y(_05079_),
    .A(_04997_),
    .B(_05078_));
 sg13g2_inv_1 _13022_ (.Y(_05080_),
    .A(_05079_));
 sg13g2_nand2_1 _13023_ (.Y(_05081_),
    .A(_05080_),
    .B(net364));
 sg13g2_inv_1 _13024_ (.Y(_05082_),
    .A(\synth.voice.genblk4[4].next_state_scan[0] ));
 sg13g2_nand2_1 _13025_ (.Y(_05083_),
    .A(_05000_),
    .B(\synth.voice.genblk4[2].next_state_scan[12] ));
 sg13g2_o21ai_1 _13026_ (.B1(_05083_),
    .Y(_05084_),
    .A1(_05039_),
    .A2(_05082_));
 sg13g2_a21oi_1 _13027_ (.A1(\synth.voice.wave_reg[4] ),
    .A2(net327),
    .Y(_05085_),
    .B1(_05084_));
 sg13g2_xnor2_1 _13028_ (.Y(_05086_),
    .A(net326),
    .B(_05085_));
 sg13g2_nand2_1 _13029_ (.Y(_05087_),
    .A(_05086_),
    .B(_05068_));
 sg13g2_nand3_1 _13030_ (.B(net367),
    .C(_05087_),
    .A(_05081_),
    .Y(_05088_));
 sg13g2_inv_1 _13031_ (.Y(_05089_),
    .A(\synth.voice.scan_outs[3][0] ));
 sg13g2_buf_1 _13032_ (.A(\synth.voice.genblk4[4].next_state_scan[2] ),
    .X(_05090_));
 sg13g2_nand2_1 _13033_ (.Y(_05091_),
    .A(_04999_),
    .B(_05090_));
 sg13g2_o21ai_1 _13034_ (.B1(_05091_),
    .Y(_05092_),
    .A1(_05089_),
    .A2(_05003_));
 sg13g2_a21oi_1 _13035_ (.A1(\synth.voice.wave_reg[6] ),
    .A2(net327),
    .Y(_05093_),
    .B1(_05092_));
 sg13g2_xnor2_1 _13036_ (.Y(_05094_),
    .A(net326),
    .B(_05093_));
 sg13g2_nand2_1 _13037_ (.Y(_05095_),
    .A(_05094_),
    .B(net368));
 sg13g2_inv_1 _13038_ (.Y(_05096_),
    .A(\synth.voice.scan_outs[3][1] ));
 sg13g2_nand2_1 _13039_ (.Y(_05097_),
    .A(_04999_),
    .B(\synth.voice.genblk4[4].next_state_scan[3] ));
 sg13g2_o21ai_1 _13040_ (.B1(_05097_),
    .Y(_05098_),
    .A1(_05003_),
    .A2(_05096_));
 sg13g2_a21oi_1 _13041_ (.A1(\synth.voice.wave_reg[7] ),
    .A2(net327),
    .Y(_05099_),
    .B1(_05098_));
 sg13g2_xnor2_1 _13042_ (.Y(_05100_),
    .A(net326),
    .B(_05099_));
 sg13g2_nand2_1 _13043_ (.Y(_05101_),
    .A(_05100_),
    .B(net369));
 sg13g2_nand3_1 _13044_ (.B(_05101_),
    .C(net362),
    .A(_05095_),
    .Y(_05102_));
 sg13g2_buf_1 _13045_ (.A(net398),
    .X(_05103_));
 sg13g2_nand3_1 _13046_ (.B(_05102_),
    .C(net361),
    .A(_05088_),
    .Y(_05104_));
 sg13g2_inv_1 _13047_ (.Y(_05105_),
    .A(_05034_));
 sg13g2_nand3_1 _13048_ (.B(_05104_),
    .C(net360),
    .A(_05074_),
    .Y(_05106_));
 sg13g2_nand2_1 _13049_ (.Y(_05107_),
    .A(_05037_),
    .B(_05106_));
 sg13g2_nor2_1 _13050_ (.A(_04996_),
    .B(_05107_),
    .Y(_05108_));
 sg13g2_buf_1 _13051_ (.A(_04988_),
    .X(_05109_));
 sg13g2_nand2_1 _13052_ (.Y(_05110_),
    .A(\synth.voice.genblk4[2].next_state_scan[7] ),
    .B(net399));
 sg13g2_inv_1 _13053_ (.Y(_05111_),
    .A(_05110_));
 sg13g2_a221oi_1 _13054_ (.B2(\synth.controller.out[5] ),
    .C1(_05111_),
    .B1(net370),
    .A1(\synth.voice.genblk4[3].next_state_scan[11] ),
    .Y(_05112_),
    .A2(net359));
 sg13g2_xnor2_1 _13055_ (.Y(_05113_),
    .A(net363),
    .B(_05018_));
 sg13g2_nand2_1 _13056_ (.Y(_05114_),
    .A(_05113_),
    .B(_05010_));
 sg13g2_xnor2_1 _13057_ (.Y(_05115_),
    .A(_04997_),
    .B(_05099_));
 sg13g2_nand2_1 _13058_ (.Y(_05116_),
    .A(_05115_),
    .B(net368));
 sg13g2_nand2_1 _13059_ (.Y(_05117_),
    .A(_05114_),
    .B(_05116_));
 sg13g2_nand2_1 _13060_ (.Y(_05118_),
    .A(_05117_),
    .B(net367));
 sg13g2_nand2_1 _13061_ (.Y(_05119_),
    .A(_05118_),
    .B(_05026_));
 sg13g2_nand2_1 _13062_ (.Y(_05120_),
    .A(_05119_),
    .B(net366));
 sg13g2_a21oi_1 _13063_ (.A1(_05120_),
    .A2(_05032_),
    .Y(_05121_),
    .B1(net360));
 sg13g2_nor2_1 _13064_ (.A(net368),
    .B(_05094_),
    .Y(_05122_));
 sg13g2_nor2_1 _13065_ (.A(net364),
    .B(_05080_),
    .Y(_05123_));
 sg13g2_o21ai_1 _13066_ (.B1(net362),
    .Y(_05124_),
    .A1(_05122_),
    .A2(_05123_));
 sg13g2_nand2_1 _13067_ (.Y(_05125_),
    .A(_05045_),
    .B(_05068_));
 sg13g2_nand2_1 _13068_ (.Y(_05126_),
    .A(_05086_),
    .B(_05011_));
 sg13g2_nand3_1 _13069_ (.B(_05126_),
    .C(net367),
    .A(_05125_),
    .Y(_05127_));
 sg13g2_nand3_1 _13070_ (.B(net398),
    .C(_05127_),
    .A(_05124_),
    .Y(_05128_));
 sg13g2_inv_1 _13071_ (.Y(_05129_),
    .A(_05061_));
 sg13g2_nand2_1 _13072_ (.Y(_05130_),
    .A(_05129_),
    .B(net325));
 sg13g2_xnor2_1 _13073_ (.Y(_05131_),
    .A(net326),
    .B(_05051_));
 sg13g2_nand2_1 _13074_ (.Y(_05132_),
    .A(_05131_),
    .B(net364));
 sg13g2_nand3_1 _13075_ (.B(_05132_),
    .C(_05055_),
    .A(_05130_),
    .Y(_05133_));
 sg13g2_nand2_1 _13076_ (.Y(_05134_),
    .A(_05067_),
    .B(_05011_));
 sg13g2_buf_1 _13077_ (.A(_05003_),
    .X(_05135_));
 sg13g2_inv_1 _13078_ (.Y(_05136_),
    .A(\synth.voice.genblk4[2].next_state_scan[7] ));
 sg13g2_buf_1 _13079_ (.A(_04999_),
    .X(_05137_));
 sg13g2_nand2_1 _13080_ (.Y(_05138_),
    .A(net358),
    .B(\synth.voice.genblk4[3].next_state_scan[11] ));
 sg13g2_o21ai_1 _13081_ (.B1(_05138_),
    .Y(_05139_),
    .A1(net322),
    .A2(_05136_));
 sg13g2_xnor2_1 _13082_ (.Y(_05140_),
    .A(net326),
    .B(_05139_));
 sg13g2_nand2_1 _13083_ (.Y(_05141_),
    .A(_05140_),
    .B(net368));
 sg13g2_nand2_1 _13084_ (.Y(_05142_),
    .A(_05134_),
    .B(_05141_));
 sg13g2_nand2_1 _13085_ (.Y(_05143_),
    .A(_05142_),
    .B(net367));
 sg13g2_nand3_1 _13086_ (.B(_05143_),
    .C(net366),
    .A(_05133_),
    .Y(_05144_));
 sg13g2_nand3_1 _13087_ (.B(net360),
    .C(_05144_),
    .A(_05128_),
    .Y(_05145_));
 sg13g2_inv_1 _13088_ (.Y(_05146_),
    .A(net397));
 sg13g2_nand3b_1 _13089_ (.B(_05145_),
    .C(_05146_),
    .Y(_05147_),
    .A_N(_05121_));
 sg13g2_nor2_1 _13090_ (.A(_05112_),
    .B(_05147_),
    .Y(_05148_));
 sg13g2_nand2_1 _13091_ (.Y(_05149_),
    .A(_05107_),
    .B(_04996_));
 sg13g2_nand2_1 _13092_ (.Y(_05150_),
    .A(_05148_),
    .B(_05149_));
 sg13g2_nand2b_1 _13093_ (.Y(_05151_),
    .B(_05150_),
    .A_N(_05108_));
 sg13g2_buf_1 _13094_ (.A(_04992_),
    .X(_05152_));
 sg13g2_nand2_1 _13095_ (.Y(_05153_),
    .A(\synth.voice.genblk4[3].next_state_scan[9] ),
    .B(net359));
 sg13g2_inv_1 _13096_ (.Y(_05154_),
    .A(_05153_));
 sg13g2_a221oi_1 _13097_ (.B2(\synth.controller.out[3] ),
    .C1(_05154_),
    .B1(net370),
    .A1(\synth.voice.genblk4[2].next_state_scan[5] ),
    .Y(_05155_),
    .A2(_05152_));
 sg13g2_buf_1 _13098_ (.A(_05155_),
    .X(_05156_));
 sg13g2_a21oi_1 _13099_ (.A1(net325),
    .A2(_05079_),
    .Y(_05157_),
    .B1(_05122_));
 sg13g2_nand2_1 _13100_ (.Y(_05158_),
    .A(_05157_),
    .B(net367));
 sg13g2_nand3_1 _13101_ (.B(_05116_),
    .C(net362),
    .A(_05114_),
    .Y(_05159_));
 sg13g2_nand3_1 _13102_ (.B(net366),
    .C(_05159_),
    .A(_05158_),
    .Y(_05160_));
 sg13g2_nand2_1 _13103_ (.Y(_05161_),
    .A(_05160_),
    .B(_05032_));
 sg13g2_nand2_1 _13104_ (.Y(_05162_),
    .A(_05161_),
    .B(net365));
 sg13g2_nand3_1 _13105_ (.B(_05132_),
    .C(net324),
    .A(_05130_),
    .Y(_05163_));
 sg13g2_buf_1 _13106_ (.A(_05022_),
    .X(_05164_));
 sg13g2_nand3_1 _13107_ (.B(_05126_),
    .C(net356),
    .A(_05125_),
    .Y(_05165_));
 sg13g2_nand3_1 _13108_ (.B(_05165_),
    .C(net398),
    .A(_05163_),
    .Y(_05166_));
 sg13g2_nand2_1 _13109_ (.Y(_05167_),
    .A(_05142_),
    .B(_05164_));
 sg13g2_inv_1 _13110_ (.Y(_05168_),
    .A(\synth.voice.genblk4[2].next_state_scan[6] ));
 sg13g2_nand2_1 _13111_ (.Y(_05169_),
    .A(net358),
    .B(\synth.voice.genblk4[3].next_state_scan[10] ));
 sg13g2_o21ai_1 _13112_ (.B1(_05169_),
    .Y(_05170_),
    .A1(net322),
    .A2(_05168_));
 sg13g2_xnor2_1 _13113_ (.Y(_05171_),
    .A(net363),
    .B(_05170_));
 sg13g2_inv_1 _13114_ (.Y(_05172_),
    .A(\synth.voice.genblk4[2].next_state_scan[5] ));
 sg13g2_nand2_1 _13115_ (.Y(_05173_),
    .A(net358),
    .B(\synth.voice.genblk4[3].next_state_scan[9] ));
 sg13g2_o21ai_1 _13116_ (.B1(_05173_),
    .Y(_05174_),
    .A1(net322),
    .A2(_05172_));
 sg13g2_xnor2_1 _13117_ (.Y(_05175_),
    .A(_04998_),
    .B(_05174_));
 sg13g2_nor2_1 _13118_ (.A(_05010_),
    .B(_05175_),
    .Y(_05176_));
 sg13g2_a21oi_1 _13119_ (.A1(net369),
    .A2(_05171_),
    .Y(_05177_),
    .B1(_05176_));
 sg13g2_nand2_1 _13120_ (.Y(_05178_),
    .A(_05177_),
    .B(net324));
 sg13g2_nand3_1 _13121_ (.B(net323),
    .C(_05178_),
    .A(_05167_),
    .Y(_05179_));
 sg13g2_nand3_1 _13122_ (.B(_05179_),
    .C(net360),
    .A(_05166_),
    .Y(_05180_));
 sg13g2_nand3_1 _13123_ (.B(_05146_),
    .C(_05180_),
    .A(_05162_),
    .Y(_05181_));
 sg13g2_nor2_1 _13124_ (.A(_05156_),
    .B(_05181_),
    .Y(_05182_));
 sg13g2_nand3_1 _13125_ (.B(_05021_),
    .C(_05022_),
    .A(_05012_),
    .Y(_05183_));
 sg13g2_nand3_1 _13126_ (.B(_05101_),
    .C(net367),
    .A(_05095_),
    .Y(_05184_));
 sg13g2_nand2_1 _13127_ (.Y(_05185_),
    .A(_05183_),
    .B(_05184_));
 sg13g2_nand2_1 _13128_ (.Y(_05186_),
    .A(_05185_),
    .B(net366));
 sg13g2_nand2_1 _13129_ (.Y(_05187_),
    .A(_05186_),
    .B(_05032_));
 sg13g2_a21oi_1 _13130_ (.A1(_05187_),
    .A2(net365),
    .Y(_05188_),
    .B1(net397));
 sg13g2_nand2_1 _13131_ (.Y(_05189_),
    .A(_05054_),
    .B(net324));
 sg13g2_nand3_1 _13132_ (.B(net356),
    .C(_05087_),
    .A(_05081_),
    .Y(_05190_));
 sg13g2_nand3_1 _13133_ (.B(net361),
    .C(_05190_),
    .A(_05189_),
    .Y(_05191_));
 sg13g2_nand3_1 _13134_ (.B(_05069_),
    .C(net362),
    .A(_05062_),
    .Y(_05192_));
 sg13g2_nor2_1 _13135_ (.A(net368),
    .B(_05140_),
    .Y(_05193_));
 sg13g2_a21oi_1 _13136_ (.A1(net325),
    .A2(_05171_),
    .Y(_05194_),
    .B1(_05193_));
 sg13g2_nand2b_1 _13137_ (.Y(_05195_),
    .B(net324),
    .A_N(_05194_));
 sg13g2_nand2_1 _13138_ (.Y(_05196_),
    .A(_05192_),
    .B(_05195_));
 sg13g2_nand2_1 _13139_ (.Y(_05197_),
    .A(_05196_),
    .B(net323));
 sg13g2_buf_1 _13140_ (.A(_05105_),
    .X(_05198_));
 sg13g2_nand3_1 _13141_ (.B(_05197_),
    .C(_05198_),
    .A(_05191_),
    .Y(_05199_));
 sg13g2_nand2_1 _13142_ (.Y(_05200_),
    .A(_05188_),
    .B(_05199_));
 sg13g2_buf_1 _13143_ (.A(_04990_),
    .X(_05201_));
 sg13g2_nand2_1 _13144_ (.Y(_05202_),
    .A(\synth.voice.genblk4[3].next_state_scan[10] ),
    .B(net359));
 sg13g2_inv_1 _13145_ (.Y(_05203_),
    .A(_05202_));
 sg13g2_a221oi_1 _13146_ (.B2(\synth.controller.out[4] ),
    .C1(_05203_),
    .B1(_05201_),
    .A1(\synth.voice.genblk4[2].next_state_scan[6] ),
    .Y(_05204_),
    .A2(net357));
 sg13g2_buf_1 _13147_ (.A(_05204_),
    .X(_05205_));
 sg13g2_nand2_1 _13148_ (.Y(_05206_),
    .A(_05200_),
    .B(_05205_));
 sg13g2_nor2_1 _13149_ (.A(_05205_),
    .B(_05200_),
    .Y(_05207_));
 sg13g2_a21oi_1 _13150_ (.A1(_05182_),
    .A2(_05206_),
    .Y(_05208_),
    .B1(_05207_));
 sg13g2_inv_1 _13151_ (.Y(_05209_),
    .A(_05208_));
 sg13g2_xnor2_1 _13152_ (.Y(_05210_),
    .A(_04996_),
    .B(_05107_));
 sg13g2_nand2_1 _13153_ (.Y(_05211_),
    .A(_05147_),
    .B(_05112_));
 sg13g2_nand2_1 _13154_ (.Y(_05212_),
    .A(_05145_),
    .B(_05146_));
 sg13g2_nor2_1 _13155_ (.A(_05121_),
    .B(_05212_),
    .Y(_05213_));
 sg13g2_nand2b_1 _13156_ (.Y(_05214_),
    .B(_05213_),
    .A_N(_05112_));
 sg13g2_nand2_1 _13157_ (.Y(_05215_),
    .A(_05211_),
    .B(_05214_));
 sg13g2_nor2_1 _13158_ (.A(_05210_),
    .B(_05215_),
    .Y(_05216_));
 sg13g2_nand2_1 _13159_ (.Y(_05217_),
    .A(_05209_),
    .B(_05216_));
 sg13g2_nand2b_1 _13160_ (.Y(_05218_),
    .B(_05217_),
    .A_N(_05151_));
 sg13g2_xnor2_1 _13161_ (.Y(_05219_),
    .A(_05205_),
    .B(_05200_));
 sg13g2_xnor2_1 _13162_ (.Y(_05220_),
    .A(_05156_),
    .B(_05181_));
 sg13g2_nor2_1 _13163_ (.A(_05219_),
    .B(_05220_),
    .Y(_05221_));
 sg13g2_nand2_1 _13164_ (.Y(_05222_),
    .A(_05216_),
    .B(_05221_));
 sg13g2_inv_1 _13165_ (.Y(_05223_),
    .A(\synth.voice.genblk4[2].next_state_scan[2] ));
 sg13g2_nand2_1 _13166_ (.Y(_05224_),
    .A(net358),
    .B(\synth.voice.genblk4[3].next_state_scan[6] ));
 sg13g2_o21ai_1 _13167_ (.B1(_05224_),
    .Y(_05225_),
    .A1(net322),
    .A2(_05223_));
 sg13g2_xnor2_1 _13168_ (.Y(_05226_),
    .A(net363),
    .B(_05225_));
 sg13g2_inv_1 _13169_ (.Y(_05227_),
    .A(\synth.voice.genblk4[2].next_state_scan[1] ));
 sg13g2_nand2_1 _13170_ (.Y(_05228_),
    .A(net358),
    .B(\synth.voice.genblk4[3].next_state_scan[5] ));
 sg13g2_o21ai_1 _13171_ (.B1(_05228_),
    .Y(_05229_),
    .A1(net322),
    .A2(_05227_));
 sg13g2_xnor2_1 _13172_ (.Y(_05230_),
    .A(net326),
    .B(_05229_));
 sg13g2_nor2_1 _13173_ (.A(net369),
    .B(_05230_),
    .Y(_05231_));
 sg13g2_a21oi_1 _13174_ (.A1(net364),
    .A2(_05226_),
    .Y(_05232_),
    .B1(_05231_));
 sg13g2_nor2_1 _13175_ (.A(net356),
    .B(_05232_),
    .Y(_05233_));
 sg13g2_inv_1 _13176_ (.Y(_05234_),
    .A(\synth.voice.genblk4[2].next_state_scan[4] ));
 sg13g2_nand2_1 _13177_ (.Y(_05235_),
    .A(net358),
    .B(\synth.voice.genblk4[3].next_state_scan[8] ));
 sg13g2_o21ai_1 _13178_ (.B1(_05235_),
    .Y(_05236_),
    .A1(_05135_),
    .A2(_05234_));
 sg13g2_xnor2_1 _13179_ (.Y(_05237_),
    .A(net363),
    .B(_05236_));
 sg13g2_inv_1 _13180_ (.Y(_05238_),
    .A(\synth.voice.genblk4[2].next_state_scan[3] ));
 sg13g2_nand2_1 _13181_ (.Y(_05239_),
    .A(_05137_),
    .B(\synth.voice.genblk4[3].next_state_scan[7] ));
 sg13g2_o21ai_1 _13182_ (.B1(_05239_),
    .Y(_05240_),
    .A1(net322),
    .A2(_05238_));
 sg13g2_xnor2_1 _13183_ (.Y(_05241_),
    .A(_05013_),
    .B(_05240_));
 sg13g2_nor2_1 _13184_ (.A(net369),
    .B(_05241_),
    .Y(_05242_));
 sg13g2_a21oi_1 _13185_ (.A1(net369),
    .A2(_05237_),
    .Y(_05243_),
    .B1(_05242_));
 sg13g2_nand2b_1 _13186_ (.Y(_05244_),
    .B(net356),
    .A_N(_05243_));
 sg13g2_nand2b_1 _13187_ (.Y(_05245_),
    .B(_05244_),
    .A_N(_05233_));
 sg13g2_a21oi_1 _13188_ (.A1(_05245_),
    .A2(net323),
    .Y(_05246_),
    .B1(_05034_));
 sg13g2_nand3_1 _13189_ (.B(net361),
    .C(_05178_),
    .A(_05167_),
    .Y(_05247_));
 sg13g2_a21oi_1 _13190_ (.A1(_05246_),
    .A2(_05247_),
    .Y(_05248_),
    .B1(net397));
 sg13g2_nand2_1 _13191_ (.Y(_05249_),
    .A(_05158_),
    .B(_05159_));
 sg13g2_nand2_1 _13192_ (.Y(_05250_),
    .A(_05249_),
    .B(net361));
 sg13g2_nand3_1 _13193_ (.B(_05165_),
    .C(net323),
    .A(_05163_),
    .Y(_05251_));
 sg13g2_nand3_1 _13194_ (.B(net365),
    .C(_05251_),
    .A(_05250_),
    .Y(_05252_));
 sg13g2_nand2_1 _13195_ (.Y(_05253_),
    .A(\synth.voice.genblk4[3].next_state_scan[5] ),
    .B(net359));
 sg13g2_nand2_1 _13196_ (.Y(_05254_),
    .A(net370),
    .B(\synth.voice.acc[3] ));
 sg13g2_nand2_1 _13197_ (.Y(_05255_),
    .A(\synth.voice.genblk4[2].next_state_scan[1] ),
    .B(net399));
 sg13g2_nand3_1 _13198_ (.B(_05254_),
    .C(_05255_),
    .A(_05253_),
    .Y(_05256_));
 sg13g2_nand3_1 _13199_ (.B(_05252_),
    .C(_05256_),
    .A(_05248_),
    .Y(_05257_));
 sg13g2_buf_1 _13200_ (.A(_05257_),
    .X(_05258_));
 sg13g2_inv_1 _13201_ (.Y(_05259_),
    .A(_05258_));
 sg13g2_nand3_1 _13202_ (.B(_05195_),
    .C(net361),
    .A(_05192_),
    .Y(_05260_));
 sg13g2_nor2_1 _13203_ (.A(_05038_),
    .B(_05226_),
    .Y(_05261_));
 sg13g2_a21oi_1 _13204_ (.A1(_05038_),
    .A2(_05241_),
    .Y(_05262_),
    .B1(_05261_));
 sg13g2_nor2_1 _13205_ (.A(net368),
    .B(_05175_),
    .Y(_05263_));
 sg13g2_a21oi_1 _13206_ (.A1(net325),
    .A2(_05237_),
    .Y(_05264_),
    .B1(_05263_));
 sg13g2_nor2_1 _13207_ (.A(_05071_),
    .B(_05264_),
    .Y(_05265_));
 sg13g2_a21oi_1 _13208_ (.A1(net324),
    .A2(_05262_),
    .Y(_05266_),
    .B1(_05265_));
 sg13g2_nand2_1 _13209_ (.Y(_05267_),
    .A(_05266_),
    .B(net323));
 sg13g2_nand2_1 _13210_ (.Y(_05268_),
    .A(_05260_),
    .B(_05267_));
 sg13g2_a21oi_1 _13211_ (.A1(_05268_),
    .A2(_05198_),
    .Y(_05269_),
    .B1(net397));
 sg13g2_nand3_1 _13212_ (.B(net323),
    .C(_05190_),
    .A(_05189_),
    .Y(_05270_));
 sg13g2_nand3_1 _13213_ (.B(_05184_),
    .C(net361),
    .A(_05183_),
    .Y(_05271_));
 sg13g2_nand3_1 _13214_ (.B(_05271_),
    .C(net365),
    .A(_05270_),
    .Y(_05272_));
 sg13g2_nand2_1 _13215_ (.Y(_05273_),
    .A(_05269_),
    .B(_05272_));
 sg13g2_nand2_1 _13216_ (.Y(_05274_),
    .A(\synth.voice.genblk4[2].next_state_scan[2] ),
    .B(net357));
 sg13g2_inv_1 _13217_ (.Y(_05275_),
    .A(_05274_));
 sg13g2_a221oi_1 _13218_ (.B2(\synth.controller.out[0] ),
    .C1(_05275_),
    .B1(net355),
    .A1(\synth.voice.genblk4[3].next_state_scan[6] ),
    .Y(_05276_),
    .A2(_04989_));
 sg13g2_buf_1 _13219_ (.A(_05276_),
    .X(_05277_));
 sg13g2_nand2_1 _13220_ (.Y(_05278_),
    .A(_05273_),
    .B(_05277_));
 sg13g2_nor2_1 _13221_ (.A(_05277_),
    .B(_05273_),
    .Y(_05279_));
 sg13g2_a21oi_1 _13222_ (.A1(_05259_),
    .A2(_05278_),
    .Y(_05280_),
    .B1(_05279_));
 sg13g2_nand2_1 _13223_ (.Y(_05281_),
    .A(\synth.voice.genblk4[2].next_state_scan[3] ),
    .B(\synth.voice.a_sel_reg[1] ));
 sg13g2_inv_1 _13224_ (.Y(_05282_),
    .A(_05281_));
 sg13g2_a221oi_1 _13225_ (.B2(\synth.controller.out[1] ),
    .C1(_05282_),
    .B1(net370),
    .A1(\synth.voice.genblk4[3].next_state_scan[7] ),
    .Y(_05283_),
    .A2(net359));
 sg13g2_buf_1 _13226_ (.A(_05283_),
    .X(_05284_));
 sg13g2_nor2_1 _13227_ (.A(net362),
    .B(_05243_),
    .Y(_05285_));
 sg13g2_nand2b_1 _13228_ (.Y(_05286_),
    .B(net362),
    .A_N(_05177_));
 sg13g2_nand2b_1 _13229_ (.Y(_05287_),
    .B(_05286_),
    .A_N(_05285_));
 sg13g2_a21oi_1 _13230_ (.A1(_05287_),
    .A2(_05073_),
    .Y(_05288_),
    .B1(_05034_));
 sg13g2_nand3_1 _13231_ (.B(_05143_),
    .C(_05028_),
    .A(_05133_),
    .Y(_05289_));
 sg13g2_a21oi_1 _13232_ (.A1(_05288_),
    .A2(_05289_),
    .Y(_05290_),
    .B1(_05036_));
 sg13g2_nand3_1 _13233_ (.B(net366),
    .C(_05127_),
    .A(_05124_),
    .Y(_05291_));
 sg13g2_nand3_1 _13234_ (.B(net398),
    .C(_05026_),
    .A(_05118_),
    .Y(_05292_));
 sg13g2_nand3_1 _13235_ (.B(_05292_),
    .C(_05034_),
    .A(_05291_),
    .Y(_05293_));
 sg13g2_nand2_1 _13236_ (.Y(_05294_),
    .A(_05290_),
    .B(_05293_));
 sg13g2_xnor2_1 _13237_ (.Y(_05295_),
    .A(_05284_),
    .B(_05294_));
 sg13g2_nand2_1 _13238_ (.Y(_05296_),
    .A(\synth.voice.genblk4[2].next_state_scan[4] ),
    .B(_04992_));
 sg13g2_inv_1 _13239_ (.Y(_05297_),
    .A(_05296_));
 sg13g2_a221oi_1 _13240_ (.B2(\synth.controller.out[2] ),
    .C1(_05297_),
    .B1(net370),
    .A1(\synth.voice.genblk4[3].next_state_scan[8] ),
    .Y(_05298_),
    .A2(_05109_));
 sg13g2_nand3_1 _13241_ (.B(_05072_),
    .C(net398),
    .A(_05056_),
    .Y(_05299_));
 sg13g2_nand2_1 _13242_ (.Y(_05300_),
    .A(_05194_),
    .B(net362));
 sg13g2_nand2_1 _13243_ (.Y(_05301_),
    .A(_05264_),
    .B(net324));
 sg13g2_nand3_1 _13244_ (.B(_05301_),
    .C(_05029_),
    .A(_05300_),
    .Y(_05302_));
 sg13g2_nand3_1 _13245_ (.B(net360),
    .C(_05302_),
    .A(_05299_),
    .Y(_05303_));
 sg13g2_nand3_1 _13246_ (.B(_05102_),
    .C(net366),
    .A(_05088_),
    .Y(_05304_));
 sg13g2_nand3_1 _13247_ (.B(net398),
    .C(_05026_),
    .A(_05024_),
    .Y(_05305_));
 sg13g2_nand3_1 _13248_ (.B(_05305_),
    .C(_05034_),
    .A(_05304_),
    .Y(_05306_));
 sg13g2_nand2_1 _13249_ (.Y(_05307_),
    .A(_05303_),
    .B(_05306_));
 sg13g2_nor2_1 _13250_ (.A(_05036_),
    .B(_05307_),
    .Y(_05308_));
 sg13g2_nand2b_1 _13251_ (.Y(_05309_),
    .B(_05308_),
    .A_N(_05298_));
 sg13g2_nand3_1 _13252_ (.B(_05306_),
    .C(_05146_),
    .A(_05303_),
    .Y(_05310_));
 sg13g2_nand2_1 _13253_ (.Y(_05311_),
    .A(_05310_),
    .B(_05298_));
 sg13g2_nand2_1 _13254_ (.Y(_05312_),
    .A(_05309_),
    .B(_05311_));
 sg13g2_nor2_1 _13255_ (.A(_05295_),
    .B(_05312_),
    .Y(_05313_));
 sg13g2_inv_1 _13256_ (.Y(_05314_),
    .A(_05313_));
 sg13g2_nor2_1 _13257_ (.A(_05284_),
    .B(_05294_),
    .Y(_05315_));
 sg13g2_nand2_1 _13258_ (.Y(_05316_),
    .A(_05311_),
    .B(_05315_));
 sg13g2_nand2_1 _13259_ (.Y(_05317_),
    .A(_05316_),
    .B(_05309_));
 sg13g2_inv_1 _13260_ (.Y(_05318_),
    .A(_05317_));
 sg13g2_o21ai_1 _13261_ (.B1(_05318_),
    .Y(_05319_),
    .A1(_05280_),
    .A2(_05314_));
 sg13g2_nand2b_1 _13262_ (.Y(_05320_),
    .B(_05319_),
    .A_N(_05222_));
 sg13g2_nand2b_1 _13263_ (.Y(_05321_),
    .B(_05320_),
    .A_N(_05218_));
 sg13g2_nand2_1 _13264_ (.Y(_05322_),
    .A(\synth.voice.scan_outs[3][0] ),
    .B(net399));
 sg13g2_nand2_1 _13265_ (.Y(_05323_),
    .A(net370),
    .B(_03327_));
 sg13g2_nand2_1 _13266_ (.Y(_05324_),
    .A(net359),
    .B(_05090_));
 sg13g2_and3_1 _13267_ (.X(_05325_),
    .A(_05322_),
    .B(_05323_),
    .C(_05324_));
 sg13g2_nand2_1 _13268_ (.Y(_05326_),
    .A(_05187_),
    .B(net321));
 sg13g2_a21oi_1 _13269_ (.A1(_05031_),
    .A2(_05034_),
    .Y(_05327_),
    .B1(net397));
 sg13g2_buf_1 _13270_ (.A(_05327_),
    .X(_05328_));
 sg13g2_nand3b_1 _13271_ (.B(_05326_),
    .C(net207),
    .Y(_05329_),
    .A_N(_05325_));
 sg13g2_buf_1 _13272_ (.A(_05329_),
    .X(_05330_));
 sg13g2_nand2_1 _13273_ (.Y(_05331_),
    .A(_05326_),
    .B(net207));
 sg13g2_nand2_1 _13274_ (.Y(_05332_),
    .A(_05331_),
    .B(_05325_));
 sg13g2_nand2_2 _13275_ (.Y(_05333_),
    .A(_05330_),
    .B(_05332_));
 sg13g2_nand2_1 _13276_ (.Y(_05334_),
    .A(_05161_),
    .B(net321));
 sg13g2_nand2_1 _13277_ (.Y(_05335_),
    .A(\synth.voice.genblk4[2].next_state_scan[13] ),
    .B(net399));
 sg13g2_inv_1 _13278_ (.Y(_05336_),
    .A(_05335_));
 sg13g2_a221oi_1 _13279_ (.B2(\synth.controller.out[11] ),
    .C1(_05336_),
    .B1(net355),
    .A1(\synth.voice.genblk4[4].next_state_scan[1] ),
    .Y(_05337_),
    .A2(net371));
 sg13g2_inv_1 _13280_ (.Y(_05338_),
    .A(_05337_));
 sg13g2_a21oi_1 _13281_ (.A1(_05334_),
    .A2(net207),
    .Y(_05339_),
    .B1(_05338_));
 sg13g2_nand3_1 _13282_ (.B(net207),
    .C(_05338_),
    .A(_05334_),
    .Y(_05340_));
 sg13g2_buf_1 _13283_ (.A(_05340_),
    .X(_05341_));
 sg13g2_nand2b_1 _13284_ (.Y(_05342_),
    .B(_05341_),
    .A_N(_05339_));
 sg13g2_nor2_1 _13285_ (.A(_05333_),
    .B(_05342_),
    .Y(_05343_));
 sg13g2_nand2_1 _13286_ (.Y(_05344_),
    .A(_05152_),
    .B(\synth.voice.scan_outs[3][1] ));
 sg13g2_inv_1 _13287_ (.Y(_05345_),
    .A(_05344_));
 sg13g2_a221oi_1 _13288_ (.B2(_03330_),
    .C1(_05345_),
    .B1(_05201_),
    .A1(_04989_),
    .Y(_05346_),
    .A2(\synth.voice.genblk4[4].next_state_scan[3] ));
 sg13g2_nand2_1 _13289_ (.Y(_05347_),
    .A(_05120_),
    .B(_05032_));
 sg13g2_nand2_1 _13290_ (.Y(_05348_),
    .A(_05347_),
    .B(net321));
 sg13g2_nand2_1 _13291_ (.Y(_05349_),
    .A(_05348_),
    .B(net207));
 sg13g2_nor2_1 _13292_ (.A(_05346_),
    .B(_05349_),
    .Y(_05350_));
 sg13g2_inv_1 _13293_ (.Y(_05351_),
    .A(_05350_));
 sg13g2_nand2_1 _13294_ (.Y(_05352_),
    .A(_05349_),
    .B(_05346_));
 sg13g2_nand2_2 _13295_ (.Y(_05353_),
    .A(_05351_),
    .B(_05352_));
 sg13g2_nand2_1 _13296_ (.Y(_05354_),
    .A(net371),
    .B(_05015_));
 sg13g2_inv_1 _13297_ (.Y(_05355_),
    .A(_05354_));
 sg13g2_a221oi_1 _13298_ (.B2(\synth.controller.out[14] ),
    .C1(_05355_),
    .B1(net355),
    .A1(net357),
    .Y(_05356_),
    .A2(\synth.voice.genblk4[3].next_state_scan[0] ));
 sg13g2_nand2_1 _13299_ (.Y(_05357_),
    .A(_05033_),
    .B(net321));
 sg13g2_nand2_1 _13300_ (.Y(_05358_),
    .A(_05357_),
    .B(net207));
 sg13g2_nor2_1 _13301_ (.A(_05356_),
    .B(_05358_),
    .Y(_05359_));
 sg13g2_nand2_1 _13302_ (.Y(_05360_),
    .A(_05358_),
    .B(_05356_));
 sg13g2_nand2b_1 _13303_ (.Y(_05361_),
    .B(_05360_),
    .A_N(_05359_));
 sg13g2_nor2_1 _13304_ (.A(_05353_),
    .B(_05361_),
    .Y(_05362_));
 sg13g2_nand2_1 _13305_ (.Y(_05363_),
    .A(_05343_),
    .B(_05362_));
 sg13g2_nand2_1 _13306_ (.Y(_05364_),
    .A(\synth.voice.genblk4[2].next_state_scan[10] ),
    .B(net357));
 sg13g2_nand2_1 _13307_ (.Y(_05365_),
    .A(net355),
    .B(_03364_));
 sg13g2_nand2_1 _13308_ (.Y(_05366_),
    .A(_05047_),
    .B(net371));
 sg13g2_nand3_1 _13309_ (.B(_05365_),
    .C(_05366_),
    .A(_05364_),
    .Y(_05367_));
 sg13g2_nand3_1 _13310_ (.B(_05271_),
    .C(net321),
    .A(_05270_),
    .Y(_05368_));
 sg13g2_nand2_1 _13311_ (.Y(_05369_),
    .A(_05368_),
    .B(_05328_));
 sg13g2_xnor2_1 _13312_ (.Y(_05370_),
    .A(_05367_),
    .B(_05369_));
 sg13g2_inv_1 _13313_ (.Y(_05371_),
    .A(_05370_));
 sg13g2_nand2_1 _13314_ (.Y(_05372_),
    .A(\synth.voice.genblk4[3].next_state_scan[13] ),
    .B(net359));
 sg13g2_inv_1 _13315_ (.Y(_05373_),
    .A(_05372_));
 sg13g2_a221oi_1 _13316_ (.B2(\synth.controller.out[7] ),
    .C1(_05373_),
    .B1(net355),
    .A1(\synth.voice.genblk4[2].next_state_scan[9] ),
    .Y(_05374_),
    .A2(net357));
 sg13g2_nand3_1 _13317_ (.B(net360),
    .C(_05251_),
    .A(_05250_),
    .Y(_05375_));
 sg13g2_nand2_1 _13318_ (.Y(_05376_),
    .A(_05375_),
    .B(_05327_));
 sg13g2_nor2_1 _13319_ (.A(_05374_),
    .B(_05376_),
    .Y(_05377_));
 sg13g2_nand2_1 _13320_ (.Y(_05378_),
    .A(_05376_),
    .B(_05374_));
 sg13g2_nand2b_1 _13321_ (.Y(_05379_),
    .B(_05378_),
    .A_N(_05377_));
 sg13g2_nor2_1 _13322_ (.A(_05371_),
    .B(_05379_),
    .Y(_05380_));
 sg13g2_nand2_1 _13323_ (.Y(_05381_),
    .A(\synth.voice.genblk4[4].next_state_scan[0] ),
    .B(net359));
 sg13g2_nand2_1 _13324_ (.Y(_05382_),
    .A(net370),
    .B(_03316_));
 sg13g2_nand2_1 _13325_ (.Y(_05383_),
    .A(\synth.voice.genblk4[2].next_state_scan[12] ),
    .B(net399));
 sg13g2_and3_1 _13326_ (.X(_05384_),
    .A(_05381_),
    .B(_05382_),
    .C(_05383_));
 sg13g2_nand3_1 _13327_ (.B(_05305_),
    .C(net321),
    .A(_05304_),
    .Y(_05385_));
 sg13g2_nand3b_1 _13328_ (.B(_05385_),
    .C(net207),
    .Y(_05386_),
    .A_N(_05384_));
 sg13g2_buf_1 _13329_ (.A(_05386_),
    .X(_05387_));
 sg13g2_nand2_1 _13330_ (.Y(_05388_),
    .A(_05385_),
    .B(net207));
 sg13g2_nand2_1 _13331_ (.Y(_05389_),
    .A(_05388_),
    .B(_05384_));
 sg13g2_nand2_1 _13332_ (.Y(_05390_),
    .A(_05387_),
    .B(_05389_));
 sg13g2_nand3_1 _13333_ (.B(_05292_),
    .C(net321),
    .A(_05291_),
    .Y(_05391_));
 sg13g2_nand2_1 _13334_ (.Y(_05392_),
    .A(_05391_),
    .B(_05328_));
 sg13g2_inv_1 _13335_ (.Y(_05393_),
    .A(_05392_));
 sg13g2_nand2_1 _13336_ (.Y(_05394_),
    .A(\synth.voice.genblk4[2].next_state_scan[11] ),
    .B(net357));
 sg13g2_nand2_1 _13337_ (.Y(_05395_),
    .A(net355),
    .B(_03366_));
 sg13g2_nand2_1 _13338_ (.Y(_05396_),
    .A(_05040_),
    .B(net371));
 sg13g2_and3_1 _13339_ (.X(_05397_),
    .A(_05394_),
    .B(_05395_),
    .C(_05396_));
 sg13g2_inv_1 _13340_ (.Y(_05398_),
    .A(_05397_));
 sg13g2_nand2_1 _13341_ (.Y(_05399_),
    .A(_05393_),
    .B(_05398_));
 sg13g2_nand2_1 _13342_ (.Y(_05400_),
    .A(_05392_),
    .B(_05397_));
 sg13g2_nand2_1 _13343_ (.Y(_05401_),
    .A(_05399_),
    .B(_05400_));
 sg13g2_nor2_1 _13344_ (.A(_05390_),
    .B(_05401_),
    .Y(_05402_));
 sg13g2_nand2_1 _13345_ (.Y(_05403_),
    .A(_05380_),
    .B(_05402_));
 sg13g2_nor2_1 _13346_ (.A(_05363_),
    .B(_05403_),
    .Y(_05404_));
 sg13g2_nand2_1 _13347_ (.Y(_05405_),
    .A(_05321_),
    .B(_05404_));
 sg13g2_inv_1 _13348_ (.Y(_05406_),
    .A(_05402_));
 sg13g2_nor2b_1 _13349_ (.A(_05369_),
    .B_N(_05367_),
    .Y(_05407_));
 sg13g2_a21oi_1 _13350_ (.A1(_05370_),
    .A2(_05377_),
    .Y(_05408_),
    .B1(_05407_));
 sg13g2_inv_1 _13351_ (.Y(_05409_),
    .A(_05389_));
 sg13g2_a21oi_1 _13352_ (.A1(_05399_),
    .A2(_05387_),
    .Y(_05410_),
    .B1(_05409_));
 sg13g2_inv_1 _13353_ (.Y(_05411_),
    .A(_05410_));
 sg13g2_o21ai_1 _13354_ (.B1(_05411_),
    .Y(_05412_),
    .A1(_05406_),
    .A2(_05408_));
 sg13g2_inv_1 _13355_ (.Y(_05413_),
    .A(_05363_));
 sg13g2_o21ai_1 _13356_ (.B1(_05330_),
    .Y(_05414_),
    .A1(_05341_),
    .A2(_05333_));
 sg13g2_inv_1 _13357_ (.Y(_05415_),
    .A(_05414_));
 sg13g2_nor2_1 _13358_ (.A(_05359_),
    .B(_05350_),
    .Y(_05416_));
 sg13g2_o21ai_1 _13359_ (.B1(_05416_),
    .Y(_05417_),
    .A1(_05353_),
    .A2(_05415_));
 sg13g2_a22oi_1 _13360_ (.Y(_05418_),
    .B1(_05360_),
    .B2(_05417_),
    .A2(_05413_),
    .A1(_05412_));
 sg13g2_nand2_1 _13361_ (.Y(_05419_),
    .A(_05248_),
    .B(_05252_));
 sg13g2_nand2b_1 _13362_ (.Y(_05420_),
    .B(_05419_),
    .A_N(_05256_));
 sg13g2_nand2_1 _13363_ (.Y(_05421_),
    .A(_05420_),
    .B(_05258_));
 sg13g2_xnor2_1 _13364_ (.Y(_05422_),
    .A(_05277_),
    .B(_05273_));
 sg13g2_nor2_1 _13365_ (.A(_05421_),
    .B(_05422_),
    .Y(_05423_));
 sg13g2_nand2_1 _13366_ (.Y(_05424_),
    .A(_05313_),
    .B(_05423_));
 sg13g2_nor2_1 _13367_ (.A(_05424_),
    .B(_05222_),
    .Y(_05425_));
 sg13g2_inv_1 _13368_ (.Y(_05426_),
    .A(\synth.voice.scan_outs[2][0] ));
 sg13g2_nand2_1 _13369_ (.Y(_05427_),
    .A(\synth.voice.genblk4[3].next_state_scan[2] ),
    .B(net358));
 sg13g2_o21ai_1 _13370_ (.B1(_05427_),
    .Y(_05428_),
    .A1(_05426_),
    .A2(net322));
 sg13g2_xnor2_1 _13371_ (.Y(_05429_),
    .A(net363),
    .B(_05428_));
 sg13g2_nand2_1 _13372_ (.Y(_05430_),
    .A(_05429_),
    .B(net325));
 sg13g2_inv_1 _13373_ (.Y(_05431_),
    .A(\synth.voice.scan_outs[2][1] ));
 sg13g2_nand2_1 _13374_ (.Y(_05432_),
    .A(net358),
    .B(\synth.voice.genblk4[3].next_state_scan[3] ));
 sg13g2_o21ai_1 _13375_ (.B1(_05432_),
    .Y(_05433_),
    .A1(net322),
    .A2(_05431_));
 sg13g2_xnor2_1 _13376_ (.Y(_05434_),
    .A(net363),
    .B(_05433_));
 sg13g2_a21oi_1 _13377_ (.A1(_05434_),
    .A2(net364),
    .Y(_05435_),
    .B1(net356));
 sg13g2_inv_1 _13378_ (.Y(_05436_),
    .A(\synth.voice.genblk4[2].next_state_scan[0] ));
 sg13g2_nand2_1 _13379_ (.Y(_05437_),
    .A(_05137_),
    .B(\synth.voice.genblk4[3].next_state_scan[4] ));
 sg13g2_o21ai_1 _13380_ (.B1(_05437_),
    .Y(_05438_),
    .A1(_05135_),
    .A2(_05436_));
 sg13g2_xnor2_1 _13381_ (.Y(_05439_),
    .A(_05013_),
    .B(_05438_));
 sg13g2_mux2_1 _13382_ (.A0(_05439_),
    .A1(_05230_),
    .S(net364),
    .X(_05440_));
 sg13g2_a22oi_1 _13383_ (.Y(_05441_),
    .B1(net356),
    .B2(_05440_),
    .A2(_05435_),
    .A1(_05430_));
 sg13g2_a21oi_1 _13384_ (.A1(_05441_),
    .A2(_05073_),
    .Y(_05442_),
    .B1(net365));
 sg13g2_nand2b_1 _13385_ (.Y(_05443_),
    .B(net361),
    .A_N(_05266_));
 sg13g2_inv_1 _13386_ (.Y(_05444_),
    .A(_00144_));
 sg13g2_a21oi_1 _13387_ (.A1(_05442_),
    .A2(_05443_),
    .Y(_05445_),
    .B1(_05444_));
 sg13g2_nand3_1 _13388_ (.B(_05197_),
    .C(net365),
    .A(_05191_),
    .Y(_05446_));
 sg13g2_nand2_1 _13389_ (.Y(_05447_),
    .A(_05445_),
    .B(_05446_));
 sg13g2_nand2_1 _13390_ (.Y(_05448_),
    .A(\synth.voice.scan_outs[2][0] ),
    .B(net357));
 sg13g2_nand2_1 _13391_ (.Y(_05449_),
    .A(\synth.voice.acc[0] ),
    .B(net355));
 sg13g2_nand2_1 _13392_ (.Y(_05450_),
    .A(\synth.voice.genblk4[3].next_state_scan[2] ),
    .B(net371));
 sg13g2_and3_1 _13393_ (.X(_05451_),
    .A(_05448_),
    .B(_05449_),
    .C(_05450_));
 sg13g2_nand2_1 _13394_ (.Y(_05452_),
    .A(_05447_),
    .B(_05451_));
 sg13g2_nor2_1 _13395_ (.A(_05020_),
    .B(_05439_),
    .Y(_05453_));
 sg13g2_a21oi_1 _13396_ (.A1(net325),
    .A2(_05434_),
    .Y(_05454_),
    .B1(_05453_));
 sg13g2_nand2b_1 _13397_ (.Y(_05455_),
    .B(net364),
    .A_N(_05429_));
 sg13g2_a21oi_1 _13398_ (.A1(net325),
    .A2(net363),
    .Y(_05456_),
    .B1(net356));
 sg13g2_a21oi_1 _13399_ (.A1(_05455_),
    .A2(_05456_),
    .Y(_05457_),
    .B1(net361));
 sg13g2_o21ai_1 _13400_ (.B1(_05457_),
    .Y(_05458_),
    .A1(net324),
    .A2(_05454_));
 sg13g2_o21ai_1 _13401_ (.B1(_05458_),
    .Y(_05459_),
    .A1(net323),
    .A2(_05245_));
 sg13g2_nand3_1 _13402_ (.B(_05179_),
    .C(net365),
    .A(_05166_),
    .Y(_05460_));
 sg13g2_nand2_1 _13403_ (.Y(_05461_),
    .A(_05460_),
    .B(_00144_));
 sg13g2_a21oi_2 _13404_ (.B1(_05461_),
    .Y(_05462_),
    .A2(_05459_),
    .A1(net321));
 sg13g2_nand3b_1 _13405_ (.B(_05445_),
    .C(_05446_),
    .Y(_05463_),
    .A_N(_05451_));
 sg13g2_buf_1 _13406_ (.A(_05463_),
    .X(_05464_));
 sg13g2_inv_1 _13407_ (.Y(_05465_),
    .A(_05464_));
 sg13g2_a21oi_2 _13408_ (.B1(_05465_),
    .Y(_05466_),
    .A2(_05462_),
    .A1(_05452_));
 sg13g2_nand2_1 _13409_ (.Y(_05467_),
    .A(\synth.voice.genblk4[3].next_state_scan[4] ),
    .B(net371));
 sg13g2_nand2_1 _13410_ (.Y(_05468_),
    .A(_04991_),
    .B(\synth.voice.acc[2] ));
 sg13g2_nand2_1 _13411_ (.Y(_05469_),
    .A(\synth.voice.genblk4[2].next_state_scan[0] ),
    .B(net399));
 sg13g2_nand3_1 _13412_ (.B(_05468_),
    .C(_05469_),
    .A(_05467_),
    .Y(_05470_));
 sg13g2_nand3_1 _13413_ (.B(_05104_),
    .C(_05035_),
    .A(_05074_),
    .Y(_05471_));
 sg13g2_nor2_1 _13414_ (.A(net356),
    .B(_05440_),
    .Y(_05472_));
 sg13g2_a21oi_1 _13415_ (.A1(_05164_),
    .A2(_05262_),
    .Y(_05473_),
    .B1(_05472_));
 sg13g2_nor2_1 _13416_ (.A(_05103_),
    .B(_05473_),
    .Y(_05474_));
 sg13g2_nand3_1 _13417_ (.B(_05301_),
    .C(_05028_),
    .A(_05300_),
    .Y(_05475_));
 sg13g2_nand2_1 _13418_ (.Y(_05476_),
    .A(_05475_),
    .B(net360));
 sg13g2_nor2_1 _13419_ (.A(_05474_),
    .B(_05476_),
    .Y(_05477_));
 sg13g2_nor2_1 _13420_ (.A(net397),
    .B(_05477_),
    .Y(_05478_));
 sg13g2_nand2_1 _13421_ (.Y(_05479_),
    .A(_05471_),
    .B(_05478_));
 sg13g2_nand2b_1 _13422_ (.Y(_05480_),
    .B(_05479_),
    .A_N(_05470_));
 sg13g2_nand3_1 _13423_ (.B(_05478_),
    .C(_05470_),
    .A(_05471_),
    .Y(_05481_));
 sg13g2_buf_1 _13424_ (.A(_05481_),
    .X(_05482_));
 sg13g2_nand2_1 _13425_ (.Y(_05483_),
    .A(_05480_),
    .B(_05482_));
 sg13g2_nand2_1 _13426_ (.Y(_05484_),
    .A(\synth.voice.genblk4[3].next_state_scan[3] ),
    .B(_05109_));
 sg13g2_nand2_1 _13427_ (.Y(_05485_),
    .A(_04991_),
    .B(\synth.voice.acc[1] ));
 sg13g2_nand2_1 _13428_ (.Y(_05486_),
    .A(\synth.voice.scan_outs[2][1] ),
    .B(net399));
 sg13g2_nand3_1 _13429_ (.B(_05485_),
    .C(_05486_),
    .A(_05484_),
    .Y(_05487_));
 sg13g2_nand2_1 _13430_ (.Y(_05488_),
    .A(_05454_),
    .B(net324));
 sg13g2_nand2_1 _13431_ (.Y(_05489_),
    .A(_05232_),
    .B(net362));
 sg13g2_nand3_1 _13432_ (.B(_05489_),
    .C(_05029_),
    .A(_05488_),
    .Y(_05490_));
 sg13g2_nand2_1 _13433_ (.Y(_05491_),
    .A(_05490_),
    .B(net360));
 sg13g2_a21oi_1 _13434_ (.A1(_05103_),
    .A2(_05287_),
    .Y(_05492_),
    .B1(_05491_));
 sg13g2_nor2_1 _13435_ (.A(net397),
    .B(_05492_),
    .Y(_05493_));
 sg13g2_nand3_1 _13436_ (.B(_05035_),
    .C(_05144_),
    .A(_05128_),
    .Y(_05494_));
 sg13g2_nand2_1 _13437_ (.Y(_05495_),
    .A(_05493_),
    .B(_05494_));
 sg13g2_nand2b_1 _13438_ (.Y(_05496_),
    .B(_05495_),
    .A_N(_05487_));
 sg13g2_nand3_1 _13439_ (.B(_05494_),
    .C(_05487_),
    .A(_05493_),
    .Y(_05497_));
 sg13g2_buf_1 _13440_ (.A(_05497_),
    .X(_05498_));
 sg13g2_nand2_1 _13441_ (.Y(_05499_),
    .A(_05496_),
    .B(_05498_));
 sg13g2_nor2_1 _13442_ (.A(_05483_),
    .B(_05499_),
    .Y(_05500_));
 sg13g2_inv_1 _13443_ (.Y(_05501_),
    .A(_05500_));
 sg13g2_inv_1 _13444_ (.Y(_05502_),
    .A(_05480_));
 sg13g2_o21ai_1 _13445_ (.B1(_05482_),
    .Y(_05503_),
    .A1(_05498_),
    .A2(_05502_));
 sg13g2_inv_1 _13446_ (.Y(_05504_),
    .A(_05503_));
 sg13g2_o21ai_1 _13447_ (.B1(_05504_),
    .Y(_05505_),
    .A1(_05466_),
    .A2(_05501_));
 sg13g2_buf_1 _13448_ (.A(_05505_),
    .X(_05506_));
 sg13g2_nand3_1 _13449_ (.B(_05506_),
    .C(_05404_),
    .A(_05425_),
    .Y(_05507_));
 sg13g2_nand2_1 _13450_ (.Y(_05508_),
    .A(net371),
    .B(_05005_));
 sg13g2_inv_1 _13451_ (.Y(_05509_),
    .A(_05508_));
 sg13g2_a221oi_1 _13452_ (.B2(\synth.controller.out[15] ),
    .C1(_05509_),
    .B1(net355),
    .A1(net357),
    .Y(_05510_),
    .A2(\synth.voice.genblk4[3].next_state_scan[1] ));
 sg13g2_nand2_1 _13453_ (.Y(_05511_),
    .A(_05009_),
    .B(_00144_));
 sg13g2_nor2_1 _13454_ (.A(_05510_),
    .B(_05511_),
    .Y(_05512_));
 sg13g2_nand4_1 _13455_ (.B(_05418_),
    .C(_05507_),
    .A(_05405_),
    .Y(_05513_),
    .D(_05512_));
 sg13g2_buf_1 _13456_ (.A(_05513_),
    .X(_05514_));
 sg13g2_buf_1 _13457_ (.A(net71),
    .X(_05515_));
 sg13g2_nand2_1 _13458_ (.Y(_05516_),
    .A(_05464_),
    .B(_05452_));
 sg13g2_xnor2_1 _13459_ (.Y(_05517_),
    .A(_05462_),
    .B(_05516_));
 sg13g2_nand2_1 _13460_ (.Y(_05518_),
    .A(net66),
    .B(_05517_));
 sg13g2_nand2_1 _13461_ (.Y(_05519_),
    .A(_05511_),
    .B(_05510_));
 sg13g2_nand3_1 _13462_ (.B(_05418_),
    .C(_05507_),
    .A(_05405_),
    .Y(_05520_));
 sg13g2_nand2b_1 _13463_ (.Y(_05521_),
    .B(_05520_),
    .A_N(_05519_));
 sg13g2_buf_1 _13464_ (.A(_05521_),
    .X(_05522_));
 sg13g2_buf_1 _13465_ (.A(net65),
    .X(_05523_));
 sg13g2_nand2_1 _13466_ (.Y(_05524_),
    .A(_05518_),
    .B(net45));
 sg13g2_nor2_1 _13467_ (.A(_04785_),
    .B(_04029_),
    .Y(_05525_));
 sg13g2_a21o_1 _13468_ (.A2(_04021_),
    .A1(_03607_),
    .B1(_05525_),
    .X(_05526_));
 sg13g2_buf_1 _13469_ (.A(_05526_),
    .X(_05527_));
 sg13g2_nor2b_2 _13470_ (.A(net242),
    .B_N(\synth.voice.target_reg[1] ),
    .Y(_05528_));
 sg13g2_nor2b_1 _13471_ (.A(net169),
    .B_N(_05528_),
    .Y(_05529_));
 sg13g2_buf_2 _13472_ (.A(_05529_),
    .X(_05530_));
 sg13g2_buf_1 _13473_ (.A(_05530_),
    .X(_05531_));
 sg13g2_nand2_1 _13474_ (.Y(_05532_),
    .A(_05524_),
    .B(net126));
 sg13g2_buf_1 _13475_ (.A(_05527_),
    .X(_05533_));
 sg13g2_nor2_1 _13476_ (.A(_05528_),
    .B(net169),
    .Y(_05534_));
 sg13g2_buf_2 _13477_ (.A(_05534_),
    .X(_05535_));
 sg13g2_buf_1 _13478_ (.A(_05535_),
    .X(_05536_));
 sg13g2_a22oi_1 _13479_ (.Y(_05537_),
    .B1(\synth.voice.scan_outs[2][0] ),
    .B2(net125),
    .A2(net152),
    .A1(\synth.voice.genblk4[2].next_state_scan[0] ));
 sg13g2_nand2_1 _13480_ (.Y(_01215_),
    .A(_05532_),
    .B(_05537_));
 sg13g2_xor2_1 _13481_ (.B(_05466_),
    .A(_05499_),
    .X(_05538_));
 sg13g2_nand2_1 _13482_ (.Y(_05539_),
    .A(net66),
    .B(_05538_));
 sg13g2_nand2_1 _13483_ (.Y(_05540_),
    .A(_05539_),
    .B(net45));
 sg13g2_nand2_1 _13484_ (.Y(_05541_),
    .A(_05540_),
    .B(_05531_));
 sg13g2_a22oi_1 _13485_ (.Y(_05542_),
    .B1(\synth.voice.scan_outs[2][1] ),
    .B2(net125),
    .A2(net152),
    .A1(\synth.voice.genblk4[2].next_state_scan[1] ));
 sg13g2_nand2_1 _13486_ (.Y(_01216_),
    .A(_05541_),
    .B(_05542_));
 sg13g2_a21oi_1 _13487_ (.A1(_05493_),
    .A2(_05494_),
    .Y(_05543_),
    .B1(_05487_));
 sg13g2_o21ai_1 _13488_ (.B1(_05498_),
    .Y(_05544_),
    .A1(_05464_),
    .A2(_05543_));
 sg13g2_nor2_1 _13489_ (.A(_05499_),
    .B(_05516_),
    .Y(_05545_));
 sg13g2_nand2_1 _13490_ (.Y(_05546_),
    .A(_05545_),
    .B(_05462_));
 sg13g2_nand2b_1 _13491_ (.Y(_05547_),
    .B(_05546_),
    .A_N(_05544_));
 sg13g2_buf_1 _13492_ (.A(_05547_),
    .X(_05548_));
 sg13g2_xnor2_1 _13493_ (.Y(_05549_),
    .A(_05483_),
    .B(_05548_));
 sg13g2_nand2_1 _13494_ (.Y(_05550_),
    .A(net66),
    .B(_05549_));
 sg13g2_nand2_1 _13495_ (.Y(_05551_),
    .A(_05550_),
    .B(net45));
 sg13g2_nand2_1 _13496_ (.Y(_05552_),
    .A(_05551_),
    .B(net126));
 sg13g2_a22oi_1 _13497_ (.Y(_05553_),
    .B1(\synth.voice.genblk4[2].next_state_scan[0] ),
    .B2(net125),
    .A2(net152),
    .A1(\synth.voice.genblk4[2].next_state_scan[2] ));
 sg13g2_nand2_1 _13498_ (.Y(_01217_),
    .A(_05552_),
    .B(_05553_));
 sg13g2_xnor2_1 _13499_ (.Y(_05554_),
    .A(_05421_),
    .B(_05506_));
 sg13g2_nand2_1 _13500_ (.Y(_05555_),
    .A(net66),
    .B(_05554_));
 sg13g2_nand2_1 _13501_ (.Y(_05556_),
    .A(_05555_),
    .B(net45));
 sg13g2_nand2_1 _13502_ (.Y(_05557_),
    .A(_05556_),
    .B(net126));
 sg13g2_a22oi_1 _13503_ (.Y(_05558_),
    .B1(\synth.voice.genblk4[2].next_state_scan[1] ),
    .B2(net125),
    .A2(net152),
    .A1(\synth.voice.genblk4[2].next_state_scan[3] ));
 sg13g2_nand2_1 _13504_ (.Y(_01218_),
    .A(_05557_),
    .B(_05558_));
 sg13g2_nor2_1 _13505_ (.A(_05483_),
    .B(_05421_),
    .Y(_05559_));
 sg13g2_nand2_1 _13506_ (.Y(_05560_),
    .A(_05548_),
    .B(_05559_));
 sg13g2_inv_1 _13507_ (.Y(_05561_),
    .A(_05420_));
 sg13g2_a21oi_1 _13508_ (.A1(_05258_),
    .A2(_05482_),
    .Y(_05562_),
    .B1(_05561_));
 sg13g2_inv_1 _13509_ (.Y(_05563_),
    .A(_05562_));
 sg13g2_nand2_1 _13510_ (.Y(_05564_),
    .A(_05560_),
    .B(_05563_));
 sg13g2_xnor2_1 _13511_ (.Y(_05565_),
    .A(_05422_),
    .B(_05564_));
 sg13g2_nand2_1 _13512_ (.Y(_05566_),
    .A(net66),
    .B(_05565_));
 sg13g2_nand2_1 _13513_ (.Y(_05567_),
    .A(_05566_),
    .B(net45));
 sg13g2_nand2_1 _13514_ (.Y(_05568_),
    .A(_05567_),
    .B(net126));
 sg13g2_a22oi_1 _13515_ (.Y(_05569_),
    .B1(\synth.voice.genblk4[2].next_state_scan[2] ),
    .B2(_05536_),
    .A2(_05533_),
    .A1(\synth.voice.genblk4[2].next_state_scan[4] ));
 sg13g2_nand2_1 _13516_ (.Y(_01219_),
    .A(_05568_),
    .B(_05569_));
 sg13g2_nand2_1 _13517_ (.Y(_05570_),
    .A(_05506_),
    .B(_05423_));
 sg13g2_nand2_1 _13518_ (.Y(_05571_),
    .A(_05570_),
    .B(_05280_));
 sg13g2_xnor2_1 _13519_ (.Y(_05572_),
    .A(_05295_),
    .B(_05571_));
 sg13g2_nand2_1 _13520_ (.Y(_05573_),
    .A(net66),
    .B(_05572_));
 sg13g2_nand2_1 _13521_ (.Y(_05574_),
    .A(_05573_),
    .B(_05523_));
 sg13g2_nand2_1 _13522_ (.Y(_05575_),
    .A(_05574_),
    .B(net126));
 sg13g2_a22oi_1 _13523_ (.Y(_05576_),
    .B1(\synth.voice.genblk4[2].next_state_scan[3] ),
    .B2(_05536_),
    .A2(_05533_),
    .A1(\synth.voice.genblk4[2].next_state_scan[5] ));
 sg13g2_nand2_1 _13524_ (.Y(_01220_),
    .A(_05575_),
    .B(_05576_));
 sg13g2_nor2_1 _13525_ (.A(_05295_),
    .B(_05422_),
    .Y(_05577_));
 sg13g2_nand2_1 _13526_ (.Y(_05578_),
    .A(_05577_),
    .B(_05562_));
 sg13g2_nand2_1 _13527_ (.Y(_05579_),
    .A(_05294_),
    .B(_05284_));
 sg13g2_a21oi_1 _13528_ (.A1(_05279_),
    .A2(_05579_),
    .Y(_05580_),
    .B1(_05315_));
 sg13g2_nand2_1 _13529_ (.Y(_05581_),
    .A(_05578_),
    .B(_05580_));
 sg13g2_nand2_1 _13530_ (.Y(_05582_),
    .A(_05577_),
    .B(_05559_));
 sg13g2_nand2b_1 _13531_ (.Y(_05583_),
    .B(_05548_),
    .A_N(_05582_));
 sg13g2_nand2b_1 _13532_ (.Y(_05584_),
    .B(_05583_),
    .A_N(_05581_));
 sg13g2_xnor2_1 _13533_ (.Y(_05585_),
    .A(_05312_),
    .B(_05584_));
 sg13g2_nand2_1 _13534_ (.Y(_05586_),
    .A(net66),
    .B(_05585_));
 sg13g2_nand2_1 _13535_ (.Y(_05587_),
    .A(_05586_),
    .B(net45));
 sg13g2_nand2_1 _13536_ (.Y(_05588_),
    .A(_05587_),
    .B(_05531_));
 sg13g2_a22oi_1 _13537_ (.Y(_05589_),
    .B1(\synth.voice.genblk4[2].next_state_scan[4] ),
    .B2(net125),
    .A2(net152),
    .A1(\synth.voice.genblk4[2].next_state_scan[6] ));
 sg13g2_nand2_1 _13538_ (.Y(_01221_),
    .A(_05588_),
    .B(_05589_));
 sg13g2_nand2b_1 _13539_ (.Y(_05590_),
    .B(_05506_),
    .A_N(_05424_));
 sg13g2_inv_1 _13540_ (.Y(_05591_),
    .A(_05319_));
 sg13g2_nand2_1 _13541_ (.Y(_05592_),
    .A(_05590_),
    .B(_05591_));
 sg13g2_xnor2_1 _13542_ (.Y(_05593_),
    .A(_05220_),
    .B(_05592_));
 sg13g2_nand2_1 _13543_ (.Y(_05594_),
    .A(_05515_),
    .B(_05593_));
 sg13g2_nand2_1 _13544_ (.Y(_05595_),
    .A(_05594_),
    .B(net45));
 sg13g2_nand2_1 _13545_ (.Y(_05596_),
    .A(_05595_),
    .B(net126));
 sg13g2_a22oi_1 _13546_ (.Y(_05597_),
    .B1(\synth.voice.genblk4[2].next_state_scan[5] ),
    .B2(net125),
    .A2(net152),
    .A1(\synth.voice.genblk4[2].next_state_scan[7] ));
 sg13g2_nand2_1 _13547_ (.Y(_01222_),
    .A(_05596_),
    .B(_05597_));
 sg13g2_nor3_1 _13548_ (.A(_03668_),
    .B(_01737_),
    .C(net242),
    .Y(_05598_));
 sg13g2_xnor2_1 _13549_ (.Y(_05599_),
    .A(_04908_),
    .B(_05598_));
 sg13g2_nor2_1 _13550_ (.A(\synth.voice.coeff_index[2] ),
    .B(_04711_),
    .Y(_05600_));
 sg13g2_a21oi_1 _13551_ (.A1(_05599_),
    .A2(_04711_),
    .Y(_01223_),
    .B1(_05600_));
 sg13g2_inv_1 _13552_ (.Y(_05601_),
    .A(_05219_));
 sg13g2_nand2_1 _13553_ (.Y(_05602_),
    .A(_05545_),
    .B(_05559_));
 sg13g2_nor2_1 _13554_ (.A(_05312_),
    .B(_05220_),
    .Y(_05603_));
 sg13g2_nand2_1 _13555_ (.Y(_05604_),
    .A(_05603_),
    .B(_05577_));
 sg13g2_nor2_1 _13556_ (.A(_05602_),
    .B(_05604_),
    .Y(_05605_));
 sg13g2_nand2_1 _13557_ (.Y(_05606_),
    .A(_05544_),
    .B(_05559_));
 sg13g2_nand2_1 _13558_ (.Y(_05607_),
    .A(_05606_),
    .B(_05563_));
 sg13g2_nand2b_1 _13559_ (.Y(_05608_),
    .B(_05607_),
    .A_N(_05604_));
 sg13g2_inv_1 _13560_ (.Y(_05609_),
    .A(_05580_));
 sg13g2_inv_1 _13561_ (.Y(_05610_),
    .A(_05309_));
 sg13g2_nand2_1 _13562_ (.Y(_05611_),
    .A(_05181_),
    .B(_05156_));
 sg13g2_nand2_1 _13563_ (.Y(_05612_),
    .A(_05610_),
    .B(_05611_));
 sg13g2_nand2b_1 _13564_ (.Y(_05613_),
    .B(_05612_),
    .A_N(_05182_));
 sg13g2_a21oi_1 _13565_ (.A1(_05603_),
    .A2(_05609_),
    .Y(_05614_),
    .B1(_05613_));
 sg13g2_nand2_1 _13566_ (.Y(_05615_),
    .A(_05608_),
    .B(_05614_));
 sg13g2_a21oi_1 _13567_ (.A1(_05462_),
    .A2(_05605_),
    .Y(_05616_),
    .B1(_05615_));
 sg13g2_xnor2_1 _13568_ (.Y(_05617_),
    .A(_05601_),
    .B(_05616_));
 sg13g2_nand2_1 _13569_ (.Y(_05618_),
    .A(net66),
    .B(_05617_));
 sg13g2_nand2_1 _13570_ (.Y(_05619_),
    .A(_05618_),
    .B(net45));
 sg13g2_nand2_1 _13571_ (.Y(_05620_),
    .A(_05619_),
    .B(net126));
 sg13g2_a22oi_1 _13572_ (.Y(_05621_),
    .B1(\synth.voice.genblk4[2].next_state_scan[6] ),
    .B2(net125),
    .A2(net152),
    .A1(\synth.voice.genblk4[2].next_state_scan[8] ));
 sg13g2_nand2_1 _13573_ (.Y(_01224_),
    .A(_05620_),
    .B(_05621_));
 sg13g2_inv_1 _13574_ (.Y(_05622_),
    .A(_05215_));
 sg13g2_inv_1 _13575_ (.Y(_05623_),
    .A(_05466_));
 sg13g2_nand2_1 _13576_ (.Y(_05624_),
    .A(_05423_),
    .B(_05500_));
 sg13g2_nand2_1 _13577_ (.Y(_05625_),
    .A(_05221_),
    .B(_05313_));
 sg13g2_nor2_1 _13578_ (.A(_05624_),
    .B(_05625_),
    .Y(_05626_));
 sg13g2_nand2_1 _13579_ (.Y(_05627_),
    .A(_05423_),
    .B(_05503_));
 sg13g2_nand2_1 _13580_ (.Y(_05628_),
    .A(_05627_),
    .B(_05280_));
 sg13g2_nand2b_1 _13581_ (.Y(_05629_),
    .B(_05628_),
    .A_N(_05625_));
 sg13g2_a21oi_1 _13582_ (.A1(_05221_),
    .A2(_05317_),
    .Y(_05630_),
    .B1(_05209_));
 sg13g2_nand2_1 _13583_ (.Y(_05631_),
    .A(_05629_),
    .B(_05630_));
 sg13g2_a21oi_1 _13584_ (.A1(_05623_),
    .A2(_05626_),
    .Y(_05632_),
    .B1(_05631_));
 sg13g2_xnor2_1 _13585_ (.Y(_05633_),
    .A(_05622_),
    .B(_05632_));
 sg13g2_nand2_1 _13586_ (.Y(_05634_),
    .A(_05515_),
    .B(_05633_));
 sg13g2_nand2_1 _13587_ (.Y(_05635_),
    .A(_05634_),
    .B(_05523_));
 sg13g2_nand2_1 _13588_ (.Y(_05636_),
    .A(_05635_),
    .B(net126));
 sg13g2_a22oi_1 _13589_ (.Y(_05637_),
    .B1(\synth.voice.genblk4[2].next_state_scan[7] ),
    .B2(net125),
    .A2(net152),
    .A1(\synth.voice.genblk4[2].next_state_scan[9] ));
 sg13g2_nand2_1 _13590_ (.Y(_01225_),
    .A(_05636_),
    .B(_05637_));
 sg13g2_nor2_1 _13591_ (.A(_05219_),
    .B(_05215_),
    .Y(_05638_));
 sg13g2_nand2_1 _13592_ (.Y(_05639_),
    .A(_05638_),
    .B(_05603_));
 sg13g2_nor2_1 _13593_ (.A(_05582_),
    .B(_05639_),
    .Y(_05640_));
 sg13g2_inv_1 _13594_ (.Y(_05641_),
    .A(_05639_));
 sg13g2_nand2_1 _13595_ (.Y(_05642_),
    .A(_05581_),
    .B(_05641_));
 sg13g2_nand2_1 _13596_ (.Y(_05643_),
    .A(_05211_),
    .B(_05207_));
 sg13g2_nand2_1 _13597_ (.Y(_05644_),
    .A(_05643_),
    .B(_05214_));
 sg13g2_a21oi_1 _13598_ (.A1(_05613_),
    .A2(_05638_),
    .Y(_05645_),
    .B1(_05644_));
 sg13g2_nand2_1 _13599_ (.Y(_05646_),
    .A(_05642_),
    .B(_05645_));
 sg13g2_a21oi_1 _13600_ (.A1(_05548_),
    .A2(_05640_),
    .Y(_05647_),
    .B1(_05646_));
 sg13g2_xor2_1 _13601_ (.B(_05647_),
    .A(_05210_),
    .X(_05648_));
 sg13g2_nand2_1 _13602_ (.Y(_05649_),
    .A(_05514_),
    .B(_05648_));
 sg13g2_nand2_1 _13603_ (.Y(_05650_),
    .A(_05649_),
    .B(_05522_));
 sg13g2_nand2_1 _13604_ (.Y(_05651_),
    .A(_05650_),
    .B(_05530_));
 sg13g2_a22oi_1 _13605_ (.Y(_05652_),
    .B1(\synth.voice.genblk4[2].next_state_scan[8] ),
    .B2(_05535_),
    .A2(net169),
    .A1(\synth.voice.genblk4[2].next_state_scan[10] ));
 sg13g2_nand2_1 _13606_ (.Y(_01226_),
    .A(_05651_),
    .B(_05652_));
 sg13g2_nand2_1 _13607_ (.Y(_05653_),
    .A(_05425_),
    .B(_05506_));
 sg13g2_nor2b_1 _13608_ (.A(_05321_),
    .B_N(_05653_),
    .Y(_05654_));
 sg13g2_xor2_1 _13609_ (.B(_05654_),
    .A(_05379_),
    .X(_05655_));
 sg13g2_nand2_1 _13610_ (.Y(_05656_),
    .A(net71),
    .B(_05655_));
 sg13g2_nand2_1 _13611_ (.Y(_05657_),
    .A(_05656_),
    .B(net65));
 sg13g2_nand2_1 _13612_ (.Y(_05658_),
    .A(_05657_),
    .B(_05530_));
 sg13g2_a22oi_1 _13613_ (.Y(_05659_),
    .B1(\synth.voice.genblk4[2].next_state_scan[9] ),
    .B2(_05535_),
    .A2(net169),
    .A1(\synth.voice.genblk4[2].next_state_scan[11] ));
 sg13g2_nand2_1 _13614_ (.Y(_01227_),
    .A(_05658_),
    .B(_05659_));
 sg13g2_nor2_1 _13615_ (.A(_05210_),
    .B(_05379_),
    .Y(_05660_));
 sg13g2_nand2_1 _13616_ (.Y(_05661_),
    .A(_05638_),
    .B(_05660_));
 sg13g2_nor2_1 _13617_ (.A(_05604_),
    .B(_05661_),
    .Y(_05662_));
 sg13g2_nand2_1 _13618_ (.Y(_05663_),
    .A(_05564_),
    .B(_05662_));
 sg13g2_nand2_1 _13619_ (.Y(_05664_),
    .A(_05108_),
    .B(_05378_));
 sg13g2_nand2b_1 _13620_ (.Y(_05665_),
    .B(_05664_),
    .A_N(_05377_));
 sg13g2_nand2_1 _13621_ (.Y(_05666_),
    .A(_05644_),
    .B(_05660_));
 sg13g2_nand2b_1 _13622_ (.Y(_05667_),
    .B(_05666_),
    .A_N(_05665_));
 sg13g2_nor2_1 _13623_ (.A(_05661_),
    .B(_05614_),
    .Y(_05668_));
 sg13g2_nor2_1 _13624_ (.A(_05667_),
    .B(_05668_),
    .Y(_05669_));
 sg13g2_nand2_1 _13625_ (.Y(_05670_),
    .A(_05663_),
    .B(_05669_));
 sg13g2_xnor2_1 _13626_ (.Y(_05671_),
    .A(_05371_),
    .B(_05670_));
 sg13g2_nand2_1 _13627_ (.Y(_05672_),
    .A(net71),
    .B(_05671_));
 sg13g2_nand2_1 _13628_ (.Y(_05673_),
    .A(_05672_),
    .B(net65));
 sg13g2_nand2_1 _13629_ (.Y(_05674_),
    .A(_05673_),
    .B(_05530_));
 sg13g2_a22oi_1 _13630_ (.Y(_05675_),
    .B1(\synth.voice.genblk4[2].next_state_scan[10] ),
    .B2(_05535_),
    .A2(net169),
    .A1(\synth.voice.genblk4[2].next_state_scan[12] ));
 sg13g2_nand2_1 _13631_ (.Y(_01228_),
    .A(_05674_),
    .B(_05675_));
 sg13g2_nand2_1 _13632_ (.Y(_05676_),
    .A(_05216_),
    .B(_05380_));
 sg13g2_nor2_1 _13633_ (.A(_05625_),
    .B(_05676_),
    .Y(_05677_));
 sg13g2_nand2_1 _13634_ (.Y(_05678_),
    .A(_05571_),
    .B(_05677_));
 sg13g2_nand2_1 _13635_ (.Y(_05679_),
    .A(_05151_),
    .B(_05380_));
 sg13g2_nand2_1 _13636_ (.Y(_05680_),
    .A(_05679_),
    .B(_05408_));
 sg13g2_nor2_1 _13637_ (.A(_05676_),
    .B(_05630_),
    .Y(_05681_));
 sg13g2_nor2_1 _13638_ (.A(_05680_),
    .B(_05681_),
    .Y(_05682_));
 sg13g2_nand2_1 _13639_ (.Y(_05683_),
    .A(_05678_),
    .B(_05682_));
 sg13g2_xnor2_1 _13640_ (.Y(_05684_),
    .A(_05401_),
    .B(_05683_));
 sg13g2_nand2_1 _13641_ (.Y(_05685_),
    .A(net71),
    .B(_05684_));
 sg13g2_nand2_1 _13642_ (.Y(_05686_),
    .A(_05685_),
    .B(net65));
 sg13g2_nand2_1 _13643_ (.Y(_05687_),
    .A(_05686_),
    .B(_05530_));
 sg13g2_a22oi_1 _13644_ (.Y(_05688_),
    .B1(\synth.voice.genblk4[2].next_state_scan[11] ),
    .B2(_05535_),
    .A2(net169),
    .A1(\synth.voice.genblk4[2].next_state_scan[13] ));
 sg13g2_nand2_1 _13645_ (.Y(_01229_),
    .A(_05687_),
    .B(_05688_));
 sg13g2_nor2_1 _13646_ (.A(_05401_),
    .B(_05371_),
    .Y(_05689_));
 sg13g2_nand2_1 _13647_ (.Y(_05690_),
    .A(_05660_),
    .B(_05689_));
 sg13g2_nor2_1 _13648_ (.A(_05690_),
    .B(_05639_),
    .Y(_05691_));
 sg13g2_nand2_1 _13649_ (.Y(_05692_),
    .A(_05584_),
    .B(_05691_));
 sg13g2_nand2_1 _13650_ (.Y(_05693_),
    .A(_05400_),
    .B(_05407_));
 sg13g2_nand2_1 _13651_ (.Y(_05694_),
    .A(_05693_),
    .B(_05399_));
 sg13g2_nand2_1 _13652_ (.Y(_05695_),
    .A(_05665_),
    .B(_05689_));
 sg13g2_nand2b_1 _13653_ (.Y(_05696_),
    .B(_05695_),
    .A_N(_05694_));
 sg13g2_nor2_1 _13654_ (.A(_05690_),
    .B(_05645_),
    .Y(_05697_));
 sg13g2_nor2_1 _13655_ (.A(_05696_),
    .B(_05697_),
    .Y(_05698_));
 sg13g2_nand2_1 _13656_ (.Y(_05699_),
    .A(_05692_),
    .B(_05698_));
 sg13g2_xnor2_1 _13657_ (.Y(_05700_),
    .A(_05390_),
    .B(_05699_));
 sg13g2_nand2_1 _13658_ (.Y(_05701_),
    .A(net71),
    .B(_05700_));
 sg13g2_nand2_1 _13659_ (.Y(_05702_),
    .A(_05701_),
    .B(net65));
 sg13g2_nand2_1 _13660_ (.Y(_05703_),
    .A(_05702_),
    .B(_05530_));
 sg13g2_a22oi_1 _13661_ (.Y(_05704_),
    .B1(\synth.voice.genblk4[2].next_state_scan[12] ),
    .B2(_05535_),
    .A2(net169),
    .A1(_03370_));
 sg13g2_nand2_1 _13662_ (.Y(_01230_),
    .A(_05703_),
    .B(_05704_));
 sg13g2_nor2_1 _13663_ (.A(_05403_),
    .B(_05222_),
    .Y(_05705_));
 sg13g2_nand2_1 _13664_ (.Y(_05706_),
    .A(_05592_),
    .B(_05705_));
 sg13g2_inv_1 _13665_ (.Y(_05707_),
    .A(_05403_));
 sg13g2_a21oi_1 _13666_ (.A1(_05218_),
    .A2(_05707_),
    .Y(_05708_),
    .B1(_05412_));
 sg13g2_nand2_1 _13667_ (.Y(_05709_),
    .A(_05706_),
    .B(_05708_));
 sg13g2_xnor2_1 _13668_ (.Y(_05710_),
    .A(_05342_),
    .B(_05709_));
 sg13g2_nand2_1 _13669_ (.Y(_05711_),
    .A(net71),
    .B(_05710_));
 sg13g2_nand2_1 _13670_ (.Y(_05712_),
    .A(_05711_),
    .B(net65));
 sg13g2_nand2_1 _13671_ (.Y(_05713_),
    .A(_05712_),
    .B(_05530_));
 sg13g2_a22oi_1 _13672_ (.Y(_05714_),
    .B1(\synth.voice.genblk4[2].next_state_scan[13] ),
    .B2(_05535_),
    .A2(net169),
    .A1(net401));
 sg13g2_nand2_1 _13673_ (.Y(_01231_),
    .A(_05713_),
    .B(_05714_));
 sg13g2_nor2_1 _13674_ (.A(_05390_),
    .B(_05342_),
    .Y(_05715_));
 sg13g2_nand2_1 _13675_ (.Y(_05716_),
    .A(_05715_),
    .B(_05689_));
 sg13g2_nor2_1 _13676_ (.A(_05716_),
    .B(_05661_),
    .Y(_05717_));
 sg13g2_nand2_1 _13677_ (.Y(_05718_),
    .A(_05615_),
    .B(_05717_));
 sg13g2_inv_1 _13678_ (.Y(_05719_),
    .A(_05716_));
 sg13g2_a21oi_1 _13679_ (.A1(_05341_),
    .A2(_05387_),
    .Y(_05720_),
    .B1(_05339_));
 sg13g2_a21o_1 _13680_ (.A2(_05694_),
    .A1(_05715_),
    .B1(_05720_),
    .X(_05721_));
 sg13g2_a21oi_1 _13681_ (.A1(_05667_),
    .A2(_05719_),
    .Y(_05722_),
    .B1(_05721_));
 sg13g2_nand3_1 _13682_ (.B(_05605_),
    .C(_05462_),
    .A(_05717_),
    .Y(_05723_));
 sg13g2_nand3_1 _13683_ (.B(_05722_),
    .C(_05723_),
    .A(_05718_),
    .Y(_05724_));
 sg13g2_nand2_1 _13684_ (.Y(_05725_),
    .A(_05724_),
    .B(_05333_));
 sg13g2_inv_1 _13685_ (.Y(_05726_),
    .A(_05333_));
 sg13g2_nand4_1 _13686_ (.B(_05722_),
    .C(_05726_),
    .A(_05718_),
    .Y(_05727_),
    .D(_05723_));
 sg13g2_nand2_1 _13687_ (.Y(_05728_),
    .A(_05725_),
    .B(_05727_));
 sg13g2_nand2_1 _13688_ (.Y(_05729_),
    .A(_05728_),
    .B(net71));
 sg13g2_nand2_1 _13689_ (.Y(_05730_),
    .A(_05729_),
    .B(net65));
 sg13g2_inv_1 _13690_ (.Y(_05731_),
    .A(_03607_));
 sg13g2_nand2_1 _13691_ (.Y(_05732_),
    .A(_03590_),
    .B(_04250_));
 sg13g2_o21ai_1 _13692_ (.B1(_05732_),
    .Y(_05733_),
    .A1(_04247_),
    .A2(_05731_));
 sg13g2_buf_1 _13693_ (.A(_05733_),
    .X(_05734_));
 sg13g2_buf_1 _13694_ (.A(_05734_),
    .X(_05735_));
 sg13g2_nor2b_1 _13695_ (.A(net168),
    .B_N(_05528_),
    .Y(_05736_));
 sg13g2_nand2_1 _13696_ (.Y(_05737_),
    .A(_05730_),
    .B(_05736_));
 sg13g2_buf_1 _13697_ (.A(net168),
    .X(_05738_));
 sg13g2_nor2_2 _13698_ (.A(_05528_),
    .B(net168),
    .Y(_05739_));
 sg13g2_a22oi_1 _13699_ (.Y(_05740_),
    .B1(\synth.voice.scan_outs[3][0] ),
    .B2(_05739_),
    .A2(net151),
    .A1(\synth.voice.genblk4[3].next_state_scan[0] ));
 sg13g2_nand2_1 _13700_ (.Y(_01232_),
    .A(_05737_),
    .B(_05740_));
 sg13g2_nand2_1 _13701_ (.Y(_05741_),
    .A(_05343_),
    .B(_05402_));
 sg13g2_nor2_1 _13702_ (.A(_05741_),
    .B(_05676_),
    .Y(_05742_));
 sg13g2_nand2_1 _13703_ (.Y(_05743_),
    .A(_05631_),
    .B(_05742_));
 sg13g2_a21oi_1 _13704_ (.A1(_05679_),
    .A2(_05408_),
    .Y(_05744_),
    .B1(_05741_));
 sg13g2_a21oi_1 _13705_ (.A1(_05343_),
    .A2(_05410_),
    .Y(_05745_),
    .B1(_05414_));
 sg13g2_nor2b_1 _13706_ (.A(_05744_),
    .B_N(_05745_),
    .Y(_05746_));
 sg13g2_nand3_1 _13707_ (.B(_05626_),
    .C(_05623_),
    .A(_05742_),
    .Y(_05747_));
 sg13g2_nand3_1 _13708_ (.B(_05746_),
    .C(_05747_),
    .A(_05743_),
    .Y(_05748_));
 sg13g2_nand2_1 _13709_ (.Y(_05749_),
    .A(_05748_),
    .B(_05353_));
 sg13g2_inv_1 _13710_ (.Y(_05750_),
    .A(_05353_));
 sg13g2_nand4_1 _13711_ (.B(_05750_),
    .C(_05746_),
    .A(_05743_),
    .Y(_05751_),
    .D(_05747_));
 sg13g2_nand2_1 _13712_ (.Y(_05752_),
    .A(_05749_),
    .B(_05751_));
 sg13g2_nand2_1 _13713_ (.Y(_05753_),
    .A(_05752_),
    .B(net71));
 sg13g2_nand2_1 _13714_ (.Y(_05754_),
    .A(_05753_),
    .B(net65));
 sg13g2_nand2_1 _13715_ (.Y(_05755_),
    .A(_05754_),
    .B(_05736_));
 sg13g2_a22oi_1 _13716_ (.Y(_05756_),
    .B1(\synth.voice.scan_outs[3][1] ),
    .B2(_05739_),
    .A2(net151),
    .A1(\synth.voice.genblk4[3].next_state_scan[1] ));
 sg13g2_nand2_1 _13717_ (.Y(_01233_),
    .A(_05755_),
    .B(_05756_));
 sg13g2_inv_1 _13718_ (.Y(_05757_),
    .A(\synth.voice.genblk4[0].next_state_scan[4] ));
 sg13g2_nor3_1 _13719_ (.A(_03668_),
    .B(_00053_),
    .C(_01737_),
    .Y(_05758_));
 sg13g2_inv_1 _13720_ (.Y(_05759_),
    .A(_05758_));
 sg13g2_inv_1 _13721_ (.Y(_05760_),
    .A(\synth.voice.coeff_index[1] ));
 sg13g2_o21ai_1 _13722_ (.B1(_05760_),
    .Y(_05761_),
    .A1(net242),
    .A2(_05759_));
 sg13g2_nor2_1 _13723_ (.A(_05760_),
    .B(_05759_),
    .Y(_05762_));
 sg13g2_nand2_1 _13724_ (.Y(_05763_),
    .A(_05762_),
    .B(_04200_));
 sg13g2_a21oi_1 _13725_ (.A1(_05761_),
    .A2(_05763_),
    .Y(_05764_),
    .B1(_03612_));
 sg13g2_a21oi_1 _13726_ (.A1(_05757_),
    .A2(_03612_),
    .Y(_01234_),
    .B1(_05764_));
 sg13g2_nor2_1 _13727_ (.A(_05333_),
    .B(_05353_),
    .Y(_05765_));
 sg13g2_nand2_1 _13728_ (.Y(_05766_),
    .A(_05715_),
    .B(_05765_));
 sg13g2_nor2_1 _13729_ (.A(_05766_),
    .B(_05690_),
    .Y(_05767_));
 sg13g2_nand2_1 _13730_ (.Y(_05768_),
    .A(_05646_),
    .B(_05767_));
 sg13g2_inv_1 _13731_ (.Y(_05769_),
    .A(_05766_));
 sg13g2_nand2_1 _13732_ (.Y(_05770_),
    .A(_05765_),
    .B(_05720_));
 sg13g2_nand2b_1 _13733_ (.Y(_05771_),
    .B(_05750_),
    .A_N(_05330_));
 sg13g2_nand3_1 _13734_ (.B(_05351_),
    .C(_05771_),
    .A(_05770_),
    .Y(_05772_));
 sg13g2_a21oi_1 _13735_ (.A1(_05696_),
    .A2(_05769_),
    .Y(_05773_),
    .B1(_05772_));
 sg13g2_nand3_1 _13736_ (.B(_05767_),
    .C(_05548_),
    .A(_05640_),
    .Y(_05774_));
 sg13g2_nand3_1 _13737_ (.B(_05773_),
    .C(_05774_),
    .A(_05768_),
    .Y(_05775_));
 sg13g2_nand2_1 _13738_ (.Y(_05776_),
    .A(_05775_),
    .B(_05361_));
 sg13g2_inv_1 _13739_ (.Y(_05777_),
    .A(_05361_));
 sg13g2_nand4_1 _13740_ (.B(_05777_),
    .C(_05773_),
    .A(_05768_),
    .Y(_05778_),
    .D(_05774_));
 sg13g2_nand2_1 _13741_ (.Y(_05779_),
    .A(_05776_),
    .B(_05778_));
 sg13g2_nand2_1 _13742_ (.Y(_05780_),
    .A(_05779_),
    .B(_05514_));
 sg13g2_nand2_1 _13743_ (.Y(_05781_),
    .A(_05780_),
    .B(_05522_));
 sg13g2_nand2_1 _13744_ (.Y(_05782_),
    .A(_05781_),
    .B(_05736_));
 sg13g2_a22oi_1 _13745_ (.Y(_05783_),
    .B1(\synth.voice.genblk4[3].next_state_scan[0] ),
    .B2(_05739_),
    .A2(net151),
    .A1(\synth.voice.genblk4[3].next_state_scan[2] ));
 sg13g2_nand2_1 _13746_ (.Y(_01235_),
    .A(_05782_),
    .B(_05783_));
 sg13g2_nand2b_1 _13747_ (.Y(_05784_),
    .B(_05520_),
    .A_N(_05512_));
 sg13g2_nand3_1 _13748_ (.B(_05519_),
    .C(_05736_),
    .A(_05784_),
    .Y(_05785_));
 sg13g2_a22oi_1 _13749_ (.Y(_05786_),
    .B1(\synth.voice.genblk4[3].next_state_scan[1] ),
    .B2(_05739_),
    .A2(net151),
    .A1(\synth.voice.genblk4[3].next_state_scan[3] ));
 sg13g2_nand2_1 _13750_ (.Y(_01236_),
    .A(_05785_),
    .B(_05786_));
 sg13g2_nor2b_1 _13751_ (.A(_03434_),
    .B_N(\synth.voice.target_reg[3] ),
    .Y(_05787_));
 sg13g2_nor2b_1 _13752_ (.A(_05734_),
    .B_N(_05787_),
    .Y(_05788_));
 sg13g2_buf_1 _13753_ (.A(_05788_),
    .X(_05789_));
 sg13g2_buf_1 _13754_ (.A(_05789_),
    .X(_05790_));
 sg13g2_nand2_1 _13755_ (.Y(_05791_),
    .A(_05524_),
    .B(net133));
 sg13g2_nor2_1 _13756_ (.A(_05787_),
    .B(net168),
    .Y(_05792_));
 sg13g2_buf_1 _13757_ (.A(_05792_),
    .X(_05793_));
 sg13g2_a22oi_1 _13758_ (.Y(_05794_),
    .B1(\synth.voice.genblk4[3].next_state_scan[2] ),
    .B2(net132),
    .A2(_05738_),
    .A1(\synth.voice.genblk4[3].next_state_scan[4] ));
 sg13g2_nand2_1 _13759_ (.Y(_01237_),
    .A(_05791_),
    .B(_05794_));
 sg13g2_nand2_1 _13760_ (.Y(_05795_),
    .A(_05540_),
    .B(net133));
 sg13g2_a22oi_1 _13761_ (.Y(_05796_),
    .B1(\synth.voice.genblk4[3].next_state_scan[3] ),
    .B2(net132),
    .A2(net151),
    .A1(\synth.voice.genblk4[3].next_state_scan[5] ));
 sg13g2_nand2_1 _13762_ (.Y(_01238_),
    .A(_05795_),
    .B(_05796_));
 sg13g2_nand2_1 _13763_ (.Y(_05797_),
    .A(_05551_),
    .B(net133));
 sg13g2_a22oi_1 _13764_ (.Y(_05798_),
    .B1(\synth.voice.genblk4[3].next_state_scan[4] ),
    .B2(net132),
    .A2(net151),
    .A1(\synth.voice.genblk4[3].next_state_scan[6] ));
 sg13g2_nand2_1 _13765_ (.Y(_01239_),
    .A(_05797_),
    .B(_05798_));
 sg13g2_nand2_1 _13766_ (.Y(_05799_),
    .A(_05556_),
    .B(net133));
 sg13g2_a22oi_1 _13767_ (.Y(_05800_),
    .B1(\synth.voice.genblk4[3].next_state_scan[5] ),
    .B2(net132),
    .A2(net151),
    .A1(\synth.voice.genblk4[3].next_state_scan[7] ));
 sg13g2_nand2_1 _13768_ (.Y(_01240_),
    .A(_05799_),
    .B(_05800_));
 sg13g2_nand2_1 _13769_ (.Y(_05801_),
    .A(_05567_),
    .B(_05790_));
 sg13g2_a22oi_1 _13770_ (.Y(_05802_),
    .B1(\synth.voice.genblk4[3].next_state_scan[6] ),
    .B2(_05793_),
    .A2(_05738_),
    .A1(\synth.voice.genblk4[3].next_state_scan[8] ));
 sg13g2_nand2_1 _13771_ (.Y(_01241_),
    .A(_05801_),
    .B(_05802_));
 sg13g2_nand2_1 _13772_ (.Y(_05803_),
    .A(_05574_),
    .B(_05790_));
 sg13g2_a22oi_1 _13773_ (.Y(_05804_),
    .B1(\synth.voice.genblk4[3].next_state_scan[7] ),
    .B2(_05793_),
    .A2(net151),
    .A1(\synth.voice.genblk4[3].next_state_scan[9] ));
 sg13g2_nand2_1 _13774_ (.Y(_01242_),
    .A(_05803_),
    .B(_05804_));
 sg13g2_nand2_1 _13775_ (.Y(_05805_),
    .A(_05587_),
    .B(net133));
 sg13g2_a22oi_1 _13776_ (.Y(_05806_),
    .B1(\synth.voice.genblk4[3].next_state_scan[8] ),
    .B2(net132),
    .A2(net168),
    .A1(\synth.voice.genblk4[3].next_state_scan[10] ));
 sg13g2_nand2_1 _13777_ (.Y(_01243_),
    .A(_05805_),
    .B(_05806_));
 sg13g2_nand2_1 _13778_ (.Y(_05807_),
    .A(_05595_),
    .B(net133));
 sg13g2_a22oi_1 _13779_ (.Y(_05808_),
    .B1(\synth.voice.genblk4[3].next_state_scan[9] ),
    .B2(net132),
    .A2(net168),
    .A1(\synth.voice.genblk4[3].next_state_scan[11] ));
 sg13g2_nand2_1 _13780_ (.Y(_01244_),
    .A(_05807_),
    .B(_05808_));
 sg13g2_inv_1 _13781_ (.Y(_05809_),
    .A(\synth.voice.coeff_index[2] ));
 sg13g2_xnor2_1 _13782_ (.Y(_05810_),
    .A(_05809_),
    .B(_05763_));
 sg13g2_nor2_1 _13783_ (.A(\synth.voice.genblk4[0].next_state_scan[5] ),
    .B(net189),
    .Y(_05811_));
 sg13g2_a21oi_1 _13784_ (.A1(_05810_),
    .A2(net189),
    .Y(_01245_),
    .B1(_05811_));
 sg13g2_nand2_1 _13785_ (.Y(_05812_),
    .A(_05619_),
    .B(net133));
 sg13g2_a22oi_1 _13786_ (.Y(_05813_),
    .B1(\synth.voice.genblk4[3].next_state_scan[10] ),
    .B2(net132),
    .A2(_05735_),
    .A1(\synth.voice.genblk4[3].next_state_scan[12] ));
 sg13g2_nand2_1 _13787_ (.Y(_01246_),
    .A(_05812_),
    .B(_05813_));
 sg13g2_nand2_1 _13788_ (.Y(_05814_),
    .A(_05635_),
    .B(net133));
 sg13g2_a22oi_1 _13789_ (.Y(_05815_),
    .B1(\synth.voice.genblk4[3].next_state_scan[11] ),
    .B2(net132),
    .A2(_05735_),
    .A1(\synth.voice.genblk4[3].next_state_scan[13] ));
 sg13g2_nand2_1 _13790_ (.Y(_01247_),
    .A(_05814_),
    .B(_05815_));
 sg13g2_nand2_1 _13791_ (.Y(_05816_),
    .A(_05650_),
    .B(_05789_));
 sg13g2_a22oi_1 _13792_ (.Y(_05817_),
    .B1(\synth.voice.genblk4[3].next_state_scan[12] ),
    .B2(_05792_),
    .A2(net168),
    .A1(_03370_));
 sg13g2_nand2_1 _13793_ (.Y(_01248_),
    .A(_05816_),
    .B(_05817_));
 sg13g2_nand2_1 _13794_ (.Y(_05818_),
    .A(_05657_),
    .B(_05789_));
 sg13g2_a22oi_1 _13795_ (.Y(_05819_),
    .B1(\synth.voice.genblk4[3].next_state_scan[13] ),
    .B2(_05792_),
    .A2(net168),
    .A1(_03379_));
 sg13g2_nand2_1 _13796_ (.Y(_01249_),
    .A(_05818_),
    .B(_05819_));
 sg13g2_inv_1 _13797_ (.Y(_05820_),
    .A(_03595_));
 sg13g2_nor2_1 _13798_ (.A(_05820_),
    .B(_04026_),
    .Y(_05821_));
 sg13g2_a21oi_1 _13799_ (.A1(_03603_),
    .A2(_04023_),
    .Y(_05822_),
    .B1(_05821_));
 sg13g2_buf_1 _13800_ (.A(_05822_),
    .X(_05823_));
 sg13g2_inv_1 _13801_ (.Y(_05824_),
    .A(_05823_));
 sg13g2_nor2b_1 _13802_ (.A(_05824_),
    .B_N(_05787_),
    .Y(_05825_));
 sg13g2_buf_2 _13803_ (.A(_05825_),
    .X(_05826_));
 sg13g2_nand2_1 _13804_ (.Y(_05827_),
    .A(_05673_),
    .B(_05826_));
 sg13g2_buf_1 _13805_ (.A(_05824_),
    .X(_05828_));
 sg13g2_buf_1 _13806_ (.A(_05828_),
    .X(_05829_));
 sg13g2_nor2_1 _13807_ (.A(_05787_),
    .B(_05824_),
    .Y(_05830_));
 sg13g2_buf_2 _13808_ (.A(_05830_),
    .X(_05831_));
 sg13g2_a22oi_1 _13809_ (.Y(_05832_),
    .B1(_05047_),
    .B2(_05831_),
    .A2(net124),
    .A1(\synth.voice.genblk4[4].next_state_scan[0] ));
 sg13g2_nand2_1 _13810_ (.Y(_01250_),
    .A(_05827_),
    .B(_05832_));
 sg13g2_nand2_1 _13811_ (.Y(_05833_),
    .A(_05686_),
    .B(_05826_));
 sg13g2_a22oi_1 _13812_ (.Y(_05834_),
    .B1(_05040_),
    .B2(_05831_),
    .A2(net124),
    .A1(\synth.voice.genblk4[4].next_state_scan[1] ));
 sg13g2_nand2_1 _13813_ (.Y(_01251_),
    .A(_05833_),
    .B(_05834_));
 sg13g2_nand2_1 _13814_ (.Y(_05835_),
    .A(_05702_),
    .B(_05826_));
 sg13g2_a22oi_1 _13815_ (.Y(_05836_),
    .B1(\synth.voice.genblk4[4].next_state_scan[0] ),
    .B2(_05831_),
    .A2(net124),
    .A1(_05090_));
 sg13g2_nand2_1 _13816_ (.Y(_01252_),
    .A(_05835_),
    .B(_05836_));
 sg13g2_nand2_1 _13817_ (.Y(_05837_),
    .A(_05712_),
    .B(_05826_));
 sg13g2_a22oi_1 _13818_ (.Y(_05838_),
    .B1(\synth.voice.genblk4[4].next_state_scan[1] ),
    .B2(_05831_),
    .A2(net124),
    .A1(\synth.voice.genblk4[4].next_state_scan[3] ));
 sg13g2_nand2_1 _13819_ (.Y(_01253_),
    .A(_05837_),
    .B(_05838_));
 sg13g2_nand2_1 _13820_ (.Y(_05839_),
    .A(_05730_),
    .B(_05826_));
 sg13g2_a22oi_1 _13821_ (.Y(_05840_),
    .B1(_05090_),
    .B2(_05831_),
    .A2(net124),
    .A1(_05015_));
 sg13g2_nand2_1 _13822_ (.Y(_01254_),
    .A(_05839_),
    .B(_05840_));
 sg13g2_nand2_1 _13823_ (.Y(_05841_),
    .A(_05754_),
    .B(_05826_));
 sg13g2_a22oi_1 _13824_ (.Y(_05842_),
    .B1(\synth.voice.genblk4[4].next_state_scan[3] ),
    .B2(_05831_),
    .A2(net124),
    .A1(_05005_));
 sg13g2_nand2_1 _13825_ (.Y(_01255_),
    .A(_05841_),
    .B(_05842_));
 sg13g2_inv_1 _13826_ (.Y(_05843_),
    .A(\synth.voice.genblk4[0].next_state_scan[6] ));
 sg13g2_nor2_1 _13827_ (.A(_05843_),
    .B(net189),
    .Y(_05844_));
 sg13g2_a21oi_1 _13828_ (.A1(_04782_),
    .A2(net189),
    .Y(_05845_),
    .B1(_05844_));
 sg13g2_nor2_1 _13829_ (.A(\synth.voice.genblk4[0].next_state_scan[4] ),
    .B(_04207_),
    .Y(_05846_));
 sg13g2_a21oi_1 _13830_ (.A1(net44),
    .A2(_05845_),
    .Y(_01256_),
    .B1(_05846_));
 sg13g2_nand2_1 _13831_ (.Y(_05847_),
    .A(_05781_),
    .B(_05826_));
 sg13g2_a22oi_1 _13832_ (.Y(_05848_),
    .B1(_05015_),
    .B2(_05831_),
    .A2(_05829_),
    .A1(\synth.voice.float_period[0][0] ));
 sg13g2_nand2_1 _13833_ (.Y(_01257_),
    .A(_05847_),
    .B(_05848_));
 sg13g2_nand3_1 _13834_ (.B(_05519_),
    .C(_05826_),
    .A(_05784_),
    .Y(_05849_));
 sg13g2_a22oi_1 _13835_ (.Y(_05850_),
    .B1(_05005_),
    .B2(_05831_),
    .A2(_05829_),
    .A1(\synth.voice.float_period[0][1] ));
 sg13g2_nand2_1 _13836_ (.Y(_01258_),
    .A(_05849_),
    .B(_05850_));
 sg13g2_nor3_1 _13837_ (.A(net400),
    .B(_03810_),
    .C(_03727_),
    .Y(_05851_));
 sg13g2_nand3_1 _13838_ (.B(_04016_),
    .C(_05851_),
    .A(_04013_),
    .Y(_05852_));
 sg13g2_buf_2 _13839_ (.A(_05852_),
    .X(_05853_));
 sg13g2_nand2_1 _13840_ (.Y(_05854_),
    .A(_05853_),
    .B(_05823_));
 sg13g2_buf_2 _13841_ (.A(_05854_),
    .X(_05855_));
 sg13g2_nand3_1 _13842_ (.B(_03735_),
    .C(_03814_),
    .A(_03834_),
    .Y(_05856_));
 sg13g2_nor2_1 _13843_ (.A(_03765_),
    .B(net328),
    .Y(_05857_));
 sg13g2_a21oi_1 _13844_ (.A1(_05856_),
    .A2(net328),
    .Y(_05858_),
    .B1(_05857_));
 sg13g2_buf_1 _13845_ (.A(_05823_),
    .X(_05859_));
 sg13g2_mux2_1 _13846_ (.A0(\synth.voice.float_period[0][2] ),
    .A1(_05858_),
    .S(net150),
    .X(_05860_));
 sg13g2_nand2_1 _13847_ (.Y(_05861_),
    .A(_05855_),
    .B(_05860_));
 sg13g2_buf_1 _13848_ (.A(_05853_),
    .X(_05862_));
 sg13g2_nand3_1 _13849_ (.B(\synth.voice.float_period[0][0] ),
    .C(net150),
    .A(net33),
    .Y(_05863_));
 sg13g2_nand2_1 _13850_ (.Y(_01259_),
    .A(_05861_),
    .B(_05863_));
 sg13g2_xnor2_1 _13851_ (.Y(_05864_),
    .A(_03814_),
    .B(_04050_));
 sg13g2_inv_1 _13852_ (.Y(_05865_),
    .A(\synth.controller.reg_wdata[1] ));
 sg13g2_nor2_1 _13853_ (.A(net328),
    .B(_05865_),
    .Y(_05866_));
 sg13g2_a21oi_1 _13854_ (.A1(_05864_),
    .A2(net328),
    .Y(_05867_),
    .B1(_05866_));
 sg13g2_nand2_1 _13855_ (.Y(_05868_),
    .A(net131),
    .B(\synth.voice.float_period[0][3] ));
 sg13g2_o21ai_1 _13856_ (.B1(_05868_),
    .Y(_05869_),
    .A1(net124),
    .A2(_05867_));
 sg13g2_nand2_1 _13857_ (.Y(_05870_),
    .A(_05855_),
    .B(_05869_));
 sg13g2_nand3_1 _13858_ (.B(\synth.voice.float_period[0][1] ),
    .C(net150),
    .A(net33),
    .Y(_05871_));
 sg13g2_nand2_1 _13859_ (.Y(_01260_),
    .A(_05870_),
    .B(_05871_));
 sg13g2_xnor2_1 _13860_ (.Y(_05872_),
    .A(_03853_),
    .B(_03859_));
 sg13g2_inv_1 _13861_ (.Y(_05873_),
    .A(_03750_));
 sg13g2_nor2_1 _13862_ (.A(net328),
    .B(_05873_),
    .Y(_05874_));
 sg13g2_a21oi_1 _13863_ (.A1(_05872_),
    .A2(net328),
    .Y(_05875_),
    .B1(_05874_));
 sg13g2_nand2_1 _13864_ (.Y(_05876_),
    .A(net131),
    .B(_03746_));
 sg13g2_o21ai_1 _13865_ (.B1(_05876_),
    .Y(_05877_),
    .A1(net124),
    .A2(_05875_));
 sg13g2_nand2_1 _13866_ (.Y(_05878_),
    .A(_05855_),
    .B(_05877_));
 sg13g2_nand3_1 _13867_ (.B(\synth.voice.float_period[0][2] ),
    .C(net150),
    .A(net33),
    .Y(_05879_));
 sg13g2_nand2_1 _13868_ (.Y(_01261_),
    .A(_05878_),
    .B(_05879_));
 sg13g2_xor2_1 _13869_ (.B(_04138_),
    .A(_03852_),
    .X(_05880_));
 sg13g2_nor2_1 _13870_ (.A(net328),
    .B(_03782_),
    .Y(_05881_));
 sg13g2_a21oi_1 _13871_ (.A1(_05880_),
    .A2(_04087_),
    .Y(_05882_),
    .B1(_05881_));
 sg13g2_nand2_1 _13872_ (.Y(_05883_),
    .A(net131),
    .B(\synth.voice.float_period[0][5] ));
 sg13g2_o21ai_1 _13873_ (.B1(_05883_),
    .Y(_05884_),
    .A1(net131),
    .A2(_05882_));
 sg13g2_nand2_1 _13874_ (.Y(_05885_),
    .A(_05855_),
    .B(_05884_));
 sg13g2_nand3_1 _13875_ (.B(\synth.voice.float_period[0][3] ),
    .C(net150),
    .A(net33),
    .Y(_05886_));
 sg13g2_nand2_1 _13876_ (.Y(_01262_),
    .A(_05885_),
    .B(_05886_));
 sg13g2_nand2_1 _13877_ (.Y(_05887_),
    .A(net131),
    .B(\synth.voice.float_period[0][6] ));
 sg13g2_o21ai_1 _13878_ (.B1(_05887_),
    .Y(_05888_),
    .A1(net131),
    .A2(_04041_));
 sg13g2_nand2_1 _13879_ (.Y(_05889_),
    .A(_05855_),
    .B(_05888_));
 sg13g2_nand3_1 _13880_ (.B(_03746_),
    .C(net150),
    .A(net33),
    .Y(_05890_));
 sg13g2_nand2_1 _13881_ (.Y(_01263_),
    .A(_05889_),
    .B(_05890_));
 sg13g2_nand2_1 _13882_ (.Y(_05891_),
    .A(_05828_),
    .B(\synth.voice.float_period[0][7] ));
 sg13g2_o21ai_1 _13883_ (.B1(_05891_),
    .Y(_05892_),
    .A1(net131),
    .A2(_04064_));
 sg13g2_nand2_1 _13884_ (.Y(_05893_),
    .A(_05855_),
    .B(_05892_));
 sg13g2_nand3_1 _13885_ (.B(\synth.voice.float_period[0][5] ),
    .C(_05859_),
    .A(_05862_),
    .Y(_05894_));
 sg13g2_nand2_1 _13886_ (.Y(_01264_),
    .A(_05893_),
    .B(_05894_));
 sg13g2_nand3_1 _13887_ (.B(_04075_),
    .C(_05823_),
    .A(_04073_),
    .Y(_05895_));
 sg13g2_o21ai_1 _13888_ (.B1(_05895_),
    .Y(_05896_),
    .A1(net377),
    .A2(net150));
 sg13g2_nand2_1 _13889_ (.Y(_05897_),
    .A(_05855_),
    .B(_05896_));
 sg13g2_nand3_1 _13890_ (.B(\synth.voice.float_period[0][6] ),
    .C(_05859_),
    .A(net33),
    .Y(_05898_));
 sg13g2_nand2_1 _13891_ (.Y(_01265_),
    .A(_05897_),
    .B(_05898_));
 sg13g2_nand3_1 _13892_ (.B(_04089_),
    .C(_05823_),
    .A(_04088_),
    .Y(_05899_));
 sg13g2_nand2_1 _13893_ (.Y(_05900_),
    .A(net131),
    .B(net401));
 sg13g2_nand2_1 _13894_ (.Y(_05901_),
    .A(_05899_),
    .B(_05900_));
 sg13g2_nand2_1 _13895_ (.Y(_05902_),
    .A(_05855_),
    .B(_05901_));
 sg13g2_nand3_1 _13896_ (.B(\synth.voice.float_period[0][7] ),
    .C(net150),
    .A(_05862_),
    .Y(_05903_));
 sg13g2_nand2_1 _13897_ (.Y(_01266_),
    .A(_05902_),
    .B(_05903_));
 sg13g2_inv_1 _13898_ (.Y(_05904_),
    .A(\synth.voice.genblk4[0].next_state_scan[7] ));
 sg13g2_nor2_1 _13899_ (.A(_05904_),
    .B(_03609_),
    .Y(_05905_));
 sg13g2_a21oi_1 _13900_ (.A1(_04825_),
    .A2(net189),
    .Y(_05906_),
    .B1(_05905_));
 sg13g2_nor2_1 _13901_ (.A(\synth.voice.genblk4[0].next_state_scan[5] ),
    .B(net43),
    .Y(_05907_));
 sg13g2_a21oi_1 _13902_ (.A1(_04206_),
    .A2(_05906_),
    .Y(_01267_),
    .B1(_05907_));
 sg13g2_nor2_1 _13903_ (.A(_04784_),
    .B(_04026_),
    .Y(_05908_));
 sg13g2_a21oi_1 _13904_ (.A1(_04023_),
    .A2(_04783_),
    .Y(_05909_),
    .B1(_05908_));
 sg13g2_buf_1 _13905_ (.A(_05909_),
    .X(_05910_));
 sg13g2_buf_1 _13906_ (.A(net167),
    .X(_05911_));
 sg13g2_nand2_2 _13907_ (.Y(_05912_),
    .A(_05853_),
    .B(net149));
 sg13g2_nand3_1 _13908_ (.B(_04100_),
    .C(net167),
    .A(_04099_),
    .Y(_05913_));
 sg13g2_inv_1 _13909_ (.Y(_05914_),
    .A(_05909_));
 sg13g2_buf_1 _13910_ (.A(net166),
    .X(_05915_));
 sg13g2_nand2_1 _13911_ (.Y(_05916_),
    .A(net148),
    .B(\synth.voice.float_period[0][10] ));
 sg13g2_nand2_1 _13912_ (.Y(_05917_),
    .A(_05913_),
    .B(_05916_));
 sg13g2_nand2_1 _13913_ (.Y(_05918_),
    .A(_05912_),
    .B(_05917_));
 sg13g2_buf_1 _13914_ (.A(net149),
    .X(_05919_));
 sg13g2_nand3_1 _13915_ (.B(\synth.voice.float_period[0][8] ),
    .C(net130),
    .A(net33),
    .Y(_05920_));
 sg13g2_nand2_1 _13916_ (.Y(_01268_),
    .A(_05918_),
    .B(_05920_));
 sg13g2_nand3_1 _13917_ (.B(_04118_),
    .C(net167),
    .A(_04117_),
    .Y(_05921_));
 sg13g2_nand2_1 _13918_ (.Y(_05922_),
    .A(net148),
    .B(\synth.voice.float_period[0][11] ));
 sg13g2_nand2_1 _13919_ (.Y(_05923_),
    .A(_05921_),
    .B(_05922_));
 sg13g2_nand2_1 _13920_ (.Y(_05924_),
    .A(_05912_),
    .B(_05923_));
 sg13g2_nand3_1 _13921_ (.B(\synth.voice.float_period[0][9] ),
    .C(net130),
    .A(net33),
    .Y(_05925_));
 sg13g2_nand2_1 _13922_ (.Y(_01269_),
    .A(_05924_),
    .B(_05925_));
 sg13g2_nand3_1 _13923_ (.B(_04128_),
    .C(_05910_),
    .A(_04127_),
    .Y(_05926_));
 sg13g2_nand2_1 _13924_ (.Y(_05927_),
    .A(net148),
    .B(\synth.voice.float_period[0][12] ));
 sg13g2_nand2_1 _13925_ (.Y(_05928_),
    .A(_05926_),
    .B(_05927_));
 sg13g2_nand2_1 _13926_ (.Y(_05929_),
    .A(_05912_),
    .B(_05928_));
 sg13g2_nand3_1 _13927_ (.B(\synth.voice.float_period[0][10] ),
    .C(net130),
    .A(_05853_),
    .Y(_05930_));
 sg13g2_nand2_1 _13928_ (.Y(_01270_),
    .A(_05929_),
    .B(_05930_));
 sg13g2_nand3_1 _13929_ (.B(_04150_),
    .C(net167),
    .A(_04148_),
    .Y(_05931_));
 sg13g2_nand2_1 _13930_ (.Y(_05932_),
    .A(net148),
    .B(\synth.voice.float_period[0][13] ));
 sg13g2_nand2_1 _13931_ (.Y(_05933_),
    .A(_05931_),
    .B(_05932_));
 sg13g2_nand2_1 _13932_ (.Y(_05934_),
    .A(_05912_),
    .B(_05933_));
 sg13g2_nand3_1 _13933_ (.B(\synth.voice.float_period[0][11] ),
    .C(net130),
    .A(_05853_),
    .Y(_05935_));
 sg13g2_nand2_1 _13934_ (.Y(_01271_),
    .A(_05934_),
    .B(_05935_));
 sg13g2_nand3_1 _13935_ (.B(_04169_),
    .C(_05910_),
    .A(_04167_),
    .Y(_05936_));
 sg13g2_nand2_1 _13936_ (.Y(_05937_),
    .A(_05915_),
    .B(\synth.voice.float_period[1][0] ));
 sg13g2_nand2_1 _13937_ (.Y(_05938_),
    .A(_05936_),
    .B(_05937_));
 sg13g2_nand2_1 _13938_ (.Y(_05939_),
    .A(_05912_),
    .B(_05938_));
 sg13g2_nand3_1 _13939_ (.B(\synth.voice.float_period[0][12] ),
    .C(net130),
    .A(_05853_),
    .Y(_05940_));
 sg13g2_nand2_1 _13940_ (.Y(_01272_),
    .A(_05939_),
    .B(_05940_));
 sg13g2_nand3_1 _13941_ (.B(_04189_),
    .C(net167),
    .A(_04187_),
    .Y(_05941_));
 sg13g2_nand2_1 _13942_ (.Y(_05942_),
    .A(_05914_),
    .B(\synth.voice.float_period[1][1] ));
 sg13g2_nand2_1 _13943_ (.Y(_05943_),
    .A(_05941_),
    .B(_05942_));
 sg13g2_nand2_1 _13944_ (.Y(_05944_),
    .A(_05912_),
    .B(_05943_));
 sg13g2_nand3_1 _13945_ (.B(\synth.voice.float_period[0][13] ),
    .C(_05919_),
    .A(_05853_),
    .Y(_05945_));
 sg13g2_nand2_1 _13946_ (.Y(_01273_),
    .A(_05944_),
    .B(_05945_));
 sg13g2_nor2_1 _13947_ (.A(_03727_),
    .B(_03426_),
    .Y(_05946_));
 sg13g2_nand3_1 _13948_ (.B(_04016_),
    .C(_05946_),
    .A(_04013_),
    .Y(_05947_));
 sg13g2_buf_2 _13949_ (.A(_05947_),
    .X(_05948_));
 sg13g2_nand2_1 _13950_ (.Y(_05949_),
    .A(_05948_),
    .B(net167));
 sg13g2_buf_1 _13951_ (.A(_05949_),
    .X(_05950_));
 sg13g2_mux2_1 _13952_ (.A0(\synth.voice.float_period[1][2] ),
    .A1(_05858_),
    .S(net149),
    .X(_05951_));
 sg13g2_nand2_1 _13953_ (.Y(_05952_),
    .A(net29),
    .B(_05951_));
 sg13g2_buf_1 _13954_ (.A(_05948_),
    .X(_05953_));
 sg13g2_nand3_1 _13955_ (.B(\synth.voice.float_period[1][0] ),
    .C(net130),
    .A(net32),
    .Y(_05954_));
 sg13g2_nand2_1 _13956_ (.Y(_01274_),
    .A(_05952_),
    .B(_05954_));
 sg13g2_nand2_1 _13957_ (.Y(_05955_),
    .A(net166),
    .B(\synth.voice.float_period[1][3] ));
 sg13g2_o21ai_1 _13958_ (.B1(_05955_),
    .Y(_05956_),
    .A1(net148),
    .A2(_05867_));
 sg13g2_nand2_1 _13959_ (.Y(_05957_),
    .A(net29),
    .B(_05956_));
 sg13g2_nand3_1 _13960_ (.B(\synth.voice.float_period[1][1] ),
    .C(net130),
    .A(net32),
    .Y(_05958_));
 sg13g2_nand2_1 _13961_ (.Y(_01275_),
    .A(_05957_),
    .B(_05958_));
 sg13g2_nand2_1 _13962_ (.Y(_05959_),
    .A(net166),
    .B(\synth.voice.float_period[1][4] ));
 sg13g2_o21ai_1 _13963_ (.B1(_05959_),
    .Y(_05960_),
    .A1(net148),
    .A2(_05875_));
 sg13g2_nand2_1 _13964_ (.Y(_05961_),
    .A(_05950_),
    .B(_05960_));
 sg13g2_nand3_1 _13965_ (.B(\synth.voice.float_period[1][2] ),
    .C(net130),
    .A(net32),
    .Y(_05962_));
 sg13g2_nand2_1 _13966_ (.Y(_01276_),
    .A(_05961_),
    .B(_05962_));
 sg13g2_nand2_1 _13967_ (.Y(_05963_),
    .A(net166),
    .B(_03732_));
 sg13g2_o21ai_1 _13968_ (.B1(_05963_),
    .Y(_05964_),
    .A1(net148),
    .A2(_05882_));
 sg13g2_nand2_1 _13969_ (.Y(_05965_),
    .A(_05950_),
    .B(_05964_));
 sg13g2_nand3_1 _13970_ (.B(\synth.voice.float_period[1][3] ),
    .C(_05919_),
    .A(net32),
    .Y(_05966_));
 sg13g2_nand2_1 _13971_ (.Y(_01277_),
    .A(_05965_),
    .B(_05966_));
 sg13g2_nand2_1 _13972_ (.Y(_05967_),
    .A(net180),
    .B(\synth.voice.genblk4[0].next_state_scan[8] ));
 sg13g2_o21ai_1 _13973_ (.B1(_05967_),
    .Y(_05968_),
    .A1(net180),
    .A2(_04843_));
 sg13g2_nand2_1 _13974_ (.Y(_05969_),
    .A(_04207_),
    .B(_05968_));
 sg13g2_o21ai_1 _13975_ (.B1(_05969_),
    .Y(_01278_),
    .A1(_05843_),
    .A2(_04206_));
 sg13g2_nand2_1 _13976_ (.Y(_05970_),
    .A(net166),
    .B(_03762_));
 sg13g2_o21ai_1 _13977_ (.B1(_05970_),
    .Y(_05971_),
    .A1(net148),
    .A2(_04041_));
 sg13g2_nand2_1 _13978_ (.Y(_05972_),
    .A(net29),
    .B(_05971_));
 sg13g2_nand3_1 _13979_ (.B(\synth.voice.float_period[1][4] ),
    .C(_05911_),
    .A(_05953_),
    .Y(_05973_));
 sg13g2_nand2_1 _13980_ (.Y(_01279_),
    .A(_05972_),
    .B(_05973_));
 sg13g2_nand2_1 _13981_ (.Y(_05974_),
    .A(_05914_),
    .B(_03863_));
 sg13g2_o21ai_1 _13982_ (.B1(_05974_),
    .Y(_05975_),
    .A1(_05915_),
    .A2(_04064_));
 sg13g2_nand2_1 _13983_ (.Y(_05976_),
    .A(net29),
    .B(_05975_));
 sg13g2_nand3_1 _13984_ (.B(_03732_),
    .C(net149),
    .A(net32),
    .Y(_05977_));
 sg13g2_nand2_1 _13985_ (.Y(_01280_),
    .A(_05976_),
    .B(_05977_));
 sg13g2_nand3_1 _13986_ (.B(_04075_),
    .C(net167),
    .A(_04073_),
    .Y(_05978_));
 sg13g2_o21ai_1 _13987_ (.B1(_05978_),
    .Y(_05979_),
    .A1(_04897_),
    .A2(_05911_));
 sg13g2_nand2_1 _13988_ (.Y(_05980_),
    .A(net29),
    .B(_05979_));
 sg13g2_nand3_1 _13989_ (.B(_03762_),
    .C(net149),
    .A(_05953_),
    .Y(_05981_));
 sg13g2_nand2_1 _13990_ (.Y(_01281_),
    .A(_05980_),
    .B(_05981_));
 sg13g2_nand3_1 _13991_ (.B(_04089_),
    .C(net167),
    .A(_04088_),
    .Y(_05982_));
 sg13g2_nand2_1 _13992_ (.Y(_05983_),
    .A(net166),
    .B(_03874_));
 sg13g2_nand2_1 _13993_ (.Y(_05984_),
    .A(_05982_),
    .B(_05983_));
 sg13g2_nand2_1 _13994_ (.Y(_05985_),
    .A(net29),
    .B(_05984_));
 sg13g2_nand3_1 _13995_ (.B(_03863_),
    .C(net149),
    .A(net32),
    .Y(_05986_));
 sg13g2_nand2_1 _13996_ (.Y(_01282_),
    .A(_05985_),
    .B(_05986_));
 sg13g2_nand2_1 _13997_ (.Y(_05987_),
    .A(net166),
    .B(_03370_));
 sg13g2_nand2_1 _13998_ (.Y(_05988_),
    .A(_05913_),
    .B(_05987_));
 sg13g2_nand2_1 _13999_ (.Y(_05989_),
    .A(net29),
    .B(_05988_));
 sg13g2_nand3_1 _14000_ (.B(\synth.voice.float_period[1][8] ),
    .C(net149),
    .A(net32),
    .Y(_05990_));
 sg13g2_nand2_1 _14001_ (.Y(_01283_),
    .A(_05989_),
    .B(_05990_));
 sg13g2_nand2_1 _14002_ (.Y(_05991_),
    .A(net166),
    .B(net401));
 sg13g2_nand2_1 _14003_ (.Y(_05992_),
    .A(_05921_),
    .B(_05991_));
 sg13g2_nand2_1 _14004_ (.Y(_05993_),
    .A(net29),
    .B(_05992_));
 sg13g2_nand3_1 _14005_ (.B(_03874_),
    .C(net149),
    .A(net32),
    .Y(_05994_));
 sg13g2_nand2_1 _14006_ (.Y(_01284_),
    .A(_05993_),
    .B(_05994_));
 sg13g2_nand2_1 _14007_ (.Y(_05995_),
    .A(_05948_),
    .B(net157));
 sg13g2_nand2_1 _14008_ (.Y(_05996_),
    .A(_04092_),
    .B(\synth.voice.float_period[1][12] ));
 sg13g2_nand2_1 _14009_ (.Y(_05997_),
    .A(_04129_),
    .B(_05996_));
 sg13g2_nand2_1 _14010_ (.Y(_05998_),
    .A(_05995_),
    .B(_05997_));
 sg13g2_nand3_1 _14011_ (.B(_03451_),
    .C(net158),
    .A(_05948_),
    .Y(_05999_));
 sg13g2_nand2_1 _14012_ (.Y(_01285_),
    .A(_05998_),
    .B(_05999_));
 sg13g2_nand2_1 _14013_ (.Y(_06000_),
    .A(_04092_),
    .B(\synth.voice.float_period[1][13] ));
 sg13g2_nand2_1 _14014_ (.Y(_06001_),
    .A(_04151_),
    .B(_06000_));
 sg13g2_nand2_1 _14015_ (.Y(_06002_),
    .A(_05995_),
    .B(_06001_));
 sg13g2_nand3_1 _14016_ (.B(\synth.voice.float_period[1][11] ),
    .C(net158),
    .A(_05948_),
    .Y(_06003_));
 sg13g2_nand2_1 _14017_ (.Y(_01286_),
    .A(_06002_),
    .B(_06003_));
 sg13g2_nand2_1 _14018_ (.Y(_06004_),
    .A(net140),
    .B(_03818_));
 sg13g2_nand2_1 _14019_ (.Y(_06005_),
    .A(_04170_),
    .B(_06004_));
 sg13g2_nand2_1 _14020_ (.Y(_06006_),
    .A(_05995_),
    .B(_06005_));
 sg13g2_nand3_1 _14021_ (.B(\synth.voice.float_period[1][12] ),
    .C(_04036_),
    .A(_05948_),
    .Y(_06007_));
 sg13g2_nand2_1 _14022_ (.Y(_01287_),
    .A(_06006_),
    .B(_06007_));
 sg13g2_nand2_1 _14023_ (.Y(_06008_),
    .A(_04091_),
    .B(\synth.voice.genblk4[6].next_state_scan[3] ));
 sg13g2_nand2_1 _14024_ (.Y(_06009_),
    .A(_04190_),
    .B(_06008_));
 sg13g2_nand2_1 _14025_ (.Y(_06010_),
    .A(_05995_),
    .B(_06009_));
 sg13g2_nand3_1 _14026_ (.B(\synth.voice.float_period[1][13] ),
    .C(_04036_),
    .A(_05948_),
    .Y(_06011_));
 sg13g2_nand2_1 _14027_ (.Y(_01288_),
    .A(_06010_),
    .B(_06011_));
 sg13g2_nand2_1 _14028_ (.Y(_06012_),
    .A(net180),
    .B(\synth.voice.genblk4[0].next_state_scan[9] ));
 sg13g2_o21ai_1 _14029_ (.B1(_06012_),
    .Y(_06013_),
    .A1(net180),
    .A2(_04853_));
 sg13g2_nand2_1 _14030_ (.Y(_06014_),
    .A(net43),
    .B(_06013_));
 sg13g2_o21ai_1 _14031_ (.B1(_06014_),
    .Y(_01289_),
    .A1(_05904_),
    .A2(net44));
 sg13g2_a21oi_1 _14032_ (.A1(_04668_),
    .A2(_04674_),
    .Y(_06015_),
    .B1(_04701_));
 sg13g2_inv_1 _14033_ (.Y(_06016_),
    .A(_06015_));
 sg13g2_xnor2_1 _14034_ (.Y(_06017_),
    .A(_04529_),
    .B(_04528_));
 sg13g2_inv_1 _14035_ (.Y(_06018_),
    .A(_04684_));
 sg13g2_nand2b_1 _14036_ (.Y(_06019_),
    .B(_06018_),
    .A_N(_04665_));
 sg13g2_a22oi_1 _14037_ (.Y(_06020_),
    .B1(_06019_),
    .B2(net34),
    .A2(_06017_),
    .A1(_04667_));
 sg13g2_nand2_1 _14038_ (.Y(_06021_),
    .A(net136),
    .B(\synth.voice.wave_reg[0] ));
 sg13g2_o21ai_1 _14039_ (.B1(_06021_),
    .Y(_01309_),
    .A1(_06016_),
    .A2(_06020_));
 sg13g2_inv_1 _14040_ (.Y(_06022_),
    .A(\synth.voice.wave_reg[1] ));
 sg13g2_inv_1 _14041_ (.Y(_06023_),
    .A(_04665_));
 sg13g2_xnor2_1 _14042_ (.Y(_06024_),
    .A(_06017_),
    .B(net34));
 sg13g2_nor2_1 _14043_ (.A(_06018_),
    .B(_04651_),
    .Y(_06025_));
 sg13g2_nor2_2 _14044_ (.A(_04667_),
    .B(_06025_),
    .Y(_06026_));
 sg13g2_o21ai_1 _14045_ (.B1(_06026_),
    .Y(_06027_),
    .A1(_06023_),
    .A2(_06024_));
 sg13g2_xor2_1 _14046_ (.B(_04625_),
    .A(_04531_),
    .X(_06028_));
 sg13g2_inv_1 _14047_ (.Y(_06029_),
    .A(_06028_));
 sg13g2_a21oi_1 _14048_ (.A1(_06029_),
    .A2(_04667_),
    .Y(_06030_),
    .B1(_06016_));
 sg13g2_nand2_1 _14049_ (.Y(_06031_),
    .A(_06027_),
    .B(_06030_));
 sg13g2_o21ai_1 _14050_ (.B1(_06031_),
    .Y(_01310_),
    .A1(_06022_),
    .A2(_04700_));
 sg13g2_inv_1 _14051_ (.Y(_06032_),
    .A(_04667_));
 sg13g2_xor2_1 _14052_ (.B(_04504_),
    .A(_04533_),
    .X(_06033_));
 sg13g2_nand2_1 _14053_ (.Y(_06034_),
    .A(_04698_),
    .B(_06028_));
 sg13g2_nand2_1 _14054_ (.Y(_06035_),
    .A(_04651_),
    .B(_06029_));
 sg13g2_nand3_1 _14055_ (.B(_06035_),
    .C(_04665_),
    .A(_06034_),
    .Y(_06036_));
 sg13g2_a21oi_1 _14056_ (.A1(_06036_),
    .A2(_06026_),
    .Y(_06037_),
    .B1(_06016_));
 sg13g2_o21ai_1 _14057_ (.B1(_06037_),
    .Y(_06038_),
    .A1(_06032_),
    .A2(_06033_));
 sg13g2_nand2_1 _14058_ (.Y(_06039_),
    .A(net136),
    .B(\synth.voice.wave_reg[2] ));
 sg13g2_nand2_1 _14059_ (.Y(_01311_),
    .A(_06038_),
    .B(_06039_));
 sg13g2_xnor2_1 _14060_ (.Y(_06040_),
    .A(_04523_),
    .B(_04676_));
 sg13g2_nand2b_1 _14061_ (.Y(_06041_),
    .B(_04651_),
    .A_N(_06033_));
 sg13g2_nand2_1 _14062_ (.Y(_06042_),
    .A(_04698_),
    .B(_06033_));
 sg13g2_nand3_1 _14063_ (.B(_06042_),
    .C(_04665_),
    .A(_06041_),
    .Y(_06043_));
 sg13g2_a21oi_1 _14064_ (.A1(_06043_),
    .A2(_06026_),
    .Y(_06044_),
    .B1(_06016_));
 sg13g2_o21ai_1 _14065_ (.B1(_06044_),
    .Y(_06045_),
    .A1(_06032_),
    .A2(_06040_));
 sg13g2_nand2_1 _14066_ (.Y(_06046_),
    .A(net136),
    .B(\synth.voice.wave_reg[3] ));
 sg13g2_nand2_1 _14067_ (.Y(_01312_),
    .A(_06045_),
    .B(_06046_));
 sg13g2_xnor2_1 _14068_ (.Y(_06047_),
    .A(_04569_),
    .B(_04540_));
 sg13g2_inv_1 _14069_ (.Y(_06048_),
    .A(_06047_));
 sg13g2_nand2b_1 _14070_ (.Y(_06049_),
    .B(_04651_),
    .A_N(_06040_));
 sg13g2_nand2_1 _14071_ (.Y(_06050_),
    .A(_04646_),
    .B(_06040_));
 sg13g2_nand3_1 _14072_ (.B(_06050_),
    .C(_04665_),
    .A(_06049_),
    .Y(_06051_));
 sg13g2_a21oi_1 _14073_ (.A1(_06051_),
    .A2(_06026_),
    .Y(_06052_),
    .B1(_06016_));
 sg13g2_o21ai_1 _14074_ (.B1(_06052_),
    .Y(_06053_),
    .A1(_06032_),
    .A2(_06048_));
 sg13g2_nand2_1 _14075_ (.Y(_06054_),
    .A(net136),
    .B(\synth.voice.wave_reg[4] ));
 sg13g2_nand2_1 _14076_ (.Y(_01313_),
    .A(_06053_),
    .B(_06054_));
 sg13g2_a21oi_1 _14077_ (.A1(_04531_),
    .A2(_04628_),
    .Y(_06055_),
    .B1(_04612_));
 sg13g2_xnor2_1 _14078_ (.Y(_06056_),
    .A(_04554_),
    .B(_06055_));
 sg13g2_nand2_1 _14079_ (.Y(_06057_),
    .A(_04651_),
    .B(_06047_));
 sg13g2_nand2_1 _14080_ (.Y(_06058_),
    .A(_04646_),
    .B(_06048_));
 sg13g2_nand3_1 _14081_ (.B(_06058_),
    .C(_04665_),
    .A(_06057_),
    .Y(_06059_));
 sg13g2_a21oi_1 _14082_ (.A1(_06059_),
    .A2(_06026_),
    .Y(_06060_),
    .B1(_06016_));
 sg13g2_o21ai_1 _14083_ (.B1(_06060_),
    .Y(_06061_),
    .A1(_06032_),
    .A2(_06056_));
 sg13g2_nand2_1 _14084_ (.Y(_06062_),
    .A(net136),
    .B(\synth.voice.wave_reg[5] ));
 sg13g2_nand2_1 _14085_ (.Y(_01314_),
    .A(_06061_),
    .B(_06062_));
 sg13g2_a21oi_1 _14086_ (.A1(net34),
    .A2(_06056_),
    .Y(_06063_),
    .B1(_06023_));
 sg13g2_o21ai_1 _14087_ (.B1(_06063_),
    .Y(_06064_),
    .A1(net34),
    .A2(_06056_));
 sg13g2_nand2_1 _14088_ (.Y(_06065_),
    .A(_04658_),
    .B(_04674_));
 sg13g2_nand3_1 _14089_ (.B(_06026_),
    .C(_06065_),
    .A(_06064_),
    .Y(_06066_));
 sg13g2_o21ai_1 _14090_ (.B1(_04597_),
    .Y(_06067_),
    .A1(_04570_),
    .A2(_04539_));
 sg13g2_nand4_1 _14091_ (.B(_04534_),
    .C(_04554_),
    .A(_04524_),
    .Y(_06068_),
    .D(_04569_));
 sg13g2_nand2b_1 _14092_ (.Y(_06069_),
    .B(_06068_),
    .A_N(_06067_));
 sg13g2_xnor2_1 _14093_ (.Y(_06070_),
    .A(_04590_),
    .B(_06069_));
 sg13g2_a21oi_1 _14094_ (.A1(_06070_),
    .A2(_04667_),
    .Y(_06071_),
    .B1(_06016_));
 sg13g2_nand2_1 _14095_ (.Y(_06072_),
    .A(_06066_),
    .B(_06071_));
 sg13g2_nand2_1 _14096_ (.Y(_06073_),
    .A(net136),
    .B(\synth.voice.wave_reg[6] ));
 sg13g2_nand2_1 _14097_ (.Y(_01315_),
    .A(_06072_),
    .B(_06073_));
 sg13g2_inv_1 _14098_ (.Y(_06074_),
    .A(\synth.voice.wave_reg[7] ));
 sg13g2_nand2_1 _14099_ (.Y(_06075_),
    .A(_04681_),
    .B(_04667_));
 sg13g2_nand3_1 _14100_ (.B(_04691_),
    .C(_06015_),
    .A(_06075_),
    .Y(_06076_));
 sg13g2_nor2_1 _14101_ (.A(_06070_),
    .B(_04651_),
    .Y(_06077_));
 sg13g2_nor2b_1 _14102_ (.A(net34),
    .B_N(_06070_),
    .Y(_06078_));
 sg13g2_nor3_1 _14103_ (.A(_06023_),
    .B(_06077_),
    .C(_06078_),
    .Y(_06079_));
 sg13g2_nor3_1 _14104_ (.A(_06025_),
    .B(_06076_),
    .C(_06079_),
    .Y(_06080_));
 sg13g2_a21oi_1 _14105_ (.A1(_06074_),
    .A2(_04702_),
    .Y(_01316_),
    .B1(_06080_));
 sg13g2_inv_1 _14106_ (.Y(_06081_),
    .A(_04606_));
 sg13g2_o21ai_1 _14107_ (.B1(_04700_),
    .Y(_06082_),
    .A1(_06032_),
    .A2(_06081_));
 sg13g2_nand2_1 _14108_ (.Y(_06083_),
    .A(_04681_),
    .B(_04665_));
 sg13g2_a21oi_1 _14109_ (.A1(_06083_),
    .A2(_06019_),
    .Y(_06084_),
    .B1(net34));
 sg13g2_a21oi_1 _14110_ (.A1(net34),
    .A2(_06083_),
    .Y(_06085_),
    .B1(_06084_));
 sg13g2_nand2_1 _14111_ (.Y(_06086_),
    .A(_04702_),
    .B(\synth.voice.wave_reg[8] ));
 sg13g2_o21ai_1 _14112_ (.B1(_06086_),
    .Y(_01317_),
    .A1(_06082_),
    .A2(_06085_));
 sg13g2_inv_1 _14113_ (.Y(_06087_),
    .A(\synth.voice.wave_reg[9] ));
 sg13g2_nand2_1 _14114_ (.Y(_06088_),
    .A(_04694_),
    .B(_04703_));
 sg13g2_o21ai_1 _14115_ (.B1(_06088_),
    .Y(_01318_),
    .A1(_06087_),
    .A2(_04700_));
 sg13g2_inv_1 _14116_ (.Y(_06089_),
    .A(_02272_));
 sg13g2_nor2_1 _14117_ (.A(net1),
    .B(net2),
    .Y(_06090_));
 sg13g2_a21oi_1 _14118_ (.A1(net1),
    .A2(_06089_),
    .Y(_00183_),
    .B1(_06090_));
 sg13g2_nor2_1 _14119_ (.A(\ppu.copper_inst.store[5] ),
    .B(\ppu.copper_inst.store[4] ),
    .Y(_06091_));
 sg13g2_nand3_1 _14120_ (.B(_02376_),
    .C(_06091_),
    .A(_02374_),
    .Y(_06092_));
 sg13g2_nor2_1 _14121_ (.A(_03085_),
    .B(_06092_),
    .Y(_06093_));
 sg13g2_nand2_1 _14122_ (.Y(_06094_),
    .A(_06093_),
    .B(_02384_));
 sg13g2_nand4_1 _14123_ (.B(_01854_),
    .C(_02376_),
    .A(_02374_),
    .Y(_06095_),
    .D(_06091_));
 sg13g2_buf_2 _14124_ (.A(_06095_),
    .X(_06096_));
 sg13g2_nand2_1 _14125_ (.Y(_06097_),
    .A(_02928_),
    .B(\ppu.depth_out_t[1] ));
 sg13g2_inv_1 _14126_ (.Y(_06098_),
    .A(\ppu.depth_out_t[0] ));
 sg13g2_nand3_1 _14127_ (.B(\ppu.depth_out_s[0] ),
    .C(_06098_),
    .A(_06097_),
    .Y(_06099_));
 sg13g2_inv_1 _14128_ (.Y(_06100_),
    .A(\ppu.depth_out_t[1] ));
 sg13g2_inv_1 _14129_ (.Y(_06101_),
    .A(\ppu.display_mask[2] ));
 sg13g2_a21oi_1 _14130_ (.A1(_06100_),
    .A2(\ppu.depth_out_s[1] ),
    .Y(_06102_),
    .B1(_06101_));
 sg13g2_nand2_1 _14131_ (.Y(_06103_),
    .A(_06099_),
    .B(_06102_));
 sg13g2_buf_2 _14132_ (.A(_06103_),
    .X(_06104_));
 sg13g2_inv_1 _14133_ (.Y(_06105_),
    .A(_02288_));
 sg13g2_inv_1 _14134_ (.Y(_06106_),
    .A(\ppu.pixel_out_t[0] ));
 sg13g2_a22oi_1 _14135_ (.Y(_06107_),
    .B1(_06106_),
    .B2(_06104_),
    .A2(net389),
    .A1(_06105_));
 sg13g2_o21ai_1 _14136_ (.B1(_06107_),
    .Y(_06108_),
    .A1(\ppu.pixel_out_s[0] ),
    .A2(_06104_));
 sg13g2_nand2_1 _14137_ (.Y(_06109_),
    .A(_06096_),
    .B(_06108_));
 sg13g2_nand3_1 _14138_ (.B(_06109_),
    .C(net343),
    .A(_06094_),
    .Y(_06110_));
 sg13g2_nand2_1 _14139_ (.Y(_06111_),
    .A(net390),
    .B(\ppu.curr_pal_addr[0] ));
 sg13g2_nand2_1 _14140_ (.Y(_06112_),
    .A(_06110_),
    .B(_06111_));
 sg13g2_buf_1 _14141_ (.A(_06112_),
    .X(_00262_));
 sg13g2_nand2_1 _14142_ (.Y(_06113_),
    .A(_06093_),
    .B(_02382_));
 sg13g2_inv_1 _14143_ (.Y(_06114_),
    .A(\ppu.pixel_out_t[1] ));
 sg13g2_a22oi_1 _14144_ (.Y(_06115_),
    .B1(_06114_),
    .B2(_06104_),
    .A2(net389),
    .A1(_06105_));
 sg13g2_o21ai_1 _14145_ (.B1(_06115_),
    .Y(_06116_),
    .A1(\ppu.pixel_out_s[1] ),
    .A2(_06104_));
 sg13g2_nand2_1 _14146_ (.Y(_06117_),
    .A(_06096_),
    .B(_06116_));
 sg13g2_nand3_1 _14147_ (.B(_06117_),
    .C(net343),
    .A(_06113_),
    .Y(_06118_));
 sg13g2_nand2_1 _14148_ (.Y(_06119_),
    .A(net390),
    .B(\ppu.curr_pal_addr[1] ));
 sg13g2_nand2_1 _14149_ (.Y(_06120_),
    .A(_06118_),
    .B(_06119_));
 sg13g2_buf_1 _14150_ (.A(_06120_),
    .X(_00263_));
 sg13g2_nand2_1 _14151_ (.Y(_06121_),
    .A(_06093_),
    .B(_02460_));
 sg13g2_inv_1 _14152_ (.Y(_06122_),
    .A(\ppu.pixel_out_t[2] ));
 sg13g2_a22oi_1 _14153_ (.Y(_06123_),
    .B1(_06122_),
    .B2(_06104_),
    .A2(net389),
    .A1(_06105_));
 sg13g2_o21ai_1 _14154_ (.B1(_06123_),
    .Y(_06124_),
    .A1(\ppu.pixel_out_s[2] ),
    .A2(_06104_));
 sg13g2_nand2_1 _14155_ (.Y(_06125_),
    .A(_06096_),
    .B(_06124_));
 sg13g2_nand3_1 _14156_ (.B(_06125_),
    .C(net343),
    .A(_06121_),
    .Y(_06126_));
 sg13g2_nand2_1 _14157_ (.Y(_06127_),
    .A(net390),
    .B(\ppu.curr_pal_addr[2] ));
 sg13g2_nand2_1 _14158_ (.Y(_06128_),
    .A(_06126_),
    .B(_06127_));
 sg13g2_buf_1 _14159_ (.A(_06128_),
    .X(_00264_));
 sg13g2_nand2_1 _14160_ (.Y(_06129_),
    .A(_06093_),
    .B(_02294_));
 sg13g2_nand2_1 _14161_ (.Y(_06130_),
    .A(_06104_),
    .B(_00042_));
 sg13g2_nand3_1 _14162_ (.B(_00041_),
    .C(_06102_),
    .A(_06099_),
    .Y(_06131_));
 sg13g2_nand2_1 _14163_ (.Y(_06132_),
    .A(_06105_),
    .B(_02285_));
 sg13g2_nand3_1 _14164_ (.B(_06131_),
    .C(_06132_),
    .A(_06130_),
    .Y(_06133_));
 sg13g2_nand2_1 _14165_ (.Y(_06134_),
    .A(_06096_),
    .B(_06133_));
 sg13g2_nand3_1 _14166_ (.B(_06134_),
    .C(net343),
    .A(_06129_),
    .Y(_06135_));
 sg13g2_nand2_1 _14167_ (.Y(_06136_),
    .A(net390),
    .B(\ppu.curr_pal_addr[3] ));
 sg13g2_nand2_1 _14168_ (.Y(_06137_),
    .A(_06135_),
    .B(_06136_));
 sg13g2_buf_1 _14169_ (.A(_06137_),
    .X(_00265_));
 sg13g2_nor2_1 _14170_ (.A(_00264_),
    .B(_00265_),
    .Y(_06138_));
 sg13g2_buf_1 _14171_ (.A(_06138_),
    .X(_06139_));
 sg13g2_nor2_1 _14172_ (.A(_00262_),
    .B(_00263_),
    .Y(_06140_));
 sg13g2_buf_2 _14173_ (.A(_06140_),
    .X(_06141_));
 sg13g2_nand2_1 _14174_ (.Y(_06142_),
    .A(_06139_),
    .B(_06141_));
 sg13g2_buf_2 _14175_ (.A(_06142_),
    .X(_06143_));
 sg13g2_mux2_1 _14176_ (.A0(\ppu.pal[0][4] ),
    .A1(\ppu.pal[0][0] ),
    .S(net70),
    .X(_00299_));
 sg13g2_mux2_1 _14177_ (.A0(\ppu.pal[0][5] ),
    .A1(\ppu.pal[0][1] ),
    .S(net70),
    .X(_00300_));
 sg13g2_mux2_1 _14178_ (.A0(\ppu.pal[0][6] ),
    .A1(\ppu.pal[0][2] ),
    .S(_06143_),
    .X(_00301_));
 sg13g2_mux2_1 _14179_ (.A0(\ppu.pal[0][7] ),
    .A1(\ppu.pal[0][3] ),
    .S(net70),
    .X(_00302_));
 sg13g2_a21oi_1 _14180_ (.A1(_06096_),
    .A2(_06133_),
    .Y(_06144_),
    .B1(net390));
 sg13g2_inv_1 _14181_ (.Y(_06145_),
    .A(_06136_));
 sg13g2_a21oi_2 _14182_ (.B1(_06145_),
    .Y(_06146_),
    .A2(_06129_),
    .A1(_06144_));
 sg13g2_nand2_1 _14183_ (.Y(_06147_),
    .A(_06146_),
    .B(_00264_));
 sg13g2_a21oi_1 _14184_ (.A1(_06096_),
    .A2(_06116_),
    .Y(_06148_),
    .B1(_02063_));
 sg13g2_inv_1 _14185_ (.Y(_06149_),
    .A(_06119_));
 sg13g2_a21oi_2 _14186_ (.B1(_06149_),
    .Y(_06150_),
    .A2(_06113_),
    .A1(_06148_));
 sg13g2_nand2_1 _14187_ (.Y(_06151_),
    .A(_06150_),
    .B(_00262_));
 sg13g2_nor2_1 _14188_ (.A(_06147_),
    .B(_06151_),
    .Y(_06152_));
 sg13g2_nand2_1 _14189_ (.Y(_06153_),
    .A(_06152_),
    .B(\ppu.pal[5][0] ));
 sg13g2_buf_1 _14190_ (.A(_06141_),
    .X(_06154_));
 sg13g2_a21oi_1 _14191_ (.A1(_06096_),
    .A2(_06124_),
    .Y(_06155_),
    .B1(net390));
 sg13g2_inv_1 _14192_ (.Y(_06156_),
    .A(_06127_));
 sg13g2_a21oi_2 _14193_ (.B1(_06156_),
    .Y(_06157_),
    .A2(_06121_),
    .A1(_06155_));
 sg13g2_nor2_1 _14194_ (.A(_00265_),
    .B(_06157_),
    .Y(_06158_));
 sg13g2_buf_2 _14195_ (.A(_06158_),
    .X(_06159_));
 sg13g2_nand3_1 _14196_ (.B(_06159_),
    .C(\ppu.pal[4][0] ),
    .A(net85),
    .Y(_06160_));
 sg13g2_nand2_1 _14197_ (.Y(_06161_),
    .A(_06153_),
    .B(_06160_));
 sg13g2_a21oi_1 _14198_ (.A1(_06096_),
    .A2(_06108_),
    .Y(_06162_),
    .B1(net390));
 sg13g2_inv_1 _14199_ (.Y(_06163_),
    .A(_06111_));
 sg13g2_a21oi_2 _14200_ (.B1(_06163_),
    .Y(_06164_),
    .A2(_06094_),
    .A1(_06162_));
 sg13g2_nand2_1 _14201_ (.Y(_06165_),
    .A(_06164_),
    .B(_00263_));
 sg13g2_nor2_1 _14202_ (.A(_06147_),
    .B(_06165_),
    .Y(_06166_));
 sg13g2_buf_1 _14203_ (.A(_06166_),
    .X(_06167_));
 sg13g2_nand2_1 _14204_ (.Y(_06168_),
    .A(net84),
    .B(\ppu.pal[6][0] ));
 sg13g2_nand2_1 _14205_ (.Y(_06169_),
    .A(_00262_),
    .B(_00263_));
 sg13g2_nor2_1 _14206_ (.A(_06147_),
    .B(_06169_),
    .Y(_06170_));
 sg13g2_buf_1 _14207_ (.A(_06170_),
    .X(_06171_));
 sg13g2_nand2_1 _14208_ (.Y(_06172_),
    .A(net83),
    .B(\ppu.pal[7][0] ));
 sg13g2_nand2_1 _14209_ (.Y(_06173_),
    .A(_06168_),
    .B(_06172_));
 sg13g2_nor2_1 _14210_ (.A(_06161_),
    .B(_06173_),
    .Y(_06174_));
 sg13g2_nor2_1 _14211_ (.A(_06164_),
    .B(_06150_),
    .Y(_06175_));
 sg13g2_buf_2 _14212_ (.A(_06175_),
    .X(_06176_));
 sg13g2_nand2_1 _14213_ (.Y(_06177_),
    .A(_06176_),
    .B(_06138_));
 sg13g2_buf_1 _14214_ (.A(_06177_),
    .X(_06178_));
 sg13g2_nor2b_1 _14215_ (.A(_06178_),
    .B_N(\ppu.pal[3][0] ),
    .Y(_06179_));
 sg13g2_nor2_2 _14216_ (.A(_00262_),
    .B(_06150_),
    .Y(_06180_));
 sg13g2_nand3_1 _14217_ (.B(_06180_),
    .C(\ppu.pal[2][0] ),
    .A(net90),
    .Y(_06181_));
 sg13g2_nor2_2 _14218_ (.A(_00263_),
    .B(_06164_),
    .Y(_06182_));
 sg13g2_nand3_1 _14219_ (.B(_06182_),
    .C(\ppu.pal[1][0] ),
    .A(net90),
    .Y(_06183_));
 sg13g2_nand2_1 _14220_ (.Y(_06184_),
    .A(_06181_),
    .B(_06183_));
 sg13g2_nor2_1 _14221_ (.A(_06179_),
    .B(_06184_),
    .Y(_06185_));
 sg13g2_nand2_1 _14222_ (.Y(_06186_),
    .A(_06174_),
    .B(_06185_));
 sg13g2_nand2_1 _14223_ (.Y(_06187_),
    .A(_06157_),
    .B(_00265_));
 sg13g2_nor2_1 _14224_ (.A(_06151_),
    .B(_06187_),
    .Y(_06188_));
 sg13g2_nand2_1 _14225_ (.Y(_06189_),
    .A(_06188_),
    .B(\ppu.pal[9][0] ));
 sg13g2_nor2_2 _14226_ (.A(_00264_),
    .B(_06146_),
    .Y(_06190_));
 sg13g2_nand3_1 _14227_ (.B(_06190_),
    .C(\ppu.pal[8][0] ),
    .A(net85),
    .Y(_06191_));
 sg13g2_nand2_1 _14228_ (.Y(_06192_),
    .A(_06189_),
    .B(_06191_));
 sg13g2_nor2_1 _14229_ (.A(_06169_),
    .B(_06187_),
    .Y(_06193_));
 sg13g2_buf_1 _14230_ (.A(_06193_),
    .X(_06194_));
 sg13g2_nand2_1 _14231_ (.Y(_06195_),
    .A(net81),
    .B(\ppu.pal[11][0] ));
 sg13g2_nor2_2 _14232_ (.A(_06165_),
    .B(_06187_),
    .Y(_06196_));
 sg13g2_buf_8 _14233_ (.A(_06196_),
    .X(_06197_));
 sg13g2_nand2_1 _14234_ (.Y(_06198_),
    .A(net80),
    .B(\ppu.pal[10][0] ));
 sg13g2_nand2_1 _14235_ (.Y(_06199_),
    .A(_06195_),
    .B(_06198_));
 sg13g2_nor2_1 _14236_ (.A(_06192_),
    .B(_06199_),
    .Y(_06200_));
 sg13g2_nand2_1 _14237_ (.Y(_06201_),
    .A(_00264_),
    .B(_00265_));
 sg13g2_nor2_1 _14238_ (.A(_06151_),
    .B(_06201_),
    .Y(_06202_));
 sg13g2_nand2_1 _14239_ (.Y(_06203_),
    .A(_06202_),
    .B(\ppu.pal[13][0] ));
 sg13g2_nor2_2 _14240_ (.A(_06157_),
    .B(_06146_),
    .Y(_06204_));
 sg13g2_nand3_1 _14241_ (.B(_06141_),
    .C(\ppu.pal[12][0] ),
    .A(_06204_),
    .Y(_06205_));
 sg13g2_nand2_1 _14242_ (.Y(_06206_),
    .A(_06203_),
    .B(_06205_));
 sg13g2_nor2_2 _14243_ (.A(_06169_),
    .B(_06201_),
    .Y(_06207_));
 sg13g2_nand2_1 _14244_ (.Y(_06208_),
    .A(_06207_),
    .B(\ppu.pal[15][0] ));
 sg13g2_nor2_1 _14245_ (.A(_06165_),
    .B(_06201_),
    .Y(_06209_));
 sg13g2_nand2_1 _14246_ (.Y(_06210_),
    .A(_06209_),
    .B(\ppu.pal[14][0] ));
 sg13g2_nand2_1 _14247_ (.Y(_06211_),
    .A(_06208_),
    .B(_06210_));
 sg13g2_nor2_1 _14248_ (.A(_06206_),
    .B(_06211_),
    .Y(_06212_));
 sg13g2_nand2_1 _14249_ (.Y(_06213_),
    .A(_06200_),
    .B(_06212_));
 sg13g2_nor2_1 _14250_ (.A(_06186_),
    .B(_06213_),
    .Y(_06214_));
 sg13g2_nor2_2 _14251_ (.A(_00122_),
    .B(_06092_),
    .Y(_06215_));
 sg13g2_inv_1 _14252_ (.Y(_06216_),
    .A(_06215_));
 sg13g2_inv_4 _14253_ (.A(net70),
    .Y(_06217_));
 sg13g2_nand2_1 _14254_ (.Y(_06218_),
    .A(_06217_),
    .B(\ppu.pal[0][0] ));
 sg13g2_nand3_1 _14255_ (.B(_06216_),
    .C(_06218_),
    .A(_06214_),
    .Y(_06219_));
 sg13g2_buf_2 _14256_ (.A(_06219_),
    .X(_06220_));
 sg13g2_buf_1 _14257_ (.A(_06220_),
    .X(_06221_));
 sg13g2_buf_1 _14258_ (.A(net390),
    .X(_06222_));
 sg13g2_nor2_1 _14259_ (.A(net320),
    .B(_02393_),
    .Y(_06223_));
 sg13g2_a21oi_1 _14260_ (.A1(net320),
    .A2(_02408_),
    .Y(_06224_),
    .B1(_06223_));
 sg13g2_nand2_1 _14261_ (.Y(_06225_),
    .A(_06215_),
    .B(_06224_));
 sg13g2_buf_2 _14262_ (.A(_06225_),
    .X(_06226_));
 sg13g2_buf_1 _14263_ (.A(_06226_),
    .X(_06227_));
 sg13g2_nand3_1 _14264_ (.B(_06217_),
    .C(net115),
    .A(net41),
    .Y(_06228_));
 sg13g2_nand2_1 _14265_ (.Y(_06229_),
    .A(net70),
    .B(\ppu.pal[0][4] ));
 sg13g2_nand2_1 _14266_ (.Y(_00303_),
    .A(_06228_),
    .B(_06229_));
 sg13g2_nand3_1 _14267_ (.B(_06159_),
    .C(\ppu.pal[4][1] ),
    .A(net85),
    .Y(_06230_));
 sg13g2_nand3_1 _14268_ (.B(_06182_),
    .C(\ppu.pal[5][1] ),
    .A(_06159_),
    .Y(_06231_));
 sg13g2_nand2_1 _14269_ (.Y(_06232_),
    .A(_06230_),
    .B(_06231_));
 sg13g2_nand2_1 _14270_ (.Y(_06233_),
    .A(_06166_),
    .B(\ppu.pal[6][1] ));
 sg13g2_nand2_1 _14271_ (.Y(_06234_),
    .A(_06170_),
    .B(\ppu.pal[7][1] ));
 sg13g2_nand2_1 _14272_ (.Y(_06235_),
    .A(_06233_),
    .B(_06234_));
 sg13g2_nor2_1 _14273_ (.A(_06232_),
    .B(_06235_),
    .Y(_06236_));
 sg13g2_nor2b_1 _14274_ (.A(_06177_),
    .B_N(\ppu.pal[3][1] ),
    .Y(_06237_));
 sg13g2_nand3_1 _14275_ (.B(_06180_),
    .C(\ppu.pal[2][1] ),
    .A(net90),
    .Y(_06238_));
 sg13g2_nand3_1 _14276_ (.B(_06182_),
    .C(\ppu.pal[1][1] ),
    .A(_06139_),
    .Y(_06239_));
 sg13g2_nand2_1 _14277_ (.Y(_06240_),
    .A(_06238_),
    .B(_06239_));
 sg13g2_nor2_1 _14278_ (.A(_06237_),
    .B(_06240_),
    .Y(_06241_));
 sg13g2_nand2_1 _14279_ (.Y(_06242_),
    .A(_06236_),
    .B(_06241_));
 sg13g2_nand2_1 _14280_ (.Y(_06243_),
    .A(_06209_),
    .B(\ppu.pal[14][1] ));
 sg13g2_nand3_1 _14281_ (.B(_06141_),
    .C(\ppu.pal[12][1] ),
    .A(_06204_),
    .Y(_06244_));
 sg13g2_nand2_1 _14282_ (.Y(_06245_),
    .A(_06243_),
    .B(_06244_));
 sg13g2_buf_1 _14283_ (.A(_06202_),
    .X(_06246_));
 sg13g2_nand2_1 _14284_ (.Y(_06247_),
    .A(net79),
    .B(\ppu.pal[13][1] ));
 sg13g2_nand2_1 _14285_ (.Y(_06248_),
    .A(_06207_),
    .B(\ppu.pal[15][1] ));
 sg13g2_nand2_1 _14286_ (.Y(_06249_),
    .A(_06247_),
    .B(_06248_));
 sg13g2_nor2_1 _14287_ (.A(_06245_),
    .B(_06249_),
    .Y(_06250_));
 sg13g2_nand2_1 _14288_ (.Y(_06251_),
    .A(_06196_),
    .B(\ppu.pal[10][1] ));
 sg13g2_nand3_1 _14289_ (.B(_06190_),
    .C(\ppu.pal[11][1] ),
    .A(_06176_),
    .Y(_06252_));
 sg13g2_nand2_1 _14290_ (.Y(_06253_),
    .A(_06251_),
    .B(_06252_));
 sg13g2_nand2_1 _14291_ (.Y(_06254_),
    .A(_06188_),
    .B(\ppu.pal[9][1] ));
 sg13g2_nand3_1 _14292_ (.B(_06190_),
    .C(\ppu.pal[8][1] ),
    .A(net85),
    .Y(_06255_));
 sg13g2_nand2_1 _14293_ (.Y(_06256_),
    .A(_06254_),
    .B(_06255_));
 sg13g2_nor2_1 _14294_ (.A(_06253_),
    .B(_06256_),
    .Y(_06257_));
 sg13g2_nand2_1 _14295_ (.Y(_06258_),
    .A(_06250_),
    .B(_06257_));
 sg13g2_nor2_1 _14296_ (.A(_06242_),
    .B(_06258_),
    .Y(_06259_));
 sg13g2_nand2_1 _14297_ (.Y(_06260_),
    .A(_06217_),
    .B(\ppu.pal[0][1] ));
 sg13g2_nand3_1 _14298_ (.B(_06216_),
    .C(_06260_),
    .A(_06259_),
    .Y(_06261_));
 sg13g2_buf_2 _14299_ (.A(_06261_),
    .X(_06262_));
 sg13g2_buf_8 _14300_ (.A(_06262_),
    .X(_06263_));
 sg13g2_nor2_1 _14301_ (.A(net320),
    .B(_02397_),
    .Y(_06264_));
 sg13g2_a21oi_1 _14302_ (.A1(net320),
    .A2(net406),
    .Y(_06265_),
    .B1(_06264_));
 sg13g2_nand2_1 _14303_ (.Y(_06266_),
    .A(_06215_),
    .B(_06265_));
 sg13g2_buf_2 _14304_ (.A(_06266_),
    .X(_06267_));
 sg13g2_buf_1 _14305_ (.A(_06267_),
    .X(_06268_));
 sg13g2_nand3_1 _14306_ (.B(_06217_),
    .C(net114),
    .A(net40),
    .Y(_06269_));
 sg13g2_nand2_1 _14307_ (.Y(_06270_),
    .A(net70),
    .B(\ppu.pal[0][5] ));
 sg13g2_nand2_1 _14308_ (.Y(_00304_),
    .A(_06269_),
    .B(_06270_));
 sg13g2_nand2_1 _14309_ (.Y(_06271_),
    .A(_06166_),
    .B(\ppu.pal[6][2] ));
 sg13g2_nand3_1 _14310_ (.B(_06159_),
    .C(\ppu.pal[7][2] ),
    .A(_06176_),
    .Y(_06272_));
 sg13g2_nand2_1 _14311_ (.Y(_06273_),
    .A(_06271_),
    .B(_06272_));
 sg13g2_buf_1 _14312_ (.A(_06152_),
    .X(_06274_));
 sg13g2_nand2_1 _14313_ (.Y(_06275_),
    .A(net78),
    .B(\ppu.pal[5][2] ));
 sg13g2_nand3_1 _14314_ (.B(_06159_),
    .C(\ppu.pal[4][2] ),
    .A(net85),
    .Y(_06276_));
 sg13g2_nand2_1 _14315_ (.Y(_06277_),
    .A(_06275_),
    .B(_06276_));
 sg13g2_nor2_1 _14316_ (.A(_06273_),
    .B(_06277_),
    .Y(_06278_));
 sg13g2_nand2_1 _14317_ (.Y(_06279_),
    .A(_06138_),
    .B(_06182_));
 sg13g2_buf_1 _14318_ (.A(_06279_),
    .X(_06280_));
 sg13g2_nor2b_1 _14319_ (.A(_06280_),
    .B_N(\ppu.pal[1][2] ),
    .Y(_06281_));
 sg13g2_nand3_1 _14320_ (.B(_06180_),
    .C(\ppu.pal[2][2] ),
    .A(net90),
    .Y(_06282_));
 sg13g2_nand3_1 _14321_ (.B(net90),
    .C(\ppu.pal[3][2] ),
    .A(_06176_),
    .Y(_06283_));
 sg13g2_nand2_1 _14322_ (.Y(_06284_),
    .A(_06282_),
    .B(_06283_));
 sg13g2_nor2_1 _14323_ (.A(_06281_),
    .B(_06284_),
    .Y(_06285_));
 sg13g2_nand2_1 _14324_ (.Y(_06286_),
    .A(_06278_),
    .B(_06285_));
 sg13g2_nand2_1 _14325_ (.Y(_06287_),
    .A(_06202_),
    .B(\ppu.pal[13][2] ));
 sg13g2_nand3_1 _14326_ (.B(_06141_),
    .C(\ppu.pal[12][2] ),
    .A(_06204_),
    .Y(_06288_));
 sg13g2_nand2_1 _14327_ (.Y(_06289_),
    .A(_06287_),
    .B(_06288_));
 sg13g2_buf_8 _14328_ (.A(_06207_),
    .X(_06290_));
 sg13g2_nand2_1 _14329_ (.Y(_06291_),
    .A(net76),
    .B(\ppu.pal[15][2] ));
 sg13g2_buf_1 _14330_ (.A(_06209_),
    .X(_06292_));
 sg13g2_nand2_1 _14331_ (.Y(_06293_),
    .A(net75),
    .B(\ppu.pal[14][2] ));
 sg13g2_nand2_1 _14332_ (.Y(_06294_),
    .A(_06291_),
    .B(_06293_));
 sg13g2_nor2_1 _14333_ (.A(_06289_),
    .B(_06294_),
    .Y(_06295_));
 sg13g2_nand2_1 _14334_ (.Y(_06296_),
    .A(_06188_),
    .B(\ppu.pal[9][2] ));
 sg13g2_nand3_1 _14335_ (.B(_06190_),
    .C(\ppu.pal[8][2] ),
    .A(_06141_),
    .Y(_06297_));
 sg13g2_nand2_1 _14336_ (.Y(_06298_),
    .A(_06296_),
    .B(_06297_));
 sg13g2_nand2_1 _14337_ (.Y(_06299_),
    .A(_06193_),
    .B(\ppu.pal[11][2] ));
 sg13g2_nand2_1 _14338_ (.Y(_06300_),
    .A(_06196_),
    .B(\ppu.pal[10][2] ));
 sg13g2_nand2_1 _14339_ (.Y(_06301_),
    .A(_06299_),
    .B(_06300_));
 sg13g2_nor2_1 _14340_ (.A(_06298_),
    .B(_06301_),
    .Y(_06302_));
 sg13g2_nand2_1 _14341_ (.Y(_06303_),
    .A(_06295_),
    .B(_06302_));
 sg13g2_nor2_1 _14342_ (.A(_06286_),
    .B(_06303_),
    .Y(_06304_));
 sg13g2_nand2_1 _14343_ (.Y(_06305_),
    .A(_06217_),
    .B(\ppu.pal[0][2] ));
 sg13g2_nand3_1 _14344_ (.B(_06216_),
    .C(_06305_),
    .A(_06304_),
    .Y(_06306_));
 sg13g2_buf_2 _14345_ (.A(_06306_),
    .X(_06307_));
 sg13g2_buf_8 _14346_ (.A(_06307_),
    .X(_06308_));
 sg13g2_nor2_1 _14347_ (.A(net320),
    .B(_02401_),
    .Y(_06309_));
 sg13g2_a21oi_1 _14348_ (.A1(net320),
    .A2(_02414_),
    .Y(_06310_),
    .B1(_06309_));
 sg13g2_nand2_1 _14349_ (.Y(_06311_),
    .A(_06215_),
    .B(_06310_));
 sg13g2_buf_2 _14350_ (.A(_06311_),
    .X(_06312_));
 sg13g2_buf_1 _14351_ (.A(_06312_),
    .X(_06313_));
 sg13g2_nand3_1 _14352_ (.B(_06217_),
    .C(net113),
    .A(net39),
    .Y(_06314_));
 sg13g2_nand2_1 _14353_ (.Y(_06315_),
    .A(net70),
    .B(\ppu.pal[0][6] ));
 sg13g2_nand2_1 _14354_ (.Y(_00305_),
    .A(_06314_),
    .B(_06315_));
 sg13g2_nand2_1 _14355_ (.Y(_06316_),
    .A(_06166_),
    .B(\ppu.pal[6][3] ));
 sg13g2_nand3_1 _14356_ (.B(_06159_),
    .C(\ppu.pal[7][3] ),
    .A(_06176_),
    .Y(_06317_));
 sg13g2_nand2_1 _14357_ (.Y(_06318_),
    .A(_06316_),
    .B(_06317_));
 sg13g2_nand2_1 _14358_ (.Y(_06319_),
    .A(_06152_),
    .B(\ppu.pal[5][3] ));
 sg13g2_nand3_1 _14359_ (.B(_06159_),
    .C(\ppu.pal[4][3] ),
    .A(net85),
    .Y(_06320_));
 sg13g2_nand2_1 _14360_ (.Y(_06321_),
    .A(_06319_),
    .B(_06320_));
 sg13g2_nor2_1 _14361_ (.A(_06318_),
    .B(_06321_),
    .Y(_06322_));
 sg13g2_nor2b_1 _14362_ (.A(_06279_),
    .B_N(\ppu.pal[1][3] ),
    .Y(_06323_));
 sg13g2_nand3_1 _14363_ (.B(net90),
    .C(\ppu.pal[3][3] ),
    .A(_06176_),
    .Y(_06324_));
 sg13g2_nand3_1 _14364_ (.B(_06180_),
    .C(\ppu.pal[2][3] ),
    .A(net90),
    .Y(_06325_));
 sg13g2_nand2_1 _14365_ (.Y(_06326_),
    .A(_06324_),
    .B(_06325_));
 sg13g2_nor2_1 _14366_ (.A(_06323_),
    .B(_06326_),
    .Y(_06327_));
 sg13g2_nand2_1 _14367_ (.Y(_06328_),
    .A(_06322_),
    .B(_06327_));
 sg13g2_nand2_1 _14368_ (.Y(_06329_),
    .A(_06193_),
    .B(\ppu.pal[11][3] ));
 sg13g2_nand3_1 _14369_ (.B(_06190_),
    .C(\ppu.pal[8][3] ),
    .A(_06154_),
    .Y(_06330_));
 sg13g2_nand2_1 _14370_ (.Y(_06331_),
    .A(_06329_),
    .B(_06330_));
 sg13g2_buf_1 _14371_ (.A(_06188_),
    .X(_06332_));
 sg13g2_nand2_1 _14372_ (.Y(_06333_),
    .A(_06332_),
    .B(\ppu.pal[9][3] ));
 sg13g2_nand2_1 _14373_ (.Y(_06334_),
    .A(_06196_),
    .B(\ppu.pal[10][3] ));
 sg13g2_nand2_1 _14374_ (.Y(_06335_),
    .A(_06333_),
    .B(_06334_));
 sg13g2_nor2_1 _14375_ (.A(_06331_),
    .B(_06335_),
    .Y(_06336_));
 sg13g2_nand2_1 _14376_ (.Y(_06337_),
    .A(_06207_),
    .B(\ppu.pal[15][3] ));
 sg13g2_nand3_1 _14377_ (.B(_06182_),
    .C(\ppu.pal[13][3] ),
    .A(_06204_),
    .Y(_06338_));
 sg13g2_nand2_1 _14378_ (.Y(_06339_),
    .A(_06337_),
    .B(_06338_));
 sg13g2_nand2_1 _14379_ (.Y(_06340_),
    .A(_06209_),
    .B(\ppu.pal[14][3] ));
 sg13g2_nand3_1 _14380_ (.B(_06141_),
    .C(\ppu.pal[12][3] ),
    .A(_06204_),
    .Y(_06341_));
 sg13g2_nand2_1 _14381_ (.Y(_06342_),
    .A(_06340_),
    .B(_06341_));
 sg13g2_nor2_1 _14382_ (.A(_06339_),
    .B(_06342_),
    .Y(_06343_));
 sg13g2_nand2_1 _14383_ (.Y(_06344_),
    .A(_06336_),
    .B(_06343_));
 sg13g2_nor2_1 _14384_ (.A(_06328_),
    .B(_06344_),
    .Y(_06345_));
 sg13g2_nand2_1 _14385_ (.Y(_06346_),
    .A(_06217_),
    .B(\ppu.pal[0][3] ));
 sg13g2_nand3_1 _14386_ (.B(_06216_),
    .C(_06346_),
    .A(_06345_),
    .Y(_06347_));
 sg13g2_buf_2 _14387_ (.A(_06347_),
    .X(_06348_));
 sg13g2_buf_1 _14388_ (.A(_06348_),
    .X(_06349_));
 sg13g2_nor2_1 _14389_ (.A(net320),
    .B(_02405_),
    .Y(_06350_));
 sg13g2_a21oi_1 _14390_ (.A1(net320),
    .A2(_02417_),
    .Y(_06351_),
    .B1(_06350_));
 sg13g2_nand2_1 _14391_ (.Y(_06352_),
    .A(_06215_),
    .B(_06351_));
 sg13g2_buf_2 _14392_ (.A(_06352_),
    .X(_06353_));
 sg13g2_buf_1 _14393_ (.A(_06353_),
    .X(_06354_));
 sg13g2_nand3_1 _14394_ (.B(_06217_),
    .C(net112),
    .A(net38),
    .Y(_06355_));
 sg13g2_nand2_1 _14395_ (.Y(_06356_),
    .A(net70),
    .B(\ppu.pal[0][7] ));
 sg13g2_nand2_1 _14396_ (.Y(_00306_),
    .A(_06355_),
    .B(_06356_));
 sg13g2_mux2_1 _14397_ (.A0(\ppu.pal[10][0] ),
    .A1(\ppu.pal[10][4] ),
    .S(net80),
    .X(_00307_));
 sg13g2_mux2_1 _14398_ (.A0(\ppu.pal[10][1] ),
    .A1(\ppu.pal[10][5] ),
    .S(_06197_),
    .X(_00308_));
 sg13g2_mux2_1 _14399_ (.A0(\ppu.pal[10][2] ),
    .A1(\ppu.pal[10][6] ),
    .S(net80),
    .X(_00309_));
 sg13g2_mux2_1 _14400_ (.A0(\ppu.pal[10][3] ),
    .A1(\ppu.pal[10][7] ),
    .S(net80),
    .X(_00310_));
 sg13g2_nand3_1 _14401_ (.B(net80),
    .C(net115),
    .A(net41),
    .Y(_06357_));
 sg13g2_inv_1 _14402_ (.Y(_06358_),
    .A(net80));
 sg13g2_nand2_1 _14403_ (.Y(_06359_),
    .A(_06358_),
    .B(\ppu.pal[10][4] ));
 sg13g2_nand2_1 _14404_ (.Y(_00311_),
    .A(_06357_),
    .B(_06359_));
 sg13g2_nand3_1 _14405_ (.B(_06197_),
    .C(net114),
    .A(net40),
    .Y(_06360_));
 sg13g2_nand2_1 _14406_ (.Y(_06361_),
    .A(_06358_),
    .B(\ppu.pal[10][5] ));
 sg13g2_nand2_1 _14407_ (.Y(_00312_),
    .A(_06360_),
    .B(_06361_));
 sg13g2_nand3_1 _14408_ (.B(net80),
    .C(net113),
    .A(net39),
    .Y(_06362_));
 sg13g2_nand2_1 _14409_ (.Y(_06363_),
    .A(_06358_),
    .B(\ppu.pal[10][6] ));
 sg13g2_nand2_1 _14410_ (.Y(_00313_),
    .A(_06362_),
    .B(_06363_));
 sg13g2_nand3_1 _14411_ (.B(net80),
    .C(net112),
    .A(net38),
    .Y(_06364_));
 sg13g2_nand2_1 _14412_ (.Y(_06365_),
    .A(_06358_),
    .B(\ppu.pal[10][7] ));
 sg13g2_nand2_1 _14413_ (.Y(_00314_),
    .A(_06364_),
    .B(_06365_));
 sg13g2_mux2_1 _14414_ (.A0(\ppu.pal[11][0] ),
    .A1(\ppu.pal[11][4] ),
    .S(net81),
    .X(_00315_));
 sg13g2_mux2_1 _14415_ (.A0(\ppu.pal[11][1] ),
    .A1(\ppu.pal[11][5] ),
    .S(net81),
    .X(_00316_));
 sg13g2_mux2_1 _14416_ (.A0(\ppu.pal[11][2] ),
    .A1(\ppu.pal[11][6] ),
    .S(_06194_),
    .X(_00317_));
 sg13g2_mux2_1 _14417_ (.A0(\ppu.pal[11][3] ),
    .A1(\ppu.pal[11][7] ),
    .S(net81),
    .X(_00318_));
 sg13g2_nand3_1 _14418_ (.B(net81),
    .C(net115),
    .A(net41),
    .Y(_06366_));
 sg13g2_inv_1 _14419_ (.Y(_06367_),
    .A(net81));
 sg13g2_nand2_1 _14420_ (.Y(_06368_),
    .A(_06367_),
    .B(\ppu.pal[11][4] ));
 sg13g2_nand2_1 _14421_ (.Y(_00319_),
    .A(_06366_),
    .B(_06368_));
 sg13g2_nand3_1 _14422_ (.B(net81),
    .C(net114),
    .A(net40),
    .Y(_06369_));
 sg13g2_nand2_1 _14423_ (.Y(_06370_),
    .A(_06367_),
    .B(\ppu.pal[11][5] ));
 sg13g2_nand2_1 _14424_ (.Y(_00320_),
    .A(_06369_),
    .B(_06370_));
 sg13g2_nand3_1 _14425_ (.B(_06194_),
    .C(net113),
    .A(net39),
    .Y(_06371_));
 sg13g2_nand2_1 _14426_ (.Y(_06372_),
    .A(_06367_),
    .B(\ppu.pal[11][6] ));
 sg13g2_nand2_1 _14427_ (.Y(_00321_),
    .A(_06371_),
    .B(_06372_));
 sg13g2_nand3_1 _14428_ (.B(net81),
    .C(net112),
    .A(net38),
    .Y(_06373_));
 sg13g2_nand2_1 _14429_ (.Y(_06374_),
    .A(_06367_),
    .B(\ppu.pal[11][7] ));
 sg13g2_nand2_1 _14430_ (.Y(_00322_),
    .A(_06373_),
    .B(_06374_));
 sg13g2_nand2_1 _14431_ (.Y(_06375_),
    .A(_06204_),
    .B(_06154_));
 sg13g2_buf_1 _14432_ (.A(_06375_),
    .X(_06376_));
 sg13g2_mux2_1 _14433_ (.A0(\ppu.pal[12][4] ),
    .A1(\ppu.pal[12][0] ),
    .S(net64),
    .X(_00323_));
 sg13g2_mux2_1 _14434_ (.A0(\ppu.pal[12][5] ),
    .A1(\ppu.pal[12][1] ),
    .S(net64),
    .X(_00324_));
 sg13g2_mux2_1 _14435_ (.A0(\ppu.pal[12][6] ),
    .A1(\ppu.pal[12][2] ),
    .S(net64),
    .X(_00325_));
 sg13g2_mux2_1 _14436_ (.A0(\ppu.pal[12][7] ),
    .A1(\ppu.pal[12][3] ),
    .S(net64),
    .X(_00326_));
 sg13g2_inv_1 _14437_ (.Y(_06377_),
    .A(net64));
 sg13g2_nand3_1 _14438_ (.B(_06377_),
    .C(_06227_),
    .A(_06221_),
    .Y(_06378_));
 sg13g2_nand2_1 _14439_ (.Y(_06379_),
    .A(_06376_),
    .B(\ppu.pal[12][4] ));
 sg13g2_nand2_1 _14440_ (.Y(_00327_),
    .A(_06378_),
    .B(_06379_));
 sg13g2_nand3_1 _14441_ (.B(_06377_),
    .C(net114),
    .A(net40),
    .Y(_06380_));
 sg13g2_nand2_1 _14442_ (.Y(_06381_),
    .A(net64),
    .B(\ppu.pal[12][5] ));
 sg13g2_nand2_1 _14443_ (.Y(_00328_),
    .A(_06380_),
    .B(_06381_));
 sg13g2_nand3_1 _14444_ (.B(_06377_),
    .C(_06313_),
    .A(_06308_),
    .Y(_06382_));
 sg13g2_nand2_1 _14445_ (.Y(_06383_),
    .A(net64),
    .B(\ppu.pal[12][6] ));
 sg13g2_nand2_1 _14446_ (.Y(_00329_),
    .A(_06382_),
    .B(_06383_));
 sg13g2_nand3_1 _14447_ (.B(_06377_),
    .C(net112),
    .A(net38),
    .Y(_06384_));
 sg13g2_nand2_1 _14448_ (.Y(_06385_),
    .A(net64),
    .B(\ppu.pal[12][7] ));
 sg13g2_nand2_1 _14449_ (.Y(_00330_),
    .A(_06384_),
    .B(_06385_));
 sg13g2_mux2_1 _14450_ (.A0(\ppu.pal[13][0] ),
    .A1(\ppu.pal[13][4] ),
    .S(net79),
    .X(_00331_));
 sg13g2_mux2_1 _14451_ (.A0(\ppu.pal[13][1] ),
    .A1(\ppu.pal[13][5] ),
    .S(net79),
    .X(_00332_));
 sg13g2_mux2_1 _14452_ (.A0(\ppu.pal[13][2] ),
    .A1(\ppu.pal[13][6] ),
    .S(_06246_),
    .X(_00333_));
 sg13g2_mux2_1 _14453_ (.A0(\ppu.pal[13][3] ),
    .A1(\ppu.pal[13][7] ),
    .S(net79),
    .X(_00334_));
 sg13g2_nand3_1 _14454_ (.B(net79),
    .C(net115),
    .A(net41),
    .Y(_06386_));
 sg13g2_inv_1 _14455_ (.Y(_06387_),
    .A(net79));
 sg13g2_nand2_1 _14456_ (.Y(_06388_),
    .A(_06387_),
    .B(\ppu.pal[13][4] ));
 sg13g2_nand2_1 _14457_ (.Y(_00335_),
    .A(_06386_),
    .B(_06388_));
 sg13g2_nand3_1 _14458_ (.B(net79),
    .C(net114),
    .A(net40),
    .Y(_06389_));
 sg13g2_nand2_1 _14459_ (.Y(_06390_),
    .A(_06387_),
    .B(\ppu.pal[13][5] ));
 sg13g2_nand2_1 _14460_ (.Y(_00336_),
    .A(_06389_),
    .B(_06390_));
 sg13g2_nand3_1 _14461_ (.B(_06246_),
    .C(net113),
    .A(net39),
    .Y(_06391_));
 sg13g2_nand2_1 _14462_ (.Y(_06392_),
    .A(_06387_),
    .B(\ppu.pal[13][6] ));
 sg13g2_nand2_1 _14463_ (.Y(_00337_),
    .A(_06391_),
    .B(_06392_));
 sg13g2_nand3_1 _14464_ (.B(net79),
    .C(net112),
    .A(net38),
    .Y(_06393_));
 sg13g2_nand2_1 _14465_ (.Y(_06394_),
    .A(_06387_),
    .B(\ppu.pal[13][7] ));
 sg13g2_nand2_1 _14466_ (.Y(_00338_),
    .A(_06393_),
    .B(_06394_));
 sg13g2_mux2_1 _14467_ (.A0(\ppu.pal[14][0] ),
    .A1(\ppu.pal[14][4] ),
    .S(_06292_),
    .X(_00339_));
 sg13g2_mux2_1 _14468_ (.A0(\ppu.pal[14][1] ),
    .A1(\ppu.pal[14][5] ),
    .S(net75),
    .X(_00340_));
 sg13g2_mux2_1 _14469_ (.A0(\ppu.pal[14][2] ),
    .A1(\ppu.pal[14][6] ),
    .S(net75),
    .X(_00341_));
 sg13g2_mux2_1 _14470_ (.A0(\ppu.pal[14][3] ),
    .A1(\ppu.pal[14][7] ),
    .S(net75),
    .X(_00342_));
 sg13g2_nand3_1 _14471_ (.B(net75),
    .C(net115),
    .A(net41),
    .Y(_06395_));
 sg13g2_inv_1 _14472_ (.Y(_06396_),
    .A(net75));
 sg13g2_nand2_1 _14473_ (.Y(_06397_),
    .A(_06396_),
    .B(\ppu.pal[14][4] ));
 sg13g2_nand2_1 _14474_ (.Y(_00343_),
    .A(_06395_),
    .B(_06397_));
 sg13g2_nand3_1 _14475_ (.B(net75),
    .C(_06268_),
    .A(_06263_),
    .Y(_06398_));
 sg13g2_nand2_1 _14476_ (.Y(_06399_),
    .A(_06396_),
    .B(\ppu.pal[14][5] ));
 sg13g2_nand2_1 _14477_ (.Y(_00344_),
    .A(_06398_),
    .B(_06399_));
 sg13g2_nand3_1 _14478_ (.B(net75),
    .C(_06313_),
    .A(_06308_),
    .Y(_06400_));
 sg13g2_nand2_1 _14479_ (.Y(_06401_),
    .A(_06396_),
    .B(\ppu.pal[14][6] ));
 sg13g2_nand2_1 _14480_ (.Y(_00345_),
    .A(_06400_),
    .B(_06401_));
 sg13g2_nand3_1 _14481_ (.B(_06292_),
    .C(_06354_),
    .A(_06349_),
    .Y(_06402_));
 sg13g2_nand2_1 _14482_ (.Y(_06403_),
    .A(_06396_),
    .B(\ppu.pal[14][7] ));
 sg13g2_nand2_1 _14483_ (.Y(_00346_),
    .A(_06402_),
    .B(_06403_));
 sg13g2_mux2_1 _14484_ (.A0(\ppu.pal[15][0] ),
    .A1(\ppu.pal[15][4] ),
    .S(net76),
    .X(_00347_));
 sg13g2_mux2_1 _14485_ (.A0(\ppu.pal[15][1] ),
    .A1(\ppu.pal[15][5] ),
    .S(_06290_),
    .X(_00348_));
 sg13g2_mux2_1 _14486_ (.A0(\ppu.pal[15][2] ),
    .A1(\ppu.pal[15][6] ),
    .S(net76),
    .X(_00349_));
 sg13g2_mux2_1 _14487_ (.A0(\ppu.pal[15][3] ),
    .A1(\ppu.pal[15][7] ),
    .S(_06290_),
    .X(_00350_));
 sg13g2_nand3_1 _14488_ (.B(net76),
    .C(_06227_),
    .A(_06221_),
    .Y(_06404_));
 sg13g2_inv_1 _14489_ (.Y(_06405_),
    .A(net76));
 sg13g2_nand2_1 _14490_ (.Y(_06406_),
    .A(_06405_),
    .B(\ppu.pal[15][4] ));
 sg13g2_nand2_1 _14491_ (.Y(_00351_),
    .A(_06404_),
    .B(_06406_));
 sg13g2_nand3_1 _14492_ (.B(net76),
    .C(_06268_),
    .A(_06263_),
    .Y(_06407_));
 sg13g2_nand2_1 _14493_ (.Y(_06408_),
    .A(_06405_),
    .B(\ppu.pal[15][5] ));
 sg13g2_nand2_1 _14494_ (.Y(_00352_),
    .A(_06407_),
    .B(_06408_));
 sg13g2_nand3_1 _14495_ (.B(net76),
    .C(net113),
    .A(net39),
    .Y(_06409_));
 sg13g2_nand2_1 _14496_ (.Y(_06410_),
    .A(_06405_),
    .B(\ppu.pal[15][6] ));
 sg13g2_nand2_1 _14497_ (.Y(_00353_),
    .A(_06409_),
    .B(_06410_));
 sg13g2_nand3_1 _14498_ (.B(net76),
    .C(_06354_),
    .A(_06349_),
    .Y(_06411_));
 sg13g2_nand2_1 _14499_ (.Y(_06412_),
    .A(_06405_),
    .B(\ppu.pal[15][7] ));
 sg13g2_nand2_1 _14500_ (.Y(_00354_),
    .A(_06411_),
    .B(_06412_));
 sg13g2_mux2_1 _14501_ (.A0(\ppu.pal[1][4] ),
    .A1(\ppu.pal[1][0] ),
    .S(net77),
    .X(_00355_));
 sg13g2_mux2_1 _14502_ (.A0(\ppu.pal[1][5] ),
    .A1(\ppu.pal[1][1] ),
    .S(net77),
    .X(_00356_));
 sg13g2_mux2_1 _14503_ (.A0(\ppu.pal[1][6] ),
    .A1(\ppu.pal[1][2] ),
    .S(net77),
    .X(_00357_));
 sg13g2_mux2_1 _14504_ (.A0(\ppu.pal[1][7] ),
    .A1(\ppu.pal[1][3] ),
    .S(net77),
    .X(_00358_));
 sg13g2_inv_1 _14505_ (.Y(_06413_),
    .A(net77));
 sg13g2_nand3_1 _14506_ (.B(_06413_),
    .C(net115),
    .A(net41),
    .Y(_06414_));
 sg13g2_nand2_1 _14507_ (.Y(_06415_),
    .A(net77),
    .B(\ppu.pal[1][4] ));
 sg13g2_nand2_1 _14508_ (.Y(_00359_),
    .A(_06414_),
    .B(_06415_));
 sg13g2_nand3_1 _14509_ (.B(_06413_),
    .C(net114),
    .A(net40),
    .Y(_06416_));
 sg13g2_nand2_1 _14510_ (.Y(_06417_),
    .A(net77),
    .B(\ppu.pal[1][5] ));
 sg13g2_nand2_1 _14511_ (.Y(_00360_),
    .A(_06416_),
    .B(_06417_));
 sg13g2_nand3_1 _14512_ (.B(_06413_),
    .C(net113),
    .A(net39),
    .Y(_06418_));
 sg13g2_nand2_1 _14513_ (.Y(_06419_),
    .A(net77),
    .B(\ppu.pal[1][6] ));
 sg13g2_nand2_1 _14514_ (.Y(_00361_),
    .A(_06418_),
    .B(_06419_));
 sg13g2_nand3_1 _14515_ (.B(_06413_),
    .C(net112),
    .A(net38),
    .Y(_06420_));
 sg13g2_nand2_1 _14516_ (.Y(_06421_),
    .A(_06280_),
    .B(\ppu.pal[1][7] ));
 sg13g2_nand2_1 _14517_ (.Y(_00362_),
    .A(_06420_),
    .B(_06421_));
 sg13g2_nand2_1 _14518_ (.Y(_06422_),
    .A(net90),
    .B(_06180_));
 sg13g2_buf_1 _14519_ (.A(_06422_),
    .X(_06423_));
 sg13g2_mux2_1 _14520_ (.A0(\ppu.pal[2][4] ),
    .A1(\ppu.pal[2][0] ),
    .S(net69),
    .X(_00363_));
 sg13g2_mux2_1 _14521_ (.A0(\ppu.pal[2][5] ),
    .A1(\ppu.pal[2][1] ),
    .S(net69),
    .X(_00364_));
 sg13g2_mux2_1 _14522_ (.A0(\ppu.pal[2][6] ),
    .A1(\ppu.pal[2][2] ),
    .S(net69),
    .X(_00365_));
 sg13g2_mux2_1 _14523_ (.A0(\ppu.pal[2][7] ),
    .A1(\ppu.pal[2][3] ),
    .S(net69),
    .X(_00366_));
 sg13g2_inv_1 _14524_ (.Y(_06424_),
    .A(net69));
 sg13g2_nand3_1 _14525_ (.B(_06424_),
    .C(net115),
    .A(net41),
    .Y(_06425_));
 sg13g2_nand2_1 _14526_ (.Y(_06426_),
    .A(net69),
    .B(\ppu.pal[2][4] ));
 sg13g2_nand2_1 _14527_ (.Y(_00367_),
    .A(_06425_),
    .B(_06426_));
 sg13g2_nand3_1 _14528_ (.B(_06424_),
    .C(net114),
    .A(net40),
    .Y(_06427_));
 sg13g2_nand2_1 _14529_ (.Y(_06428_),
    .A(net69),
    .B(\ppu.pal[2][5] ));
 sg13g2_nand2_1 _14530_ (.Y(_00368_),
    .A(_06427_),
    .B(_06428_));
 sg13g2_nand3_1 _14531_ (.B(_06424_),
    .C(net113),
    .A(net39),
    .Y(_06429_));
 sg13g2_nand2_1 _14532_ (.Y(_06430_),
    .A(net69),
    .B(\ppu.pal[2][6] ));
 sg13g2_nand2_1 _14533_ (.Y(_00369_),
    .A(_06429_),
    .B(_06430_));
 sg13g2_nand3_1 _14534_ (.B(_06424_),
    .C(net112),
    .A(net38),
    .Y(_06431_));
 sg13g2_nand2_1 _14535_ (.Y(_06432_),
    .A(_06423_),
    .B(\ppu.pal[2][7] ));
 sg13g2_nand2_1 _14536_ (.Y(_00370_),
    .A(_06431_),
    .B(_06432_));
 sg13g2_mux2_1 _14537_ (.A0(\ppu.pal[3][4] ),
    .A1(\ppu.pal[3][0] ),
    .S(net82),
    .X(_00371_));
 sg13g2_mux2_1 _14538_ (.A0(\ppu.pal[3][5] ),
    .A1(\ppu.pal[3][1] ),
    .S(net82),
    .X(_00372_));
 sg13g2_mux2_1 _14539_ (.A0(\ppu.pal[3][6] ),
    .A1(\ppu.pal[3][2] ),
    .S(net82),
    .X(_00373_));
 sg13g2_mux2_1 _14540_ (.A0(\ppu.pal[3][7] ),
    .A1(\ppu.pal[3][3] ),
    .S(net82),
    .X(_00374_));
 sg13g2_inv_1 _14541_ (.Y(_06433_),
    .A(net82));
 sg13g2_nand3_1 _14542_ (.B(_06433_),
    .C(net115),
    .A(net41),
    .Y(_06434_));
 sg13g2_nand2_1 _14543_ (.Y(_06435_),
    .A(net82),
    .B(\ppu.pal[3][4] ));
 sg13g2_nand2_1 _14544_ (.Y(_00375_),
    .A(_06434_),
    .B(_06435_));
 sg13g2_nand3_1 _14545_ (.B(_06433_),
    .C(net114),
    .A(net40),
    .Y(_06436_));
 sg13g2_nand2_1 _14546_ (.Y(_06437_),
    .A(_06178_),
    .B(\ppu.pal[3][5] ));
 sg13g2_nand2_1 _14547_ (.Y(_00376_),
    .A(_06436_),
    .B(_06437_));
 sg13g2_nand3_1 _14548_ (.B(_06433_),
    .C(net113),
    .A(net39),
    .Y(_06438_));
 sg13g2_nand2_1 _14549_ (.Y(_06439_),
    .A(net82),
    .B(\ppu.pal[3][6] ));
 sg13g2_nand2_1 _14550_ (.Y(_00377_),
    .A(_06438_),
    .B(_06439_));
 sg13g2_nand3_1 _14551_ (.B(_06433_),
    .C(net112),
    .A(net38),
    .Y(_06440_));
 sg13g2_nand2_1 _14552_ (.Y(_06441_),
    .A(net82),
    .B(\ppu.pal[3][7] ));
 sg13g2_nand2_1 _14553_ (.Y(_00378_),
    .A(_06440_),
    .B(_06441_));
 sg13g2_nand2_1 _14554_ (.Y(_06442_),
    .A(net85),
    .B(_06159_));
 sg13g2_buf_1 _14555_ (.A(_06442_),
    .X(_06443_));
 sg13g2_mux2_1 _14556_ (.A0(\ppu.pal[4][4] ),
    .A1(\ppu.pal[4][0] ),
    .S(net63),
    .X(_00379_));
 sg13g2_mux2_1 _14557_ (.A0(\ppu.pal[4][5] ),
    .A1(\ppu.pal[4][1] ),
    .S(net63),
    .X(_00380_));
 sg13g2_mux2_1 _14558_ (.A0(\ppu.pal[4][6] ),
    .A1(\ppu.pal[4][2] ),
    .S(net63),
    .X(_00381_));
 sg13g2_mux2_1 _14559_ (.A0(\ppu.pal[4][7] ),
    .A1(\ppu.pal[4][3] ),
    .S(net63),
    .X(_00382_));
 sg13g2_inv_1 _14560_ (.Y(_06444_),
    .A(_06443_));
 sg13g2_nand3_1 _14561_ (.B(_06444_),
    .C(_06226_),
    .A(_06220_),
    .Y(_06445_));
 sg13g2_nand2_1 _14562_ (.Y(_06446_),
    .A(net63),
    .B(\ppu.pal[4][4] ));
 sg13g2_nand2_1 _14563_ (.Y(_00383_),
    .A(_06445_),
    .B(_06446_));
 sg13g2_nand3_1 _14564_ (.B(_06444_),
    .C(_06267_),
    .A(_06262_),
    .Y(_06447_));
 sg13g2_nand2_1 _14565_ (.Y(_06448_),
    .A(net63),
    .B(\ppu.pal[4][5] ));
 sg13g2_nand2_1 _14566_ (.Y(_00384_),
    .A(_06447_),
    .B(_06448_));
 sg13g2_nand3_1 _14567_ (.B(_06444_),
    .C(_06312_),
    .A(_06307_),
    .Y(_06449_));
 sg13g2_nand2_1 _14568_ (.Y(_06450_),
    .A(net63),
    .B(\ppu.pal[4][6] ));
 sg13g2_nand2_1 _14569_ (.Y(_00385_),
    .A(_06449_),
    .B(_06450_));
 sg13g2_nand3_1 _14570_ (.B(_06444_),
    .C(_06353_),
    .A(_06348_),
    .Y(_06451_));
 sg13g2_nand2_1 _14571_ (.Y(_06452_),
    .A(net63),
    .B(\ppu.pal[4][7] ));
 sg13g2_nand2_1 _14572_ (.Y(_00386_),
    .A(_06451_),
    .B(_06452_));
 sg13g2_mux2_1 _14573_ (.A0(\ppu.pal[5][0] ),
    .A1(\ppu.pal[5][4] ),
    .S(net78),
    .X(_00387_));
 sg13g2_mux2_1 _14574_ (.A0(\ppu.pal[5][1] ),
    .A1(\ppu.pal[5][5] ),
    .S(net78),
    .X(_00388_));
 sg13g2_mux2_1 _14575_ (.A0(\ppu.pal[5][2] ),
    .A1(\ppu.pal[5][6] ),
    .S(net78),
    .X(_00389_));
 sg13g2_mux2_1 _14576_ (.A0(\ppu.pal[5][3] ),
    .A1(\ppu.pal[5][7] ),
    .S(net78),
    .X(_00390_));
 sg13g2_nand3_1 _14577_ (.B(_06274_),
    .C(_06226_),
    .A(_06220_),
    .Y(_06453_));
 sg13g2_inv_1 _14578_ (.Y(_06454_),
    .A(_06274_));
 sg13g2_nand2_1 _14579_ (.Y(_06455_),
    .A(_06454_),
    .B(\ppu.pal[5][4] ));
 sg13g2_nand2_1 _14580_ (.Y(_00391_),
    .A(_06453_),
    .B(_06455_));
 sg13g2_nand3_1 _14581_ (.B(net78),
    .C(_06267_),
    .A(_06262_),
    .Y(_06456_));
 sg13g2_nand2_1 _14582_ (.Y(_06457_),
    .A(_06454_),
    .B(\ppu.pal[5][5] ));
 sg13g2_nand2_1 _14583_ (.Y(_00392_),
    .A(_06456_),
    .B(_06457_));
 sg13g2_nand3_1 _14584_ (.B(net78),
    .C(_06312_),
    .A(_06307_),
    .Y(_06458_));
 sg13g2_nand2_1 _14585_ (.Y(_06459_),
    .A(_06454_),
    .B(\ppu.pal[5][6] ));
 sg13g2_nand2_1 _14586_ (.Y(_00393_),
    .A(_06458_),
    .B(_06459_));
 sg13g2_nand3_1 _14587_ (.B(net78),
    .C(_06353_),
    .A(_06348_),
    .Y(_06460_));
 sg13g2_nand2_1 _14588_ (.Y(_06461_),
    .A(_06454_),
    .B(\ppu.pal[5][7] ));
 sg13g2_nand2_1 _14589_ (.Y(_00394_),
    .A(_06460_),
    .B(_06461_));
 sg13g2_mux2_1 _14590_ (.A0(\ppu.pal[6][0] ),
    .A1(\ppu.pal[6][4] ),
    .S(net84),
    .X(_00395_));
 sg13g2_mux2_1 _14591_ (.A0(\ppu.pal[6][1] ),
    .A1(\ppu.pal[6][5] ),
    .S(_06167_),
    .X(_00396_));
 sg13g2_mux2_1 _14592_ (.A0(\ppu.pal[6][2] ),
    .A1(\ppu.pal[6][6] ),
    .S(net84),
    .X(_00397_));
 sg13g2_mux2_1 _14593_ (.A0(\ppu.pal[6][3] ),
    .A1(\ppu.pal[6][7] ),
    .S(net84),
    .X(_00398_));
 sg13g2_nand3_1 _14594_ (.B(net84),
    .C(_06226_),
    .A(_06220_),
    .Y(_06462_));
 sg13g2_inv_1 _14595_ (.Y(_06463_),
    .A(net84));
 sg13g2_nand2_1 _14596_ (.Y(_06464_),
    .A(_06463_),
    .B(\ppu.pal[6][4] ));
 sg13g2_nand2_1 _14597_ (.Y(_00399_),
    .A(_06462_),
    .B(_06464_));
 sg13g2_nand3_1 _14598_ (.B(net84),
    .C(_06267_),
    .A(_06262_),
    .Y(_06465_));
 sg13g2_nand2_1 _14599_ (.Y(_06466_),
    .A(_06463_),
    .B(\ppu.pal[6][5] ));
 sg13g2_nand2_1 _14600_ (.Y(_00400_),
    .A(_06465_),
    .B(_06466_));
 sg13g2_nand3_1 _14601_ (.B(net84),
    .C(_06312_),
    .A(_06307_),
    .Y(_06467_));
 sg13g2_nand2_1 _14602_ (.Y(_06468_),
    .A(_06463_),
    .B(\ppu.pal[6][6] ));
 sg13g2_nand2_1 _14603_ (.Y(_00401_),
    .A(_06467_),
    .B(_06468_));
 sg13g2_nand3_1 _14604_ (.B(_06167_),
    .C(_06353_),
    .A(_06348_),
    .Y(_06469_));
 sg13g2_nand2_1 _14605_ (.Y(_06470_),
    .A(_06463_),
    .B(\ppu.pal[6][7] ));
 sg13g2_nand2_1 _14606_ (.Y(_00402_),
    .A(_06469_),
    .B(_06470_));
 sg13g2_mux2_1 _14607_ (.A0(\ppu.pal[7][0] ),
    .A1(\ppu.pal[7][4] ),
    .S(net83),
    .X(_00403_));
 sg13g2_mux2_1 _14608_ (.A0(\ppu.pal[7][1] ),
    .A1(\ppu.pal[7][5] ),
    .S(net83),
    .X(_00404_));
 sg13g2_mux2_1 _14609_ (.A0(\ppu.pal[7][2] ),
    .A1(\ppu.pal[7][6] ),
    .S(_06171_),
    .X(_00405_));
 sg13g2_mux2_1 _14610_ (.A0(\ppu.pal[7][3] ),
    .A1(\ppu.pal[7][7] ),
    .S(_06171_),
    .X(_00406_));
 sg13g2_nand3_1 _14611_ (.B(net83),
    .C(_06226_),
    .A(_06220_),
    .Y(_06471_));
 sg13g2_inv_1 _14612_ (.Y(_06472_),
    .A(net83));
 sg13g2_nand2_1 _14613_ (.Y(_06473_),
    .A(_06472_),
    .B(\ppu.pal[7][4] ));
 sg13g2_nand2_1 _14614_ (.Y(_00407_),
    .A(_06471_),
    .B(_06473_));
 sg13g2_nand3_1 _14615_ (.B(net83),
    .C(_06267_),
    .A(_06262_),
    .Y(_06474_));
 sg13g2_nand2_1 _14616_ (.Y(_06475_),
    .A(_06472_),
    .B(\ppu.pal[7][5] ));
 sg13g2_nand2_1 _14617_ (.Y(_00408_),
    .A(_06474_),
    .B(_06475_));
 sg13g2_nand3_1 _14618_ (.B(net83),
    .C(_06312_),
    .A(_06307_),
    .Y(_06476_));
 sg13g2_nand2_1 _14619_ (.Y(_06477_),
    .A(_06472_),
    .B(\ppu.pal[7][6] ));
 sg13g2_nand2_1 _14620_ (.Y(_00409_),
    .A(_06476_),
    .B(_06477_));
 sg13g2_nand3_1 _14621_ (.B(net83),
    .C(_06353_),
    .A(_06348_),
    .Y(_06478_));
 sg13g2_nand2_1 _14622_ (.Y(_06479_),
    .A(_06472_),
    .B(\ppu.pal[7][7] ));
 sg13g2_nand2_1 _14623_ (.Y(_00410_),
    .A(_06478_),
    .B(_06479_));
 sg13g2_nand2_1 _14624_ (.Y(_06480_),
    .A(net85),
    .B(_06190_));
 sg13g2_buf_1 _14625_ (.A(_06480_),
    .X(_06481_));
 sg13g2_mux2_1 _14626_ (.A0(\ppu.pal[8][4] ),
    .A1(\ppu.pal[8][0] ),
    .S(net62),
    .X(_00411_));
 sg13g2_mux2_1 _14627_ (.A0(\ppu.pal[8][5] ),
    .A1(\ppu.pal[8][1] ),
    .S(net62),
    .X(_00412_));
 sg13g2_mux2_1 _14628_ (.A0(\ppu.pal[8][6] ),
    .A1(\ppu.pal[8][2] ),
    .S(_06481_),
    .X(_00413_));
 sg13g2_mux2_1 _14629_ (.A0(\ppu.pal[8][7] ),
    .A1(\ppu.pal[8][3] ),
    .S(net62),
    .X(_00414_));
 sg13g2_inv_1 _14630_ (.Y(_06482_),
    .A(net62));
 sg13g2_nand3_1 _14631_ (.B(_06482_),
    .C(_06226_),
    .A(_06220_),
    .Y(_06483_));
 sg13g2_nand2_1 _14632_ (.Y(_06484_),
    .A(net62),
    .B(\ppu.pal[8][4] ));
 sg13g2_nand2_1 _14633_ (.Y(_00415_),
    .A(_06483_),
    .B(_06484_));
 sg13g2_nand3_1 _14634_ (.B(_06482_),
    .C(_06267_),
    .A(_06262_),
    .Y(_06485_));
 sg13g2_nand2_1 _14635_ (.Y(_06486_),
    .A(net62),
    .B(\ppu.pal[8][5] ));
 sg13g2_nand2_1 _14636_ (.Y(_00416_),
    .A(_06485_),
    .B(_06486_));
 sg13g2_nand3_1 _14637_ (.B(_06482_),
    .C(_06312_),
    .A(_06307_),
    .Y(_06487_));
 sg13g2_nand2_1 _14638_ (.Y(_06488_),
    .A(net62),
    .B(\ppu.pal[8][6] ));
 sg13g2_nand2_1 _14639_ (.Y(_00417_),
    .A(_06487_),
    .B(_06488_));
 sg13g2_nand3_1 _14640_ (.B(_06482_),
    .C(_06353_),
    .A(_06348_),
    .Y(_06489_));
 sg13g2_nand2_1 _14641_ (.Y(_06490_),
    .A(net62),
    .B(\ppu.pal[8][7] ));
 sg13g2_nand2_1 _14642_ (.Y(_00418_),
    .A(_06489_),
    .B(_06490_));
 sg13g2_mux2_1 _14643_ (.A0(\ppu.pal[9][0] ),
    .A1(\ppu.pal[9][4] ),
    .S(net74),
    .X(_00419_));
 sg13g2_mux2_1 _14644_ (.A0(\ppu.pal[9][1] ),
    .A1(\ppu.pal[9][5] ),
    .S(net74),
    .X(_00420_));
 sg13g2_mux2_1 _14645_ (.A0(\ppu.pal[9][2] ),
    .A1(\ppu.pal[9][6] ),
    .S(_06332_),
    .X(_00421_));
 sg13g2_mux2_1 _14646_ (.A0(\ppu.pal[9][3] ),
    .A1(\ppu.pal[9][7] ),
    .S(net74),
    .X(_00422_));
 sg13g2_nand3_1 _14647_ (.B(net74),
    .C(_06226_),
    .A(_06220_),
    .Y(_06491_));
 sg13g2_inv_1 _14648_ (.Y(_06492_),
    .A(net74));
 sg13g2_nand2_1 _14649_ (.Y(_06493_),
    .A(_06492_),
    .B(\ppu.pal[9][4] ));
 sg13g2_nand2_1 _14650_ (.Y(_00423_),
    .A(_06491_),
    .B(_06493_));
 sg13g2_nand3_1 _14651_ (.B(net74),
    .C(_06267_),
    .A(_06262_),
    .Y(_06494_));
 sg13g2_nand2_1 _14652_ (.Y(_06495_),
    .A(_06492_),
    .B(\ppu.pal[9][5] ));
 sg13g2_nand2_1 _14653_ (.Y(_00424_),
    .A(_06494_),
    .B(_06495_));
 sg13g2_nand3_1 _14654_ (.B(net74),
    .C(_06312_),
    .A(_06307_),
    .Y(_06496_));
 sg13g2_nand2_1 _14655_ (.Y(_06497_),
    .A(_06492_),
    .B(\ppu.pal[9][6] ));
 sg13g2_nand2_1 _14656_ (.Y(_00425_),
    .A(_06496_),
    .B(_06497_));
 sg13g2_nand3_1 _14657_ (.B(net74),
    .C(_06353_),
    .A(_06348_),
    .Y(_06498_));
 sg13g2_nand2_1 _14658_ (.Y(_06499_),
    .A(_06492_),
    .B(\ppu.pal[9][7] ));
 sg13g2_nand2_1 _14659_ (.Y(_00426_),
    .A(_06498_),
    .B(_06499_));
 sg13g2_nand2_1 _14660_ (.Y(\ppu.pal_data_out[2] ),
    .A(_06304_),
    .B(_06305_));
 sg13g2_buf_1 _14661_ (.A(\ppu.dither_r.u[1] ),
    .X(_06500_));
 sg13g2_buf_1 _14662_ (.A(_02234_),
    .X(_06501_));
 sg13g2_mux2_1 _14663_ (.A0(_06500_),
    .A1(\ppu.pal_data_out[2] ),
    .S(_06501_),
    .X(_00441_));
 sg13g2_nand2_1 _14664_ (.Y(\ppu.pal_data_out[3] ),
    .A(_06345_),
    .B(_06346_));
 sg13g2_inv_1 _14665_ (.Y(_06502_),
    .A(\ppu.dither_r.u[2] ));
 sg13g2_buf_1 _14666_ (.A(net264),
    .X(_06503_));
 sg13g2_buf_1 _14667_ (.A(net264),
    .X(_06504_));
 sg13g2_nor2_1 _14668_ (.A(net240),
    .B(\ppu.pal_data_out[3] ),
    .Y(_06505_));
 sg13g2_a21oi_1 _14669_ (.A1(_06502_),
    .A2(net241),
    .Y(_00442_),
    .B1(_06505_));
 sg13g2_buf_1 _14670_ (.A(\ppu.b0_out[2] ),
    .X(_06506_));
 sg13g2_inv_1 _14671_ (.Y(_06507_),
    .A(_06506_));
 sg13g2_nor2_1 _14672_ (.A(\ppu.pal_out[0] ),
    .B(net241),
    .Y(_06508_));
 sg13g2_a21oi_1 _14673_ (.A1(_06507_),
    .A2(net241),
    .Y(_00443_),
    .B1(_06508_));
 sg13g2_inv_1 _14674_ (.Y(_06509_),
    .A(\ppu.b0_out[3] ));
 sg13g2_nor2_1 _14675_ (.A(\ppu.pal_out[1] ),
    .B(net240),
    .Y(_06510_));
 sg13g2_a21oi_1 _14676_ (.A1(_06509_),
    .A2(net241),
    .Y(_00444_),
    .B1(_06510_));
 sg13g2_buf_1 _14677_ (.A(\ppu.dither_g.u[0] ),
    .X(_06511_));
 sg13g2_inv_1 _14678_ (.Y(_06512_),
    .A(_06511_));
 sg13g2_nor2_1 _14679_ (.A(\ppu.pal_out[2] ),
    .B(net240),
    .Y(_06513_));
 sg13g2_a21oi_1 _14680_ (.A1(_06512_),
    .A2(net241),
    .Y(_00445_),
    .B1(_06513_));
 sg13g2_buf_1 _14681_ (.A(\ppu.dither_g.u[1] ),
    .X(_06514_));
 sg13g2_inv_1 _14682_ (.Y(_06515_),
    .A(_06514_));
 sg13g2_nor2_1 _14683_ (.A(\ppu.pal_out[3] ),
    .B(net240),
    .Y(_06516_));
 sg13g2_a21oi_1 _14684_ (.A1(_06515_),
    .A2(net241),
    .Y(_00446_),
    .B1(_06516_));
 sg13g2_nand2_1 _14685_ (.Y(\ppu.pal_data_out[0] ),
    .A(_06214_),
    .B(_06218_));
 sg13g2_inv_1 _14686_ (.Y(_06517_),
    .A(\ppu.dither_g.u[2] ));
 sg13g2_nor2_1 _14687_ (.A(net240),
    .B(\ppu.pal_data_out[0] ),
    .Y(_06518_));
 sg13g2_a21oi_1 _14688_ (.A1(_06517_),
    .A2(net241),
    .Y(_00447_),
    .B1(_06518_));
 sg13g2_nand2_1 _14689_ (.Y(\ppu.pal_data_out[1] ),
    .A(_06259_),
    .B(_06260_));
 sg13g2_buf_1 _14690_ (.A(\ppu.b0_out[1] ),
    .X(_06519_));
 sg13g2_inv_1 _14691_ (.Y(_06520_),
    .A(net396));
 sg13g2_nor2_1 _14692_ (.A(net240),
    .B(\ppu.pal_data_out[1] ),
    .Y(_06521_));
 sg13g2_a21oi_1 _14693_ (.A1(_06520_),
    .A2(net241),
    .Y(_00448_),
    .B1(_06521_));
 sg13g2_inv_1 _14694_ (.Y(_06522_),
    .A(\ppu.sprite_buffer.oam_load_sprite_valid ));
 sg13g2_inv_1 _14695_ (.Y(_06523_),
    .A(_02588_));
 sg13g2_nor3_2 _14696_ (.A(_00028_),
    .B(_06523_),
    .C(_02884_),
    .Y(_06524_));
 sg13g2_xor2_1 _14697_ (.B(_06524_),
    .A(_00151_),
    .X(_06525_));
 sg13g2_inv_1 _14698_ (.Y(_06526_),
    .A(\ppu.sprite_buffer.valid_sprites[2] ));
 sg13g2_nand2b_1 _14699_ (.Y(_06527_),
    .B(_06524_),
    .A_N(_00151_));
 sg13g2_xnor2_1 _14700_ (.Y(_06528_),
    .A(_00077_),
    .B(_06527_));
 sg13g2_a21oi_1 _14701_ (.A1(_06525_),
    .A2(_06526_),
    .Y(_06529_),
    .B1(_06528_));
 sg13g2_o21ai_1 _14702_ (.B1(_06529_),
    .Y(_06530_),
    .A1(\ppu.sprite_buffer.valid_sprites[3] ),
    .A2(_06525_));
 sg13g2_inv_1 _14703_ (.Y(_06531_),
    .A(\ppu.sprite_buffer.valid_sprites[0] ));
 sg13g2_o21ai_1 _14704_ (.B1(_06528_),
    .Y(_06532_),
    .A1(\ppu.sprite_buffer.valid_sprites[1] ),
    .A2(_06525_));
 sg13g2_a21oi_1 _14705_ (.A1(_06531_),
    .A2(_06525_),
    .Y(_06533_),
    .B1(_06532_));
 sg13g2_nor2_1 _14706_ (.A(net240),
    .B(_06533_),
    .Y(_06534_));
 sg13g2_a22oi_1 _14707_ (.Y(_00635_),
    .B1(_06530_),
    .B2(_06534_),
    .A2(_06503_),
    .A1(_06522_));
 sg13g2_inv_1 _14708_ (.Y(_06535_),
    .A(_02813_));
 sg13g2_inv_1 _14709_ (.Y(_06536_),
    .A(_02810_));
 sg13g2_nand2_1 _14710_ (.Y(_06537_),
    .A(_02243_),
    .B(_02807_));
 sg13g2_a21oi_1 _14711_ (.A1(_02246_),
    .A2(_06536_),
    .Y(_06538_),
    .B1(_06537_));
 sg13g2_a221oi_1 _14712_ (.B2(_02810_),
    .C1(_06538_),
    .B1(_02245_),
    .A1(\ppu.rs2.y_scan.counter[3] ),
    .Y(_06539_),
    .A2(_02813_));
 sg13g2_a21oi_1 _14713_ (.A1(_02342_),
    .A2(_06535_),
    .Y(_06540_),
    .B1(_06539_));
 sg13g2_xor2_1 _14714_ (.B(_02816_),
    .A(_02242_),
    .X(_06541_));
 sg13g2_nand2b_1 _14715_ (.Y(_06542_),
    .B(_06541_),
    .A_N(_06540_));
 sg13g2_o21ai_1 _14716_ (.B1(_06542_),
    .Y(_06543_),
    .A1(_02242_),
    .A2(_02816_));
 sg13g2_xor2_1 _14717_ (.B(\data_pins[0] ),
    .A(_02241_),
    .X(_06544_));
 sg13g2_nand2_1 _14718_ (.Y(_06545_),
    .A(_06543_),
    .B(_06544_));
 sg13g2_or2_1 _14719_ (.X(_06546_),
    .B(_06543_),
    .A(_06544_));
 sg13g2_xnor2_1 _14720_ (.Y(_06547_),
    .A(_02321_),
    .B(net408));
 sg13g2_o21ai_1 _14721_ (.B1(_06545_),
    .Y(_06548_),
    .A1(_02241_),
    .A2(net405));
 sg13g2_xor2_1 _14722_ (.B(net403),
    .A(_02240_),
    .X(_06549_));
 sg13g2_nand2_1 _14723_ (.Y(_06550_),
    .A(_06548_),
    .B(_06549_));
 sg13g2_o21ai_1 _14724_ (.B1(_06550_),
    .Y(_06551_),
    .A1(_02240_),
    .A2(net403));
 sg13g2_xor2_1 _14725_ (.B(_02489_),
    .A(_02239_),
    .X(_06552_));
 sg13g2_nand2_1 _14726_ (.Y(_06553_),
    .A(_06551_),
    .B(_06552_));
 sg13g2_o21ai_1 _14727_ (.B1(_06553_),
    .Y(_06554_),
    .A1(_02239_),
    .A2(_02489_));
 sg13g2_nor2_1 _14728_ (.A(_06547_),
    .B(_06554_),
    .Y(_06555_));
 sg13g2_a21oi_1 _14729_ (.A1(_06545_),
    .A2(_06546_),
    .Y(_06556_),
    .B1(_06555_));
 sg13g2_nand2_1 _14730_ (.Y(_06557_),
    .A(_06554_),
    .B(_06547_));
 sg13g2_xnor2_1 _14731_ (.Y(_06558_),
    .A(_06552_),
    .B(_06551_));
 sg13g2_nand2b_1 _14732_ (.Y(_06559_),
    .B(_06540_),
    .A_N(_06541_));
 sg13g2_or2_1 _14733_ (.X(_06560_),
    .B(_06548_),
    .A(_06549_));
 sg13g2_nand2_1 _14734_ (.Y(_06561_),
    .A(_01863_),
    .B(net235));
 sg13g2_a221oi_1 _14735_ (.B2(_06550_),
    .C1(_06561_),
    .B1(_06560_),
    .A1(_06542_),
    .Y(_06562_),
    .A2(_06559_));
 sg13g2_nand4_1 _14736_ (.B(_06557_),
    .C(_06558_),
    .A(_06556_),
    .Y(_06563_),
    .D(_06562_));
 sg13g2_o21ai_1 _14737_ (.B1(_06563_),
    .Y(_00821_),
    .A1(_01868_),
    .A2(net235));
 sg13g2_nor4_1 _14738_ (.A(_03198_),
    .B(_03196_),
    .C(_03202_),
    .D(_03200_),
    .Y(_06564_));
 sg13g2_nand2b_1 _14739_ (.Y(_06565_),
    .B(_03210_),
    .A_N(_06564_));
 sg13g2_buf_1 _14740_ (.A(\ppu.display_mask[0] ),
    .X(_06566_));
 sg13g2_nand2_1 _14741_ (.Y(_06567_),
    .A(_06566_),
    .B(\ppu.tilemap.map_pixels[0][1] ));
 sg13g2_nand2_1 _14742_ (.Y(_06568_),
    .A(_06566_),
    .B(\ppu.tilemap.map_pixels[0][0] ));
 sg13g2_nand2_1 _14743_ (.Y(_06569_),
    .A(_06567_),
    .B(_06568_));
 sg13g2_a21oi_1 _14744_ (.A1(_06565_),
    .A2(_06569_),
    .Y(_06570_),
    .B1(\ppu.tilemap.attr[0][0] ));
 sg13g2_nand2_1 _14745_ (.Y(_06571_),
    .A(_06566_),
    .B(\ppu.tilemap.map_pixels[0][3] ));
 sg13g2_nand2_1 _14746_ (.Y(_06572_),
    .A(_06566_),
    .B(\ppu.tilemap.map_pixels[0][2] ));
 sg13g2_nand2_1 _14747_ (.Y(_06573_),
    .A(_06571_),
    .B(_06572_));
 sg13g2_o21ai_1 _14748_ (.B1(_06573_),
    .Y(_06574_),
    .A1(_03210_),
    .A2(_06564_));
 sg13g2_nand2_1 _14749_ (.Y(_06575_),
    .A(_06570_),
    .B(_06574_));
 sg13g2_buf_2 _14750_ (.A(_06575_),
    .X(_06576_));
 sg13g2_nand2_1 _14751_ (.Y(_06577_),
    .A(_06576_),
    .B(_03189_));
 sg13g2_o21ai_1 _14752_ (.B1(_06577_),
    .Y(_06578_),
    .A1(_03248_),
    .A2(_06576_));
 sg13g2_buf_1 _14753_ (.A(\ppu.display_mask[1] ),
    .X(_06579_));
 sg13g2_buf_1 _14754_ (.A(_06576_),
    .X(_06580_));
 sg13g2_a21oi_1 _14755_ (.A1(_06579_),
    .A2(\ppu.tilemap.map_pixels[1][0] ),
    .Y(_06581_),
    .B1(net185));
 sg13g2_nand2_1 _14756_ (.Y(_06582_),
    .A(net185),
    .B(_06568_));
 sg13g2_nand2b_1 _14757_ (.Y(_06583_),
    .B(_06582_),
    .A_N(_06581_));
 sg13g2_inv_1 _14758_ (.Y(_06584_),
    .A(_06576_));
 sg13g2_nor2b_1 _14759_ (.A(_06584_),
    .B_N(_06572_),
    .Y(_06585_));
 sg13g2_a21o_1 _14760_ (.A2(\ppu.tilemap.map_pixels[1][2] ),
    .A1(_06579_),
    .B1(_06576_),
    .X(_06586_));
 sg13g2_nand2b_1 _14761_ (.Y(_06587_),
    .B(_06586_),
    .A_N(_06585_));
 sg13g2_inv_1 _14762_ (.Y(_06588_),
    .A(_06587_));
 sg13g2_nor2_1 _14763_ (.A(_06578_),
    .B(_06588_),
    .Y(_06589_));
 sg13g2_a21o_1 _14764_ (.A2(_06583_),
    .A1(_06578_),
    .B1(_06589_),
    .X(_06590_));
 sg13g2_nor2b_1 _14765_ (.A(_06584_),
    .B_N(_06571_),
    .Y(_06591_));
 sg13g2_a21o_1 _14766_ (.A2(\ppu.tilemap.map_pixels[1][3] ),
    .A1(_06579_),
    .B1(_06576_),
    .X(_06592_));
 sg13g2_nand2b_1 _14767_ (.Y(_06593_),
    .B(_06592_),
    .A_N(_06591_));
 sg13g2_a21oi_1 _14768_ (.A1(_06579_),
    .A2(\ppu.tilemap.map_pixels[1][1] ),
    .Y(_06594_),
    .B1(_06576_));
 sg13g2_nand2_1 _14769_ (.Y(_06595_),
    .A(net185),
    .B(_06567_));
 sg13g2_nand2b_1 _14770_ (.Y(_06596_),
    .B(_06595_),
    .A_N(_06594_));
 sg13g2_mux2_1 _14771_ (.A0(_06593_),
    .A1(_06596_),
    .S(_06578_),
    .X(_06597_));
 sg13g2_buf_1 _14772_ (.A(_06597_),
    .X(_06598_));
 sg13g2_a21oi_1 _14773_ (.A1(_06584_),
    .A2(\ppu.tilemap.attr[1][0] ),
    .Y(_06599_),
    .B1(\ppu.tilemap.attr[0][0] ));
 sg13g2_nand3_1 _14774_ (.B(_06598_),
    .C(_06599_),
    .A(_06590_),
    .Y(_06600_));
 sg13g2_inv_1 _14775_ (.Y(_06601_),
    .A(_06600_));
 sg13g2_nor2_1 _14776_ (.A(\ppu.tilemap.attr[1][2] ),
    .B(_06580_),
    .Y(_06602_));
 sg13g2_a21o_1 _14777_ (.A2(net185),
    .A1(_03198_),
    .B1(_06602_),
    .X(_06603_));
 sg13g2_inv_1 _14778_ (.Y(_06604_),
    .A(_06603_));
 sg13g2_nor2_1 _14779_ (.A(\ppu.tilemap.attr[1][3] ),
    .B(net185),
    .Y(_06605_));
 sg13g2_a21o_1 _14780_ (.A2(net185),
    .A1(_03200_),
    .B1(_06605_),
    .X(_06606_));
 sg13g2_inv_1 _14781_ (.Y(_06607_),
    .A(_06606_));
 sg13g2_nor2_1 _14782_ (.A(\ppu.tilemap.attr[1][1] ),
    .B(_06576_),
    .Y(_06608_));
 sg13g2_a21o_1 _14783_ (.A2(net185),
    .A1(_03196_),
    .B1(_06608_),
    .X(_06609_));
 sg13g2_buf_1 _14784_ (.A(_06609_),
    .X(_06610_));
 sg13g2_inv_1 _14785_ (.Y(_06611_),
    .A(_06610_));
 sg13g2_nor2b_1 _14786_ (.A(net185),
    .B_N(_00162_),
    .Y(_06612_));
 sg13g2_a21oi_1 _14787_ (.A1(_00161_),
    .A2(_06580_),
    .Y(_06613_),
    .B1(_06612_));
 sg13g2_nand4_1 _14788_ (.B(_06607_),
    .C(_06611_),
    .A(_06604_),
    .Y(_06614_),
    .D(_06613_));
 sg13g2_nor2b_1 _14789_ (.A(_06588_),
    .B_N(_06583_),
    .Y(_06615_));
 sg13g2_nand3_1 _14790_ (.B(_06593_),
    .C(_06599_),
    .A(_06615_),
    .Y(_06616_));
 sg13g2_inv_2 _14791_ (.Y(_06617_),
    .A(_06614_));
 sg13g2_nand2_1 _14792_ (.Y(_06618_),
    .A(_06617_),
    .B(_06596_));
 sg13g2_nor2_1 _14793_ (.A(_06616_),
    .B(_06618_),
    .Y(_06619_));
 sg13g2_a21oi_1 _14794_ (.A1(_06601_),
    .A2(_06614_),
    .Y(_06620_),
    .B1(_06619_));
 sg13g2_nand3_1 _14795_ (.B(net206),
    .C(_06584_),
    .A(_06620_),
    .Y(_06621_));
 sg13g2_o21ai_1 _14796_ (.B1(_06621_),
    .Y(_00835_),
    .A1(_06098_),
    .A2(net206));
 sg13g2_nand3b_1 _14797_ (.B(net206),
    .C(_06584_),
    .Y(_06622_),
    .A_N(_06620_));
 sg13g2_o21ai_1 _14798_ (.B1(_06622_),
    .Y(_00836_),
    .A1(_06100_),
    .A2(net206));
 sg13g2_o21ai_1 _14799_ (.B1(_06606_),
    .Y(_06623_),
    .A1(_06603_),
    .A2(_06598_));
 sg13g2_nor2_1 _14800_ (.A(_06603_),
    .B(_06598_),
    .Y(_06624_));
 sg13g2_nand2_1 _14801_ (.Y(_06625_),
    .A(_06624_),
    .B(_06607_));
 sg13g2_nand3_1 _14802_ (.B(_06623_),
    .C(_06625_),
    .A(_06600_),
    .Y(_06626_));
 sg13g2_inv_1 _14803_ (.Y(_06627_),
    .A(_06590_));
 sg13g2_a21oi_1 _14804_ (.A1(_06627_),
    .A2(_06610_),
    .Y(_06628_),
    .B1(_06617_));
 sg13g2_o21ai_1 _14805_ (.B1(_06628_),
    .Y(_06629_),
    .A1(_06610_),
    .A2(_06626_));
 sg13g2_a21oi_1 _14806_ (.A1(_06617_),
    .A2(_06583_),
    .Y(_06630_),
    .B1(net240));
 sg13g2_nand2_1 _14807_ (.Y(_06631_),
    .A(_06629_),
    .B(_06630_));
 sg13g2_o21ai_1 _14808_ (.B1(_06631_),
    .Y(_00879_),
    .A1(_06106_),
    .A2(net206));
 sg13g2_xnor2_1 _14809_ (.Y(_06632_),
    .A(_06613_),
    .B(_06625_));
 sg13g2_nand2_1 _14810_ (.Y(_06633_),
    .A(_06632_),
    .B(_06600_));
 sg13g2_nor2b_1 _14811_ (.A(_06604_),
    .B_N(_06598_),
    .Y(_06634_));
 sg13g2_nor3_1 _14812_ (.A(_06624_),
    .B(_06634_),
    .C(_06601_),
    .Y(_06635_));
 sg13g2_a21oi_1 _14813_ (.A1(_06635_),
    .A2(_06610_),
    .Y(_06636_),
    .B1(_06617_));
 sg13g2_o21ai_1 _14814_ (.B1(_06636_),
    .Y(_06637_),
    .A1(_06610_),
    .A2(_06633_));
 sg13g2_nand3_1 _14815_ (.B(net206),
    .C(_06618_),
    .A(_06637_),
    .Y(_06638_));
 sg13g2_o21ai_1 _14816_ (.B1(_06638_),
    .Y(_00880_),
    .A1(_06114_),
    .A2(net206));
 sg13g2_a21oi_1 _14817_ (.A1(_06627_),
    .A2(_06611_),
    .Y(_06639_),
    .B1(_06617_));
 sg13g2_o21ai_1 _14818_ (.B1(_06639_),
    .Y(_06640_),
    .A1(_06611_),
    .A2(_06626_));
 sg13g2_a21oi_1 _14819_ (.A1(_06617_),
    .A2(_06587_),
    .Y(_06641_),
    .B1(_06504_));
 sg13g2_nand2_1 _14820_ (.Y(_06642_),
    .A(_06640_),
    .B(_06641_));
 sg13g2_o21ai_1 _14821_ (.B1(_06642_),
    .Y(_00881_),
    .A1(_06122_),
    .A2(net206));
 sg13g2_inv_1 _14822_ (.Y(_06643_),
    .A(\ppu.pixel_out_t[3] ));
 sg13g2_a21oi_1 _14823_ (.A1(_06635_),
    .A2(_06611_),
    .Y(_06644_),
    .B1(_06617_));
 sg13g2_o21ai_1 _14824_ (.B1(_06644_),
    .Y(_06645_),
    .A1(_06611_),
    .A2(_06633_));
 sg13g2_a21oi_1 _14825_ (.A1(_06617_),
    .A2(_06593_),
    .Y(_06646_),
    .B1(net264));
 sg13g2_nand2_1 _14826_ (.Y(_06647_),
    .A(_06645_),
    .B(_06646_));
 sg13g2_o21ai_1 _14827_ (.B1(_06647_),
    .Y(_00882_),
    .A1(_06643_),
    .A2(_06501_));
 sg13g2_nand2_1 _14828_ (.Y(_06648_),
    .A(_03401_),
    .B(_03400_));
 sg13g2_nor2_1 _14829_ (.A(_03403_),
    .B(_06648_),
    .Y(_06649_));
 sg13g2_nand2_1 _14830_ (.Y(_06650_),
    .A(_03586_),
    .B(_06649_));
 sg13g2_nor2_1 _14831_ (.A(_01789_),
    .B(_06650_),
    .Y(_06651_));
 sg13g2_xnor2_1 _14832_ (.Y(_06652_),
    .A(\synth.controller.read_index_reg[0] ),
    .B(_06651_));
 sg13g2_inv_2 _14833_ (.Y(_06653_),
    .A(\synth.voice.coeff_index[4] ));
 sg13g2_o21ai_1 _14834_ (.B1(_01720_),
    .Y(_06654_),
    .A1(_00049_),
    .A2(_06653_));
 sg13g2_buf_8 _14835_ (.A(_06654_),
    .X(_06655_));
 sg13g2_xnor2_1 _14836_ (.Y(_06656_),
    .A(_05760_),
    .B(_06655_));
 sg13g2_xnor2_1 _14837_ (.Y(_06657_),
    .A(_04908_),
    .B(_06655_));
 sg13g2_nand2_2 _14838_ (.Y(_06658_),
    .A(_06656_),
    .B(_06657_));
 sg13g2_inv_1 _14839_ (.Y(_06659_),
    .A(\synth.voice.coeff_index[3] ));
 sg13g2_xnor2_1 _14840_ (.Y(_06660_),
    .A(_06659_),
    .B(_06655_));
 sg13g2_xnor2_1 _14841_ (.Y(_06661_),
    .A(_05809_),
    .B(_06655_));
 sg13g2_nor2b_1 _14842_ (.A(_06660_),
    .B_N(_06661_),
    .Y(_06662_));
 sg13g2_buf_2 _14843_ (.A(_06662_),
    .X(_06663_));
 sg13g2_inv_2 _14844_ (.Y(_06664_),
    .A(_06663_));
 sg13g2_nor2_1 _14845_ (.A(_06658_),
    .B(_06664_),
    .Y(_06665_));
 sg13g2_inv_1 _14846_ (.Y(_06666_),
    .A(_00049_));
 sg13g2_inv_1 _14847_ (.Y(_06667_),
    .A(_00050_));
 sg13g2_xnor2_1 _14848_ (.Y(_06668_),
    .A(_06667_),
    .B(_06655_));
 sg13g2_inv_2 _14849_ (.Y(_06669_),
    .A(_06668_));
 sg13g2_nor2_1 _14850_ (.A(_06666_),
    .B(_06669_),
    .Y(_06670_));
 sg13g2_buf_2 _14851_ (.A(_06670_),
    .X(_06671_));
 sg13g2_nand2_1 _14852_ (.Y(_06672_),
    .A(_06665_),
    .B(_06671_));
 sg13g2_nor2_2 _14853_ (.A(_06660_),
    .B(_06661_),
    .Y(_06673_));
 sg13g2_inv_4 _14854_ (.A(_06673_),
    .Y(_06674_));
 sg13g2_inv_4 _14855_ (.A(_06656_),
    .Y(_06675_));
 sg13g2_nor2_1 _14856_ (.A(_06657_),
    .B(_06675_),
    .Y(_06676_));
 sg13g2_inv_2 _14857_ (.Y(_06677_),
    .A(_06676_));
 sg13g2_nor2_1 _14858_ (.A(_06674_),
    .B(_06677_),
    .Y(_06678_));
 sg13g2_nand2_1 _14859_ (.Y(_06679_),
    .A(_06678_),
    .B(_06671_));
 sg13g2_inv_1 _14860_ (.Y(_06680_),
    .A(_06660_));
 sg13g2_nor2_2 _14861_ (.A(_06661_),
    .B(_06680_),
    .Y(_06681_));
 sg13g2_inv_4 _14862_ (.A(_06681_),
    .Y(_06682_));
 sg13g2_nor2_1 _14863_ (.A(_06675_),
    .B(_06682_),
    .Y(_06683_));
 sg13g2_nand2_1 _14864_ (.Y(_06684_),
    .A(_06683_),
    .B(_06671_));
 sg13g2_nand3_1 _14865_ (.B(_06679_),
    .C(_06684_),
    .A(_06672_),
    .Y(_06685_));
 sg13g2_nand2_2 _14866_ (.Y(_06686_),
    .A(_06660_),
    .B(_06661_));
 sg13g2_xor2_1 _14867_ (.B(_06655_),
    .A(_04908_),
    .X(_06687_));
 sg13g2_nand2_2 _14868_ (.Y(_06688_),
    .A(_06675_),
    .B(_06687_));
 sg13g2_nor2_1 _14869_ (.A(_06686_),
    .B(_06688_),
    .Y(_06689_));
 sg13g2_nand2_1 _14870_ (.Y(_06690_),
    .A(_06689_),
    .B(_06671_));
 sg13g2_nor2_2 _14871_ (.A(_06686_),
    .B(_06658_),
    .Y(_06691_));
 sg13g2_nand2_2 _14872_ (.Y(_06692_),
    .A(_06691_),
    .B(_06671_));
 sg13g2_nand2_1 _14873_ (.Y(_06693_),
    .A(_06690_),
    .B(_06692_));
 sg13g2_nor2_2 _14874_ (.A(_06656_),
    .B(_06687_),
    .Y(_06694_));
 sg13g2_inv_4 _14875_ (.A(_06694_),
    .Y(_06695_));
 sg13g2_nor2_1 _14876_ (.A(_06674_),
    .B(_06695_),
    .Y(_06696_));
 sg13g2_buf_1 _14877_ (.A(_06671_),
    .X(_06697_));
 sg13g2_nand2_1 _14878_ (.Y(_06698_),
    .A(_06696_),
    .B(net205));
 sg13g2_nor2_1 _14879_ (.A(_06658_),
    .B(_06674_),
    .Y(_06699_));
 sg13g2_nand2_1 _14880_ (.Y(_06700_),
    .A(_06699_),
    .B(net205));
 sg13g2_nand2_1 _14881_ (.Y(_06701_),
    .A(_06669_),
    .B(_01750_));
 sg13g2_buf_1 _14882_ (.A(_06701_),
    .X(_06702_));
 sg13g2_inv_2 _14883_ (.Y(_06703_),
    .A(net219));
 sg13g2_nand2_2 _14884_ (.Y(_06704_),
    .A(_06691_),
    .B(net204));
 sg13g2_nand3_1 _14885_ (.B(_06700_),
    .C(_06704_),
    .A(_06698_),
    .Y(_06705_));
 sg13g2_nor2_1 _14886_ (.A(_01750_),
    .B(_06669_),
    .Y(_06706_));
 sg13g2_nand3_1 _14887_ (.B(_06706_),
    .C(_06656_),
    .A(_06663_),
    .Y(_06707_));
 sg13g2_nor2_1 _14888_ (.A(_06687_),
    .B(_06707_),
    .Y(_06708_));
 sg13g2_nor2_1 _14889_ (.A(_06658_),
    .B(_06682_),
    .Y(_06709_));
 sg13g2_buf_1 _14890_ (.A(_06706_),
    .X(_06710_));
 sg13g2_nand2_1 _14891_ (.Y(_06711_),
    .A(_06709_),
    .B(net218));
 sg13g2_inv_4 _14892_ (.A(_06688_),
    .Y(_06712_));
 sg13g2_nand3_1 _14893_ (.B(_06663_),
    .C(net218),
    .A(_06712_),
    .Y(_06713_));
 sg13g2_nand2_1 _14894_ (.Y(_06714_),
    .A(_06711_),
    .B(_06713_));
 sg13g2_nor2_1 _14895_ (.A(_06708_),
    .B(_06714_),
    .Y(_06715_));
 sg13g2_nor3_1 _14896_ (.A(net219),
    .B(_06695_),
    .C(_06682_),
    .Y(_06716_));
 sg13g2_nor3_2 _14897_ (.A(_06675_),
    .B(net219),
    .C(_06664_),
    .Y(_06717_));
 sg13g2_nor2_1 _14898_ (.A(_06716_),
    .B(_06717_),
    .Y(_06718_));
 sg13g2_nand2_1 _14899_ (.Y(_06719_),
    .A(_06715_),
    .B(_06718_));
 sg13g2_nor4_2 _14900_ (.A(_06685_),
    .B(_06693_),
    .C(_06705_),
    .Y(_06720_),
    .D(_06719_));
 sg13g2_nor2_1 _14901_ (.A(_06686_),
    .B(_06677_),
    .Y(_06721_));
 sg13g2_nand2_1 _14902_ (.Y(_06722_),
    .A(_06721_),
    .B(net205));
 sg13g2_nand2_1 _14903_ (.Y(_06723_),
    .A(_06696_),
    .B(net204));
 sg13g2_nand2_2 _14904_ (.Y(_06724_),
    .A(_06722_),
    .B(_06723_));
 sg13g2_nor2_1 _14905_ (.A(_06688_),
    .B(_06682_),
    .Y(_06725_));
 sg13g2_nand2_1 _14906_ (.Y(_06726_),
    .A(_06725_),
    .B(_06697_));
 sg13g2_inv_1 _14907_ (.Y(_06727_),
    .A(_06726_));
 sg13g2_inv_1 _14908_ (.Y(_06728_),
    .A(_06671_));
 sg13g2_nand2_1 _14909_ (.Y(_06729_),
    .A(_06712_),
    .B(_06663_));
 sg13g2_nor2_1 _14910_ (.A(_06728_),
    .B(_06729_),
    .Y(_06730_));
 sg13g2_nand2_1 _14911_ (.Y(_06731_),
    .A(_06663_),
    .B(_06676_));
 sg13g2_nor2_1 _14912_ (.A(_06728_),
    .B(_06731_),
    .Y(_06732_));
 sg13g2_nand2_1 _14913_ (.Y(_06733_),
    .A(_06712_),
    .B(_06673_));
 sg13g2_nor2_1 _14914_ (.A(_06728_),
    .B(_06733_),
    .Y(_06734_));
 sg13g2_nor2_1 _14915_ (.A(_06732_),
    .B(_06734_),
    .Y(_06735_));
 sg13g2_inv_1 _14916_ (.Y(_06736_),
    .A(_06731_));
 sg13g2_nand2_1 _14917_ (.Y(_06737_),
    .A(_06736_),
    .B(net218));
 sg13g2_nand2_1 _14918_ (.Y(_06738_),
    .A(_06735_),
    .B(_06737_));
 sg13g2_nor4_1 _14919_ (.A(_06724_),
    .B(_06727_),
    .C(_06730_),
    .D(_06738_),
    .Y(_06739_));
 sg13g2_a21oi_1 _14920_ (.A1(_06720_),
    .A2(_06739_),
    .Y(_06740_),
    .B1(_01716_));
 sg13g2_inv_1 _14921_ (.Y(_06741_),
    .A(_01716_));
 sg13g2_nand2_1 _14922_ (.Y(_06742_),
    .A(_06720_),
    .B(_06739_));
 sg13g2_nor2_1 _14923_ (.A(_06741_),
    .B(_06742_),
    .Y(_06743_));
 sg13g2_buf_2 _14924_ (.A(\synth.voice.fir_table.i_term[2] ),
    .X(_06744_));
 sg13g2_inv_2 _14925_ (.Y(_06745_),
    .A(net218));
 sg13g2_inv_2 _14926_ (.Y(_06746_),
    .A(_06699_));
 sg13g2_nor2_1 _14927_ (.A(_06745_),
    .B(_06746_),
    .Y(_06747_));
 sg13g2_nor3_1 _14928_ (.A(_06745_),
    .B(_06674_),
    .C(_06677_),
    .Y(_06748_));
 sg13g2_nor2_1 _14929_ (.A(_06747_),
    .B(_06748_),
    .Y(_06749_));
 sg13g2_inv_1 _14930_ (.Y(_06750_),
    .A(_06749_));
 sg13g2_nor2_1 _14931_ (.A(net219),
    .B(_06733_),
    .Y(_06751_));
 sg13g2_nor2_1 _14932_ (.A(net219),
    .B(_06729_),
    .Y(_06752_));
 sg13g2_nor2_1 _14933_ (.A(net219),
    .B(_06746_),
    .Y(_06753_));
 sg13g2_nor3_1 _14934_ (.A(_06751_),
    .B(_06752_),
    .C(_06753_),
    .Y(_06754_));
 sg13g2_nand2_1 _14935_ (.Y(_06755_),
    .A(_06663_),
    .B(_06694_));
 sg13g2_inv_1 _14936_ (.Y(_06756_),
    .A(_06755_));
 sg13g2_o21ai_1 _14937_ (.B1(net204),
    .Y(_06757_),
    .A1(_06678_),
    .A2(_06756_));
 sg13g2_buf_1 _14938_ (.A(_06757_),
    .X(_06758_));
 sg13g2_nand2_1 _14939_ (.Y(_06759_),
    .A(_06754_),
    .B(_06758_));
 sg13g2_nor2_1 _14940_ (.A(_06750_),
    .B(_06759_),
    .Y(_06760_));
 sg13g2_nand2_1 _14941_ (.Y(_06761_),
    .A(_06696_),
    .B(_06710_));
 sg13g2_nand2_1 _14942_ (.Y(_06762_),
    .A(_06689_),
    .B(net204));
 sg13g2_nand2_1 _14943_ (.Y(_06763_),
    .A(_06761_),
    .B(_06762_));
 sg13g2_nand2_1 _14944_ (.Y(_06764_),
    .A(_06676_),
    .B(_06681_));
 sg13g2_nor2_1 _14945_ (.A(_06745_),
    .B(_06764_),
    .Y(_06765_));
 sg13g2_nor2_1 _14946_ (.A(_06745_),
    .B(_06755_),
    .Y(_06766_));
 sg13g2_nor2_1 _14947_ (.A(_06765_),
    .B(_06766_),
    .Y(_06767_));
 sg13g2_nand2_1 _14948_ (.Y(_06768_),
    .A(_06725_),
    .B(_06710_));
 sg13g2_nor2_1 _14949_ (.A(_06695_),
    .B(_06682_),
    .Y(_06769_));
 sg13g2_nand2_1 _14950_ (.Y(_06770_),
    .A(_06769_),
    .B(net218));
 sg13g2_nand3_1 _14951_ (.B(_06768_),
    .C(_06770_),
    .A(_06767_),
    .Y(_06771_));
 sg13g2_nor2_1 _14952_ (.A(_06763_),
    .B(_06771_),
    .Y(_06772_));
 sg13g2_nand2_1 _14953_ (.Y(_06773_),
    .A(_06769_),
    .B(net205));
 sg13g2_nor2_1 _14954_ (.A(_06686_),
    .B(_06695_),
    .Y(_06774_));
 sg13g2_nand2_1 _14955_ (.Y(_06775_),
    .A(_06774_),
    .B(net205));
 sg13g2_nand2_1 _14956_ (.Y(_06776_),
    .A(_06773_),
    .B(_06775_));
 sg13g2_nand2_1 _14957_ (.Y(_06777_),
    .A(_06725_),
    .B(net204));
 sg13g2_nand2_1 _14958_ (.Y(_06778_),
    .A(_06683_),
    .B(net204));
 sg13g2_nand2_1 _14959_ (.Y(_06779_),
    .A(_06777_),
    .B(_06778_));
 sg13g2_nand2_1 _14960_ (.Y(_06780_),
    .A(_06774_),
    .B(net218));
 sg13g2_nand2_1 _14961_ (.Y(_06781_),
    .A(_06689_),
    .B(net218));
 sg13g2_nand2_1 _14962_ (.Y(_06782_),
    .A(_06691_),
    .B(net218));
 sg13g2_nand3_1 _14963_ (.B(_06781_),
    .C(_06782_),
    .A(_06780_),
    .Y(_06783_));
 sg13g2_nor3_1 _14964_ (.A(_06776_),
    .B(_06779_),
    .C(_06783_),
    .Y(_06784_));
 sg13g2_nor2_1 _14965_ (.A(_06745_),
    .B(_06733_),
    .Y(_06785_));
 sg13g2_inv_1 _14966_ (.Y(_06786_),
    .A(_06785_));
 sg13g2_nand2_1 _14967_ (.Y(_06787_),
    .A(_06721_),
    .B(net204));
 sg13g2_nand2_1 _14968_ (.Y(_06788_),
    .A(_06786_),
    .B(_06787_));
 sg13g2_inv_1 _14969_ (.Y(_06789_),
    .A(_06721_));
 sg13g2_nor2_1 _14970_ (.A(_06745_),
    .B(_06789_),
    .Y(_06790_));
 sg13g2_inv_1 _14971_ (.Y(_06791_),
    .A(_06790_));
 sg13g2_nand2_1 _14972_ (.Y(_06792_),
    .A(_06774_),
    .B(net204));
 sg13g2_nand2_1 _14973_ (.Y(_06793_),
    .A(_06791_),
    .B(_06792_));
 sg13g2_nor2_1 _14974_ (.A(_06788_),
    .B(_06793_),
    .Y(_06794_));
 sg13g2_nand4_1 _14975_ (.B(_06772_),
    .C(_06784_),
    .A(_06760_),
    .Y(_06795_),
    .D(_06794_));
 sg13g2_nor2b_1 _14976_ (.A(_06744_),
    .B_N(_06795_),
    .Y(_06796_));
 sg13g2_inv_1 _14977_ (.Y(_06797_),
    .A(_06744_));
 sg13g2_o21ai_1 _14978_ (.B1(_01732_),
    .Y(_06798_),
    .A1(_06797_),
    .A2(_06795_));
 sg13g2_nor4_2 _14979_ (.A(_06740_),
    .B(_06743_),
    .C(_06796_),
    .Y(_06799_),
    .D(_06798_));
 sg13g2_and2_1 _14980_ (.A(_06720_),
    .B(_06794_),
    .X(_06800_));
 sg13g2_o21ai_1 _14981_ (.B1(_06800_),
    .Y(_06801_),
    .A1(_06742_),
    .A2(_06795_));
 sg13g2_xor2_1 _14982_ (.B(_06801_),
    .A(_00048_),
    .X(_06802_));
 sg13g2_nand2_2 _14983_ (.Y(_06803_),
    .A(_06799_),
    .B(_06802_));
 sg13g2_o21ai_1 _14984_ (.B1(_01732_),
    .Y(_06804_),
    .A1(_01722_),
    .A2(_06803_));
 sg13g2_inv_1 _14985_ (.Y(_06805_),
    .A(_03432_));
 sg13g2_nand2_1 _14986_ (.Y(_06806_),
    .A(_06805_),
    .B(_03429_));
 sg13g2_nand2_1 _14987_ (.Y(_06807_),
    .A(_06804_),
    .B(_06806_));
 sg13g2_inv_1 _14988_ (.Y(_06808_),
    .A(\synth.controller.write_index_reg[0] ));
 sg13g2_nor2_1 _14989_ (.A(_03376_),
    .B(_03600_),
    .Y(_06809_));
 sg13g2_inv_1 _14990_ (.Y(_06810_),
    .A(_06809_));
 sg13g2_nor2_1 _14991_ (.A(_06808_),
    .B(_06810_),
    .Y(_06811_));
 sg13g2_nand2_1 _14992_ (.Y(_06812_),
    .A(_06811_),
    .B(_03596_));
 sg13g2_nor3_2 _14993_ (.A(_03430_),
    .B(_01725_),
    .C(_01756_),
    .Y(_06813_));
 sg13g2_o21ai_1 _14994_ (.B1(_06813_),
    .Y(_06814_),
    .A1(_04716_),
    .A2(_06812_));
 sg13g2_nor2b_1 _14995_ (.A(_06807_),
    .B_N(_06814_),
    .Y(_06815_));
 sg13g2_buf_2 _14996_ (.A(_06815_),
    .X(_06816_));
 sg13g2_nand2_1 _14997_ (.Y(_06817_),
    .A(_06816_),
    .B(_03443_));
 sg13g2_nor2_1 _14998_ (.A(_01789_),
    .B(_06817_),
    .Y(_06818_));
 sg13g2_buf_2 _14999_ (.A(_06818_),
    .X(_06819_));
 sg13g2_nor2_1 _15000_ (.A(_06652_),
    .B(_06819_),
    .Y(_00910_));
 sg13g2_nor4_2 _15001_ (.A(_01789_),
    .B(_00057_),
    .C(_04027_),
    .Y(_06820_),
    .D(_06650_));
 sg13g2_a21oi_1 _15002_ (.A1(_06651_),
    .A2(_03592_),
    .Y(_06821_),
    .B1(_03591_));
 sg13g2_nor3_1 _15003_ (.A(_06820_),
    .B(_06821_),
    .C(_06819_),
    .Y(_00911_));
 sg13g2_nand2_1 _15004_ (.Y(_06822_),
    .A(_06820_),
    .B(\synth.controller.read_index_reg[2] ));
 sg13g2_inv_1 _15005_ (.Y(_06823_),
    .A(_06822_));
 sg13g2_nor2_1 _15006_ (.A(\synth.controller.read_index_reg[2] ),
    .B(_06820_),
    .Y(_06824_));
 sg13g2_nor3_1 _15007_ (.A(_06823_),
    .B(_06824_),
    .C(_06819_),
    .Y(_00912_));
 sg13g2_xor2_1 _15008_ (.B(_06822_),
    .A(\synth.controller.read_index_reg[3] ),
    .X(_06825_));
 sg13g2_nor2_1 _15009_ (.A(_06825_),
    .B(_06819_),
    .Y(_00913_));
 sg13g2_buf_1 _15010_ (.A(net402),
    .X(_06826_));
 sg13g2_buf_1 _15011_ (.A(net402),
    .X(_06827_));
 sg13g2_nand2_1 _15012_ (.Y(_06828_),
    .A(_06827_),
    .B(_03765_));
 sg13g2_o21ai_1 _15013_ (.B1(_06828_),
    .Y(_00914_),
    .A1(_06826_),
    .A2(_05873_));
 sg13g2_nand2_1 _15014_ (.Y(_06829_),
    .A(net353),
    .B(_03930_));
 sg13g2_o21ai_1 _15015_ (.B1(_06829_),
    .Y(_00915_),
    .A1(net354),
    .A2(_04168_));
 sg13g2_nand2_1 _15016_ (.Y(_06830_),
    .A(net353),
    .B(\synth.controller.reg_waddr[3] ));
 sg13g2_o21ai_1 _15017_ (.B1(_06830_),
    .Y(_00916_),
    .A1(net354),
    .A2(_04188_));
 sg13g2_buf_1 _15018_ (.A(net402),
    .X(_06831_));
 sg13g2_nand2_1 _15019_ (.Y(_06832_),
    .A(net352),
    .B(\synth.controller.rx_buffer[12] ));
 sg13g2_o21ai_1 _15020_ (.B1(_06832_),
    .Y(_00917_),
    .A1(net354),
    .A2(_04074_));
 sg13g2_nor2_1 _15021_ (.A(net402),
    .B(\synth.controller.rx_buffer[15] ),
    .Y(_06833_));
 sg13g2_a21oi_1 _15022_ (.A1(net354),
    .A2(_04188_),
    .Y(_00918_),
    .B1(_06833_));
 sg13g2_nand2_1 _15023_ (.Y(_06834_),
    .A(net352),
    .B(net328));
 sg13g2_o21ai_1 _15024_ (.B1(_06834_),
    .Y(_00919_),
    .A1(net354),
    .A2(_03371_));
 sg13g2_nand2_1 _15025_ (.Y(_06835_),
    .A(net352),
    .B(\synth.controller.rx_buffer[15] ));
 sg13g2_o21ai_1 _15026_ (.B1(_06835_),
    .Y(_00920_),
    .A1(net354),
    .A2(_03383_));
 sg13g2_nand2_1 _15027_ (.Y(_06836_),
    .A(net352),
    .B(\synth.controller.reg_wdata[1] ));
 sg13g2_o21ai_1 _15028_ (.B1(_06836_),
    .Y(_00921_),
    .A1(net354),
    .A2(_03782_));
 sg13g2_nand2_1 _15029_ (.Y(_06837_),
    .A(net352),
    .B(_03750_));
 sg13g2_o21ai_1 _15030_ (.B1(_06837_),
    .Y(_00922_),
    .A1(net354),
    .A2(_03806_));
 sg13g2_nand2_1 _15031_ (.Y(_06838_),
    .A(net352),
    .B(\synth.controller.reg_wdata[3] ));
 sg13g2_o21ai_1 _15032_ (.B1(_06838_),
    .Y(_00923_),
    .A1(net353),
    .A2(_04062_));
 sg13g2_nand2_1 _15033_ (.Y(_06839_),
    .A(net352),
    .B(\synth.controller.reg_wdata[4] ));
 sg13g2_o21ai_1 _15034_ (.B1(_06839_),
    .Y(_00924_),
    .A1(net353),
    .A2(_03947_));
 sg13g2_nand2_1 _15035_ (.Y(_06840_),
    .A(net352),
    .B(\synth.controller.reg_wdata[5] ));
 sg13g2_o21ai_1 _15036_ (.B1(_06840_),
    .Y(_00925_),
    .A1(net353),
    .A2(_03978_));
 sg13g2_nand2_1 _15037_ (.Y(_06841_),
    .A(_06831_),
    .B(net374));
 sg13g2_o21ai_1 _15038_ (.B1(_06841_),
    .Y(_00926_),
    .A1(_06827_),
    .A2(_03960_));
 sg13g2_nand2_1 _15039_ (.Y(_06842_),
    .A(_06831_),
    .B(_03956_));
 sg13g2_o21ai_1 _15040_ (.B1(_06842_),
    .Y(_00927_),
    .A1(net353),
    .A2(_04007_));
 sg13g2_nand2_1 _15041_ (.Y(_06843_),
    .A(net402),
    .B(_03959_));
 sg13g2_o21ai_1 _15042_ (.B1(_06843_),
    .Y(_00928_),
    .A1(net353),
    .A2(_03933_));
 sg13g2_nand2_1 _15043_ (.Y(_06844_),
    .A(net402),
    .B(_03945_));
 sg13g2_o21ai_1 _15044_ (.B1(_06844_),
    .Y(_00929_),
    .A1(net353),
    .A2(_04149_));
 sg13g2_buf_1 _15045_ (.A(_01798_),
    .X(_06845_));
 sg13g2_buf_1 _15046_ (.A(_06845_),
    .X(_06846_));
 sg13g2_xnor2_1 _15047_ (.Y(_06847_),
    .A(_00111_),
    .B(_06809_));
 sg13g2_nand3_1 _15048_ (.B(net319),
    .C(_06847_),
    .A(_06817_),
    .Y(_06848_));
 sg13g2_o21ai_1 _15049_ (.B1(_06848_),
    .Y(_00961_),
    .A1(net290),
    .A2(_06808_));
 sg13g2_a21oi_1 _15050_ (.A1(_06811_),
    .A2(net319),
    .Y(_06849_),
    .B1(_03596_));
 sg13g2_nor2_1 _15051_ (.A(_01789_),
    .B(_06812_),
    .Y(_06850_));
 sg13g2_nor3_1 _15052_ (.A(_06849_),
    .B(_06850_),
    .C(_06819_),
    .Y(_00962_));
 sg13g2_nor3_1 _15053_ (.A(_01789_),
    .B(_04022_),
    .C(_06812_),
    .Y(_06851_));
 sg13g2_nor2_1 _15054_ (.A(_03604_),
    .B(_06850_),
    .Y(_06852_));
 sg13g2_nor3_1 _15055_ (.A(_06851_),
    .B(_06852_),
    .C(_06819_),
    .Y(_00963_));
 sg13g2_xnor2_1 _15056_ (.Y(_06853_),
    .A(\synth.controller.write_index_reg[3] ),
    .B(_06851_));
 sg13g2_nor2_1 _15057_ (.A(_06853_),
    .B(_06819_),
    .Y(_00964_));
 sg13g2_buf_1 _15058_ (.A(_04358_),
    .X(_06854_));
 sg13g2_mux2_1 _15059_ (.A0(\synth.voice.genblk4[8].next_state_scan[6] ),
    .A1(\synth.voice.genblk4[8].next_state_scan[8] ),
    .S(net147),
    .X(_01138_));
 sg13g2_mux2_1 _15060_ (.A0(\synth.voice.genblk4[8].next_state_scan[7] ),
    .A1(\synth.voice.genblk4[8].next_state_scan[9] ),
    .S(net147),
    .X(_01139_));
 sg13g2_mux2_1 _15061_ (.A0(\synth.voice.genblk4[8].next_state_scan[8] ),
    .A1(\synth.voice.genblk4[8].next_state_scan[10] ),
    .S(net147),
    .X(_01140_));
 sg13g2_mux2_1 _15062_ (.A0(\synth.voice.genblk4[8].next_state_scan[9] ),
    .A1(\synth.voice.genblk4[8].next_state_scan[11] ),
    .S(_06854_),
    .X(_01141_));
 sg13g2_mux2_1 _15063_ (.A0(\synth.voice.genblk4[8].next_state_scan[10] ),
    .A1(\synth.voice.genblk4[8].next_state_scan[12] ),
    .S(net147),
    .X(_01143_));
 sg13g2_mux2_1 _15064_ (.A0(\synth.voice.genblk4[8].next_state_scan[11] ),
    .A1(\synth.voice.genblk4[8].next_state_scan[13] ),
    .S(_06854_),
    .X(_01144_));
 sg13g2_nor2_1 _15065_ (.A(\synth.voice.genblk4[8].next_state_scan[12] ),
    .B(net147),
    .Y(_06855_));
 sg13g2_a21oi_1 _15066_ (.A1(net377),
    .A2(net147),
    .Y(_01145_),
    .B1(_06855_));
 sg13g2_nor2_1 _15067_ (.A(\synth.voice.genblk4[8].next_state_scan[13] ),
    .B(net147),
    .Y(_06856_));
 sg13g2_a21oi_1 _15068_ (.A1(_03383_),
    .A2(net147),
    .Y(_01146_),
    .B1(_06856_));
 sg13g2_inv_1 _15069_ (.Y(_06857_),
    .A(_02579_));
 sg13g2_nor4_2 _15070_ (.A(net297),
    .B(_02586_),
    .C(_06857_),
    .Y(_06858_),
    .D(_02602_));
 sg13g2_xor2_1 _15071_ (.B(_06858_),
    .A(_00131_),
    .X(_06859_));
 sg13g2_nand2_1 _15072_ (.Y(_06860_),
    .A(_02461_),
    .B(_02452_));
 sg13g2_o21ai_1 _15073_ (.B1(_02270_),
    .Y(_06861_),
    .A1(\ppu.copper_inst.cmp[1] ),
    .A2(_06860_));
 sg13g2_a21oi_1 _15074_ (.A1(_06859_),
    .A2(_06860_),
    .Y(_00217_),
    .B1(_06861_));
 sg13g2_inv_1 _15075_ (.Y(_06862_),
    .A(_06860_));
 sg13g2_buf_1 _15076_ (.A(_06862_),
    .X(_06863_));
 sg13g2_buf_1 _15077_ (.A(\ppu.copper_inst.addr[10] ),
    .X(_06864_));
 sg13g2_nand2_2 _15078_ (.Y(_06865_),
    .A(_06858_),
    .B(\ppu.copper_inst.addr[0] ));
 sg13g2_nor2_2 _15079_ (.A(_00132_),
    .B(_06865_),
    .Y(_06866_));
 sg13g2_inv_1 _15080_ (.Y(_06867_),
    .A(\ppu.copper_inst.addr[6] ));
 sg13g2_inv_1 _15081_ (.Y(_06868_),
    .A(\ppu.copper_inst.addr[7] ));
 sg13g2_inv_1 _15082_ (.Y(_06869_),
    .A(\ppu.copper_inst.addr[8] ));
 sg13g2_inv_1 _15083_ (.Y(_06870_),
    .A(\ppu.copper_inst.addr[9] ));
 sg13g2_nor4_1 _15084_ (.A(_06867_),
    .B(_06868_),
    .C(_06869_),
    .D(_06870_),
    .Y(_06871_));
 sg13g2_buf_1 _15085_ (.A(\ppu.copper_inst.addr[2] ),
    .X(_06872_));
 sg13g2_inv_1 _15086_ (.Y(_06873_),
    .A(_06872_));
 sg13g2_buf_1 _15087_ (.A(\ppu.copper_inst.addr[3] ),
    .X(_06874_));
 sg13g2_inv_1 _15088_ (.Y(_06875_),
    .A(_06874_));
 sg13g2_inv_1 _15089_ (.Y(_06876_),
    .A(\ppu.copper_inst.addr[4] ));
 sg13g2_inv_1 _15090_ (.Y(_06877_),
    .A(\ppu.copper_inst.addr[5] ));
 sg13g2_nor4_2 _15091_ (.A(_06873_),
    .B(_06875_),
    .C(_06876_),
    .Y(_06878_),
    .D(_06877_));
 sg13g2_nand3_1 _15092_ (.B(_06871_),
    .C(_06878_),
    .A(_06866_),
    .Y(_06879_));
 sg13g2_xor2_1 _15093_ (.B(_06879_),
    .A(_06864_),
    .X(_06880_));
 sg13g2_buf_1 _15094_ (.A(_06862_),
    .X(_06881_));
 sg13g2_inv_2 _15095_ (.Y(_06882_),
    .A(_02270_));
 sg13g2_buf_1 _15096_ (.A(_06882_),
    .X(_06883_));
 sg13g2_a21oi_1 _15097_ (.A1(net95),
    .A2(_02400_),
    .Y(_06884_),
    .B1(net68));
 sg13g2_o21ai_1 _15098_ (.B1(_06884_),
    .Y(_00218_),
    .A1(_06863_),
    .A2(_06880_));
 sg13g2_inv_1 _15099_ (.Y(_06885_),
    .A(\ppu.copper_inst.addr[11] ));
 sg13g2_nand2_1 _15100_ (.Y(_06886_),
    .A(\ppu.copper_inst.addr[1] ),
    .B(_06872_));
 sg13g2_nor2_2 _15101_ (.A(_06886_),
    .B(_06865_),
    .Y(_06887_));
 sg13g2_nand2_1 _15102_ (.Y(_06888_),
    .A(_06874_),
    .B(\ppu.copper_inst.addr[4] ));
 sg13g2_nand2_1 _15103_ (.Y(_06889_),
    .A(\ppu.copper_inst.addr[9] ),
    .B(_06864_));
 sg13g2_nand2_1 _15104_ (.Y(_06890_),
    .A(\ppu.copper_inst.addr[7] ),
    .B(\ppu.copper_inst.addr[8] ));
 sg13g2_nand2_1 _15105_ (.Y(_06891_),
    .A(\ppu.copper_inst.addr[5] ),
    .B(\ppu.copper_inst.addr[6] ));
 sg13g2_nor4_1 _15106_ (.A(_06888_),
    .B(_06889_),
    .C(_06890_),
    .D(_06891_),
    .Y(_06892_));
 sg13g2_nand2_1 _15107_ (.Y(_06893_),
    .A(_06887_),
    .B(_06892_));
 sg13g2_xnor2_1 _15108_ (.Y(_06894_),
    .A(_06885_),
    .B(_06893_));
 sg13g2_a21oi_1 _15109_ (.A1(net95),
    .A2(_02404_),
    .Y(_06895_),
    .B1(net68));
 sg13g2_o21ai_1 _15110_ (.B1(_06895_),
    .Y(_00219_),
    .A1(_06863_),
    .A2(_06894_));
 sg13g2_inv_1 _15111_ (.Y(_06896_),
    .A(\ppu.copper_inst.addr[12] ));
 sg13g2_nand3_1 _15112_ (.B(_06872_),
    .C(_06874_),
    .A(_06866_),
    .Y(_06897_));
 sg13g2_inv_1 _15113_ (.Y(_06898_),
    .A(_06897_));
 sg13g2_nand2_1 _15114_ (.Y(_06899_),
    .A(_06864_),
    .B(\ppu.copper_inst.addr[11] ));
 sg13g2_nor3_1 _15115_ (.A(_06869_),
    .B(_06870_),
    .C(_06899_),
    .Y(_06900_));
 sg13g2_nor4_1 _15116_ (.A(_06876_),
    .B(_06877_),
    .C(_06867_),
    .D(_06868_),
    .Y(_06901_));
 sg13g2_nand3_1 _15117_ (.B(_06900_),
    .C(_06901_),
    .A(_06898_),
    .Y(_06902_));
 sg13g2_xnor2_1 _15118_ (.Y(_06903_),
    .A(_06896_),
    .B(_06902_));
 sg13g2_a21oi_1 _15119_ (.A1(net95),
    .A2(_02408_),
    .Y(_06904_),
    .B1(net68));
 sg13g2_o21ai_1 _15120_ (.B1(_06904_),
    .Y(_00220_),
    .A1(net96),
    .A2(_06903_));
 sg13g2_inv_1 _15121_ (.Y(_06905_),
    .A(\ppu.copper_inst.addr[13] ));
 sg13g2_inv_1 _15122_ (.Y(_06906_),
    .A(_06865_));
 sg13g2_nor2_1 _15123_ (.A(_06888_),
    .B(_06886_),
    .Y(_06907_));
 sg13g2_nand2_1 _15124_ (.Y(_06908_),
    .A(\ppu.copper_inst.addr[11] ),
    .B(\ppu.copper_inst.addr[12] ));
 sg13g2_nor2_1 _15125_ (.A(_06889_),
    .B(_06908_),
    .Y(_06909_));
 sg13g2_nor2_1 _15126_ (.A(_06890_),
    .B(_06891_),
    .Y(_06910_));
 sg13g2_nand4_1 _15127_ (.B(_06907_),
    .C(_06909_),
    .A(_06906_),
    .Y(_06911_),
    .D(_06910_));
 sg13g2_xnor2_1 _15128_ (.Y(_06912_),
    .A(_06905_),
    .B(_06911_));
 sg13g2_a21oi_1 _15129_ (.A1(net95),
    .A2(_02411_),
    .Y(_06913_),
    .B1(net68));
 sg13g2_o21ai_1 _15130_ (.B1(_06913_),
    .Y(_00221_),
    .A1(net96),
    .A2(_06912_));
 sg13g2_inv_1 _15131_ (.Y(_06914_),
    .A(\ppu.copper_inst.addr[14] ));
 sg13g2_nor3_1 _15132_ (.A(_06896_),
    .B(_06905_),
    .C(_06899_),
    .Y(_06915_));
 sg13g2_nand4_1 _15133_ (.B(_06871_),
    .C(_06878_),
    .A(_06866_),
    .Y(_06916_),
    .D(_06915_));
 sg13g2_xnor2_1 _15134_ (.Y(_06917_),
    .A(_06914_),
    .B(_06916_));
 sg13g2_a21oi_1 _15135_ (.A1(net95),
    .A2(_02414_),
    .Y(_06918_),
    .B1(net68));
 sg13g2_o21ai_1 _15136_ (.B1(_06918_),
    .Y(_00222_),
    .A1(net96),
    .A2(_06917_));
 sg13g2_nor2_1 _15137_ (.A(_06888_),
    .B(_06891_),
    .Y(_06919_));
 sg13g2_nand2_1 _15138_ (.Y(_06920_),
    .A(\ppu.copper_inst.addr[13] ),
    .B(\ppu.copper_inst.addr[14] ));
 sg13g2_nor4_1 _15139_ (.A(_06889_),
    .B(_06890_),
    .C(_06908_),
    .D(_06920_),
    .Y(_06921_));
 sg13g2_nand3_1 _15140_ (.B(_06919_),
    .C(_06921_),
    .A(_06887_),
    .Y(_06922_));
 sg13g2_xor2_1 _15141_ (.B(_06922_),
    .A(\ppu.copper_inst.addr[15] ),
    .X(_06923_));
 sg13g2_buf_1 _15142_ (.A(_06862_),
    .X(_06924_));
 sg13g2_a21oi_1 _15143_ (.A1(net94),
    .A2(_02417_),
    .Y(_06925_),
    .B1(net68));
 sg13g2_o21ai_1 _15144_ (.B1(_06925_),
    .Y(_00223_),
    .A1(net96),
    .A2(_06923_));
 sg13g2_xor2_1 _15145_ (.B(_06865_),
    .A(\ppu.copper_inst.addr[1] ),
    .X(_06926_));
 sg13g2_a21oi_1 _15146_ (.A1(net94),
    .A2(\ppu.copper_inst.cmp[2] ),
    .Y(_06927_),
    .B1(net68));
 sg13g2_o21ai_1 _15147_ (.B1(_06927_),
    .Y(_00224_),
    .A1(net96),
    .A2(_06926_));
 sg13g2_xnor2_1 _15148_ (.Y(_06928_),
    .A(_06872_),
    .B(_06866_));
 sg13g2_a21oi_1 _15149_ (.A1(net94),
    .A2(\ppu.copper_inst.cmp[3] ),
    .Y(_06929_),
    .B1(_06883_));
 sg13g2_o21ai_1 _15150_ (.B1(_06929_),
    .Y(_00225_),
    .A1(net96),
    .A2(_06928_));
 sg13g2_xnor2_1 _15151_ (.Y(_06930_),
    .A(_06874_),
    .B(_06887_));
 sg13g2_a21oi_1 _15152_ (.A1(_06924_),
    .A2(_02348_),
    .Y(_06931_),
    .B1(_06883_));
 sg13g2_o21ai_1 _15153_ (.B1(_06931_),
    .Y(_00226_),
    .A1(net96),
    .A2(_06930_));
 sg13g2_xnor2_1 _15154_ (.Y(_06932_),
    .A(_06876_),
    .B(_06897_));
 sg13g2_a21oi_1 _15155_ (.A1(net94),
    .A2(_02304_),
    .Y(_06933_),
    .B1(_06882_));
 sg13g2_o21ai_1 _15156_ (.B1(_06933_),
    .Y(_00227_),
    .A1(net96),
    .A2(_06932_));
 sg13g2_nand2_1 _15157_ (.Y(_06934_),
    .A(_06906_),
    .B(_06907_));
 sg13g2_xnor2_1 _15158_ (.Y(_06935_),
    .A(_06877_),
    .B(_06934_));
 sg13g2_a21oi_1 _15159_ (.A1(net94),
    .A2(\ppu.copper_inst.cmp[6] ),
    .Y(_06936_),
    .B1(_06882_));
 sg13g2_o21ai_1 _15160_ (.B1(_06936_),
    .Y(_00228_),
    .A1(net95),
    .A2(_06935_));
 sg13g2_nand2_1 _15161_ (.Y(_06937_),
    .A(_06866_),
    .B(_06878_));
 sg13g2_xnor2_1 _15162_ (.Y(_06938_),
    .A(_06867_),
    .B(_06937_));
 sg13g2_a21oi_1 _15163_ (.A1(net94),
    .A2(_02315_),
    .Y(_06939_),
    .B1(_06882_));
 sg13g2_o21ai_1 _15164_ (.B1(_06939_),
    .Y(_00229_),
    .A1(net95),
    .A2(_06938_));
 sg13g2_nand2_1 _15165_ (.Y(_06940_),
    .A(_06887_),
    .B(_06919_));
 sg13g2_xnor2_1 _15166_ (.Y(_06941_),
    .A(_06868_),
    .B(_06940_));
 sg13g2_a21oi_1 _15167_ (.A1(_06924_),
    .A2(\ppu.copper_inst.cmp[8] ),
    .Y(_06942_),
    .B1(_06882_));
 sg13g2_o21ai_1 _15168_ (.B1(_06942_),
    .Y(_00230_),
    .A1(net95),
    .A2(_06941_));
 sg13g2_nand2_1 _15169_ (.Y(_06943_),
    .A(_06898_),
    .B(_06901_));
 sg13g2_xnor2_1 _15170_ (.Y(_06944_),
    .A(_06869_),
    .B(_06943_));
 sg13g2_a21oi_1 _15171_ (.A1(net94),
    .A2(_02392_),
    .Y(_06945_),
    .B1(_06882_));
 sg13g2_o21ai_1 _15172_ (.B1(_06945_),
    .Y(_00231_),
    .A1(_06881_),
    .A2(_06944_));
 sg13g2_nand3_1 _15173_ (.B(_06907_),
    .C(_06910_),
    .A(_06906_),
    .Y(_06946_));
 sg13g2_xnor2_1 _15174_ (.Y(_06947_),
    .A(_06870_),
    .B(_06946_));
 sg13g2_a21oi_1 _15175_ (.A1(net94),
    .A2(_02396_),
    .Y(_06948_),
    .B1(_06882_));
 sg13g2_o21ai_1 _15176_ (.B1(_06948_),
    .Y(_00232_),
    .A1(_06881_),
    .A2(_06947_));
 sg13g2_a22oi_1 _15177_ (.Y(_06949_),
    .B1(_02382_),
    .B2(_02461_),
    .A2(_02379_),
    .A1(\ppu.copper_inst.cmp_on ));
 sg13g2_nor2_1 _15178_ (.A(net68),
    .B(_06949_),
    .Y(_00242_));
 sg13g2_nand2_1 _15179_ (.Y(_06950_),
    .A(\ppu.copper_inst.x_cmp[2] ),
    .B(_01836_));
 sg13g2_nand2_1 _15180_ (.Y(_06951_),
    .A(_02210_),
    .B(_01816_));
 sg13g2_nor3_1 _15181_ (.A(_01804_),
    .B(_06950_),
    .C(_06951_),
    .Y(_06952_));
 sg13g2_xnor2_1 _15182_ (.Y(_06953_),
    .A(_01830_),
    .B(_06952_));
 sg13g2_nand2_1 _15183_ (.Y(_00452_),
    .A(_02216_),
    .B(_06953_));
 sg13g2_nor2_1 _15184_ (.A(_06950_),
    .B(_02226_),
    .Y(_06954_));
 sg13g2_inv_1 _15185_ (.Y(_06955_),
    .A(_02549_));
 sg13g2_nand2_1 _15186_ (.Y(_06956_),
    .A(_06954_),
    .B(_06955_));
 sg13g2_xnor2_1 _15187_ (.Y(_06957_),
    .A(_01812_),
    .B(_06956_));
 sg13g2_nand2_1 _15188_ (.Y(_00453_),
    .A(_02216_),
    .B(_06957_));
 sg13g2_nor2_1 _15189_ (.A(_01844_),
    .B(_06951_),
    .Y(_06958_));
 sg13g2_nand3_1 _15190_ (.B(_01836_),
    .C(_02550_),
    .A(_06958_),
    .Y(_06959_));
 sg13g2_xor2_1 _15191_ (.B(_06959_),
    .A(_02075_),
    .X(_06960_));
 sg13g2_nor2_1 _15192_ (.A(_06960_),
    .B(_02217_),
    .Y(_00454_));
 sg13g2_nand4_1 _15193_ (.B(_01811_),
    .C(_02075_),
    .A(_06954_),
    .Y(_06961_),
    .D(_06955_));
 sg13g2_xor2_1 _15194_ (.B(_06961_),
    .A(_01827_),
    .X(_06962_));
 sg13g2_nor2_1 _15195_ (.A(_06962_),
    .B(_02217_),
    .Y(_00455_));
 sg13g2_buf_1 _15196_ (.A(net146),
    .X(_06963_));
 sg13g2_nor2_1 _15197_ (.A(_00178_),
    .B(_02876_),
    .Y(_06964_));
 sg13g2_xnor2_1 _15198_ (.Y(_06965_),
    .A(_02866_),
    .B(_06964_));
 sg13g2_nor2_1 _15199_ (.A(net123),
    .B(_06965_),
    .Y(_00600_));
 sg13g2_inv_1 _15200_ (.Y(_06966_),
    .A(\ppu.sprite_buffer.extra_sorted_addr_bits[1] ));
 sg13g2_o21ai_1 _15201_ (.B1(_01853_),
    .Y(_06967_),
    .A1(_06966_),
    .A2(_02878_));
 sg13g2_a21oi_1 _15202_ (.A1(_06966_),
    .A2(_02878_),
    .Y(_00601_),
    .B1(_06967_));
 sg13g2_inv_1 _15203_ (.Y(_06968_),
    .A(\ppu.sprite_buffer.extra_sorted_addr_bits[2] ));
 sg13g2_nand3_1 _15204_ (.B(\ppu.sprite_buffer.extra_sorted_addr_bits[1] ),
    .C(_02866_),
    .A(_06964_),
    .Y(_06969_));
 sg13g2_o21ai_1 _15205_ (.B1(_01853_),
    .Y(_06970_),
    .A1(_06968_),
    .A2(_06969_));
 sg13g2_a21oi_1 _15206_ (.A1(_06968_),
    .A2(_06969_),
    .Y(_00602_),
    .B1(_06970_));
 sg13g2_nand2_1 _15207_ (.Y(_06971_),
    .A(_02851_),
    .B(_01863_));
 sg13g2_inv_1 _15208_ (.Y(_06972_),
    .A(_06971_));
 sg13g2_a21oi_1 _15209_ (.A1(_02803_),
    .A2(_01863_),
    .Y(_06973_),
    .B1(_01871_));
 sg13g2_nor3_1 _15210_ (.A(_06972_),
    .B(_06973_),
    .C(_06963_),
    .Y(_00627_));
 sg13g2_nor2_1 _15211_ (.A(_01872_),
    .B(_06972_),
    .Y(_06974_));
 sg13g2_nor2_1 _15212_ (.A(_01873_),
    .B(_06971_),
    .Y(_06975_));
 sg13g2_nor3_1 _15213_ (.A(_06974_),
    .B(_06975_),
    .C(net123),
    .Y(_00628_));
 sg13g2_nand2_1 _15214_ (.Y(_06976_),
    .A(_02670_),
    .B(net254));
 sg13g2_xnor2_1 _15215_ (.Y(_06977_),
    .A(_02672_),
    .B(_06976_));
 sg13g2_nor2_1 _15216_ (.A(_06977_),
    .B(net123),
    .Y(_00629_));
 sg13g2_nor2_1 _15217_ (.A(_00061_),
    .B(_06976_),
    .Y(_06978_));
 sg13g2_nand2_1 _15218_ (.Y(_06979_),
    .A(_06978_),
    .B(_02566_));
 sg13g2_inv_1 _15219_ (.Y(_06980_),
    .A(_06979_));
 sg13g2_nor2_1 _15220_ (.A(_02566_),
    .B(_06978_),
    .Y(_06981_));
 sg13g2_nor3_1 _15221_ (.A(_06980_),
    .B(_06981_),
    .C(net146),
    .Y(_00630_));
 sg13g2_xor2_1 _15222_ (.B(_06979_),
    .A(_02568_),
    .X(_06982_));
 sg13g2_nor2_1 _15223_ (.A(_06982_),
    .B(net123),
    .Y(_00631_));
 sg13g2_nor2_1 _15224_ (.A(_01908_),
    .B(_01906_),
    .Y(_06983_));
 sg13g2_nor2_1 _15225_ (.A(\ppu.sprite_buffer.final_pixels_in ),
    .B(_01907_),
    .Y(_06984_));
 sg13g2_nor3_1 _15226_ (.A(_06983_),
    .B(_06984_),
    .C(net146),
    .Y(_00632_));
 sg13g2_nand2_1 _15227_ (.Y(_06985_),
    .A(_06983_),
    .B(_01909_));
 sg13g2_inv_1 _15228_ (.Y(_06986_),
    .A(_06985_));
 sg13g2_nor2_1 _15229_ (.A(_01909_),
    .B(_06983_),
    .Y(_06987_));
 sg13g2_nor3_1 _15230_ (.A(_06986_),
    .B(_06987_),
    .C(net146),
    .Y(_00633_));
 sg13g2_xnor2_1 _15231_ (.Y(_06988_),
    .A(_02157_),
    .B(_06985_));
 sg13g2_nor2_1 _15232_ (.A(_06988_),
    .B(net123),
    .Y(_00634_));
 sg13g2_buf_1 _15233_ (.A(_02883_),
    .X(_06989_));
 sg13g2_a21oi_1 _15234_ (.A1(net104),
    .A2(_02588_),
    .Y(_06990_),
    .B1(\ppu.sprite_buffer.oam_req_step ));
 sg13g2_nor3_1 _15235_ (.A(net146),
    .B(_06990_),
    .C(_06524_),
    .Y(_00636_));
 sg13g2_xor2_1 _15236_ (.B(_02871_),
    .A(\ppu.sprite_buffer.out_counters[0][0] ),
    .X(_06991_));
 sg13g2_nor2_1 _15237_ (.A(net123),
    .B(_06991_),
    .Y(_00637_));
 sg13g2_nor2_1 _15238_ (.A(_02873_),
    .B(_02872_),
    .Y(_06992_));
 sg13g2_nor3_1 _15239_ (.A(net146),
    .B(_06992_),
    .C(_02875_),
    .Y(_00638_));
 sg13g2_a21oi_1 _15240_ (.A1(_02876_),
    .A2(_00178_),
    .Y(_06993_),
    .B1(net146));
 sg13g2_nor2b_1 _15241_ (.A(_06964_),
    .B_N(_06993_),
    .Y(_00639_));
 sg13g2_nor2_1 _15242_ (.A(net123),
    .B(_06525_),
    .Y(_00640_));
 sg13g2_nor2_1 _15243_ (.A(net123),
    .B(_06528_),
    .Y(_00641_));
 sg13g2_nor2_1 _15244_ (.A(_02579_),
    .B(_02603_),
    .Y(_06994_));
 sg13g2_buf_2 _15245_ (.A(_06994_),
    .X(_06995_));
 sg13g2_buf_1 _15246_ (.A(_06995_),
    .X(_06996_));
 sg13g2_nand2_1 _15247_ (.Y(_06997_),
    .A(_06996_),
    .B(net254));
 sg13g2_xnor2_1 _15248_ (.Y(_06998_),
    .A(_00160_),
    .B(_06997_));
 sg13g2_nor2_1 _15249_ (.A(_06963_),
    .B(_06998_),
    .Y(_00642_));
 sg13g2_buf_1 _15250_ (.A(\ppu.sprite_buffer.out_counters[2][1] ),
    .X(_06999_));
 sg13g2_buf_1 _15251_ (.A(net395),
    .X(_07000_));
 sg13g2_nor2b_1 _15252_ (.A(_06997_),
    .B_N(\ppu.sprite_buffer.out_counters[2][0] ),
    .Y(_07001_));
 sg13g2_nor2_1 _15253_ (.A(net351),
    .B(_07001_),
    .Y(_07002_));
 sg13g2_nand2_1 _15254_ (.Y(_07003_),
    .A(_07001_),
    .B(net351));
 sg13g2_inv_1 _15255_ (.Y(_07004_),
    .A(_07003_));
 sg13g2_nor3_1 _15256_ (.A(_01913_),
    .B(_07002_),
    .C(_07004_),
    .Y(_00643_));
 sg13g2_nor2b_1 _15257_ (.A(_07003_),
    .B_N(\ppu.sprite_buffer.out_counters[2][2] ),
    .Y(_07005_));
 sg13g2_nor2_1 _15258_ (.A(\ppu.sprite_buffer.out_counters[2][2] ),
    .B(_07004_),
    .Y(_07006_));
 sg13g2_nor3_1 _15259_ (.A(_01913_),
    .B(_07005_),
    .C(_07006_),
    .Y(_00644_));
 sg13g2_a22oi_1 _15260_ (.Y(_07007_),
    .B1(_02069_),
    .B2(_02079_),
    .A2(_02068_),
    .A1(_01827_));
 sg13g2_nand2_1 _15261_ (.Y(_07008_),
    .A(_02092_),
    .B(_02277_));
 sg13g2_nor2_1 _15262_ (.A(_07007_),
    .B(_07008_),
    .Y(_07009_));
 sg13g2_a21o_1 _15263_ (.A2(net216),
    .A1(_07009_),
    .B1(_06531_),
    .X(_07010_));
 sg13g2_nor2_1 _15264_ (.A(_02207_),
    .B(_01853_),
    .Y(_07011_));
 sg13g2_a21oi_1 _15265_ (.A1(_07010_),
    .A2(_02178_),
    .Y(_00817_),
    .B1(_07011_));
 sg13g2_nand2_1 _15266_ (.Y(_07012_),
    .A(_07009_),
    .B(net235));
 sg13g2_nand2_1 _15267_ (.Y(_07013_),
    .A(_07012_),
    .B(\ppu.sprite_buffer.valid_sprites[1] ));
 sg13g2_a21oi_1 _15268_ (.A1(_07013_),
    .A2(_02159_),
    .Y(_00818_),
    .B1(_07011_));
 sg13g2_a21o_1 _15269_ (.A2(net251),
    .A1(_07009_),
    .B1(_06526_),
    .X(_07014_));
 sg13g2_inv_1 _15270_ (.Y(_07015_),
    .A(_02143_));
 sg13g2_a21oi_1 _15271_ (.A1(_07014_),
    .A2(_07015_),
    .Y(_00819_),
    .B1(_07011_));
 sg13g2_nand2_1 _15272_ (.Y(_07016_),
    .A(_07009_),
    .B(_02234_));
 sg13g2_a21oi_1 _15273_ (.A1(_07016_),
    .A2(\ppu.sprite_buffer.valid_sprites[3] ),
    .Y(_07017_),
    .B1(_01911_));
 sg13g2_nor2_1 _15274_ (.A(_07011_),
    .B(_07017_),
    .Y(_00820_));
 sg13g2_inv_1 _15275_ (.Y(_07018_),
    .A(_06813_));
 sg13g2_nor3_1 _15276_ (.A(_04716_),
    .B(_07018_),
    .C(_06812_),
    .Y(_07019_));
 sg13g2_nand3_1 _15277_ (.B(_06806_),
    .C(_07019_),
    .A(_06804_),
    .Y(_07020_));
 sg13g2_buf_2 _15278_ (.A(_07020_),
    .X(_07021_));
 sg13g2_nand2_1 _15279_ (.Y(_07022_),
    .A(_01736_),
    .B(_03412_));
 sg13g2_xor2_1 _15280_ (.B(_07022_),
    .A(_00052_),
    .X(_07023_));
 sg13g2_nand3_1 _15281_ (.B(\synth.voice.coeff_index[2] ),
    .C(_07023_),
    .A(_05762_),
    .Y(_07024_));
 sg13g2_o21ai_1 _15282_ (.B1(_07024_),
    .Y(_07025_),
    .A1(_06659_),
    .A2(_07022_));
 sg13g2_nand2_1 _15283_ (.Y(_07026_),
    .A(_07025_),
    .B(_06667_));
 sg13g2_o21ai_1 _15284_ (.B1(_01736_),
    .Y(_07027_),
    .A1(_01792_),
    .A2(_07026_));
 sg13g2_nand2_1 _15285_ (.Y(_07028_),
    .A(_07021_),
    .B(_07027_));
 sg13g2_buf_8 _15286_ (.A(_06816_),
    .X(_07029_));
 sg13g2_nand2_1 _15287_ (.Y(_07030_),
    .A(net67),
    .B(_01754_));
 sg13g2_inv_1 _15288_ (.Y(_07031_),
    .A(_07029_));
 sg13g2_a21oi_1 _15289_ (.A1(_07031_),
    .A2(_01727_),
    .Y(_07032_),
    .B1(net394));
 sg13g2_o21ai_1 _15290_ (.B1(_07032_),
    .Y(_00883_),
    .A1(_07028_),
    .A2(_07030_));
 sg13g2_nor2_1 _15291_ (.A(_01776_),
    .B(_07031_),
    .Y(_07033_));
 sg13g2_nand2_1 _15292_ (.Y(_07034_),
    .A(_07028_),
    .B(net67));
 sg13g2_inv_1 _15293_ (.Y(_07035_),
    .A(_07034_));
 sg13g2_o21ai_1 _15294_ (.B1(_06845_),
    .Y(_07036_),
    .A1(_01728_),
    .A2(net67));
 sg13g2_nor3_1 _15295_ (.A(_07033_),
    .B(_07035_),
    .C(_07036_),
    .Y(_00884_));
 sg13g2_a21oi_1 _15296_ (.A1(net67),
    .A2(_01773_),
    .Y(_07037_),
    .B1(_01725_));
 sg13g2_nand3_1 _15297_ (.B(_01725_),
    .C(net299),
    .A(net67),
    .Y(_07038_));
 sg13g2_nand2_1 _15298_ (.Y(_07039_),
    .A(_07038_),
    .B(_07034_));
 sg13g2_o21ai_1 _15299_ (.B1(net290),
    .Y(_00885_),
    .A1(_07037_),
    .A2(_07039_));
 sg13g2_nor3_1 _15300_ (.A(_00150_),
    .B(_01742_),
    .C(_01734_),
    .Y(_07040_));
 sg13g2_nand2_1 _15301_ (.Y(_07041_),
    .A(net67),
    .B(_07040_));
 sg13g2_xnor2_1 _15302_ (.Y(_07042_),
    .A(_03430_),
    .B(_07041_));
 sg13g2_nor3_1 _15303_ (.A(net394),
    .B(_07035_),
    .C(_07042_),
    .Y(_00886_));
 sg13g2_nand2_1 _15304_ (.Y(_07043_),
    .A(_07029_),
    .B(_06813_));
 sg13g2_xnor2_1 _15305_ (.Y(_07044_),
    .A(_00146_),
    .B(_07043_));
 sg13g2_buf_1 _15306_ (.A(_01789_),
    .X(_07045_));
 sg13g2_a21oi_1 _15307_ (.A1(_07031_),
    .A2(\synth.controller.curr_voice[0] ),
    .Y(_07046_),
    .B1(net350));
 sg13g2_o21ai_1 _15308_ (.B1(_07046_),
    .Y(_00887_),
    .A1(_07031_),
    .A2(_07044_));
 sg13g2_inv_1 _15309_ (.Y(_07047_),
    .A(\synth.controller.curr_voice[1] ));
 sg13g2_nand4_1 _15310_ (.B(\synth.controller.curr_voice[0] ),
    .C(_06806_),
    .A(_06804_),
    .Y(_07048_),
    .D(_07019_));
 sg13g2_nor2_2 _15311_ (.A(_07047_),
    .B(_07048_),
    .Y(_07049_));
 sg13g2_inv_4 _15312_ (.A(_07049_),
    .Y(_07050_));
 sg13g2_nand2_1 _15313_ (.Y(_07051_),
    .A(_07048_),
    .B(_07047_));
 sg13g2_buf_1 _15314_ (.A(_07045_),
    .X(_07052_));
 sg13g2_a21o_1 _15315_ (.A2(_07051_),
    .A1(_07050_),
    .B1(net318),
    .X(_00888_));
 sg13g2_nand2_1 _15316_ (.Y(_07053_),
    .A(_06649_),
    .B(_03404_));
 sg13g2_o21ai_1 _15317_ (.B1(_03385_),
    .Y(_07054_),
    .A1(_03309_),
    .A2(_07053_));
 sg13g2_buf_1 _15318_ (.A(net350),
    .X(_07055_));
 sg13g2_a21oi_1 _15319_ (.A1(_07054_),
    .A2(_03319_),
    .Y(_00905_),
    .B1(_07055_));
 sg13g2_inv_1 _15320_ (.Y(_07056_),
    .A(\ppu_ctrl[0] ));
 sg13g2_nor2_1 _15321_ (.A(_03930_),
    .B(\synth.controller.reg_waddr[3] ),
    .Y(_07057_));
 sg13g2_inv_1 _15322_ (.Y(_07058_),
    .A(_07057_));
 sg13g2_nor3_1 _15323_ (.A(_03382_),
    .B(_03598_),
    .C(_04014_),
    .Y(_07059_));
 sg13g2_inv_1 _15324_ (.Y(_07060_),
    .A(_07059_));
 sg13g2_nor4_1 _15325_ (.A(_03959_),
    .B(_04007_),
    .C(_07058_),
    .D(_07060_),
    .Y(_07061_));
 sg13g2_buf_2 _15326_ (.A(_07061_),
    .X(_07062_));
 sg13g2_a21oi_1 _15327_ (.A1(_07062_),
    .A2(_03765_),
    .Y(_07063_),
    .B1(net350));
 sg13g2_o21ai_1 _15328_ (.B1(_07063_),
    .Y(_00906_),
    .A1(_07056_),
    .A2(_07062_));
 sg13g2_buf_1 _15329_ (.A(net319),
    .X(_07064_));
 sg13g2_o21ai_1 _15330_ (.B1(net289),
    .Y(_07065_),
    .A1(\ppu_ctrl[2] ),
    .A2(_07062_));
 sg13g2_a21oi_1 _15331_ (.A1(_05873_),
    .A2(_07062_),
    .Y(_00907_),
    .B1(_07065_));
 sg13g2_buf_2 _15332_ (.A(dither_out),
    .X(_07066_));
 sg13g2_inv_2 _15333_ (.Y(_07067_),
    .A(_07066_));
 sg13g2_a21oi_1 _15334_ (.A1(_07062_),
    .A2(\synth.controller.reg_wdata[3] ),
    .Y(_07068_),
    .B1(net350));
 sg13g2_o21ai_1 _15335_ (.B1(_07068_),
    .Y(_00908_),
    .A1(_07067_),
    .A2(_07062_));
 sg13g2_o21ai_1 _15336_ (.B1(_07064_),
    .Y(_07069_),
    .A1(\ppu_ctrl[4] ),
    .A2(_07062_));
 sg13g2_a21oi_1 _15337_ (.A1(_03806_),
    .A2(_07062_),
    .Y(_00909_),
    .B1(_07069_));
 sg13g2_nor3_1 _15338_ (.A(net394),
    .B(_06826_),
    .C(_03376_),
    .Y(_00930_));
 sg13g2_inv_1 _15339_ (.Y(_07070_),
    .A(_07026_));
 sg13g2_a21oi_1 _15340_ (.A1(net67),
    .A2(_07070_),
    .Y(_07071_),
    .B1(\synth.controller.sample_counter[0] ));
 sg13g2_and3_1 _15341_ (.X(_07072_),
    .A(net67),
    .B(\synth.controller.sample_counter[0] ),
    .C(_07070_));
 sg13g2_nor3_1 _15342_ (.A(net394),
    .B(_07071_),
    .C(_07072_),
    .Y(_00933_));
 sg13g2_xnor2_1 _15343_ (.Y(_07073_),
    .A(\synth.controller.sample_counter[1] ),
    .B(_07072_));
 sg13g2_nor2_1 _15344_ (.A(net317),
    .B(_07073_),
    .Y(_00934_));
 sg13g2_nor4_2 _15345_ (.A(_03959_),
    .B(_03945_),
    .C(_07058_),
    .Y(_07074_),
    .D(_07060_));
 sg13g2_nor2_1 _15346_ (.A(\synth.controller.sample_credits[0] ),
    .B(_03319_),
    .Y(_07075_));
 sg13g2_nor2b_1 _15347_ (.A(_03300_),
    .B_N(\synth.controller.sample_credits[0] ),
    .Y(_07076_));
 sg13g2_nor2_1 _15348_ (.A(_07075_),
    .B(_07076_),
    .Y(_07077_));
 sg13g2_a21oi_1 _15349_ (.A1(_07074_),
    .A2(_03765_),
    .Y(_07078_),
    .B1(_07045_));
 sg13g2_o21ai_1 _15350_ (.B1(_07078_),
    .Y(_00935_),
    .A1(_07074_),
    .A2(_07077_));
 sg13g2_xor2_1 _15351_ (.B(_07075_),
    .A(\synth.controller.sample_credits[1] ),
    .X(_07079_));
 sg13g2_o21ai_1 _15352_ (.B1(net289),
    .Y(_07080_),
    .A1(_07079_),
    .A2(_07074_));
 sg13g2_a21oi_1 _15353_ (.A1(_05865_),
    .A2(_07074_),
    .Y(_00936_),
    .B1(_07080_));
 sg13g2_inv_1 _15354_ (.Y(_07081_),
    .A(\synth.controller.sbio_credits[0] ));
 sg13g2_nor4_1 _15355_ (.A(_03960_),
    .B(_03945_),
    .C(_07058_),
    .D(_07060_),
    .Y(_07082_));
 sg13g2_buf_1 _15356_ (.A(_07082_),
    .X(_07083_));
 sg13g2_a21oi_1 _15357_ (.A1(_07083_),
    .A2(_03765_),
    .Y(_07084_),
    .B1(net350));
 sg13g2_o21ai_1 _15358_ (.B1(_07084_),
    .Y(_00937_),
    .A1(_07081_),
    .A2(_07083_));
 sg13g2_o21ai_1 _15359_ (.B1(net289),
    .Y(_07085_),
    .A1(\synth.controller.sbio_credits[1] ),
    .A2(_07083_));
 sg13g2_a21oi_1 _15360_ (.A1(_05865_),
    .A2(_07083_),
    .Y(_00938_),
    .B1(_07085_));
 sg13g2_o21ai_1 _15361_ (.B1(net289),
    .Y(_07086_),
    .A1(\synth.controller.sbio_credits[2] ),
    .A2(_07083_));
 sg13g2_a21oi_1 _15362_ (.A1(_05873_),
    .A2(_07083_),
    .Y(_00939_),
    .B1(_07086_));
 sg13g2_inv_1 _15363_ (.Y(_07087_),
    .A(_03376_));
 sg13g2_o21ai_1 _15364_ (.B1(_03372_),
    .Y(_07088_),
    .A1(_03370_),
    .A2(net401));
 sg13g2_a21oi_2 _15365_ (.B1(net350),
    .Y(_07089_),
    .A2(_07088_),
    .A1(_07087_));
 sg13g2_nand2b_1 _15366_ (.Y(_00940_),
    .B(_07089_),
    .A_N(_00181_));
 sg13g2_nor2_1 _15367_ (.A(\synth.controller.rx_counter[1] ),
    .B(\synth.controller.rx_counter[0] ),
    .Y(_07090_));
 sg13g2_o21ai_1 _15368_ (.B1(_07089_),
    .Y(_00941_),
    .A1(_03375_),
    .A2(_07090_));
 sg13g2_nor2_1 _15369_ (.A(\synth.controller.rx_counter[2] ),
    .B(_03375_),
    .Y(_07091_));
 sg13g2_o21ai_1 _15370_ (.B1(_07089_),
    .Y(_00942_),
    .A1(_07087_),
    .A2(_07091_));
 sg13g2_o21ai_1 _15371_ (.B1(_07089_),
    .Y(_00943_),
    .A1(_03373_),
    .A2(_07087_));
 sg13g2_inv_1 _15372_ (.Y(_07092_),
    .A(_07053_));
 sg13g2_inv_1 _15373_ (.Y(_07093_),
    .A(_03405_));
 sg13g2_nor2_1 _15374_ (.A(_07093_),
    .B(_03399_),
    .Y(_07094_));
 sg13g2_nor3_2 _15375_ (.A(net350),
    .B(_07092_),
    .C(_07094_),
    .Y(_07095_));
 sg13g2_and2_1 _15376_ (.A(_07095_),
    .B(_00182_),
    .X(_00944_));
 sg13g2_inv_1 _15377_ (.Y(_07096_),
    .A(_06648_));
 sg13g2_nor2_1 _15378_ (.A(_03401_),
    .B(_03400_),
    .Y(_07097_));
 sg13g2_o21ai_1 _15379_ (.B1(_07095_),
    .Y(_00945_),
    .A1(_07096_),
    .A2(_07097_));
 sg13g2_nor2_1 _15380_ (.A(\synth.controller.sbio_tx.counter[2] ),
    .B(_07096_),
    .Y(_07098_));
 sg13g2_o21ai_1 _15381_ (.B1(_07095_),
    .Y(_00946_),
    .A1(_06649_),
    .A2(_07098_));
 sg13g2_o21ai_1 _15382_ (.B1(_07095_),
    .Y(_00947_),
    .A1(_03404_),
    .A2(_06649_));
 sg13g2_nand3_1 _15383_ (.B(_03591_),
    .C(\synth.controller.read_index_reg[0] ),
    .A(_04351_),
    .Y(_07099_));
 sg13g2_o21ai_1 _15384_ (.B1(\synth.controller.scanning_out ),
    .Y(_07100_),
    .A1(_06650_),
    .A2(_07099_));
 sg13g2_a21oi_1 _15385_ (.A1(_06817_),
    .A2(_07100_),
    .Y(_00948_),
    .B1(_07055_));
 sg13g2_o21ai_1 _15386_ (.B1(_07035_),
    .Y(_07101_),
    .A1(_06805_),
    .A2(_07070_));
 sg13g2_a21oi_1 _15387_ (.A1(_07034_),
    .A2(\synth.controller.step_sample ),
    .Y(_07102_),
    .B1(net394));
 sg13g2_nand2_1 _15388_ (.Y(_00949_),
    .A(_07101_),
    .B(_07102_));
 sg13g2_nor2_1 _15389_ (.A(_03306_),
    .B(_03408_),
    .Y(_07103_));
 sg13g2_nand2_1 _15390_ (.Y(_07104_),
    .A(_07092_),
    .B(_07103_));
 sg13g2_nand2_1 _15391_ (.Y(_07105_),
    .A(_07104_),
    .B(_00149_));
 sg13g2_nor2_1 _15392_ (.A(_00149_),
    .B(_07104_),
    .Y(_07106_));
 sg13g2_inv_1 _15393_ (.Y(_07107_),
    .A(_07106_));
 sg13g2_nand3_1 _15394_ (.B(_07105_),
    .C(_07107_),
    .A(_07021_),
    .Y(_07108_));
 sg13g2_nand2_1 _15395_ (.Y(_00950_),
    .A(_07108_),
    .B(_06846_));
 sg13g2_nor2_1 _15396_ (.A(_03393_),
    .B(_07107_),
    .Y(_07109_));
 sg13g2_nor2_1 _15397_ (.A(\synth.controller.sweep_addr_index[1] ),
    .B(_07106_),
    .Y(_07110_));
 sg13g2_nand2_1 _15398_ (.Y(_07111_),
    .A(_07021_),
    .B(_00080_));
 sg13g2_nor3_1 _15399_ (.A(_07109_),
    .B(_07110_),
    .C(_07111_),
    .Y(_00951_));
 sg13g2_xor2_1 _15400_ (.B(_07109_),
    .A(\synth.controller.sweep_addr_index[2] ),
    .X(_07112_));
 sg13g2_a21o_1 _15401_ (.A2(_07112_),
    .A1(_07021_),
    .B1(net318),
    .X(_00952_));
 sg13g2_nand2b_1 _15402_ (.Y(_07113_),
    .B(_00148_),
    .A_N(_04016_));
 sg13g2_nor2b_1 _15403_ (.A(_00148_),
    .B_N(_04016_),
    .Y(_07114_));
 sg13g2_inv_1 _15404_ (.Y(_07115_),
    .A(_07114_));
 sg13g2_nand3_1 _15405_ (.B(_07113_),
    .C(_07115_),
    .A(_07021_),
    .Y(_07116_));
 sg13g2_nand2_1 _15406_ (.Y(_00953_),
    .A(_07116_),
    .B(net290));
 sg13g2_xnor2_1 _15407_ (.Y(_07117_),
    .A(_03423_),
    .B(_07114_));
 sg13g2_nor2_1 _15408_ (.A(_07117_),
    .B(_07111_),
    .Y(_00954_));
 sg13g2_nor2_1 _15409_ (.A(_00120_),
    .B(_07115_),
    .Y(_07118_));
 sg13g2_xnor2_1 _15410_ (.Y(_07119_),
    .A(_00051_),
    .B(_07118_));
 sg13g2_a21o_1 _15411_ (.A2(_07119_),
    .A1(_07021_),
    .B1(net318),
    .X(_00955_));
 sg13g2_o21ai_1 _15412_ (.B1(_03384_),
    .Y(_07120_),
    .A1(_03371_),
    .A2(_03383_));
 sg13g2_xor2_1 _15413_ (.B(_03407_),
    .A(_07120_),
    .X(_07121_));
 sg13g2_nor2_1 _15414_ (.A(_03388_),
    .B(_07121_),
    .Y(_07122_));
 sg13g2_inv_1 _15415_ (.Y(_07123_),
    .A(_07122_));
 sg13g2_nand2_1 _15416_ (.Y(_07124_),
    .A(_07123_),
    .B(_06846_));
 sg13g2_a21oi_1 _15417_ (.A1(_03388_),
    .A2(_07121_),
    .Y(_00956_),
    .B1(_07124_));
 sg13g2_nor3_1 _15418_ (.A(\synth.controller.tx_outstanding[1] ),
    .B(_07120_),
    .C(_03407_),
    .Y(_07125_));
 sg13g2_nor2_1 _15419_ (.A(_07120_),
    .B(_03407_),
    .Y(_07126_));
 sg13g2_nor2_1 _15420_ (.A(_03386_),
    .B(_07126_),
    .Y(_07127_));
 sg13g2_nor2_1 _15421_ (.A(_07125_),
    .B(_07127_),
    .Y(_07128_));
 sg13g2_o21ai_1 _15422_ (.B1(net289),
    .Y(_07129_),
    .A1(_07128_),
    .A2(_07123_));
 sg13g2_a21oi_1 _15423_ (.A1(_07123_),
    .A2(_07128_),
    .Y(_00957_),
    .B1(_07129_));
 sg13g2_inv_1 _15424_ (.Y(_07130_),
    .A(_07127_));
 sg13g2_nand2_1 _15425_ (.Y(_07131_),
    .A(_07125_),
    .B(_03388_));
 sg13g2_o21ai_1 _15426_ (.B1(_07131_),
    .Y(_07132_),
    .A1(_07130_),
    .A2(_07123_));
 sg13g2_o21ai_1 _15427_ (.B1(net289),
    .Y(_07133_),
    .A1(\synth.controller.tx_outstanding[2] ),
    .A2(_07132_));
 sg13g2_a21oi_1 _15428_ (.A1(\synth.controller.tx_outstanding[2] ),
    .A2(_07132_),
    .Y(_00958_),
    .B1(_07133_));
 sg13g2_buf_1 _15429_ (.A(\synth.voice.scan_accs_reg ),
    .X(_07134_));
 sg13g2_nor2b_1 _15430_ (.A(_07134_),
    .B_N(\synth.voice.target_reg[2] ),
    .Y(_07135_));
 sg13g2_buf_1 _15431_ (.A(_07135_),
    .X(_07136_));
 sg13g2_buf_1 _15432_ (.A(_07136_),
    .X(_07137_));
 sg13g2_nand2_1 _15433_ (.Y(_07138_),
    .A(_05524_),
    .B(_07137_));
 sg13g2_buf_1 _15434_ (.A(_07134_),
    .X(_07139_));
 sg13g2_buf_1 _15435_ (.A(_07139_),
    .X(_07140_));
 sg13g2_nor2_1 _15436_ (.A(\synth.voice.target_reg[2] ),
    .B(_07134_),
    .Y(_07141_));
 sg13g2_buf_1 _15437_ (.A(_07141_),
    .X(_07142_));
 sg13g2_a22oi_1 _15438_ (.Y(_07143_),
    .B1(\synth.voice.acc[0] ),
    .B2(net315),
    .A2(\synth.voice.accs[5][0] ),
    .A1(net316));
 sg13g2_a21oi_1 _15439_ (.A1(_07138_),
    .A2(_07143_),
    .Y(_00965_),
    .B1(net317));
 sg13g2_nand2_1 _15440_ (.Y(_07144_),
    .A(_05650_),
    .B(_07137_));
 sg13g2_a22oi_1 _15441_ (.Y(_07145_),
    .B1(\synth.controller.out[6] ),
    .B2(net315),
    .A2(\synth.voice.accs[5][10] ),
    .A1(net316));
 sg13g2_a21oi_1 _15442_ (.A1(_07144_),
    .A2(_07145_),
    .Y(_00966_),
    .B1(net317));
 sg13g2_nand2_1 _15443_ (.Y(_07146_),
    .A(_05657_),
    .B(net288));
 sg13g2_a22oi_1 _15444_ (.Y(_07147_),
    .B1(\synth.controller.out[7] ),
    .B2(net315),
    .A2(\synth.voice.accs[5][11] ),
    .A1(net316));
 sg13g2_a21oi_1 _15445_ (.A1(_07146_),
    .A2(_07147_),
    .Y(_00967_),
    .B1(net317));
 sg13g2_nand2_1 _15446_ (.Y(_07148_),
    .A(_05673_),
    .B(net288));
 sg13g2_a22oi_1 _15447_ (.Y(_07149_),
    .B1(_03364_),
    .B2(net315),
    .A2(\synth.voice.accs[5][12] ),
    .A1(net316));
 sg13g2_a21oi_1 _15448_ (.A1(_07148_),
    .A2(_07149_),
    .Y(_00968_),
    .B1(net317));
 sg13g2_nand2_1 _15449_ (.Y(_07150_),
    .A(_05686_),
    .B(net288));
 sg13g2_a22oi_1 _15450_ (.Y(_07151_),
    .B1(_03366_),
    .B2(net315),
    .A2(\synth.voice.accs[5][13] ),
    .A1(net316));
 sg13g2_a21oi_1 _15451_ (.A1(_07150_),
    .A2(_07151_),
    .Y(_00969_),
    .B1(net317));
 sg13g2_nand2_1 _15452_ (.Y(_07152_),
    .A(_05702_),
    .B(net288));
 sg13g2_a22oi_1 _15453_ (.Y(_07153_),
    .B1(_03316_),
    .B2(net315),
    .A2(\synth.voice.accs[5][14] ),
    .A1(net316));
 sg13g2_a21oi_1 _15454_ (.A1(_07152_),
    .A2(_07153_),
    .Y(_00970_),
    .B1(net317));
 sg13g2_nand2_1 _15455_ (.Y(_07154_),
    .A(_05712_),
    .B(net288));
 sg13g2_a22oi_1 _15456_ (.Y(_07155_),
    .B1(\synth.controller.out[11] ),
    .B2(net315),
    .A2(\synth.voice.accs[5][15] ),
    .A1(net316));
 sg13g2_a21oi_1 _15457_ (.A1(_07154_),
    .A2(_07155_),
    .Y(_00971_),
    .B1(net317));
 sg13g2_nand2_1 _15458_ (.Y(_07156_),
    .A(_05730_),
    .B(net288));
 sg13g2_buf_1 _15459_ (.A(_07139_),
    .X(_07157_));
 sg13g2_a22oi_1 _15460_ (.Y(_07158_),
    .B1(_03327_),
    .B2(net315),
    .A2(\synth.voice.accs[5][16] ),
    .A1(net314));
 sg13g2_buf_1 _15461_ (.A(net350),
    .X(_07159_));
 sg13g2_a21oi_1 _15462_ (.A1(_07156_),
    .A2(_07158_),
    .Y(_00972_),
    .B1(net313));
 sg13g2_nand2_1 _15463_ (.Y(_07160_),
    .A(_05754_),
    .B(net288));
 sg13g2_a22oi_1 _15464_ (.Y(_07161_),
    .B1(_03330_),
    .B2(_07142_),
    .A2(\synth.voice.accs[5][17] ),
    .A1(net314));
 sg13g2_a21oi_1 _15465_ (.A1(_07160_),
    .A2(_07161_),
    .Y(_00973_),
    .B1(net313));
 sg13g2_nand2_1 _15466_ (.Y(_07162_),
    .A(_05781_),
    .B(net288));
 sg13g2_a22oi_1 _15467_ (.Y(_07163_),
    .B1(\synth.controller.out[14] ),
    .B2(_07142_),
    .A2(\synth.voice.accs[5][18] ),
    .A1(net314));
 sg13g2_a21oi_1 _15468_ (.A1(_07162_),
    .A2(_07163_),
    .Y(_00974_),
    .B1(net313));
 sg13g2_buf_1 _15469_ (.A(_07136_),
    .X(_07164_));
 sg13g2_nand3_1 _15470_ (.B(_05519_),
    .C(net287),
    .A(_05784_),
    .Y(_07165_));
 sg13g2_buf_1 _15471_ (.A(_07141_),
    .X(_07166_));
 sg13g2_a22oi_1 _15472_ (.Y(_07167_),
    .B1(\synth.controller.out[15] ),
    .B2(net312),
    .A2(\synth.voice.accs[5][19] ),
    .A1(net314));
 sg13g2_a21oi_1 _15473_ (.A1(_07165_),
    .A2(_07167_),
    .Y(_00975_),
    .B1(net313));
 sg13g2_nand2_1 _15474_ (.Y(_07168_),
    .A(_05540_),
    .B(net287));
 sg13g2_a22oi_1 _15475_ (.Y(_07169_),
    .B1(\synth.voice.acc[1] ),
    .B2(net312),
    .A2(\synth.voice.accs[5][1] ),
    .A1(net314));
 sg13g2_a21oi_1 _15476_ (.A1(_07168_),
    .A2(_07169_),
    .Y(_00976_),
    .B1(net313));
 sg13g2_nand2_1 _15477_ (.Y(_07170_),
    .A(_05551_),
    .B(net287));
 sg13g2_a22oi_1 _15478_ (.Y(_07171_),
    .B1(\synth.voice.acc[2] ),
    .B2(net312),
    .A2(\synth.voice.accs[5][2] ),
    .A1(net314));
 sg13g2_a21oi_1 _15479_ (.A1(_07170_),
    .A2(_07171_),
    .Y(_00977_),
    .B1(net313));
 sg13g2_nand2_1 _15480_ (.Y(_07172_),
    .A(_05556_),
    .B(net287));
 sg13g2_a22oi_1 _15481_ (.Y(_07173_),
    .B1(\synth.voice.acc[3] ),
    .B2(net312),
    .A2(\synth.voice.accs[5][3] ),
    .A1(net314));
 sg13g2_a21oi_1 _15482_ (.A1(_07172_),
    .A2(_07173_),
    .Y(_00978_),
    .B1(net313));
 sg13g2_nand2_1 _15483_ (.Y(_07174_),
    .A(_05567_),
    .B(net287));
 sg13g2_a22oi_1 _15484_ (.Y(_07175_),
    .B1(\synth.controller.out[0] ),
    .B2(net312),
    .A2(\synth.voice.accs[5][4] ),
    .A1(net314));
 sg13g2_a21oi_1 _15485_ (.A1(_07174_),
    .A2(_07175_),
    .Y(_00979_),
    .B1(net313));
 sg13g2_nand2_1 _15486_ (.Y(_07176_),
    .A(_05574_),
    .B(_07164_));
 sg13g2_a22oi_1 _15487_ (.Y(_07177_),
    .B1(\synth.controller.out[1] ),
    .B2(_07166_),
    .A2(\synth.voice.accs[5][5] ),
    .A1(_07157_));
 sg13g2_a21oi_1 _15488_ (.A1(_07176_),
    .A2(_07177_),
    .Y(_00980_),
    .B1(_07159_));
 sg13g2_nand2_1 _15489_ (.Y(_07178_),
    .A(_05587_),
    .B(_07164_));
 sg13g2_a22oi_1 _15490_ (.Y(_07179_),
    .B1(\synth.controller.out[2] ),
    .B2(_07166_),
    .A2(\synth.voice.accs[5][6] ),
    .A1(_07157_));
 sg13g2_a21oi_1 _15491_ (.A1(_07178_),
    .A2(_07179_),
    .Y(_00981_),
    .B1(_07159_));
 sg13g2_nand2_1 _15492_ (.Y(_07180_),
    .A(_05595_),
    .B(net287));
 sg13g2_buf_1 _15493_ (.A(_07134_),
    .X(_07181_));
 sg13g2_a22oi_1 _15494_ (.Y(_07182_),
    .B1(\synth.controller.out[3] ),
    .B2(net312),
    .A2(\synth.voice.accs[5][7] ),
    .A1(net349));
 sg13g2_a21oi_1 _15495_ (.A1(_07180_),
    .A2(_07182_),
    .Y(_00982_),
    .B1(net318));
 sg13g2_nand2_1 _15496_ (.Y(_07183_),
    .A(_05619_),
    .B(net287));
 sg13g2_a22oi_1 _15497_ (.Y(_07184_),
    .B1(\synth.controller.out[4] ),
    .B2(net312),
    .A2(\synth.voice.accs[5][8] ),
    .A1(net349));
 sg13g2_a21oi_1 _15498_ (.A1(_07183_),
    .A2(_07184_),
    .Y(_00983_),
    .B1(net318));
 sg13g2_nand2_1 _15499_ (.Y(_07185_),
    .A(_05635_),
    .B(net287));
 sg13g2_a22oi_1 _15500_ (.Y(_07186_),
    .B1(\synth.controller.out[5] ),
    .B2(net312),
    .A2(\synth.voice.accs[5][9] ),
    .A1(net349));
 sg13g2_a21oi_1 _15501_ (.A1(_07185_),
    .A2(_07186_),
    .Y(_00984_),
    .B1(net318));
 sg13g2_buf_1 _15502_ (.A(_07139_),
    .X(_07187_));
 sg13g2_buf_1 _15503_ (.A(_07187_),
    .X(_07188_));
 sg13g2_inv_1 _15504_ (.Y(_07189_),
    .A(\synth.voice.acc[0] ));
 sg13g2_buf_1 _15505_ (.A(net349),
    .X(_07190_));
 sg13g2_buf_1 _15506_ (.A(net319),
    .X(_07191_));
 sg13g2_o21ai_1 _15507_ (.B1(_07191_),
    .Y(_07192_),
    .A1(_07190_),
    .A2(\synth.voice.accs[1][0] ));
 sg13g2_a21oi_1 _15508_ (.A1(net286),
    .A2(_07189_),
    .Y(_00985_),
    .B1(_07192_));
 sg13g2_inv_1 _15509_ (.Y(_07193_),
    .A(\synth.controller.out[6] ));
 sg13g2_o21ai_1 _15510_ (.B1(net285),
    .Y(_07194_),
    .A1(net311),
    .A2(\synth.voice.accs[1][10] ));
 sg13g2_a21oi_1 _15511_ (.A1(net286),
    .A2(_07193_),
    .Y(_00986_),
    .B1(_07194_));
 sg13g2_inv_1 _15512_ (.Y(_07195_),
    .A(\synth.controller.out[7] ));
 sg13g2_o21ai_1 _15513_ (.B1(net285),
    .Y(_07196_),
    .A1(net311),
    .A2(\synth.voice.accs[1][11] ));
 sg13g2_a21oi_1 _15514_ (.A1(_07188_),
    .A2(_07195_),
    .Y(_00987_),
    .B1(_07196_));
 sg13g2_inv_1 _15515_ (.Y(_07197_),
    .A(_03364_));
 sg13g2_o21ai_1 _15516_ (.B1(net285),
    .Y(_07198_),
    .A1(net311),
    .A2(\synth.voice.accs[1][12] ));
 sg13g2_a21oi_1 _15517_ (.A1(net286),
    .A2(_07197_),
    .Y(_00988_),
    .B1(_07198_));
 sg13g2_inv_1 _15518_ (.Y(_07199_),
    .A(_03366_));
 sg13g2_o21ai_1 _15519_ (.B1(net285),
    .Y(_07200_),
    .A1(net311),
    .A2(\synth.voice.accs[1][13] ));
 sg13g2_a21oi_1 _15520_ (.A1(net286),
    .A2(_07199_),
    .Y(_00989_),
    .B1(_07200_));
 sg13g2_inv_1 _15521_ (.Y(_07201_),
    .A(_03316_));
 sg13g2_o21ai_1 _15522_ (.B1(net285),
    .Y(_07202_),
    .A1(net311),
    .A2(\synth.voice.accs[1][14] ));
 sg13g2_a21oi_1 _15523_ (.A1(net286),
    .A2(_07201_),
    .Y(_00990_),
    .B1(_07202_));
 sg13g2_o21ai_1 _15524_ (.B1(net285),
    .Y(_07203_),
    .A1(net311),
    .A2(\synth.voice.accs[1][15] ));
 sg13g2_a21oi_1 _15525_ (.A1(net286),
    .A2(_03322_),
    .Y(_00991_),
    .B1(_07203_));
 sg13g2_inv_1 _15526_ (.Y(_07204_),
    .A(_03327_));
 sg13g2_o21ai_1 _15527_ (.B1(net285),
    .Y(_07205_),
    .A1(net311),
    .A2(\synth.voice.accs[1][16] ));
 sg13g2_a21oi_1 _15528_ (.A1(net286),
    .A2(_07204_),
    .Y(_00992_),
    .B1(_07205_));
 sg13g2_inv_1 _15529_ (.Y(_07206_),
    .A(_03330_));
 sg13g2_o21ai_1 _15530_ (.B1(_07191_),
    .Y(_07207_),
    .A1(_07190_),
    .A2(\synth.voice.accs[1][17] ));
 sg13g2_a21oi_1 _15531_ (.A1(_07188_),
    .A2(_07206_),
    .Y(_00993_),
    .B1(_07207_));
 sg13g2_o21ai_1 _15532_ (.B1(net285),
    .Y(_07208_),
    .A1(net311),
    .A2(\synth.voice.accs[1][18] ));
 sg13g2_a21oi_1 _15533_ (.A1(net286),
    .A2(_03333_),
    .Y(_00994_),
    .B1(_07208_));
 sg13g2_buf_1 _15534_ (.A(_07187_),
    .X(_07209_));
 sg13g2_buf_1 _15535_ (.A(_07181_),
    .X(_07210_));
 sg13g2_buf_1 _15536_ (.A(net319),
    .X(_07211_));
 sg13g2_o21ai_1 _15537_ (.B1(net283),
    .Y(_07212_),
    .A1(net310),
    .A2(\synth.voice.accs[1][19] ));
 sg13g2_a21oi_1 _15538_ (.A1(net284),
    .A2(_03335_),
    .Y(_00995_),
    .B1(_07212_));
 sg13g2_inv_1 _15539_ (.Y(_07213_),
    .A(\synth.voice.acc[1] ));
 sg13g2_o21ai_1 _15540_ (.B1(net283),
    .Y(_07214_),
    .A1(net310),
    .A2(\synth.voice.accs[1][1] ));
 sg13g2_a21oi_1 _15541_ (.A1(net284),
    .A2(_07213_),
    .Y(_00996_),
    .B1(_07214_));
 sg13g2_inv_1 _15542_ (.Y(_07215_),
    .A(\synth.voice.acc[2] ));
 sg13g2_o21ai_1 _15543_ (.B1(_07211_),
    .Y(_07216_),
    .A1(_07210_),
    .A2(\synth.voice.accs[1][2] ));
 sg13g2_a21oi_1 _15544_ (.A1(net284),
    .A2(_07215_),
    .Y(_00997_),
    .B1(_07216_));
 sg13g2_inv_1 _15545_ (.Y(_07217_),
    .A(\synth.voice.acc[3] ));
 sg13g2_o21ai_1 _15546_ (.B1(_07211_),
    .Y(_07218_),
    .A1(_07210_),
    .A2(\synth.voice.accs[1][3] ));
 sg13g2_a21oi_1 _15547_ (.A1(_07209_),
    .A2(_07217_),
    .Y(_00998_),
    .B1(_07218_));
 sg13g2_inv_1 _15548_ (.Y(_07219_),
    .A(\synth.controller.out[0] ));
 sg13g2_o21ai_1 _15549_ (.B1(net283),
    .Y(_07220_),
    .A1(net310),
    .A2(\synth.voice.accs[1][4] ));
 sg13g2_a21oi_1 _15550_ (.A1(net284),
    .A2(_07219_),
    .Y(_00999_),
    .B1(_07220_));
 sg13g2_inv_1 _15551_ (.Y(_07221_),
    .A(\synth.controller.out[1] ));
 sg13g2_o21ai_1 _15552_ (.B1(net283),
    .Y(_07222_),
    .A1(net310),
    .A2(\synth.voice.accs[1][5] ));
 sg13g2_a21oi_1 _15553_ (.A1(_07209_),
    .A2(_07221_),
    .Y(_01000_),
    .B1(_07222_));
 sg13g2_inv_1 _15554_ (.Y(_07223_),
    .A(\synth.controller.out[2] ));
 sg13g2_o21ai_1 _15555_ (.B1(net283),
    .Y(_07224_),
    .A1(net310),
    .A2(\synth.voice.accs[1][6] ));
 sg13g2_a21oi_1 _15556_ (.A1(net284),
    .A2(_07223_),
    .Y(_01001_),
    .B1(_07224_));
 sg13g2_inv_1 _15557_ (.Y(_07225_),
    .A(\synth.controller.out[3] ));
 sg13g2_o21ai_1 _15558_ (.B1(net283),
    .Y(_07226_),
    .A1(net310),
    .A2(\synth.voice.accs[1][7] ));
 sg13g2_a21oi_1 _15559_ (.A1(net284),
    .A2(_07225_),
    .Y(_01002_),
    .B1(_07226_));
 sg13g2_inv_1 _15560_ (.Y(_07227_),
    .A(\synth.controller.out[4] ));
 sg13g2_o21ai_1 _15561_ (.B1(net283),
    .Y(_07228_),
    .A1(net310),
    .A2(\synth.voice.accs[1][8] ));
 sg13g2_a21oi_1 _15562_ (.A1(net284),
    .A2(_07227_),
    .Y(_01003_),
    .B1(_07228_));
 sg13g2_inv_1 _15563_ (.Y(_07229_),
    .A(\synth.controller.out[5] ));
 sg13g2_o21ai_1 _15564_ (.B1(net283),
    .Y(_07230_),
    .A1(net310),
    .A2(\synth.voice.accs[1][9] ));
 sg13g2_a21oi_1 _15565_ (.A1(net284),
    .A2(_07229_),
    .Y(_01004_),
    .B1(_07230_));
 sg13g2_buf_1 _15566_ (.A(_07187_),
    .X(_07231_));
 sg13g2_inv_1 _15567_ (.Y(_07232_),
    .A(\synth.voice.accs[1][0] ));
 sg13g2_buf_1 _15568_ (.A(net349),
    .X(_07233_));
 sg13g2_buf_1 _15569_ (.A(net319),
    .X(_07234_));
 sg13g2_o21ai_1 _15570_ (.B1(net281),
    .Y(_07235_),
    .A1(net309),
    .A2(\synth.voice.accs[2][0] ));
 sg13g2_a21oi_1 _15571_ (.A1(net282),
    .A2(_07232_),
    .Y(_01005_),
    .B1(_07235_));
 sg13g2_inv_1 _15572_ (.Y(_07236_),
    .A(\synth.voice.accs[1][10] ));
 sg13g2_o21ai_1 _15573_ (.B1(net281),
    .Y(_07237_),
    .A1(net309),
    .A2(\synth.voice.accs[2][10] ));
 sg13g2_a21oi_1 _15574_ (.A1(net282),
    .A2(_07236_),
    .Y(_01006_),
    .B1(_07237_));
 sg13g2_inv_1 _15575_ (.Y(_07238_),
    .A(\synth.voice.accs[1][11] ));
 sg13g2_o21ai_1 _15576_ (.B1(net281),
    .Y(_07239_),
    .A1(net309),
    .A2(\synth.voice.accs[2][11] ));
 sg13g2_a21oi_1 _15577_ (.A1(net282),
    .A2(_07238_),
    .Y(_01007_),
    .B1(_07239_));
 sg13g2_inv_1 _15578_ (.Y(_07240_),
    .A(\synth.voice.accs[1][12] ));
 sg13g2_o21ai_1 _15579_ (.B1(net281),
    .Y(_07241_),
    .A1(net309),
    .A2(\synth.voice.accs[2][12] ));
 sg13g2_a21oi_1 _15580_ (.A1(net282),
    .A2(_07240_),
    .Y(_01008_),
    .B1(_07241_));
 sg13g2_inv_1 _15581_ (.Y(_07242_),
    .A(\synth.voice.accs[1][13] ));
 sg13g2_o21ai_1 _15582_ (.B1(net281),
    .Y(_07243_),
    .A1(net309),
    .A2(\synth.voice.accs[2][13] ));
 sg13g2_a21oi_1 _15583_ (.A1(net282),
    .A2(_07242_),
    .Y(_01009_),
    .B1(_07243_));
 sg13g2_inv_1 _15584_ (.Y(_07244_),
    .A(\synth.voice.accs[1][14] ));
 sg13g2_o21ai_1 _15585_ (.B1(net281),
    .Y(_07245_),
    .A1(net309),
    .A2(\synth.voice.accs[2][14] ));
 sg13g2_a21oi_1 _15586_ (.A1(net282),
    .A2(_07244_),
    .Y(_01010_),
    .B1(_07245_));
 sg13g2_inv_1 _15587_ (.Y(_07246_),
    .A(\synth.voice.accs[1][15] ));
 sg13g2_o21ai_1 _15588_ (.B1(_07234_),
    .Y(_07247_),
    .A1(_07233_),
    .A2(\synth.voice.accs[2][15] ));
 sg13g2_a21oi_1 _15589_ (.A1(_07231_),
    .A2(_07246_),
    .Y(_01011_),
    .B1(_07247_));
 sg13g2_inv_1 _15590_ (.Y(_07248_),
    .A(\synth.voice.accs[1][16] ));
 sg13g2_o21ai_1 _15591_ (.B1(net281),
    .Y(_07249_),
    .A1(net309),
    .A2(\synth.voice.accs[2][16] ));
 sg13g2_a21oi_1 _15592_ (.A1(net282),
    .A2(_07248_),
    .Y(_01012_),
    .B1(_07249_));
 sg13g2_inv_1 _15593_ (.Y(_07250_),
    .A(\synth.voice.accs[1][17] ));
 sg13g2_o21ai_1 _15594_ (.B1(net281),
    .Y(_07251_),
    .A1(net309),
    .A2(\synth.voice.accs[2][17] ));
 sg13g2_a21oi_1 _15595_ (.A1(net282),
    .A2(_07250_),
    .Y(_01013_),
    .B1(_07251_));
 sg13g2_inv_1 _15596_ (.Y(_07252_),
    .A(\synth.voice.accs[1][18] ));
 sg13g2_o21ai_1 _15597_ (.B1(_07234_),
    .Y(_07253_),
    .A1(_07233_),
    .A2(\synth.voice.accs[2][18] ));
 sg13g2_a21oi_1 _15598_ (.A1(_07231_),
    .A2(_07252_),
    .Y(_01014_),
    .B1(_07253_));
 sg13g2_buf_1 _15599_ (.A(_07187_),
    .X(_07254_));
 sg13g2_inv_1 _15600_ (.Y(_07255_),
    .A(\synth.voice.accs[1][19] ));
 sg13g2_buf_1 _15601_ (.A(net349),
    .X(_07256_));
 sg13g2_buf_1 _15602_ (.A(_01798_),
    .X(_07257_));
 sg13g2_buf_1 _15603_ (.A(_07257_),
    .X(_07258_));
 sg13g2_o21ai_1 _15604_ (.B1(net279),
    .Y(_07259_),
    .A1(net308),
    .A2(\synth.voice.accs[2][19] ));
 sg13g2_a21oi_1 _15605_ (.A1(net280),
    .A2(_07255_),
    .Y(_01015_),
    .B1(_07259_));
 sg13g2_inv_1 _15606_ (.Y(_07260_),
    .A(\synth.voice.accs[1][1] ));
 sg13g2_o21ai_1 _15607_ (.B1(net279),
    .Y(_07261_),
    .A1(net308),
    .A2(\synth.voice.accs[2][1] ));
 sg13g2_a21oi_1 _15608_ (.A1(_07254_),
    .A2(_07260_),
    .Y(_01016_),
    .B1(_07261_));
 sg13g2_inv_1 _15609_ (.Y(_07262_),
    .A(\synth.voice.accs[1][2] ));
 sg13g2_o21ai_1 _15610_ (.B1(_07258_),
    .Y(_07263_),
    .A1(_07256_),
    .A2(\synth.voice.accs[2][2] ));
 sg13g2_a21oi_1 _15611_ (.A1(_07254_),
    .A2(_07262_),
    .Y(_01017_),
    .B1(_07263_));
 sg13g2_inv_1 _15612_ (.Y(_07264_),
    .A(\synth.voice.accs[1][3] ));
 sg13g2_o21ai_1 _15613_ (.B1(net279),
    .Y(_07265_),
    .A1(net308),
    .A2(\synth.voice.accs[2][3] ));
 sg13g2_a21oi_1 _15614_ (.A1(net280),
    .A2(_07264_),
    .Y(_01018_),
    .B1(_07265_));
 sg13g2_inv_1 _15615_ (.Y(_07266_),
    .A(\synth.voice.accs[1][4] ));
 sg13g2_o21ai_1 _15616_ (.B1(_07258_),
    .Y(_07267_),
    .A1(_07256_),
    .A2(\synth.voice.accs[2][4] ));
 sg13g2_a21oi_1 _15617_ (.A1(net280),
    .A2(_07266_),
    .Y(_01019_),
    .B1(_07267_));
 sg13g2_inv_1 _15618_ (.Y(_07268_),
    .A(\synth.voice.accs[1][5] ));
 sg13g2_o21ai_1 _15619_ (.B1(net279),
    .Y(_07269_),
    .A1(net308),
    .A2(\synth.voice.accs[2][5] ));
 sg13g2_a21oi_1 _15620_ (.A1(net280),
    .A2(_07268_),
    .Y(_01020_),
    .B1(_07269_));
 sg13g2_inv_1 _15621_ (.Y(_07270_),
    .A(\synth.voice.accs[1][6] ));
 sg13g2_o21ai_1 _15622_ (.B1(net279),
    .Y(_07271_),
    .A1(net308),
    .A2(\synth.voice.accs[2][6] ));
 sg13g2_a21oi_1 _15623_ (.A1(net280),
    .A2(_07270_),
    .Y(_01021_),
    .B1(_07271_));
 sg13g2_inv_1 _15624_ (.Y(_07272_),
    .A(\synth.voice.accs[1][7] ));
 sg13g2_o21ai_1 _15625_ (.B1(net279),
    .Y(_07273_),
    .A1(net308),
    .A2(\synth.voice.accs[2][7] ));
 sg13g2_a21oi_1 _15626_ (.A1(net280),
    .A2(_07272_),
    .Y(_01022_),
    .B1(_07273_));
 sg13g2_inv_1 _15627_ (.Y(_07274_),
    .A(\synth.voice.accs[1][8] ));
 sg13g2_o21ai_1 _15628_ (.B1(net279),
    .Y(_07275_),
    .A1(net308),
    .A2(\synth.voice.accs[2][8] ));
 sg13g2_a21oi_1 _15629_ (.A1(net280),
    .A2(_07274_),
    .Y(_01023_),
    .B1(_07275_));
 sg13g2_inv_1 _15630_ (.Y(_07276_),
    .A(\synth.voice.accs[1][9] ));
 sg13g2_o21ai_1 _15631_ (.B1(net279),
    .Y(_07277_),
    .A1(net308),
    .A2(\synth.voice.accs[2][9] ));
 sg13g2_a21oi_1 _15632_ (.A1(net280),
    .A2(_07276_),
    .Y(_01024_),
    .B1(_07277_));
 sg13g2_buf_1 _15633_ (.A(_07187_),
    .X(_07278_));
 sg13g2_inv_1 _15634_ (.Y(_07279_),
    .A(\synth.voice.accs[2][0] ));
 sg13g2_buf_1 _15635_ (.A(net349),
    .X(_07280_));
 sg13g2_buf_1 _15636_ (.A(_07257_),
    .X(_07281_));
 sg13g2_o21ai_1 _15637_ (.B1(net277),
    .Y(_07282_),
    .A1(net307),
    .A2(\synth.voice.accs[3][0] ));
 sg13g2_a21oi_1 _15638_ (.A1(net278),
    .A2(_07279_),
    .Y(_01025_),
    .B1(_07282_));
 sg13g2_inv_1 _15639_ (.Y(_07283_),
    .A(\synth.voice.accs[2][10] ));
 sg13g2_o21ai_1 _15640_ (.B1(net277),
    .Y(_07284_),
    .A1(net307),
    .A2(\synth.voice.accs[3][10] ));
 sg13g2_a21oi_1 _15641_ (.A1(net278),
    .A2(_07283_),
    .Y(_01026_),
    .B1(_07284_));
 sg13g2_inv_1 _15642_ (.Y(_07285_),
    .A(\synth.voice.accs[2][11] ));
 sg13g2_o21ai_1 _15643_ (.B1(_07281_),
    .Y(_07286_),
    .A1(_07280_),
    .A2(\synth.voice.accs[3][11] ));
 sg13g2_a21oi_1 _15644_ (.A1(net278),
    .A2(_07285_),
    .Y(_01027_),
    .B1(_07286_));
 sg13g2_inv_1 _15645_ (.Y(_07287_),
    .A(\synth.voice.accs[2][12] ));
 sg13g2_o21ai_1 _15646_ (.B1(net277),
    .Y(_07288_),
    .A1(net307),
    .A2(\synth.voice.accs[3][12] ));
 sg13g2_a21oi_1 _15647_ (.A1(net278),
    .A2(_07287_),
    .Y(_01028_),
    .B1(_07288_));
 sg13g2_inv_1 _15648_ (.Y(_07289_),
    .A(\synth.voice.accs[2][13] ));
 sg13g2_o21ai_1 _15649_ (.B1(net277),
    .Y(_07290_),
    .A1(net307),
    .A2(\synth.voice.accs[3][13] ));
 sg13g2_a21oi_1 _15650_ (.A1(net278),
    .A2(_07289_),
    .Y(_01029_),
    .B1(_07290_));
 sg13g2_inv_1 _15651_ (.Y(_07291_),
    .A(\synth.voice.accs[2][14] ));
 sg13g2_o21ai_1 _15652_ (.B1(net277),
    .Y(_07292_),
    .A1(net307),
    .A2(\synth.voice.accs[3][14] ));
 sg13g2_a21oi_1 _15653_ (.A1(net278),
    .A2(_07291_),
    .Y(_01030_),
    .B1(_07292_));
 sg13g2_inv_1 _15654_ (.Y(_07293_),
    .A(\synth.voice.accs[2][15] ));
 sg13g2_o21ai_1 _15655_ (.B1(_07281_),
    .Y(_07294_),
    .A1(_07280_),
    .A2(\synth.voice.accs[3][15] ));
 sg13g2_a21oi_1 _15656_ (.A1(_07278_),
    .A2(_07293_),
    .Y(_01031_),
    .B1(_07294_));
 sg13g2_inv_1 _15657_ (.Y(_07295_),
    .A(\synth.voice.accs[2][16] ));
 sg13g2_o21ai_1 _15658_ (.B1(net277),
    .Y(_07296_),
    .A1(net307),
    .A2(\synth.voice.accs[3][16] ));
 sg13g2_a21oi_1 _15659_ (.A1(net278),
    .A2(_07295_),
    .Y(_01032_),
    .B1(_07296_));
 sg13g2_inv_1 _15660_ (.Y(_07297_),
    .A(\synth.voice.accs[2][17] ));
 sg13g2_o21ai_1 _15661_ (.B1(net277),
    .Y(_07298_),
    .A1(net307),
    .A2(\synth.voice.accs[3][17] ));
 sg13g2_a21oi_1 _15662_ (.A1(net278),
    .A2(_07297_),
    .Y(_01033_),
    .B1(_07298_));
 sg13g2_inv_1 _15663_ (.Y(_07299_),
    .A(\synth.voice.accs[2][18] ));
 sg13g2_o21ai_1 _15664_ (.B1(net277),
    .Y(_07300_),
    .A1(net307),
    .A2(\synth.voice.accs[3][18] ));
 sg13g2_a21oi_1 _15665_ (.A1(_07278_),
    .A2(_07299_),
    .Y(_01034_),
    .B1(_07300_));
 sg13g2_buf_1 _15666_ (.A(_07187_),
    .X(_07301_));
 sg13g2_inv_1 _15667_ (.Y(_07302_),
    .A(\synth.voice.accs[2][19] ));
 sg13g2_buf_1 _15668_ (.A(net349),
    .X(_07303_));
 sg13g2_buf_1 _15669_ (.A(_07257_),
    .X(_07304_));
 sg13g2_o21ai_1 _15670_ (.B1(net275),
    .Y(_07305_),
    .A1(net306),
    .A2(\synth.voice.accs[3][19] ));
 sg13g2_a21oi_1 _15671_ (.A1(net276),
    .A2(_07302_),
    .Y(_01035_),
    .B1(_07305_));
 sg13g2_inv_1 _15672_ (.Y(_07306_),
    .A(\synth.voice.accs[2][1] ));
 sg13g2_o21ai_1 _15673_ (.B1(_07304_),
    .Y(_07307_),
    .A1(_07303_),
    .A2(\synth.voice.accs[3][1] ));
 sg13g2_a21oi_1 _15674_ (.A1(_07301_),
    .A2(_07306_),
    .Y(_01036_),
    .B1(_07307_));
 sg13g2_inv_1 _15675_ (.Y(_07308_),
    .A(\synth.voice.accs[2][2] ));
 sg13g2_o21ai_1 _15676_ (.B1(_07304_),
    .Y(_07309_),
    .A1(_07303_),
    .A2(\synth.voice.accs[3][2] ));
 sg13g2_a21oi_1 _15677_ (.A1(_07301_),
    .A2(_07308_),
    .Y(_01037_),
    .B1(_07309_));
 sg13g2_inv_1 _15678_ (.Y(_07310_),
    .A(\synth.voice.accs[2][3] ));
 sg13g2_o21ai_1 _15679_ (.B1(net275),
    .Y(_07311_),
    .A1(net306),
    .A2(\synth.voice.accs[3][3] ));
 sg13g2_a21oi_1 _15680_ (.A1(net276),
    .A2(_07310_),
    .Y(_01038_),
    .B1(_07311_));
 sg13g2_inv_1 _15681_ (.Y(_07312_),
    .A(\synth.voice.accs[2][4] ));
 sg13g2_o21ai_1 _15682_ (.B1(net275),
    .Y(_07313_),
    .A1(net306),
    .A2(\synth.voice.accs[3][4] ));
 sg13g2_a21oi_1 _15683_ (.A1(net276),
    .A2(_07312_),
    .Y(_01039_),
    .B1(_07313_));
 sg13g2_inv_1 _15684_ (.Y(_07314_),
    .A(\synth.voice.accs[2][5] ));
 sg13g2_o21ai_1 _15685_ (.B1(net275),
    .Y(_07315_),
    .A1(net306),
    .A2(\synth.voice.accs[3][5] ));
 sg13g2_a21oi_1 _15686_ (.A1(net276),
    .A2(_07314_),
    .Y(_01040_),
    .B1(_07315_));
 sg13g2_inv_1 _15687_ (.Y(_07316_),
    .A(\synth.voice.accs[2][6] ));
 sg13g2_o21ai_1 _15688_ (.B1(net275),
    .Y(_07317_),
    .A1(net306),
    .A2(\synth.voice.accs[3][6] ));
 sg13g2_a21oi_1 _15689_ (.A1(net276),
    .A2(_07316_),
    .Y(_01041_),
    .B1(_07317_));
 sg13g2_inv_1 _15690_ (.Y(_07318_),
    .A(\synth.voice.accs[2][7] ));
 sg13g2_o21ai_1 _15691_ (.B1(net275),
    .Y(_07319_),
    .A1(net306),
    .A2(\synth.voice.accs[3][7] ));
 sg13g2_a21oi_1 _15692_ (.A1(net276),
    .A2(_07318_),
    .Y(_01042_),
    .B1(_07319_));
 sg13g2_inv_1 _15693_ (.Y(_07320_),
    .A(\synth.voice.accs[2][8] ));
 sg13g2_o21ai_1 _15694_ (.B1(net275),
    .Y(_07321_),
    .A1(net306),
    .A2(\synth.voice.accs[3][8] ));
 sg13g2_a21oi_1 _15695_ (.A1(net276),
    .A2(_07320_),
    .Y(_01043_),
    .B1(_07321_));
 sg13g2_inv_1 _15696_ (.Y(_07322_),
    .A(\synth.voice.accs[2][9] ));
 sg13g2_o21ai_1 _15697_ (.B1(net275),
    .Y(_07323_),
    .A1(net306),
    .A2(\synth.voice.accs[3][9] ));
 sg13g2_a21oi_1 _15698_ (.A1(net276),
    .A2(_07322_),
    .Y(_01044_),
    .B1(_07323_));
 sg13g2_buf_1 _15699_ (.A(_07187_),
    .X(_07324_));
 sg13g2_inv_1 _15700_ (.Y(_07325_),
    .A(\synth.voice.accs[3][0] ));
 sg13g2_buf_1 _15701_ (.A(_07139_),
    .X(_07326_));
 sg13g2_buf_1 _15702_ (.A(_07257_),
    .X(_07327_));
 sg13g2_o21ai_1 _15703_ (.B1(net273),
    .Y(_07328_),
    .A1(net305),
    .A2(\synth.voice.accs[4][0] ));
 sg13g2_a21oi_1 _15704_ (.A1(net274),
    .A2(_07325_),
    .Y(_01045_),
    .B1(_07328_));
 sg13g2_inv_1 _15705_ (.Y(_07329_),
    .A(\synth.voice.accs[3][10] ));
 sg13g2_o21ai_1 _15706_ (.B1(net273),
    .Y(_07330_),
    .A1(net305),
    .A2(\synth.voice.accs[4][10] ));
 sg13g2_a21oi_1 _15707_ (.A1(net274),
    .A2(_07329_),
    .Y(_01046_),
    .B1(_07330_));
 sg13g2_inv_1 _15708_ (.Y(_07331_),
    .A(\synth.voice.accs[3][11] ));
 sg13g2_o21ai_1 _15709_ (.B1(net273),
    .Y(_07332_),
    .A1(net305),
    .A2(\synth.voice.accs[4][11] ));
 sg13g2_a21oi_1 _15710_ (.A1(_07324_),
    .A2(_07331_),
    .Y(_01047_),
    .B1(_07332_));
 sg13g2_inv_1 _15711_ (.Y(_07333_),
    .A(\synth.voice.accs[3][12] ));
 sg13g2_o21ai_1 _15712_ (.B1(_07327_),
    .Y(_07334_),
    .A1(_07326_),
    .A2(\synth.voice.accs[4][12] ));
 sg13g2_a21oi_1 _15713_ (.A1(net274),
    .A2(_07333_),
    .Y(_01048_),
    .B1(_07334_));
 sg13g2_inv_1 _15714_ (.Y(_07335_),
    .A(\synth.voice.accs[3][13] ));
 sg13g2_o21ai_1 _15715_ (.B1(_07327_),
    .Y(_07336_),
    .A1(_07326_),
    .A2(\synth.voice.accs[4][13] ));
 sg13g2_a21oi_1 _15716_ (.A1(net274),
    .A2(_07335_),
    .Y(_01049_),
    .B1(_07336_));
 sg13g2_inv_1 _15717_ (.Y(_07337_),
    .A(\synth.voice.accs[3][14] ));
 sg13g2_o21ai_1 _15718_ (.B1(net273),
    .Y(_07338_),
    .A1(net305),
    .A2(\synth.voice.accs[4][14] ));
 sg13g2_a21oi_1 _15719_ (.A1(net274),
    .A2(_07337_),
    .Y(_01050_),
    .B1(_07338_));
 sg13g2_inv_1 _15720_ (.Y(_07339_),
    .A(\synth.voice.accs[3][15] ));
 sg13g2_o21ai_1 _15721_ (.B1(net273),
    .Y(_07340_),
    .A1(net305),
    .A2(\synth.voice.accs[4][15] ));
 sg13g2_a21oi_1 _15722_ (.A1(net274),
    .A2(_07339_),
    .Y(_01051_),
    .B1(_07340_));
 sg13g2_inv_1 _15723_ (.Y(_07341_),
    .A(\synth.voice.accs[3][16] ));
 sg13g2_o21ai_1 _15724_ (.B1(net273),
    .Y(_07342_),
    .A1(net305),
    .A2(\synth.voice.accs[4][16] ));
 sg13g2_a21oi_1 _15725_ (.A1(net274),
    .A2(_07341_),
    .Y(_01052_),
    .B1(_07342_));
 sg13g2_inv_1 _15726_ (.Y(_07343_),
    .A(\synth.voice.accs[3][17] ));
 sg13g2_o21ai_1 _15727_ (.B1(net273),
    .Y(_07344_),
    .A1(net305),
    .A2(\synth.voice.accs[4][17] ));
 sg13g2_a21oi_1 _15728_ (.A1(net274),
    .A2(_07343_),
    .Y(_01053_),
    .B1(_07344_));
 sg13g2_inv_1 _15729_ (.Y(_07345_),
    .A(\synth.voice.accs[3][18] ));
 sg13g2_o21ai_1 _15730_ (.B1(net273),
    .Y(_07346_),
    .A1(net305),
    .A2(\synth.voice.accs[4][18] ));
 sg13g2_a21oi_1 _15731_ (.A1(_07324_),
    .A2(_07345_),
    .Y(_01054_),
    .B1(_07346_));
 sg13g2_buf_1 _15732_ (.A(_07140_),
    .X(_07347_));
 sg13g2_inv_1 _15733_ (.Y(_07348_),
    .A(\synth.voice.accs[3][19] ));
 sg13g2_buf_1 _15734_ (.A(_07139_),
    .X(_07349_));
 sg13g2_buf_1 _15735_ (.A(_07257_),
    .X(_07350_));
 sg13g2_o21ai_1 _15736_ (.B1(net271),
    .Y(_07351_),
    .A1(net304),
    .A2(\synth.voice.accs[4][19] ));
 sg13g2_a21oi_1 _15737_ (.A1(net272),
    .A2(_07348_),
    .Y(_01055_),
    .B1(_07351_));
 sg13g2_inv_1 _15738_ (.Y(_07352_),
    .A(\synth.voice.accs[3][1] ));
 sg13g2_o21ai_1 _15739_ (.B1(_07350_),
    .Y(_07353_),
    .A1(_07349_),
    .A2(\synth.voice.accs[4][1] ));
 sg13g2_a21oi_1 _15740_ (.A1(_07347_),
    .A2(_07352_),
    .Y(_01056_),
    .B1(_07353_));
 sg13g2_inv_1 _15741_ (.Y(_07354_),
    .A(\synth.voice.accs[3][2] ));
 sg13g2_o21ai_1 _15742_ (.B1(_07350_),
    .Y(_07355_),
    .A1(_07349_),
    .A2(\synth.voice.accs[4][2] ));
 sg13g2_a21oi_1 _15743_ (.A1(_07347_),
    .A2(_07354_),
    .Y(_01057_),
    .B1(_07355_));
 sg13g2_inv_1 _15744_ (.Y(_07356_),
    .A(\synth.voice.accs[3][3] ));
 sg13g2_o21ai_1 _15745_ (.B1(net271),
    .Y(_07357_),
    .A1(net304),
    .A2(\synth.voice.accs[4][3] ));
 sg13g2_a21oi_1 _15746_ (.A1(net272),
    .A2(_07356_),
    .Y(_01058_),
    .B1(_07357_));
 sg13g2_inv_1 _15747_ (.Y(_07358_),
    .A(\synth.voice.accs[3][4] ));
 sg13g2_o21ai_1 _15748_ (.B1(net271),
    .Y(_07359_),
    .A1(net304),
    .A2(\synth.voice.accs[4][4] ));
 sg13g2_a21oi_1 _15749_ (.A1(net272),
    .A2(_07358_),
    .Y(_01059_),
    .B1(_07359_));
 sg13g2_inv_1 _15750_ (.Y(_07360_),
    .A(\synth.voice.accs[3][5] ));
 sg13g2_o21ai_1 _15751_ (.B1(net271),
    .Y(_07361_),
    .A1(net304),
    .A2(\synth.voice.accs[4][5] ));
 sg13g2_a21oi_1 _15752_ (.A1(net272),
    .A2(_07360_),
    .Y(_01060_),
    .B1(_07361_));
 sg13g2_inv_1 _15753_ (.Y(_07362_),
    .A(\synth.voice.accs[3][6] ));
 sg13g2_o21ai_1 _15754_ (.B1(net271),
    .Y(_07363_),
    .A1(net304),
    .A2(\synth.voice.accs[4][6] ));
 sg13g2_a21oi_1 _15755_ (.A1(net272),
    .A2(_07362_),
    .Y(_01061_),
    .B1(_07363_));
 sg13g2_inv_1 _15756_ (.Y(_07364_),
    .A(\synth.voice.accs[3][7] ));
 sg13g2_o21ai_1 _15757_ (.B1(net271),
    .Y(_07365_),
    .A1(net304),
    .A2(\synth.voice.accs[4][7] ));
 sg13g2_a21oi_1 _15758_ (.A1(net272),
    .A2(_07364_),
    .Y(_01062_),
    .B1(_07365_));
 sg13g2_inv_1 _15759_ (.Y(_07366_),
    .A(\synth.voice.accs[3][8] ));
 sg13g2_o21ai_1 _15760_ (.B1(net271),
    .Y(_07367_),
    .A1(net304),
    .A2(\synth.voice.accs[4][8] ));
 sg13g2_a21oi_1 _15761_ (.A1(net272),
    .A2(_07366_),
    .Y(_01063_),
    .B1(_07367_));
 sg13g2_inv_1 _15762_ (.Y(_07368_),
    .A(\synth.voice.accs[3][9] ));
 sg13g2_o21ai_1 _15763_ (.B1(net271),
    .Y(_07369_),
    .A1(net304),
    .A2(\synth.voice.accs[4][9] ));
 sg13g2_a21oi_1 _15764_ (.A1(net272),
    .A2(_07368_),
    .Y(_01064_),
    .B1(_07369_));
 sg13g2_buf_1 _15765_ (.A(net316),
    .X(_07370_));
 sg13g2_inv_1 _15766_ (.Y(_07371_),
    .A(\synth.voice.accs[4][0] ));
 sg13g2_buf_1 _15767_ (.A(_07139_),
    .X(_07372_));
 sg13g2_buf_1 _15768_ (.A(_07257_),
    .X(_07373_));
 sg13g2_o21ai_1 _15769_ (.B1(net269),
    .Y(_07374_),
    .A1(net303),
    .A2(\synth.voice.accs[5][0] ));
 sg13g2_a21oi_1 _15770_ (.A1(net270),
    .A2(_07371_),
    .Y(_01065_),
    .B1(_07374_));
 sg13g2_inv_1 _15771_ (.Y(_07375_),
    .A(\synth.voice.accs[4][10] ));
 sg13g2_o21ai_1 _15772_ (.B1(_07373_),
    .Y(_07376_),
    .A1(_07372_),
    .A2(\synth.voice.accs[5][10] ));
 sg13g2_a21oi_1 _15773_ (.A1(net270),
    .A2(_07375_),
    .Y(_01066_),
    .B1(_07376_));
 sg13g2_inv_1 _15774_ (.Y(_07377_),
    .A(\synth.voice.accs[4][11] ));
 sg13g2_o21ai_1 _15775_ (.B1(net269),
    .Y(_07378_),
    .A1(net303),
    .A2(\synth.voice.accs[5][11] ));
 sg13g2_a21oi_1 _15776_ (.A1(net270),
    .A2(_07377_),
    .Y(_01067_),
    .B1(_07378_));
 sg13g2_inv_1 _15777_ (.Y(_07379_),
    .A(\synth.voice.accs[4][12] ));
 sg13g2_o21ai_1 _15778_ (.B1(net269),
    .Y(_07380_),
    .A1(net303),
    .A2(\synth.voice.accs[5][12] ));
 sg13g2_a21oi_1 _15779_ (.A1(net270),
    .A2(_07379_),
    .Y(_01068_),
    .B1(_07380_));
 sg13g2_inv_1 _15780_ (.Y(_07381_),
    .A(\synth.voice.accs[4][13] ));
 sg13g2_o21ai_1 _15781_ (.B1(net269),
    .Y(_07382_),
    .A1(net303),
    .A2(\synth.voice.accs[5][13] ));
 sg13g2_a21oi_1 _15782_ (.A1(net270),
    .A2(_07381_),
    .Y(_01069_),
    .B1(_07382_));
 sg13g2_inv_1 _15783_ (.Y(_07383_),
    .A(\synth.voice.accs[4][14] ));
 sg13g2_o21ai_1 _15784_ (.B1(net269),
    .Y(_07384_),
    .A1(net303),
    .A2(\synth.voice.accs[5][14] ));
 sg13g2_a21oi_1 _15785_ (.A1(net270),
    .A2(_07383_),
    .Y(_01070_),
    .B1(_07384_));
 sg13g2_inv_1 _15786_ (.Y(_07385_),
    .A(\synth.voice.accs[4][15] ));
 sg13g2_o21ai_1 _15787_ (.B1(net269),
    .Y(_07386_),
    .A1(net303),
    .A2(\synth.voice.accs[5][15] ));
 sg13g2_a21oi_1 _15788_ (.A1(net270),
    .A2(_07385_),
    .Y(_01071_),
    .B1(_07386_));
 sg13g2_inv_1 _15789_ (.Y(_07387_),
    .A(\synth.voice.accs[4][16] ));
 sg13g2_o21ai_1 _15790_ (.B1(net269),
    .Y(_07388_),
    .A1(net303),
    .A2(\synth.voice.accs[5][16] ));
 sg13g2_a21oi_1 _15791_ (.A1(net270),
    .A2(_07387_),
    .Y(_01072_),
    .B1(_07388_));
 sg13g2_inv_1 _15792_ (.Y(_07389_),
    .A(\synth.voice.accs[4][17] ));
 sg13g2_o21ai_1 _15793_ (.B1(_07373_),
    .Y(_07390_),
    .A1(_07372_),
    .A2(\synth.voice.accs[5][17] ));
 sg13g2_a21oi_1 _15794_ (.A1(_07370_),
    .A2(_07389_),
    .Y(_01073_),
    .B1(_07390_));
 sg13g2_inv_1 _15795_ (.Y(_07391_),
    .A(\synth.voice.accs[4][18] ));
 sg13g2_o21ai_1 _15796_ (.B1(net269),
    .Y(_07392_),
    .A1(net303),
    .A2(\synth.voice.accs[5][18] ));
 sg13g2_a21oi_1 _15797_ (.A1(_07370_),
    .A2(_07391_),
    .Y(_01074_),
    .B1(_07392_));
 sg13g2_buf_1 _15798_ (.A(_07140_),
    .X(_07393_));
 sg13g2_inv_1 _15799_ (.Y(_07394_),
    .A(\synth.voice.accs[4][19] ));
 sg13g2_buf_1 _15800_ (.A(_07139_),
    .X(_07395_));
 sg13g2_buf_1 _15801_ (.A(_07257_),
    .X(_07396_));
 sg13g2_o21ai_1 _15802_ (.B1(net267),
    .Y(_07397_),
    .A1(net302),
    .A2(\synth.voice.accs[5][19] ));
 sg13g2_a21oi_1 _15803_ (.A1(net268),
    .A2(_07394_),
    .Y(_01075_),
    .B1(_07397_));
 sg13g2_inv_1 _15804_ (.Y(_07398_),
    .A(\synth.voice.accs[4][1] ));
 sg13g2_o21ai_1 _15805_ (.B1(net267),
    .Y(_07399_),
    .A1(net302),
    .A2(\synth.voice.accs[5][1] ));
 sg13g2_a21oi_1 _15806_ (.A1(net268),
    .A2(_07398_),
    .Y(_01076_),
    .B1(_07399_));
 sg13g2_inv_1 _15807_ (.Y(_07400_),
    .A(\synth.voice.accs[4][2] ));
 sg13g2_o21ai_1 _15808_ (.B1(net267),
    .Y(_07401_),
    .A1(net302),
    .A2(\synth.voice.accs[5][2] ));
 sg13g2_a21oi_1 _15809_ (.A1(net268),
    .A2(_07400_),
    .Y(_01077_),
    .B1(_07401_));
 sg13g2_inv_1 _15810_ (.Y(_07402_),
    .A(\synth.voice.accs[4][3] ));
 sg13g2_o21ai_1 _15811_ (.B1(net267),
    .Y(_07403_),
    .A1(net302),
    .A2(\synth.voice.accs[5][3] ));
 sg13g2_a21oi_1 _15812_ (.A1(net268),
    .A2(_07402_),
    .Y(_01078_),
    .B1(_07403_));
 sg13g2_inv_1 _15813_ (.Y(_07404_),
    .A(\synth.voice.accs[4][4] ));
 sg13g2_o21ai_1 _15814_ (.B1(net267),
    .Y(_07405_),
    .A1(net302),
    .A2(\synth.voice.accs[5][4] ));
 sg13g2_a21oi_1 _15815_ (.A1(net268),
    .A2(_07404_),
    .Y(_01079_),
    .B1(_07405_));
 sg13g2_inv_1 _15816_ (.Y(_07406_),
    .A(\synth.voice.accs[4][5] ));
 sg13g2_o21ai_1 _15817_ (.B1(_07396_),
    .Y(_07407_),
    .A1(_07395_),
    .A2(\synth.voice.accs[5][5] ));
 sg13g2_a21oi_1 _15818_ (.A1(_07393_),
    .A2(_07406_),
    .Y(_01080_),
    .B1(_07407_));
 sg13g2_inv_1 _15819_ (.Y(_07408_),
    .A(\synth.voice.accs[4][6] ));
 sg13g2_o21ai_1 _15820_ (.B1(_07396_),
    .Y(_07409_),
    .A1(_07395_),
    .A2(\synth.voice.accs[5][6] ));
 sg13g2_a21oi_1 _15821_ (.A1(_07393_),
    .A2(_07408_),
    .Y(_01081_),
    .B1(_07409_));
 sg13g2_inv_1 _15822_ (.Y(_07410_),
    .A(\synth.voice.accs[4][7] ));
 sg13g2_o21ai_1 _15823_ (.B1(net267),
    .Y(_07411_),
    .A1(net302),
    .A2(\synth.voice.accs[5][7] ));
 sg13g2_a21oi_1 _15824_ (.A1(net268),
    .A2(_07410_),
    .Y(_01082_),
    .B1(_07411_));
 sg13g2_inv_1 _15825_ (.Y(_07412_),
    .A(\synth.voice.accs[4][8] ));
 sg13g2_o21ai_1 _15826_ (.B1(net267),
    .Y(_07413_),
    .A1(net302),
    .A2(\synth.voice.accs[5][8] ));
 sg13g2_a21oi_1 _15827_ (.A1(net268),
    .A2(_07412_),
    .Y(_01083_),
    .B1(_07413_));
 sg13g2_inv_1 _15828_ (.Y(_07414_),
    .A(\synth.voice.accs[4][9] ));
 sg13g2_o21ai_1 _15829_ (.B1(net267),
    .Y(_07415_),
    .A1(net302),
    .A2(\synth.voice.accs[5][9] ));
 sg13g2_a21oi_1 _15830_ (.A1(net268),
    .A2(_07414_),
    .Y(_01084_),
    .B1(_07415_));
 sg13g2_a21oi_1 _15831_ (.A1(_05762_),
    .A2(\synth.voice.coeff_index[2] ),
    .Y(_07416_),
    .B1(_07023_));
 sg13g2_nand2b_1 _15832_ (.Y(_07417_),
    .B(_07024_),
    .A_N(_07416_));
 sg13g2_xor2_1 _15833_ (.B(_07417_),
    .A(_00052_),
    .X(_07418_));
 sg13g2_xnor2_1 _15834_ (.Y(_07419_),
    .A(\synth.voice.coeff_index[4] ),
    .B(_07025_));
 sg13g2_nor2_1 _15835_ (.A(_06667_),
    .B(_07419_),
    .Y(_07420_));
 sg13g2_nor3_1 _15836_ (.A(net183),
    .B(_07418_),
    .C(_07420_),
    .Y(_07421_));
 sg13g2_nand2_1 _15837_ (.Y(_07422_),
    .A(_07419_),
    .B(_06667_));
 sg13g2_nand2_1 _15838_ (.Y(_07423_),
    .A(_07421_),
    .B(_07422_));
 sg13g2_buf_2 _15839_ (.A(_07423_),
    .X(_07424_));
 sg13g2_nand2_1 _15840_ (.Y(_07425_),
    .A(net183),
    .B(_03441_));
 sg13g2_nand3b_1 _15841_ (.B(_07424_),
    .C(_07425_),
    .Y(_07426_),
    .A_N(_03449_));
 sg13g2_inv_1 _15842_ (.Y(_07427_),
    .A(_07424_));
 sg13g2_nand2_1 _15843_ (.Y(_07428_),
    .A(_07427_),
    .B(\synth.voice.oct_counter[0] ));
 sg13g2_a21oi_1 _15844_ (.A1(_07426_),
    .A2(_07428_),
    .Y(_01087_),
    .B1(net318));
 sg13g2_nand2_1 _15845_ (.Y(_07429_),
    .A(_03553_),
    .B(_03554_));
 sg13g2_buf_1 _15846_ (.A(_07424_),
    .X(_07430_));
 sg13g2_buf_2 _15847_ (.A(_01798_),
    .X(_07431_));
 sg13g2_o21ai_1 _15848_ (.B1(net301),
    .Y(_07432_),
    .A1(\synth.voice.oct_counter[10] ),
    .A2(net111));
 sg13g2_a21oi_1 _15849_ (.A1(_07429_),
    .A2(net111),
    .Y(_01088_),
    .B1(_07432_));
 sg13g2_xnor2_1 _15850_ (.Y(_07433_),
    .A(_03460_),
    .B(_03449_));
 sg13g2_o21ai_1 _15851_ (.B1(_07431_),
    .Y(_07434_),
    .A1(\synth.voice.oct_counter[1] ),
    .A2(net111));
 sg13g2_a21oi_1 _15852_ (.A1(net111),
    .A2(_07433_),
    .Y(_01089_),
    .B1(_07434_));
 sg13g2_o21ai_1 _15853_ (.B1(net301),
    .Y(_07435_),
    .A1(\synth.voice.oct_counter[2] ),
    .A2(_07424_));
 sg13g2_a21oi_1 _15854_ (.A1(_03469_),
    .A2(net111),
    .Y(_01090_),
    .B1(_07435_));
 sg13g2_inv_1 _15855_ (.Y(_07436_),
    .A(_03492_));
 sg13g2_o21ai_1 _15856_ (.B1(net301),
    .Y(_07437_),
    .A1(_03464_),
    .A2(_07427_));
 sg13g2_a21oi_1 _15857_ (.A1(_07436_),
    .A2(_07427_),
    .Y(_01091_),
    .B1(_07437_));
 sg13g2_o21ai_1 _15858_ (.B1(net301),
    .Y(_07438_),
    .A1(_03489_),
    .A2(_07424_));
 sg13g2_a21oi_1 _15859_ (.A1(_03524_),
    .A2(net111),
    .Y(_01092_),
    .B1(_07438_));
 sg13g2_o21ai_1 _15860_ (.B1(net301),
    .Y(_07439_),
    .A1(_03527_),
    .A2(_07427_));
 sg13g2_a21oi_1 _15861_ (.A1(_03495_),
    .A2(_07427_),
    .Y(_01093_),
    .B1(_07439_));
 sg13g2_nand2_1 _15862_ (.Y(_07440_),
    .A(_03518_),
    .B(_03520_));
 sg13g2_o21ai_1 _15863_ (.B1(net301),
    .Y(_07441_),
    .A1(\synth.voice.oct_counter[6] ),
    .A2(_07424_));
 sg13g2_a21oi_1 _15864_ (.A1(_07440_),
    .A2(net111),
    .Y(_01094_),
    .B1(_07441_));
 sg13g2_inv_1 _15865_ (.Y(_07442_),
    .A(_03504_));
 sg13g2_o21ai_1 _15866_ (.B1(net301),
    .Y(_07443_),
    .A1(_03482_),
    .A2(_07424_));
 sg13g2_a21oi_1 _15867_ (.A1(_07442_),
    .A2(_07430_),
    .Y(_01095_),
    .B1(_07443_));
 sg13g2_a21oi_1 _15868_ (.A1(_03577_),
    .A2(_03578_),
    .Y(_07444_),
    .B1(_07427_));
 sg13g2_o21ai_1 _15869_ (.B1(_07064_),
    .Y(_07445_),
    .A1(_03540_),
    .A2(_07430_));
 sg13g2_nor2_1 _15870_ (.A(_07444_),
    .B(_07445_),
    .Y(_01096_));
 sg13g2_o21ai_1 _15871_ (.B1(net301),
    .Y(_07446_),
    .A1(_03535_),
    .A2(_07424_));
 sg13g2_a21oi_1 _15872_ (.A1(_03571_),
    .A2(net111),
    .Y(_01097_),
    .B1(_07446_));
 sg13g2_inv_1 _15873_ (.Y(_07447_),
    .A(\synth.voice.next_sweep_oct_counter[0] ));
 sg13g2_buf_8 _15874_ (.A(_07049_),
    .X(_07448_));
 sg13g2_o21ai_1 _15875_ (.B1(_07431_),
    .Y(_07449_),
    .A1(_03948_),
    .A2(net73));
 sg13g2_a21oi_1 _15876_ (.A1(_07447_),
    .A2(net73),
    .Y(_01290_),
    .B1(_07449_));
 sg13g2_nor2_1 _15877_ (.A(_03992_),
    .B(_07050_),
    .Y(_07450_));
 sg13g2_nor3_1 _15878_ (.A(_03987_),
    .B(_04003_),
    .C(_03989_),
    .Y(_07451_));
 sg13g2_a21oi_1 _15879_ (.A1(net73),
    .A2(_07451_),
    .Y(_07452_),
    .B1(\synth.voice.sweep_oct_counter[10] ));
 sg13g2_nor3_1 _15880_ (.A(net394),
    .B(_07450_),
    .C(_07452_),
    .Y(_01291_));
 sg13g2_nand2_1 _15881_ (.Y(_07453_),
    .A(net73),
    .B(_03996_));
 sg13g2_nand2_1 _15882_ (.Y(_07454_),
    .A(_07453_),
    .B(net290));
 sg13g2_nor2_1 _15883_ (.A(_03982_),
    .B(_07450_),
    .Y(_07455_));
 sg13g2_nor2_1 _15884_ (.A(_07454_),
    .B(_07455_),
    .Y(_01292_));
 sg13g2_a21oi_1 _15885_ (.A1(net73),
    .A2(_03996_),
    .Y(_07456_),
    .B1(\synth.voice.sweep_oct_counter[12] ));
 sg13g2_nor2_1 _15886_ (.A(_03983_),
    .B(_07453_),
    .Y(_07457_));
 sg13g2_nor3_1 _15887_ (.A(_01790_),
    .B(_07456_),
    .C(_07457_),
    .Y(_01293_));
 sg13g2_nand4_1 _15888_ (.B(\synth.controller.curr_voice[1] ),
    .C(\synth.controller.curr_voice[0] ),
    .A(_06816_),
    .Y(_07458_),
    .D(_06813_));
 sg13g2_buf_2 _15889_ (.A(_07458_),
    .X(_07459_));
 sg13g2_inv_4 _15890_ (.A(_07459_),
    .Y(_07460_));
 sg13g2_nand2_1 _15891_ (.Y(_07461_),
    .A(\synth.voice.sweep_oct_counter[9] ),
    .B(\synth.voice.sweep_oct_counter[10] ));
 sg13g2_nand2_1 _15892_ (.Y(_07462_),
    .A(_03982_),
    .B(\synth.voice.sweep_oct_counter[12] ));
 sg13g2_nand4_1 _15893_ (.B(_03961_),
    .C(_03988_),
    .A(\synth.voice.sweep_oct_counter[5] ),
    .Y(_07463_),
    .D(\synth.voice.sweep_oct_counter[8] ));
 sg13g2_nor4_1 _15894_ (.A(_07461_),
    .B(_07462_),
    .C(_07463_),
    .D(_03970_),
    .Y(_07464_));
 sg13g2_xnor2_1 _15895_ (.Y(_07465_),
    .A(_03994_),
    .B(_07464_));
 sg13g2_nand2_1 _15896_ (.Y(_07466_),
    .A(_07460_),
    .B(_07465_));
 sg13g2_nand2_1 _15897_ (.Y(_07467_),
    .A(_07459_),
    .B(\synth.voice.sweep_oct_counter[13] ));
 sg13g2_a21oi_1 _15898_ (.A1(_07466_),
    .A2(_07467_),
    .Y(_01294_),
    .B1(net318));
 sg13g2_nand2_1 _15899_ (.Y(_07468_),
    .A(_07049_),
    .B(_03951_));
 sg13g2_nand2_1 _15900_ (.Y(_07469_),
    .A(_07468_),
    .B(net290));
 sg13g2_a21oi_1 _15901_ (.A1(net73),
    .A2(_03948_),
    .Y(_07470_),
    .B1(\synth.voice.sweep_oct_counter[1] ));
 sg13g2_nor2_1 _15902_ (.A(_07469_),
    .B(_07470_),
    .Y(_01295_));
 sg13g2_a21oi_1 _15903_ (.A1(net73),
    .A2(_03951_),
    .Y(_07471_),
    .B1(\synth.voice.sweep_oct_counter[2] ));
 sg13g2_nor2_1 _15904_ (.A(_03953_),
    .B(_07468_),
    .Y(_07472_));
 sg13g2_nor3_1 _15905_ (.A(_01790_),
    .B(_07471_),
    .C(_07472_),
    .Y(_01296_));
 sg13g2_xnor2_1 _15906_ (.Y(_07473_),
    .A(_03964_),
    .B(_03965_));
 sg13g2_nand2_1 _15907_ (.Y(_07474_),
    .A(_07460_),
    .B(_07473_));
 sg13g2_nand2_1 _15908_ (.Y(_07475_),
    .A(_07459_),
    .B(\synth.voice.sweep_oct_counter[3] ));
 sg13g2_a21oi_1 _15909_ (.A1(_07474_),
    .A2(_07475_),
    .Y(_01297_),
    .B1(_07052_));
 sg13g2_xnor2_1 _15910_ (.Y(_07476_),
    .A(_03963_),
    .B(_03967_));
 sg13g2_nand2_1 _15911_ (.Y(_07477_),
    .A(_07460_),
    .B(_07476_));
 sg13g2_nand2_1 _15912_ (.Y(_07478_),
    .A(_07459_),
    .B(\synth.voice.sweep_oct_counter[4] ));
 sg13g2_a21oi_1 _15913_ (.A1(_07477_),
    .A2(_07478_),
    .Y(_01298_),
    .B1(_07052_));
 sg13g2_nand2_1 _15914_ (.Y(_07479_),
    .A(_07460_),
    .B(_03969_));
 sg13g2_o21ai_1 _15915_ (.B1(net319),
    .Y(_07480_),
    .A1(_03972_),
    .A2(_07050_));
 sg13g2_a21oi_1 _15916_ (.A1(_07479_),
    .A2(_03962_),
    .Y(_01299_),
    .B1(_07480_));
 sg13g2_nor2_1 _15917_ (.A(_03972_),
    .B(_07050_),
    .Y(_07481_));
 sg13g2_nor2_1 _15918_ (.A(_03961_),
    .B(_07481_),
    .Y(_07482_));
 sg13g2_nand2_1 _15919_ (.Y(_07483_),
    .A(_07481_),
    .B(_03961_));
 sg13g2_nand2_1 _15920_ (.Y(_07484_),
    .A(_07483_),
    .B(net290));
 sg13g2_nor2_1 _15921_ (.A(_07482_),
    .B(_07484_),
    .Y(_01300_));
 sg13g2_inv_1 _15922_ (.Y(_07485_),
    .A(_03988_));
 sg13g2_nand2b_1 _15923_ (.Y(_07486_),
    .B(net73),
    .A_N(_03989_));
 sg13g2_nand2_1 _15924_ (.Y(_07487_),
    .A(_07486_),
    .B(net290));
 sg13g2_a21oi_1 _15925_ (.A1(_07483_),
    .A2(_07485_),
    .Y(_01301_),
    .B1(_07487_));
 sg13g2_nand2_1 _15926_ (.Y(_07488_),
    .A(_07448_),
    .B(_03990_));
 sg13g2_nand2_1 _15927_ (.Y(_07489_),
    .A(_07488_),
    .B(net289));
 sg13g2_a21oi_1 _15928_ (.A1(_03987_),
    .A2(_07486_),
    .Y(_01302_),
    .B1(_07489_));
 sg13g2_nand2_1 _15929_ (.Y(_07490_),
    .A(_07448_),
    .B(_07451_));
 sg13g2_nand2_1 _15930_ (.Y(_07491_),
    .A(_07490_),
    .B(net289));
 sg13g2_a21oi_1 _15931_ (.A1(_04003_),
    .A2(_07488_),
    .Y(_01303_),
    .B1(_07491_));
 sg13g2_a21oi_1 _15932_ (.A1(_06799_),
    .A2(_06802_),
    .Y(_07492_),
    .B1(_06666_));
 sg13g2_a21oi_1 _15933_ (.A1(_00049_),
    .A2(_01722_),
    .Y(_07493_),
    .B1(_06803_));
 sg13g2_nor3_1 _15934_ (.A(net394),
    .B(_07492_),
    .C(_07493_),
    .Y(_01304_));
 sg13g2_o21ai_1 _15935_ (.B1(net319),
    .Y(_07494_),
    .A1(_01751_),
    .A2(_06803_));
 sg13g2_a21oi_1 _15936_ (.A1(_01720_),
    .A2(_06803_),
    .Y(_01305_),
    .B1(_07494_));
 sg13g2_xnor2_1 _15937_ (.Y(_07495_),
    .A(_00048_),
    .B(_01731_));
 sg13g2_nand2_1 _15938_ (.Y(_07496_),
    .A(_06803_),
    .B(_00080_));
 sg13g2_nor2_1 _15939_ (.A(_07495_),
    .B(_07496_),
    .Y(_01306_));
 sg13g2_nor3_1 _15940_ (.A(_01793_),
    .B(_06741_),
    .C(_01731_),
    .Y(_07497_));
 sg13g2_a21oi_1 _15941_ (.A1(_01732_),
    .A2(_01715_),
    .Y(_07498_),
    .B1(_01716_));
 sg13g2_nor3_1 _15942_ (.A(_07497_),
    .B(_07498_),
    .C(_07496_),
    .Y(_01307_));
 sg13g2_xnor2_1 _15943_ (.Y(_07499_),
    .A(_06744_),
    .B(_07497_));
 sg13g2_nor2_1 _15944_ (.A(_07499_),
    .B(_07496_),
    .Y(_01308_));
 sg13g2_inv_1 _15945_ (.Y(_07500_),
    .A(_07103_));
 sg13g2_inv_1 _15946_ (.Y(_07501_),
    .A(_03400_));
 sg13g2_nand2_1 _15947_ (.Y(_07502_),
    .A(_03400_),
    .B(_00146_));
 sg13g2_nand3_1 _15948_ (.B(_03402_),
    .C(_03403_),
    .A(_07502_),
    .Y(_07503_));
 sg13g2_a21oi_1 _15949_ (.A1(_03393_),
    .A2(_07501_),
    .Y(_07504_),
    .B1(_07503_));
 sg13g2_nor2_1 _15950_ (.A(_03595_),
    .B(_04785_),
    .Y(_07505_));
 sg13g2_nor3_1 _15951_ (.A(_04025_),
    .B(_04812_),
    .C(_07505_),
    .Y(_07506_));
 sg13g2_nor2_1 _15952_ (.A(_05096_),
    .B(_05732_),
    .Y(_07507_));
 sg13g2_a221oi_1 _15953_ (.B2(_05525_),
    .C1(_07507_),
    .B1(\synth.voice.scan_outs[2][1] ),
    .A1(_04786_),
    .Y(_07508_),
    .A2(_04491_));
 sg13g2_a22oi_1 _15954_ (.Y(_07509_),
    .B1(_05040_),
    .B2(_05821_),
    .A2(\synth.voice.float_period[0][9] ),
    .A1(_05908_));
 sg13g2_inv_1 _15955_ (.Y(_07510_),
    .A(_04251_));
 sg13g2_a22oi_1 _15956_ (.Y(_07511_),
    .B1(_03437_),
    .B2(_04030_),
    .A2(\synth.voice.mods[1][3] ),
    .A1(_07510_));
 sg13g2_nor2_1 _15957_ (.A(_00081_),
    .B(_04718_),
    .Y(_07512_));
 sg13g2_nor2b_1 _15958_ (.A(_04813_),
    .B_N(_01765_),
    .Y(_07513_));
 sg13g2_nor2_1 _15959_ (.A(_00147_),
    .B(_04352_),
    .Y(_07514_));
 sg13g2_and3_1 _15960_ (.X(_07515_),
    .A(_04028_),
    .B(\synth.voice.params[25] ),
    .C(_04812_));
 sg13g2_nor4_1 _15961_ (.A(_07512_),
    .B(_07513_),
    .C(_07514_),
    .D(_07515_),
    .Y(_07516_));
 sg13g2_nand4_1 _15962_ (.B(_07509_),
    .C(_07511_),
    .A(_07508_),
    .Y(_07517_),
    .D(_07516_));
 sg13g2_a21oi_1 _15963_ (.A1(\synth.voice.delayed_p[0] ),
    .A2(_07506_),
    .Y(_07518_),
    .B1(_07517_));
 sg13g2_a21oi_1 _15964_ (.A1(_03308_),
    .A2(\synth.controller.out_reg[1] ),
    .Y(_07519_),
    .B1(_07103_));
 sg13g2_o21ai_1 _15965_ (.B1(_07519_),
    .Y(_07520_),
    .A1(_03308_),
    .A2(_07518_));
 sg13g2_o21ai_1 _15966_ (.B1(_07520_),
    .Y(_07521_),
    .A1(_07500_),
    .A2(_07504_));
 sg13g2_o21ai_1 _15967_ (.B1(_07093_),
    .Y(_07522_),
    .A1(_03404_),
    .A2(_03305_));
 sg13g2_a21oi_1 _15968_ (.A1(_07521_),
    .A2(_03404_),
    .Y(_01319_),
    .B1(_07522_));
 sg13g2_buf_1 _15969_ (.A(_02220_),
    .X(_07523_));
 sg13g2_nand2_1 _15970_ (.Y(_07524_),
    .A(_02269_),
    .B(net239));
 sg13g2_nand2_1 _15971_ (.Y(_07525_),
    .A(_03306_),
    .B(_03305_));
 sg13g2_o21ai_1 _15972_ (.B1(\synth.controller.ext_tx_request ),
    .Y(_07526_),
    .A1(_07525_),
    .A2(_07053_));
 sg13g2_nand2_1 _15973_ (.Y(_07527_),
    .A(net290),
    .B(\ppu_ctrl[2] ));
 sg13g2_a21oi_1 _15974_ (.A1(_07524_),
    .A2(_07526_),
    .Y(_01320_),
    .B1(_07527_));
 sg13g2_nor4_2 _15975_ (.A(_02420_),
    .B(_02451_),
    .C(_02476_),
    .Y(_07528_),
    .D(_02379_));
 sg13g2_inv_1 _15976_ (.Y(_07529_),
    .A(_07528_));
 sg13g2_o21ai_1 _15977_ (.B1(_07523_),
    .Y(_07530_),
    .A1(_02290_),
    .A2(net110));
 sg13g2_a21o_1 _15978_ (.A2(net110),
    .A1(_06566_),
    .B1(_07530_),
    .X(_00266_));
 sg13g2_o21ai_1 _15979_ (.B1(_07523_),
    .Y(_07531_),
    .A1(net340),
    .A2(net110));
 sg13g2_a21o_1 _15980_ (.A2(net110),
    .A1(_06579_),
    .B1(_07531_),
    .X(_00267_));
 sg13g2_a21oi_1 _15981_ (.A1(_07528_),
    .A2(_02396_),
    .Y(_07532_),
    .B1(net250));
 sg13g2_o21ai_1 _15982_ (.B1(_07532_),
    .Y(_00268_),
    .A1(_06101_),
    .A2(_07528_));
 sg13g2_a21oi_1 _15983_ (.A1(net110),
    .A2(\ppu.display_mask[3] ),
    .Y(_07533_),
    .B1(_02198_));
 sg13g2_o21ai_1 _15984_ (.B1(_07533_),
    .Y(_00269_),
    .A1(net338),
    .A2(net110));
 sg13g2_a21oi_1 _15985_ (.A1(net110),
    .A2(\ppu.display_mask[4] ),
    .Y(_07534_),
    .B1(_02198_));
 sg13g2_o21ai_1 _15986_ (.B1(_07534_),
    .Y(_00270_),
    .A1(_02406_),
    .A2(net110));
 sg13g2_o21ai_1 _15987_ (.B1(net239),
    .Y(_07535_),
    .A1(net387),
    .A2(_07529_));
 sg13g2_a21o_1 _15988_ (.A2(_07529_),
    .A1(\ppu.display_mask[5] ),
    .B1(_07535_),
    .X(_00271_));
 sg13g2_nand2_1 _15989_ (.Y(_07536_),
    .A(_02605_),
    .B(_02477_));
 sg13g2_buf_1 _15990_ (.A(_07536_),
    .X(_07537_));
 sg13g2_buf_1 _15991_ (.A(_07537_),
    .X(_07538_));
 sg13g2_o21ai_1 _15992_ (.B1(_02221_),
    .Y(_07539_),
    .A1(\ppu.copper_inst.store[7] ),
    .A2(_07537_));
 sg13g2_a21oi_1 _15993_ (.A1(_02201_),
    .A2(_07538_),
    .Y(_00272_),
    .B1(_07539_));
 sg13g2_inv_1 _15994_ (.Y(_07540_),
    .A(_07537_));
 sg13g2_o21ai_1 _15995_ (.B1(net249),
    .Y(_07541_),
    .A1(\ppu.gfxmode1[1] ),
    .A2(_07540_));
 sg13g2_a21oi_1 _15996_ (.A1(net340),
    .A2(_07540_),
    .Y(_00273_),
    .B1(_07541_));
 sg13g2_o21ai_1 _15997_ (.B1(_02221_),
    .Y(_07542_),
    .A1(_02396_),
    .A2(_07537_));
 sg13g2_a21oi_1 _15998_ (.A1(_02219_),
    .A2(_07538_),
    .Y(_00274_),
    .B1(_07542_));
 sg13g2_a21oi_1 _15999_ (.A1(net92),
    .A2(\ppu.gfxmode1[3] ),
    .Y(_07543_),
    .B1(net250));
 sg13g2_o21ai_1 _16000_ (.B1(_07543_),
    .Y(_00275_),
    .A1(net338),
    .A2(net92));
 sg13g2_a21oi_1 _16001_ (.A1(net92),
    .A2(\ppu.gfxmode1[4] ),
    .Y(_07544_),
    .B1(net250));
 sg13g2_o21ai_1 _16002_ (.B1(_07544_),
    .Y(_00276_),
    .A1(net337),
    .A2(net92));
 sg13g2_a21oi_1 _16003_ (.A1(net92),
    .A2(\ppu.gfxmode1[5] ),
    .Y(_07545_),
    .B1(net250));
 sg13g2_o21ai_1 _16004_ (.B1(_07545_),
    .Y(_00277_),
    .A1(net387),
    .A2(net92));
 sg13g2_a21oi_1 _16005_ (.A1(net92),
    .A2(\ppu.gfxmode1[6] ),
    .Y(_07546_),
    .B1(net250));
 sg13g2_o21ai_1 _16006_ (.B1(_07546_),
    .Y(_00278_),
    .A1(_02412_),
    .A2(net92));
 sg13g2_o21ai_1 _16007_ (.B1(net249),
    .Y(_07547_),
    .A1(\ppu.gfxmode1[7] ),
    .A2(_07540_));
 sg13g2_a21oi_1 _16008_ (.A1(net386),
    .A2(_07540_),
    .Y(_00279_),
    .B1(_07547_));
 sg13g2_buf_1 _16009_ (.A(net298),
    .X(_07548_));
 sg13g2_a21oi_1 _16010_ (.A1(_07540_),
    .A2(_02417_),
    .Y(_07549_),
    .B1(net257));
 sg13g2_o21ai_1 _16011_ (.B1(_07549_),
    .Y(_00280_),
    .A1(_01832_),
    .A2(_07540_));
 sg13g2_nand2_1 _16012_ (.Y(_07550_),
    .A(_02625_),
    .B(_02477_));
 sg13g2_inv_2 _16013_ (.Y(_07551_),
    .A(_07550_));
 sg13g2_buf_1 _16014_ (.A(_02220_),
    .X(_07552_));
 sg13g2_o21ai_1 _16015_ (.B1(net238),
    .Y(_07553_),
    .A1(\ppu.gfxmode2[0] ),
    .A2(_07551_));
 sg13g2_a21oi_1 _16016_ (.A1(net388),
    .A2(_07551_),
    .Y(_00281_),
    .B1(_07553_));
 sg13g2_o21ai_1 _16017_ (.B1(net238),
    .Y(_07554_),
    .A1(\ppu.gfxmode2[1] ),
    .A2(_07551_));
 sg13g2_a21oi_1 _16018_ (.A1(net340),
    .A2(_07551_),
    .Y(_00282_),
    .B1(_07554_));
 sg13g2_o21ai_1 _16019_ (.B1(net238),
    .Y(_07555_),
    .A1(\ppu.gfxmode2[2] ),
    .A2(_07551_));
 sg13g2_a21oi_1 _16020_ (.A1(net339),
    .A2(_07551_),
    .Y(_00283_),
    .B1(_07555_));
 sg13g2_buf_1 _16021_ (.A(_07550_),
    .X(_07556_));
 sg13g2_a21oi_1 _16022_ (.A1(net103),
    .A2(\ppu.gfxmode2[3] ),
    .Y(_07557_),
    .B1(net257));
 sg13g2_o21ai_1 _16023_ (.B1(_07557_),
    .Y(_00284_),
    .A1(net338),
    .A2(net103));
 sg13g2_o21ai_1 _16024_ (.B1(net238),
    .Y(_07558_),
    .A1(\ppu.gfxmode2[4] ),
    .A2(_07551_));
 sg13g2_a21oi_1 _16025_ (.A1(net337),
    .A2(_07551_),
    .Y(_00285_),
    .B1(_07558_));
 sg13g2_buf_1 _16026_ (.A(\ppu.gfxmode2[5] ),
    .X(_07559_));
 sg13g2_inv_1 _16027_ (.Y(_07560_),
    .A(_07559_));
 sg13g2_o21ai_1 _16028_ (.B1(net238),
    .Y(_07561_),
    .A1(_02408_),
    .A2(net103));
 sg13g2_a21oi_1 _16029_ (.A1(_07560_),
    .A2(net103),
    .Y(_00286_),
    .B1(_07561_));
 sg13g2_buf_1 _16030_ (.A(\ppu.gfxmode2[6] ),
    .X(_07562_));
 sg13g2_inv_1 _16031_ (.Y(_07563_),
    .A(_07562_));
 sg13g2_o21ai_1 _16032_ (.B1(net238),
    .Y(_07564_),
    .A1(net406),
    .A2(net103));
 sg13g2_a21oi_1 _16033_ (.A1(_07563_),
    .A2(net103),
    .Y(_00287_),
    .B1(_07564_));
 sg13g2_o21ai_1 _16034_ (.B1(net239),
    .Y(_07565_),
    .A1(net386),
    .A2(net103));
 sg13g2_a21o_1 _16035_ (.A2(net103),
    .A1(\ppu.gfxmode2[7] ),
    .B1(_07565_),
    .X(_00288_));
 sg13g2_o21ai_1 _16036_ (.B1(net239),
    .Y(_07566_),
    .A1(net385),
    .A2(_07556_));
 sg13g2_a21o_1 _16037_ (.A2(_07556_),
    .A1(\ppu.gfxmode2[8] ),
    .B1(_07566_),
    .X(_00289_));
 sg13g2_nand4_1 _16038_ (.B(_02387_),
    .C(_02434_),
    .A(_02378_),
    .Y(_07567_),
    .D(_02477_));
 sg13g2_buf_1 _16039_ (.A(_07567_),
    .X(_07568_));
 sg13g2_buf_1 _16040_ (.A(net118),
    .X(_07569_));
 sg13g2_a21oi_1 _16041_ (.A1(net109),
    .A2(\ppu.gfxmode3[0] ),
    .Y(_07570_),
    .B1(net257));
 sg13g2_o21ai_1 _16042_ (.B1(_07570_),
    .Y(_00290_),
    .A1(net388),
    .A2(net109));
 sg13g2_o21ai_1 _16043_ (.B1(net239),
    .Y(_07571_),
    .A1(_02393_),
    .A2(net118));
 sg13g2_a21o_1 _16044_ (.A2(_07569_),
    .A1(\ppu.gfxmode3[1] ),
    .B1(_07571_),
    .X(_00291_));
 sg13g2_a21oi_1 _16045_ (.A1(net118),
    .A2(\ppu.gfxmode3[2] ),
    .Y(_07572_),
    .B1(net257));
 sg13g2_o21ai_1 _16046_ (.B1(_07572_),
    .Y(_00292_),
    .A1(net339),
    .A2(net109));
 sg13g2_a21oi_1 _16047_ (.A1(net118),
    .A2(\ppu.gfxmode3[3] ),
    .Y(_07573_),
    .B1(net257));
 sg13g2_o21ai_1 _16048_ (.B1(_07573_),
    .Y(_00293_),
    .A1(_02401_),
    .A2(net109));
 sg13g2_a21oi_1 _16049_ (.A1(_07568_),
    .A2(\ppu.gfxmode3[4] ),
    .Y(_07574_),
    .B1(net257));
 sg13g2_o21ai_1 _16050_ (.B1(_07574_),
    .Y(_00294_),
    .A1(_02405_),
    .A2(_07569_));
 sg13g2_a21oi_1 _16051_ (.A1(net118),
    .A2(\ppu.gfxmode3[5] ),
    .Y(_07575_),
    .B1(net257));
 sg13g2_o21ai_1 _16052_ (.B1(_07575_),
    .Y(_00295_),
    .A1(net387),
    .A2(net109));
 sg13g2_inv_1 _16053_ (.Y(_07576_),
    .A(\ppu.gfxmode3[6] ));
 sg13g2_o21ai_1 _16054_ (.B1(net238),
    .Y(_07577_),
    .A1(net406),
    .A2(net118));
 sg13g2_a21oi_1 _16055_ (.A1(_07576_),
    .A2(net109),
    .Y(_00296_),
    .B1(_07577_));
 sg13g2_o21ai_1 _16056_ (.B1(_02220_),
    .Y(_07578_),
    .A1(net386),
    .A2(net118));
 sg13g2_a21o_1 _16057_ (.A2(net109),
    .A1(\ppu.gfxmode3[7] ),
    .B1(_07578_),
    .X(_00297_));
 sg13g2_o21ai_1 _16058_ (.B1(_02220_),
    .Y(_07579_),
    .A1(net385),
    .A2(net118));
 sg13g2_a21o_1 _16059_ (.A2(net109),
    .A1(\ppu.gfxmode3[8] ),
    .B1(_07579_),
    .X(_00298_));
 sg13g2_inv_1 _16060_ (.Y(_07580_),
    .A(\ppu.ram_on ));
 sg13g2_a21oi_1 _16061_ (.A1(_06503_),
    .A2(_07580_),
    .Y(_00427_),
    .B1(net247));
 sg13g2_nand2_1 _16062_ (.Y(_07581_),
    .A(net236),
    .B(\ppu.ram_on ));
 sg13g2_nand2_1 _16063_ (.Y(_07582_),
    .A(_06504_),
    .B(_02526_));
 sg13g2_a21oi_1 _16064_ (.A1(_07581_),
    .A2(_07582_),
    .Y(_00428_),
    .B1(net247));
 sg13g2_inv_1 _16065_ (.Y(_07583_),
    .A(_02267_));
 sg13g2_nor2_2 _16066_ (.A(net347),
    .B(_02199_),
    .Y(_07584_));
 sg13g2_o21ai_1 _16067_ (.B1(_07552_),
    .Y(_07585_),
    .A1(\ppu.rs2.vsync0 ),
    .A2(_07584_));
 sg13g2_a21oi_1 _16068_ (.A1(_07583_),
    .A2(_07584_),
    .Y(_00449_),
    .B1(_07585_));
 sg13g2_nor2_1 _16069_ (.A(\ppu.gfxmode2[3] ),
    .B(net257),
    .Y(_07586_));
 sg13g2_xnor2_1 _16070_ (.Y(_07587_),
    .A(_01836_),
    .B(_06958_));
 sg13g2_a22oi_1 _16071_ (.Y(_00450_),
    .B1(_07587_),
    .B2(_02216_),
    .A2(_07586_),
    .A1(_07584_));
 sg13g2_nor2_1 _16072_ (.A(\ppu.gfxmode2[4] ),
    .B(net258),
    .Y(_07588_));
 sg13g2_xnor2_1 _16073_ (.Y(_07589_),
    .A(_01803_),
    .B(_06954_));
 sg13g2_a22oi_1 _16074_ (.Y(_00451_),
    .B1(_07589_),
    .B2(_02216_),
    .A2(_07588_),
    .A1(_07584_));
 sg13g2_buf_1 _16075_ (.A(_02261_),
    .X(_07590_));
 sg13g2_nor2_1 _16076_ (.A(net347),
    .B(_02200_),
    .Y(_07591_));
 sg13g2_nor3_1 _16077_ (.A(net247),
    .B(_07590_),
    .C(_07591_),
    .Y(_00456_));
 sg13g2_nand2_1 _16078_ (.Y(_07592_),
    .A(_07559_),
    .B(_07562_));
 sg13g2_inv_1 _16079_ (.Y(_07593_),
    .A(_00044_));
 sg13g2_nand2_2 _16080_ (.Y(_07594_),
    .A(_02265_),
    .B(net407));
 sg13g2_inv_1 _16081_ (.Y(_07595_),
    .A(_07594_));
 sg13g2_nor2_2 _16082_ (.A(_07593_),
    .B(_07595_),
    .Y(_07596_));
 sg13g2_inv_1 _16083_ (.Y(_07597_),
    .A(_07596_));
 sg13g2_nor2_1 _16084_ (.A(_07592_),
    .B(_07597_),
    .Y(_07598_));
 sg13g2_inv_1 _16085_ (.Y(_07599_),
    .A(_07598_));
 sg13g2_nor2_1 _16086_ (.A(net407),
    .B(_07599_),
    .Y(_07600_));
 sg13g2_nand2_1 _16087_ (.Y(_07601_),
    .A(_07600_),
    .B(_02265_));
 sg13g2_nor2_2 _16088_ (.A(net341),
    .B(_07595_),
    .Y(_07602_));
 sg13g2_inv_1 _16089_ (.Y(_07603_),
    .A(_07602_));
 sg13g2_nor2_1 _16090_ (.A(_07562_),
    .B(_07560_),
    .Y(_07604_));
 sg13g2_nand2_1 _16091_ (.Y(_07605_),
    .A(_07597_),
    .B(_07604_));
 sg13g2_nand3_1 _16092_ (.B(_07603_),
    .C(_07605_),
    .A(_07599_),
    .Y(_07606_));
 sg13g2_nor2_1 _16093_ (.A(_07604_),
    .B(_07596_),
    .Y(_07607_));
 sg13g2_nand2_1 _16094_ (.Y(_07608_),
    .A(_07607_),
    .B(net407));
 sg13g2_nand4_1 _16095_ (.B(_07606_),
    .C(_07594_),
    .A(_07601_),
    .Y(_07609_),
    .D(_07608_));
 sg13g2_nor2b_1 _16096_ (.A(net122),
    .B_N(_00036_),
    .Y(_07610_));
 sg13g2_a21oi_1 _16097_ (.A1(_07609_),
    .A2(_02259_),
    .Y(_07611_),
    .B1(_07610_));
 sg13g2_o21ai_1 _16098_ (.B1(_07552_),
    .Y(_07612_),
    .A1(_01865_),
    .A2(net165));
 sg13g2_a21oi_1 _16099_ (.A1(net165),
    .A2(_07611_),
    .Y(_00457_),
    .B1(_07612_));
 sg13g2_inv_1 _16100_ (.Y(_07613_),
    .A(_02243_));
 sg13g2_inv_1 _16101_ (.Y(_07614_),
    .A(_02244_));
 sg13g2_nand2_1 _16102_ (.Y(_07615_),
    .A(_02243_),
    .B(_01865_));
 sg13g2_nand2_1 _16103_ (.Y(_07616_),
    .A(_07563_),
    .B(_00044_));
 sg13g2_nand2_1 _16104_ (.Y(_07617_),
    .A(net341),
    .B(_07592_));
 sg13g2_inv_1 _16105_ (.Y(_07618_),
    .A(_07617_));
 sg13g2_inv_1 _16106_ (.Y(_07619_),
    .A(_07592_));
 sg13g2_nor2_1 _16107_ (.A(_07619_),
    .B(_07596_),
    .Y(_07620_));
 sg13g2_inv_1 _16108_ (.Y(_07621_),
    .A(_07620_));
 sg13g2_a21oi_1 _16109_ (.A1(_07560_),
    .A2(_07563_),
    .Y(_07622_),
    .B1(net407));
 sg13g2_nand2_1 _16110_ (.Y(_07623_),
    .A(_07621_),
    .B(_07622_));
 sg13g2_o21ai_1 _16111_ (.B1(_07623_),
    .Y(_07624_),
    .A1(_07594_),
    .A2(_07619_));
 sg13g2_a22oi_1 _16112_ (.Y(_07625_),
    .B1(_02287_),
    .B2(_07624_),
    .A2(_07618_),
    .A1(_07616_));
 sg13g2_a22oi_1 _16113_ (.Y(_07626_),
    .B1(_07625_),
    .B2(net122),
    .A2(_07615_),
    .A1(_07614_));
 sg13g2_o21ai_1 _16114_ (.B1(net238),
    .Y(_07627_),
    .A1(_07626_),
    .A2(net184));
 sg13g2_a21oi_1 _16115_ (.A1(_07613_),
    .A2(net184),
    .Y(_00458_),
    .B1(_07627_));
 sg13g2_nand2_1 _16116_ (.Y(_07628_),
    .A(_07622_),
    .B(_07593_));
 sg13g2_nor2_1 _16117_ (.A(_07559_),
    .B(_07596_),
    .Y(_07629_));
 sg13g2_a21oi_1 _16118_ (.A1(_07629_),
    .A2(_07562_),
    .Y(_07630_),
    .B1(_07598_));
 sg13g2_a22oi_1 _16119_ (.Y(_07631_),
    .B1(_02266_),
    .B2(_07630_),
    .A2(_07628_),
    .A1(_07602_));
 sg13g2_xnor2_1 _16120_ (.Y(_07632_),
    .A(_02246_),
    .B(_02244_));
 sg13g2_o21ai_1 _16121_ (.B1(_07632_),
    .Y(_07633_),
    .A1(_07631_),
    .A2(_02260_));
 sg13g2_o21ai_1 _16122_ (.B1(net239),
    .Y(_07634_),
    .A1(_02245_),
    .A2(net165));
 sg13g2_a21oi_1 _16123_ (.A1(net165),
    .A2(_07633_),
    .Y(_00459_),
    .B1(_07634_));
 sg13g2_a21oi_1 _16124_ (.A1(_02244_),
    .A2(_02246_),
    .Y(_07635_),
    .B1(_02342_));
 sg13g2_nand2_1 _16125_ (.Y(_07636_),
    .A(_07596_),
    .B(_07559_));
 sg13g2_a21oi_1 _16126_ (.A1(_07621_),
    .A2(_07636_),
    .Y(_07637_),
    .B1(_02287_));
 sg13g2_nor2_1 _16127_ (.A(_07603_),
    .B(_07600_),
    .Y(_07638_));
 sg13g2_o21ai_1 _16128_ (.B1(net122),
    .Y(_07639_),
    .A1(_07637_),
    .A2(_07638_));
 sg13g2_o21ai_1 _16129_ (.B1(_07639_),
    .Y(_07640_),
    .A1(_02248_),
    .A2(_07635_));
 sg13g2_a21o_1 _16130_ (.A2(_07640_),
    .A1(net165),
    .B1(_02197_),
    .X(_07641_));
 sg13g2_a21oi_1 _16131_ (.A1(_02342_),
    .A2(_02262_),
    .Y(_00460_),
    .B1(_07641_));
 sg13g2_inv_1 _16132_ (.Y(_07642_),
    .A(_02242_));
 sg13g2_nor2_1 _16133_ (.A(_07642_),
    .B(_02248_),
    .Y(_07643_));
 sg13g2_a21oi_1 _16134_ (.A1(_07560_),
    .A2(_07562_),
    .Y(_07644_),
    .B1(_07594_));
 sg13g2_a221oi_1 _16135_ (.B2(net341),
    .C1(_07644_),
    .B1(_07629_),
    .A1(_02267_),
    .Y(_07645_),
    .A2(_07619_));
 sg13g2_a21oi_1 _16136_ (.A1(net122),
    .A2(_07645_),
    .Y(_07646_),
    .B1(net184));
 sg13g2_o21ai_1 _16137_ (.B1(_07646_),
    .Y(_07647_),
    .A1(_02250_),
    .A2(_07643_));
 sg13g2_nand2_1 _16138_ (.Y(_07648_),
    .A(net184),
    .B(_02242_));
 sg13g2_a21oi_1 _16139_ (.A1(_07647_),
    .A2(_07648_),
    .Y(_00461_),
    .B1(net247));
 sg13g2_inv_1 _16140_ (.Y(_07649_),
    .A(_07629_));
 sg13g2_inv_1 _16141_ (.Y(_07650_),
    .A(_07604_));
 sg13g2_nand3b_1 _16142_ (.B(_07649_),
    .C(_07650_),
    .Y(_07651_),
    .A_N(net407));
 sg13g2_nor2_1 _16143_ (.A(_07602_),
    .B(_07598_),
    .Y(_07652_));
 sg13g2_nand4_1 _16144_ (.B(_07636_),
    .C(net407),
    .A(_07649_),
    .Y(_07653_),
    .D(_07563_));
 sg13g2_a22oi_1 _16145_ (.Y(_07654_),
    .B1(_07652_),
    .B2(_07653_),
    .A2(_07602_),
    .A1(_07651_));
 sg13g2_nand2_1 _16146_ (.Y(_07655_),
    .A(_02251_),
    .B(_02241_));
 sg13g2_a21oi_1 _16147_ (.A1(_02253_),
    .A2(_07655_),
    .Y(_07656_),
    .B1(net122));
 sg13g2_a21oi_1 _16148_ (.A1(net122),
    .A2(_07654_),
    .Y(_07657_),
    .B1(_07656_));
 sg13g2_a21o_1 _16149_ (.A2(_07657_),
    .A1(_02261_),
    .B1(net258),
    .X(_07658_));
 sg13g2_a21oi_1 _16150_ (.A1(_02307_),
    .A2(net184),
    .Y(_00462_),
    .B1(_07658_));
 sg13g2_nor3_1 _16151_ (.A(_00044_),
    .B(_07592_),
    .C(_02287_),
    .Y(_07659_));
 sg13g2_a221oi_1 _16152_ (.B2(_02267_),
    .C1(_07659_),
    .B1(_07607_),
    .A1(_07650_),
    .Y(_07660_),
    .A2(_07644_));
 sg13g2_nor2_1 _16153_ (.A(_07660_),
    .B(_02260_),
    .Y(_07661_));
 sg13g2_nand2_1 _16154_ (.Y(_07662_),
    .A(_02253_),
    .B(_02240_));
 sg13g2_a21oi_1 _16155_ (.A1(_02255_),
    .A2(_07662_),
    .Y(_07663_),
    .B1(net122));
 sg13g2_nor2_1 _16156_ (.A(_07661_),
    .B(_07663_),
    .Y(_07664_));
 sg13g2_o21ai_1 _16157_ (.B1(net239),
    .Y(_07665_),
    .A1(_02240_),
    .A2(net165));
 sg13g2_a21oi_1 _16158_ (.A1(net165),
    .A2(_07664_),
    .Y(_00463_),
    .B1(_07665_));
 sg13g2_o21ai_1 _16159_ (.B1(_02239_),
    .Y(_07666_),
    .A1(_02255_),
    .A2(net184));
 sg13g2_o21ai_1 _16160_ (.B1(_02237_),
    .Y(_07667_),
    .A1(_07559_),
    .A2(_07594_));
 sg13g2_nand3_1 _16161_ (.B(_02256_),
    .C(_07667_),
    .A(_07590_),
    .Y(_07668_));
 sg13g2_a21oi_1 _16162_ (.A1(_07666_),
    .A2(_07668_),
    .Y(_00464_),
    .B1(net247));
 sg13g2_a21oi_1 _16163_ (.A1(net165),
    .A2(_02256_),
    .Y(_07669_),
    .B1(_02321_));
 sg13g2_nand2_1 _16164_ (.Y(_07670_),
    .A(net407),
    .B(_02237_));
 sg13g2_a21oi_1 _16165_ (.A1(_07604_),
    .A2(_02265_),
    .Y(_07671_),
    .B1(_07670_));
 sg13g2_o21ai_1 _16166_ (.B1(_07671_),
    .Y(_07672_),
    .A1(_02265_),
    .A2(_07598_));
 sg13g2_o21ai_1 _16167_ (.B1(_07672_),
    .Y(_07673_),
    .A1(_02321_),
    .A2(_02237_));
 sg13g2_nor3_1 _16168_ (.A(_02257_),
    .B(_07673_),
    .C(net184),
    .Y(_07674_));
 sg13g2_nor3_1 _16169_ (.A(net247),
    .B(_07669_),
    .C(_07674_),
    .Y(_00465_));
 sg13g2_o21ai_1 _16170_ (.B1(net239),
    .Y(_07675_),
    .A1(_02264_),
    .A2(_02263_));
 sg13g2_a21oi_1 _16171_ (.A1(_02263_),
    .A2(_07597_),
    .Y(_00466_),
    .B1(_07675_));
 sg13g2_a21oi_1 _16172_ (.A1(_02263_),
    .A2(_07602_),
    .Y(_07676_),
    .B1(_07548_));
 sg13g2_o21ai_1 _16173_ (.B1(_07676_),
    .Y(_00467_),
    .A1(_02266_),
    .A2(_02263_));
 sg13g2_inv_1 _16174_ (.Y(_07677_),
    .A(_00179_));
 sg13g2_nor2_1 _16175_ (.A(_07677_),
    .B(_02881_),
    .Y(_00504_));
 sg13g2_nor2_1 _16176_ (.A(net235),
    .B(net259),
    .Y(_07678_));
 sg13g2_nor2_1 _16177_ (.A(_02881_),
    .B(_07678_),
    .Y(_00505_));
 sg13g2_nand2_1 _16178_ (.Y(_07679_),
    .A(\ppu.sync_delay[0] ),
    .B(\ppu.sync_delay[1] ));
 sg13g2_xnor2_1 _16179_ (.Y(_07680_),
    .A(\ppu.vsync ),
    .B(_02282_));
 sg13g2_nor3_1 _16180_ (.A(_02274_),
    .B(_07679_),
    .C(_07680_),
    .Y(_07681_));
 sg13g2_o21ai_1 _16181_ (.B1(_07681_),
    .Y(_07682_),
    .A1(hsync),
    .A2(_02280_));
 sg13g2_nand2_1 _16182_ (.Y(_07683_),
    .A(_02288_),
    .B(_02284_));
 sg13g2_a22oi_1 _16183_ (.Y(_07684_),
    .B1(_07683_),
    .B2(_06132_),
    .A2(hsync),
    .A1(_02280_));
 sg13g2_nand2b_1 _16184_ (.Y(_07685_),
    .B(_07684_),
    .A_N(_07682_));
 sg13g2_nand3_1 _16185_ (.B(\ppu.sync_delay[0] ),
    .C(net249),
    .A(_07685_),
    .Y(_00822_));
 sg13g2_nand3b_1 _16186_ (.B(net249),
    .C(_07679_),
    .Y(_00823_),
    .A_N(_02273_));
 sg13g2_o21ai_1 _16187_ (.B1(_02276_),
    .Y(_00824_),
    .A1(_02274_),
    .A2(_02273_));
 sg13g2_nor2_1 _16188_ (.A(net242),
    .B(_07417_),
    .Y(_01085_));
 sg13g2_nor2_1 _16189_ (.A(net242),
    .B(_07419_),
    .Y(_01086_));
 sg13g2_buf_1 _16190_ (.A(net395),
    .X(_07686_));
 sg13g2_nand2_1 _16191_ (.Y(_07687_),
    .A(net348),
    .B(\ppu.sprite_buffer.attr_y[1][12] ));
 sg13g2_o21ai_1 _16192_ (.B1(_07687_),
    .Y(_07688_),
    .A1(net351),
    .A2(_02759_));
 sg13g2_a22oi_1 _16193_ (.Y(_07689_),
    .B1(_07688_),
    .B2(net93),
    .A2(net121),
    .A1(\ppu.base_addr_regs[0][6] ));
 sg13g2_nand2_1 _16194_ (.Y(_07690_),
    .A(net104),
    .B(\ppu.base_addr_regs[1][5] ));
 sg13g2_nand2_1 _16195_ (.Y(_07691_),
    .A(_07689_),
    .B(_07690_));
 sg13g2_buf_1 _16196_ (.A(_02531_),
    .X(_07692_));
 sg13g2_nand2_1 _16197_ (.Y(_07693_),
    .A(_07691_),
    .B(net217));
 sg13g2_buf_1 _16198_ (.A(_02532_),
    .X(_07694_));
 sg13g2_a21oi_1 _16199_ (.A1(net203),
    .A2(\ppu.copper_inst.addr[12] ),
    .Y(_07695_),
    .B1(_01891_));
 sg13g2_nand2_1 _16200_ (.Y(_07696_),
    .A(_07686_),
    .B(\ppu.sprite_buffer.attr_y[1][8] ));
 sg13g2_o21ai_1 _16201_ (.B1(_07696_),
    .Y(_07697_),
    .A1(net351),
    .A2(_02778_));
 sg13g2_nand2_1 _16202_ (.Y(_07698_),
    .A(net93),
    .B(_07697_));
 sg13g2_nand2_1 _16203_ (.Y(_07699_),
    .A(net104),
    .B(\ppu.base_addr_regs[1][1] ));
 sg13g2_a21oi_1 _16204_ (.A1(_02579_),
    .A2(\ppu.base_addr_regs[0][2] ),
    .Y(_07700_),
    .B1(net234));
 sg13g2_nand3_1 _16205_ (.B(_07699_),
    .C(_07700_),
    .A(_07698_),
    .Y(_07701_));
 sg13g2_o21ai_1 _16206_ (.B1(_07701_),
    .Y(_07702_),
    .A1(\ppu.copper_inst.addr[8] ),
    .A2(net217));
 sg13g2_a22oi_1 _16207_ (.Y(_07703_),
    .B1(_02140_),
    .B2(_07702_),
    .A2(_07695_),
    .A1(_07693_));
 sg13g2_a22oi_1 _16208_ (.Y(_07704_),
    .B1(\ppu.sprite_buffer.id_buffer[1][3] ),
    .B2(_02898_),
    .A2(\ppu.sprite_buffer.id_buffer[2][3] ),
    .A1(_02908_));
 sg13g2_a22oi_1 _16209_ (.Y(_07705_),
    .B1(\ppu.sprite_buffer.id_buffer[3][3] ),
    .B2(_02918_),
    .A2(\ppu.sprite_buffer.id_buffer[0][3] ),
    .A1(_02887_));
 sg13g2_nand2_1 _16210_ (.Y(_07706_),
    .A(_07704_),
    .B(_07705_));
 sg13g2_nand2_1 _16211_ (.Y(_07707_),
    .A(net395),
    .B(\ppu.sprite_buffer.attr_y[1][4] ));
 sg13g2_o21ai_1 _16212_ (.B1(_07707_),
    .Y(_07708_),
    .A1(net348),
    .A2(_02770_));
 sg13g2_a22oi_1 _16213_ (.Y(_07709_),
    .B1(_07708_),
    .B2(_06995_),
    .A2(_07706_),
    .A1(_02883_));
 sg13g2_o21ai_1 _16214_ (.B1(_07709_),
    .Y(_07710_),
    .A1(_06966_),
    .A2(_06857_));
 sg13g2_nand2_1 _16215_ (.Y(_07711_),
    .A(_07710_),
    .B(_07692_));
 sg13g2_a21oi_1 _16216_ (.A1(net203),
    .A2(\ppu.copper_inst.addr[4] ),
    .Y(_07712_),
    .B1(_02042_));
 sg13g2_nor2b_1 _16217_ (.A(_06857_),
    .B_N(_00079_),
    .Y(_07713_));
 sg13g2_nor2_1 _16218_ (.A(\ppu.sprite_buffer.oam_req_step ),
    .B(_02884_),
    .Y(_07714_));
 sg13g2_nor2_1 _16219_ (.A(_07713_),
    .B(_07714_),
    .Y(_07715_));
 sg13g2_nand2_1 _16220_ (.Y(_07716_),
    .A(net395),
    .B(\ppu.sprite_buffer.attr_y[1][0] ));
 sg13g2_o21ai_1 _16221_ (.B1(_07716_),
    .Y(_07717_),
    .A1(net395),
    .A2(_02749_));
 sg13g2_xnor2_1 _16222_ (.Y(_07718_),
    .A(_07613_),
    .B(_07717_));
 sg13g2_a21oi_1 _16223_ (.A1(net93),
    .A2(_07718_),
    .Y(_07719_),
    .B1(net234));
 sg13g2_o21ai_1 _16224_ (.B1(net237),
    .Y(_07720_),
    .A1(_00131_),
    .A2(_02531_));
 sg13g2_a21oi_1 _16225_ (.A1(_07715_),
    .A2(_07719_),
    .Y(_07721_),
    .B1(_07720_));
 sg13g2_a21oi_1 _16226_ (.A1(_07711_),
    .A2(_07712_),
    .Y(_07722_),
    .B1(_07721_));
 sg13g2_nand2_1 _16227_ (.Y(_07723_),
    .A(_07703_),
    .B(_07722_));
 sg13g2_inv_1 _16228_ (.Y(_07724_),
    .A(_02585_));
 sg13g2_nand2_1 _16229_ (.Y(_07725_),
    .A(_07723_),
    .B(_07724_));
 sg13g2_buf_1 _16230_ (.A(net343),
    .X(_07726_));
 sg13g2_buf_1 _16231_ (.A(net293),
    .X(_07727_));
 sg13g2_nand2_1 _16232_ (.Y(_07728_),
    .A(net256),
    .B(\ppu.scroll_regs[2][7] ));
 sg13g2_o21ai_1 _16233_ (.B1(_07728_),
    .Y(_07729_),
    .A1(net256),
    .A2(_02621_));
 sg13g2_xnor2_1 _16234_ (.Y(_07730_),
    .A(_00030_),
    .B(_07729_));
 sg13g2_nand2_1 _16235_ (.Y(_07731_),
    .A(_02545_),
    .B(_02534_));
 sg13g2_nand2_1 _16236_ (.Y(_07732_),
    .A(_02533_),
    .B(\ppu.copper_inst.x_cmp[2] ));
 sg13g2_nand2_1 _16237_ (.Y(_07733_),
    .A(_07731_),
    .B(_07732_));
 sg13g2_nand2_1 _16238_ (.Y(_07734_),
    .A(net392),
    .B(\ppu.scroll_regs[2][3] ));
 sg13g2_o21ai_1 _16239_ (.B1(_07734_),
    .Y(_07735_),
    .A1(net392),
    .A2(_02613_));
 sg13g2_xnor2_1 _16240_ (.Y(_07736_),
    .A(_00037_),
    .B(_07735_));
 sg13g2_nand2_1 _16241_ (.Y(_07737_),
    .A(_07733_),
    .B(_07736_));
 sg13g2_nand2_1 _16242_ (.Y(_07738_),
    .A(_07735_),
    .B(_01836_));
 sg13g2_nand2_1 _16243_ (.Y(_07739_),
    .A(_07737_),
    .B(_07738_));
 sg13g2_nand2_1 _16244_ (.Y(_07740_),
    .A(net346),
    .B(\ppu.scroll_regs[2][4] ));
 sg13g2_o21ai_1 _16245_ (.B1(_07740_),
    .Y(_07741_),
    .A1(net346),
    .A2(_02615_));
 sg13g2_xnor2_1 _16246_ (.Y(_07742_),
    .A(_00038_),
    .B(_07741_));
 sg13g2_nand2_1 _16247_ (.Y(_07743_),
    .A(_07739_),
    .B(_07742_));
 sg13g2_nand2_1 _16248_ (.Y(_07744_),
    .A(_07741_),
    .B(_01803_));
 sg13g2_nand2_1 _16249_ (.Y(_07745_),
    .A(_07743_),
    .B(_07744_));
 sg13g2_nand2_1 _16250_ (.Y(_07746_),
    .A(net346),
    .B(\ppu.scroll_regs[2][5] ));
 sg13g2_o21ai_1 _16251_ (.B1(_07746_),
    .Y(_07747_),
    .A1(net346),
    .A2(_02617_));
 sg13g2_xnor2_1 _16252_ (.Y(_07748_),
    .A(_00067_),
    .B(_07747_));
 sg13g2_nand2_1 _16253_ (.Y(_07749_),
    .A(_07745_),
    .B(_07748_));
 sg13g2_nand2_1 _16254_ (.Y(_07750_),
    .A(_07747_),
    .B(_01830_));
 sg13g2_nand2_1 _16255_ (.Y(_07751_),
    .A(_07749_),
    .B(_07750_));
 sg13g2_nand2_1 _16256_ (.Y(_07752_),
    .A(net293),
    .B(\ppu.scroll_regs[2][6] ));
 sg13g2_o21ai_1 _16257_ (.B1(_07752_),
    .Y(_07753_),
    .A1(net293),
    .A2(_02619_));
 sg13g2_xnor2_1 _16258_ (.Y(_07754_),
    .A(_00065_),
    .B(_07753_));
 sg13g2_nand2_1 _16259_ (.Y(_07755_),
    .A(_07751_),
    .B(_07754_));
 sg13g2_nand2_1 _16260_ (.Y(_07756_),
    .A(_07753_),
    .B(_01811_));
 sg13g2_nand2_1 _16261_ (.Y(_07757_),
    .A(_07755_),
    .B(_07756_));
 sg13g2_xnor2_1 _16262_ (.Y(_07758_),
    .A(_07730_),
    .B(_07757_));
 sg13g2_xor2_1 _16263_ (.B(_07733_),
    .A(_07736_),
    .X(_07759_));
 sg13g2_a21oi_1 _16264_ (.A1(_07759_),
    .A2(net266),
    .Y(_07760_),
    .B1(_01854_));
 sg13g2_o21ai_1 _16265_ (.B1(_07760_),
    .Y(_07761_),
    .A1(net266),
    .A2(_07758_));
 sg13g2_nand2_1 _16266_ (.Y(_07762_),
    .A(net293),
    .B(\ppu.scroll_regs[3][5] ));
 sg13g2_o21ai_1 _16267_ (.B1(_07762_),
    .Y(_07763_),
    .A1(net293),
    .A2(_02638_));
 sg13g2_xnor2_1 _16268_ (.Y(_07764_),
    .A(_02240_),
    .B(_07763_));
 sg13g2_nand2_1 _16269_ (.Y(_07765_),
    .A(net392),
    .B(\ppu.scroll_regs[3][3] ));
 sg13g2_o21ai_1 _16270_ (.B1(_07765_),
    .Y(_07766_),
    .A1(net346),
    .A2(_02634_));
 sg13g2_xnor2_1 _16271_ (.Y(_07767_),
    .A(_02242_),
    .B(_07766_));
 sg13g2_inv_1 _16272_ (.Y(_07768_),
    .A(_07767_));
 sg13g2_nand2_1 _16273_ (.Y(_07769_),
    .A(_01821_),
    .B(\ppu.scroll_regs[3][1] ));
 sg13g2_o21ai_1 _16274_ (.B1(_07769_),
    .Y(_07770_),
    .A1(net392),
    .A2(_02630_));
 sg13g2_xnor2_1 _16275_ (.Y(_07771_),
    .A(_02245_),
    .B(_07770_));
 sg13g2_nor2b_1 _16276_ (.A(net392),
    .B_N(\ppu.scroll_regs[1][0] ),
    .Y(_07772_));
 sg13g2_a21oi_1 _16277_ (.A1(_01822_),
    .A2(\ppu.scroll_regs[3][0] ),
    .Y(_07773_),
    .B1(_07772_));
 sg13g2_nor2_1 _16278_ (.A(_02243_),
    .B(_07773_),
    .Y(_07774_));
 sg13g2_nor2b_1 _16279_ (.A(_02245_),
    .B_N(_07770_),
    .Y(_07775_));
 sg13g2_a21oi_1 _16280_ (.A1(_07771_),
    .A2(_07774_),
    .Y(_07776_),
    .B1(_07775_));
 sg13g2_nand2_1 _16281_ (.Y(_07777_),
    .A(_01822_),
    .B(\ppu.scroll_regs[3][2] ));
 sg13g2_o21ai_1 _16282_ (.B1(_07777_),
    .Y(_07778_),
    .A1(net346),
    .A2(_02632_));
 sg13g2_nand2_1 _16283_ (.Y(_07779_),
    .A(_07778_),
    .B(_02342_));
 sg13g2_nor2_1 _16284_ (.A(_02342_),
    .B(_07778_),
    .Y(_07780_));
 sg13g2_a21o_1 _16285_ (.A2(_07779_),
    .A1(_07776_),
    .B1(_07780_),
    .X(_07781_));
 sg13g2_nor2_1 _16286_ (.A(_07768_),
    .B(_07781_),
    .Y(_07782_));
 sg13g2_nand2_1 _16287_ (.Y(_07783_),
    .A(_07766_),
    .B(_07642_));
 sg13g2_nor2b_1 _16288_ (.A(_07782_),
    .B_N(_07783_),
    .Y(_07784_));
 sg13g2_nand2_1 _16289_ (.Y(_07785_),
    .A(_01823_),
    .B(\ppu.scroll_regs[3][4] ));
 sg13g2_o21ai_1 _16290_ (.B1(_07785_),
    .Y(_07786_),
    .A1(_01823_),
    .A2(_02636_));
 sg13g2_nand2_1 _16291_ (.Y(_07787_),
    .A(_07786_),
    .B(_02307_));
 sg13g2_nor2_1 _16292_ (.A(_02307_),
    .B(_07786_),
    .Y(_07788_));
 sg13g2_a21oi_1 _16293_ (.A1(_07784_),
    .A2(_07787_),
    .Y(_07789_),
    .B1(_07788_));
 sg13g2_xnor2_1 _16294_ (.Y(_07790_),
    .A(_07764_),
    .B(_07789_));
 sg13g2_nand2_1 _16295_ (.Y(_07791_),
    .A(_07790_),
    .B(_07726_));
 sg13g2_a21oi_1 _16296_ (.A1(_02209_),
    .A2(\ppu.base_addr_regs[2][1] ),
    .Y(_07792_),
    .B1(net266));
 sg13g2_o21ai_1 _16297_ (.B1(_07792_),
    .Y(_07793_),
    .A1(_02209_),
    .A2(_02444_));
 sg13g2_a21o_1 _16298_ (.A2(_07793_),
    .A1(_07791_),
    .B1(net294),
    .X(_07794_));
 sg13g2_nand3_1 _16299_ (.B(_02583_),
    .C(_07794_),
    .A(_07761_),
    .Y(_07795_));
 sg13g2_inv_1 _16300_ (.Y(_07796_),
    .A(_00159_));
 sg13g2_xnor2_1 _16301_ (.Y(_07797_),
    .A(_07796_),
    .B(_07773_));
 sg13g2_o21ai_1 _16302_ (.B1(net295),
    .Y(_07798_),
    .A1(_02810_),
    .A2(net216));
 sg13g2_a21oi_1 _16303_ (.A1(_07797_),
    .A2(net216),
    .Y(_07799_),
    .B1(_07798_));
 sg13g2_nor2_1 _16304_ (.A(_07799_),
    .B(_07724_),
    .Y(_07800_));
 sg13g2_inv_1 _16305_ (.Y(_07801_),
    .A(_02526_));
 sg13g2_a21oi_1 _16306_ (.A1(_07795_),
    .A2(_07800_),
    .Y(_07802_),
    .B1(_07801_));
 sg13g2_nand2_1 _16307_ (.Y(_07803_),
    .A(_07725_),
    .B(_07802_));
 sg13g2_nor2_1 _16308_ (.A(_02526_),
    .B(_07580_),
    .Y(_07804_));
 sg13g2_a21oi_1 _16309_ (.A1(net216),
    .A2(_07804_),
    .Y(_07805_),
    .B1(net258));
 sg13g2_nor2_1 _16310_ (.A(net405),
    .B(net249),
    .Y(_07806_));
 sg13g2_a21oi_1 _16311_ (.A1(_07803_),
    .A2(_07805_),
    .Y(\addr_pins_out[0] ),
    .B1(_07806_));
 sg13g2_nand2_1 _16312_ (.Y(_07807_),
    .A(net256),
    .B(\ppu.scroll_regs[2][8] ));
 sg13g2_o21ai_1 _16313_ (.B1(_07807_),
    .Y(_07808_),
    .A1(net256),
    .A2(_02623_));
 sg13g2_xor2_1 _16314_ (.B(_07808_),
    .A(_01827_),
    .X(_07809_));
 sg13g2_a22oi_1 _16315_ (.Y(_07810_),
    .B1(_07730_),
    .B2(_07757_),
    .A2(_07729_),
    .A1(_02075_));
 sg13g2_xnor2_1 _16316_ (.Y(_07811_),
    .A(_07809_),
    .B(_07810_));
 sg13g2_xnor2_1 _16317_ (.Y(_07812_),
    .A(_07742_),
    .B(_07739_));
 sg13g2_nand2_1 _16318_ (.Y(_07813_),
    .A(_07812_),
    .B(net343));
 sg13g2_o21ai_1 _16319_ (.B1(_07813_),
    .Y(_07814_),
    .A1(net266),
    .A2(_07811_));
 sg13g2_nand2_1 _16320_ (.Y(_07815_),
    .A(_07814_),
    .B(net294));
 sg13g2_nand2_1 _16321_ (.Y(_07816_),
    .A(net293),
    .B(\ppu.scroll_regs[3][6] ));
 sg13g2_o21ai_1 _16322_ (.B1(_07816_),
    .Y(_07817_),
    .A1(net293),
    .A2(_02640_));
 sg13g2_xnor2_1 _16323_ (.Y(_07818_),
    .A(_02239_),
    .B(_07817_));
 sg13g2_nand2_1 _16324_ (.Y(_07819_),
    .A(_07789_),
    .B(_07764_));
 sg13g2_nand2b_1 _16325_ (.Y(_07820_),
    .B(_07763_),
    .A_N(_02240_));
 sg13g2_nand2_1 _16326_ (.Y(_07821_),
    .A(_07819_),
    .B(_07820_));
 sg13g2_xnor2_1 _16327_ (.Y(_07822_),
    .A(_07818_),
    .B(_07821_));
 sg13g2_nand2_1 _16328_ (.Y(_07823_),
    .A(_07822_),
    .B(_07726_));
 sg13g2_a21oi_1 _16329_ (.A1(_02209_),
    .A2(\ppu.base_addr_regs[2][2] ),
    .Y(_07824_),
    .B1(net343));
 sg13g2_o21ai_1 _16330_ (.B1(_07824_),
    .Y(_07825_),
    .A1(_02209_),
    .A2(_02446_));
 sg13g2_a21o_1 _16331_ (.A2(_07825_),
    .A1(_07823_),
    .B1(net294),
    .X(_07826_));
 sg13g2_nand3_1 _16332_ (.B(_02583_),
    .C(_07826_),
    .A(_07815_),
    .Y(_07827_));
 sg13g2_xor2_1 _16333_ (.B(_07771_),
    .A(_07774_),
    .X(_07828_));
 sg13g2_a21oi_1 _16334_ (.A1(_06535_),
    .A2(net262),
    .Y(_07829_),
    .B1(_02583_));
 sg13g2_o21ai_1 _16335_ (.B1(_07829_),
    .Y(_07830_),
    .A1(net262),
    .A2(_07828_));
 sg13g2_nand2_1 _16336_ (.Y(_07831_),
    .A(_07827_),
    .B(_07830_));
 sg13g2_nand2_1 _16337_ (.Y(_07832_),
    .A(_07831_),
    .B(_02585_));
 sg13g2_a22oi_1 _16338_ (.Y(_07833_),
    .B1(\ppu.sprite_buffer.id_buffer[3][0] ),
    .B2(_02918_),
    .A2(\ppu.sprite_buffer.id_buffer[0][0] ),
    .A1(_02887_));
 sg13g2_a22oi_1 _16339_ (.Y(_07834_),
    .B1(\ppu.sprite_buffer.id_buffer[1][0] ),
    .B2(_02898_),
    .A2(\ppu.sprite_buffer.id_buffer[2][0] ),
    .A1(_02908_));
 sg13g2_nand3_1 _16340_ (.B(_07833_),
    .C(_07834_),
    .A(net104),
    .Y(_07835_));
 sg13g2_nand2_1 _16341_ (.Y(_07836_),
    .A(_07717_),
    .B(_07796_));
 sg13g2_nand2_1 _16342_ (.Y(_07837_),
    .A(_06999_),
    .B(\ppu.sprite_buffer.attr_y[1][1] ));
 sg13g2_o21ai_1 _16343_ (.B1(_07837_),
    .Y(_07838_),
    .A1(net395),
    .A2(_02766_));
 sg13g2_xnor2_1 _16344_ (.Y(_07839_),
    .A(_02246_),
    .B(_07838_));
 sg13g2_xnor2_1 _16345_ (.Y(_07840_),
    .A(_07836_),
    .B(_07839_));
 sg13g2_nand2_1 _16346_ (.Y(_07841_),
    .A(net93),
    .B(_07840_));
 sg13g2_a21oi_1 _16347_ (.A1(net121),
    .A2(_00078_),
    .Y(_07842_),
    .B1(net234));
 sg13g2_nand3_1 _16348_ (.B(_07841_),
    .C(_07842_),
    .A(_07835_),
    .Y(_07843_));
 sg13g2_inv_1 _16349_ (.Y(_07844_),
    .A(_00132_));
 sg13g2_a21oi_1 _16350_ (.A1(net203),
    .A2(_07844_),
    .Y(_07845_),
    .B1(_01921_));
 sg13g2_nand2_1 _16351_ (.Y(_07846_),
    .A(net348),
    .B(\ppu.sprite_buffer.attr_y[1][9] ));
 sg13g2_o21ai_1 _16352_ (.B1(_07846_),
    .Y(_07847_),
    .A1(_07000_),
    .A2(_02780_));
 sg13g2_nand2_1 _16353_ (.Y(_07848_),
    .A(_06995_),
    .B(_07847_));
 sg13g2_nand2_1 _16354_ (.Y(_07849_),
    .A(_02883_),
    .B(\ppu.base_addr_regs[1][2] ));
 sg13g2_a21oi_1 _16355_ (.A1(_02579_),
    .A2(\ppu.base_addr_regs[0][3] ),
    .Y(_07850_),
    .B1(net234));
 sg13g2_nand3_1 _16356_ (.B(_07849_),
    .C(_07850_),
    .A(_07848_),
    .Y(_07851_));
 sg13g2_nand2_1 _16357_ (.Y(_07852_),
    .A(net203),
    .B(_06870_));
 sg13g2_nand2_1 _16358_ (.Y(_07853_),
    .A(_07851_),
    .B(_07852_));
 sg13g2_a22oi_1 _16359_ (.Y(_07854_),
    .B1(net259),
    .B2(_07853_),
    .A2(_07845_),
    .A1(_07843_));
 sg13g2_nand2_1 _16360_ (.Y(_07855_),
    .A(net348),
    .B(\ppu.sprite_buffer.attr_y[1][13] ));
 sg13g2_o21ai_1 _16361_ (.B1(_07855_),
    .Y(_07856_),
    .A1(_07000_),
    .A2(_02762_));
 sg13g2_a22oi_1 _16362_ (.Y(_07857_),
    .B1(_07856_),
    .B2(net93),
    .A2(net121),
    .A1(\ppu.base_addr_regs[0][7] ));
 sg13g2_nand2_1 _16363_ (.Y(_07858_),
    .A(net104),
    .B(\ppu.base_addr_regs[1][6] ));
 sg13g2_a21oi_1 _16364_ (.A1(_07857_),
    .A2(_07858_),
    .Y(_07859_),
    .B1(net203));
 sg13g2_a21oi_1 _16365_ (.A1(net203),
    .A2(\ppu.copper_inst.addr[13] ),
    .Y(_07860_),
    .B1(_01891_));
 sg13g2_nand2b_1 _16366_ (.Y(_07861_),
    .B(_07860_),
    .A_N(_07859_));
 sg13g2_a22oi_1 _16367_ (.Y(_07862_),
    .B1(\ppu.sprite_buffer.id_buffer[1][4] ),
    .B2(_02898_),
    .A2(\ppu.sprite_buffer.id_buffer[3][4] ),
    .A1(_02918_));
 sg13g2_a22oi_1 _16368_ (.Y(_07863_),
    .B1(\ppu.sprite_buffer.id_buffer[2][4] ),
    .B2(_02908_),
    .A2(\ppu.sprite_buffer.id_buffer[0][4] ),
    .A1(_02887_));
 sg13g2_nand2_1 _16369_ (.Y(_07864_),
    .A(_07862_),
    .B(_07863_));
 sg13g2_a22oi_1 _16370_ (.Y(_07865_),
    .B1(_07864_),
    .B2(_02883_),
    .A2(_02579_),
    .A1(\ppu.sprite_buffer.extra_sorted_addr_bits[2] ));
 sg13g2_nand2_1 _16371_ (.Y(_07866_),
    .A(_06999_),
    .B(\ppu.sprite_buffer.attr_y[1][5] ));
 sg13g2_o21ai_1 _16372_ (.B1(_07866_),
    .Y(_07867_),
    .A1(net348),
    .A2(_02772_));
 sg13g2_nand2_1 _16373_ (.Y(_07868_),
    .A(_06995_),
    .B(_07867_));
 sg13g2_nand2_1 _16374_ (.Y(_07869_),
    .A(_07865_),
    .B(_07868_));
 sg13g2_nand2_1 _16375_ (.Y(_07870_),
    .A(_07869_),
    .B(_07692_));
 sg13g2_a21oi_1 _16376_ (.A1(_07694_),
    .A2(\ppu.copper_inst.addr[5] ),
    .Y(_07871_),
    .B1(_02042_));
 sg13g2_a21oi_1 _16377_ (.A1(_07870_),
    .A2(_07871_),
    .Y(_07872_),
    .B1(_02585_));
 sg13g2_nand3_1 _16378_ (.B(_07861_),
    .C(_07872_),
    .A(_07854_),
    .Y(_07873_));
 sg13g2_nand2_1 _16379_ (.Y(_07874_),
    .A(_07832_),
    .B(_07873_));
 sg13g2_nand2_1 _16380_ (.Y(_07875_),
    .A(_07874_),
    .B(_02526_));
 sg13g2_a21oi_1 _16381_ (.A1(net235),
    .A2(_07804_),
    .Y(_07876_),
    .B1(net258));
 sg13g2_nor2_1 _16382_ (.A(net403),
    .B(net249),
    .Y(_07877_));
 sg13g2_a21oi_1 _16383_ (.A1(_07875_),
    .A2(_07876_),
    .Y(\addr_pins_out[1] ),
    .B1(_07877_));
 sg13g2_a21oi_1 _16384_ (.A1(net251),
    .A2(_07804_),
    .Y(_07878_),
    .B1(_07548_));
 sg13g2_a22oi_1 _16385_ (.Y(_07879_),
    .B1(\ppu.base_addr_regs[1][7] ),
    .B2(net104),
    .A2(net121),
    .A1(\ppu.base_addr_regs[0][8] ));
 sg13g2_nand2_1 _16386_ (.Y(_07880_),
    .A(_06995_),
    .B(\ppu.base_addr_regs[3][3] ));
 sg13g2_nand2_1 _16387_ (.Y(_07881_),
    .A(_07879_),
    .B(_07880_));
 sg13g2_o21ai_1 _16388_ (.B1(net254),
    .Y(_07882_),
    .A1(_06914_),
    .A2(_02531_));
 sg13g2_a21oi_1 _16389_ (.A1(_07881_),
    .A2(net217),
    .Y(_07883_),
    .B1(_07882_));
 sg13g2_a22oi_1 _16390_ (.Y(_07884_),
    .B1(\ppu.sprite_buffer.id_buffer[1][1] ),
    .B2(_02898_),
    .A2(\ppu.sprite_buffer.id_buffer[2][1] ),
    .A1(_02908_));
 sg13g2_a22oi_1 _16391_ (.Y(_07885_),
    .B1(\ppu.sprite_buffer.id_buffer[3][1] ),
    .B2(_02918_),
    .A2(\ppu.sprite_buffer.id_buffer[0][1] ),
    .A1(_02887_));
 sg13g2_nand2_1 _16392_ (.Y(_07886_),
    .A(_07884_),
    .B(_07885_));
 sg13g2_a22oi_1 _16393_ (.Y(_07887_),
    .B1(_07886_),
    .B2(net104),
    .A2(_02580_),
    .A1(\ppu.sprite_buffer.out_counters[0][2] ));
 sg13g2_nand2_1 _16394_ (.Y(_07888_),
    .A(net395),
    .B(\ppu.sprite_buffer.attr_y[1][2] ));
 sg13g2_o21ai_1 _16395_ (.B1(_07888_),
    .Y(_07889_),
    .A1(net395),
    .A2(_02768_));
 sg13g2_xnor2_1 _16396_ (.Y(_07890_),
    .A(_02342_),
    .B(_07889_));
 sg13g2_nor2_1 _16397_ (.A(_02245_),
    .B(_07838_),
    .Y(_07891_));
 sg13g2_a21oi_1 _16398_ (.A1(_07839_),
    .A2(_07836_),
    .Y(_07892_),
    .B1(_07891_));
 sg13g2_xnor2_1 _16399_ (.Y(_07893_),
    .A(_07890_),
    .B(_07892_));
 sg13g2_nand2_1 _16400_ (.Y(_07894_),
    .A(net93),
    .B(_07893_));
 sg13g2_nand2_1 _16401_ (.Y(_07895_),
    .A(_07887_),
    .B(_07894_));
 sg13g2_o21ai_1 _16402_ (.B1(_02481_),
    .Y(_07896_),
    .A1(_06873_),
    .A2(_02531_));
 sg13g2_a21oi_1 _16403_ (.A1(_07895_),
    .A2(net217),
    .Y(_07897_),
    .B1(_07896_));
 sg13g2_nor2_1 _16404_ (.A(_07883_),
    .B(_07897_),
    .Y(_07898_));
 sg13g2_a22oi_1 _16405_ (.Y(_07899_),
    .B1(\ppu.sprite_buffer.id_buffer[1][5] ),
    .B2(_02898_),
    .A2(\ppu.sprite_buffer.id_buffer[2][5] ),
    .A1(_02908_));
 sg13g2_a22oi_1 _16406_ (.Y(_07900_),
    .B1(\ppu.sprite_buffer.id_buffer[3][5] ),
    .B2(_02918_),
    .A2(\ppu.sprite_buffer.id_buffer[0][5] ),
    .A1(_02887_));
 sg13g2_nand2_1 _16407_ (.Y(_07901_),
    .A(_07899_),
    .B(_07900_));
 sg13g2_a22oi_1 _16408_ (.Y(_07902_),
    .B1(_07901_),
    .B2(net104),
    .A2(_02580_),
    .A1(\ppu.base_addr_regs[0][0] ));
 sg13g2_nand2_1 _16409_ (.Y(_07903_),
    .A(_07686_),
    .B(\ppu.sprite_buffer.attr_y[1][6] ));
 sg13g2_o21ai_1 _16410_ (.B1(_07903_),
    .Y(_07904_),
    .A1(net351),
    .A2(_02774_));
 sg13g2_nand2_1 _16411_ (.Y(_07905_),
    .A(_06996_),
    .B(_07904_));
 sg13g2_nand2_1 _16412_ (.Y(_07906_),
    .A(_07902_),
    .B(_07905_));
 sg13g2_nand2_1 _16413_ (.Y(_07907_),
    .A(_07906_),
    .B(net217));
 sg13g2_a21oi_1 _16414_ (.A1(_07694_),
    .A2(\ppu.copper_inst.addr[6] ),
    .Y(_07908_),
    .B1(_02042_));
 sg13g2_a21oi_1 _16415_ (.A1(_07907_),
    .A2(_07908_),
    .Y(_07909_),
    .B1(_02585_));
 sg13g2_nand2_1 _16416_ (.Y(_07910_),
    .A(net348),
    .B(\ppu.sprite_buffer.attr_y[1][10] ));
 sg13g2_o21ai_1 _16417_ (.B1(_07910_),
    .Y(_07911_),
    .A1(net351),
    .A2(_02755_));
 sg13g2_nand2_1 _16418_ (.Y(_07912_),
    .A(net93),
    .B(_07911_));
 sg13g2_nand2_1 _16419_ (.Y(_07913_),
    .A(_06989_),
    .B(\ppu.base_addr_regs[1][3] ));
 sg13g2_a21oi_1 _16420_ (.A1(net121),
    .A2(\ppu.base_addr_regs[0][4] ),
    .Y(_07914_),
    .B1(net234));
 sg13g2_nand3_1 _16421_ (.B(_07913_),
    .C(_07914_),
    .A(_07912_),
    .Y(_07915_));
 sg13g2_o21ai_1 _16422_ (.B1(_07915_),
    .Y(_07916_),
    .A1(_06864_),
    .A2(net217));
 sg13g2_nand2_1 _16423_ (.Y(_07917_),
    .A(_07916_),
    .B(_02140_));
 sg13g2_nand3_1 _16424_ (.B(_07909_),
    .C(_07917_),
    .A(_07898_),
    .Y(_07918_));
 sg13g2_nor2b_1 _16425_ (.A(_02239_),
    .B_N(_07817_),
    .Y(_07919_));
 sg13g2_nand2_1 _16426_ (.Y(_07920_),
    .A(_07821_),
    .B(_07818_));
 sg13g2_nand2b_1 _16427_ (.Y(_07921_),
    .B(_07920_),
    .A_N(_07919_));
 sg13g2_nand2_1 _16428_ (.Y(_07922_),
    .A(_03247_),
    .B(\ppu.scroll_regs[3][7] ));
 sg13g2_o21ai_1 _16429_ (.B1(_07922_),
    .Y(_07923_),
    .A1(_03247_),
    .A2(_02642_));
 sg13g2_xnor2_1 _16430_ (.Y(_07924_),
    .A(_02321_),
    .B(_07923_));
 sg13g2_nand2b_1 _16431_ (.Y(_07925_),
    .B(_07924_),
    .A_N(_07921_));
 sg13g2_inv_1 _16432_ (.Y(_07926_),
    .A(_07924_));
 sg13g2_nand2_1 _16433_ (.Y(_07927_),
    .A(_07921_),
    .B(_07926_));
 sg13g2_nand3_1 _16434_ (.B(net266),
    .C(_07927_),
    .A(_07925_),
    .Y(_07928_));
 sg13g2_a21oi_1 _16435_ (.A1(net256),
    .A2(\ppu.base_addr_regs[2][7] ),
    .Y(_07929_),
    .B1(net266));
 sg13g2_o21ai_1 _16436_ (.B1(_07929_),
    .Y(_07930_),
    .A1(net256),
    .A2(_02440_));
 sg13g2_a21oi_1 _16437_ (.A1(_07928_),
    .A2(_07930_),
    .Y(_07931_),
    .B1(net294));
 sg13g2_xnor2_1 _16438_ (.Y(_07932_),
    .A(_07768_),
    .B(_07781_));
 sg13g2_xnor2_1 _16439_ (.Y(_07933_),
    .A(_07748_),
    .B(_07745_));
 sg13g2_a22oi_1 _16440_ (.Y(_07934_),
    .B1(net216),
    .B2(_07933_),
    .A2(_07932_),
    .A1(net235));
 sg13g2_nor2b_1 _16441_ (.A(_07931_),
    .B_N(_07934_),
    .Y(_07935_));
 sg13g2_nor2b_1 _16442_ (.A(_07678_),
    .B_N(_02816_),
    .Y(_07936_));
 sg13g2_nor2_1 _16443_ (.A(_02450_),
    .B(net297),
    .Y(_07937_));
 sg13g2_nand2b_1 _16444_ (.Y(_07938_),
    .B(_07779_),
    .A_N(_07780_));
 sg13g2_o21ai_1 _16445_ (.B1(net237),
    .Y(_07939_),
    .A1(_07938_),
    .A2(_07776_));
 sg13g2_a21oi_1 _16446_ (.A1(_07776_),
    .A2(_07938_),
    .Y(_07940_),
    .B1(_07939_));
 sg13g2_nor4_1 _16447_ (.A(_02583_),
    .B(_07936_),
    .C(_07937_),
    .D(_07940_),
    .Y(_07941_));
 sg13g2_nor2_1 _16448_ (.A(_07941_),
    .B(_07724_),
    .Y(_07942_));
 sg13g2_o21ai_1 _16449_ (.B1(_07942_),
    .Y(_07943_),
    .A1(net295),
    .A2(_07935_));
 sg13g2_nand2_1 _16450_ (.Y(_07944_),
    .A(_07918_),
    .B(_07943_));
 sg13g2_nand2_1 _16451_ (.Y(_07945_),
    .A(_07944_),
    .B(_02526_));
 sg13g2_a22oi_1 _16452_ (.Y(\addr_pins_out[2] ),
    .B1(_07878_),
    .B2(_07945_),
    .A2(net247),
    .A1(_02686_));
 sg13g2_a22oi_1 _16453_ (.Y(_07946_),
    .B1(\ppu.sprite_buffer.id_buffer[1][2] ),
    .B2(_02898_),
    .A2(\ppu.sprite_buffer.id_buffer[3][2] ),
    .A1(_02918_));
 sg13g2_a22oi_1 _16454_ (.Y(_07947_),
    .B1(\ppu.sprite_buffer.id_buffer[2][2] ),
    .B2(_02908_),
    .A2(\ppu.sprite_buffer.id_buffer[0][2] ),
    .A1(_02887_));
 sg13g2_a21oi_1 _16455_ (.A1(_07946_),
    .A2(_07947_),
    .Y(_07948_),
    .B1(_02884_));
 sg13g2_inv_1 _16456_ (.Y(_07949_),
    .A(_00160_));
 sg13g2_a22oi_1 _16457_ (.Y(_07950_),
    .B1(_07949_),
    .B2(net93),
    .A2(net121),
    .A1(_02866_));
 sg13g2_nand2b_1 _16458_ (.Y(_07951_),
    .B(_07950_),
    .A_N(_07948_));
 sg13g2_o21ai_1 _16459_ (.B1(_02481_),
    .Y(_07952_),
    .A1(_06875_),
    .A2(_02531_));
 sg13g2_a21oi_1 _16460_ (.A1(_07951_),
    .A2(net217),
    .Y(_07953_),
    .B1(_07952_));
 sg13g2_nor2_1 _16461_ (.A(_06885_),
    .B(_02531_),
    .Y(_07954_));
 sg13g2_nand2_1 _16462_ (.Y(_07955_),
    .A(net348),
    .B(\ppu.sprite_buffer.attr_y[1][11] ));
 sg13g2_o21ai_1 _16463_ (.B1(_07955_),
    .Y(_07956_),
    .A1(net351),
    .A2(_02757_));
 sg13g2_a22oi_1 _16464_ (.Y(_07957_),
    .B1(_07956_),
    .B2(_06995_),
    .A2(net121),
    .A1(\ppu.base_addr_regs[0][5] ));
 sg13g2_nand2_1 _16465_ (.Y(_07958_),
    .A(_06989_),
    .B(\ppu.base_addr_regs[1][4] ));
 sg13g2_a21oi_1 _16466_ (.A1(_07957_),
    .A2(_07958_),
    .Y(_07959_),
    .B1(net203));
 sg13g2_nor3_1 _16467_ (.A(_02028_),
    .B(_07954_),
    .C(_07959_),
    .Y(_07960_));
 sg13g2_nor2_1 _16468_ (.A(_07953_),
    .B(_07960_),
    .Y(_07961_));
 sg13g2_a22oi_1 _16469_ (.Y(_07962_),
    .B1(\ppu.base_addr_regs[3][4] ),
    .B2(_06995_),
    .A2(\ppu.base_addr_regs[1][8] ),
    .A1(_02883_));
 sg13g2_a21oi_1 _16470_ (.A1(net234),
    .A2(\ppu.copper_inst.addr[15] ),
    .Y(_07963_),
    .B1(net297));
 sg13g2_o21ai_1 _16471_ (.B1(_07963_),
    .Y(_07964_),
    .A1(net203),
    .A2(_07962_));
 sg13g2_nand2_1 _16472_ (.Y(_07965_),
    .A(_07964_),
    .B(_07724_));
 sg13g2_inv_1 _16473_ (.Y(_07966_),
    .A(\ppu.base_addr_regs[0][1] ));
 sg13g2_nand2_1 _16474_ (.Y(_07967_),
    .A(net348),
    .B(\ppu.sprite_buffer.attr_y[1][7] ));
 sg13g2_o21ai_1 _16475_ (.B1(_07967_),
    .Y(_07968_),
    .A1(net351),
    .A2(_02776_));
 sg13g2_a22oi_1 _16476_ (.Y(_07969_),
    .B1(_07968_),
    .B2(_06995_),
    .A2(\ppu.base_addr_regs[1][0] ),
    .A1(_02883_));
 sg13g2_o21ai_1 _16477_ (.B1(_07969_),
    .Y(_07970_),
    .A1(_07966_),
    .A2(_06857_));
 sg13g2_o21ai_1 _16478_ (.B1(_02501_),
    .Y(_07971_),
    .A1(_06868_),
    .A2(_02531_));
 sg13g2_a21oi_1 _16479_ (.A1(_07970_),
    .A2(net217),
    .Y(_07972_),
    .B1(_07971_));
 sg13g2_nor2_1 _16480_ (.A(_07965_),
    .B(_07972_),
    .Y(_07973_));
 sg13g2_nand2_1 _16481_ (.Y(_07974_),
    .A(_07961_),
    .B(_07973_));
 sg13g2_xor2_1 _16482_ (.B(_07751_),
    .A(_07754_),
    .X(_07975_));
 sg13g2_nor2b_1 _16483_ (.A(_07788_),
    .B_N(_07787_),
    .Y(_07976_));
 sg13g2_nor2b_1 _16484_ (.A(_07784_),
    .B_N(_07976_),
    .Y(_07977_));
 sg13g2_nor2b_1 _16485_ (.A(_07976_),
    .B_N(_07784_),
    .Y(_07978_));
 sg13g2_o21ai_1 _16486_ (.B1(_06222_),
    .Y(_07979_),
    .A1(_07977_),
    .A2(_07978_));
 sg13g2_o21ai_1 _16487_ (.B1(_07979_),
    .Y(_07980_),
    .A1(_06222_),
    .A2(_07975_));
 sg13g2_a21o_1 _16488_ (.A2(_03085_),
    .A1(_07980_),
    .B1(_02576_),
    .X(_07981_));
 sg13g2_nor2b_1 _16489_ (.A(net256),
    .B_N(\ppu.scroll_regs[1][8] ),
    .Y(_07982_));
 sg13g2_a21oi_1 _16490_ (.A1(_07727_),
    .A2(\ppu.scroll_regs[3][8] ),
    .Y(_07983_),
    .B1(_07982_));
 sg13g2_a22oi_1 _16491_ (.Y(_07984_),
    .B1(_07919_),
    .B2(_07924_),
    .A2(_07923_),
    .A1(_02237_));
 sg13g2_o21ai_1 _16492_ (.B1(_07984_),
    .Y(_07985_),
    .A1(_07926_),
    .A2(_07920_));
 sg13g2_nor2_1 _16493_ (.A(_07983_),
    .B(_07985_),
    .Y(_07986_));
 sg13g2_nand2_1 _16494_ (.Y(_07987_),
    .A(_07985_),
    .B(_07983_));
 sg13g2_nand3b_1 _16495_ (.B(net266),
    .C(_07987_),
    .Y(_07988_),
    .A_N(_07986_));
 sg13g2_a21oi_1 _16496_ (.A1(net256),
    .A2(\ppu.base_addr_regs[2][8] ),
    .Y(_07989_),
    .B1(net266));
 sg13g2_o21ai_1 _16497_ (.B1(_07989_),
    .Y(_07990_),
    .A1(_07727_),
    .A2(_02442_));
 sg13g2_a21oi_1 _16498_ (.A1(_07988_),
    .A2(_07990_),
    .Y(_07991_),
    .B1(net294));
 sg13g2_a21oi_1 _16499_ (.A1(_02456_),
    .A2(_01905_),
    .Y(_07992_),
    .B1(_02583_));
 sg13g2_o21ai_1 _16500_ (.B1(_07992_),
    .Y(_07993_),
    .A1(net405),
    .A2(_01905_));
 sg13g2_o21ai_1 _16501_ (.B1(_07993_),
    .Y(_07994_),
    .A1(_07981_),
    .A2(_07991_));
 sg13g2_nand2_1 _16502_ (.Y(_07995_),
    .A(_07994_),
    .B(_02585_));
 sg13g2_nand3_1 _16503_ (.B(_02526_),
    .C(_07995_),
    .A(_07974_),
    .Y(_07996_));
 sg13g2_a21oi_1 _16504_ (.A1(_07581_),
    .A2(_07801_),
    .Y(_01321_),
    .B1(_02197_));
 sg13g2_nand2_1 _16505_ (.Y(_01322_),
    .A(_07996_),
    .B(_01321_));
 sg13g2_nand2_1 _16506_ (.Y(_01323_),
    .A(net250),
    .B(_01866_));
 sg13g2_nand2_1 _16507_ (.Y(\addr_pins_out[3] ),
    .A(_01322_),
    .B(_01323_));
 sg13g2_nand2_1 _16508_ (.Y(_01324_),
    .A(_03309_),
    .B(_07500_));
 sg13g2_nor2_1 _16509_ (.A(_05089_),
    .B(_05732_),
    .Y(_01325_));
 sg13g2_a221oi_1 _16510_ (.B2(_05525_),
    .C1(_01325_),
    .B1(\synth.voice.scan_outs[2][0] ),
    .A1(_04786_),
    .Y(_01326_),
    .A2(_03660_));
 sg13g2_nor2_1 _16511_ (.A(_00058_),
    .B(_04718_),
    .Y(_01327_));
 sg13g2_nor2_1 _16512_ (.A(_01766_),
    .B(_04813_),
    .Y(_01328_));
 sg13g2_nor2_1 _16513_ (.A(_00059_),
    .B(_04352_),
    .Y(_01329_));
 sg13g2_inv_1 _16514_ (.Y(_01330_),
    .A(\synth.voice.params[24] ));
 sg13g2_nor4_1 _16515_ (.A(_01330_),
    .B(_03587_),
    .C(_04350_),
    .D(_04029_),
    .Y(_01331_));
 sg13g2_nor4_1 _16516_ (.A(_01327_),
    .B(_01328_),
    .C(_01329_),
    .D(_01331_),
    .Y(_01332_));
 sg13g2_a22oi_1 _16517_ (.Y(_01333_),
    .B1(_05047_),
    .B2(_05821_),
    .A2(\synth.voice.float_period[0][8] ),
    .A1(_05908_));
 sg13g2_a22oi_1 _16518_ (.Y(_01334_),
    .B1(_03451_),
    .B2(_04030_),
    .A2(\synth.voice.mods[1][2] ),
    .A1(_07510_));
 sg13g2_nand4_1 _16519_ (.B(_01332_),
    .C(_01333_),
    .A(_01326_),
    .Y(_01335_),
    .D(_01334_));
 sg13g2_nand2_1 _16520_ (.Y(_01336_),
    .A(_07506_),
    .B(_03668_));
 sg13g2_o21ai_1 _16521_ (.B1(_01336_),
    .Y(_01337_),
    .A1(_07506_),
    .A2(_01335_));
 sg13g2_o21ai_1 _16522_ (.B1(_03404_),
    .Y(_01338_),
    .A1(_00056_),
    .A2(_03309_));
 sg13g2_nand2_1 _16523_ (.Y(_01339_),
    .A(\synth.controller.curr_voice[1] ),
    .B(_00182_));
 sg13g2_a21oi_1 _16524_ (.A1(\synth.controller.sweep_addr_index[2] ),
    .A2(_03400_),
    .Y(_01340_),
    .B1(_03401_));
 sg13g2_nand2_1 _16525_ (.Y(_01341_),
    .A(_07501_),
    .B(\synth.controller.sweep_addr_index[0] ));
 sg13g2_nand2_1 _16526_ (.Y(_01342_),
    .A(_07103_),
    .B(_03403_));
 sg13g2_a221oi_1 _16527_ (.B2(_01341_),
    .C1(_01342_),
    .B1(_01340_),
    .A1(_03401_),
    .Y(_01343_),
    .A2(_01339_));
 sg13g2_nor2_1 _16528_ (.A(_01338_),
    .B(_01343_),
    .Y(_01344_));
 sg13g2_o21ai_1 _16529_ (.B1(_01344_),
    .Y(_01345_),
    .A1(_01324_),
    .A2(_01337_));
 sg13g2_nand2_1 _16530_ (.Y(_01346_),
    .A(_03304_),
    .B(_00055_));
 sg13g2_nand3_1 _16531_ (.B(_07093_),
    .C(_01346_),
    .A(_01345_),
    .Y(_01347_));
 sg13g2_nand2_1 _16532_ (.Y(\synth.controller.sbio_tx.start_present ),
    .A(_01347_),
    .B(_03406_));
 sg13g2_nor2b_1 _16533_ (.A(_01747_),
    .B_N(_01759_),
    .Y(_01348_));
 sg13g2_nand2b_1 _16534_ (.Y(_01349_),
    .B(_04391_),
    .A_N(_01783_));
 sg13g2_nand2_1 _16535_ (.Y(_01350_),
    .A(_01783_),
    .B(\synth.voice.genblk4[8].next_state_scan[5] ));
 sg13g2_nand3_1 _16536_ (.B(_01758_),
    .C(_01350_),
    .A(_01349_),
    .Y(_01351_));
 sg13g2_xnor2_1 _16537_ (.Y(_01352_),
    .A(_01348_),
    .B(_01351_));
 sg13g2_nor2_1 _16538_ (.A(\synth.voice.flip_sign_fir ),
    .B(net201),
    .Y(_01353_));
 sg13g2_a21oi_1 _16539_ (.A1(_01352_),
    .A2(net201),
    .Y(\synth.voice.flip_sign ),
    .B1(_01353_));
 sg13g2_nor3_1 _16540_ (.A(_01793_),
    .B(_06741_),
    .C(_01794_),
    .Y(_01354_));
 sg13g2_inv_1 _16541_ (.Y(_01355_),
    .A(_01354_));
 sg13g2_nor3_2 _16542_ (.A(_01715_),
    .B(_06741_),
    .C(_01794_),
    .Y(_01356_));
 sg13g2_nor2_1 _16543_ (.A(_01356_),
    .B(_06713_),
    .Y(_01357_));
 sg13g2_a21oi_1 _16544_ (.A1(_06766_),
    .A2(_01355_),
    .Y(_01358_),
    .B1(_01357_));
 sg13g2_nor2_1 _16545_ (.A(_01719_),
    .B(_01358_),
    .Y(_01359_));
 sg13g2_nand2_1 _16546_ (.Y(_01360_),
    .A(_01717_),
    .B(_06744_));
 sg13g2_a21oi_1 _16547_ (.A1(_01355_),
    .A2(_01360_),
    .Y(_01361_),
    .B1(_06792_));
 sg13g2_inv_2 _16548_ (.Y(_01362_),
    .A(_01356_));
 sg13g2_nor2_1 _16549_ (.A(_01362_),
    .B(_06711_),
    .Y(_01363_));
 sg13g2_nor2_1 _16550_ (.A(_06752_),
    .B(_06750_),
    .Y(_01364_));
 sg13g2_inv_1 _16551_ (.Y(_01365_),
    .A(_06780_));
 sg13g2_inv_1 _16552_ (.Y(_01366_),
    .A(_06777_));
 sg13g2_nor3_1 _16553_ (.A(_06765_),
    .B(_01365_),
    .C(_01366_),
    .Y(_01367_));
 sg13g2_a21oi_1 _16554_ (.A1(_01364_),
    .A2(_01367_),
    .Y(_01368_),
    .B1(_01355_));
 sg13g2_nor4_1 _16555_ (.A(_01359_),
    .B(_01361_),
    .C(_01363_),
    .D(_01368_),
    .Y(_01369_));
 sg13g2_inv_1 _16556_ (.Y(_01370_),
    .A(_06722_));
 sg13g2_o21ai_1 _16557_ (.B1(_01796_),
    .Y(_01371_),
    .A1(_01370_),
    .A2(_06738_));
 sg13g2_nand2_1 _16558_ (.Y(_01372_),
    .A(_06781_),
    .B(_06782_));
 sg13g2_nor2_1 _16559_ (.A(_06689_),
    .B(_06678_),
    .Y(_01373_));
 sg13g2_inv_1 _16560_ (.Y(_01374_),
    .A(_06709_));
 sg13g2_a21oi_1 _16561_ (.A1(_01373_),
    .A2(_01374_),
    .Y(_01375_),
    .B1(net219));
 sg13g2_nor2_1 _16562_ (.A(_06744_),
    .B(_06741_),
    .Y(_01376_));
 sg13g2_buf_2 _16563_ (.A(_01376_),
    .X(_01377_));
 sg13g2_o21ai_1 _16564_ (.B1(_01377_),
    .Y(_01378_),
    .A1(_01372_),
    .A2(_01375_));
 sg13g2_inv_1 _16565_ (.Y(_01379_),
    .A(_06708_));
 sg13g2_nand3b_1 _16566_ (.B(_01379_),
    .C(_06692_),
    .Y(_01380_),
    .A_N(_06717_));
 sg13g2_inv_1 _16567_ (.Y(_01381_),
    .A(_01364_));
 sg13g2_nand2_1 _16568_ (.Y(_01382_),
    .A(net265),
    .B(_01362_));
 sg13g2_buf_2 _16569_ (.A(_01382_),
    .X(_01383_));
 sg13g2_o21ai_1 _16570_ (.B1(_01383_),
    .Y(_01384_),
    .A1(_01380_),
    .A2(_01381_));
 sg13g2_nand4_1 _16571_ (.B(_01371_),
    .C(_01378_),
    .A(_01369_),
    .Y(\synth.voice.fir_table.sign ),
    .D(_01384_));
 sg13g2_inv_1 _16572_ (.Y(_01385_),
    .A(_01377_));
 sg13g2_o21ai_1 _16573_ (.B1(_01385_),
    .Y(_01386_),
    .A1(_01365_),
    .A2(_06748_));
 sg13g2_nand2_1 _16574_ (.Y(_01387_),
    .A(_06724_),
    .B(net265));
 sg13g2_nand2_1 _16575_ (.Y(_01388_),
    .A(_06732_),
    .B(_01796_));
 sg13g2_nand3_1 _16576_ (.B(_01387_),
    .C(_01388_),
    .A(_01386_),
    .Y(_01389_));
 sg13g2_nor2_1 _16577_ (.A(_01796_),
    .B(_01354_),
    .Y(_01390_));
 sg13g2_nor2_1 _16578_ (.A(_01390_),
    .B(_06762_),
    .Y(_01391_));
 sg13g2_nor2_1 _16579_ (.A(_01377_),
    .B(_01796_),
    .Y(_01392_));
 sg13g2_inv_2 _16580_ (.Y(_01393_),
    .A(_01383_));
 sg13g2_nor2_1 _16581_ (.A(_01392_),
    .B(_01393_),
    .Y(_01394_));
 sg13g2_nor2b_1 _16582_ (.A(_06777_),
    .B_N(_01394_),
    .Y(_01395_));
 sg13g2_nor2_1 _16583_ (.A(_01354_),
    .B(_01392_),
    .Y(_01396_));
 sg13g2_nor2_1 _16584_ (.A(_01396_),
    .B(_06768_),
    .Y(_01397_));
 sg13g2_nor2_1 _16585_ (.A(_01794_),
    .B(_01717_),
    .Y(_01398_));
 sg13g2_inv_1 _16586_ (.Y(_01399_),
    .A(_01360_));
 sg13g2_nor2_1 _16587_ (.A(_01398_),
    .B(_01399_),
    .Y(_01400_));
 sg13g2_nor2_1 _16588_ (.A(_01400_),
    .B(_06786_),
    .Y(_01401_));
 sg13g2_nor4_1 _16589_ (.A(_01391_),
    .B(_01395_),
    .C(_01397_),
    .D(_01401_),
    .Y(_01402_));
 sg13g2_inv_1 _16590_ (.Y(_01403_),
    .A(_01392_));
 sg13g2_nor2_1 _16591_ (.A(_01403_),
    .B(_06782_),
    .Y(_01404_));
 sg13g2_nor2_1 _16592_ (.A(_01796_),
    .B(_06692_),
    .Y(_01405_));
 sg13g2_nor3_1 _16593_ (.A(_01716_),
    .B(_06744_),
    .C(_01793_),
    .Y(_01406_));
 sg13g2_inv_1 _16594_ (.Y(_01407_),
    .A(_01406_));
 sg13g2_nor2_1 _16595_ (.A(_01407_),
    .B(_06761_),
    .Y(_01408_));
 sg13g2_a21oi_1 _16596_ (.A1(_01360_),
    .A2(_01390_),
    .Y(_01409_),
    .B1(_06787_));
 sg13g2_nor4_1 _16597_ (.A(_01404_),
    .B(_01405_),
    .C(_01408_),
    .D(_01409_),
    .Y(_01410_));
 sg13g2_nand2_1 _16598_ (.Y(_01411_),
    .A(_01402_),
    .B(_01410_));
 sg13g2_nor2_1 _16599_ (.A(_01385_),
    .B(_06775_),
    .Y(_01412_));
 sg13g2_nor2_1 _16600_ (.A(net265),
    .B(_06726_),
    .Y(_01413_));
 sg13g2_inv_1 _16601_ (.Y(_01414_),
    .A(_06751_));
 sg13g2_nor2_1 _16602_ (.A(_01396_),
    .B(_01414_),
    .Y(_01415_));
 sg13g2_nor4_1 _16603_ (.A(_01412_),
    .B(_01357_),
    .C(_01413_),
    .D(_01415_),
    .Y(_01416_));
 sg13g2_nor2_1 _16604_ (.A(_01393_),
    .B(_06702_),
    .Y(_01417_));
 sg13g2_o21ai_1 _16605_ (.B1(_01417_),
    .Y(_01418_),
    .A1(_06691_),
    .A2(_06736_));
 sg13g2_nor2_1 _16606_ (.A(_06728_),
    .B(_06755_),
    .Y(_01419_));
 sg13g2_nor2_1 _16607_ (.A(_01419_),
    .B(_06730_),
    .Y(_01420_));
 sg13g2_nand4_1 _16608_ (.B(_06711_),
    .C(_01418_),
    .A(_01416_),
    .Y(_01421_),
    .D(_01420_));
 sg13g2_nor3_1 _16609_ (.A(_01389_),
    .B(_01411_),
    .C(_01421_),
    .Y(_01422_));
 sg13g2_nand2_1 _16610_ (.Y(_01423_),
    .A(_06709_),
    .B(_01383_));
 sg13g2_o21ai_1 _16611_ (.B1(_01423_),
    .Y(_01424_),
    .A1(_06764_),
    .A2(_01362_));
 sg13g2_nand2_1 _16612_ (.Y(_01425_),
    .A(_06770_),
    .B(_06781_));
 sg13g2_inv_1 _16613_ (.Y(_01426_),
    .A(_01425_));
 sg13g2_nand2_1 _16614_ (.Y(_01427_),
    .A(_01426_),
    .B(_06707_));
 sg13g2_inv_1 _16615_ (.Y(_01428_),
    .A(_06747_));
 sg13g2_a22oi_1 _16616_ (.Y(_01429_),
    .B1(_01428_),
    .B2(_06758_),
    .A2(_01403_),
    .A1(_01362_));
 sg13g2_a221oi_1 _16617_ (.B2(_01427_),
    .C1(_01429_),
    .B1(net265),
    .A1(net205),
    .Y(_01430_),
    .A2(_01424_));
 sg13g2_nand3_1 _16618_ (.B(_06703_),
    .C(_01403_),
    .A(_06683_),
    .Y(_01431_));
 sg13g2_a21oi_1 _16619_ (.A1(_01431_),
    .A2(_06792_),
    .Y(_01432_),
    .B1(_01362_));
 sg13g2_a21oi_1 _16620_ (.A1(_01393_),
    .A2(_01403_),
    .Y(_01433_),
    .B1(_06767_));
 sg13g2_inv_1 _16621_ (.Y(_01434_),
    .A(_06690_));
 sg13g2_nand2_1 _16622_ (.Y(_01435_),
    .A(_06679_),
    .B(_06700_));
 sg13g2_nor3_1 _16623_ (.A(_01434_),
    .B(_06752_),
    .C(_01435_),
    .Y(_01436_));
 sg13g2_nor2_1 _16624_ (.A(_01407_),
    .B(_01436_),
    .Y(_01437_));
 sg13g2_inv_1 _16625_ (.Y(_01438_),
    .A(_06773_));
 sg13g2_o21ai_1 _16626_ (.B1(_01438_),
    .Y(_01439_),
    .A1(_01385_),
    .A2(_01383_));
 sg13g2_a21oi_1 _16627_ (.A1(_01716_),
    .A2(_00045_),
    .Y(_01440_),
    .B1(_01399_));
 sg13g2_nand2_1 _16628_ (.Y(_01441_),
    .A(_06790_),
    .B(_01440_));
 sg13g2_nand3_1 _16629_ (.B(net205),
    .C(_01393_),
    .A(_06665_),
    .Y(_01442_));
 sg13g2_nand2_1 _16630_ (.Y(_01443_),
    .A(_01390_),
    .B(_01377_));
 sg13g2_nand2_1 _16631_ (.Y(_01444_),
    .A(_06753_),
    .B(_01443_));
 sg13g2_nand4_1 _16632_ (.B(_01441_),
    .C(_01442_),
    .A(_01439_),
    .Y(_01445_),
    .D(_01444_));
 sg13g2_nor4_1 _16633_ (.A(_01432_),
    .B(_01433_),
    .C(_01437_),
    .D(_01445_),
    .Y(_01446_));
 sg13g2_nand3_1 _16634_ (.B(_01430_),
    .C(_01446_),
    .A(_01422_),
    .Y(\synth.voice.fir_table.exp[0] ));
 sg13g2_nor2b_1 _16635_ (.A(_06779_),
    .B_N(_06758_),
    .Y(_01447_));
 sg13g2_nand2_1 _16636_ (.Y(_01448_),
    .A(_01447_),
    .B(_06700_));
 sg13g2_nor2_1 _16637_ (.A(_06788_),
    .B(_06750_),
    .Y(_01449_));
 sg13g2_inv_1 _16638_ (.Y(_01450_),
    .A(_06793_));
 sg13g2_nand4_1 _16639_ (.B(_01450_),
    .C(_06707_),
    .A(_01449_),
    .Y(_01451_),
    .D(_06704_));
 sg13g2_nor3_1 _16640_ (.A(_06717_),
    .B(_06716_),
    .C(_06724_),
    .Y(_01452_));
 sg13g2_nor2_1 _16641_ (.A(_06693_),
    .B(_06779_),
    .Y(_01453_));
 sg13g2_nand4_1 _16642_ (.B(_06754_),
    .C(_06758_),
    .A(_01452_),
    .Y(_01454_),
    .D(_01453_));
 sg13g2_nor4_1 _16643_ (.A(_06714_),
    .B(_06783_),
    .C(_01451_),
    .D(_01454_),
    .Y(_01455_));
 sg13g2_nand4_1 _16644_ (.B(_06672_),
    .C(_06700_),
    .A(_06679_),
    .Y(_01456_),
    .D(_06684_));
 sg13g2_nand4_1 _16645_ (.B(_06775_),
    .C(_06773_),
    .A(_01420_),
    .Y(_01457_),
    .D(_06726_));
 sg13g2_nor4_1 _16646_ (.A(_06732_),
    .B(_06734_),
    .C(_01456_),
    .D(_01457_),
    .Y(_01458_));
 sg13g2_and3_1 _16647_ (.X(_01459_),
    .A(_01455_),
    .B(_06772_),
    .C(_01458_));
 sg13g2_buf_1 _16648_ (.A(_01459_),
    .X(_01460_));
 sg13g2_o21ai_1 _16649_ (.B1(net265),
    .Y(_01461_),
    .A1(_01448_),
    .A2(_01460_));
 sg13g2_nand3b_1 _16650_ (.B(_06692_),
    .C(_06704_),
    .Y(_01462_),
    .A_N(_06717_));
 sg13g2_nand2_1 _16651_ (.Y(_01463_),
    .A(_01462_),
    .B(_01362_));
 sg13g2_o21ai_1 _16652_ (.B1(_06787_),
    .Y(_01464_),
    .A1(_01356_),
    .A2(_06786_));
 sg13g2_nand3_1 _16653_ (.B(_06684_),
    .C(_06768_),
    .A(_01379_),
    .Y(_01465_));
 sg13g2_a22oi_1 _16654_ (.Y(_01466_),
    .B1(_01406_),
    .B2(_01465_),
    .A2(_01360_),
    .A1(_01464_));
 sg13g2_nor3_1 _16655_ (.A(_06765_),
    .B(_06766_),
    .C(_01365_),
    .Y(_01467_));
 sg13g2_nand2_1 _16656_ (.Y(_01468_),
    .A(_06770_),
    .B(_06775_));
 sg13g2_nand2_1 _16657_ (.Y(_01469_),
    .A(_01428_),
    .B(_06782_));
 sg13g2_nor2_1 _16658_ (.A(_06744_),
    .B(_01355_),
    .Y(_01470_));
 sg13g2_inv_1 _16659_ (.Y(_01471_),
    .A(_01388_));
 sg13g2_a221oi_1 _16660_ (.B2(_01470_),
    .C1(_01471_),
    .B1(_01469_),
    .A1(_01468_),
    .Y(_01472_),
    .A2(_01394_));
 sg13g2_o21ai_1 _16661_ (.B1(_01472_),
    .Y(_01473_),
    .A1(_01385_),
    .A2(_01467_));
 sg13g2_inv_1 _16662_ (.Y(_01474_),
    .A(_01390_));
 sg13g2_nor4_1 _16663_ (.A(_06744_),
    .B(_06745_),
    .C(_01362_),
    .D(_01373_),
    .Y(_01475_));
 sg13g2_a221oi_1 _16664_ (.B2(_01474_),
    .C1(_01475_),
    .B1(_01438_),
    .A1(_06751_),
    .Y(_01476_),
    .A2(_01385_));
 sg13g2_nor3_1 _16665_ (.A(net265),
    .B(_06728_),
    .C(_06729_),
    .Y(_01477_));
 sg13g2_nor2_1 _16666_ (.A(_01398_),
    .B(_06792_),
    .Y(_01478_));
 sg13g2_a21oi_1 _16667_ (.A1(_01393_),
    .A2(_01403_),
    .Y(_01479_),
    .B1(_06762_));
 sg13g2_a21oi_1 _16668_ (.A1(_01793_),
    .A2(_01377_),
    .Y(_01480_),
    .B1(_01399_));
 sg13g2_nor3_1 _16669_ (.A(_01400_),
    .B(_01480_),
    .C(_06791_),
    .Y(_01481_));
 sg13g2_nor4_1 _16670_ (.A(_01477_),
    .B(_01478_),
    .C(_01479_),
    .D(_01481_),
    .Y(_01482_));
 sg13g2_nor2_1 _16671_ (.A(_01393_),
    .B(_06672_),
    .Y(_01483_));
 sg13g2_nor2_1 _16672_ (.A(_06734_),
    .B(_06716_),
    .Y(_01484_));
 sg13g2_nand3_1 _16673_ (.B(_06679_),
    .C(_06761_),
    .A(_01484_),
    .Y(_01485_));
 sg13g2_nor3_1 _16674_ (.A(_06724_),
    .B(_01483_),
    .C(_01485_),
    .Y(_01486_));
 sg13g2_nor3_1 _16675_ (.A(net219),
    .B(_01403_),
    .C(_06746_),
    .Y(_01487_));
 sg13g2_inv_1 _16676_ (.Y(_01488_),
    .A(_01396_));
 sg13g2_o21ai_1 _16677_ (.B1(_01488_),
    .Y(_01489_),
    .A1(_06752_),
    .A2(_01487_));
 sg13g2_nand4_1 _16678_ (.B(_01482_),
    .C(_01486_),
    .A(_01476_),
    .Y(_01490_),
    .D(_01489_));
 sg13g2_nor2_1 _16679_ (.A(_01473_),
    .B(_01490_),
    .Y(_01491_));
 sg13g2_nand4_1 _16680_ (.B(_01463_),
    .C(_01466_),
    .A(_01461_),
    .Y(\synth.voice.fir_table.exp[1] ),
    .D(_01491_));
 sg13g2_nand2_1 _16681_ (.Y(_01492_),
    .A(_06768_),
    .B(_06723_));
 sg13g2_nor2_1 _16682_ (.A(_01492_),
    .B(_01469_),
    .Y(_01493_));
 sg13g2_nand4_1 _16683_ (.B(_06754_),
    .C(_06718_),
    .A(_01493_),
    .Y(_01494_),
    .D(_06715_));
 sg13g2_nand3_1 _16684_ (.B(_06722_),
    .C(_06704_),
    .A(_06737_),
    .Y(_01495_));
 sg13g2_a22oi_1 _16685_ (.Y(_01496_),
    .B1(_01377_),
    .B2(_01438_),
    .A2(_01796_),
    .A1(_06734_));
 sg13g2_nand3_1 _16686_ (.B(_06697_),
    .C(_01383_),
    .A(_06699_),
    .Y(_01497_));
 sg13g2_nand3_1 _16687_ (.B(net205),
    .C(_01470_),
    .A(_06774_),
    .Y(_01498_));
 sg13g2_nand3_1 _16688_ (.B(_01497_),
    .C(_01498_),
    .A(_01496_),
    .Y(_01499_));
 sg13g2_nor4_1 _16689_ (.A(_01413_),
    .B(_01405_),
    .C(_01495_),
    .D(_01499_),
    .Y(_01500_));
 sg13g2_o21ai_1 _16690_ (.B1(_01356_),
    .Y(_01501_),
    .A1(_01434_),
    .A2(_06685_));
 sg13g2_nor2_1 _16691_ (.A(_01383_),
    .B(_01450_),
    .Y(_01502_));
 sg13g2_a221oi_1 _16692_ (.B2(_01443_),
    .C1(_01502_),
    .B1(_06763_),
    .A1(_06788_),
    .Y(_01503_),
    .A2(_01385_));
 sg13g2_nand3_1 _16693_ (.B(_01501_),
    .C(_01503_),
    .A(_01500_),
    .Y(_01504_));
 sg13g2_a21oi_1 _16694_ (.A1(net265),
    .A2(_01494_),
    .Y(_01505_),
    .B1(_01504_));
 sg13g2_nor2_1 _16695_ (.A(_06748_),
    .B(_01425_),
    .Y(_01506_));
 sg13g2_nand3_1 _16696_ (.B(_01467_),
    .C(_01506_),
    .A(_01447_),
    .Y(_01507_));
 sg13g2_a21oi_1 _16697_ (.A1(_01488_),
    .A2(_01507_),
    .Y(_01508_),
    .B1(_01460_));
 sg13g2_a22oi_1 _16698_ (.Y(\synth.voice.fir_table.exp[2] ),
    .B1(_01505_),
    .B2(_01508_),
    .A2(_01460_),
    .A1(_01393_));
 sg13g2_nor3_1 _16699_ (.A(_06783_),
    .B(_01366_),
    .C(_06771_),
    .Y(_01509_));
 sg13g2_a21oi_1 _16700_ (.A1(_01509_),
    .A2(_06760_),
    .Y(_01510_),
    .B1(_01392_));
 sg13g2_nor2_1 _16701_ (.A(_01510_),
    .B(_01460_),
    .Y(_01511_));
 sg13g2_o21ai_1 _16702_ (.B1(_06692_),
    .Y(_01512_),
    .A1(net265),
    .A2(_06737_));
 sg13g2_o21ai_1 _16703_ (.B1(_01383_),
    .Y(_01513_),
    .A1(_01512_),
    .A2(_06719_));
 sg13g2_nor2_1 _16704_ (.A(_01362_),
    .B(_06704_),
    .Y(_01514_));
 sg13g2_nand2_1 _16705_ (.Y(_01515_),
    .A(_01431_),
    .B(_06690_));
 sg13g2_inv_1 _16706_ (.Y(_01516_),
    .A(_01400_));
 sg13g2_a22oi_1 _16707_ (.Y(_01517_),
    .B1(_01516_),
    .B2(_06793_),
    .A2(_01377_),
    .A1(_06763_));
 sg13g2_inv_1 _16708_ (.Y(_01518_),
    .A(_01440_));
 sg13g2_a22oi_1 _16709_ (.Y(_01519_),
    .B1(_01518_),
    .B2(_06788_),
    .A2(_01796_),
    .A1(_06724_));
 sg13g2_nand2_1 _16710_ (.Y(_01520_),
    .A(_01517_),
    .B(_01519_));
 sg13g2_nor3_1 _16711_ (.A(_01514_),
    .B(_01515_),
    .C(_01520_),
    .Y(_01521_));
 sg13g2_nand4_1 _16712_ (.B(_01458_),
    .C(_01513_),
    .A(_01511_),
    .Y(\synth.voice.fir_table.exp[3] ),
    .D(_01521_));
 sg13g2_inv_1 _16713_ (.Y(_01522_),
    .A(_00170_));
 sg13g2_nand2_1 _16714_ (.Y(_01523_),
    .A(_01752_),
    .B(_01766_));
 sg13g2_nand3_1 _16715_ (.B(_01765_),
    .C(_01751_),
    .A(_01749_),
    .Y(_01524_));
 sg13g2_nand2_1 _16716_ (.Y(_01525_),
    .A(_01749_),
    .B(_01767_));
 sg13g2_nand3_1 _16717_ (.B(_01524_),
    .C(_01525_),
    .A(_01523_),
    .Y(_01526_));
 sg13g2_nand2_1 _16718_ (.Y(_01527_),
    .A(_01526_),
    .B(_04699_));
 sg13g2_buf_8 _16719_ (.A(_01527_),
    .X(_01528_));
 sg13g2_inv_4 _16720_ (.A(_01528_),
    .Y(_01529_));
 sg13g2_nand3b_1 _16721_ (.B(_01766_),
    .C(_01765_),
    .Y(_01530_),
    .A_N(_00150_));
 sg13g2_nand2_1 _16722_ (.Y(_01531_),
    .A(_01758_),
    .B(_01530_));
 sg13g2_buf_2 _16723_ (.A(_01531_),
    .X(_01532_));
 sg13g2_buf_8 _16724_ (.A(_01532_),
    .X(_01533_));
 sg13g2_inv_1 _16725_ (.Y(_01534_),
    .A(net164));
 sg13g2_nor2_1 _16726_ (.A(_01534_),
    .B(_01529_),
    .Y(_01535_));
 sg13g2_a22oi_1 _16727_ (.Y(_01536_),
    .B1(_03757_),
    .B2(_01535_),
    .A2(_01534_),
    .A1(\synth.voice.genblk4[7].next_state_scan[12] ));
 sg13g2_nand2_1 _16728_ (.Y(_01537_),
    .A(_01536_),
    .B(_01739_));
 sg13g2_a21oi_1 _16729_ (.A1(_01522_),
    .A2(_01529_),
    .Y(_01538_),
    .B1(_01537_));
 sg13g2_a21oi_1 _16730_ (.A1(_00169_),
    .A2(net202),
    .Y(_01539_),
    .B1(_01538_));
 sg13g2_nand2_1 _16731_ (.Y(_01540_),
    .A(_01529_),
    .B(_00166_));
 sg13g2_nand2_1 _16732_ (.Y(_01541_),
    .A(_01532_),
    .B(_03772_));
 sg13g2_o21ai_1 _16733_ (.B1(_01541_),
    .Y(_01542_),
    .A1(_03773_),
    .A2(_01532_));
 sg13g2_nand2_1 _16734_ (.Y(_01543_),
    .A(_01528_),
    .B(_01542_));
 sg13g2_nand2_1 _16735_ (.Y(_01544_),
    .A(_01540_),
    .B(_01543_));
 sg13g2_nor2_1 _16736_ (.A(_04956_),
    .B(_01544_),
    .Y(_01545_));
 sg13g2_buf_8 _16737_ (.A(_01528_),
    .X(_01546_));
 sg13g2_nor2b_1 _16738_ (.A(net129),
    .B_N(_00167_),
    .Y(_01547_));
 sg13g2_nor2b_1 _16739_ (.A(_01532_),
    .B_N(\synth.voice.genblk4[7].next_state_scan[8] ),
    .Y(_01548_));
 sg13g2_a21oi_1 _16740_ (.A1(\synth.voice.mods[1][2] ),
    .A2(net164),
    .Y(_01549_),
    .B1(_01548_));
 sg13g2_nor2b_1 _16741_ (.A(_01529_),
    .B_N(_01549_),
    .Y(_01550_));
 sg13g2_nor3_1 _16742_ (.A(_04968_),
    .B(_01547_),
    .C(_01550_),
    .Y(_01551_));
 sg13g2_nand2b_1 _16743_ (.Y(_01552_),
    .B(_01544_),
    .A_N(_00140_));
 sg13g2_nand3_1 _16744_ (.B(_01543_),
    .C(_00140_),
    .A(_01540_),
    .Y(_01553_));
 sg13g2_nand3_1 _16745_ (.B(_01552_),
    .C(_01553_),
    .A(_01551_),
    .Y(_01554_));
 sg13g2_nand2b_1 _16746_ (.Y(_01555_),
    .B(_01554_),
    .A_N(_01545_));
 sg13g2_nor2_1 _16747_ (.A(\synth.voice.genblk4[7].next_state_scan[10] ),
    .B(net164),
    .Y(_01556_));
 sg13g2_a21o_1 _16748_ (.A2(net164),
    .A1(_04257_),
    .B1(_01556_),
    .X(_01557_));
 sg13g2_nor2b_1 _16749_ (.A(net129),
    .B_N(_00165_),
    .Y(_01558_));
 sg13g2_a21oi_2 _16750_ (.B1(_01558_),
    .Y(_01559_),
    .A2(net129),
    .A1(_01557_));
 sg13g2_xnor2_1 _16751_ (.Y(_01560_),
    .A(_04960_),
    .B(_01559_));
 sg13g2_nand2b_1 _16752_ (.Y(_01561_),
    .B(_01529_),
    .A_N(_00164_));
 sg13g2_inv_1 _16753_ (.Y(_01562_),
    .A(\synth.voice.genblk4[7].next_state_scan[1] ));
 sg13g2_nor2_1 _16754_ (.A(\synth.voice.genblk4[7].next_state_scan[11] ),
    .B(_01532_),
    .Y(_01563_));
 sg13g2_a21oi_1 _16755_ (.A1(_01562_),
    .A2(_01532_),
    .Y(_01564_),
    .B1(_01563_));
 sg13g2_nand2_1 _16756_ (.Y(_01565_),
    .A(_01528_),
    .B(_01564_));
 sg13g2_nand2_1 _16757_ (.Y(_01566_),
    .A(_01561_),
    .B(_01565_));
 sg13g2_nor2_1 _16758_ (.A(_04934_),
    .B(_01566_),
    .Y(_01567_));
 sg13g2_nand2_1 _16759_ (.Y(_01568_),
    .A(_01566_),
    .B(_04934_));
 sg13g2_nand2b_1 _16760_ (.Y(_01569_),
    .B(_01568_),
    .A_N(_01567_));
 sg13g2_nor2_1 _16761_ (.A(_01560_),
    .B(_01569_),
    .Y(_01570_));
 sg13g2_nand2_1 _16762_ (.Y(_01571_),
    .A(_01559_),
    .B(_04941_));
 sg13g2_o21ai_1 _16763_ (.B1(_01568_),
    .Y(_01572_),
    .A1(_01567_),
    .A2(_01571_));
 sg13g2_a21oi_1 _16764_ (.A1(_01555_),
    .A2(_01570_),
    .Y(_01573_),
    .B1(_01572_));
 sg13g2_nand2_1 _16765_ (.Y(_01574_),
    .A(_01552_),
    .B(_01553_));
 sg13g2_nor2_1 _16766_ (.A(_01547_),
    .B(_01550_),
    .Y(_01575_));
 sg13g2_nor2_1 _16767_ (.A(_00141_),
    .B(_01575_),
    .Y(_01576_));
 sg13g2_nor2_1 _16768_ (.A(_01551_),
    .B(_01576_),
    .Y(_01577_));
 sg13g2_nand2b_1 _16769_ (.Y(_01578_),
    .B(_01577_),
    .A_N(_01574_));
 sg13g2_xor2_1 _16770_ (.B(_01559_),
    .A(_04960_),
    .X(_01579_));
 sg13g2_nor2b_1 _16771_ (.A(_01567_),
    .B_N(_01568_),
    .Y(_01580_));
 sg13g2_nand2_1 _16772_ (.Y(_01581_),
    .A(_01579_),
    .B(_01580_));
 sg13g2_nor2_1 _16773_ (.A(_01578_),
    .B(_01581_),
    .Y(_01582_));
 sg13g2_nand2_1 _16774_ (.Y(_01583_),
    .A(net164),
    .B(_03816_));
 sg13g2_o21ai_1 _16775_ (.B1(_01583_),
    .Y(_01584_),
    .A1(_03817_),
    .A2(net164));
 sg13g2_nor2_1 _16776_ (.A(_03818_),
    .B(net129),
    .Y(_01585_));
 sg13g2_a21oi_1 _16777_ (.A1(net129),
    .A2(_01584_),
    .Y(_01586_),
    .B1(_01585_));
 sg13g2_nor2_1 _16778_ (.A(_00143_),
    .B(_01586_),
    .Y(_01587_));
 sg13g2_nor2b_1 _16779_ (.A(_01533_),
    .B_N(\synth.voice.genblk4[7].next_state_scan[7] ),
    .Y(_01588_));
 sg13g2_a21oi_1 _16780_ (.A1(\synth.voice.genblk4[6].next_state_scan[13] ),
    .A2(_01533_),
    .Y(_01589_),
    .B1(_01588_));
 sg13g2_inv_1 _16781_ (.Y(_01590_),
    .A(_01589_));
 sg13g2_nor2_1 _16782_ (.A(_00168_),
    .B(net129),
    .Y(_01591_));
 sg13g2_a21oi_1 _16783_ (.A1(net129),
    .A2(_01590_),
    .Y(_01592_),
    .B1(_01591_));
 sg13g2_xnor2_1 _16784_ (.Y(_01593_),
    .A(_04979_),
    .B(_01592_));
 sg13g2_or2_1 _16785_ (.X(_01594_),
    .B(_01592_),
    .A(\synth.voice.genblk4[1].next_state_scan[12] ));
 sg13g2_o21ai_1 _16786_ (.B1(_01594_),
    .Y(_01595_),
    .A1(_01587_),
    .A2(_01593_));
 sg13g2_nand2_1 _16787_ (.Y(_01596_),
    .A(_01582_),
    .B(_01595_));
 sg13g2_nand2_1 _16788_ (.Y(_01597_),
    .A(_01573_),
    .B(_01596_));
 sg13g2_xor2_1 _16789_ (.B(_01586_),
    .A(\synth.voice.genblk4[1].next_state_scan[13] ),
    .X(_01598_));
 sg13g2_nor3_1 _16790_ (.A(_01593_),
    .B(_01598_),
    .C(_01578_),
    .Y(_01599_));
 sg13g2_nand2_1 _16791_ (.Y(_01600_),
    .A(_01599_),
    .B(_01570_));
 sg13g2_nand2_1 _16792_ (.Y(_01601_),
    .A(_01597_),
    .B(_01600_));
 sg13g2_nand2_1 _16793_ (.Y(_01602_),
    .A(_01601_),
    .B(_01779_));
 sg13g2_nand3_1 _16794_ (.B(_01780_),
    .C(_01600_),
    .A(_01597_),
    .Y(_01603_));
 sg13g2_nand3_1 _16795_ (.B(_01603_),
    .C(_01739_),
    .A(_01602_),
    .Y(_01604_));
 sg13g2_nand2b_1 _16796_ (.Y(_01605_),
    .B(net202),
    .A_N(_00163_));
 sg13g2_a21oi_1 _16797_ (.A1(_01604_),
    .A2(_01605_),
    .Y(_01606_),
    .B1(_03411_));
 sg13g2_nand3_1 _16798_ (.B(_03411_),
    .C(_01605_),
    .A(_01604_),
    .Y(_01607_));
 sg13g2_inv_1 _16799_ (.Y(_01608_),
    .A(_01607_));
 sg13g2_nor2_1 _16800_ (.A(_01606_),
    .B(_01608_),
    .Y(_01609_));
 sg13g2_xnor2_1 _16801_ (.Y(\synth.voice.rshift[0] ),
    .A(_01539_),
    .B(_01609_));
 sg13g2_nor2b_1 _16802_ (.A(_01609_),
    .B_N(_01539_),
    .Y(_01610_));
 sg13g2_nand2_1 _16803_ (.Y(_01611_),
    .A(_01786_),
    .B(_01758_));
 sg13g2_nand2_1 _16804_ (.Y(_01612_),
    .A(_01603_),
    .B(_01611_));
 sg13g2_inv_1 _16805_ (.Y(_01613_),
    .A(_01611_));
 sg13g2_nand4_1 _16806_ (.B(_01780_),
    .C(_01600_),
    .A(_01597_),
    .Y(_01614_),
    .D(_01613_));
 sg13g2_nand2_1 _16807_ (.Y(_01615_),
    .A(_01612_),
    .B(_01614_));
 sg13g2_nand2_1 _16808_ (.Y(_01616_),
    .A(_01615_),
    .B(_01739_));
 sg13g2_nand2_1 _16809_ (.Y(_01617_),
    .A(net202),
    .B(_00171_));
 sg13g2_nand2_1 _16810_ (.Y(_01618_),
    .A(_01616_),
    .B(_01617_));
 sg13g2_nand2_1 _16811_ (.Y(_01619_),
    .A(_01608_),
    .B(_01618_));
 sg13g2_inv_1 _16812_ (.Y(_01620_),
    .A(_01617_));
 sg13g2_a21oi_1 _16813_ (.A1(_01615_),
    .A2(_01764_),
    .Y(_01621_),
    .B1(_01620_));
 sg13g2_nand2_1 _16814_ (.Y(_01622_),
    .A(_01621_),
    .B(_01607_));
 sg13g2_inv_1 _16815_ (.Y(_01623_),
    .A(_00172_));
 sg13g2_nand2_1 _16816_ (.Y(_01624_),
    .A(_01529_),
    .B(_00173_));
 sg13g2_a22oi_1 _16817_ (.Y(_01625_),
    .B1(_03917_),
    .B2(_01535_),
    .A2(_01534_),
    .A1(\synth.voice.genblk4[7].next_state_scan[13] ));
 sg13g2_a21oi_1 _16818_ (.A1(_01625_),
    .A2(_01546_),
    .Y(_01626_),
    .B1(net202));
 sg13g2_a22oi_1 _16819_ (.Y(_01627_),
    .B1(_01624_),
    .B2(_01626_),
    .A2(net202),
    .A1(_01623_));
 sg13g2_a21oi_1 _16820_ (.A1(_01619_),
    .A2(_01622_),
    .Y(_01628_),
    .B1(_01627_));
 sg13g2_nand3_1 _16821_ (.B(_01622_),
    .C(_01627_),
    .A(_01619_),
    .Y(_01629_));
 sg13g2_nor2b_1 _16822_ (.A(_01628_),
    .B_N(_01629_),
    .Y(_01630_));
 sg13g2_xor2_1 _16823_ (.B(_01630_),
    .A(_01610_),
    .X(\synth.voice.rshift[1] ));
 sg13g2_a21oi_1 _16824_ (.A1(_01604_),
    .A2(_01605_),
    .Y(_01631_),
    .B1(_03412_));
 sg13g2_nand2_1 _16825_ (.Y(_01632_),
    .A(_01631_),
    .B(_01618_));
 sg13g2_nand2b_1 _16826_ (.Y(_01633_),
    .B(_01764_),
    .A_N(_01614_));
 sg13g2_nand3_1 _16827_ (.B(_03669_),
    .C(_01617_),
    .A(_01616_),
    .Y(_01634_));
 sg13g2_nand3_1 _16828_ (.B(_01633_),
    .C(_01634_),
    .A(_01632_),
    .Y(_01635_));
 sg13g2_nor2b_1 _16829_ (.A(net201),
    .B_N(_00174_),
    .Y(_01636_));
 sg13g2_inv_1 _16830_ (.Y(_01637_),
    .A(_00059_));
 sg13g2_a22oi_1 _16831_ (.Y(_01638_),
    .B1(_03902_),
    .B2(_01535_),
    .A2(_01534_),
    .A1(_01637_));
 sg13g2_nand2b_1 _16832_ (.Y(_01639_),
    .B(_01529_),
    .A_N(_00175_));
 sg13g2_nand3_1 _16833_ (.B(_01739_),
    .C(_01639_),
    .A(_01638_),
    .Y(_01640_));
 sg13g2_nand2b_1 _16834_ (.Y(_01641_),
    .B(_01640_),
    .A_N(_01636_));
 sg13g2_inv_1 _16835_ (.Y(_01642_),
    .A(_01641_));
 sg13g2_nand2_1 _16836_ (.Y(_01643_),
    .A(_01635_),
    .B(_01642_));
 sg13g2_nand4_1 _16837_ (.B(_01634_),
    .C(_01633_),
    .A(_01632_),
    .Y(_01644_),
    .D(_01641_));
 sg13g2_nand2_1 _16838_ (.Y(_01645_),
    .A(_01643_),
    .B(_01644_));
 sg13g2_a21oi_1 _16839_ (.A1(_01629_),
    .A2(_01610_),
    .Y(_01646_),
    .B1(_01628_));
 sg13g2_xor2_1 _16840_ (.B(_01646_),
    .A(_01645_),
    .X(\synth.voice.rshift[2] ));
 sg13g2_inv_1 _16841_ (.Y(_01647_),
    .A(_00177_));
 sg13g2_nor2_1 _16842_ (.A(_00147_),
    .B(net164),
    .Y(_01648_));
 sg13g2_a21oi_1 _16843_ (.A1(\synth.voice.genblk4[7].next_state_scan[5] ),
    .A2(net164),
    .Y(_01649_),
    .B1(_01648_));
 sg13g2_a21oi_1 _16844_ (.A1(_01546_),
    .A2(_01649_),
    .Y(_01650_),
    .B1(net202));
 sg13g2_o21ai_1 _16845_ (.B1(_01650_),
    .Y(_01651_),
    .A1(_01647_),
    .A2(net129));
 sg13g2_o21ai_1 _16846_ (.B1(_01651_),
    .Y(_01652_),
    .A1(_00176_),
    .A2(net201));
 sg13g2_nor2b_1 _16847_ (.A(_01645_),
    .B_N(_01652_),
    .Y(_01653_));
 sg13g2_nand2b_1 _16848_ (.Y(_01654_),
    .B(_01653_),
    .A_N(_01646_));
 sg13g2_inv_1 _16849_ (.Y(_01655_),
    .A(_01643_));
 sg13g2_nand2_1 _16850_ (.Y(_01656_),
    .A(_01655_),
    .B(_01652_));
 sg13g2_nand2_1 _16851_ (.Y(\synth.voice.zero_shifter_out ),
    .A(_01654_),
    .B(_01656_));
 sg13g2_nor2_1 _16852_ (.A(_01645_),
    .B(_01646_),
    .Y(_01657_));
 sg13g2_nor3_1 _16853_ (.A(_01655_),
    .B(_01652_),
    .C(_01657_),
    .Y(_01658_));
 sg13g2_nor2_1 _16854_ (.A(\synth.voice.zero_shifter_out ),
    .B(_01658_),
    .Y(\synth.voice.rshift[3] ));
 sg13g2_nand2_1 _16855_ (.Y(_01659_),
    .A(_01749_),
    .B(_01791_));
 sg13g2_nand2_1 _16856_ (.Y(_01660_),
    .A(_01735_),
    .B(_01726_));
 sg13g2_nand3_1 _16857_ (.B(_01659_),
    .C(_01660_),
    .A(net192),
    .Y(\synth.voice.scan_accs ));
 sg13g2_nand2_1 _16858_ (.Y(_01661_),
    .A(_06511_),
    .B(_02272_));
 sg13g2_a21oi_1 _16859_ (.A1(_01661_),
    .A2(\ppu_ctrl[4] ),
    .Y(\uio_out0[6] ),
    .B1(net389));
 sg13g2_nand3_1 _16860_ (.B(_06519_),
    .C(\ppu_ctrl[4] ),
    .A(_02284_),
    .Y(_01662_));
 sg13g2_nand2b_1 _16861_ (.Y(_01663_),
    .B(_07677_),
    .A_N(\ppu_ctrl[4] ));
 sg13g2_a21oi_1 _16862_ (.A1(_01662_),
    .A2(_01663_),
    .Y(\uio_out0[7] ),
    .B1(_06089_));
 sg13g2_inv_1 _16863_ (.Y(_01664_),
    .A(_00157_));
 sg13g2_o21ai_1 _16864_ (.B1(_00152_),
    .Y(_01665_),
    .A1(\ppu.b0_out[1] ),
    .A2(_01664_));
 sg13g2_a21oi_1 _16865_ (.A1(_01665_),
    .A2(_06500_),
    .Y(_01666_),
    .B1(\ppu.dither_r.u[2] ));
 sg13g2_inv_1 _16866_ (.Y(_01667_),
    .A(_01666_));
 sg13g2_nor2_1 _16867_ (.A(_06519_),
    .B(_06500_),
    .Y(_01668_));
 sg13g2_inv_1 _16868_ (.Y(_01669_),
    .A(_01668_));
 sg13g2_nand2_1 _16869_ (.Y(_01670_),
    .A(net396),
    .B(_06500_));
 sg13g2_nand3_1 _16870_ (.B(_01669_),
    .C(_01670_),
    .A(_01667_),
    .Y(_01671_));
 sg13g2_o21ai_1 _16871_ (.B1(_01671_),
    .Y(_01672_),
    .A1(_01664_),
    .A2(_01667_));
 sg13g2_inv_1 _16872_ (.Y(_01673_),
    .A(_01865_));
 sg13g2_nand3_1 _16873_ (.B(_01673_),
    .C(net396),
    .A(net294),
    .Y(_01674_));
 sg13g2_xor2_1 _16874_ (.B(_01865_),
    .A(_01854_),
    .X(_01675_));
 sg13g2_buf_1 _16875_ (.A(_01675_),
    .X(_01676_));
 sg13g2_nand2_1 _16876_ (.Y(_01677_),
    .A(_01673_),
    .B(net396));
 sg13g2_a22oi_1 _16877_ (.Y(_01678_),
    .B1(_01676_),
    .B2(_01677_),
    .A2(_00158_),
    .A1(_01674_));
 sg13g2_nor3_1 _16878_ (.A(net396),
    .B(_01676_),
    .C(_01666_),
    .Y(_01679_));
 sg13g2_a21o_1 _16879_ (.A2(_01678_),
    .A1(_01666_),
    .B1(_01679_),
    .X(_01680_));
 sg13g2_nand2b_1 _16880_ (.Y(_01681_),
    .B(_01680_),
    .A_N(_01672_));
 sg13g2_a21oi_1 _16881_ (.A1(_01669_),
    .A2(\ppu.dither_r.u[2] ),
    .Y(_01682_),
    .B1(_07067_));
 sg13g2_a221oi_1 _16882_ (.B2(_01682_),
    .C1(net389),
    .B1(_01681_),
    .A1(_06502_),
    .Y(\uo_out0[0] ),
    .A2(_07067_));
 sg13g2_nor2_1 _16883_ (.A(\ppu.dither_g.u[2] ),
    .B(_06514_),
    .Y(_01683_));
 sg13g2_nor3_1 _16884_ (.A(_06511_),
    .B(_01683_),
    .C(_01676_),
    .Y(_01684_));
 sg13g2_o21ai_1 _16885_ (.B1(_01676_),
    .Y(_01685_),
    .A1(_01865_),
    .A2(_06512_));
 sg13g2_nand3_1 _16886_ (.B(_01673_),
    .C(_06511_),
    .A(net294),
    .Y(_01686_));
 sg13g2_nand2_1 _16887_ (.Y(_01687_),
    .A(_01686_),
    .B(_00156_));
 sg13g2_nand3_1 _16888_ (.B(_01683_),
    .C(_01687_),
    .A(_01685_),
    .Y(_01688_));
 sg13g2_nand2b_1 _16889_ (.Y(_01689_),
    .B(_01688_),
    .A_N(_01684_));
 sg13g2_nand2_1 _16890_ (.Y(_01690_),
    .A(_06511_),
    .B(_06514_));
 sg13g2_a21oi_1 _16891_ (.A1(_06512_),
    .A2(_06515_),
    .Y(_01691_),
    .B1(_01683_));
 sg13g2_a22oi_1 _16892_ (.Y(_01692_),
    .B1(_01690_),
    .B2(_01691_),
    .A2(_01683_),
    .A1(_00155_));
 sg13g2_a21oi_1 _16893_ (.A1(_01689_),
    .A2(_01692_),
    .Y(_01693_),
    .B1(_07067_));
 sg13g2_o21ai_1 _16894_ (.B1(\ppu.dither_g.u[2] ),
    .Y(_01694_),
    .A1(_06511_),
    .A2(_06514_));
 sg13g2_a221oi_1 _16895_ (.B2(_01694_),
    .C1(net389),
    .B1(_01693_),
    .A1(_06517_),
    .Y(\uo_out0[1] ),
    .A2(_07067_));
 sg13g2_inv_1 _16896_ (.Y(_01695_),
    .A(_00153_));
 sg13g2_o21ai_1 _16897_ (.B1(_00152_),
    .Y(_01696_),
    .A1(net396),
    .A2(_01695_));
 sg13g2_a21oi_2 _16898_ (.B1(\ppu.b0_out[3] ),
    .Y(_01697_),
    .A2(_06506_),
    .A1(_01696_));
 sg13g2_inv_1 _16899_ (.Y(_01698_),
    .A(_01697_));
 sg13g2_o21ai_1 _16900_ (.B1(_01698_),
    .Y(_01699_),
    .A1(net396),
    .A2(_01676_));
 sg13g2_nand3_1 _16901_ (.B(_00154_),
    .C(_01677_),
    .A(_01697_),
    .Y(_01700_));
 sg13g2_o21ai_1 _16902_ (.B1(_01676_),
    .Y(_01701_),
    .A1(_00154_),
    .A2(_01677_));
 sg13g2_nand3_1 _16903_ (.B(_01700_),
    .C(_01701_),
    .A(_01699_),
    .Y(_01702_));
 sg13g2_xnor2_1 _16904_ (.Y(_01703_),
    .A(net396),
    .B(_06506_));
 sg13g2_nor2_1 _16905_ (.A(_01703_),
    .B(_01697_),
    .Y(_01704_));
 sg13g2_a21oi_1 _16906_ (.A1(_00153_),
    .A2(_01697_),
    .Y(_01705_),
    .B1(_01704_));
 sg13g2_nand2b_1 _16907_ (.Y(_01706_),
    .B(_01705_),
    .A_N(_01702_));
 sg13g2_nand2_1 _16908_ (.Y(_01707_),
    .A(_06520_),
    .B(_06507_));
 sg13g2_a21oi_1 _16909_ (.A1(_01707_),
    .A2(\ppu.b0_out[3] ),
    .Y(_01708_),
    .B1(_07067_));
 sg13g2_a221oi_1 _16910_ (.B2(_01708_),
    .C1(net389),
    .B1(_01706_),
    .A1(_06509_),
    .Y(\uo_out0[2] ),
    .A2(_07067_));
 sg13g2_xor2_1 _16911_ (.B(_01680_),
    .A(_01672_),
    .X(_01709_));
 sg13g2_o21ai_1 _16912_ (.B1(_02284_),
    .Y(_01710_),
    .A1(_06500_),
    .A2(_07066_));
 sg13g2_a21oi_1 _16913_ (.A1(_01709_),
    .A2(_07066_),
    .Y(\uo_out0[4] ),
    .B1(_01710_));
 sg13g2_xnor2_1 _16914_ (.Y(_01711_),
    .A(_01692_),
    .B(_01689_));
 sg13g2_o21ai_1 _16915_ (.B1(_02284_),
    .Y(_01712_),
    .A1(_06514_),
    .A2(_07066_));
 sg13g2_a21oi_1 _16916_ (.A1(_01711_),
    .A2(_07066_),
    .Y(\uo_out0[5] ),
    .B1(_01712_));
 sg13g2_xor2_1 _16917_ (.B(_01702_),
    .A(_01705_),
    .X(_01713_));
 sg13g2_o21ai_1 _16918_ (.B1(_02284_),
    .Y(_01714_),
    .A1(_06506_),
    .A2(_07066_));
 sg13g2_a21oi_1 _16919_ (.A1(_01713_),
    .A2(_07066_),
    .Y(\uo_out0[6] ),
    .B1(_01714_));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_1 _16921_ (.A(net410),
    .X(uio_oe[0]));
 sg13g2_buf_1 _16922_ (.A(net411),
    .X(uio_oe[1]));
 sg13g2_buf_1 _16923_ (.A(net412),
    .X(uio_oe[2]));
 sg13g2_buf_1 _16924_ (.A(net413),
    .X(uio_oe[3]));
 sg13g2_buf_1 _16925_ (.A(net414),
    .X(uio_oe[4]));
 sg13g2_buf_1 _16926_ (.A(net415),
    .X(uio_oe[5]));
 sg13g2_buf_1 _16927_ (.A(drive_uio_76),
    .X(net10));
 sg13g2_buf_1 _16928_ (.A(drive_uio_76),
    .X(net11));
 sg13g2_dfrbp_1 \cfg[0]$_DFFE_PN_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net416),
    .D(_00183_),
    .Q_N(_08992_),
    .Q(drive_uio_76));
 sg13g2_dfrbp_1 \ppu.avhsync_delayed[0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net417),
    .D(_00184_),
    .Q_N(_08991_),
    .Q(hsync));
 sg13g2_dfrbp_1 \ppu.avhsync_delayed[1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net418),
    .D(_00185_),
    .Q_N(_08990_),
    .Q(\ppu.vsync ));
 sg13g2_dfrbp_1 \ppu.avhsync_delayed[2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net419),
    .D(_00186_),
    .Q_N(_08989_),
    .Q(active));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net420),
    .D(_00187_),
    .Q_N(_08988_),
    .Q(\ppu.base_addr_regs[0][0] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net421),
    .D(_00188_),
    .Q_N(_08987_),
    .Q(\ppu.base_addr_regs[0][1] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net422),
    .D(_00189_),
    .Q_N(_08986_),
    .Q(\ppu.base_addr_regs[0][2] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net423),
    .D(_00190_),
    .Q_N(_08985_),
    .Q(\ppu.base_addr_regs[0][3] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net424),
    .D(_00191_),
    .Q_N(_08984_),
    .Q(\ppu.base_addr_regs[0][4] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net425),
    .D(_00192_),
    .Q_N(_08983_),
    .Q(\ppu.base_addr_regs[0][5] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net426),
    .D(_00193_),
    .Q_N(_08982_),
    .Q(\ppu.base_addr_regs[0][6] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net427),
    .D(_00194_),
    .Q_N(_08981_),
    .Q(\ppu.base_addr_regs[0][7] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net428),
    .D(_00195_),
    .Q_N(_08980_),
    .Q(\ppu.base_addr_regs[0][8] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net429),
    .D(_00196_),
    .Q_N(_08979_),
    .Q(\ppu.base_addr_regs[1][0] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net430),
    .D(_00197_),
    .Q_N(_08978_),
    .Q(\ppu.base_addr_regs[1][1] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net431),
    .D(_00198_),
    .Q_N(_08977_),
    .Q(\ppu.base_addr_regs[1][2] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net432),
    .D(_00199_),
    .Q_N(_08976_),
    .Q(\ppu.base_addr_regs[1][3] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net433),
    .D(_00200_),
    .Q_N(_08975_),
    .Q(\ppu.base_addr_regs[1][4] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net434),
    .D(_00201_),
    .Q_N(_08974_),
    .Q(\ppu.base_addr_regs[1][5] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net435),
    .D(_00202_),
    .Q_N(_08973_),
    .Q(\ppu.base_addr_regs[1][6] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net436),
    .D(_00203_),
    .Q_N(_08972_),
    .Q(\ppu.base_addr_regs[1][7] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net437),
    .D(_00204_),
    .Q_N(_08971_),
    .Q(\ppu.base_addr_regs[1][8] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net438),
    .D(_00205_),
    .Q_N(_08970_),
    .Q(\ppu.base_addr_regs[2][1] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net439),
    .D(_00206_),
    .Q_N(_08969_),
    .Q(\ppu.base_addr_regs[2][2] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net440),
    .D(_00207_),
    .Q_N(_08968_),
    .Q(\ppu.base_addr_regs[2][3] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net441),
    .D(_00208_),
    .Q_N(_08967_),
    .Q(\ppu.base_addr_regs[2][4] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net442),
    .D(_00209_),
    .Q_N(_08966_),
    .Q(\ppu.base_addr_regs[2][5] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net443),
    .D(_00210_),
    .Q_N(_08965_),
    .Q(\ppu.base_addr_regs[2][6] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net444),
    .D(_00211_),
    .Q_N(_08964_),
    .Q(\ppu.base_addr_regs[2][7] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net445),
    .D(_00212_),
    .Q_N(_08963_),
    .Q(\ppu.base_addr_regs[2][8] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net446),
    .D(_00213_),
    .Q_N(_08962_),
    .Q(\ppu.base_addr_regs[3][1] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net447),
    .D(_00214_),
    .Q_N(_08961_),
    .Q(\ppu.base_addr_regs[3][2] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net448),
    .D(_00215_),
    .Q_N(_08960_),
    .Q(\ppu.base_addr_regs[3][3] ));
 sg13g2_dfrbp_1 \ppu.base_addr_regs[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net449),
    .D(_00216_),
    .Q_N(_08959_),
    .Q(\ppu.base_addr_regs[3][4] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[0]$_SDFF_PP0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net450),
    .D(_00217_),
    .Q_N(_00131_),
    .Q(\ppu.copper_inst.addr[0] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[10]$_SDFF_PP1_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net451),
    .D(_00218_),
    .Q_N(_08958_),
    .Q(\ppu.copper_inst.addr[10] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[11]$_SDFF_PP1_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net452),
    .D(_00219_),
    .Q_N(_08957_),
    .Q(\ppu.copper_inst.addr[11] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[12]$_SDFF_PP1_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net453),
    .D(_00220_),
    .Q_N(_08956_),
    .Q(\ppu.copper_inst.addr[12] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[13]$_SDFF_PP1_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net454),
    .D(_00221_),
    .Q_N(_08955_),
    .Q(\ppu.copper_inst.addr[13] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[14]$_SDFF_PP1_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net455),
    .D(_00222_),
    .Q_N(_08954_),
    .Q(\ppu.copper_inst.addr[14] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[15]$_SDFF_PP1_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net456),
    .D(_00223_),
    .Q_N(_08953_),
    .Q(\ppu.copper_inst.addr[15] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[1]$_SDFF_PP1_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net457),
    .D(_00224_),
    .Q_N(_00132_),
    .Q(\ppu.copper_inst.addr[1] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[2]$_SDFF_PP1_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net458),
    .D(_00225_),
    .Q_N(_08952_),
    .Q(\ppu.copper_inst.addr[2] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[3]$_SDFF_PP1_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net459),
    .D(_00226_),
    .Q_N(_08951_),
    .Q(\ppu.copper_inst.addr[3] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[4]$_SDFF_PP1_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net460),
    .D(_00227_),
    .Q_N(_08950_),
    .Q(\ppu.copper_inst.addr[4] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[5]$_SDFF_PP1_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net461),
    .D(_00228_),
    .Q_N(_08949_),
    .Q(\ppu.copper_inst.addr[5] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[6]$_SDFF_PP1_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net462),
    .D(_00229_),
    .Q_N(_08948_),
    .Q(\ppu.copper_inst.addr[6] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[7]$_SDFF_PP1_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net463),
    .D(_00230_),
    .Q_N(_08947_),
    .Q(\ppu.copper_inst.addr[7] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[8]$_SDFF_PP1_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net464),
    .D(_00231_),
    .Q_N(_08946_),
    .Q(\ppu.copper_inst.addr[8] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.addr_reg[9]$_SDFF_PP1_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net465),
    .D(_00232_),
    .Q_N(_08945_),
    .Q(\ppu.copper_inst.addr[9] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net466),
    .D(_00233_),
    .Q_N(_08944_),
    .Q(\ppu.copper_inst.cmp[0] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net467),
    .D(_00234_),
    .Q_N(_08943_),
    .Q(\ppu.copper_inst.cmp[1] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net468),
    .D(_00235_),
    .Q_N(_08942_),
    .Q(\ppu.copper_inst.cmp[2] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net469),
    .D(_00236_),
    .Q_N(_08941_),
    .Q(\ppu.copper_inst.cmp[3] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net470),
    .D(_00237_),
    .Q_N(_08940_),
    .Q(\ppu.copper_inst.cmp[4] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net471),
    .D(_00238_),
    .Q_N(_08939_),
    .Q(\ppu.copper_inst.cmp[5] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net472),
    .D(_00239_),
    .Q_N(_08938_),
    .Q(\ppu.copper_inst.cmp[6] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net473),
    .D(_00240_),
    .Q_N(_08937_),
    .Q(\ppu.copper_inst.cmp[7] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net474),
    .D(_00241_),
    .Q_N(_00039_),
    .Q(\ppu.copper_inst.cmp[8] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp_on$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net475),
    .D(_00242_),
    .Q_N(_08936_),
    .Q(\ppu.copper_inst.cmp_on ));
 sg13g2_dfrbp_1 \ppu.copper_inst.cmp_type$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net476),
    .D(_00243_),
    .Q_N(_08993_),
    .Q(\ppu.copper_inst.cmp_type ));
 sg13g2_dfrbp_1 \ppu.copper_inst.fast_mode$_DFF_P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net477),
    .D(_00014_),
    .Q_N(_08935_),
    .Q(\ppu.copper_inst.fast_mode ));
 sg13g2_dfrbp_1 \ppu.copper_inst.on$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net478),
    .D(_00244_),
    .Q_N(_08934_),
    .Q(\ppu.copper_inst.on ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net479),
    .D(_00245_),
    .Q_N(_08933_),
    .Q(\ppu.copper_inst.store[0] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[10]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net480),
    .D(_00246_),
    .Q_N(_08932_),
    .Q(\ppu.copper_inst.store[10] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[11]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net481),
    .D(_00247_),
    .Q_N(_08931_),
    .Q(\ppu.copper_inst.store[11] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[12]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net482),
    .D(_00248_),
    .Q_N(_08930_),
    .Q(\ppu.copper_inst.store[12] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[13]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net483),
    .D(_00249_),
    .Q_N(_08929_),
    .Q(\ppu.copper_inst.store[13] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[14]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net484),
    .D(_00250_),
    .Q_N(_08928_),
    .Q(\ppu.copper_inst.store[14] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[15]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net485),
    .D(_00251_),
    .Q_N(_08927_),
    .Q(\ppu.copper_inst.store[15] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[1]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net486),
    .D(_00252_),
    .Q_N(_08926_),
    .Q(\ppu.copper_inst.store[1] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net487),
    .D(_00253_),
    .Q_N(_08925_),
    .Q(\ppu.copper_inst.store[2] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[3]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net488),
    .D(_00254_),
    .Q_N(_08924_),
    .Q(\ppu.copper_inst.store[3] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[4]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net489),
    .D(_00255_),
    .Q_N(_08923_),
    .Q(\ppu.copper_inst.store[4] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[5]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net490),
    .D(_00256_),
    .Q_N(_08922_),
    .Q(\ppu.copper_inst.store[5] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[6]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net491),
    .D(_00257_),
    .Q_N(_08921_),
    .Q(\ppu.copper_inst.store[6] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[7]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net492),
    .D(_00258_),
    .Q_N(_08920_),
    .Q(\ppu.copper_inst.store[7] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[8]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net493),
    .D(_00259_),
    .Q_N(_08919_),
    .Q(\ppu.copper_inst.store[8] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store[9]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net494),
    .D(_00260_),
    .Q_N(_08918_),
    .Q(\ppu.copper_inst.store[9] ));
 sg13g2_dfrbp_1 \ppu.copper_inst.store_valid$_SDFFCE_PP0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net495),
    .D(_00261_),
    .Q_N(_00076_),
    .Q(\ppu.copper_inst.store_valid ));
 sg13g2_dfrbp_1 \ppu.curr_pal_addr[0]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net496),
    .D(_00262_),
    .Q_N(_08917_),
    .Q(\ppu.curr_pal_addr[0] ));
 sg13g2_dfrbp_1 \ppu.curr_pal_addr[1]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net497),
    .D(_00263_),
    .Q_N(_08916_),
    .Q(\ppu.curr_pal_addr[1] ));
 sg13g2_dfrbp_1 \ppu.curr_pal_addr[2]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net498),
    .D(_00264_),
    .Q_N(_08915_),
    .Q(\ppu.curr_pal_addr[2] ));
 sg13g2_dfrbp_1 \ppu.curr_pal_addr[3]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net499),
    .D(_00265_),
    .Q_N(_08914_),
    .Q(\ppu.curr_pal_addr[3] ));
 sg13g2_dfrbp_1 \ppu.display_mask[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net500),
    .D(_00266_),
    .Q_N(_08913_),
    .Q(\ppu.display_mask[0] ));
 sg13g2_dfrbp_1 \ppu.display_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net501),
    .D(_00267_),
    .Q_N(_08912_),
    .Q(\ppu.display_mask[1] ));
 sg13g2_dfrbp_1 \ppu.display_mask[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net502),
    .D(_00268_),
    .Q_N(_08911_),
    .Q(\ppu.display_mask[2] ));
 sg13g2_dfrbp_1 \ppu.display_mask[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net503),
    .D(_00269_),
    .Q_N(_08910_),
    .Q(\ppu.display_mask[3] ));
 sg13g2_dfrbp_1 \ppu.display_mask[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net504),
    .D(_00270_),
    .Q_N(_08909_),
    .Q(\ppu.display_mask[4] ));
 sg13g2_dfrbp_1 \ppu.display_mask[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net505),
    .D(_00271_),
    .Q_N(_08908_),
    .Q(\ppu.display_mask[5] ));
 sg13g2_dfrbp_1 \ppu.gfxmode1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net506),
    .D(_00272_),
    .Q_N(_08907_),
    .Q(\ppu.gfxmode1[0] ));
 sg13g2_dfrbp_1 \ppu.gfxmode1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net507),
    .D(_00273_),
    .Q_N(_08906_),
    .Q(\ppu.gfxmode1[1] ));
 sg13g2_dfrbp_1 \ppu.gfxmode1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net508),
    .D(_00274_),
    .Q_N(_08905_),
    .Q(\ppu.gfxmode1[2] ));
 sg13g2_dfrbp_1 \ppu.gfxmode1[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net509),
    .D(_00275_),
    .Q_N(_08904_),
    .Q(\ppu.gfxmode1[3] ));
 sg13g2_dfrbp_1 \ppu.gfxmode1[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net510),
    .D(_00276_),
    .Q_N(_08903_),
    .Q(\ppu.gfxmode1[4] ));
 sg13g2_dfrbp_1 \ppu.gfxmode1[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net511),
    .D(_00277_),
    .Q_N(_08902_),
    .Q(\ppu.gfxmode1[5] ));
 sg13g2_dfrbp_1 \ppu.gfxmode1[6]$_SDFFE_PN1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net512),
    .D(_00278_),
    .Q_N(_08901_),
    .Q(\ppu.gfxmode1[6] ));
 sg13g2_dfrbp_1 \ppu.gfxmode1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net513),
    .D(_00279_),
    .Q_N(_08900_),
    .Q(\ppu.gfxmode1[7] ));
 sg13g2_dfrbp_1 \ppu.gfxmode1[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net514),
    .D(_00280_),
    .Q_N(_08899_),
    .Q(\ppu.gfxmode1[8] ));
 sg13g2_dfrbp_1 \ppu.gfxmode2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net515),
    .D(_00281_),
    .Q_N(_08898_),
    .Q(\ppu.gfxmode2[0] ));
 sg13g2_dfrbp_1 \ppu.gfxmode2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net516),
    .D(_00282_),
    .Q_N(_08897_),
    .Q(\ppu.gfxmode2[1] ));
 sg13g2_dfrbp_1 \ppu.gfxmode2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net517),
    .D(_00283_),
    .Q_N(_08896_),
    .Q(\ppu.gfxmode2[2] ));
 sg13g2_dfrbp_1 \ppu.gfxmode2[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net518),
    .D(_00284_),
    .Q_N(_08895_),
    .Q(\ppu.gfxmode2[3] ));
 sg13g2_dfrbp_1 \ppu.gfxmode2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net519),
    .D(_00285_),
    .Q_N(_08894_),
    .Q(\ppu.gfxmode2[4] ));
 sg13g2_dfrbp_1 \ppu.gfxmode2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net520),
    .D(_00286_),
    .Q_N(_08893_),
    .Q(\ppu.gfxmode2[5] ));
 sg13g2_dfrbp_1 \ppu.gfxmode2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net521),
    .D(_00287_),
    .Q_N(_08892_),
    .Q(\ppu.gfxmode2[6] ));
 sg13g2_dfrbp_1 \ppu.gfxmode2[7]$_SDFFE_PN1P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net522),
    .D(_00288_),
    .Q_N(_08891_),
    .Q(\ppu.gfxmode2[7] ));
 sg13g2_dfrbp_1 \ppu.gfxmode2[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net523),
    .D(_00289_),
    .Q_N(_08890_),
    .Q(\ppu.gfxmode2[8] ));
 sg13g2_dfrbp_1 \ppu.gfxmode3[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net524),
    .D(_00290_),
    .Q_N(_08889_),
    .Q(\ppu.gfxmode3[0] ));
 sg13g2_dfrbp_1 \ppu.gfxmode3[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net525),
    .D(_00291_),
    .Q_N(_08888_),
    .Q(\ppu.gfxmode3[1] ));
 sg13g2_dfrbp_1 \ppu.gfxmode3[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net526),
    .D(_00292_),
    .Q_N(_08887_),
    .Q(\ppu.gfxmode3[2] ));
 sg13g2_dfrbp_1 \ppu.gfxmode3[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net527),
    .D(_00293_),
    .Q_N(_08886_),
    .Q(\ppu.gfxmode3[3] ));
 sg13g2_dfrbp_1 \ppu.gfxmode3[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net528),
    .D(_00294_),
    .Q_N(_08885_),
    .Q(\ppu.gfxmode3[4] ));
 sg13g2_dfrbp_1 \ppu.gfxmode3[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net529),
    .D(_00295_),
    .Q_N(_08884_),
    .Q(\ppu.gfxmode3[5] ));
 sg13g2_dfrbp_1 \ppu.gfxmode3[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net530),
    .D(_00296_),
    .Q_N(_08883_),
    .Q(\ppu.gfxmode3[6] ));
 sg13g2_dfrbp_1 \ppu.gfxmode3[7]$_SDFFE_PN1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net531),
    .D(_00297_),
    .Q_N(_08882_),
    .Q(\ppu.gfxmode3[7] ));
 sg13g2_dfrbp_1 \ppu.gfxmode3[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net532),
    .D(_00298_),
    .Q_N(_08881_),
    .Q(\ppu.gfxmode3[8] ));
 sg13g2_dfrbp_1 \ppu.pal[0][0]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net533),
    .D(_00299_),
    .Q_N(_08880_),
    .Q(\ppu.pal[0][0] ));
 sg13g2_dfrbp_1 \ppu.pal[0][1]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net534),
    .D(_00300_),
    .Q_N(_08879_),
    .Q(\ppu.pal[0][1] ));
 sg13g2_dfrbp_1 \ppu.pal[0][2]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net535),
    .D(_00301_),
    .Q_N(_08878_),
    .Q(\ppu.pal[0][2] ));
 sg13g2_dfrbp_1 \ppu.pal[0][3]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net536),
    .D(_00302_),
    .Q_N(_08877_),
    .Q(\ppu.pal[0][3] ));
 sg13g2_dfrbp_1 \ppu.pal[0][4]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net537),
    .D(_00303_),
    .Q_N(_08876_),
    .Q(\ppu.pal[0][4] ));
 sg13g2_dfrbp_1 \ppu.pal[0][5]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net538),
    .D(_00304_),
    .Q_N(_08875_),
    .Q(\ppu.pal[0][5] ));
 sg13g2_dfrbp_1 \ppu.pal[0][6]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net539),
    .D(_00305_),
    .Q_N(_08874_),
    .Q(\ppu.pal[0][6] ));
 sg13g2_dfrbp_1 \ppu.pal[0][7]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net540),
    .D(_00306_),
    .Q_N(_08873_),
    .Q(\ppu.pal[0][7] ));
 sg13g2_dfrbp_1 \ppu.pal[10][0]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net541),
    .D(_00307_),
    .Q_N(_08872_),
    .Q(\ppu.pal[10][0] ));
 sg13g2_dfrbp_1 \ppu.pal[10][1]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net542),
    .D(_00308_),
    .Q_N(_08871_),
    .Q(\ppu.pal[10][1] ));
 sg13g2_dfrbp_1 \ppu.pal[10][2]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net543),
    .D(_00309_),
    .Q_N(_08870_),
    .Q(\ppu.pal[10][2] ));
 sg13g2_dfrbp_1 \ppu.pal[10][3]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net544),
    .D(_00310_),
    .Q_N(_08869_),
    .Q(\ppu.pal[10][3] ));
 sg13g2_dfrbp_1 \ppu.pal[10][4]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net545),
    .D(_00311_),
    .Q_N(_08868_),
    .Q(\ppu.pal[10][4] ));
 sg13g2_dfrbp_1 \ppu.pal[10][5]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net546),
    .D(_00312_),
    .Q_N(_08867_),
    .Q(\ppu.pal[10][5] ));
 sg13g2_dfrbp_1 \ppu.pal[10][6]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net547),
    .D(_00313_),
    .Q_N(_08866_),
    .Q(\ppu.pal[10][6] ));
 sg13g2_dfrbp_1 \ppu.pal[10][7]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net548),
    .D(_00314_),
    .Q_N(_08865_),
    .Q(\ppu.pal[10][7] ));
 sg13g2_dfrbp_1 \ppu.pal[11][0]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net549),
    .D(_00315_),
    .Q_N(_08864_),
    .Q(\ppu.pal[11][0] ));
 sg13g2_dfrbp_1 \ppu.pal[11][1]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net550),
    .D(_00316_),
    .Q_N(_08863_),
    .Q(\ppu.pal[11][1] ));
 sg13g2_dfrbp_1 \ppu.pal[11][2]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net551),
    .D(_00317_),
    .Q_N(_08862_),
    .Q(\ppu.pal[11][2] ));
 sg13g2_dfrbp_1 \ppu.pal[11][3]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net552),
    .D(_00318_),
    .Q_N(_08861_),
    .Q(\ppu.pal[11][3] ));
 sg13g2_dfrbp_1 \ppu.pal[11][4]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net553),
    .D(_00319_),
    .Q_N(_08860_),
    .Q(\ppu.pal[11][4] ));
 sg13g2_dfrbp_1 \ppu.pal[11][5]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net554),
    .D(_00320_),
    .Q_N(_08859_),
    .Q(\ppu.pal[11][5] ));
 sg13g2_dfrbp_1 \ppu.pal[11][6]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net555),
    .D(_00321_),
    .Q_N(_08858_),
    .Q(\ppu.pal[11][6] ));
 sg13g2_dfrbp_1 \ppu.pal[11][7]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net556),
    .D(_00322_),
    .Q_N(_08857_),
    .Q(\ppu.pal[11][7] ));
 sg13g2_dfrbp_1 \ppu.pal[12][0]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net557),
    .D(_00323_),
    .Q_N(_08856_),
    .Q(\ppu.pal[12][0] ));
 sg13g2_dfrbp_1 \ppu.pal[12][1]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net558),
    .D(_00324_),
    .Q_N(_08855_),
    .Q(\ppu.pal[12][1] ));
 sg13g2_dfrbp_1 \ppu.pal[12][2]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net559),
    .D(_00325_),
    .Q_N(_08854_),
    .Q(\ppu.pal[12][2] ));
 sg13g2_dfrbp_1 \ppu.pal[12][3]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net560),
    .D(_00326_),
    .Q_N(_08853_),
    .Q(\ppu.pal[12][3] ));
 sg13g2_dfrbp_1 \ppu.pal[12][4]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net561),
    .D(_00327_),
    .Q_N(_08852_),
    .Q(\ppu.pal[12][4] ));
 sg13g2_dfrbp_1 \ppu.pal[12][5]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net562),
    .D(_00328_),
    .Q_N(_08851_),
    .Q(\ppu.pal[12][5] ));
 sg13g2_dfrbp_1 \ppu.pal[12][6]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net563),
    .D(_00329_),
    .Q_N(_08850_),
    .Q(\ppu.pal[12][6] ));
 sg13g2_dfrbp_1 \ppu.pal[12][7]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net564),
    .D(_00330_),
    .Q_N(_08849_),
    .Q(\ppu.pal[12][7] ));
 sg13g2_dfrbp_1 \ppu.pal[13][0]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net565),
    .D(_00331_),
    .Q_N(_08848_),
    .Q(\ppu.pal[13][0] ));
 sg13g2_dfrbp_1 \ppu.pal[13][1]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net566),
    .D(_00332_),
    .Q_N(_08847_),
    .Q(\ppu.pal[13][1] ));
 sg13g2_dfrbp_1 \ppu.pal[13][2]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net567),
    .D(_00333_),
    .Q_N(_08846_),
    .Q(\ppu.pal[13][2] ));
 sg13g2_dfrbp_1 \ppu.pal[13][3]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net568),
    .D(_00334_),
    .Q_N(_08845_),
    .Q(\ppu.pal[13][3] ));
 sg13g2_dfrbp_1 \ppu.pal[13][4]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net569),
    .D(_00335_),
    .Q_N(_08844_),
    .Q(\ppu.pal[13][4] ));
 sg13g2_dfrbp_1 \ppu.pal[13][5]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net570),
    .D(_00336_),
    .Q_N(_08843_),
    .Q(\ppu.pal[13][5] ));
 sg13g2_dfrbp_1 \ppu.pal[13][6]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net571),
    .D(_00337_),
    .Q_N(_08842_),
    .Q(\ppu.pal[13][6] ));
 sg13g2_dfrbp_1 \ppu.pal[13][7]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net572),
    .D(_00338_),
    .Q_N(_08841_),
    .Q(\ppu.pal[13][7] ));
 sg13g2_dfrbp_1 \ppu.pal[14][0]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net573),
    .D(_00339_),
    .Q_N(_08840_),
    .Q(\ppu.pal[14][0] ));
 sg13g2_dfrbp_1 \ppu.pal[14][1]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net574),
    .D(_00340_),
    .Q_N(_08839_),
    .Q(\ppu.pal[14][1] ));
 sg13g2_dfrbp_1 \ppu.pal[14][2]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net575),
    .D(_00341_),
    .Q_N(_08838_),
    .Q(\ppu.pal[14][2] ));
 sg13g2_dfrbp_1 \ppu.pal[14][3]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net576),
    .D(_00342_),
    .Q_N(_08837_),
    .Q(\ppu.pal[14][3] ));
 sg13g2_dfrbp_1 \ppu.pal[14][4]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net577),
    .D(_00343_),
    .Q_N(_08836_),
    .Q(\ppu.pal[14][4] ));
 sg13g2_dfrbp_1 \ppu.pal[14][5]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net578),
    .D(_00344_),
    .Q_N(_08835_),
    .Q(\ppu.pal[14][5] ));
 sg13g2_dfrbp_1 \ppu.pal[14][6]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net579),
    .D(_00345_),
    .Q_N(_08834_),
    .Q(\ppu.pal[14][6] ));
 sg13g2_dfrbp_1 \ppu.pal[14][7]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net580),
    .D(_00346_),
    .Q_N(_08833_),
    .Q(\ppu.pal[14][7] ));
 sg13g2_dfrbp_1 \ppu.pal[15][0]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net581),
    .D(_00347_),
    .Q_N(_08832_),
    .Q(\ppu.pal[15][0] ));
 sg13g2_dfrbp_1 \ppu.pal[15][1]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net582),
    .D(_00348_),
    .Q_N(_08831_),
    .Q(\ppu.pal[15][1] ));
 sg13g2_dfrbp_1 \ppu.pal[15][2]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net583),
    .D(_00349_),
    .Q_N(_08830_),
    .Q(\ppu.pal[15][2] ));
 sg13g2_dfrbp_1 \ppu.pal[15][3]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net584),
    .D(_00350_),
    .Q_N(_08829_),
    .Q(\ppu.pal[15][3] ));
 sg13g2_dfrbp_1 \ppu.pal[15][4]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net585),
    .D(_00351_),
    .Q_N(_08828_),
    .Q(\ppu.pal[15][4] ));
 sg13g2_dfrbp_1 \ppu.pal[15][5]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net586),
    .D(_00352_),
    .Q_N(_08827_),
    .Q(\ppu.pal[15][5] ));
 sg13g2_dfrbp_1 \ppu.pal[15][6]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net587),
    .D(_00353_),
    .Q_N(_08826_),
    .Q(\ppu.pal[15][6] ));
 sg13g2_dfrbp_1 \ppu.pal[15][7]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net588),
    .D(_00354_),
    .Q_N(_08825_),
    .Q(\ppu.pal[15][7] ));
 sg13g2_dfrbp_1 \ppu.pal[1][0]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net589),
    .D(_00355_),
    .Q_N(_08824_),
    .Q(\ppu.pal[1][0] ));
 sg13g2_dfrbp_1 \ppu.pal[1][1]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net590),
    .D(_00356_),
    .Q_N(_08823_),
    .Q(\ppu.pal[1][1] ));
 sg13g2_dfrbp_1 \ppu.pal[1][2]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net591),
    .D(_00357_),
    .Q_N(_08822_),
    .Q(\ppu.pal[1][2] ));
 sg13g2_dfrbp_1 \ppu.pal[1][3]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net592),
    .D(_00358_),
    .Q_N(_08821_),
    .Q(\ppu.pal[1][3] ));
 sg13g2_dfrbp_1 \ppu.pal[1][4]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net593),
    .D(_00359_),
    .Q_N(_08820_),
    .Q(\ppu.pal[1][4] ));
 sg13g2_dfrbp_1 \ppu.pal[1][5]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net594),
    .D(_00360_),
    .Q_N(_08819_),
    .Q(\ppu.pal[1][5] ));
 sg13g2_dfrbp_1 \ppu.pal[1][6]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net595),
    .D(_00361_),
    .Q_N(_08818_),
    .Q(\ppu.pal[1][6] ));
 sg13g2_dfrbp_1 \ppu.pal[1][7]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net596),
    .D(_00362_),
    .Q_N(_08817_),
    .Q(\ppu.pal[1][7] ));
 sg13g2_dfrbp_1 \ppu.pal[2][0]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net597),
    .D(_00363_),
    .Q_N(_08816_),
    .Q(\ppu.pal[2][0] ));
 sg13g2_dfrbp_1 \ppu.pal[2][1]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net598),
    .D(_00364_),
    .Q_N(_08815_),
    .Q(\ppu.pal[2][1] ));
 sg13g2_dfrbp_1 \ppu.pal[2][2]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net599),
    .D(_00365_),
    .Q_N(_08814_),
    .Q(\ppu.pal[2][2] ));
 sg13g2_dfrbp_1 \ppu.pal[2][3]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net600),
    .D(_00366_),
    .Q_N(_08813_),
    .Q(\ppu.pal[2][3] ));
 sg13g2_dfrbp_1 \ppu.pal[2][4]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net601),
    .D(_00367_),
    .Q_N(_08812_),
    .Q(\ppu.pal[2][4] ));
 sg13g2_dfrbp_1 \ppu.pal[2][5]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net602),
    .D(_00368_),
    .Q_N(_08811_),
    .Q(\ppu.pal[2][5] ));
 sg13g2_dfrbp_1 \ppu.pal[2][6]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net603),
    .D(_00369_),
    .Q_N(_08810_),
    .Q(\ppu.pal[2][6] ));
 sg13g2_dfrbp_1 \ppu.pal[2][7]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net604),
    .D(_00370_),
    .Q_N(_08809_),
    .Q(\ppu.pal[2][7] ));
 sg13g2_dfrbp_1 \ppu.pal[3][0]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net605),
    .D(_00371_),
    .Q_N(_08808_),
    .Q(\ppu.pal[3][0] ));
 sg13g2_dfrbp_1 \ppu.pal[3][1]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net606),
    .D(_00372_),
    .Q_N(_08807_),
    .Q(\ppu.pal[3][1] ));
 sg13g2_dfrbp_1 \ppu.pal[3][2]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net607),
    .D(_00373_),
    .Q_N(_08806_),
    .Q(\ppu.pal[3][2] ));
 sg13g2_dfrbp_1 \ppu.pal[3][3]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net608),
    .D(_00374_),
    .Q_N(_08805_),
    .Q(\ppu.pal[3][3] ));
 sg13g2_dfrbp_1 \ppu.pal[3][4]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net609),
    .D(_00375_),
    .Q_N(_08804_),
    .Q(\ppu.pal[3][4] ));
 sg13g2_dfrbp_1 \ppu.pal[3][5]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net610),
    .D(_00376_),
    .Q_N(_08803_),
    .Q(\ppu.pal[3][5] ));
 sg13g2_dfrbp_1 \ppu.pal[3][6]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net611),
    .D(_00377_),
    .Q_N(_08802_),
    .Q(\ppu.pal[3][6] ));
 sg13g2_dfrbp_1 \ppu.pal[3][7]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net612),
    .D(_00378_),
    .Q_N(_08801_),
    .Q(\ppu.pal[3][7] ));
 sg13g2_dfrbp_1 \ppu.pal[4][0]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net613),
    .D(_00379_),
    .Q_N(_08800_),
    .Q(\ppu.pal[4][0] ));
 sg13g2_dfrbp_1 \ppu.pal[4][1]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net614),
    .D(_00380_),
    .Q_N(_08799_),
    .Q(\ppu.pal[4][1] ));
 sg13g2_dfrbp_1 \ppu.pal[4][2]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net615),
    .D(_00381_),
    .Q_N(_08798_),
    .Q(\ppu.pal[4][2] ));
 sg13g2_dfrbp_1 \ppu.pal[4][3]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net616),
    .D(_00382_),
    .Q_N(_08797_),
    .Q(\ppu.pal[4][3] ));
 sg13g2_dfrbp_1 \ppu.pal[4][4]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net617),
    .D(_00383_),
    .Q_N(_08796_),
    .Q(\ppu.pal[4][4] ));
 sg13g2_dfrbp_1 \ppu.pal[4][5]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net618),
    .D(_00384_),
    .Q_N(_08795_),
    .Q(\ppu.pal[4][5] ));
 sg13g2_dfrbp_1 \ppu.pal[4][6]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net619),
    .D(_00385_),
    .Q_N(_08794_),
    .Q(\ppu.pal[4][6] ));
 sg13g2_dfrbp_1 \ppu.pal[4][7]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net620),
    .D(_00386_),
    .Q_N(_08793_),
    .Q(\ppu.pal[4][7] ));
 sg13g2_dfrbp_1 \ppu.pal[5][0]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net621),
    .D(_00387_),
    .Q_N(_08792_),
    .Q(\ppu.pal[5][0] ));
 sg13g2_dfrbp_1 \ppu.pal[5][1]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net622),
    .D(_00388_),
    .Q_N(_08791_),
    .Q(\ppu.pal[5][1] ));
 sg13g2_dfrbp_1 \ppu.pal[5][2]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net623),
    .D(_00389_),
    .Q_N(_08790_),
    .Q(\ppu.pal[5][2] ));
 sg13g2_dfrbp_1 \ppu.pal[5][3]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net624),
    .D(_00390_),
    .Q_N(_08789_),
    .Q(\ppu.pal[5][3] ));
 sg13g2_dfrbp_1 \ppu.pal[5][4]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net625),
    .D(_00391_),
    .Q_N(_08788_),
    .Q(\ppu.pal[5][4] ));
 sg13g2_dfrbp_1 \ppu.pal[5][5]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net626),
    .D(_00392_),
    .Q_N(_08787_),
    .Q(\ppu.pal[5][5] ));
 sg13g2_dfrbp_1 \ppu.pal[5][6]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net627),
    .D(_00393_),
    .Q_N(_08786_),
    .Q(\ppu.pal[5][6] ));
 sg13g2_dfrbp_1 \ppu.pal[5][7]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net628),
    .D(_00394_),
    .Q_N(_08785_),
    .Q(\ppu.pal[5][7] ));
 sg13g2_dfrbp_1 \ppu.pal[6][0]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net629),
    .D(_00395_),
    .Q_N(_08784_),
    .Q(\ppu.pal[6][0] ));
 sg13g2_dfrbp_1 \ppu.pal[6][1]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net630),
    .D(_00396_),
    .Q_N(_08783_),
    .Q(\ppu.pal[6][1] ));
 sg13g2_dfrbp_1 \ppu.pal[6][2]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net631),
    .D(_00397_),
    .Q_N(_08782_),
    .Q(\ppu.pal[6][2] ));
 sg13g2_dfrbp_1 \ppu.pal[6][3]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net632),
    .D(_00398_),
    .Q_N(_08781_),
    .Q(\ppu.pal[6][3] ));
 sg13g2_dfrbp_1 \ppu.pal[6][4]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net633),
    .D(_00399_),
    .Q_N(_08780_),
    .Q(\ppu.pal[6][4] ));
 sg13g2_dfrbp_1 \ppu.pal[6][5]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net634),
    .D(_00400_),
    .Q_N(_08779_),
    .Q(\ppu.pal[6][5] ));
 sg13g2_dfrbp_1 \ppu.pal[6][6]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net635),
    .D(_00401_),
    .Q_N(_08778_),
    .Q(\ppu.pal[6][6] ));
 sg13g2_dfrbp_1 \ppu.pal[6][7]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net636),
    .D(_00402_),
    .Q_N(_08777_),
    .Q(\ppu.pal[6][7] ));
 sg13g2_dfrbp_1 \ppu.pal[7][0]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net637),
    .D(_00403_),
    .Q_N(_08776_),
    .Q(\ppu.pal[7][0] ));
 sg13g2_dfrbp_1 \ppu.pal[7][1]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net638),
    .D(_00404_),
    .Q_N(_08775_),
    .Q(\ppu.pal[7][1] ));
 sg13g2_dfrbp_1 \ppu.pal[7][2]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net639),
    .D(_00405_),
    .Q_N(_08774_),
    .Q(\ppu.pal[7][2] ));
 sg13g2_dfrbp_1 \ppu.pal[7][3]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net640),
    .D(_00406_),
    .Q_N(_08773_),
    .Q(\ppu.pal[7][3] ));
 sg13g2_dfrbp_1 \ppu.pal[7][4]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net641),
    .D(_00407_),
    .Q_N(_08772_),
    .Q(\ppu.pal[7][4] ));
 sg13g2_dfrbp_1 \ppu.pal[7][5]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net642),
    .D(_00408_),
    .Q_N(_08771_),
    .Q(\ppu.pal[7][5] ));
 sg13g2_dfrbp_1 \ppu.pal[7][6]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net643),
    .D(_00409_),
    .Q_N(_08770_),
    .Q(\ppu.pal[7][6] ));
 sg13g2_dfrbp_1 \ppu.pal[7][7]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net644),
    .D(_00410_),
    .Q_N(_08769_),
    .Q(\ppu.pal[7][7] ));
 sg13g2_dfrbp_1 \ppu.pal[8][0]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net645),
    .D(_00411_),
    .Q_N(_08768_),
    .Q(\ppu.pal[8][0] ));
 sg13g2_dfrbp_1 \ppu.pal[8][1]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net646),
    .D(_00412_),
    .Q_N(_08767_),
    .Q(\ppu.pal[8][1] ));
 sg13g2_dfrbp_1 \ppu.pal[8][2]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net647),
    .D(_00413_),
    .Q_N(_08766_),
    .Q(\ppu.pal[8][2] ));
 sg13g2_dfrbp_1 \ppu.pal[8][3]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net648),
    .D(_00414_),
    .Q_N(_08765_),
    .Q(\ppu.pal[8][3] ));
 sg13g2_dfrbp_1 \ppu.pal[8][4]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net649),
    .D(_00415_),
    .Q_N(_08764_),
    .Q(\ppu.pal[8][4] ));
 sg13g2_dfrbp_1 \ppu.pal[8][5]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net650),
    .D(_00416_),
    .Q_N(_08763_),
    .Q(\ppu.pal[8][5] ));
 sg13g2_dfrbp_1 \ppu.pal[8][6]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net651),
    .D(_00417_),
    .Q_N(_08762_),
    .Q(\ppu.pal[8][6] ));
 sg13g2_dfrbp_1 \ppu.pal[8][7]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net652),
    .D(_00418_),
    .Q_N(_08761_),
    .Q(\ppu.pal[8][7] ));
 sg13g2_dfrbp_1 \ppu.pal[9][0]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net653),
    .D(_00419_),
    .Q_N(_08760_),
    .Q(\ppu.pal[9][0] ));
 sg13g2_dfrbp_1 \ppu.pal[9][1]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net654),
    .D(_00420_),
    .Q_N(_08759_),
    .Q(\ppu.pal[9][1] ));
 sg13g2_dfrbp_1 \ppu.pal[9][2]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net655),
    .D(_00421_),
    .Q_N(_08758_),
    .Q(\ppu.pal[9][2] ));
 sg13g2_dfrbp_1 \ppu.pal[9][3]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net656),
    .D(_00422_),
    .Q_N(_08757_),
    .Q(\ppu.pal[9][3] ));
 sg13g2_dfrbp_1 \ppu.pal[9][4]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net657),
    .D(_00423_),
    .Q_N(_08756_),
    .Q(\ppu.pal[9][4] ));
 sg13g2_dfrbp_1 \ppu.pal[9][5]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net658),
    .D(_00424_),
    .Q_N(_08755_),
    .Q(\ppu.pal[9][5] ));
 sg13g2_dfrbp_1 \ppu.pal[9][6]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net659),
    .D(_00425_),
    .Q_N(_08754_),
    .Q(\ppu.pal[9][6] ));
 sg13g2_dfrbp_1 \ppu.pal[9][7]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net660),
    .D(_00426_),
    .Q_N(_08994_),
    .Q(\ppu.pal[9][7] ));
 sg13g2_dfrbp_1 \ppu.pal_temp[4]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net661),
    .D(\ppu.pal_data_out[0] ),
    .Q_N(_08995_),
    .Q(\ppu.pal_out[0] ));
 sg13g2_dfrbp_1 \ppu.pal_temp[5]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net662),
    .D(\ppu.pal_data_out[1] ),
    .Q_N(_08996_),
    .Q(\ppu.pal_out[1] ));
 sg13g2_dfrbp_1 \ppu.pal_temp[6]$_DFF_P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net663),
    .D(\ppu.pal_data_out[2] ),
    .Q_N(_08997_),
    .Q(\ppu.pal_out[2] ));
 sg13g2_dfrbp_1 \ppu.pal_temp[7]$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net664),
    .D(\ppu.pal_data_out[3] ),
    .Q_N(_08753_),
    .Q(\ppu.pal_out[3] ));
 sg13g2_dfrbp_1 \ppu.ram_on$_SDFFE_PN0N_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net665),
    .D(_00427_),
    .Q_N(_08752_),
    .Q(\ppu.ram_on ));
 sg13g2_dfrbp_1 \ppu.ram_running$_SDFFE_PN0N_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net666),
    .D(_00428_),
    .Q_N(_00029_),
    .Q(\ppu.ram_running ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net667),
    .D(_00429_),
    .Q_N(_08751_),
    .Q(\ppu.copper_inst.dt_out[0] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[10]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net668),
    .D(_00430_),
    .Q_N(_08750_),
    .Q(\ppu.copper_inst.dt_sreg[10] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[11]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net669),
    .D(_00431_),
    .Q_N(_08749_),
    .Q(\ppu.copper_inst.dt_sreg[11] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[1]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net670),
    .D(_00432_),
    .Q_N(_08748_),
    .Q(\ppu.copper_inst.dt_out[1] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[2]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net671),
    .D(_00433_),
    .Q_N(_00031_),
    .Q(\ppu.copper_inst.dt_out[2] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net672),
    .D(_00434_),
    .Q_N(_08747_),
    .Q(\ppu.copper_inst.dt_sreg[3] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[4]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net673),
    .D(_00435_),
    .Q_N(_08746_),
    .Q(\ppu.copper_inst.dt_sreg[4] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[5]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net674),
    .D(_00436_),
    .Q_N(_00035_),
    .Q(\ppu.copper_inst.dt_sreg[5] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[6]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net675),
    .D(_00437_),
    .Q_N(_08745_),
    .Q(\ppu.copper_inst.dt_sreg[6] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[7]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net676),
    .D(_00438_),
    .Q_N(_08744_),
    .Q(\ppu.copper_inst.dt_sreg[7] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[8]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net677),
    .D(_00439_),
    .Q_N(_08743_),
    .Q(\ppu.copper_inst.dt_sreg[8] ));
 sg13g2_dfrbp_1 \ppu.rcoord.levels_sreg[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net678),
    .D(_00440_),
    .Q_N(_08742_),
    .Q(\ppu.copper_inst.dt_sreg[9] ));
 sg13g2_dfrbp_1 \ppu.rgb_out_reg[10]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net679),
    .D(_00441_),
    .Q_N(_00158_),
    .Q(\ppu.dither_r.u[1] ));
 sg13g2_dfrbp_1 \ppu.rgb_out_reg[11]$_DFFE_PN_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net680),
    .D(_00442_),
    .Q_N(_00157_),
    .Q(\ppu.dither_r.u[2] ));
 sg13g2_dfrbp_1 \ppu.rgb_out_reg[2]$_DFFE_PN_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net681),
    .D(_00443_),
    .Q_N(_00154_),
    .Q(\ppu.b0_out[2] ));
 sg13g2_dfrbp_1 \ppu.rgb_out_reg[3]$_DFFE_PN_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net682),
    .D(_00444_),
    .Q_N(_00153_),
    .Q(\ppu.b0_out[3] ));
 sg13g2_dfrbp_1 \ppu.rgb_out_reg[5]$_DFFE_PN_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net683),
    .D(_00445_),
    .Q_N(_08741_),
    .Q(\ppu.dither_g.u[0] ));
 sg13g2_dfrbp_1 \ppu.rgb_out_reg[6]$_DFFE_PN_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net684),
    .D(_00446_),
    .Q_N(_00156_),
    .Q(\ppu.dither_g.u[1] ));
 sg13g2_dfrbp_1 \ppu.rgb_out_reg[7]$_DFFE_PN_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net685),
    .D(_00447_),
    .Q_N(_00155_),
    .Q(\ppu.dither_g.u[2] ));
 sg13g2_dfrbp_1 \ppu.rgb_out_reg[9]$_DFFE_PN_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net686),
    .D(_00448_),
    .Q_N(_00152_),
    .Q(\ppu.b0_out[1] ));
 sg13g2_dfrbp_1 \ppu.rs2.vsync0$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net687),
    .D(_00449_),
    .Q_N(_08998_),
    .Q(\ppu.rs2.vsync0 ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.counter[0]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net688),
    .D(_00011_),
    .Q_N(_00032_),
    .Q(\ppu.copper_inst.x_cmp[0] ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.counter[1]$_DFF_P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net689),
    .D(_00012_),
    .Q_N(_00033_),
    .Q(\ppu.copper_inst.x_cmp[1] ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.counter[2]$_DFF_P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net690),
    .D(_00013_),
    .Q_N(_00034_),
    .Q(\ppu.copper_inst.x_cmp[2] ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.counter[3]$_SDFF_PN1_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net691),
    .D(_00450_),
    .Q_N(_00037_),
    .Q(\ppu.copper_inst.x_cmp[3] ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.counter[4]$_SDFF_PN1_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net692),
    .D(_00451_),
    .Q_N(_00038_),
    .Q(\ppu.copper_inst.x_cmp[4] ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.counter[5]$_SDFF_PP1_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net693),
    .D(_00452_),
    .Q_N(_00067_),
    .Q(\ppu.rs2.x0[5] ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.counter[6]$_SDFF_PP1_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net694),
    .D(_00453_),
    .Q_N(_00065_),
    .Q(\ppu.rs2.x0[6] ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.counter[7]$_SDFF_PP0_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net695),
    .D(_00454_),
    .Q_N(_00030_),
    .Q(\ppu.rs2.x0[7] ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.counter[8]$_SDFF_PP0_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net696),
    .D(_00455_),
    .Q_N(_00040_),
    .Q(\ppu.copper_inst.x_cmp[8] ));
 sg13g2_dfrbp_1 \ppu.rs2.x_scan.phase$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net697),
    .D(_00456_),
    .Q_N(_00180_),
    .Q(\ppu.rs2.phase_x ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.counter[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net698),
    .D(_00457_),
    .Q_N(_00036_),
    .Q(\ppu.rs2.y_scan.counter[0] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.counter[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net699),
    .D(_00458_),
    .Q_N(_00159_),
    .Q(\ppu.rs2.y_scan.counter[1] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.counter[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net700),
    .D(_00459_),
    .Q_N(_08740_),
    .Q(\ppu.rs2.y_scan.counter[2] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.counter[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net701),
    .D(_00460_),
    .Q_N(_08739_),
    .Q(\ppu.rs2.y_scan.counter[3] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.counter[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net702),
    .D(_00461_),
    .Q_N(_08738_),
    .Q(\ppu.rs2.y_scan.counter[4] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.counter[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net703),
    .D(_00462_),
    .Q_N(_08737_),
    .Q(\ppu.rs2.y_scan.counter[5] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.counter[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net704),
    .D(_00463_),
    .Q_N(_08736_),
    .Q(\ppu.rs2.y_scan.counter[6] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.counter[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net705),
    .D(_00464_),
    .Q_N(_08735_),
    .Q(\ppu.rs2.y_scan.counter[7] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.counter[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net706),
    .D(_00465_),
    .Q_N(_00043_),
    .Q(\ppu.rs2.y_scan.counter[8] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.phase[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net707),
    .D(_00466_),
    .Q_N(_00044_),
    .Q(\ppu.rs2.phase_y[0] ));
 sg13g2_dfrbp_1 \ppu.rs2.y_scan.phase[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net708),
    .D(_00467_),
    .Q_N(_08734_),
    .Q(\ppu.rs2.phase_y[1] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net709),
    .D(_00468_),
    .Q_N(_08733_),
    .Q(\ppu.scroll_regs[0][0] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net710),
    .D(_00469_),
    .Q_N(_08732_),
    .Q(\ppu.scroll_regs[0][1] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net711),
    .D(_00470_),
    .Q_N(_08731_),
    .Q(\ppu.scroll_regs[0][2] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net712),
    .D(_00471_),
    .Q_N(_08730_),
    .Q(\ppu.scroll_regs[0][3] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net713),
    .D(_00472_),
    .Q_N(_08729_),
    .Q(\ppu.scroll_regs[0][4] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net714),
    .D(_00473_),
    .Q_N(_08728_),
    .Q(\ppu.scroll_regs[0][5] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net715),
    .D(_00474_),
    .Q_N(_08727_),
    .Q(\ppu.scroll_regs[0][6] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net716),
    .D(_00475_),
    .Q_N(_08726_),
    .Q(\ppu.scroll_regs[0][7] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net717),
    .D(_00476_),
    .Q_N(_08725_),
    .Q(\ppu.scroll_regs[0][8] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net718),
    .D(_00477_),
    .Q_N(_08724_),
    .Q(\ppu.scroll_regs[1][0] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net719),
    .D(_00478_),
    .Q_N(_08723_),
    .Q(\ppu.scroll_regs[1][1] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net720),
    .D(_00479_),
    .Q_N(_08722_),
    .Q(\ppu.scroll_regs[1][2] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net721),
    .D(_00480_),
    .Q_N(_08721_),
    .Q(\ppu.scroll_regs[1][3] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net722),
    .D(_00481_),
    .Q_N(_08720_),
    .Q(\ppu.scroll_regs[1][4] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net723),
    .D(_00482_),
    .Q_N(_08719_),
    .Q(\ppu.scroll_regs[1][5] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net724),
    .D(_00483_),
    .Q_N(_08718_),
    .Q(\ppu.scroll_regs[1][6] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net725),
    .D(_00484_),
    .Q_N(_08717_),
    .Q(\ppu.scroll_regs[1][7] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net726),
    .D(_00485_),
    .Q_N(_08716_),
    .Q(\ppu.scroll_regs[1][8] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net727),
    .D(_00486_),
    .Q_N(_08715_),
    .Q(\ppu.scroll_regs[2][0] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net728),
    .D(_00487_),
    .Q_N(_08714_),
    .Q(\ppu.scroll_regs[2][1] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net729),
    .D(_00488_),
    .Q_N(_08713_),
    .Q(\ppu.scroll_regs[2][2] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net730),
    .D(_00489_),
    .Q_N(_08712_),
    .Q(\ppu.scroll_regs[2][3] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net731),
    .D(_00490_),
    .Q_N(_08711_),
    .Q(\ppu.scroll_regs[2][4] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net732),
    .D(_00491_),
    .Q_N(_08710_),
    .Q(\ppu.scroll_regs[2][5] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net733),
    .D(_00492_),
    .Q_N(_08709_),
    .Q(\ppu.scroll_regs[2][6] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net734),
    .D(_00493_),
    .Q_N(_08708_),
    .Q(\ppu.scroll_regs[2][7] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net735),
    .D(_00494_),
    .Q_N(_08707_),
    .Q(\ppu.scroll_regs[2][8] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net736),
    .D(_00495_),
    .Q_N(_08706_),
    .Q(\ppu.scroll_regs[3][0] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net737),
    .D(_00496_),
    .Q_N(_08705_),
    .Q(\ppu.scroll_regs[3][1] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net738),
    .D(_00497_),
    .Q_N(_08704_),
    .Q(\ppu.scroll_regs[3][2] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net739),
    .D(_00498_),
    .Q_N(_08703_),
    .Q(\ppu.scroll_regs[3][3] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net740),
    .D(_00499_),
    .Q_N(_08702_),
    .Q(\ppu.scroll_regs[3][4] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net741),
    .D(_00500_),
    .Q_N(_08701_),
    .Q(\ppu.scroll_regs[3][5] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net742),
    .D(_00501_),
    .Q_N(_08700_),
    .Q(\ppu.scroll_regs[3][6] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net743),
    .D(_00502_),
    .Q_N(_08699_),
    .Q(\ppu.scroll_regs[3][7] ));
 sg13g2_dfrbp_1 \ppu.scroll_regs[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net744),
    .D(_00503_),
    .Q_N(_08698_),
    .Q(\ppu.scroll_regs[3][8] ));
 sg13g2_dfrbp_1 \ppu.serial_counter[0]$_SDFF_PN0_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net745),
    .D(_00504_),
    .Q_N(_00179_),
    .Q(\ppu.copper_inst.serial_counter[0] ));
 sg13g2_dfrbp_1 \ppu.serial_counter[1]$_SDFF_PN0_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net746),
    .D(_00505_),
    .Q_N(_00122_),
    .Q(\ppu.copper_inst.serial_counter[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net747),
    .D(_00506_),
    .Q_N(_00072_),
    .Q(\ppu.sprite_buffer.attr_x[0][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net748),
    .D(_00507_),
    .Q_N(_08697_),
    .Q(\ppu.sprite_buffer.attr_x[0][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net749),
    .D(_00508_),
    .Q_N(_00123_),
    .Q(\ppu.sprite_buffer.attr_x[0][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net750),
    .D(_00509_),
    .Q_N(_08696_),
    .Q(\ppu.sprite_buffer.attr_x[0][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net751),
    .D(_00510_),
    .Q_N(_00073_),
    .Q(\ppu.sprite_buffer.attr_x[0][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net752),
    .D(_00511_),
    .Q_N(_00074_),
    .Q(\ppu.sprite_buffer.attr_x[0][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net753),
    .D(_00512_),
    .Q_N(_00075_),
    .Q(\ppu.sprite_buffer.attr_x[0][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net754),
    .D(_00513_),
    .Q_N(_00071_),
    .Q(\ppu.sprite_buffer.attr_x[0][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net755),
    .D(_00514_),
    .Q_N(_00070_),
    .Q(\ppu.sprite_buffer.attr_x[0][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net756),
    .D(_00515_),
    .Q_N(_00069_),
    .Q(\ppu.sprite_buffer.attr_x[0][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net757),
    .D(_00516_),
    .Q_N(_00068_),
    .Q(\ppu.sprite_buffer.attr_x[0][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net758),
    .D(_00517_),
    .Q_N(_00066_),
    .Q(\ppu.sprite_buffer.attr_x[0][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net759),
    .D(_00518_),
    .Q_N(_00064_),
    .Q(\ppu.sprite_buffer.attr_x[0][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net760),
    .D(_00519_),
    .Q_N(_00063_),
    .Q(\ppu.sprite_buffer.attr_x[0][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net761),
    .D(_00520_),
    .Q_N(_00062_),
    .Q(\ppu.sprite_buffer.attr_x[0][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net762),
    .D(_00521_),
    .Q_N(_08695_),
    .Q(\ppu.sprite_buffer.attr_x[0][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net763),
    .D(_00522_),
    .Q_N(_08694_),
    .Q(\ppu.sprite_buffer.attr_x[1][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net764),
    .D(_00523_),
    .Q_N(_08693_),
    .Q(\ppu.sprite_buffer.attr_x[1][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net765),
    .D(_00524_),
    .Q_N(_08692_),
    .Q(\ppu.sprite_buffer.attr_x[1][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net766),
    .D(_00525_),
    .Q_N(_08691_),
    .Q(\ppu.sprite_buffer.attr_x[1][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net767),
    .D(_00526_),
    .Q_N(_08690_),
    .Q(\ppu.sprite_buffer.attr_x[1][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net768),
    .D(_00527_),
    .Q_N(_08689_),
    .Q(\ppu.sprite_buffer.attr_x[1][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net769),
    .D(_00528_),
    .Q_N(_08688_),
    .Q(\ppu.sprite_buffer.attr_x[1][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net770),
    .D(_00529_),
    .Q_N(_08687_),
    .Q(\ppu.sprite_buffer.attr_x[1][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net771),
    .D(_00530_),
    .Q_N(_08686_),
    .Q(\ppu.sprite_buffer.attr_x[1][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net772),
    .D(_00531_),
    .Q_N(_08685_),
    .Q(\ppu.sprite_buffer.attr_x[1][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net773),
    .D(_00532_),
    .Q_N(_08684_),
    .Q(\ppu.sprite_buffer.attr_x[1][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net774),
    .D(_00533_),
    .Q_N(_08683_),
    .Q(\ppu.sprite_buffer.attr_x[1][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net775),
    .D(_00534_),
    .Q_N(_08682_),
    .Q(\ppu.sprite_buffer.attr_x[1][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net776),
    .D(_00535_),
    .Q_N(_08681_),
    .Q(\ppu.sprite_buffer.attr_x[1][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net777),
    .D(_00536_),
    .Q_N(_08680_),
    .Q(\ppu.sprite_buffer.attr_x[1][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net778),
    .D(_00537_),
    .Q_N(_08679_),
    .Q(\ppu.sprite_buffer.attr_x[1][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net779),
    .D(_00538_),
    .Q_N(_08678_),
    .Q(\ppu.sprite_buffer.attr_x[2][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net780),
    .D(_00539_),
    .Q_N(_08677_),
    .Q(\ppu.sprite_buffer.attr_x[2][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net781),
    .D(_00540_),
    .Q_N(_08676_),
    .Q(\ppu.sprite_buffer.attr_x[2][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net782),
    .D(_00541_),
    .Q_N(_08675_),
    .Q(\ppu.sprite_buffer.attr_x[2][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net783),
    .D(_00542_),
    .Q_N(_08674_),
    .Q(\ppu.sprite_buffer.attr_x[2][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net784),
    .D(_00543_),
    .Q_N(_08673_),
    .Q(\ppu.sprite_buffer.attr_x[2][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net785),
    .D(_00544_),
    .Q_N(_08672_),
    .Q(\ppu.sprite_buffer.attr_x[2][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net786),
    .D(_00545_),
    .Q_N(_08671_),
    .Q(\ppu.sprite_buffer.attr_x[2][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net787),
    .D(_00546_),
    .Q_N(_08670_),
    .Q(\ppu.sprite_buffer.attr_x[2][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net788),
    .D(_00547_),
    .Q_N(_08669_),
    .Q(\ppu.sprite_buffer.attr_x[2][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net789),
    .D(_00548_),
    .Q_N(_08668_),
    .Q(\ppu.sprite_buffer.attr_x[2][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net790),
    .D(_00549_),
    .Q_N(_08667_),
    .Q(\ppu.sprite_buffer.attr_x[2][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net791),
    .D(_00550_),
    .Q_N(_08666_),
    .Q(\ppu.sprite_buffer.attr_x[2][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net792),
    .D(_00551_),
    .Q_N(_08665_),
    .Q(\ppu.sprite_buffer.attr_x[2][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net793),
    .D(_00552_),
    .Q_N(_08664_),
    .Q(\ppu.sprite_buffer.attr_x[2][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net794),
    .D(_00553_),
    .Q_N(_08663_),
    .Q(\ppu.sprite_buffer.attr_x[2][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net795),
    .D(_00554_),
    .Q_N(_08662_),
    .Q(\ppu.sprite_buffer.attr_x[3][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net796),
    .D(_00555_),
    .Q_N(_08661_),
    .Q(\ppu.sprite_buffer.attr_x[3][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net797),
    .D(_00556_),
    .Q_N(_08660_),
    .Q(\ppu.sprite_buffer.attr_x[3][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net798),
    .D(_00557_),
    .Q_N(_08659_),
    .Q(\ppu.sprite_buffer.attr_x[3][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net799),
    .D(_00558_),
    .Q_N(_08658_),
    .Q(\ppu.sprite_buffer.attr_x[3][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net800),
    .D(_00559_),
    .Q_N(_08657_),
    .Q(\ppu.sprite_buffer.attr_x[3][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net801),
    .D(_00560_),
    .Q_N(_08656_),
    .Q(\ppu.sprite_buffer.attr_x[3][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net802),
    .D(_00561_),
    .Q_N(_08655_),
    .Q(\ppu.sprite_buffer.attr_x[3][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net803),
    .D(_00562_),
    .Q_N(_08654_),
    .Q(\ppu.sprite_buffer.attr_x[3][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net804),
    .D(_00563_),
    .Q_N(_08653_),
    .Q(\ppu.sprite_buffer.attr_x[3][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net805),
    .D(_00564_),
    .Q_N(_08652_),
    .Q(\ppu.sprite_buffer.attr_x[3][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net806),
    .D(_00565_),
    .Q_N(_08651_),
    .Q(\ppu.sprite_buffer.attr_x[3][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net807),
    .D(_00566_),
    .Q_N(_08650_),
    .Q(\ppu.sprite_buffer.attr_x[3][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net808),
    .D(_00567_),
    .Q_N(_08649_),
    .Q(\ppu.sprite_buffer.attr_x[3][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net809),
    .D(_00568_),
    .Q_N(_08648_),
    .Q(\ppu.sprite_buffer.attr_x[3][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_x[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net810),
    .D(_00569_),
    .Q_N(_08647_),
    .Q(\ppu.sprite_buffer.attr_x[3][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net811),
    .D(_00570_),
    .Q_N(_08646_),
    .Q(\ppu.sprite_buffer.attr_y[0][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net812),
    .D(_00571_),
    .Q_N(_08645_),
    .Q(\ppu.sprite_buffer.attr_y[0][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net813),
    .D(_00572_),
    .Q_N(_08644_),
    .Q(\ppu.sprite_buffer.attr_y[0][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net814),
    .D(_00573_),
    .Q_N(_08643_),
    .Q(\ppu.sprite_buffer.attr_y[0][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net815),
    .D(_00574_),
    .Q_N(_08642_),
    .Q(\ppu.sprite_buffer.attr_y[0][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net816),
    .D(_00575_),
    .Q_N(_08641_),
    .Q(\ppu.sprite_buffer.attr_y[0][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net817),
    .D(_00576_),
    .Q_N(_08640_),
    .Q(\ppu.sprite_buffer.attr_y[0][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net818),
    .D(_00577_),
    .Q_N(_08639_),
    .Q(\ppu.sprite_buffer.attr_y[0][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net819),
    .D(_00578_),
    .Q_N(_08638_),
    .Q(\ppu.sprite_buffer.attr_y[0][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net820),
    .D(_00579_),
    .Q_N(_08637_),
    .Q(\ppu.sprite_buffer.attr_y[0][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net821),
    .D(_00580_),
    .Q_N(_08636_),
    .Q(\ppu.sprite_buffer.attr_y[0][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net822),
    .D(_00581_),
    .Q_N(_08635_),
    .Q(\ppu.sprite_buffer.attr_y[0][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net823),
    .D(_00582_),
    .Q_N(_08634_),
    .Q(\ppu.sprite_buffer.attr_y[0][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net824),
    .D(_00583_),
    .Q_N(_08633_),
    .Q(\ppu.sprite_buffer.attr_y[0][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net825),
    .D(_00584_),
    .Q_N(_08632_),
    .Q(\ppu.sprite_buffer.attr_y[0][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net826),
    .D(_00585_),
    .Q_N(_08631_),
    .Q(\ppu.sprite_buffer.attr_y[1][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net827),
    .D(_00586_),
    .Q_N(_08630_),
    .Q(\ppu.sprite_buffer.attr_y[1][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net828),
    .D(_00587_),
    .Q_N(_08629_),
    .Q(\ppu.sprite_buffer.attr_y[1][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net829),
    .D(_00588_),
    .Q_N(_08628_),
    .Q(\ppu.sprite_buffer.attr_y[1][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net830),
    .D(_00589_),
    .Q_N(_08627_),
    .Q(\ppu.sprite_buffer.attr_y[1][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net831),
    .D(_00590_),
    .Q_N(_08626_),
    .Q(\ppu.sprite_buffer.attr_y[1][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net832),
    .D(_00591_),
    .Q_N(_08625_),
    .Q(\ppu.sprite_buffer.attr_y[1][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net833),
    .D(_00592_),
    .Q_N(_08624_),
    .Q(\ppu.sprite_buffer.attr_y[1][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net834),
    .D(_00593_),
    .Q_N(_08623_),
    .Q(\ppu.sprite_buffer.attr_y[1][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net835),
    .D(_00594_),
    .Q_N(_08622_),
    .Q(\ppu.sprite_buffer.attr_y[1][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net836),
    .D(_00595_),
    .Q_N(_08621_),
    .Q(\ppu.sprite_buffer.attr_y[1][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net837),
    .D(_00596_),
    .Q_N(_08620_),
    .Q(\ppu.sprite_buffer.attr_y[1][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net838),
    .D(_00597_),
    .Q_N(_08619_),
    .Q(\ppu.sprite_buffer.attr_y[1][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net839),
    .D(_00598_),
    .Q_N(_08618_),
    .Q(\ppu.sprite_buffer.attr_y[1][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.attr_y[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net840),
    .D(_00599_),
    .Q_N(_08617_),
    .Q(\ppu.sprite_buffer.attr_y[1][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.extra_sorted_addr_bits[0]$_SDFF_PP0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net841),
    .D(_00600_),
    .Q_N(_08616_),
    .Q(\ppu.sprite_buffer.extra_sorted_addr_bits[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.extra_sorted_addr_bits[1]$_SDFF_PP0_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net842),
    .D(_00601_),
    .Q_N(_08615_),
    .Q(\ppu.sprite_buffer.extra_sorted_addr_bits[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.extra_sorted_addr_bits[2]$_SDFF_PP0_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net843),
    .D(_00602_),
    .Q_N(_08614_),
    .Q(\ppu.sprite_buffer.extra_sorted_addr_bits[2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net844),
    .D(_00603_),
    .Q_N(_08613_),
    .Q(\ppu.sprite_buffer.id_buffer[0][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net845),
    .D(_00604_),
    .Q_N(_08612_),
    .Q(\ppu.sprite_buffer.id_buffer[0][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net846),
    .D(_00605_),
    .Q_N(_08611_),
    .Q(\ppu.sprite_buffer.id_buffer[0][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net847),
    .D(_00606_),
    .Q_N(_08610_),
    .Q(\ppu.sprite_buffer.id_buffer[0][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net848),
    .D(_00607_),
    .Q_N(_08609_),
    .Q(\ppu.sprite_buffer.id_buffer[0][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net849),
    .D(_00608_),
    .Q_N(_08608_),
    .Q(\ppu.sprite_buffer.id_buffer[0][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net850),
    .D(_00609_),
    .Q_N(_08607_),
    .Q(\ppu.sprite_buffer.id_buffer[1][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net851),
    .D(_00610_),
    .Q_N(_08606_),
    .Q(\ppu.sprite_buffer.id_buffer[1][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net852),
    .D(_00611_),
    .Q_N(_08605_),
    .Q(\ppu.sprite_buffer.id_buffer[1][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net853),
    .D(_00612_),
    .Q_N(_08604_),
    .Q(\ppu.sprite_buffer.id_buffer[1][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net854),
    .D(_00613_),
    .Q_N(_08603_),
    .Q(\ppu.sprite_buffer.id_buffer[1][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net855),
    .D(_00614_),
    .Q_N(_08602_),
    .Q(\ppu.sprite_buffer.id_buffer[1][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net856),
    .D(_00615_),
    .Q_N(_08601_),
    .Q(\ppu.sprite_buffer.id_buffer[2][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net857),
    .D(_00616_),
    .Q_N(_08600_),
    .Q(\ppu.sprite_buffer.id_buffer[2][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net858),
    .D(_00617_),
    .Q_N(_08599_),
    .Q(\ppu.sprite_buffer.id_buffer[2][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net859),
    .D(_00618_),
    .Q_N(_08598_),
    .Q(\ppu.sprite_buffer.id_buffer[2][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net860),
    .D(_00619_),
    .Q_N(_08597_),
    .Q(\ppu.sprite_buffer.id_buffer[2][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net861),
    .D(_00620_),
    .Q_N(_08596_),
    .Q(\ppu.sprite_buffer.id_buffer[2][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net862),
    .D(_00621_),
    .Q_N(_08595_),
    .Q(\ppu.sprite_buffer.id_buffer[3][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net863),
    .D(_00622_),
    .Q_N(_08594_),
    .Q(\ppu.sprite_buffer.id_buffer[3][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net864),
    .D(_00623_),
    .Q_N(_08593_),
    .Q(\ppu.sprite_buffer.id_buffer[3][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net865),
    .D(_00624_),
    .Q_N(_08592_),
    .Q(\ppu.sprite_buffer.id_buffer[3][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net866),
    .D(_00625_),
    .Q_N(_08591_),
    .Q(\ppu.sprite_buffer.id_buffer[3][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.id_buffer[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net867),
    .D(_00626_),
    .Q_N(_08590_),
    .Q(\ppu.sprite_buffer.id_buffer[3][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.in_counters[0][0]$_SDFF_PP0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net868),
    .D(_00627_),
    .Q_N(_08589_),
    .Q(\ppu.sprite_buffer.in_counter_idy[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.in_counters[0][1]$_SDFF_PP0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net869),
    .D(_00628_),
    .Q_N(_08588_),
    .Q(\ppu.sprite_buffer.in_counter_idy[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.in_counters[1][0]$_SDFF_PP0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net870),
    .D(_00629_),
    .Q_N(_00061_),
    .Q(\ppu.sprite_buffer.in_counters[1][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.in_counters[1][1]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net871),
    .D(_00630_),
    .Q_N(_08587_),
    .Q(\ppu.sprite_buffer.in_counters[1][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.in_counters[1][2]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net872),
    .D(_00631_),
    .Q_N(_08586_),
    .Q(\ppu.sprite_buffer.in_counters[1][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.in_counters[2][0]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net873),
    .D(_00632_),
    .Q_N(_08585_),
    .Q(\ppu.sprite_buffer.final_pixels_in ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.in_counters[2][1]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net874),
    .D(_00633_),
    .Q_N(_08584_),
    .Q(\ppu.sprite_buffer.in_counters[2][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.in_counters[2][2]$_SDFF_PP0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net875),
    .D(_00634_),
    .Q_N(_08999_),
    .Q(\ppu.sprite_buffer.in_counters[2][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.last_data_pins[0]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net876),
    .D(\data_pins[0] ),
    .Q_N(_09000_),
    .Q(\ppu.sprite_buffer.data8[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.last_data_pins[1]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net877),
    .D(\data_pins[1] ),
    .Q_N(_09001_),
    .Q(\ppu.sprite_buffer.data8[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.last_data_pins[2]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net878),
    .D(\data_pins[2] ),
    .Q_N(_09002_),
    .Q(\ppu.sprite_buffer.data8[2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.last_data_pins[3]$_DFF_P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net879),
    .D(\data_pins[3] ),
    .Q_N(_08583_),
    .Q(\ppu.sprite_buffer.data8[3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.oam_load_sprite_valid$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net880),
    .D(_00635_),
    .Q_N(_08582_),
    .Q(\ppu.sprite_buffer.oam_load_sprite_valid ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.oam_req_step$_SDFFE_PP0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net881),
    .D(_00636_),
    .Q_N(_00028_),
    .Q(\ppu.sprite_buffer.oam_req_step ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.out_counters[0][0]$_SDFF_PP0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net882),
    .D(_00637_),
    .Q_N(_00079_),
    .Q(\ppu.sprite_buffer.out_counters[0][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.out_counters[0][1]$_SDFF_PP0_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net883),
    .D(_00638_),
    .Q_N(_00078_),
    .Q(\ppu.sprite_buffer.out_counters[0][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.out_counters[0][2]$_SDFF_PP0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net884),
    .D(_00639_),
    .Q_N(_00178_),
    .Q(\ppu.sprite_buffer.out_counters[0][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.out_counters[1][0]$_SDFF_PP0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net885),
    .D(_00640_),
    .Q_N(_00151_),
    .Q(\ppu.sprite_buffer.out_counter_oam[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.out_counters[1][1]$_SDFF_PP0_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net886),
    .D(_00641_),
    .Q_N(_00077_),
    .Q(\ppu.sprite_buffer.out_counter_oam[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.out_counters[2][0]$_SDFF_PP0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net887),
    .D(_00642_),
    .Q_N(_00160_),
    .Q(\ppu.sprite_buffer.out_counters[2][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.out_counters[2][1]$_SDFF_PP0_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net888),
    .D(_00643_),
    .Q_N(_08581_),
    .Q(\ppu.sprite_buffer.out_counters[2][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.out_counters[2][2]$_SDFF_PP0_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net889),
    .D(_00644_),
    .Q_N(_08580_),
    .Q(\ppu.sprite_buffer.out_counters[2][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.scan_enabled$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net890),
    .D(_00645_),
    .Q_N(_09003_),
    .Q(\ppu.sprite_buffer.scan_enabled ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.scan_on$_DFF_P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net891),
    .D(_00015_),
    .Q_N(_09004_),
    .Q(\ppu.sprite_buffer.scan_on ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[0][0]$_DFF_P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net892),
    .D(_00016_),
    .Q_N(_00130_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[0][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[0][1]$_DFF_P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net893),
    .D(_00017_),
    .Q_N(_09005_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[0][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[0][2]$_DFF_P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net894),
    .D(_00018_),
    .Q_N(_09006_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[0][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[1][0]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net895),
    .D(_00019_),
    .Q_N(_00129_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[1][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[1][1]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net896),
    .D(_00020_),
    .Q_N(_09007_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[1][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[1][2]$_DFF_P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net897),
    .D(_00021_),
    .Q_N(_09008_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[1][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[2][0]$_DFF_P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net898),
    .D(_00022_),
    .Q_N(_00128_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[2][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[2][1]$_DFF_P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net899),
    .D(_00023_),
    .Q_N(_09009_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[2][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[2][2]$_DFF_P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net900),
    .D(_00024_),
    .Q_N(_09010_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[2][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[3][0]$_DFF_P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net901),
    .D(_00025_),
    .Q_N(_00127_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[3][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[3][1]$_DFF_P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net902),
    .D(_00026_),
    .Q_N(_09011_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[3][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_catch_up_counters[3][2]$_DFF_P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net903),
    .D(_00027_),
    .Q_N(_08579_),
    .Q(\ppu.sprite_buffer.sprite_catch_up_counters[3][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net904),
    .D(_00646_),
    .Q_N(_08578_),
    .Q(\ppu.sprite_buffer.sprite_ids[0][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net905),
    .D(_00647_),
    .Q_N(_08577_),
    .Q(\ppu.sprite_buffer.sprite_ids[0][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net906),
    .D(_00648_),
    .Q_N(_08576_),
    .Q(\ppu.sprite_buffer.sprite_ids[0][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net907),
    .D(_00649_),
    .Q_N(_08575_),
    .Q(\ppu.sprite_buffer.sprite_ids[0][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net908),
    .D(_00650_),
    .Q_N(_08574_),
    .Q(\ppu.sprite_buffer.sprite_ids[0][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net909),
    .D(_00651_),
    .Q_N(_08573_),
    .Q(\ppu.sprite_buffer.sprite_ids[0][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net910),
    .D(_00652_),
    .Q_N(_08572_),
    .Q(\ppu.sprite_buffer.sprite_ids[1][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net911),
    .D(_00653_),
    .Q_N(_08571_),
    .Q(\ppu.sprite_buffer.sprite_ids[1][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net912),
    .D(_00654_),
    .Q_N(_08570_),
    .Q(\ppu.sprite_buffer.sprite_ids[1][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net913),
    .D(_00655_),
    .Q_N(_08569_),
    .Q(\ppu.sprite_buffer.sprite_ids[1][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net914),
    .D(_00656_),
    .Q_N(_08568_),
    .Q(\ppu.sprite_buffer.sprite_ids[1][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net915),
    .D(_00657_),
    .Q_N(_08567_),
    .Q(\ppu.sprite_buffer.sprite_ids[1][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net916),
    .D(_00658_),
    .Q_N(_08566_),
    .Q(\ppu.sprite_buffer.sprite_ids[2][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net917),
    .D(_00659_),
    .Q_N(_08565_),
    .Q(\ppu.sprite_buffer.sprite_ids[2][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net918),
    .D(_00660_),
    .Q_N(_08564_),
    .Q(\ppu.sprite_buffer.sprite_ids[2][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net919),
    .D(_00661_),
    .Q_N(_08563_),
    .Q(\ppu.sprite_buffer.sprite_ids[2][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net920),
    .D(_00662_),
    .Q_N(_08562_),
    .Q(\ppu.sprite_buffer.sprite_ids[2][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net921),
    .D(_00663_),
    .Q_N(_08561_),
    .Q(\ppu.sprite_buffer.sprite_ids[2][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net922),
    .D(_00664_),
    .Q_N(_08560_),
    .Q(\ppu.sprite_buffer.sprite_ids[3][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net923),
    .D(_00665_),
    .Q_N(_08559_),
    .Q(\ppu.sprite_buffer.sprite_ids[3][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net924),
    .D(_00666_),
    .Q_N(_08558_),
    .Q(\ppu.sprite_buffer.sprite_ids[3][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net925),
    .D(_00667_),
    .Q_N(_08557_),
    .Q(\ppu.sprite_buffer.sprite_ids[3][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net926),
    .D(_00668_),
    .Q_N(_08556_),
    .Q(\ppu.sprite_buffer.sprite_ids[3][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_ids[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net927),
    .D(_00669_),
    .Q_N(_08555_),
    .Q(\ppu.sprite_buffer.sprite_ids[3][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_out_color[0]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net928),
    .D(_00670_),
    .Q_N(_08554_),
    .Q(\ppu.pixel_out_s[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_out_color[1]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net929),
    .D(_00671_),
    .Q_N(_08553_),
    .Q(\ppu.pixel_out_s[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_out_color[2]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net930),
    .D(_00672_),
    .Q_N(_08552_),
    .Q(\ppu.pixel_out_s[2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_out_color[3]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net931),
    .D(_00673_),
    .Q_N(_00041_),
    .Q(\ppu.pixel_out_s[3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_out_depth[0]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net932),
    .D(_00674_),
    .Q_N(_08551_),
    .Q(\ppu.depth_out_s[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_out_depth[1]$_DFFE_PP_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net933),
    .D(_00675_),
    .Q_N(_08550_),
    .Q(\ppu.depth_out_s[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net934),
    .D(_00676_),
    .Q_N(_08549_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net935),
    .D(_00677_),
    .Q_N(_08548_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net936),
    .D(_00678_),
    .Q_N(_08547_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net937),
    .D(_00679_),
    .Q_N(_08546_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net938),
    .D(_00680_),
    .Q_N(_08545_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net939),
    .D(_00681_),
    .Q_N(_08544_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net940),
    .D(_00682_),
    .Q_N(_08543_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net941),
    .D(_00683_),
    .Q_N(_08542_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][16] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net942),
    .D(_00684_),
    .Q_N(_08541_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][17] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net943),
    .D(_00685_),
    .Q_N(_08540_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][18] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net944),
    .D(_00686_),
    .Q_N(_08539_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][19] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net945),
    .D(_00687_),
    .Q_N(_00124_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net946),
    .D(_00688_),
    .Q_N(_08538_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][20] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net947),
    .D(_00689_),
    .Q_N(_08537_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][21] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net948),
    .D(_00690_),
    .Q_N(_08536_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][22] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net949),
    .D(_00691_),
    .Q_N(_08535_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][23] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net950),
    .D(_00692_),
    .Q_N(_08534_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][24] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net951),
    .D(_00693_),
    .Q_N(_08533_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][25] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net952),
    .D(_00694_),
    .Q_N(_08532_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][26] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net953),
    .D(_00695_),
    .Q_N(_08531_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][27] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net954),
    .D(_00696_),
    .Q_N(_08530_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][28] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net955),
    .D(_00697_),
    .Q_N(_08529_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][29] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net956),
    .D(_00698_),
    .Q_N(_08528_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net957),
    .D(_00699_),
    .Q_N(_08527_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][30] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net958),
    .D(_00700_),
    .Q_N(_08526_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][31] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net959),
    .D(_00701_),
    .Q_N(_00125_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net960),
    .D(_00702_),
    .Q_N(_08525_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net961),
    .D(_00703_),
    .Q_N(_08524_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net962),
    .D(_00704_),
    .Q_N(_08523_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net963),
    .D(_00705_),
    .Q_N(_08522_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net964),
    .D(_00706_),
    .Q_N(_08521_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net965),
    .D(_00707_),
    .Q_N(_08520_),
    .Q(\ppu.sprite_buffer.sprite_pixels[0][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net966),
    .D(_00708_),
    .Q_N(_08519_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net967),
    .D(_00709_),
    .Q_N(_08518_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net968),
    .D(_00710_),
    .Q_N(_08517_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net969),
    .D(_00711_),
    .Q_N(_08516_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net970),
    .D(_00712_),
    .Q_N(_08515_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net971),
    .D(_00713_),
    .Q_N(_08514_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net972),
    .D(_00714_),
    .Q_N(_08513_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net973),
    .D(_00715_),
    .Q_N(_08512_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][16] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net974),
    .D(_00716_),
    .Q_N(_08511_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][17] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net975),
    .D(_00717_),
    .Q_N(_08510_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][18] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net976),
    .D(_00718_),
    .Q_N(_08509_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][19] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net977),
    .D(_00719_),
    .Q_N(_08508_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net978),
    .D(_00720_),
    .Q_N(_08507_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][20] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net979),
    .D(_00721_),
    .Q_N(_08506_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][21] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net980),
    .D(_00722_),
    .Q_N(_08505_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][22] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net981),
    .D(_00723_),
    .Q_N(_08504_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][23] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net982),
    .D(_00724_),
    .Q_N(_08503_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][24] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net983),
    .D(_00725_),
    .Q_N(_08502_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][25] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net984),
    .D(_00726_),
    .Q_N(_08501_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][26] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net985),
    .D(_00727_),
    .Q_N(_08500_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][27] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net986),
    .D(_00728_),
    .Q_N(_08499_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][28] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net987),
    .D(_00729_),
    .Q_N(_08498_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][29] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net988),
    .D(_00730_),
    .Q_N(_08497_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net989),
    .D(_00731_),
    .Q_N(_08496_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][30] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net990),
    .D(_00732_),
    .Q_N(_08495_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][31] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net991),
    .D(_00733_),
    .Q_N(_08494_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net992),
    .D(_00734_),
    .Q_N(_08493_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net993),
    .D(_00735_),
    .Q_N(_08492_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net994),
    .D(_00736_),
    .Q_N(_08491_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net995),
    .D(_00737_),
    .Q_N(_08490_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net996),
    .D(_00738_),
    .Q_N(_08489_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net997),
    .D(_00739_),
    .Q_N(_08488_),
    .Q(\ppu.sprite_buffer.sprite_pixels[1][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net998),
    .D(_00740_),
    .Q_N(_08487_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net999),
    .D(_00741_),
    .Q_N(_08486_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1000),
    .D(_00742_),
    .Q_N(_08485_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1001),
    .D(_00743_),
    .Q_N(_08484_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1002),
    .D(_00744_),
    .Q_N(_08483_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1003),
    .D(_00745_),
    .Q_N(_08482_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1004),
    .D(_00746_),
    .Q_N(_08481_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1005),
    .D(_00747_),
    .Q_N(_08480_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][16] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1006),
    .D(_00748_),
    .Q_N(_08479_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][17] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1007),
    .D(_00749_),
    .Q_N(_08478_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][18] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1008),
    .D(_00750_),
    .Q_N(_08477_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][19] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1009),
    .D(_00751_),
    .Q_N(_08476_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1010),
    .D(_00752_),
    .Q_N(_08475_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][20] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1011),
    .D(_00753_),
    .Q_N(_08474_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][21] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1012),
    .D(_00754_),
    .Q_N(_08473_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][22] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1013),
    .D(_00755_),
    .Q_N(_08472_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][23] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1014),
    .D(_00756_),
    .Q_N(_08471_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][24] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1015),
    .D(_00757_),
    .Q_N(_08470_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][25] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1016),
    .D(_00758_),
    .Q_N(_08469_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][26] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1017),
    .D(_00759_),
    .Q_N(_08468_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][27] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1018),
    .D(_00760_),
    .Q_N(_08467_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][28] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1019),
    .D(_00761_),
    .Q_N(_08466_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][29] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1020),
    .D(_00762_),
    .Q_N(_08465_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1021),
    .D(_00763_),
    .Q_N(_08464_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][30] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1022),
    .D(_00764_),
    .Q_N(_08463_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][31] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1023),
    .D(_00765_),
    .Q_N(_08462_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1024),
    .D(_00766_),
    .Q_N(_08461_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1025),
    .D(_00767_),
    .Q_N(_08460_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1026),
    .D(_00768_),
    .Q_N(_08459_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1027),
    .D(_00769_),
    .Q_N(_08458_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1028),
    .D(_00770_),
    .Q_N(_08457_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1029),
    .D(_00771_),
    .Q_N(_08456_),
    .Q(\ppu.sprite_buffer.sprite_pixels[2][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1030),
    .D(_00772_),
    .Q_N(_08455_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1031),
    .D(_00773_),
    .Q_N(_08454_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][10] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1032),
    .D(_00774_),
    .Q_N(_08453_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][11] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1033),
    .D(_00775_),
    .Q_N(_08452_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][12] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1034),
    .D(_00776_),
    .Q_N(_08451_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][13] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1035),
    .D(_00777_),
    .Q_N(_08450_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][14] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1036),
    .D(_00778_),
    .Q_N(_08449_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][15] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1037),
    .D(_00779_),
    .Q_N(_08448_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][16] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1038),
    .D(_00780_),
    .Q_N(_08447_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][17] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1039),
    .D(_00781_),
    .Q_N(_08446_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][18] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1040),
    .D(_00782_),
    .Q_N(_08445_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][19] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1041),
    .D(_00783_),
    .Q_N(_08444_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1042),
    .D(_00784_),
    .Q_N(_08443_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][20] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1043),
    .D(_00785_),
    .Q_N(_08442_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][21] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1044),
    .D(_00786_),
    .Q_N(_08441_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][22] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1045),
    .D(_00787_),
    .Q_N(_08440_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][23] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1046),
    .D(_00788_),
    .Q_N(_08439_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][24] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1047),
    .D(_00789_),
    .Q_N(_08438_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][25] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1048),
    .D(_00790_),
    .Q_N(_08437_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][26] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1049),
    .D(_00791_),
    .Q_N(_08436_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][27] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1050),
    .D(_00792_),
    .Q_N(_08435_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][28] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1051),
    .D(_00793_),
    .Q_N(_08434_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][29] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1052),
    .D(_00794_),
    .Q_N(_08433_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1053),
    .D(_00795_),
    .Q_N(_08432_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][30] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1054),
    .D(_00796_),
    .Q_N(_08431_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][31] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1055),
    .D(_00797_),
    .Q_N(_08430_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1056),
    .D(_00798_),
    .Q_N(_08429_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1057),
    .D(_00799_),
    .Q_N(_08428_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1058),
    .D(_00800_),
    .Q_N(_08427_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1059),
    .D(_00801_),
    .Q_N(_08426_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][7] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1060),
    .D(_00802_),
    .Q_N(_08425_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][8] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.sprite_pixels[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1061),
    .D(_00803_),
    .Q_N(_08424_),
    .Q(\ppu.sprite_buffer.sprite_pixels[3][9] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_color[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1062),
    .D(_00804_),
    .Q_N(_08423_),
    .Q(\ppu.sprite_buffer.top_color[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_color[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1063),
    .D(_00805_),
    .Q_N(_08422_),
    .Q(\ppu.sprite_buffer.top_color[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_color[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1064),
    .D(_00806_),
    .Q_N(_08421_),
    .Q(\ppu.sprite_buffer.top_color[2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_color[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1065),
    .D(_00807_),
    .Q_N(_08420_),
    .Q(\ppu.sprite_buffer.top_color[3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_depth[0]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1066),
    .D(_00808_),
    .Q_N(_08419_),
    .Q(\ppu.sprite_buffer.top_depth[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_depth[1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1067),
    .D(_00809_),
    .Q_N(_08418_),
    .Q(\ppu.sprite_buffer.top_depth[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_prio[0]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1068),
    .D(_00810_),
    .Q_N(_08417_),
    .Q(\ppu.sprite_buffer.top_prio[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_prio[1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1069),
    .D(_00811_),
    .Q_N(_08416_),
    .Q(\ppu.sprite_buffer.top_prio[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_prio[2]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1070),
    .D(_00812_),
    .Q_N(_08415_),
    .Q(\ppu.sprite_buffer.top_prio[2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_prio[3]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1071),
    .D(_00813_),
    .Q_N(_08414_),
    .Q(\ppu.sprite_buffer.top_prio[3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_prio[4]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1072),
    .D(_00814_),
    .Q_N(_08413_),
    .Q(\ppu.sprite_buffer.top_prio[4] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_prio[5]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1073),
    .D(_00815_),
    .Q_N(_08412_),
    .Q(\ppu.sprite_buffer.top_prio[5] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.top_prio[6]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1074),
    .D(_00816_),
    .Q_N(_00126_),
    .Q(\ppu.sprite_buffer.top_prio[6] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.valid_sprites[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1075),
    .D(_00817_),
    .Q_N(_08411_),
    .Q(\ppu.sprite_buffer.valid_sprites[0] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.valid_sprites[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1076),
    .D(_00818_),
    .Q_N(_08410_),
    .Q(\ppu.sprite_buffer.valid_sprites[1] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.valid_sprites[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1077),
    .D(_00819_),
    .Q_N(_08409_),
    .Q(\ppu.sprite_buffer.valid_sprites[2] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.valid_sprites[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1078),
    .D(_00820_),
    .Q_N(_08408_),
    .Q(\ppu.sprite_buffer.valid_sprites[3] ));
 sg13g2_dfrbp_1 \ppu.sprite_buffer.y_matched0$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1079),
    .D(_00821_),
    .Q_N(_08407_),
    .Q(\ppu.sprite_buffer.y_matched0 ));
 sg13g2_dfrbp_1 \ppu.sync_delay[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1080),
    .D(_00822_),
    .Q_N(_08406_),
    .Q(\ppu.sync_delay[0] ));
 sg13g2_dfrbp_1 \ppu.sync_delay[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1081),
    .D(_00823_),
    .Q_N(_08405_),
    .Q(\ppu.sync_delay[1] ));
 sg13g2_dfrbp_1 \ppu.sync_delay[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1082),
    .D(_00824_),
    .Q_N(_08404_),
    .Q(\ppu.sync_delay[2] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1083),
    .D(_00825_),
    .Q_N(_08403_),
    .Q(\ppu.tilemap.attr[0][0] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1084),
    .D(_00826_),
    .Q_N(_08402_),
    .Q(\ppu.tilemap.attr[0][1] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1085),
    .D(_00827_),
    .Q_N(_08401_),
    .Q(\ppu.tilemap.attr[0][2] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1086),
    .D(_00828_),
    .Q_N(_08400_),
    .Q(\ppu.tilemap.attr[0][3] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1087),
    .D(_00829_),
    .Q_N(_00161_),
    .Q(\ppu.tilemap.attr[0][4] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1088),
    .D(_00830_),
    .Q_N(_08399_),
    .Q(\ppu.tilemap.attr[1][0] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1089),
    .D(_00831_),
    .Q_N(_08398_),
    .Q(\ppu.tilemap.attr[1][1] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1090),
    .D(_00832_),
    .Q_N(_08397_),
    .Q(\ppu.tilemap.attr[1][2] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1091),
    .D(_00833_),
    .Q_N(_08396_),
    .Q(\ppu.tilemap.attr[1][3] ));
 sg13g2_dfrbp_1 \ppu.tilemap.attr[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1092),
    .D(_00834_),
    .Q_N(_00162_),
    .Q(\ppu.tilemap.attr[1][4] ));
 sg13g2_dfrbp_1 \ppu.tilemap.depth_out_reg[0]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1093),
    .D(_00835_),
    .Q_N(_08395_),
    .Q(\ppu.depth_out_t[0] ));
 sg13g2_dfrbp_1 \ppu.tilemap.depth_out_reg[1]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1094),
    .D(_00836_),
    .Q_N(_08394_),
    .Q(\ppu.depth_out_t[1] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1095),
    .D(_00837_),
    .Q_N(_08393_),
    .Q(\ppu.tilemap.map_pixels[0][0] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1096),
    .D(_00838_),
    .Q_N(_08392_),
    .Q(\ppu.tilemap.map_pixels[0][10] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1097),
    .D(_00839_),
    .Q_N(_08391_),
    .Q(\ppu.tilemap.map_pixels[0][11] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1098),
    .D(_00840_),
    .Q_N(_08390_),
    .Q(\ppu.tilemap.map_pixels[0][12] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1099),
    .D(_00841_),
    .Q_N(_08389_),
    .Q(\ppu.tilemap.map_pixels[0][13] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1100),
    .D(_00842_),
    .Q_N(_08388_),
    .Q(\ppu.tilemap.map_pixels[0][14] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1101),
    .D(_00843_),
    .Q_N(_08387_),
    .Q(\ppu.tilemap.map_pixels[0][15] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1102),
    .D(_00844_),
    .Q_N(_08386_),
    .Q(\ppu.tilemap.map_pixels[0][1] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1103),
    .D(_00845_),
    .Q_N(_08385_),
    .Q(\ppu.tilemap.map_pixels[0][2] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1104),
    .D(_00846_),
    .Q_N(_08384_),
    .Q(\ppu.tilemap.map_pixels[0][3] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1105),
    .D(_00847_),
    .Q_N(_08383_),
    .Q(\ppu.tilemap.map_pixels[0][4] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1106),
    .D(_00848_),
    .Q_N(_08382_),
    .Q(\ppu.tilemap.map_pixels[0][5] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1107),
    .D(_00849_),
    .Q_N(_08381_),
    .Q(\ppu.tilemap.map_pixels[0][6] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1108),
    .D(_00850_),
    .Q_N(_08380_),
    .Q(\ppu.tilemap.map_pixels[0][7] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1109),
    .D(_00851_),
    .Q_N(_08379_),
    .Q(\ppu.tilemap.map_pixels[0][8] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1110),
    .D(_00852_),
    .Q_N(_08378_),
    .Q(\ppu.tilemap.map_pixels[0][9] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1111),
    .D(_00853_),
    .Q_N(_08377_),
    .Q(\ppu.tilemap.map_pixels[1][0] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1112),
    .D(_00854_),
    .Q_N(_08376_),
    .Q(\ppu.tilemap.map_pixels[1][10] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1113),
    .D(_00855_),
    .Q_N(_08375_),
    .Q(\ppu.tilemap.map_pixels[1][11] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1114),
    .D(_00856_),
    .Q_N(_08374_),
    .Q(\ppu.tilemap.map_pixels[1][12] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1115),
    .D(_00857_),
    .Q_N(_08373_),
    .Q(\ppu.tilemap.map_pixels[1][13] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1116),
    .D(_00858_),
    .Q_N(_08372_),
    .Q(\ppu.tilemap.map_pixels[1][14] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1117),
    .D(_00859_),
    .Q_N(_08371_),
    .Q(\ppu.tilemap.map_pixels[1][15] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1118),
    .D(_00860_),
    .Q_N(_08370_),
    .Q(\ppu.tilemap.map_pixels[1][1] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1119),
    .D(_00861_),
    .Q_N(_08369_),
    .Q(\ppu.tilemap.map_pixels[1][2] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1120),
    .D(_00862_),
    .Q_N(_08368_),
    .Q(\ppu.tilemap.map_pixels[1][3] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1121),
    .D(_00863_),
    .Q_N(_08367_),
    .Q(\ppu.tilemap.map_pixels[1][4] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1122),
    .D(_00864_),
    .Q_N(_08366_),
    .Q(\ppu.tilemap.map_pixels[1][5] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1123),
    .D(_00865_),
    .Q_N(_08365_),
    .Q(\ppu.tilemap.map_pixels[1][6] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1124),
    .D(_00866_),
    .Q_N(_08364_),
    .Q(\ppu.tilemap.map_pixels[1][7] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1125),
    .D(_00867_),
    .Q_N(_08363_),
    .Q(\ppu.tilemap.map_pixels[1][8] ));
 sg13g2_dfrbp_1 \ppu.tilemap.map_pixels[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1126),
    .D(_00868_),
    .Q_N(_08362_),
    .Q(\ppu.tilemap.map_pixels[1][9] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1127),
    .D(_00869_),
    .Q_N(_08361_),
    .Q(\ppu.tilemap.next_attr[0][0] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1128),
    .D(_00870_),
    .Q_N(_08360_),
    .Q(\ppu.tilemap.next_attr[0][1] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1129),
    .D(_00871_),
    .Q_N(_08359_),
    .Q(\ppu.tilemap.next_attr[0][2] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1130),
    .D(_00872_),
    .Q_N(_08358_),
    .Q(\ppu.tilemap.next_attr[0][3] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1131),
    .D(_00873_),
    .Q_N(_08357_),
    .Q(\ppu.tilemap.next_attr[0][4] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1132),
    .D(_00874_),
    .Q_N(_08356_),
    .Q(\ppu.tilemap.next_attr[1][0] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1133),
    .D(_00875_),
    .Q_N(_08355_),
    .Q(\ppu.tilemap.next_attr[1][1] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1134),
    .D(_00876_),
    .Q_N(_08354_),
    .Q(\ppu.tilemap.next_attr[1][2] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1135),
    .D(_00877_),
    .Q_N(_08353_),
    .Q(\ppu.tilemap.next_attr[1][3] ));
 sg13g2_dfrbp_1 \ppu.tilemap.next_attr[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1136),
    .D(_00878_),
    .Q_N(_08352_),
    .Q(\ppu.tilemap.next_attr[1][4] ));
 sg13g2_dfrbp_1 \ppu.tilemap.temp_out[0]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1137),
    .D(_00879_),
    .Q_N(_08351_),
    .Q(\ppu.pixel_out_t[0] ));
 sg13g2_dfrbp_1 \ppu.tilemap.temp_out[1]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1138),
    .D(_00880_),
    .Q_N(_08350_),
    .Q(\ppu.pixel_out_t[1] ));
 sg13g2_dfrbp_1 \ppu.tilemap.temp_out[2]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1139),
    .D(_00881_),
    .Q_N(_08349_),
    .Q(\ppu.pixel_out_t[2] ));
 sg13g2_dfrbp_1 \ppu.tilemap.temp_out[3]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1140),
    .D(_00882_),
    .Q_N(_00042_),
    .Q(\ppu.pixel_out_t[3] ));
 sg13g2_dfrbp_1 \reset$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1141),
    .D(_00000_),
    .Q_N(_00080_),
    .Q(reset));
 sg13g2_dfrbp_1 \rx_in_reg[0]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1142),
    .D(_00001_),
    .Q_N(_09012_),
    .Q(\rx_in_reg[0] ));
 sg13g2_dfrbp_1 \rx_in_reg[1]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1143),
    .D(_00002_),
    .Q_N(_08348_),
    .Q(\rx_in_reg[1] ));
 sg13g2_dfrbp_1 \synth.controller.counter[0]$_SDFFE_PP1N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1144),
    .D(_00883_),
    .Q_N(_00150_),
    .Q(\synth.controller.counter[0] ));
 sg13g2_dfrbp_1 \synth.controller.counter[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1145),
    .D(_00884_),
    .Q_N(_00047_),
    .Q(\synth.controller.counter[1] ));
 sg13g2_dfrbp_1 \synth.controller.counter[2]$_SDFFE_PP1N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1146),
    .D(_00885_),
    .Q_N(_08347_),
    .Q(\synth.controller.counter[2] ));
 sg13g2_dfrbp_1 \synth.controller.counter[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1147),
    .D(_00886_),
    .Q_N(_08346_),
    .Q(\synth.controller.counter[3] ));
 sg13g2_dfrbp_1 \synth.controller.curr_voice[0]$_SDFFE_PP1N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1148),
    .D(_00887_),
    .Q_N(_00146_),
    .Q(\synth.controller.curr_voice[0] ));
 sg13g2_dfrbp_1 \synth.controller.curr_voice[1]$_SDFFE_PP1N_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1149),
    .D(_00888_),
    .Q_N(_08345_),
    .Q(\synth.controller.curr_voice[1] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1150),
    .D(_00889_),
    .Q_N(_00056_),
    .Q(\synth.controller.out_reg[0] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[10]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1151),
    .D(_00890_),
    .Q_N(_08344_),
    .Q(\synth.controller.out_reg[10] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[11]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1152),
    .D(_00891_),
    .Q_N(_08343_),
    .Q(\synth.controller.out_reg[11] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[12]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1153),
    .D(_00892_),
    .Q_N(_08342_),
    .Q(\synth.controller.out_reg[12] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[13]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1154),
    .D(_00893_),
    .Q_N(_08341_),
    .Q(\synth.controller.out_reg[13] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[14]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1155),
    .D(_00894_),
    .Q_N(_08340_),
    .Q(\synth.controller.out_reg[14] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[15]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1156),
    .D(_00895_),
    .Q_N(_08339_),
    .Q(\synth.controller.out_reg[15] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[1]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1157),
    .D(_00896_),
    .Q_N(_08338_),
    .Q(\synth.controller.out_reg[1] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[2]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1158),
    .D(_00897_),
    .Q_N(_08337_),
    .Q(\synth.controller.out_reg[2] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[3]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1159),
    .D(_00898_),
    .Q_N(_08336_),
    .Q(\synth.controller.out_reg[3] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[4]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1160),
    .D(_00899_),
    .Q_N(_08335_),
    .Q(\synth.controller.out_reg[4] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[5]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1161),
    .D(_00900_),
    .Q_N(_08334_),
    .Q(\synth.controller.out_reg[5] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[6]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1162),
    .D(_00901_),
    .Q_N(_08333_),
    .Q(\synth.controller.out_reg[6] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[7]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1163),
    .D(_00902_),
    .Q_N(_08332_),
    .Q(\synth.controller.out_reg[7] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1164),
    .D(_00903_),
    .Q_N(_08331_),
    .Q(\synth.controller.out_reg[8] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg[9]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1165),
    .D(_00904_),
    .Q_N(_08330_),
    .Q(\synth.controller.out_reg[9] ));
 sg13g2_dfrbp_1 \synth.controller.out_reg_valid$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1166),
    .D(_00905_),
    .Q_N(_08329_),
    .Q(\synth.controller.out_reg_valid ));
 sg13g2_dfrbp_1 \synth.controller.ppu_ctrl_reg[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1167),
    .D(_00906_),
    .Q_N(_08328_),
    .Q(\ppu_ctrl[0] ));
 sg13g2_dfrbp_1 \synth.controller.ppu_ctrl_reg[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1168),
    .D(_00907_),
    .Q_N(_08327_),
    .Q(\ppu_ctrl[2] ));
 sg13g2_dfrbp_1 \synth.controller.ppu_ctrl_reg[3]$_SDFFE_PP1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1169),
    .D(_00908_),
    .Q_N(_08326_),
    .Q(dither_out));
 sg13g2_dfrbp_1 \synth.controller.ppu_ctrl_reg[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1170),
    .D(_00909_),
    .Q_N(_08325_),
    .Q(\ppu_ctrl[4] ));
 sg13g2_dfrbp_1 \synth.controller.read_index_reg[0]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1171),
    .D(_00910_),
    .Q_N(_00057_),
    .Q(\synth.controller.read_index_reg[0] ));
 sg13g2_dfrbp_1 \synth.controller.read_index_reg[1]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1172),
    .D(_00911_),
    .Q_N(_08324_),
    .Q(\synth.controller.read_index_reg[1] ));
 sg13g2_dfrbp_1 \synth.controller.read_index_reg[2]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1173),
    .D(_00912_),
    .Q_N(_08323_),
    .Q(\synth.controller.read_index_reg[2] ));
 sg13g2_dfrbp_1 \synth.controller.read_index_reg[3]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1174),
    .D(_00913_),
    .Q_N(_08322_),
    .Q(\synth.controller.read_index_reg[3] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[0]$_DFFE_PN_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1175),
    .D(_00914_),
    .Q_N(_08321_),
    .Q(\synth.controller.reg_wdata[0] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[10]$_DFFE_PN_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1176),
    .D(_00915_),
    .Q_N(_00119_),
    .Q(\synth.controller.reg_waddr[2] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[11]$_DFFE_PN_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1177),
    .D(_00916_),
    .Q_N(_08320_),
    .Q(\synth.controller.reg_waddr[3] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[12]$_DFFE_PN_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1178),
    .D(_00917_),
    .Q_N(_08319_),
    .Q(\synth.controller.rx_buffer[12] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[13]$_DFFE_PN_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1179),
    .D(_00918_),
    .Q_N(_08318_),
    .Q(\synth.controller.rx_buffer[13] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[14]$_DFFE_PN_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1180),
    .D(_00919_),
    .Q_N(_08317_),
    .Q(\synth.controller.rx_buffer[14] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[15]$_DFFE_PN_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1181),
    .D(_00920_),
    .Q_N(_08316_),
    .Q(\synth.controller.rx_buffer[15] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[1]$_DFFE_PN_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1182),
    .D(_00921_),
    .Q_N(_08315_),
    .Q(\synth.controller.reg_wdata[1] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[2]$_DFFE_PN_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1183),
    .D(_00922_),
    .Q_N(_08314_),
    .Q(\synth.controller.reg_wdata[2] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[3]$_DFFE_PN_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1184),
    .D(_00923_),
    .Q_N(_08313_),
    .Q(\synth.controller.reg_wdata[3] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[4]$_DFFE_PN_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1185),
    .D(_00924_),
    .Q_N(_08312_),
    .Q(\synth.controller.reg_wdata[4] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[5]$_DFFE_PN_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1186),
    .D(_00925_),
    .Q_N(_00121_),
    .Q(\synth.controller.reg_wdata[5] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[6]$_DFFE_PN_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1187),
    .D(_00926_),
    .Q_N(_00118_),
    .Q(\synth.controller.reg_wdata[6] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[7]$_DFFE_PN_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1188),
    .D(_00927_),
    .Q_N(_08311_),
    .Q(\synth.controller.reg_wdata[7] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[8]$_DFFE_PN_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1189),
    .D(_00928_),
    .Q_N(_08310_),
    .Q(\synth.controller.reg_waddr[0] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer[9]$_DFFE_PN_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1190),
    .D(_00929_),
    .Q_N(_08309_),
    .Q(\synth.controller.reg_waddr[1] ));
 sg13g2_dfrbp_1 \synth.controller.rx_buffer_valid$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1191),
    .D(_00930_),
    .Q_N(_08308_),
    .Q(\synth.controller.rx_buffer_valid ));
 sg13g2_dfrbp_1 \synth.controller.rx_sbs[0]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1192),
    .D(_00931_),
    .Q_N(_08307_),
    .Q(\synth.controller.rx_sbs[0] ));
 sg13g2_dfrbp_1 \synth.controller.rx_sbs[1]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1193),
    .D(_00932_),
    .Q_N(_08306_),
    .Q(\synth.controller.rx_sbs[1] ));
 sg13g2_dfrbp_1 \synth.controller.sample_counter[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1194),
    .D(_00933_),
    .Q_N(_08305_),
    .Q(\synth.controller.sample_counter[0] ));
 sg13g2_dfrbp_1 \synth.controller.sample_counter[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1195),
    .D(_00934_),
    .Q_N(_08304_),
    .Q(\synth.controller.sample_counter[1] ));
 sg13g2_dfrbp_1 \synth.controller.sample_credits[0]$_SDFF_PP1_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1196),
    .D(_00935_),
    .Q_N(_08303_),
    .Q(\synth.controller.sample_credits[0] ));
 sg13g2_dfrbp_1 \synth.controller.sample_credits[1]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1197),
    .D(_00936_),
    .Q_N(_08302_),
    .Q(\synth.controller.sample_credits[1] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_credits[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1198),
    .D(_00937_),
    .Q_N(_08301_),
    .Q(\synth.controller.sbio_credits[0] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_credits[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1199),
    .D(_00938_),
    .Q_N(_08300_),
    .Q(\synth.controller.sbio_credits[1] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_credits[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1200),
    .D(_00939_),
    .Q_N(_08299_),
    .Q(\synth.controller.sbio_credits[2] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_rx.counter[0]$_SDFF_PP1_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1201),
    .D(_00940_),
    .Q_N(_00181_),
    .Q(\synth.controller.rx_counter[0] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_rx.counter[1]$_SDFF_PP1_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1202),
    .D(_00941_),
    .Q_N(_08298_),
    .Q(\synth.controller.rx_counter[1] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_rx.counter[2]$_SDFF_PP1_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1203),
    .D(_00942_),
    .Q_N(_08297_),
    .Q(\synth.controller.rx_counter[2] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_rx.counter[3]$_SDFF_PP1_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1204),
    .D(_00943_),
    .Q_N(_08296_),
    .Q(\synth.controller.rx_counter[3] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_tx.counter[0]$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1205),
    .D(_00944_),
    .Q_N(_00182_),
    .Q(\synth.controller.sbio_tx.counter[0] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_tx.counter[1]$_SDFF_PP1_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1206),
    .D(_00945_),
    .Q_N(_08295_),
    .Q(\synth.controller.sbio_tx.counter[1] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_tx.counter[2]$_SDFF_PP1_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1207),
    .D(_00946_),
    .Q_N(_08294_),
    .Q(\synth.controller.sbio_tx.counter[2] ));
 sg13g2_dfrbp_1 \synth.controller.sbio_tx.counter[3]$_SDFF_PP1_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1208),
    .D(_00947_),
    .Q_N(_08293_),
    .Q(\synth.controller.sbio_tx.counter[3] ));
 sg13g2_dfrbp_1 \synth.controller.scanning_out$_SDFFE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1209),
    .D(_00948_),
    .Q_N(_08292_),
    .Q(\synth.controller.scanning_out ));
 sg13g2_dfrbp_1 \synth.controller.step_sample_reg$_SDFFE_PP1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1210),
    .D(_00949_),
    .Q_N(_08291_),
    .Q(\synth.controller.step_sample ));
 sg13g2_dfrbp_1 \synth.controller.sweep_addr_index[0]$_SDFF_PP1_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1211),
    .D(_00950_),
    .Q_N(_00149_),
    .Q(\synth.controller.sweep_addr_index[0] ));
 sg13g2_dfrbp_1 \synth.controller.sweep_addr_index[1]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1212),
    .D(_00951_),
    .Q_N(_08290_),
    .Q(\synth.controller.sweep_addr_index[1] ));
 sg13g2_dfrbp_1 \synth.controller.sweep_addr_index[2]$_SDFF_PP1_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1213),
    .D(_00952_),
    .Q_N(_08289_),
    .Q(\synth.controller.sweep_addr_index[2] ));
 sg13g2_dfrbp_1 \synth.controller.sweep_data_index[0]$_SDFF_PP1_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1214),
    .D(_00953_),
    .Q_N(_00148_),
    .Q(\synth.controller.sweep_data_index[0] ));
 sg13g2_dfrbp_1 \synth.controller.sweep_data_index[1]$_SDFF_PP0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1215),
    .D(_00954_),
    .Q_N(_00120_),
    .Q(\synth.controller.sweep_data_index[1] ));
 sg13g2_dfrbp_1 \synth.controller.sweep_data_index[2]$_SDFF_PP1_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1216),
    .D(_00955_),
    .Q_N(_00051_),
    .Q(\synth.controller.sweep_data_index[2] ));
 sg13g2_dfrbp_1 \synth.controller.tx_outstanding[0]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1217),
    .D(_00956_),
    .Q_N(_08288_),
    .Q(\synth.controller.tx_outstanding[0] ));
 sg13g2_dfrbp_1 \synth.controller.tx_outstanding[1]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1218),
    .D(_00957_),
    .Q_N(_08287_),
    .Q(\synth.controller.tx_outstanding[1] ));
 sg13g2_dfrbp_1 \synth.controller.tx_outstanding[2]$_SDFF_PP0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1219),
    .D(_00958_),
    .Q_N(_08286_),
    .Q(\synth.controller.tx_outstanding[2] ));
 sg13g2_dfrbp_1 \synth.controller.tx_source[0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1220),
    .D(_00959_),
    .Q_N(_00055_),
    .Q(\synth.controller.tx_source[0] ));
 sg13g2_dfrbp_1 \synth.controller.tx_source[1]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1221),
    .D(_00960_),
    .Q_N(_08285_),
    .Q(\synth.controller.tx_source[1] ));
 sg13g2_dfrbp_1 \synth.controller.write_index_reg[0]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1222),
    .D(_00961_),
    .Q_N(_00111_),
    .Q(\synth.controller.write_index_reg[0] ));
 sg13g2_dfrbp_1 \synth.controller.write_index_reg[1]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1223),
    .D(_00962_),
    .Q_N(_08284_),
    .Q(\synth.controller.write_index_reg[1] ));
 sg13g2_dfrbp_1 \synth.controller.write_index_reg[2]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1224),
    .D(_00963_),
    .Q_N(_08283_),
    .Q(\synth.controller.write_index_reg[2] ));
 sg13g2_dfrbp_1 \synth.controller.write_index_reg[3]$_SDFFCE_PP0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1225),
    .D(_00964_),
    .Q_N(_09013_),
    .Q(\synth.controller.write_index_reg[3] ));
 sg13g2_dfrbp_1 \synth.voice.a_sel_reg[1]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1226),
    .D(_00003_),
    .Q_N(_09014_),
    .Q(\synth.voice.a_sel_reg[1] ));
 sg13g2_dfrbp_1 \synth.voice.a_sel_reg[2]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1227),
    .D(_00004_),
    .Q_N(_09015_),
    .Q(\synth.voice.a_sel_reg[2] ));
 sg13g2_dfrbp_1 \synth.voice.a_sel_reg[3]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1228),
    .D(_00005_),
    .Q_N(_08282_),
    .Q(\synth.voice.a_sel_reg[3] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1229),
    .D(_00965_),
    .Q_N(_08281_),
    .Q(\synth.voice.acc[0] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1230),
    .D(_00966_),
    .Q_N(_08280_),
    .Q(\synth.controller.out[6] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1231),
    .D(_00967_),
    .Q_N(_08279_),
    .Q(\synth.controller.out[7] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1232),
    .D(_00968_),
    .Q_N(_08278_),
    .Q(\synth.controller.out[8] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1233),
    .D(_00969_),
    .Q_N(_08277_),
    .Q(\synth.controller.out[9] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1234),
    .D(_00970_),
    .Q_N(_08276_),
    .Q(\synth.controller.out[10] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1235),
    .D(_00971_),
    .Q_N(_08275_),
    .Q(\synth.controller.out[11] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1236),
    .D(_00972_),
    .Q_N(_08274_),
    .Q(\synth.controller.out[12] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1237),
    .D(_00973_),
    .Q_N(_08273_),
    .Q(\synth.controller.out[13] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1238),
    .D(_00974_),
    .Q_N(_08272_),
    .Q(\synth.controller.out[14] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1239),
    .D(_00975_),
    .Q_N(_08271_),
    .Q(\synth.controller.out[15] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1240),
    .D(_00976_),
    .Q_N(_08270_),
    .Q(\synth.voice.acc[1] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1241),
    .D(_00977_),
    .Q_N(_08269_),
    .Q(\synth.voice.acc[2] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1242),
    .D(_00978_),
    .Q_N(_08268_),
    .Q(\synth.voice.acc[3] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1243),
    .D(_00979_),
    .Q_N(_08267_),
    .Q(\synth.controller.out[0] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1244),
    .D(_00980_),
    .Q_N(_08266_),
    .Q(\synth.controller.out[1] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1245),
    .D(_00981_),
    .Q_N(_08265_),
    .Q(\synth.controller.out[2] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1246),
    .D(_00982_),
    .Q_N(_08264_),
    .Q(\synth.controller.out[3] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1247),
    .D(_00983_),
    .Q_N(_08263_),
    .Q(\synth.controller.out[4] ));
 sg13g2_dfrbp_1 \synth.voice.accs[0][9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1248),
    .D(_00984_),
    .Q_N(_08262_),
    .Q(\synth.controller.out[5] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1249),
    .D(_00985_),
    .Q_N(_08261_),
    .Q(\synth.voice.accs[1][0] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1250),
    .D(_00986_),
    .Q_N(_08260_),
    .Q(\synth.voice.accs[1][10] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1251),
    .D(_00987_),
    .Q_N(_08259_),
    .Q(\synth.voice.accs[1][11] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1252),
    .D(_00988_),
    .Q_N(_08258_),
    .Q(\synth.voice.accs[1][12] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1253),
    .D(_00989_),
    .Q_N(_08257_),
    .Q(\synth.voice.accs[1][13] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1254),
    .D(_00990_),
    .Q_N(_08256_),
    .Q(\synth.voice.accs[1][14] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1255),
    .D(_00991_),
    .Q_N(_08255_),
    .Q(\synth.voice.accs[1][15] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1256),
    .D(_00992_),
    .Q_N(_08254_),
    .Q(\synth.voice.accs[1][16] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1257),
    .D(_00993_),
    .Q_N(_08253_),
    .Q(\synth.voice.accs[1][17] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1258),
    .D(_00994_),
    .Q_N(_08252_),
    .Q(\synth.voice.accs[1][18] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1259),
    .D(_00995_),
    .Q_N(_08251_),
    .Q(\synth.voice.accs[1][19] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1260),
    .D(_00996_),
    .Q_N(_08250_),
    .Q(\synth.voice.accs[1][1] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1261),
    .D(_00997_),
    .Q_N(_08249_),
    .Q(\synth.voice.accs[1][2] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1262),
    .D(_00998_),
    .Q_N(_08248_),
    .Q(\synth.voice.accs[1][3] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1263),
    .D(_00999_),
    .Q_N(_08247_),
    .Q(\synth.voice.accs[1][4] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1264),
    .D(_01000_),
    .Q_N(_08246_),
    .Q(\synth.voice.accs[1][5] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1265),
    .D(_01001_),
    .Q_N(_08245_),
    .Q(\synth.voice.accs[1][6] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1266),
    .D(_01002_),
    .Q_N(_08244_),
    .Q(\synth.voice.accs[1][7] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1267),
    .D(_01003_),
    .Q_N(_08243_),
    .Q(\synth.voice.accs[1][8] ));
 sg13g2_dfrbp_1 \synth.voice.accs[1][9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1268),
    .D(_01004_),
    .Q_N(_08242_),
    .Q(\synth.voice.accs[1][9] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1269),
    .D(_01005_),
    .Q_N(_08241_),
    .Q(\synth.voice.accs[2][0] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1270),
    .D(_01006_),
    .Q_N(_08240_),
    .Q(\synth.voice.accs[2][10] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1271),
    .D(_01007_),
    .Q_N(_08239_),
    .Q(\synth.voice.accs[2][11] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1272),
    .D(_01008_),
    .Q_N(_08238_),
    .Q(\synth.voice.accs[2][12] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1273),
    .D(_01009_),
    .Q_N(_08237_),
    .Q(\synth.voice.accs[2][13] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1274),
    .D(_01010_),
    .Q_N(_08236_),
    .Q(\synth.voice.accs[2][14] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1275),
    .D(_01011_),
    .Q_N(_08235_),
    .Q(\synth.voice.accs[2][15] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1276),
    .D(_01012_),
    .Q_N(_08234_),
    .Q(\synth.voice.accs[2][16] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1277),
    .D(_01013_),
    .Q_N(_08233_),
    .Q(\synth.voice.accs[2][17] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1278),
    .D(_01014_),
    .Q_N(_08232_),
    .Q(\synth.voice.accs[2][18] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1279),
    .D(_01015_),
    .Q_N(_08231_),
    .Q(\synth.voice.accs[2][19] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1280),
    .D(_01016_),
    .Q_N(_08230_),
    .Q(\synth.voice.accs[2][1] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1281),
    .D(_01017_),
    .Q_N(_08229_),
    .Q(\synth.voice.accs[2][2] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1282),
    .D(_01018_),
    .Q_N(_08228_),
    .Q(\synth.voice.accs[2][3] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1283),
    .D(_01019_),
    .Q_N(_08227_),
    .Q(\synth.voice.accs[2][4] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1284),
    .D(_01020_),
    .Q_N(_08226_),
    .Q(\synth.voice.accs[2][5] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1285),
    .D(_01021_),
    .Q_N(_08225_),
    .Q(\synth.voice.accs[2][6] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1286),
    .D(_01022_),
    .Q_N(_08224_),
    .Q(\synth.voice.accs[2][7] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1287),
    .D(_01023_),
    .Q_N(_08223_),
    .Q(\synth.voice.accs[2][8] ));
 sg13g2_dfrbp_1 \synth.voice.accs[2][9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1288),
    .D(_01024_),
    .Q_N(_08222_),
    .Q(\synth.voice.accs[2][9] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1289),
    .D(_01025_),
    .Q_N(_08221_),
    .Q(\synth.voice.accs[3][0] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1290),
    .D(_01026_),
    .Q_N(_08220_),
    .Q(\synth.voice.accs[3][10] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1291),
    .D(_01027_),
    .Q_N(_08219_),
    .Q(\synth.voice.accs[3][11] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1292),
    .D(_01028_),
    .Q_N(_08218_),
    .Q(\synth.voice.accs[3][12] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1293),
    .D(_01029_),
    .Q_N(_08217_),
    .Q(\synth.voice.accs[3][13] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1294),
    .D(_01030_),
    .Q_N(_08216_),
    .Q(\synth.voice.accs[3][14] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1295),
    .D(_01031_),
    .Q_N(_08215_),
    .Q(\synth.voice.accs[3][15] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1296),
    .D(_01032_),
    .Q_N(_08214_),
    .Q(\synth.voice.accs[3][16] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1297),
    .D(_01033_),
    .Q_N(_08213_),
    .Q(\synth.voice.accs[3][17] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1298),
    .D(_01034_),
    .Q_N(_08212_),
    .Q(\synth.voice.accs[3][18] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1299),
    .D(_01035_),
    .Q_N(_08211_),
    .Q(\synth.voice.accs[3][19] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1300),
    .D(_01036_),
    .Q_N(_08210_),
    .Q(\synth.voice.accs[3][1] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1301),
    .D(_01037_),
    .Q_N(_08209_),
    .Q(\synth.voice.accs[3][2] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1302),
    .D(_01038_),
    .Q_N(_08208_),
    .Q(\synth.voice.accs[3][3] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1303),
    .D(_01039_),
    .Q_N(_08207_),
    .Q(\synth.voice.accs[3][4] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1304),
    .D(_01040_),
    .Q_N(_08206_),
    .Q(\synth.voice.accs[3][5] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1305),
    .D(_01041_),
    .Q_N(_08205_),
    .Q(\synth.voice.accs[3][6] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1306),
    .D(_01042_),
    .Q_N(_08204_),
    .Q(\synth.voice.accs[3][7] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1307),
    .D(_01043_),
    .Q_N(_08203_),
    .Q(\synth.voice.accs[3][8] ));
 sg13g2_dfrbp_1 \synth.voice.accs[3][9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1308),
    .D(_01044_),
    .Q_N(_08202_),
    .Q(\synth.voice.accs[3][9] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1309),
    .D(_01045_),
    .Q_N(_08201_),
    .Q(\synth.voice.accs[4][0] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1310),
    .D(_01046_),
    .Q_N(_08200_),
    .Q(\synth.voice.accs[4][10] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1311),
    .D(_01047_),
    .Q_N(_08199_),
    .Q(\synth.voice.accs[4][11] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1312),
    .D(_01048_),
    .Q_N(_08198_),
    .Q(\synth.voice.accs[4][12] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1313),
    .D(_01049_),
    .Q_N(_08197_),
    .Q(\synth.voice.accs[4][13] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1314),
    .D(_01050_),
    .Q_N(_08196_),
    .Q(\synth.voice.accs[4][14] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1315),
    .D(_01051_),
    .Q_N(_08195_),
    .Q(\synth.voice.accs[4][15] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1316),
    .D(_01052_),
    .Q_N(_08194_),
    .Q(\synth.voice.accs[4][16] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1317),
    .D(_01053_),
    .Q_N(_08193_),
    .Q(\synth.voice.accs[4][17] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1318),
    .D(_01054_),
    .Q_N(_08192_),
    .Q(\synth.voice.accs[4][18] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1319),
    .D(_01055_),
    .Q_N(_08191_),
    .Q(\synth.voice.accs[4][19] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1320),
    .D(_01056_),
    .Q_N(_08190_),
    .Q(\synth.voice.accs[4][1] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1321),
    .D(_01057_),
    .Q_N(_08189_),
    .Q(\synth.voice.accs[4][2] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1322),
    .D(_01058_),
    .Q_N(_08188_),
    .Q(\synth.voice.accs[4][3] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1323),
    .D(_01059_),
    .Q_N(_08187_),
    .Q(\synth.voice.accs[4][4] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1324),
    .D(_01060_),
    .Q_N(_08186_),
    .Q(\synth.voice.accs[4][5] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1325),
    .D(_01061_),
    .Q_N(_08185_),
    .Q(\synth.voice.accs[4][6] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1326),
    .D(_01062_),
    .Q_N(_08184_),
    .Q(\synth.voice.accs[4][7] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1327),
    .D(_01063_),
    .Q_N(_08183_),
    .Q(\synth.voice.accs[4][8] ));
 sg13g2_dfrbp_1 \synth.voice.accs[4][9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1328),
    .D(_01064_),
    .Q_N(_08182_),
    .Q(\synth.voice.accs[4][9] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1329),
    .D(_01065_),
    .Q_N(_08181_),
    .Q(\synth.voice.accs[5][0] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1330),
    .D(_01066_),
    .Q_N(_08180_),
    .Q(\synth.voice.accs[5][10] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1331),
    .D(_01067_),
    .Q_N(_08179_),
    .Q(\synth.voice.accs[5][11] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1332),
    .D(_01068_),
    .Q_N(_08178_),
    .Q(\synth.voice.accs[5][12] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1333),
    .D(_01069_),
    .Q_N(_08177_),
    .Q(\synth.voice.accs[5][13] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][14]$_SDFFE_PP0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1334),
    .D(_01070_),
    .Q_N(_08176_),
    .Q(\synth.voice.accs[5][14] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][15]$_SDFFE_PP0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1335),
    .D(_01071_),
    .Q_N(_08175_),
    .Q(\synth.voice.accs[5][15] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][16]$_SDFFE_PP0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1336),
    .D(_01072_),
    .Q_N(_08174_),
    .Q(\synth.voice.accs[5][16] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][17]$_SDFFE_PP0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1337),
    .D(_01073_),
    .Q_N(_08173_),
    .Q(\synth.voice.accs[5][17] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][18]$_SDFFE_PP0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1338),
    .D(_01074_),
    .Q_N(_08172_),
    .Q(\synth.voice.accs[5][18] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][19]$_SDFFE_PP0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1339),
    .D(_01075_),
    .Q_N(_08171_),
    .Q(\synth.voice.accs[5][19] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1340),
    .D(_01076_),
    .Q_N(_08170_),
    .Q(\synth.voice.accs[5][1] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1341),
    .D(_01077_),
    .Q_N(_08169_),
    .Q(\synth.voice.accs[5][2] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1342),
    .D(_01078_),
    .Q_N(_08168_),
    .Q(\synth.voice.accs[5][3] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1343),
    .D(_01079_),
    .Q_N(_08167_),
    .Q(\synth.voice.accs[5][4] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1344),
    .D(_01080_),
    .Q_N(_08166_),
    .Q(\synth.voice.accs[5][5] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1345),
    .D(_01081_),
    .Q_N(_08165_),
    .Q(\synth.voice.accs[5][6] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1346),
    .D(_01082_),
    .Q_N(_08164_),
    .Q(\synth.voice.accs[5][7] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1347),
    .D(_01083_),
    .Q_N(_08163_),
    .Q(\synth.voice.accs[5][8] ));
 sg13g2_dfrbp_1 \synth.voice.accs[5][9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1348),
    .D(_01084_),
    .Q_N(_09016_),
    .Q(\synth.voice.accs[5][9] ));
 sg13g2_dfrbp_1 \synth.voice.b_sel_reg[0]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1349),
    .D(_00006_),
    .Q_N(_09017_),
    .Q(\synth.voice.b_sel_reg[0] ));
 sg13g2_dfrbp_1 \synth.voice.b_sel_reg[2]$_DFF_P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1350),
    .D(_00007_),
    .Q_N(_08162_),
    .Q(\synth.voice.b_sel_reg[2] ));
 sg13g2_dfrbp_1 \synth.voice.fir_offset_msbs[0]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1351),
    .D(_01085_),
    .Q_N(_00052_),
    .Q(\synth.voice.coeff_index[3] ));
 sg13g2_dfrbp_1 \synth.voice.fir_offset_msbs[1]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1352),
    .D(_01086_),
    .Q_N(_00050_),
    .Q(\synth.voice.coeff_index[4] ));
 sg13g2_dfrbp_1 \synth.voice.flip_sign_fir$_DFF_P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1353),
    .D(\synth.voice.fir_table.sign ),
    .Q_N(_09018_),
    .Q(\synth.voice.flip_sign_fir ));
 sg13g2_dfrbp_1 \synth.voice.flip_sign_reg$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1354),
    .D(\synth.voice.flip_sign ),
    .Q_N(_00145_),
    .Q(\synth.voice.flip_sign_reg ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1355),
    .D(_01087_),
    .Q_N(_00112_),
    .Q(\synth.voice.oct_counter[0] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1356),
    .D(_01088_),
    .Q_N(_08161_),
    .Q(\synth.voice.oct_counter[10] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1357),
    .D(_01089_),
    .Q_N(_00113_),
    .Q(\synth.voice.oct_counter[1] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1358),
    .D(_01090_),
    .Q_N(_00116_),
    .Q(\synth.voice.oct_counter[2] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1359),
    .D(_01091_),
    .Q_N(_00117_),
    .Q(\synth.voice.oct_counter[3] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1360),
    .D(_01092_),
    .Q_N(_08160_),
    .Q(\synth.voice.oct_counter[4] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1361),
    .D(_01093_),
    .Q_N(_08159_),
    .Q(\synth.voice.oct_counter[5] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1362),
    .D(_01094_),
    .Q_N(_08158_),
    .Q(\synth.voice.oct_counter[6] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1363),
    .D(_01095_),
    .Q_N(_08157_),
    .Q(\synth.voice.oct_counter[7] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1364),
    .D(_01096_),
    .Q_N(_08156_),
    .Q(\synth.voice.oct_counter[8] ));
 sg13g2_dfrbp_1 \synth.voice.oct_counter[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1365),
    .D(_01097_),
    .Q_N(_09019_),
    .Q(\synth.voice.oct_counter[9] ));
 sg13g2_dfrbp_1 \synth.voice.restart_acc_reg$_DFF_P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1366),
    .D(\synth.voice.restart_acc ),
    .Q_N(_09020_),
    .Q(\synth.controller.out_valid ));
 sg13g2_dfrbp_1 \synth.voice.rshift_reg0[0]$_DFF_P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1367),
    .D(\synth.voice.fir_table.exp[0] ),
    .Q_N(_00169_),
    .Q(\synth.voice.rshift_reg0[0] ));
 sg13g2_dfrbp_1 \synth.voice.rshift_reg0[1]$_DFF_P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1368),
    .D(\synth.voice.fir_table.exp[1] ),
    .Q_N(_00172_),
    .Q(\synth.voice.rshift_reg0[1] ));
 sg13g2_dfrbp_1 \synth.voice.rshift_reg0[2]$_DFF_P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1369),
    .D(\synth.voice.fir_table.exp[2] ),
    .Q_N(_00174_),
    .Q(\synth.voice.rshift_reg0[2] ));
 sg13g2_dfrbp_1 \synth.voice.rshift_reg0[3]$_DFF_P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1370),
    .D(\synth.voice.fir_table.exp[3] ),
    .Q_N(_00176_),
    .Q(\synth.voice.rshift_reg0[3] ));
 sg13g2_dfrbp_1 \synth.voice.rshift_reg[0]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1371),
    .D(\synth.voice.rshift[0] ),
    .Q_N(_09021_),
    .Q(\synth.voice.rshift_reg[0] ));
 sg13g2_dfrbp_1 \synth.voice.rshift_reg[1]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1372),
    .D(\synth.voice.rshift[1] ),
    .Q_N(_09022_),
    .Q(\synth.voice.rshift_reg[1] ));
 sg13g2_dfrbp_1 \synth.voice.rshift_reg[2]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1373),
    .D(\synth.voice.rshift[2] ),
    .Q_N(_09023_),
    .Q(\synth.voice.rshift_reg[2] ));
 sg13g2_dfrbp_1 \synth.voice.rshift_reg[3]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1374),
    .D(\synth.voice.rshift[3] ),
    .Q_N(_09024_),
    .Q(\synth.voice.rshift_reg[3] ));
 sg13g2_dfrbp_1 \synth.voice.scan_accs_reg$_DFF_P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1375),
    .D(\synth.voice.scan_accs ),
    .Q_N(_08155_),
    .Q(\synth.voice.scan_accs_reg ));
 sg13g2_dfrbp_1 \synth.voice.state[0]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1376),
    .D(_01098_),
    .Q_N(_00054_),
    .Q(\synth.voice.delayed_s ));
 sg13g2_dfrbp_1 \synth.voice.state[100]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1377),
    .D(_01099_),
    .Q_N(_08154_),
    .Q(\synth.voice.genblk4[6].next_state_scan[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[101]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1378),
    .D(_01100_),
    .Q_N(_00168_),
    .Q(\synth.voice.genblk4[6].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[102]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1379),
    .D(_01101_),
    .Q_N(_00167_),
    .Q(\synth.voice.genblk4[6].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[103]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1380),
    .D(_01102_),
    .Q_N(_00166_),
    .Q(\synth.voice.genblk4[6].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[104]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1381),
    .D(_01103_),
    .Q_N(_00165_),
    .Q(\synth.voice.genblk4[6].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[105]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1382),
    .D(_01104_),
    .Q_N(_00164_),
    .Q(\synth.voice.genblk4[6].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.state[106]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1383),
    .D(_01105_),
    .Q_N(_00170_),
    .Q(\synth.voice.genblk4[6].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[107]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1384),
    .D(_01106_),
    .Q_N(_00173_),
    .Q(\synth.voice.genblk4[6].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[108]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1385),
    .D(_01107_),
    .Q_N(_00175_),
    .Q(\synth.voice.genblk4[6].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[109]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1386),
    .D(_01108_),
    .Q_N(_00177_),
    .Q(\synth.voice.genblk4[6].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1387),
    .D(_01109_),
    .Q_N(_00100_),
    .Q(\synth.voice.genblk4[0].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[110]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1388),
    .D(_01110_),
    .Q_N(_08153_),
    .Q(\synth.voice.genblk4[6].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[111]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1389),
    .D(_01111_),
    .Q_N(_08152_),
    .Q(\synth.voice.genblk4[6].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[112]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1390),
    .D(_01112_),
    .Q_N(_08151_),
    .Q(\synth.voice.mods[1][2] ));
 sg13g2_dfrbp_1 \synth.voice.state[113]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1391),
    .D(_01113_),
    .Q_N(_08150_),
    .Q(\synth.voice.mods[1][3] ));
 sg13g2_dfrbp_1 \synth.voice.state[114]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1392),
    .D(_01114_),
    .Q_N(_08149_),
    .Q(\synth.voice.genblk4[7].next_state_scan[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[115]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1393),
    .D(_01115_),
    .Q_N(_08148_),
    .Q(\synth.voice.genblk4[7].next_state_scan[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[116]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1394),
    .D(_01116_),
    .Q_N(_08147_),
    .Q(\synth.voice.genblk4[7].next_state_scan[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[117]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1395),
    .D(_01117_),
    .Q_N(_08146_),
    .Q(\synth.voice.genblk4[7].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[118]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1396),
    .D(_01118_),
    .Q_N(_08145_),
    .Q(\synth.voice.genblk4[7].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[119]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1397),
    .D(_01119_),
    .Q_N(_08144_),
    .Q(\synth.voice.genblk4[7].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[11]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1398),
    .D(_01120_),
    .Q_N(_00098_),
    .Q(\synth.voice.genblk4[0].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[120]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1399),
    .D(_01121_),
    .Q_N(_08143_),
    .Q(\synth.voice.genblk4[7].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[121]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1400),
    .D(_01122_),
    .Q_N(_08142_),
    .Q(\synth.voice.genblk4[7].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.state[122]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1401),
    .D(_01123_),
    .Q_N(_08141_),
    .Q(\synth.voice.genblk4[7].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[123]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1402),
    .D(_01124_),
    .Q_N(_08140_),
    .Q(\synth.voice.genblk4[7].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[124]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1403),
    .D(_01125_),
    .Q_N(_08139_),
    .Q(\synth.voice.genblk4[7].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[125]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1404),
    .D(_01126_),
    .Q_N(_08138_),
    .Q(\synth.voice.genblk4[7].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[126]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1405),
    .D(_01127_),
    .Q_N(_08137_),
    .Q(\synth.voice.genblk4[7].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[127]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1406),
    .D(_01128_),
    .Q_N(_08136_),
    .Q(\synth.voice.genblk4[7].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[128]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1407),
    .D(_01129_),
    .Q_N(_00059_),
    .Q(\synth.voice.mods[2][8] ));
 sg13g2_dfrbp_1 \synth.voice.state[129]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1408),
    .D(_01130_),
    .Q_N(_00147_),
    .Q(\synth.voice.mods[2][9] ));
 sg13g2_dfrbp_1 \synth.voice.state[12]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1409),
    .D(_01131_),
    .Q_N(_00096_),
    .Q(\synth.voice.genblk4[0].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[130]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1410),
    .D(_01132_),
    .Q_N(_08135_),
    .Q(\synth.voice.genblk4[8].next_state_scan[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[131]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1411),
    .D(_01133_),
    .Q_N(_08134_),
    .Q(\synth.voice.genblk4[8].next_state_scan[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[132]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1412),
    .D(_01134_),
    .Q_N(_08133_),
    .Q(\synth.voice.genblk4[8].next_state_scan[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[133]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1413),
    .D(_01135_),
    .Q_N(_08132_),
    .Q(\synth.voice.genblk4[8].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[134]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1414),
    .D(_01136_),
    .Q_N(_08131_),
    .Q(\synth.voice.genblk4[8].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[135]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1415),
    .D(_01137_),
    .Q_N(_08130_),
    .Q(\synth.voice.genblk4[8].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[136]$_DFFE_PN_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1416),
    .D(_01138_),
    .Q_N(_00108_),
    .Q(\synth.voice.genblk4[8].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[137]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1417),
    .D(_01139_),
    .Q_N(_00109_),
    .Q(\synth.voice.genblk4[8].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.state[138]$_DFFE_PN_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1418),
    .D(_01140_),
    .Q_N(_00110_),
    .Q(\synth.voice.genblk4[8].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[139]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1419),
    .D(_01141_),
    .Q_N(_00092_),
    .Q(\synth.voice.genblk4[8].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[13]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1420),
    .D(_01142_),
    .Q_N(_00095_),
    .Q(\synth.voice.genblk4[0].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[140]$_DFFE_PN_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1421),
    .D(_01143_),
    .Q_N(_00094_),
    .Q(\synth.voice.genblk4[8].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[141]$_DFFE_PN_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1422),
    .D(_01144_),
    .Q_N(_00086_),
    .Q(\synth.voice.genblk4[8].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[142]$_DFFE_PN_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1423),
    .D(_01145_),
    .Q_N(_00088_),
    .Q(\synth.voice.genblk4[8].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[143]$_DFFE_PN_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1424),
    .D(_01146_),
    .Q_N(_00085_),
    .Q(\synth.voice.genblk4[8].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[144]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1425),
    .D(_01147_),
    .Q_N(_00058_),
    .Q(\synth.voice.params[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[145]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1426),
    .D(_01148_),
    .Q_N(_00081_),
    .Q(\synth.voice.params[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[146]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1427),
    .D(_01149_),
    .Q_N(_00082_),
    .Q(\synth.voice.genblk4[9].next_state_scan[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[147]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1428),
    .D(_01150_),
    .Q_N(_00083_),
    .Q(\synth.voice.genblk4[9].next_state_scan[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[148]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1429),
    .D(_01151_),
    .Q_N(_08129_),
    .Q(\synth.voice.genblk4[9].next_state_scan[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[149]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1430),
    .D(_01152_),
    .Q_N(_08128_),
    .Q(\synth.voice.genblk4[9].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[14]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1431),
    .D(_01153_),
    .Q_N(_00093_),
    .Q(\synth.voice.genblk4[0].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[150]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1432),
    .D(_01154_),
    .Q_N(_08127_),
    .Q(\synth.voice.genblk4[9].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[151]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1433),
    .D(_01155_),
    .Q_N(_08126_),
    .Q(\synth.voice.genblk4[9].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[152]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1434),
    .D(_01156_),
    .Q_N(_08125_),
    .Q(\synth.voice.genblk4[9].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[153]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1435),
    .D(_01157_),
    .Q_N(_08124_),
    .Q(\synth.voice.genblk4[9].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.state[154]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1436),
    .D(_01158_),
    .Q_N(_08123_),
    .Q(\synth.voice.genblk4[9].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[155]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1437),
    .D(_01159_),
    .Q_N(_08122_),
    .Q(\synth.voice.genblk4[9].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[156]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1438),
    .D(_01160_),
    .Q_N(_08121_),
    .Q(\synth.voice.genblk4[9].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[157]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1439),
    .D(_01161_),
    .Q_N(_08120_),
    .Q(\synth.voice.genblk4[9].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[158]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1440),
    .D(_01162_),
    .Q_N(_08119_),
    .Q(\synth.voice.genblk4[9].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[159]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1441),
    .D(_01163_),
    .Q_N(_08118_),
    .Q(\synth.voice.genblk4[9].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[15]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1442),
    .D(_01164_),
    .Q_N(_00091_),
    .Q(\synth.voice.genblk4[0].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[160]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1443),
    .D(_01165_),
    .Q_N(_08117_),
    .Q(\synth.voice.params[24] ));
 sg13g2_dfrbp_1 \synth.voice.state[161]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1444),
    .D(_01166_),
    .Q_N(_08116_),
    .Q(\synth.voice.params[25] ));
 sg13g2_dfrbp_1 \synth.voice.state[162]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1445),
    .D(_01167_),
    .Q_N(_08115_),
    .Q(\synth.voice.genblk4[10].next_state_scan[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[163]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1446),
    .D(_01168_),
    .Q_N(_08114_),
    .Q(\synth.voice.genblk4[10].next_state_scan[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[164]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1447),
    .D(_01169_),
    .Q_N(_08113_),
    .Q(\synth.voice.genblk4[10].next_state_scan[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[165]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1448),
    .D(_01170_),
    .Q_N(_08112_),
    .Q(\synth.voice.genblk4[10].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[166]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1449),
    .D(_01171_),
    .Q_N(_08111_),
    .Q(\synth.voice.genblk4[10].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[167]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1450),
    .D(_01172_),
    .Q_N(_08110_),
    .Q(\synth.voice.genblk4[10].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[168]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1451),
    .D(_01173_),
    .Q_N(_08109_),
    .Q(\synth.voice.genblk4[10].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[169]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1452),
    .D(_01174_),
    .Q_N(_08108_),
    .Q(\synth.voice.genblk4[10].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.state[16]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1453),
    .D(_01175_),
    .Q_N(_00060_),
    .Q(\synth.voice.lfsr[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[170]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1454),
    .D(_01176_),
    .Q_N(_08107_),
    .Q(\synth.voice.genblk4[10].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[171]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1455),
    .D(_01177_),
    .Q_N(_08106_),
    .Q(\synth.voice.genblk4[10].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[172]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1456),
    .D(_01178_),
    .Q_N(_08105_),
    .Q(\synth.voice.genblk4[10].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[173]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1457),
    .D(_01179_),
    .Q_N(_08104_),
    .Q(\synth.voice.genblk4[10].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[174]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1458),
    .D(_01180_),
    .Q_N(_08103_),
    .Q(\synth.voice.genblk4[10].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[175]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1459),
    .D(_01181_),
    .Q_N(_08102_),
    .Q(\synth.voice.genblk4[10].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[176]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1460),
    .D(_01182_),
    .Q_N(_00046_),
    .Q(\synth.voice.scan_outs[11][0] ));
 sg13g2_dfrbp_1 \synth.voice.state[177]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1461),
    .D(_01183_),
    .Q_N(_08101_),
    .Q(\synth.voice.scan_outs[11][1] ));
 sg13g2_dfrbp_1 \synth.voice.state[178]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1462),
    .D(_01184_),
    .Q_N(_08100_),
    .Q(\synth.voice.bpf_en[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[179]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1463),
    .D(_01185_),
    .Q_N(_08099_),
    .Q(\synth.voice.bpf_en[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[17]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1464),
    .D(_01186_),
    .Q_N(_00105_),
    .Q(\synth.voice.lfsr[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[180]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1465),
    .D(_01187_),
    .Q_N(_08098_),
    .Q(\synth.voice.bpf_en[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[181]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1466),
    .D(_01188_),
    .Q_N(_08097_),
    .Q(\synth.voice.genblk4[11].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[182]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1467),
    .D(_01189_),
    .Q_N(_08096_),
    .Q(\synth.voice.genblk4[11].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[183]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1468),
    .D(_01190_),
    .Q_N(_08095_),
    .Q(\synth.voice.genblk4[11].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[184]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1469),
    .D(_01191_),
    .Q_N(_08094_),
    .Q(\synth.voice.genblk4[11].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[185]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1470),
    .D(_01192_),
    .Q_N(_08093_),
    .Q(\synth.voice.genblk4[11].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.state[186]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1471),
    .D(_01193_),
    .Q_N(_00163_),
    .Q(\synth.voice.genblk4[11].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[187]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1472),
    .D(_01194_),
    .Q_N(_00171_),
    .Q(\synth.voice.genblk4[11].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[188]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1473),
    .D(_01195_),
    .Q_N(_08092_),
    .Q(\synth.voice.genblk4[11].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[189]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1474),
    .D(_01196_),
    .Q_N(_08091_),
    .Q(\synth.voice.genblk4[11].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[18]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1475),
    .D(_01197_),
    .Q_N(_00103_),
    .Q(\synth.voice.genblk4[1].next_state_scan[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[190]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1476),
    .D(_01198_),
    .Q_N(_08090_),
    .Q(\synth.voice.genblk4[11].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[191]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1477),
    .D(_01199_),
    .Q_N(_08089_),
    .Q(\synth.voice.genblk4[11].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[19]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1478),
    .D(_01200_),
    .Q_N(_00101_),
    .Q(\synth.voice.genblk4[1].next_state_scan[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[1]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1479),
    .D(_01201_),
    .Q_N(_08088_),
    .Q(\synth.voice.delayed_p[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[20]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1480),
    .D(_01202_),
    .Q_N(_00099_),
    .Q(\synth.voice.genblk4[1].next_state_scan[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[21]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1481),
    .D(_01203_),
    .Q_N(_00097_),
    .Q(\synth.voice.genblk4[1].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[22]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1482),
    .D(_01204_),
    .Q_N(_00090_),
    .Q(\synth.voice.genblk4[1].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[23]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1483),
    .D(_01205_),
    .Q_N(_00089_),
    .Q(\synth.voice.genblk4[1].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[24]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1484),
    .D(_01206_),
    .Q_N(_00087_),
    .Q(\synth.voice.genblk4[1].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[25]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1485),
    .D(_01207_),
    .Q_N(_00084_),
    .Q(\synth.voice.genblk4[1].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.state[26]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1486),
    .D(_01208_),
    .Q_N(_08087_),
    .Q(\synth.voice.genblk4[1].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[27]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1487),
    .D(_01209_),
    .Q_N(_00139_),
    .Q(\synth.voice.genblk4[1].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[28]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1488),
    .D(_01210_),
    .Q_N(_00140_),
    .Q(\synth.voice.genblk4[1].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[29]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1489),
    .D(_01211_),
    .Q_N(_00141_),
    .Q(\synth.voice.genblk4[1].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1490),
    .D(_01212_),
    .Q_N(_08086_),
    .Q(\synth.voice.delayed_p[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[30]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1491),
    .D(_01213_),
    .Q_N(_00142_),
    .Q(\synth.voice.genblk4[1].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[31]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1492),
    .D(_01214_),
    .Q_N(_00143_),
    .Q(\synth.voice.genblk4[1].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[32]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1493),
    .D(_01215_),
    .Q_N(_08085_),
    .Q(\synth.voice.scan_outs[2][0] ));
 sg13g2_dfrbp_1 \synth.voice.state[33]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1494),
    .D(_01216_),
    .Q_N(_08084_),
    .Q(\synth.voice.scan_outs[2][1] ));
 sg13g2_dfrbp_1 \synth.voice.state[34]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1495),
    .D(_01217_),
    .Q_N(_08083_),
    .Q(\synth.voice.genblk4[2].next_state_scan[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[35]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1496),
    .D(_01218_),
    .Q_N(_08082_),
    .Q(\synth.voice.genblk4[2].next_state_scan[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[36]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1497),
    .D(_01219_),
    .Q_N(_08081_),
    .Q(\synth.voice.genblk4[2].next_state_scan[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[37]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1498),
    .D(_01220_),
    .Q_N(_08080_),
    .Q(\synth.voice.genblk4[2].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[38]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1499),
    .D(_01221_),
    .Q_N(_08079_),
    .Q(\synth.voice.genblk4[2].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[39]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1500),
    .D(_01222_),
    .Q_N(_08078_),
    .Q(\synth.voice.genblk4[2].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[3]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1501),
    .D(_01223_),
    .Q_N(_00053_),
    .Q(\synth.voice.coeff_index[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[40]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1502),
    .D(_01224_),
    .Q_N(_08077_),
    .Q(\synth.voice.genblk4[2].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[41]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1503),
    .D(_01225_),
    .Q_N(_08076_),
    .Q(\synth.voice.genblk4[2].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.state[42]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1504),
    .D(_01226_),
    .Q_N(_08075_),
    .Q(\synth.voice.genblk4[2].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[43]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1505),
    .D(_01227_),
    .Q_N(_08074_),
    .Q(\synth.voice.genblk4[2].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[44]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1506),
    .D(_01228_),
    .Q_N(_08073_),
    .Q(\synth.voice.genblk4[2].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[45]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1507),
    .D(_01229_),
    .Q_N(_08072_),
    .Q(\synth.voice.genblk4[2].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[46]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1508),
    .D(_01230_),
    .Q_N(_08071_),
    .Q(\synth.voice.genblk4[2].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[47]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1509),
    .D(_01231_),
    .Q_N(_08070_),
    .Q(\synth.voice.genblk4[2].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[48]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1510),
    .D(_01232_),
    .Q_N(_08069_),
    .Q(\synth.voice.scan_outs[3][0] ));
 sg13g2_dfrbp_1 \synth.voice.state[49]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1511),
    .D(_01233_),
    .Q_N(_08068_),
    .Q(\synth.voice.scan_outs[3][1] ));
 sg13g2_dfrbp_1 \synth.voice.state[4]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1512),
    .D(_01234_),
    .Q_N(_08067_),
    .Q(\synth.voice.coeff_index[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[50]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1513),
    .D(_01235_),
    .Q_N(_08066_),
    .Q(\synth.voice.genblk4[3].next_state_scan[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[51]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1514),
    .D(_01236_),
    .Q_N(_08065_),
    .Q(\synth.voice.genblk4[3].next_state_scan[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[52]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1515),
    .D(_01237_),
    .Q_N(_08064_),
    .Q(\synth.voice.genblk4[3].next_state_scan[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[53]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1516),
    .D(_01238_),
    .Q_N(_08063_),
    .Q(\synth.voice.genblk4[3].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[54]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1517),
    .D(_01239_),
    .Q_N(_08062_),
    .Q(\synth.voice.genblk4[3].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[55]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1518),
    .D(_01240_),
    .Q_N(_08061_),
    .Q(\synth.voice.genblk4[3].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[56]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1519),
    .D(_01241_),
    .Q_N(_08060_),
    .Q(\synth.voice.genblk4[3].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[57]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1520),
    .D(_01242_),
    .Q_N(_08059_),
    .Q(\synth.voice.genblk4[3].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.state[58]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1521),
    .D(_01243_),
    .Q_N(_08058_),
    .Q(\synth.voice.genblk4[3].next_state_scan[8] ));
 sg13g2_dfrbp_1 \synth.voice.state[59]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1522),
    .D(_01244_),
    .Q_N(_08057_),
    .Q(\synth.voice.genblk4[3].next_state_scan[9] ));
 sg13g2_dfrbp_1 \synth.voice.state[5]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1523),
    .D(_01245_),
    .Q_N(_08056_),
    .Q(\synth.voice.coeff_index[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[60]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1524),
    .D(_01246_),
    .Q_N(_08055_),
    .Q(\synth.voice.genblk4[3].next_state_scan[10] ));
 sg13g2_dfrbp_1 \synth.voice.state[61]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1525),
    .D(_01247_),
    .Q_N(_08054_),
    .Q(\synth.voice.genblk4[3].next_state_scan[11] ));
 sg13g2_dfrbp_1 \synth.voice.state[62]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1526),
    .D(_01248_),
    .Q_N(_08053_),
    .Q(\synth.voice.genblk4[3].next_state_scan[12] ));
 sg13g2_dfrbp_1 \synth.voice.state[63]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1527),
    .D(_01249_),
    .Q_N(_08052_),
    .Q(\synth.voice.genblk4[3].next_state_scan[13] ));
 sg13g2_dfrbp_1 \synth.voice.state[64]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1528),
    .D(_01250_),
    .Q_N(_08051_),
    .Q(\synth.voice.scan_outs[4][0] ));
 sg13g2_dfrbp_1 \synth.voice.state[65]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1529),
    .D(_01251_),
    .Q_N(_08050_),
    .Q(\synth.voice.scan_outs[4][1] ));
 sg13g2_dfrbp_1 \synth.voice.state[66]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1530),
    .D(_01252_),
    .Q_N(_08049_),
    .Q(\synth.voice.genblk4[4].next_state_scan[0] ));
 sg13g2_dfrbp_1 \synth.voice.state[67]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1531),
    .D(_01253_),
    .Q_N(_08048_),
    .Q(\synth.voice.genblk4[4].next_state_scan[1] ));
 sg13g2_dfrbp_1 \synth.voice.state[68]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1532),
    .D(_01254_),
    .Q_N(_08047_),
    .Q(\synth.voice.genblk4[4].next_state_scan[2] ));
 sg13g2_dfrbp_1 \synth.voice.state[69]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1533),
    .D(_01255_),
    .Q_N(_08046_),
    .Q(\synth.voice.genblk4[4].next_state_scan[3] ));
 sg13g2_dfrbp_1 \synth.voice.state[6]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1534),
    .D(_01256_),
    .Q_N(_00107_),
    .Q(\synth.voice.genblk4[0].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[70]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1535),
    .D(_01257_),
    .Q_N(_08045_),
    .Q(\synth.voice.genblk4[4].next_state_scan[4] ));
 sg13g2_dfrbp_1 \synth.voice.state[71]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1536),
    .D(_01258_),
    .Q_N(_08044_),
    .Q(\synth.voice.genblk4[4].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[72]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1537),
    .D(_01259_),
    .Q_N(_00137_),
    .Q(\synth.voice.float_period[0][0] ));
 sg13g2_dfrbp_1 \synth.voice.state[73]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1538),
    .D(_01260_),
    .Q_N(_00135_),
    .Q(\synth.voice.float_period[0][1] ));
 sg13g2_dfrbp_1 \synth.voice.state[74]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1539),
    .D(_01261_),
    .Q_N(_00133_),
    .Q(\synth.voice.float_period[0][2] ));
 sg13g2_dfrbp_1 \synth.voice.state[75]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1540),
    .D(_01262_),
    .Q_N(_08043_),
    .Q(\synth.voice.float_period[0][3] ));
 sg13g2_dfrbp_1 \synth.voice.state[76]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1541),
    .D(_01263_),
    .Q_N(_08042_),
    .Q(\synth.voice.float_period[0][4] ));
 sg13g2_dfrbp_1 \synth.voice.state[77]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1542),
    .D(_01264_),
    .Q_N(_08041_),
    .Q(\synth.voice.float_period[0][5] ));
 sg13g2_dfrbp_1 \synth.voice.state[78]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1543),
    .D(_01265_),
    .Q_N(_08040_),
    .Q(\synth.voice.float_period[0][6] ));
 sg13g2_dfrbp_1 \synth.voice.state[79]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1544),
    .D(_01266_),
    .Q_N(_08039_),
    .Q(\synth.voice.float_period[0][7] ));
 sg13g2_dfrbp_1 \synth.voice.state[7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1545),
    .D(_01267_),
    .Q_N(_00106_),
    .Q(\synth.voice.genblk4[0].next_state_scan[5] ));
 sg13g2_dfrbp_1 \synth.voice.state[80]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1546),
    .D(_01268_),
    .Q_N(_08038_),
    .Q(\synth.voice.float_period[0][8] ));
 sg13g2_dfrbp_1 \synth.voice.state[81]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1547),
    .D(_01269_),
    .Q_N(_08037_),
    .Q(\synth.voice.float_period[0][9] ));
 sg13g2_dfrbp_1 \synth.voice.state[82]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1548),
    .D(_01270_),
    .Q_N(_08036_),
    .Q(\synth.voice.float_period[0][10] ));
 sg13g2_dfrbp_1 \synth.voice.state[83]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1549),
    .D(_01271_),
    .Q_N(_00114_),
    .Q(\synth.voice.float_period[0][11] ));
 sg13g2_dfrbp_1 \synth.voice.state[84]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1550),
    .D(_01272_),
    .Q_N(_08035_),
    .Q(\synth.voice.float_period[0][12] ));
 sg13g2_dfrbp_1 \synth.voice.state[85]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1551),
    .D(_01273_),
    .Q_N(_08034_),
    .Q(\synth.voice.float_period[0][13] ));
 sg13g2_dfrbp_1 \synth.voice.state[86]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1552),
    .D(_01274_),
    .Q_N(_00138_),
    .Q(\synth.voice.float_period[1][0] ));
 sg13g2_dfrbp_1 \synth.voice.state[87]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1553),
    .D(_01275_),
    .Q_N(_00136_),
    .Q(\synth.voice.float_period[1][1] ));
 sg13g2_dfrbp_1 \synth.voice.state[88]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1554),
    .D(_01276_),
    .Q_N(_00134_),
    .Q(\synth.voice.float_period[1][2] ));
 sg13g2_dfrbp_1 \synth.voice.state[89]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1555),
    .D(_01277_),
    .Q_N(_08033_),
    .Q(\synth.voice.float_period[1][3] ));
 sg13g2_dfrbp_1 \synth.voice.state[8]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1556),
    .D(_01278_),
    .Q_N(_00104_),
    .Q(\synth.voice.genblk4[0].next_state_scan[6] ));
 sg13g2_dfrbp_1 \synth.voice.state[90]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1557),
    .D(_01279_),
    .Q_N(_08032_),
    .Q(\synth.voice.float_period[1][4] ));
 sg13g2_dfrbp_1 \synth.voice.state[91]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1558),
    .D(_01280_),
    .Q_N(_08031_),
    .Q(\synth.voice.float_period[1][5] ));
 sg13g2_dfrbp_1 \synth.voice.state[92]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1559),
    .D(_01281_),
    .Q_N(_08030_),
    .Q(\synth.voice.float_period[1][6] ));
 sg13g2_dfrbp_1 \synth.voice.state[93]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1560),
    .D(_01282_),
    .Q_N(_08029_),
    .Q(\synth.voice.float_period[1][7] ));
 sg13g2_dfrbp_1 \synth.voice.state[94]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1561),
    .D(_01283_),
    .Q_N(_08028_),
    .Q(\synth.voice.float_period[1][8] ));
 sg13g2_dfrbp_1 \synth.voice.state[95]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1562),
    .D(_01284_),
    .Q_N(_08027_),
    .Q(\synth.voice.float_period[1][9] ));
 sg13g2_dfrbp_1 \synth.voice.state[96]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1563),
    .D(_01285_),
    .Q_N(_08026_),
    .Q(\synth.voice.float_period[1][10] ));
 sg13g2_dfrbp_1 \synth.voice.state[97]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1564),
    .D(_01286_),
    .Q_N(_00115_),
    .Q(\synth.voice.float_period[1][11] ));
 sg13g2_dfrbp_1 \synth.voice.state[98]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1565),
    .D(_01287_),
    .Q_N(_08025_),
    .Q(\synth.voice.float_period[1][12] ));
 sg13g2_dfrbp_1 \synth.voice.state[99]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1566),
    .D(_01288_),
    .Q_N(_08024_),
    .Q(\synth.voice.float_period[1][13] ));
 sg13g2_dfrbp_1 \synth.voice.state[9]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1567),
    .D(_01289_),
    .Q_N(_00102_),
    .Q(\synth.voice.genblk4[0].next_state_scan[7] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1568),
    .D(_01290_),
    .Q_N(\synth.voice.next_sweep_oct_counter[0] ),
    .Q(\synth.voice.sweep_oct_counter[0] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1569),
    .D(_01291_),
    .Q_N(_08023_),
    .Q(\synth.voice.sweep_oct_counter[10] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1570),
    .D(_01292_),
    .Q_N(_08022_),
    .Q(\synth.voice.sweep_oct_counter[11] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[12]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1571),
    .D(_01293_),
    .Q_N(_08021_),
    .Q(\synth.voice.sweep_oct_counter[12] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[13]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1572),
    .D(_01294_),
    .Q_N(_08020_),
    .Q(\synth.voice.sweep_oct_counter[13] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1573),
    .D(_01295_),
    .Q_N(_08019_),
    .Q(\synth.voice.sweep_oct_counter[1] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1574),
    .D(_01296_),
    .Q_N(_08018_),
    .Q(\synth.voice.sweep_oct_counter[2] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1575),
    .D(_01297_),
    .Q_N(_08017_),
    .Q(\synth.voice.sweep_oct_counter[3] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1576),
    .D(_01298_),
    .Q_N(_08016_),
    .Q(\synth.voice.sweep_oct_counter[4] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1577),
    .D(_01299_),
    .Q_N(_08015_),
    .Q(\synth.voice.sweep_oct_counter[5] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1578),
    .D(_01300_),
    .Q_N(_08014_),
    .Q(\synth.voice.sweep_oct_counter[6] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1579),
    .D(_01301_),
    .Q_N(_08013_),
    .Q(\synth.voice.sweep_oct_counter[7] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1580),
    .D(_01302_),
    .Q_N(_08012_),
    .Q(\synth.voice.sweep_oct_counter[8] ));
 sg13g2_dfrbp_1 \synth.voice.sweep_oct_counter[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1581),
    .D(_01303_),
    .Q_N(_08011_),
    .Q(\synth.voice.sweep_oct_counter[9] ));
 sg13g2_dfrbp_1 \synth.voice.tap[0]$_SDFF_PP0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1582),
    .D(_01304_),
    .Q_N(_00049_),
    .Q(\synth.controller.tap_pos[0] ));
 sg13g2_dfrbp_1 \synth.voice.tap[1]$_SDFF_PP0_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1583),
    .D(_01305_),
    .Q_N(_09025_),
    .Q(\synth.controller.tap_pos[1] ));
 sg13g2_dfrbp_1 \synth.voice.target_reg[1]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1584),
    .D(_00008_),
    .Q_N(_09026_),
    .Q(\synth.voice.target_reg[1] ));
 sg13g2_dfrbp_1 \synth.voice.target_reg[2]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1585),
    .D(_00009_),
    .Q_N(_09027_),
    .Q(\synth.voice.target_reg[2] ));
 sg13g2_dfrbp_1 \synth.voice.target_reg[3]$_DFF_P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1586),
    .D(_00010_),
    .Q_N(_08010_),
    .Q(\synth.voice.target_reg[3] ));
 sg13g2_dfrbp_1 \synth.voice.term_index[0]$_SDFF_PP0_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1587),
    .D(_01306_),
    .Q_N(_00048_),
    .Q(\synth.voice.fir_table.i_term[0] ));
 sg13g2_dfrbp_1 \synth.voice.term_index[1]$_SDFF_PP0_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1588),
    .D(_01307_),
    .Q_N(_08009_),
    .Q(\synth.voice.fir_table.i_term[1] ));
 sg13g2_dfrbp_1 \synth.voice.term_index[2]$_SDFF_PP0_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1589),
    .D(_01308_),
    .Q_N(_00045_),
    .Q(\synth.voice.fir_table.i_term[2] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1590),
    .D(_01309_),
    .Q_N(_08008_),
    .Q(\synth.voice.wave_reg[0] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1591),
    .D(_01310_),
    .Q_N(_08007_),
    .Q(\synth.voice.wave_reg[1] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1592),
    .D(_01311_),
    .Q_N(_08006_),
    .Q(\synth.voice.wave_reg[2] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1593),
    .D(_01312_),
    .Q_N(_08005_),
    .Q(\synth.voice.wave_reg[3] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[4]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1594),
    .D(_01313_),
    .Q_N(_08004_),
    .Q(\synth.voice.wave_reg[4] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[5]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1595),
    .D(_01314_),
    .Q_N(_08003_),
    .Q(\synth.voice.wave_reg[5] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[6]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1596),
    .D(_01315_),
    .Q_N(_08002_),
    .Q(\synth.voice.wave_reg[6] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1597),
    .D(_01316_),
    .Q_N(_08001_),
    .Q(\synth.voice.wave_reg[7] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1598),
    .D(_01317_),
    .Q_N(_08000_),
    .Q(\synth.voice.wave_reg[8] ));
 sg13g2_dfrbp_1 \synth.voice.wave_reg[9]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1599),
    .D(_01318_),
    .Q_N(_09028_),
    .Q(\synth.voice.wave_reg[9] ));
 sg13g2_dfrbp_1 \synth.voice.zero_shifter_out_reg$_DFF_P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1600),
    .D(\synth.voice.zero_shifter_out ),
    .Q_N(_00144_),
    .Q(\synth.voice.zero_shifter_out_reg ));
 sg13g2_dfrbp_1 \ui_in_reg[0]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1601),
    .D(net2),
    .Q_N(_09029_),
    .Q(\data_pins[0] ));
 sg13g2_dfrbp_1 \ui_in_reg[1]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1602),
    .D(net3),
    .Q_N(_09030_),
    .Q(\data_pins[1] ));
 sg13g2_dfrbp_1 \ui_in_reg[2]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1603),
    .D(net4),
    .Q_N(_09031_),
    .Q(\data_pins[2] ));
 sg13g2_dfrbp_1 \ui_in_reg[3]$_DFF_P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1604),
    .D(net5),
    .Q_N(_09032_),
    .Q(\data_pins[3] ));
 sg13g2_dfrbp_1 \uio_out_reg[0]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1605),
    .D(\addr_pins_out[0] ),
    .Q_N(_09033_),
    .Q(net12));
 sg13g2_dfrbp_1 \uio_out_reg[1]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1606),
    .D(\addr_pins_out[1] ),
    .Q_N(_09034_),
    .Q(net13));
 sg13g2_dfrbp_1 \uio_out_reg[2]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1607),
    .D(\addr_pins_out[2] ),
    .Q_N(_09035_),
    .Q(net14));
 sg13g2_dfrbp_1 \uio_out_reg[3]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1608),
    .D(\addr_pins_out[3] ),
    .Q_N(_09036_),
    .Q(net15));
 sg13g2_dfrbp_1 \uio_out_reg[4]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1609),
    .D(\synth.controller.sbio_tx.start_present ),
    .Q_N(_07999_),
    .Q(net16));
 sg13g2_dfrbp_1 \uio_out_reg[5]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1610),
    .D(_01319_),
    .Q_N(_09037_),
    .Q(net17));
 sg13g2_dfrbp_1 \uio_out_reg[6]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1611),
    .D(\uio_out0[6] ),
    .Q_N(_09038_),
    .Q(net18));
 sg13g2_dfrbp_1 \uio_out_reg[7]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1612),
    .D(\uio_out0[7] ),
    .Q_N(_09039_),
    .Q(net19));
 sg13g2_dfrbp_1 \uo_out_reg[0]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1613),
    .D(\uo_out0[0] ),
    .Q_N(_09040_),
    .Q(net20));
 sg13g2_dfrbp_1 \uo_out_reg[1]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1614),
    .D(\uo_out0[1] ),
    .Q_N(_09041_),
    .Q(net21));
 sg13g2_dfrbp_1 \uo_out_reg[2]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1615),
    .D(\uo_out0[2] ),
    .Q_N(_09042_),
    .Q(net22));
 sg13g2_dfrbp_1 \uo_out_reg[3]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1616),
    .D(\ppu.vsync ),
    .Q_N(_09043_),
    .Q(net23));
 sg13g2_dfrbp_1 \uo_out_reg[4]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1617),
    .D(\uo_out0[4] ),
    .Q_N(_09044_),
    .Q(net24));
 sg13g2_dfrbp_1 \uo_out_reg[5]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1618),
    .D(\uo_out0[5] ),
    .Q_N(_09045_),
    .Q(net25));
 sg13g2_dfrbp_1 \uo_out_reg[6]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1619),
    .D(\uo_out0[6] ),
    .Q_N(_09046_),
    .Q(net26));
 sg13g2_dfrbp_1 \uo_out_reg[7]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1620),
    .D(hsync),
    .Q_N(_07998_),
    .Q(net27));
 sg13g2_dfrbp_1 \vblank_pending$_SDFF_PP0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1621),
    .D(_01320_),
    .Q_N(_07997_),
    .Q(\synth.controller.ext_tx_request ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[7]),
    .X(net9));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[6]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[7]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[0]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[1]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[2]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[4]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[5]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[6]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[7]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[0]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[1]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[2]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[3]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[4]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[5]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[6]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout28 (.A(_03125_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_05950_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_04034_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_03138_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_05953_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_05862_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_04698_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_04317_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_04240_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_04046_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_06349_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_06308_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_06263_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_06221_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_04797_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_04207_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_04206_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_05523_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_03001_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_03000_),
    .X(net47));
 sg13g2_buf_4 fanout48 (.X(net48),
    .A(_02999_));
 sg13g2_buf_2 fanout49 (.A(_02998_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_02979_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_02978_),
    .X(net51));
 sg13g2_buf_4 fanout52 (.X(net52),
    .A(_02977_));
 sg13g2_buf_2 fanout53 (.A(_02976_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_02957_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_02956_),
    .X(net55));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(_02955_));
 sg13g2_buf_2 fanout57 (.A(_02954_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_02935_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_02934_),
    .X(net59));
 sg13g2_buf_4 fanout60 (.X(net60),
    .A(_02933_));
 sg13g2_buf_2 fanout61 (.A(_02932_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_06481_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_06443_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_06376_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_05522_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_05515_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_07029_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_06883_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_06423_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_06143_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_05514_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_03059_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_07448_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_06332_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_06292_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_06290_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_06280_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_06274_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_06246_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_06197_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_06194_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_06178_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_06171_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_06167_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_06154_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_02920_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_02910_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_02900_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_02889_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_06139_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_02424_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_07538_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_06996_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_06924_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_06881_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_06863_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_02628_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_02609_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_02464_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_02437_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_02423_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_02390_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_07556_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_06989_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_02627_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_02608_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_02463_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_02389_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_07569_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_07529_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_07430_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_06354_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_06313_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_06268_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_06227_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_02659_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_02647_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_07568_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_02658_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_02646_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_02580_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_02259_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_06963_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_05829_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_05536_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_05531_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_04803_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_04440_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_01546_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_05919_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_05828_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_05793_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_05790_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_04802_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_04708_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_04702_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_04412_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_04262_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_04212_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_04092_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_04047_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_03629_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_03422_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_02806_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_02058_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_01913_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_06854_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_05915_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_05911_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_05859_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_05738_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_05533_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_04799_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_04438_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_04433_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_04258_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_04042_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_04036_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_03628_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_03615_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_02853_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_02838_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_02824_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_01533_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_07590_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_05914_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_05910_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_05735_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_05527_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_04763_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_04760_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_04759_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_04474_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_04456_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_04450_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_04358_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_04355_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_04265_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_04254_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_04230_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_04210_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_03612_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_03448_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_02262_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_06580_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_04817_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_04816_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_04723_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_04711_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_04462_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_04421_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_03456_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_03419_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_03253_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_03218_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_03217_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_03207_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_02518_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_02517_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_02236_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_01764_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_01740_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_07694_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_06703_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_06697_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_06501_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_05328_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_04815_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_04722_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_04721_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_03418_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_03325_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_03313_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_03260_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_03195_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_02481_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_07692_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_06710_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_06702_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_03417_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_02786_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_02784_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_02760_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_02753_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_02752_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_02737_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_02735_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_02717_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_02715_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_02698_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_02696_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_02678_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_02676_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_02532_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_02501_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_02234_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_02182_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_07552_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_07523_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_06504_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_06503_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_03434_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_03416_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_03193_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_03161_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_02927_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_02881_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_02714_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_02221_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_02198_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_02140_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_02108_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_02051_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_01905_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_01775_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_07727_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_07548_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_02197_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_02109_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_01944_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_01927_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_01921_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_01904_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_01891_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_01797_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_07726_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_07396_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_07393_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_07373_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_07370_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_07350_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_07347_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_07327_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_07324_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_07304_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_07301_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_07281_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_07278_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_07258_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_07254_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_07234_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_07231_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_07211_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_07209_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_07191_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_07188_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_07164_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_07137_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_07064_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_06846_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_03809_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_03739_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_03247_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_03085_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_02576_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_01926_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_01890_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_01800_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_01773_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_01745_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_07431_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_07395_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_07372_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_07349_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_07326_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_07303_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_07280_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_07256_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_07233_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_07210_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_07190_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_07166_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_07159_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_07157_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_07142_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_07140_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_07055_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_07052_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_06845_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_06222_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_05198_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_05135_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_05073_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_05071_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_05068_),
    .X(net325));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_05013_));
 sg13g2_buf_2 fanout327 (.A(_05002_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_04087_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_03889_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_03810_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_03801_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_03742_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_03735_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_03729_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_02688_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_02686_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_02406_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_02402_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_02398_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_02394_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_02306_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_02299_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_02053_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_01933_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_01857_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_01823_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_01817_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_07686_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_07181_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_07045_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_07000_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_06831_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_06827_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_06826_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_05201_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_05164_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_05152_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_05137_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_05109_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_05105_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_05103_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_05055_),
    .X(net362));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(_05046_));
 sg13g2_buf_2 fanout364 (.A(_05038_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_05035_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_05029_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_05023_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_05020_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_05011_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_04991_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_04989_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_04074_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_04039_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_03952_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_03835_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_03723_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_03371_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_03319_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_03315_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_03300_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_02721_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_02505_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_02494_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_02485_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_02418_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_02415_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_02409_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_02291_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_02285_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_02063_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_01918_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_01822_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_01805_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_01790_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_06999_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_06519_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_05036_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_05028_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_04992_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_03423_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_03379_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_03372_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_02493_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_02489_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_02484_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_02411_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_02264_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_01866_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_01821_),
    .X(net409));
 sg13g2_tiehi _16921__410 (.L_HI(net410));
 sg13g2_tiehi _16922__411 (.L_HI(net411));
 sg13g2_tiehi _16923__412 (.L_HI(net412));
 sg13g2_tiehi _16924__413 (.L_HI(net413));
 sg13g2_tiehi _16925__414 (.L_HI(net414));
 sg13g2_tiehi _16926__415 (.L_HI(net415));
 sg13g2_tiehi \cfg[0]$_DFFE_PN__416  (.L_HI(net416));
 sg13g2_tiehi \ppu.avhsync_delayed[0]$_DFFE_PP__417  (.L_HI(net417));
 sg13g2_tiehi \ppu.avhsync_delayed[1]$_DFFE_PP__418  (.L_HI(net418));
 sg13g2_tiehi \ppu.avhsync_delayed[2]$_DFFE_PP__419  (.L_HI(net419));
 sg13g2_tiehi \ppu.base_addr_regs[0][0]$_DFFE_PP__420  (.L_HI(net420));
 sg13g2_tiehi \ppu.base_addr_regs[0][1]$_DFFE_PP__421  (.L_HI(net421));
 sg13g2_tiehi \ppu.base_addr_regs[0][2]$_DFFE_PP__422  (.L_HI(net422));
 sg13g2_tiehi \ppu.base_addr_regs[0][3]$_DFFE_PP__423  (.L_HI(net423));
 sg13g2_tiehi \ppu.base_addr_regs[0][4]$_DFFE_PP__424  (.L_HI(net424));
 sg13g2_tiehi \ppu.base_addr_regs[0][5]$_DFFE_PP__425  (.L_HI(net425));
 sg13g2_tiehi \ppu.base_addr_regs[0][6]$_DFFE_PP__426  (.L_HI(net426));
 sg13g2_tiehi \ppu.base_addr_regs[0][7]$_DFFE_PP__427  (.L_HI(net427));
 sg13g2_tiehi \ppu.base_addr_regs[0][8]$_DFFE_PP__428  (.L_HI(net428));
 sg13g2_tiehi \ppu.base_addr_regs[1][0]$_DFFE_PP__429  (.L_HI(net429));
 sg13g2_tiehi \ppu.base_addr_regs[1][1]$_DFFE_PP__430  (.L_HI(net430));
 sg13g2_tiehi \ppu.base_addr_regs[1][2]$_DFFE_PP__431  (.L_HI(net431));
 sg13g2_tiehi \ppu.base_addr_regs[1][3]$_DFFE_PP__432  (.L_HI(net432));
 sg13g2_tiehi \ppu.base_addr_regs[1][4]$_DFFE_PP__433  (.L_HI(net433));
 sg13g2_tiehi \ppu.base_addr_regs[1][5]$_DFFE_PP__434  (.L_HI(net434));
 sg13g2_tiehi \ppu.base_addr_regs[1][6]$_DFFE_PP__435  (.L_HI(net435));
 sg13g2_tiehi \ppu.base_addr_regs[1][7]$_DFFE_PP__436  (.L_HI(net436));
 sg13g2_tiehi \ppu.base_addr_regs[1][8]$_DFFE_PP__437  (.L_HI(net437));
 sg13g2_tiehi \ppu.base_addr_regs[2][1]$_DFFE_PP__438  (.L_HI(net438));
 sg13g2_tiehi \ppu.base_addr_regs[2][2]$_DFFE_PP__439  (.L_HI(net439));
 sg13g2_tiehi \ppu.base_addr_regs[2][3]$_DFFE_PP__440  (.L_HI(net440));
 sg13g2_tiehi \ppu.base_addr_regs[2][4]$_DFFE_PP__441  (.L_HI(net441));
 sg13g2_tiehi \ppu.base_addr_regs[2][5]$_DFFE_PP__442  (.L_HI(net442));
 sg13g2_tiehi \ppu.base_addr_regs[2][6]$_DFFE_PP__443  (.L_HI(net443));
 sg13g2_tiehi \ppu.base_addr_regs[2][7]$_DFFE_PP__444  (.L_HI(net444));
 sg13g2_tiehi \ppu.base_addr_regs[2][8]$_DFFE_PP__445  (.L_HI(net445));
 sg13g2_tiehi \ppu.base_addr_regs[3][1]$_DFFE_PP__446  (.L_HI(net446));
 sg13g2_tiehi \ppu.base_addr_regs[3][2]$_DFFE_PP__447  (.L_HI(net447));
 sg13g2_tiehi \ppu.base_addr_regs[3][3]$_DFFE_PP__448  (.L_HI(net448));
 sg13g2_tiehi \ppu.base_addr_regs[3][4]$_DFFE_PP__449  (.L_HI(net449));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[0]$_SDFF_PP0__450  (.L_HI(net450));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[10]$_SDFF_PP1__451  (.L_HI(net451));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[11]$_SDFF_PP1__452  (.L_HI(net452));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[12]$_SDFF_PP1__453  (.L_HI(net453));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[13]$_SDFF_PP1__454  (.L_HI(net454));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[14]$_SDFF_PP1__455  (.L_HI(net455));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[15]$_SDFF_PP1__456  (.L_HI(net456));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[1]$_SDFF_PP1__457  (.L_HI(net457));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[2]$_SDFF_PP1__458  (.L_HI(net458));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[3]$_SDFF_PP1__459  (.L_HI(net459));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[4]$_SDFF_PP1__460  (.L_HI(net460));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[5]$_SDFF_PP1__461  (.L_HI(net461));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[6]$_SDFF_PP1__462  (.L_HI(net462));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[7]$_SDFF_PP1__463  (.L_HI(net463));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[8]$_SDFF_PP1__464  (.L_HI(net464));
 sg13g2_tiehi \ppu.copper_inst.addr_reg[9]$_SDFF_PP1__465  (.L_HI(net465));
 sg13g2_tiehi \ppu.copper_inst.cmp[0]$_DFFE_PP__466  (.L_HI(net466));
 sg13g2_tiehi \ppu.copper_inst.cmp[1]$_DFFE_PP__467  (.L_HI(net467));
 sg13g2_tiehi \ppu.copper_inst.cmp[2]$_DFFE_PP__468  (.L_HI(net468));
 sg13g2_tiehi \ppu.copper_inst.cmp[3]$_DFFE_PP__469  (.L_HI(net469));
 sg13g2_tiehi \ppu.copper_inst.cmp[4]$_DFFE_PP__470  (.L_HI(net470));
 sg13g2_tiehi \ppu.copper_inst.cmp[5]$_DFFE_PP__471  (.L_HI(net471));
 sg13g2_tiehi \ppu.copper_inst.cmp[6]$_DFFE_PP__472  (.L_HI(net472));
 sg13g2_tiehi \ppu.copper_inst.cmp[7]$_DFFE_PP__473  (.L_HI(net473));
 sg13g2_tiehi \ppu.copper_inst.cmp[8]$_DFFE_PP__474  (.L_HI(net474));
 sg13g2_tiehi \ppu.copper_inst.cmp_on$_SDFFE_PP0P__475  (.L_HI(net475));
 sg13g2_tiehi \ppu.copper_inst.cmp_type$_DFFE_PP__476  (.L_HI(net476));
 sg13g2_tiehi \ppu.copper_inst.fast_mode$_DFF_P__477  (.L_HI(net477));
 sg13g2_tiehi \ppu.copper_inst.on$_DFFE_PP__478  (.L_HI(net478));
 sg13g2_tiehi \ppu.copper_inst.store[0]$_DFFE_PP__479  (.L_HI(net479));
 sg13g2_tiehi \ppu.copper_inst.store[10]$_DFFE_PP__480  (.L_HI(net480));
 sg13g2_tiehi \ppu.copper_inst.store[11]$_DFFE_PP__481  (.L_HI(net481));
 sg13g2_tiehi \ppu.copper_inst.store[12]$_DFFE_PP__482  (.L_HI(net482));
 sg13g2_tiehi \ppu.copper_inst.store[13]$_DFFE_PP__483  (.L_HI(net483));
 sg13g2_tiehi \ppu.copper_inst.store[14]$_DFFE_PP__484  (.L_HI(net484));
 sg13g2_tiehi \ppu.copper_inst.store[15]$_DFFE_PP__485  (.L_HI(net485));
 sg13g2_tiehi \ppu.copper_inst.store[1]$_DFFE_PP__486  (.L_HI(net486));
 sg13g2_tiehi \ppu.copper_inst.store[2]$_DFFE_PP__487  (.L_HI(net487));
 sg13g2_tiehi \ppu.copper_inst.store[3]$_DFFE_PP__488  (.L_HI(net488));
 sg13g2_tiehi \ppu.copper_inst.store[4]$_DFFE_PP__489  (.L_HI(net489));
 sg13g2_tiehi \ppu.copper_inst.store[5]$_DFFE_PP__490  (.L_HI(net490));
 sg13g2_tiehi \ppu.copper_inst.store[6]$_DFFE_PP__491  (.L_HI(net491));
 sg13g2_tiehi \ppu.copper_inst.store[7]$_DFFE_PP__492  (.L_HI(net492));
 sg13g2_tiehi \ppu.copper_inst.store[8]$_DFFE_PP__493  (.L_HI(net493));
 sg13g2_tiehi \ppu.copper_inst.store[9]$_DFFE_PP__494  (.L_HI(net494));
 sg13g2_tiehi \ppu.copper_inst.store_valid$_SDFFCE_PP0P__495  (.L_HI(net495));
 sg13g2_tiehi \ppu.curr_pal_addr[0]$_DFFE_PN__496  (.L_HI(net496));
 sg13g2_tiehi \ppu.curr_pal_addr[1]$_DFFE_PN__497  (.L_HI(net497));
 sg13g2_tiehi \ppu.curr_pal_addr[2]$_DFFE_PN__498  (.L_HI(net498));
 sg13g2_tiehi \ppu.curr_pal_addr[3]$_DFFE_PN__499  (.L_HI(net499));
 sg13g2_tiehi \ppu.display_mask[0]$_SDFFE_PN1P__500  (.L_HI(net500));
 sg13g2_tiehi \ppu.display_mask[1]$_SDFFE_PN1P__501  (.L_HI(net501));
 sg13g2_tiehi \ppu.display_mask[2]$_SDFFE_PN1P__502  (.L_HI(net502));
 sg13g2_tiehi \ppu.display_mask[3]$_SDFFE_PN1P__503  (.L_HI(net503));
 sg13g2_tiehi \ppu.display_mask[4]$_SDFFE_PN1P__504  (.L_HI(net504));
 sg13g2_tiehi \ppu.display_mask[5]$_SDFFE_PN1P__505  (.L_HI(net505));
 sg13g2_tiehi \ppu.gfxmode1[0]$_SDFFE_PN0P__506  (.L_HI(net506));
 sg13g2_tiehi \ppu.gfxmode1[1]$_SDFFE_PN0P__507  (.L_HI(net507));
 sg13g2_tiehi \ppu.gfxmode1[2]$_SDFFE_PN0P__508  (.L_HI(net508));
 sg13g2_tiehi \ppu.gfxmode1[3]$_SDFFE_PN1P__509  (.L_HI(net509));
 sg13g2_tiehi \ppu.gfxmode1[4]$_SDFFE_PN1P__510  (.L_HI(net510));
 sg13g2_tiehi \ppu.gfxmode1[5]$_SDFFE_PN1P__511  (.L_HI(net511));
 sg13g2_tiehi \ppu.gfxmode1[6]$_SDFFE_PN1P__512  (.L_HI(net512));
 sg13g2_tiehi \ppu.gfxmode1[7]$_SDFFE_PN0P__513  (.L_HI(net513));
 sg13g2_tiehi \ppu.gfxmode1[8]$_SDFFE_PN1P__514  (.L_HI(net514));
 sg13g2_tiehi \ppu.gfxmode2[0]$_SDFFE_PN0P__515  (.L_HI(net515));
 sg13g2_tiehi \ppu.gfxmode2[1]$_SDFFE_PN0P__516  (.L_HI(net516));
 sg13g2_tiehi \ppu.gfxmode2[2]$_SDFFE_PN0P__517  (.L_HI(net517));
 sg13g2_tiehi \ppu.gfxmode2[3]$_SDFFE_PN1P__518  (.L_HI(net518));
 sg13g2_tiehi \ppu.gfxmode2[4]$_SDFFE_PN0P__519  (.L_HI(net519));
 sg13g2_tiehi \ppu.gfxmode2[5]$_SDFFE_PN0P__520  (.L_HI(net520));
 sg13g2_tiehi \ppu.gfxmode2[6]$_SDFFE_PN0P__521  (.L_HI(net521));
 sg13g2_tiehi \ppu.gfxmode2[7]$_SDFFE_PN1P__522  (.L_HI(net522));
 sg13g2_tiehi \ppu.gfxmode2[8]$_SDFFE_PN1P__523  (.L_HI(net523));
 sg13g2_tiehi \ppu.gfxmode3[0]$_SDFFE_PN1P__524  (.L_HI(net524));
 sg13g2_tiehi \ppu.gfxmode3[1]$_SDFFE_PN1P__525  (.L_HI(net525));
 sg13g2_tiehi \ppu.gfxmode3[2]$_SDFFE_PN1P__526  (.L_HI(net526));
 sg13g2_tiehi \ppu.gfxmode3[3]$_SDFFE_PN1P__527  (.L_HI(net527));
 sg13g2_tiehi \ppu.gfxmode3[4]$_SDFFE_PN1P__528  (.L_HI(net528));
 sg13g2_tiehi \ppu.gfxmode3[5]$_SDFFE_PN1P__529  (.L_HI(net529));
 sg13g2_tiehi \ppu.gfxmode3[6]$_SDFFE_PN0P__530  (.L_HI(net530));
 sg13g2_tiehi \ppu.gfxmode3[7]$_SDFFE_PN1P__531  (.L_HI(net531));
 sg13g2_tiehi \ppu.gfxmode3[8]$_SDFFE_PN1P__532  (.L_HI(net532));
 sg13g2_tiehi \ppu.pal[0][0]$_DFFE_PN__533  (.L_HI(net533));
 sg13g2_tiehi \ppu.pal[0][1]$_DFFE_PN__534  (.L_HI(net534));
 sg13g2_tiehi \ppu.pal[0][2]$_DFFE_PN__535  (.L_HI(net535));
 sg13g2_tiehi \ppu.pal[0][3]$_DFFE_PN__536  (.L_HI(net536));
 sg13g2_tiehi \ppu.pal[0][4]$_DFFE_PN__537  (.L_HI(net537));
 sg13g2_tiehi \ppu.pal[0][5]$_DFFE_PN__538  (.L_HI(net538));
 sg13g2_tiehi \ppu.pal[0][6]$_DFFE_PN__539  (.L_HI(net539));
 sg13g2_tiehi \ppu.pal[0][7]$_DFFE_PN__540  (.L_HI(net540));
 sg13g2_tiehi \ppu.pal[10][0]$_DFFE_PN__541  (.L_HI(net541));
 sg13g2_tiehi \ppu.pal[10][1]$_DFFE_PN__542  (.L_HI(net542));
 sg13g2_tiehi \ppu.pal[10][2]$_DFFE_PN__543  (.L_HI(net543));
 sg13g2_tiehi \ppu.pal[10][3]$_DFFE_PN__544  (.L_HI(net544));
 sg13g2_tiehi \ppu.pal[10][4]$_DFFE_PN__545  (.L_HI(net545));
 sg13g2_tiehi \ppu.pal[10][5]$_DFFE_PN__546  (.L_HI(net546));
 sg13g2_tiehi \ppu.pal[10][6]$_DFFE_PN__547  (.L_HI(net547));
 sg13g2_tiehi \ppu.pal[10][7]$_DFFE_PN__548  (.L_HI(net548));
 sg13g2_tiehi \ppu.pal[11][0]$_DFFE_PN__549  (.L_HI(net549));
 sg13g2_tiehi \ppu.pal[11][1]$_DFFE_PN__550  (.L_HI(net550));
 sg13g2_tiehi \ppu.pal[11][2]$_DFFE_PN__551  (.L_HI(net551));
 sg13g2_tiehi \ppu.pal[11][3]$_DFFE_PN__552  (.L_HI(net552));
 sg13g2_tiehi \ppu.pal[11][4]$_DFFE_PN__553  (.L_HI(net553));
 sg13g2_tiehi \ppu.pal[11][5]$_DFFE_PN__554  (.L_HI(net554));
 sg13g2_tiehi \ppu.pal[11][6]$_DFFE_PN__555  (.L_HI(net555));
 sg13g2_tiehi \ppu.pal[11][7]$_DFFE_PN__556  (.L_HI(net556));
 sg13g2_tiehi \ppu.pal[12][0]$_DFFE_PN__557  (.L_HI(net557));
 sg13g2_tiehi \ppu.pal[12][1]$_DFFE_PN__558  (.L_HI(net558));
 sg13g2_tiehi \ppu.pal[12][2]$_DFFE_PN__559  (.L_HI(net559));
 sg13g2_tiehi \ppu.pal[12][3]$_DFFE_PN__560  (.L_HI(net560));
 sg13g2_tiehi \ppu.pal[12][4]$_DFFE_PN__561  (.L_HI(net561));
 sg13g2_tiehi \ppu.pal[12][5]$_DFFE_PN__562  (.L_HI(net562));
 sg13g2_tiehi \ppu.pal[12][6]$_DFFE_PN__563  (.L_HI(net563));
 sg13g2_tiehi \ppu.pal[12][7]$_DFFE_PN__564  (.L_HI(net564));
 sg13g2_tiehi \ppu.pal[13][0]$_DFFE_PN__565  (.L_HI(net565));
 sg13g2_tiehi \ppu.pal[13][1]$_DFFE_PN__566  (.L_HI(net566));
 sg13g2_tiehi \ppu.pal[13][2]$_DFFE_PN__567  (.L_HI(net567));
 sg13g2_tiehi \ppu.pal[13][3]$_DFFE_PN__568  (.L_HI(net568));
 sg13g2_tiehi \ppu.pal[13][4]$_DFFE_PN__569  (.L_HI(net569));
 sg13g2_tiehi \ppu.pal[13][5]$_DFFE_PN__570  (.L_HI(net570));
 sg13g2_tiehi \ppu.pal[13][6]$_DFFE_PN__571  (.L_HI(net571));
 sg13g2_tiehi \ppu.pal[13][7]$_DFFE_PN__572  (.L_HI(net572));
 sg13g2_tiehi \ppu.pal[14][0]$_DFFE_PN__573  (.L_HI(net573));
 sg13g2_tiehi \ppu.pal[14][1]$_DFFE_PN__574  (.L_HI(net574));
 sg13g2_tiehi \ppu.pal[14][2]$_DFFE_PN__575  (.L_HI(net575));
 sg13g2_tiehi \ppu.pal[14][3]$_DFFE_PN__576  (.L_HI(net576));
 sg13g2_tiehi \ppu.pal[14][4]$_DFFE_PN__577  (.L_HI(net577));
 sg13g2_tiehi \ppu.pal[14][5]$_DFFE_PN__578  (.L_HI(net578));
 sg13g2_tiehi \ppu.pal[14][6]$_DFFE_PN__579  (.L_HI(net579));
 sg13g2_tiehi \ppu.pal[14][7]$_DFFE_PN__580  (.L_HI(net580));
 sg13g2_tiehi \ppu.pal[15][0]$_DFFE_PN__581  (.L_HI(net581));
 sg13g2_tiehi \ppu.pal[15][1]$_DFFE_PN__582  (.L_HI(net582));
 sg13g2_tiehi \ppu.pal[15][2]$_DFFE_PN__583  (.L_HI(net583));
 sg13g2_tiehi \ppu.pal[15][3]$_DFFE_PN__584  (.L_HI(net584));
 sg13g2_tiehi \ppu.pal[15][4]$_DFFE_PN__585  (.L_HI(net585));
 sg13g2_tiehi \ppu.pal[15][5]$_DFFE_PN__586  (.L_HI(net586));
 sg13g2_tiehi \ppu.pal[15][6]$_DFFE_PN__587  (.L_HI(net587));
 sg13g2_tiehi \ppu.pal[15][7]$_DFFE_PN__588  (.L_HI(net588));
 sg13g2_tiehi \ppu.pal[1][0]$_DFFE_PN__589  (.L_HI(net589));
 sg13g2_tiehi \ppu.pal[1][1]$_DFFE_PN__590  (.L_HI(net590));
 sg13g2_tiehi \ppu.pal[1][2]$_DFFE_PN__591  (.L_HI(net591));
 sg13g2_tiehi \ppu.pal[1][3]$_DFFE_PN__592  (.L_HI(net592));
 sg13g2_tiehi \ppu.pal[1][4]$_DFFE_PN__593  (.L_HI(net593));
 sg13g2_tiehi \ppu.pal[1][5]$_DFFE_PN__594  (.L_HI(net594));
 sg13g2_tiehi \ppu.pal[1][6]$_DFFE_PN__595  (.L_HI(net595));
 sg13g2_tiehi \ppu.pal[1][7]$_DFFE_PN__596  (.L_HI(net596));
 sg13g2_tiehi \ppu.pal[2][0]$_DFFE_PN__597  (.L_HI(net597));
 sg13g2_tiehi \ppu.pal[2][1]$_DFFE_PN__598  (.L_HI(net598));
 sg13g2_tiehi \ppu.pal[2][2]$_DFFE_PN__599  (.L_HI(net599));
 sg13g2_tiehi \ppu.pal[2][3]$_DFFE_PN__600  (.L_HI(net600));
 sg13g2_tiehi \ppu.pal[2][4]$_DFFE_PN__601  (.L_HI(net601));
 sg13g2_tiehi \ppu.pal[2][5]$_DFFE_PN__602  (.L_HI(net602));
 sg13g2_tiehi \ppu.pal[2][6]$_DFFE_PN__603  (.L_HI(net603));
 sg13g2_tiehi \ppu.pal[2][7]$_DFFE_PN__604  (.L_HI(net604));
 sg13g2_tiehi \ppu.pal[3][0]$_DFFE_PN__605  (.L_HI(net605));
 sg13g2_tiehi \ppu.pal[3][1]$_DFFE_PN__606  (.L_HI(net606));
 sg13g2_tiehi \ppu.pal[3][2]$_DFFE_PN__607  (.L_HI(net607));
 sg13g2_tiehi \ppu.pal[3][3]$_DFFE_PN__608  (.L_HI(net608));
 sg13g2_tiehi \ppu.pal[3][4]$_DFFE_PN__609  (.L_HI(net609));
 sg13g2_tiehi \ppu.pal[3][5]$_DFFE_PN__610  (.L_HI(net610));
 sg13g2_tiehi \ppu.pal[3][6]$_DFFE_PN__611  (.L_HI(net611));
 sg13g2_tiehi \ppu.pal[3][7]$_DFFE_PN__612  (.L_HI(net612));
 sg13g2_tiehi \ppu.pal[4][0]$_DFFE_PN__613  (.L_HI(net613));
 sg13g2_tiehi \ppu.pal[4][1]$_DFFE_PN__614  (.L_HI(net614));
 sg13g2_tiehi \ppu.pal[4][2]$_DFFE_PN__615  (.L_HI(net615));
 sg13g2_tiehi \ppu.pal[4][3]$_DFFE_PN__616  (.L_HI(net616));
 sg13g2_tiehi \ppu.pal[4][4]$_DFFE_PN__617  (.L_HI(net617));
 sg13g2_tiehi \ppu.pal[4][5]$_DFFE_PN__618  (.L_HI(net618));
 sg13g2_tiehi \ppu.pal[4][6]$_DFFE_PN__619  (.L_HI(net619));
 sg13g2_tiehi \ppu.pal[4][7]$_DFFE_PN__620  (.L_HI(net620));
 sg13g2_tiehi \ppu.pal[5][0]$_DFFE_PN__621  (.L_HI(net621));
 sg13g2_tiehi \ppu.pal[5][1]$_DFFE_PN__622  (.L_HI(net622));
 sg13g2_tiehi \ppu.pal[5][2]$_DFFE_PN__623  (.L_HI(net623));
 sg13g2_tiehi \ppu.pal[5][3]$_DFFE_PN__624  (.L_HI(net624));
 sg13g2_tiehi \ppu.pal[5][4]$_DFFE_PN__625  (.L_HI(net625));
 sg13g2_tiehi \ppu.pal[5][5]$_DFFE_PN__626  (.L_HI(net626));
 sg13g2_tiehi \ppu.pal[5][6]$_DFFE_PN__627  (.L_HI(net627));
 sg13g2_tiehi \ppu.pal[5][7]$_DFFE_PN__628  (.L_HI(net628));
 sg13g2_tiehi \ppu.pal[6][0]$_DFFE_PN__629  (.L_HI(net629));
 sg13g2_tiehi \ppu.pal[6][1]$_DFFE_PN__630  (.L_HI(net630));
 sg13g2_tiehi \ppu.pal[6][2]$_DFFE_PN__631  (.L_HI(net631));
 sg13g2_tiehi \ppu.pal[6][3]$_DFFE_PN__632  (.L_HI(net632));
 sg13g2_tiehi \ppu.pal[6][4]$_DFFE_PN__633  (.L_HI(net633));
 sg13g2_tiehi \ppu.pal[6][5]$_DFFE_PN__634  (.L_HI(net634));
 sg13g2_tiehi \ppu.pal[6][6]$_DFFE_PN__635  (.L_HI(net635));
 sg13g2_tiehi \ppu.pal[6][7]$_DFFE_PN__636  (.L_HI(net636));
 sg13g2_tiehi \ppu.pal[7][0]$_DFFE_PN__637  (.L_HI(net637));
 sg13g2_tiehi \ppu.pal[7][1]$_DFFE_PN__638  (.L_HI(net638));
 sg13g2_tiehi \ppu.pal[7][2]$_DFFE_PN__639  (.L_HI(net639));
 sg13g2_tiehi \ppu.pal[7][3]$_DFFE_PN__640  (.L_HI(net640));
 sg13g2_tiehi \ppu.pal[7][4]$_DFFE_PN__641  (.L_HI(net641));
 sg13g2_tiehi \ppu.pal[7][5]$_DFFE_PN__642  (.L_HI(net642));
 sg13g2_tiehi \ppu.pal[7][6]$_DFFE_PN__643  (.L_HI(net643));
 sg13g2_tiehi \ppu.pal[7][7]$_DFFE_PN__644  (.L_HI(net644));
 sg13g2_tiehi \ppu.pal[8][0]$_DFFE_PN__645  (.L_HI(net645));
 sg13g2_tiehi \ppu.pal[8][1]$_DFFE_PN__646  (.L_HI(net646));
 sg13g2_tiehi \ppu.pal[8][2]$_DFFE_PN__647  (.L_HI(net647));
 sg13g2_tiehi \ppu.pal[8][3]$_DFFE_PN__648  (.L_HI(net648));
 sg13g2_tiehi \ppu.pal[8][4]$_DFFE_PN__649  (.L_HI(net649));
 sg13g2_tiehi \ppu.pal[8][5]$_DFFE_PN__650  (.L_HI(net650));
 sg13g2_tiehi \ppu.pal[8][6]$_DFFE_PN__651  (.L_HI(net651));
 sg13g2_tiehi \ppu.pal[8][7]$_DFFE_PN__652  (.L_HI(net652));
 sg13g2_tiehi \ppu.pal[9][0]$_DFFE_PN__653  (.L_HI(net653));
 sg13g2_tiehi \ppu.pal[9][1]$_DFFE_PN__654  (.L_HI(net654));
 sg13g2_tiehi \ppu.pal[9][2]$_DFFE_PN__655  (.L_HI(net655));
 sg13g2_tiehi \ppu.pal[9][3]$_DFFE_PN__656  (.L_HI(net656));
 sg13g2_tiehi \ppu.pal[9][4]$_DFFE_PN__657  (.L_HI(net657));
 sg13g2_tiehi \ppu.pal[9][5]$_DFFE_PN__658  (.L_HI(net658));
 sg13g2_tiehi \ppu.pal[9][6]$_DFFE_PN__659  (.L_HI(net659));
 sg13g2_tiehi \ppu.pal[9][7]$_DFFE_PN__660  (.L_HI(net660));
 sg13g2_tiehi \ppu.pal_temp[4]$_DFF_P__661  (.L_HI(net661));
 sg13g2_tiehi \ppu.pal_temp[5]$_DFF_P__662  (.L_HI(net662));
 sg13g2_tiehi \ppu.pal_temp[6]$_DFF_P__663  (.L_HI(net663));
 sg13g2_tiehi \ppu.pal_temp[7]$_DFF_P__664  (.L_HI(net664));
 sg13g2_tiehi \ppu.ram_on$_SDFFE_PN0N__665  (.L_HI(net665));
 sg13g2_tiehi \ppu.ram_running$_SDFFE_PN0N__666  (.L_HI(net666));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[0]$_DFFE_PP__667  (.L_HI(net667));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[10]$_SDFFCE_PN0P__668  (.L_HI(net668));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[11]$_SDFFCE_PN0P__669  (.L_HI(net669));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[1]$_DFFE_PP__670  (.L_HI(net670));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[2]$_DFFE_PP__671  (.L_HI(net671));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[3]$_DFFE_PP__672  (.L_HI(net672));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[4]$_DFFE_PP__673  (.L_HI(net673));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[5]$_DFFE_PP__674  (.L_HI(net674));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[6]$_DFFE_PP__675  (.L_HI(net675));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[7]$_DFFE_PP__676  (.L_HI(net676));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[8]$_DFFE_PP__677  (.L_HI(net677));
 sg13g2_tiehi \ppu.rcoord.levels_sreg[9]$_SDFFCE_PN0P__678  (.L_HI(net678));
 sg13g2_tiehi \ppu.rgb_out_reg[10]$_DFFE_PN__679  (.L_HI(net679));
 sg13g2_tiehi \ppu.rgb_out_reg[11]$_DFFE_PN__680  (.L_HI(net680));
 sg13g2_tiehi \ppu.rgb_out_reg[2]$_DFFE_PN__681  (.L_HI(net681));
 sg13g2_tiehi \ppu.rgb_out_reg[3]$_DFFE_PN__682  (.L_HI(net682));
 sg13g2_tiehi \ppu.rgb_out_reg[5]$_DFFE_PN__683  (.L_HI(net683));
 sg13g2_tiehi \ppu.rgb_out_reg[6]$_DFFE_PN__684  (.L_HI(net684));
 sg13g2_tiehi \ppu.rgb_out_reg[7]$_DFFE_PN__685  (.L_HI(net685));
 sg13g2_tiehi \ppu.rgb_out_reg[9]$_DFFE_PN__686  (.L_HI(net686));
 sg13g2_tiehi \ppu.rs2.vsync0$_SDFFE_PN0P__687  (.L_HI(net687));
 sg13g2_tiehi \ppu.rs2.x_scan.counter[0]$_DFF_P__688  (.L_HI(net688));
 sg13g2_tiehi \ppu.rs2.x_scan.counter[1]$_DFF_P__689  (.L_HI(net689));
 sg13g2_tiehi \ppu.rs2.x_scan.counter[2]$_DFF_P__690  (.L_HI(net690));
 sg13g2_tiehi \ppu.rs2.x_scan.counter[3]$_SDFF_PN1__691  (.L_HI(net691));
 sg13g2_tiehi \ppu.rs2.x_scan.counter[4]$_SDFF_PN1__692  (.L_HI(net692));
 sg13g2_tiehi \ppu.rs2.x_scan.counter[5]$_SDFF_PP1__693  (.L_HI(net693));
 sg13g2_tiehi \ppu.rs2.x_scan.counter[6]$_SDFF_PP1__694  (.L_HI(net694));
 sg13g2_tiehi \ppu.rs2.x_scan.counter[7]$_SDFF_PP0__695  (.L_HI(net695));
 sg13g2_tiehi \ppu.rs2.x_scan.counter[8]$_SDFF_PP0__696  (.L_HI(net696));
 sg13g2_tiehi \ppu.rs2.x_scan.phase$_SDFFE_PN0P__697  (.L_HI(net697));
 sg13g2_tiehi \ppu.rs2.y_scan.counter[0]$_SDFFE_PN0P__698  (.L_HI(net698));
 sg13g2_tiehi \ppu.rs2.y_scan.counter[1]$_SDFFE_PN0P__699  (.L_HI(net699));
 sg13g2_tiehi \ppu.rs2.y_scan.counter[2]$_SDFFE_PN0P__700  (.L_HI(net700));
 sg13g2_tiehi \ppu.rs2.y_scan.counter[3]$_SDFFE_PN0P__701  (.L_HI(net701));
 sg13g2_tiehi \ppu.rs2.y_scan.counter[4]$_SDFFE_PN0P__702  (.L_HI(net702));
 sg13g2_tiehi \ppu.rs2.y_scan.counter[5]$_SDFFE_PN0P__703  (.L_HI(net703));
 sg13g2_tiehi \ppu.rs2.y_scan.counter[6]$_SDFFE_PN0P__704  (.L_HI(net704));
 sg13g2_tiehi \ppu.rs2.y_scan.counter[7]$_SDFFE_PN0P__705  (.L_HI(net705));
 sg13g2_tiehi \ppu.rs2.y_scan.counter[8]$_SDFFE_PN0P__706  (.L_HI(net706));
 sg13g2_tiehi \ppu.rs2.y_scan.phase[0]$_SDFFE_PN0P__707  (.L_HI(net707));
 sg13g2_tiehi \ppu.rs2.y_scan.phase[1]$_SDFFE_PN1P__708  (.L_HI(net708));
 sg13g2_tiehi \ppu.scroll_regs[0][0]$_DFFE_PP__709  (.L_HI(net709));
 sg13g2_tiehi \ppu.scroll_regs[0][1]$_DFFE_PP__710  (.L_HI(net710));
 sg13g2_tiehi \ppu.scroll_regs[0][2]$_DFFE_PP__711  (.L_HI(net711));
 sg13g2_tiehi \ppu.scroll_regs[0][3]$_DFFE_PP__712  (.L_HI(net712));
 sg13g2_tiehi \ppu.scroll_regs[0][4]$_DFFE_PP__713  (.L_HI(net713));
 sg13g2_tiehi \ppu.scroll_regs[0][5]$_DFFE_PP__714  (.L_HI(net714));
 sg13g2_tiehi \ppu.scroll_regs[0][6]$_DFFE_PP__715  (.L_HI(net715));
 sg13g2_tiehi \ppu.scroll_regs[0][7]$_DFFE_PP__716  (.L_HI(net716));
 sg13g2_tiehi \ppu.scroll_regs[0][8]$_DFFE_PP__717  (.L_HI(net717));
 sg13g2_tiehi \ppu.scroll_regs[1][0]$_DFFE_PP__718  (.L_HI(net718));
 sg13g2_tiehi \ppu.scroll_regs[1][1]$_DFFE_PP__719  (.L_HI(net719));
 sg13g2_tiehi \ppu.scroll_regs[1][2]$_DFFE_PP__720  (.L_HI(net720));
 sg13g2_tiehi \ppu.scroll_regs[1][3]$_DFFE_PP__721  (.L_HI(net721));
 sg13g2_tiehi \ppu.scroll_regs[1][4]$_DFFE_PP__722  (.L_HI(net722));
 sg13g2_tiehi \ppu.scroll_regs[1][5]$_DFFE_PP__723  (.L_HI(net723));
 sg13g2_tiehi \ppu.scroll_regs[1][6]$_DFFE_PP__724  (.L_HI(net724));
 sg13g2_tiehi \ppu.scroll_regs[1][7]$_DFFE_PP__725  (.L_HI(net725));
 sg13g2_tiehi \ppu.scroll_regs[1][8]$_DFFE_PP__726  (.L_HI(net726));
 sg13g2_tiehi \ppu.scroll_regs[2][0]$_DFFE_PP__727  (.L_HI(net727));
 sg13g2_tiehi \ppu.scroll_regs[2][1]$_DFFE_PP__728  (.L_HI(net728));
 sg13g2_tiehi \ppu.scroll_regs[2][2]$_DFFE_PP__729  (.L_HI(net729));
 sg13g2_tiehi \ppu.scroll_regs[2][3]$_DFFE_PP__730  (.L_HI(net730));
 sg13g2_tiehi \ppu.scroll_regs[2][4]$_DFFE_PP__731  (.L_HI(net731));
 sg13g2_tiehi \ppu.scroll_regs[2][5]$_DFFE_PP__732  (.L_HI(net732));
 sg13g2_tiehi \ppu.scroll_regs[2][6]$_DFFE_PP__733  (.L_HI(net733));
 sg13g2_tiehi \ppu.scroll_regs[2][7]$_DFFE_PP__734  (.L_HI(net734));
 sg13g2_tiehi \ppu.scroll_regs[2][8]$_DFFE_PP__735  (.L_HI(net735));
 sg13g2_tiehi \ppu.scroll_regs[3][0]$_DFFE_PP__736  (.L_HI(net736));
 sg13g2_tiehi \ppu.scroll_regs[3][1]$_DFFE_PP__737  (.L_HI(net737));
 sg13g2_tiehi \ppu.scroll_regs[3][2]$_DFFE_PP__738  (.L_HI(net738));
 sg13g2_tiehi \ppu.scroll_regs[3][3]$_DFFE_PP__739  (.L_HI(net739));
 sg13g2_tiehi \ppu.scroll_regs[3][4]$_DFFE_PP__740  (.L_HI(net740));
 sg13g2_tiehi \ppu.scroll_regs[3][5]$_DFFE_PP__741  (.L_HI(net741));
 sg13g2_tiehi \ppu.scroll_regs[3][6]$_DFFE_PP__742  (.L_HI(net742));
 sg13g2_tiehi \ppu.scroll_regs[3][7]$_DFFE_PP__743  (.L_HI(net743));
 sg13g2_tiehi \ppu.scroll_regs[3][8]$_DFFE_PP__744  (.L_HI(net744));
 sg13g2_tiehi \ppu.serial_counter[0]$_SDFF_PN0__745  (.L_HI(net745));
 sg13g2_tiehi \ppu.serial_counter[1]$_SDFF_PN0__746  (.L_HI(net746));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][0]$_DFFE_PP__747  (.L_HI(net747));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][10]$_DFFE_PP__748  (.L_HI(net748));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][11]$_DFFE_PP__749  (.L_HI(net749));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][12]$_DFFE_PP__750  (.L_HI(net750));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][13]$_DFFE_PP__751  (.L_HI(net751));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][14]$_DFFE_PP__752  (.L_HI(net752));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][15]$_DFFE_PP__753  (.L_HI(net753));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][1]$_DFFE_PP__754  (.L_HI(net754));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][2]$_DFFE_PP__755  (.L_HI(net755));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][3]$_DFFE_PP__756  (.L_HI(net756));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][4]$_DFFE_PP__757  (.L_HI(net757));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][5]$_DFFE_PP__758  (.L_HI(net758));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][6]$_DFFE_PP__759  (.L_HI(net759));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][7]$_DFFE_PP__760  (.L_HI(net760));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][8]$_DFFE_PP__761  (.L_HI(net761));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[0][9]$_DFFE_PP__762  (.L_HI(net762));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][0]$_DFFE_PP__763  (.L_HI(net763));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][10]$_DFFE_PP__764  (.L_HI(net764));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][11]$_DFFE_PP__765  (.L_HI(net765));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][12]$_DFFE_PP__766  (.L_HI(net766));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][13]$_DFFE_PP__767  (.L_HI(net767));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][14]$_DFFE_PP__768  (.L_HI(net768));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][15]$_DFFE_PP__769  (.L_HI(net769));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][1]$_DFFE_PP__770  (.L_HI(net770));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][2]$_DFFE_PP__771  (.L_HI(net771));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][3]$_DFFE_PP__772  (.L_HI(net772));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][4]$_DFFE_PP__773  (.L_HI(net773));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][5]$_DFFE_PP__774  (.L_HI(net774));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][6]$_DFFE_PP__775  (.L_HI(net775));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][7]$_DFFE_PP__776  (.L_HI(net776));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][8]$_DFFE_PP__777  (.L_HI(net777));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[1][9]$_DFFE_PP__778  (.L_HI(net778));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][0]$_DFFE_PP__779  (.L_HI(net779));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][10]$_DFFE_PP__780  (.L_HI(net780));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][11]$_DFFE_PP__781  (.L_HI(net781));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][12]$_DFFE_PP__782  (.L_HI(net782));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][13]$_DFFE_PP__783  (.L_HI(net783));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][14]$_DFFE_PP__784  (.L_HI(net784));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][15]$_DFFE_PP__785  (.L_HI(net785));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][1]$_DFFE_PP__786  (.L_HI(net786));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][2]$_DFFE_PP__787  (.L_HI(net787));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][3]$_DFFE_PP__788  (.L_HI(net788));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][4]$_DFFE_PP__789  (.L_HI(net789));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][5]$_DFFE_PP__790  (.L_HI(net790));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][6]$_DFFE_PP__791  (.L_HI(net791));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][7]$_DFFE_PP__792  (.L_HI(net792));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][8]$_DFFE_PP__793  (.L_HI(net793));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[2][9]$_DFFE_PP__794  (.L_HI(net794));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][0]$_DFFE_PP__795  (.L_HI(net795));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][10]$_DFFE_PP__796  (.L_HI(net796));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][11]$_DFFE_PP__797  (.L_HI(net797));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][12]$_DFFE_PP__798  (.L_HI(net798));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][13]$_DFFE_PP__799  (.L_HI(net799));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][14]$_DFFE_PP__800  (.L_HI(net800));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][15]$_DFFE_PP__801  (.L_HI(net801));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][1]$_DFFE_PP__802  (.L_HI(net802));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][2]$_DFFE_PP__803  (.L_HI(net803));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][3]$_DFFE_PP__804  (.L_HI(net804));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][4]$_DFFE_PP__805  (.L_HI(net805));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][5]$_DFFE_PP__806  (.L_HI(net806));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][6]$_DFFE_PP__807  (.L_HI(net807));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][7]$_DFFE_PP__808  (.L_HI(net808));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][8]$_DFFE_PP__809  (.L_HI(net809));
 sg13g2_tiehi \ppu.sprite_buffer.attr_x[3][9]$_DFFE_PP__810  (.L_HI(net810));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][0]$_DFFE_PP__811  (.L_HI(net811));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][10]$_DFFE_PP__812  (.L_HI(net812));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][11]$_DFFE_PP__813  (.L_HI(net813));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][12]$_DFFE_PP__814  (.L_HI(net814));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][13]$_DFFE_PP__815  (.L_HI(net815));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][14]$_DFFE_PP__816  (.L_HI(net816));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][15]$_DFFE_PP__817  (.L_HI(net817));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][1]$_DFFE_PP__818  (.L_HI(net818));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][2]$_DFFE_PP__819  (.L_HI(net819));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][4]$_DFFE_PP__820  (.L_HI(net820));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][5]$_DFFE_PP__821  (.L_HI(net821));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][6]$_DFFE_PP__822  (.L_HI(net822));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][7]$_DFFE_PP__823  (.L_HI(net823));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][8]$_DFFE_PP__824  (.L_HI(net824));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[0][9]$_DFFE_PP__825  (.L_HI(net825));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][0]$_DFFE_PP__826  (.L_HI(net826));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][10]$_DFFE_PP__827  (.L_HI(net827));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][11]$_DFFE_PP__828  (.L_HI(net828));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][12]$_DFFE_PP__829  (.L_HI(net829));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][13]$_DFFE_PP__830  (.L_HI(net830));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][14]$_DFFE_PP__831  (.L_HI(net831));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][15]$_DFFE_PP__832  (.L_HI(net832));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][1]$_DFFE_PP__833  (.L_HI(net833));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][2]$_DFFE_PP__834  (.L_HI(net834));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][4]$_DFFE_PP__835  (.L_HI(net835));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][5]$_DFFE_PP__836  (.L_HI(net836));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][6]$_DFFE_PP__837  (.L_HI(net837));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][7]$_DFFE_PP__838  (.L_HI(net838));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][8]$_DFFE_PP__839  (.L_HI(net839));
 sg13g2_tiehi \ppu.sprite_buffer.attr_y[1][9]$_DFFE_PP__840  (.L_HI(net840));
 sg13g2_tiehi \ppu.sprite_buffer.extra_sorted_addr_bits[0]$_SDFF_PP0__841  (.L_HI(net841));
 sg13g2_tiehi \ppu.sprite_buffer.extra_sorted_addr_bits[1]$_SDFF_PP0__842  (.L_HI(net842));
 sg13g2_tiehi \ppu.sprite_buffer.extra_sorted_addr_bits[2]$_SDFF_PP0__843  (.L_HI(net843));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[0][0]$_DFFE_PP__844  (.L_HI(net844));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[0][1]$_DFFE_PP__845  (.L_HI(net845));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[0][2]$_DFFE_PP__846  (.L_HI(net846));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[0][3]$_DFFE_PP__847  (.L_HI(net847));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[0][4]$_DFFE_PP__848  (.L_HI(net848));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[0][5]$_DFFE_PP__849  (.L_HI(net849));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[1][0]$_DFFE_PP__850  (.L_HI(net850));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[1][1]$_DFFE_PP__851  (.L_HI(net851));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[1][2]$_DFFE_PP__852  (.L_HI(net852));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[1][3]$_DFFE_PP__853  (.L_HI(net853));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[1][4]$_DFFE_PP__854  (.L_HI(net854));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[1][5]$_DFFE_PP__855  (.L_HI(net855));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[2][0]$_DFFE_PP__856  (.L_HI(net856));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[2][1]$_DFFE_PP__857  (.L_HI(net857));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[2][2]$_DFFE_PP__858  (.L_HI(net858));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[2][3]$_DFFE_PP__859  (.L_HI(net859));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[2][4]$_DFFE_PP__860  (.L_HI(net860));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[2][5]$_DFFE_PP__861  (.L_HI(net861));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[3][0]$_DFFE_PP__862  (.L_HI(net862));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[3][1]$_DFFE_PP__863  (.L_HI(net863));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[3][2]$_DFFE_PP__864  (.L_HI(net864));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[3][3]$_DFFE_PP__865  (.L_HI(net865));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[3][4]$_DFFE_PP__866  (.L_HI(net866));
 sg13g2_tiehi \ppu.sprite_buffer.id_buffer[3][5]$_DFFE_PP__867  (.L_HI(net867));
 sg13g2_tiehi \ppu.sprite_buffer.in_counters[0][0]$_SDFF_PP0__868  (.L_HI(net868));
 sg13g2_tiehi \ppu.sprite_buffer.in_counters[0][1]$_SDFF_PP0__869  (.L_HI(net869));
 sg13g2_tiehi \ppu.sprite_buffer.in_counters[1][0]$_SDFF_PP0__870  (.L_HI(net870));
 sg13g2_tiehi \ppu.sprite_buffer.in_counters[1][1]$_SDFF_PP0__871  (.L_HI(net871));
 sg13g2_tiehi \ppu.sprite_buffer.in_counters[1][2]$_SDFF_PP0__872  (.L_HI(net872));
 sg13g2_tiehi \ppu.sprite_buffer.in_counters[2][0]$_SDFF_PP0__873  (.L_HI(net873));
 sg13g2_tiehi \ppu.sprite_buffer.in_counters[2][1]$_SDFF_PP0__874  (.L_HI(net874));
 sg13g2_tiehi \ppu.sprite_buffer.in_counters[2][2]$_SDFF_PP0__875  (.L_HI(net875));
 sg13g2_tiehi \ppu.sprite_buffer.last_data_pins[0]$_DFF_P__876  (.L_HI(net876));
 sg13g2_tiehi \ppu.sprite_buffer.last_data_pins[1]$_DFF_P__877  (.L_HI(net877));
 sg13g2_tiehi \ppu.sprite_buffer.last_data_pins[2]$_DFF_P__878  (.L_HI(net878));
 sg13g2_tiehi \ppu.sprite_buffer.last_data_pins[3]$_DFF_P__879  (.L_HI(net879));
 sg13g2_tiehi \ppu.sprite_buffer.oam_load_sprite_valid$_DFFE_PN__880  (.L_HI(net880));
 sg13g2_tiehi \ppu.sprite_buffer.oam_req_step$_SDFFE_PP0P__881  (.L_HI(net881));
 sg13g2_tiehi \ppu.sprite_buffer.out_counters[0][0]$_SDFF_PP0__882  (.L_HI(net882));
 sg13g2_tiehi \ppu.sprite_buffer.out_counters[0][1]$_SDFF_PP0__883  (.L_HI(net883));
 sg13g2_tiehi \ppu.sprite_buffer.out_counters[0][2]$_SDFF_PP0__884  (.L_HI(net884));
 sg13g2_tiehi \ppu.sprite_buffer.out_counters[1][0]$_SDFF_PP0__885  (.L_HI(net885));
 sg13g2_tiehi \ppu.sprite_buffer.out_counters[1][1]$_SDFF_PP0__886  (.L_HI(net886));
 sg13g2_tiehi \ppu.sprite_buffer.out_counters[2][0]$_SDFF_PP0__887  (.L_HI(net887));
 sg13g2_tiehi \ppu.sprite_buffer.out_counters[2][1]$_SDFF_PP0__888  (.L_HI(net888));
 sg13g2_tiehi \ppu.sprite_buffer.out_counters[2][2]$_SDFF_PP0__889  (.L_HI(net889));
 sg13g2_tiehi \ppu.sprite_buffer.scan_enabled$_DFFE_PP__890  (.L_HI(net890));
 sg13g2_tiehi \ppu.sprite_buffer.scan_on$_DFF_P__891  (.L_HI(net891));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[0][0]$_DFF_P__892  (.L_HI(net892));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[0][1]$_DFF_P__893  (.L_HI(net893));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[0][2]$_DFF_P__894  (.L_HI(net894));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[1][0]$_DFF_P__895  (.L_HI(net895));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[1][1]$_DFF_P__896  (.L_HI(net896));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[1][2]$_DFF_P__897  (.L_HI(net897));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[2][0]$_DFF_P__898  (.L_HI(net898));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[2][1]$_DFF_P__899  (.L_HI(net899));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[2][2]$_DFF_P__900  (.L_HI(net900));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[3][0]$_DFF_P__901  (.L_HI(net901));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[3][1]$_DFF_P__902  (.L_HI(net902));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_catch_up_counters[3][2]$_DFF_P__903  (.L_HI(net903));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[0][0]$_DFFE_PP__904  (.L_HI(net904));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[0][1]$_DFFE_PP__905  (.L_HI(net905));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[0][2]$_DFFE_PP__906  (.L_HI(net906));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[0][3]$_DFFE_PP__907  (.L_HI(net907));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[0][4]$_DFFE_PP__908  (.L_HI(net908));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[0][5]$_DFFE_PP__909  (.L_HI(net909));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[1][0]$_DFFE_PP__910  (.L_HI(net910));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[1][1]$_DFFE_PP__911  (.L_HI(net911));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[1][2]$_DFFE_PP__912  (.L_HI(net912));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[1][3]$_DFFE_PP__913  (.L_HI(net913));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[1][4]$_DFFE_PP__914  (.L_HI(net914));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[1][5]$_DFFE_PP__915  (.L_HI(net915));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[2][0]$_DFFE_PP__916  (.L_HI(net916));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[2][1]$_DFFE_PP__917  (.L_HI(net917));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[2][2]$_DFFE_PP__918  (.L_HI(net918));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[2][3]$_DFFE_PP__919  (.L_HI(net919));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[2][4]$_DFFE_PP__920  (.L_HI(net920));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[2][5]$_DFFE_PP__921  (.L_HI(net921));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[3][0]$_DFFE_PP__922  (.L_HI(net922));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[3][1]$_DFFE_PP__923  (.L_HI(net923));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[3][2]$_DFFE_PP__924  (.L_HI(net924));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[3][3]$_DFFE_PP__925  (.L_HI(net925));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[3][4]$_DFFE_PP__926  (.L_HI(net926));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_ids[3][5]$_DFFE_PP__927  (.L_HI(net927));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_out_color[0]$_DFFE_PP__928  (.L_HI(net928));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_out_color[1]$_DFFE_PP__929  (.L_HI(net929));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_out_color[2]$_DFFE_PP__930  (.L_HI(net930));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_out_color[3]$_DFFE_PP__931  (.L_HI(net931));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_out_depth[0]$_DFFE_PP__932  (.L_HI(net932));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_out_depth[1]$_DFFE_PP__933  (.L_HI(net933));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][0]$_DFFE_PP__934  (.L_HI(net934));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][10]$_DFFE_PP__935  (.L_HI(net935));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][11]$_DFFE_PP__936  (.L_HI(net936));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][12]$_DFFE_PP__937  (.L_HI(net937));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][13]$_DFFE_PP__938  (.L_HI(net938));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][14]$_DFFE_PP__939  (.L_HI(net939));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][15]$_DFFE_PP__940  (.L_HI(net940));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][16]$_DFFE_PP__941  (.L_HI(net941));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][17]$_DFFE_PP__942  (.L_HI(net942));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][18]$_DFFE_PP__943  (.L_HI(net943));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][19]$_DFFE_PP__944  (.L_HI(net944));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][1]$_DFFE_PP__945  (.L_HI(net945));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][20]$_DFFE_PP__946  (.L_HI(net946));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][21]$_DFFE_PP__947  (.L_HI(net947));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][22]$_DFFE_PP__948  (.L_HI(net948));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][23]$_DFFE_PP__949  (.L_HI(net949));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][24]$_DFFE_PP__950  (.L_HI(net950));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][25]$_DFFE_PP__951  (.L_HI(net951));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][26]$_DFFE_PP__952  (.L_HI(net952));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][27]$_DFFE_PP__953  (.L_HI(net953));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][28]$_DFFE_PP__954  (.L_HI(net954));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][29]$_DFFE_PP__955  (.L_HI(net955));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][2]$_DFFE_PP__956  (.L_HI(net956));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][30]$_DFFE_PP__957  (.L_HI(net957));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][31]$_DFFE_PP__958  (.L_HI(net958));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][3]$_DFFE_PP__959  (.L_HI(net959));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][4]$_DFFE_PP__960  (.L_HI(net960));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][5]$_DFFE_PP__961  (.L_HI(net961));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][6]$_DFFE_PP__962  (.L_HI(net962));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][7]$_DFFE_PP__963  (.L_HI(net963));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][8]$_DFFE_PP__964  (.L_HI(net964));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[0][9]$_DFFE_PP__965  (.L_HI(net965));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][0]$_DFFE_PP__966  (.L_HI(net966));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][10]$_DFFE_PP__967  (.L_HI(net967));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][11]$_DFFE_PP__968  (.L_HI(net968));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][12]$_DFFE_PP__969  (.L_HI(net969));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][13]$_DFFE_PP__970  (.L_HI(net970));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][14]$_DFFE_PP__971  (.L_HI(net971));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][15]$_DFFE_PP__972  (.L_HI(net972));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][16]$_DFFE_PP__973  (.L_HI(net973));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][17]$_DFFE_PP__974  (.L_HI(net974));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][18]$_DFFE_PP__975  (.L_HI(net975));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][19]$_DFFE_PP__976  (.L_HI(net976));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][1]$_DFFE_PP__977  (.L_HI(net977));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][20]$_DFFE_PP__978  (.L_HI(net978));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][21]$_DFFE_PP__979  (.L_HI(net979));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][22]$_DFFE_PP__980  (.L_HI(net980));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][23]$_DFFE_PP__981  (.L_HI(net981));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][24]$_DFFE_PP__982  (.L_HI(net982));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][25]$_DFFE_PP__983  (.L_HI(net983));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][26]$_DFFE_PP__984  (.L_HI(net984));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][27]$_DFFE_PP__985  (.L_HI(net985));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][28]$_DFFE_PP__986  (.L_HI(net986));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][29]$_DFFE_PP__987  (.L_HI(net987));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][2]$_DFFE_PP__988  (.L_HI(net988));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][30]$_DFFE_PP__989  (.L_HI(net989));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][31]$_DFFE_PP__990  (.L_HI(net990));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][3]$_DFFE_PP__991  (.L_HI(net991));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][4]$_DFFE_PP__992  (.L_HI(net992));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][5]$_DFFE_PP__993  (.L_HI(net993));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][6]$_DFFE_PP__994  (.L_HI(net994));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][7]$_DFFE_PP__995  (.L_HI(net995));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][8]$_DFFE_PP__996  (.L_HI(net996));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[1][9]$_DFFE_PP__997  (.L_HI(net997));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][0]$_DFFE_PP__998  (.L_HI(net998));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][10]$_DFFE_PP__999  (.L_HI(net999));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][11]$_DFFE_PP__1000  (.L_HI(net1000));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][12]$_DFFE_PP__1001  (.L_HI(net1001));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][13]$_DFFE_PP__1002  (.L_HI(net1002));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][14]$_DFFE_PP__1003  (.L_HI(net1003));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][15]$_DFFE_PP__1004  (.L_HI(net1004));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][16]$_DFFE_PP__1005  (.L_HI(net1005));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][17]$_DFFE_PP__1006  (.L_HI(net1006));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][18]$_DFFE_PP__1007  (.L_HI(net1007));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][19]$_DFFE_PP__1008  (.L_HI(net1008));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][1]$_DFFE_PP__1009  (.L_HI(net1009));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][20]$_DFFE_PP__1010  (.L_HI(net1010));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][21]$_DFFE_PP__1011  (.L_HI(net1011));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][22]$_DFFE_PP__1012  (.L_HI(net1012));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][23]$_DFFE_PP__1013  (.L_HI(net1013));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][24]$_DFFE_PP__1014  (.L_HI(net1014));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][25]$_DFFE_PP__1015  (.L_HI(net1015));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][26]$_DFFE_PP__1016  (.L_HI(net1016));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][27]$_DFFE_PP__1017  (.L_HI(net1017));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][28]$_DFFE_PP__1018  (.L_HI(net1018));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][29]$_DFFE_PP__1019  (.L_HI(net1019));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][2]$_DFFE_PP__1020  (.L_HI(net1020));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][30]$_DFFE_PP__1021  (.L_HI(net1021));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][31]$_DFFE_PP__1022  (.L_HI(net1022));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][3]$_DFFE_PP__1023  (.L_HI(net1023));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][4]$_DFFE_PP__1024  (.L_HI(net1024));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][5]$_DFFE_PP__1025  (.L_HI(net1025));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][6]$_DFFE_PP__1026  (.L_HI(net1026));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][7]$_DFFE_PP__1027  (.L_HI(net1027));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][8]$_DFFE_PP__1028  (.L_HI(net1028));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[2][9]$_DFFE_PP__1029  (.L_HI(net1029));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][0]$_DFFE_PP__1030  (.L_HI(net1030));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][10]$_DFFE_PP__1031  (.L_HI(net1031));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][11]$_DFFE_PP__1032  (.L_HI(net1032));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][12]$_DFFE_PP__1033  (.L_HI(net1033));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][13]$_DFFE_PP__1034  (.L_HI(net1034));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][14]$_DFFE_PP__1035  (.L_HI(net1035));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][15]$_DFFE_PP__1036  (.L_HI(net1036));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][16]$_DFFE_PP__1037  (.L_HI(net1037));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][17]$_DFFE_PP__1038  (.L_HI(net1038));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][18]$_DFFE_PP__1039  (.L_HI(net1039));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][19]$_DFFE_PP__1040  (.L_HI(net1040));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][1]$_DFFE_PP__1041  (.L_HI(net1041));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][20]$_DFFE_PP__1042  (.L_HI(net1042));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][21]$_DFFE_PP__1043  (.L_HI(net1043));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][22]$_DFFE_PP__1044  (.L_HI(net1044));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][23]$_DFFE_PP__1045  (.L_HI(net1045));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][24]$_DFFE_PP__1046  (.L_HI(net1046));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][25]$_DFFE_PP__1047  (.L_HI(net1047));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][26]$_DFFE_PP__1048  (.L_HI(net1048));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][27]$_DFFE_PP__1049  (.L_HI(net1049));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][28]$_DFFE_PP__1050  (.L_HI(net1050));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][29]$_DFFE_PP__1051  (.L_HI(net1051));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][2]$_DFFE_PP__1052  (.L_HI(net1052));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][30]$_DFFE_PP__1053  (.L_HI(net1053));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][31]$_DFFE_PP__1054  (.L_HI(net1054));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][3]$_DFFE_PP__1055  (.L_HI(net1055));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][4]$_DFFE_PP__1056  (.L_HI(net1056));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][5]$_DFFE_PP__1057  (.L_HI(net1057));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][6]$_DFFE_PP__1058  (.L_HI(net1058));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][7]$_DFFE_PP__1059  (.L_HI(net1059));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][8]$_DFFE_PP__1060  (.L_HI(net1060));
 sg13g2_tiehi \ppu.sprite_buffer.sprite_pixels[3][9]$_DFFE_PP__1061  (.L_HI(net1061));
 sg13g2_tiehi \ppu.sprite_buffer.top_color[0]$_SDFFCE_PN0P__1062  (.L_HI(net1062));
 sg13g2_tiehi \ppu.sprite_buffer.top_color[1]$_SDFFCE_PN0P__1063  (.L_HI(net1063));
 sg13g2_tiehi \ppu.sprite_buffer.top_color[2]$_SDFFCE_PN0P__1064  (.L_HI(net1064));
 sg13g2_tiehi \ppu.sprite_buffer.top_color[3]$_SDFFCE_PN0P__1065  (.L_HI(net1065));
 sg13g2_tiehi \ppu.sprite_buffer.top_depth[0]$_SDFFCE_PN1P__1066  (.L_HI(net1066));
 sg13g2_tiehi \ppu.sprite_buffer.top_depth[1]$_SDFFCE_PN1P__1067  (.L_HI(net1067));
 sg13g2_tiehi \ppu.sprite_buffer.top_prio[0]$_DFFE_PP__1068  (.L_HI(net1068));
 sg13g2_tiehi \ppu.sprite_buffer.top_prio[1]$_DFFE_PP__1069  (.L_HI(net1069));
 sg13g2_tiehi \ppu.sprite_buffer.top_prio[2]$_DFFE_PP__1070  (.L_HI(net1070));
 sg13g2_tiehi \ppu.sprite_buffer.top_prio[3]$_DFFE_PP__1071  (.L_HI(net1071));
 sg13g2_tiehi \ppu.sprite_buffer.top_prio[4]$_DFFE_PP__1072  (.L_HI(net1072));
 sg13g2_tiehi \ppu.sprite_buffer.top_prio[5]$_DFFE_PP__1073  (.L_HI(net1073));
 sg13g2_tiehi \ppu.sprite_buffer.top_prio[6]$_DFFE_PP__1074  (.L_HI(net1074));
 sg13g2_tiehi \ppu.sprite_buffer.valid_sprites[0]$_SDFFE_PP0P__1075  (.L_HI(net1075));
 sg13g2_tiehi \ppu.sprite_buffer.valid_sprites[1]$_SDFFE_PP0P__1076  (.L_HI(net1076));
 sg13g2_tiehi \ppu.sprite_buffer.valid_sprites[2]$_SDFFE_PP0P__1077  (.L_HI(net1077));
 sg13g2_tiehi \ppu.sprite_buffer.valid_sprites[3]$_SDFFE_PP0P__1078  (.L_HI(net1078));
 sg13g2_tiehi \ppu.sprite_buffer.y_matched0$_DFFE_PN__1079  (.L_HI(net1079));
 sg13g2_tiehi \ppu.sync_delay[0]$_SDFFE_PN1P__1080  (.L_HI(net1080));
 sg13g2_tiehi \ppu.sync_delay[1]$_SDFFE_PN1P__1081  (.L_HI(net1081));
 sg13g2_tiehi \ppu.sync_delay[2]$_SDFFE_PN1P__1082  (.L_HI(net1082));
 sg13g2_tiehi \ppu.tilemap.attr[0][0]$_DFFE_PP__1083  (.L_HI(net1083));
 sg13g2_tiehi \ppu.tilemap.attr[0][1]$_DFFE_PP__1084  (.L_HI(net1084));
 sg13g2_tiehi \ppu.tilemap.attr[0][2]$_DFFE_PP__1085  (.L_HI(net1085));
 sg13g2_tiehi \ppu.tilemap.attr[0][3]$_DFFE_PP__1086  (.L_HI(net1086));
 sg13g2_tiehi \ppu.tilemap.attr[0][4]$_DFFE_PP__1087  (.L_HI(net1087));
 sg13g2_tiehi \ppu.tilemap.attr[1][0]$_DFFE_PP__1088  (.L_HI(net1088));
 sg13g2_tiehi \ppu.tilemap.attr[1][1]$_DFFE_PP__1089  (.L_HI(net1089));
 sg13g2_tiehi \ppu.tilemap.attr[1][2]$_DFFE_PP__1090  (.L_HI(net1090));
 sg13g2_tiehi \ppu.tilemap.attr[1][3]$_DFFE_PP__1091  (.L_HI(net1091));
 sg13g2_tiehi \ppu.tilemap.attr[1][4]$_DFFE_PP__1092  (.L_HI(net1092));
 sg13g2_tiehi \ppu.tilemap.depth_out_reg[0]$_SDFFCE_PP0N__1093  (.L_HI(net1093));
 sg13g2_tiehi \ppu.tilemap.depth_out_reg[1]$_SDFFCE_PP0N__1094  (.L_HI(net1094));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][0]$_DFFE_PP__1095  (.L_HI(net1095));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][10]$_DFFE_PP__1096  (.L_HI(net1096));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][11]$_DFFE_PP__1097  (.L_HI(net1097));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][12]$_DFFE_PP__1098  (.L_HI(net1098));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][13]$_DFFE_PP__1099  (.L_HI(net1099));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][14]$_DFFE_PP__1100  (.L_HI(net1100));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][15]$_DFFE_PP__1101  (.L_HI(net1101));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][1]$_DFFE_PP__1102  (.L_HI(net1102));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][2]$_DFFE_PP__1103  (.L_HI(net1103));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][3]$_DFFE_PP__1104  (.L_HI(net1104));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][4]$_DFFE_PP__1105  (.L_HI(net1105));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][5]$_DFFE_PP__1106  (.L_HI(net1106));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][6]$_DFFE_PP__1107  (.L_HI(net1107));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][7]$_DFFE_PP__1108  (.L_HI(net1108));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][8]$_DFFE_PP__1109  (.L_HI(net1109));
 sg13g2_tiehi \ppu.tilemap.map_pixels[0][9]$_DFFE_PP__1110  (.L_HI(net1110));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][0]$_DFFE_PP__1111  (.L_HI(net1111));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][10]$_DFFE_PP__1112  (.L_HI(net1112));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][11]$_DFFE_PP__1113  (.L_HI(net1113));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][12]$_DFFE_PP__1114  (.L_HI(net1114));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][13]$_DFFE_PP__1115  (.L_HI(net1115));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][14]$_DFFE_PP__1116  (.L_HI(net1116));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][15]$_DFFE_PP__1117  (.L_HI(net1117));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][1]$_DFFE_PP__1118  (.L_HI(net1118));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][2]$_DFFE_PP__1119  (.L_HI(net1119));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][3]$_DFFE_PP__1120  (.L_HI(net1120));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][4]$_DFFE_PP__1121  (.L_HI(net1121));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][5]$_DFFE_PP__1122  (.L_HI(net1122));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][6]$_DFFE_PP__1123  (.L_HI(net1123));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][7]$_DFFE_PP__1124  (.L_HI(net1124));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][8]$_DFFE_PP__1125  (.L_HI(net1125));
 sg13g2_tiehi \ppu.tilemap.map_pixels[1][9]$_DFFE_PP__1126  (.L_HI(net1126));
 sg13g2_tiehi \ppu.tilemap.next_attr[0][0]$_DFFE_PP__1127  (.L_HI(net1127));
 sg13g2_tiehi \ppu.tilemap.next_attr[0][1]$_DFFE_PP__1128  (.L_HI(net1128));
 sg13g2_tiehi \ppu.tilemap.next_attr[0][2]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \ppu.tilemap.next_attr[0][3]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \ppu.tilemap.next_attr[0][4]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \ppu.tilemap.next_attr[1][0]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \ppu.tilemap.next_attr[1][1]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \ppu.tilemap.next_attr[1][2]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \ppu.tilemap.next_attr[1][3]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \ppu.tilemap.next_attr[1][4]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \ppu.tilemap.temp_out[0]$_DFFE_PN__1137  (.L_HI(net1137));
 sg13g2_tiehi \ppu.tilemap.temp_out[1]$_DFFE_PN__1138  (.L_HI(net1138));
 sg13g2_tiehi \ppu.tilemap.temp_out[2]$_DFFE_PN__1139  (.L_HI(net1139));
 sg13g2_tiehi \ppu.tilemap.temp_out[3]$_DFFE_PN__1140  (.L_HI(net1140));
 sg13g2_tiehi \reset$_DFF_P__1141  (.L_HI(net1141));
 sg13g2_tiehi \rx_in_reg[0]$_DFF_P__1142  (.L_HI(net1142));
 sg13g2_tiehi \rx_in_reg[1]$_DFF_P__1143  (.L_HI(net1143));
 sg13g2_tiehi \synth.controller.counter[0]$_SDFFE_PP1N__1144  (.L_HI(net1144));
 sg13g2_tiehi \synth.controller.counter[1]$_SDFFE_PP0N__1145  (.L_HI(net1145));
 sg13g2_tiehi \synth.controller.counter[2]$_SDFFE_PP1N__1146  (.L_HI(net1146));
 sg13g2_tiehi \synth.controller.counter[3]$_SDFFE_PP0N__1147  (.L_HI(net1147));
 sg13g2_tiehi \synth.controller.curr_voice[0]$_SDFFE_PP1N__1148  (.L_HI(net1148));
 sg13g2_tiehi \synth.controller.curr_voice[1]$_SDFFE_PP1N__1149  (.L_HI(net1149));
 sg13g2_tiehi \synth.controller.out_reg[0]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \synth.controller.out_reg[10]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \synth.controller.out_reg[11]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \synth.controller.out_reg[12]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \synth.controller.out_reg[13]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \synth.controller.out_reg[14]$_SDFFCE_PN0P__1155  (.L_HI(net1155));
 sg13g2_tiehi \synth.controller.out_reg[15]$_SDFFCE_PN0P__1156  (.L_HI(net1156));
 sg13g2_tiehi \synth.controller.out_reg[1]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \synth.controller.out_reg[2]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \synth.controller.out_reg[3]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \synth.controller.out_reg[4]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \synth.controller.out_reg[5]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \synth.controller.out_reg[6]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \synth.controller.out_reg[7]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \synth.controller.out_reg[8]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \synth.controller.out_reg[9]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \synth.controller.out_reg_valid$_SDFFE_PP0P__1166  (.L_HI(net1166));
 sg13g2_tiehi \synth.controller.ppu_ctrl_reg[0]$_SDFFE_PP1P__1167  (.L_HI(net1167));
 sg13g2_tiehi \synth.controller.ppu_ctrl_reg[2]$_SDFFE_PP0P__1168  (.L_HI(net1168));
 sg13g2_tiehi \synth.controller.ppu_ctrl_reg[3]$_SDFFE_PP1P__1169  (.L_HI(net1169));
 sg13g2_tiehi \synth.controller.ppu_ctrl_reg[4]$_SDFFE_PP0P__1170  (.L_HI(net1170));
 sg13g2_tiehi \synth.controller.read_index_reg[0]$_SDFFCE_PP0N__1171  (.L_HI(net1171));
 sg13g2_tiehi \synth.controller.read_index_reg[1]$_SDFFCE_PP0N__1172  (.L_HI(net1172));
 sg13g2_tiehi \synth.controller.read_index_reg[2]$_SDFFCE_PP0N__1173  (.L_HI(net1173));
 sg13g2_tiehi \synth.controller.read_index_reg[3]$_SDFFCE_PP0N__1174  (.L_HI(net1174));
 sg13g2_tiehi \synth.controller.rx_buffer[0]$_DFFE_PN__1175  (.L_HI(net1175));
 sg13g2_tiehi \synth.controller.rx_buffer[10]$_DFFE_PN__1176  (.L_HI(net1176));
 sg13g2_tiehi \synth.controller.rx_buffer[11]$_DFFE_PN__1177  (.L_HI(net1177));
 sg13g2_tiehi \synth.controller.rx_buffer[12]$_DFFE_PN__1178  (.L_HI(net1178));
 sg13g2_tiehi \synth.controller.rx_buffer[13]$_DFFE_PN__1179  (.L_HI(net1179));
 sg13g2_tiehi \synth.controller.rx_buffer[14]$_DFFE_PN__1180  (.L_HI(net1180));
 sg13g2_tiehi \synth.controller.rx_buffer[15]$_DFFE_PN__1181  (.L_HI(net1181));
 sg13g2_tiehi \synth.controller.rx_buffer[1]$_DFFE_PN__1182  (.L_HI(net1182));
 sg13g2_tiehi \synth.controller.rx_buffer[2]$_DFFE_PN__1183  (.L_HI(net1183));
 sg13g2_tiehi \synth.controller.rx_buffer[3]$_DFFE_PN__1184  (.L_HI(net1184));
 sg13g2_tiehi \synth.controller.rx_buffer[4]$_DFFE_PN__1185  (.L_HI(net1185));
 sg13g2_tiehi \synth.controller.rx_buffer[5]$_DFFE_PN__1186  (.L_HI(net1186));
 sg13g2_tiehi \synth.controller.rx_buffer[6]$_DFFE_PN__1187  (.L_HI(net1187));
 sg13g2_tiehi \synth.controller.rx_buffer[7]$_DFFE_PN__1188  (.L_HI(net1188));
 sg13g2_tiehi \synth.controller.rx_buffer[8]$_DFFE_PN__1189  (.L_HI(net1189));
 sg13g2_tiehi \synth.controller.rx_buffer[9]$_DFFE_PN__1190  (.L_HI(net1190));
 sg13g2_tiehi \synth.controller.rx_buffer_valid$_SDFF_PP0__1191  (.L_HI(net1191));
 sg13g2_tiehi \synth.controller.rx_sbs[0]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \synth.controller.rx_sbs[1]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \synth.controller.sample_counter[0]$_SDFFE_PP0N__1194  (.L_HI(net1194));
 sg13g2_tiehi \synth.controller.sample_counter[1]$_SDFFE_PP0N__1195  (.L_HI(net1195));
 sg13g2_tiehi \synth.controller.sample_credits[0]$_SDFF_PP1__1196  (.L_HI(net1196));
 sg13g2_tiehi \synth.controller.sample_credits[1]$_SDFF_PP0__1197  (.L_HI(net1197));
 sg13g2_tiehi \synth.controller.sbio_credits[0]$_SDFFE_PP1P__1198  (.L_HI(net1198));
 sg13g2_tiehi \synth.controller.sbio_credits[1]$_SDFFE_PP0P__1199  (.L_HI(net1199));
 sg13g2_tiehi \synth.controller.sbio_credits[2]$_SDFFE_PP0P__1200  (.L_HI(net1200));
 sg13g2_tiehi \synth.controller.sbio_rx.counter[0]$_SDFF_PP1__1201  (.L_HI(net1201));
 sg13g2_tiehi \synth.controller.sbio_rx.counter[1]$_SDFF_PP1__1202  (.L_HI(net1202));
 sg13g2_tiehi \synth.controller.sbio_rx.counter[2]$_SDFF_PP1__1203  (.L_HI(net1203));
 sg13g2_tiehi \synth.controller.sbio_rx.counter[3]$_SDFF_PP1__1204  (.L_HI(net1204));
 sg13g2_tiehi \synth.controller.sbio_tx.counter[0]$_SDFF_PP0__1205  (.L_HI(net1205));
 sg13g2_tiehi \synth.controller.sbio_tx.counter[1]$_SDFF_PP1__1206  (.L_HI(net1206));
 sg13g2_tiehi \synth.controller.sbio_tx.counter[2]$_SDFF_PP1__1207  (.L_HI(net1207));
 sg13g2_tiehi \synth.controller.sbio_tx.counter[3]$_SDFF_PP1__1208  (.L_HI(net1208));
 sg13g2_tiehi \synth.controller.scanning_out$_SDFFE_PP0P__1209  (.L_HI(net1209));
 sg13g2_tiehi \synth.controller.step_sample_reg$_SDFFE_PP1P__1210  (.L_HI(net1210));
 sg13g2_tiehi \synth.controller.sweep_addr_index[0]$_SDFF_PP1__1211  (.L_HI(net1211));
 sg13g2_tiehi \synth.controller.sweep_addr_index[1]$_SDFF_PP0__1212  (.L_HI(net1212));
 sg13g2_tiehi \synth.controller.sweep_addr_index[2]$_SDFF_PP1__1213  (.L_HI(net1213));
 sg13g2_tiehi \synth.controller.sweep_data_index[0]$_SDFF_PP1__1214  (.L_HI(net1214));
 sg13g2_tiehi \synth.controller.sweep_data_index[1]$_SDFF_PP0__1215  (.L_HI(net1215));
 sg13g2_tiehi \synth.controller.sweep_data_index[2]$_SDFF_PP1__1216  (.L_HI(net1216));
 sg13g2_tiehi \synth.controller.tx_outstanding[0]$_SDFF_PP0__1217  (.L_HI(net1217));
 sg13g2_tiehi \synth.controller.tx_outstanding[1]$_SDFF_PP0__1218  (.L_HI(net1218));
 sg13g2_tiehi \synth.controller.tx_outstanding[2]$_SDFF_PP0__1219  (.L_HI(net1219));
 sg13g2_tiehi \synth.controller.tx_source[0]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \synth.controller.tx_source[1]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \synth.controller.write_index_reg[0]$_SDFFCE_PP0N__1222  (.L_HI(net1222));
 sg13g2_tiehi \synth.controller.write_index_reg[1]$_SDFFCE_PP0N__1223  (.L_HI(net1223));
 sg13g2_tiehi \synth.controller.write_index_reg[2]$_SDFFCE_PP0N__1224  (.L_HI(net1224));
 sg13g2_tiehi \synth.controller.write_index_reg[3]$_SDFFCE_PP0N__1225  (.L_HI(net1225));
 sg13g2_tiehi \synth.voice.a_sel_reg[1]$_DFF_P__1226  (.L_HI(net1226));
 sg13g2_tiehi \synth.voice.a_sel_reg[2]$_DFF_P__1227  (.L_HI(net1227));
 sg13g2_tiehi \synth.voice.a_sel_reg[3]$_DFF_P__1228  (.L_HI(net1228));
 sg13g2_tiehi \synth.voice.accs[0][0]$_SDFFE_PP0P__1229  (.L_HI(net1229));
 sg13g2_tiehi \synth.voice.accs[0][10]$_SDFFE_PP0P__1230  (.L_HI(net1230));
 sg13g2_tiehi \synth.voice.accs[0][11]$_SDFFE_PP0P__1231  (.L_HI(net1231));
 sg13g2_tiehi \synth.voice.accs[0][12]$_SDFFE_PP0P__1232  (.L_HI(net1232));
 sg13g2_tiehi \synth.voice.accs[0][13]$_SDFFE_PP0P__1233  (.L_HI(net1233));
 sg13g2_tiehi \synth.voice.accs[0][14]$_SDFFE_PP0P__1234  (.L_HI(net1234));
 sg13g2_tiehi \synth.voice.accs[0][15]$_SDFFE_PP0P__1235  (.L_HI(net1235));
 sg13g2_tiehi \synth.voice.accs[0][16]$_SDFFE_PP0P__1236  (.L_HI(net1236));
 sg13g2_tiehi \synth.voice.accs[0][17]$_SDFFE_PP0P__1237  (.L_HI(net1237));
 sg13g2_tiehi \synth.voice.accs[0][18]$_SDFFE_PP0P__1238  (.L_HI(net1238));
 sg13g2_tiehi \synth.voice.accs[0][19]$_SDFFE_PP0P__1239  (.L_HI(net1239));
 sg13g2_tiehi \synth.voice.accs[0][1]$_SDFFE_PP0P__1240  (.L_HI(net1240));
 sg13g2_tiehi \synth.voice.accs[0][2]$_SDFFE_PP0P__1241  (.L_HI(net1241));
 sg13g2_tiehi \synth.voice.accs[0][3]$_SDFFE_PP0P__1242  (.L_HI(net1242));
 sg13g2_tiehi \synth.voice.accs[0][4]$_SDFFE_PP0P__1243  (.L_HI(net1243));
 sg13g2_tiehi \synth.voice.accs[0][5]$_SDFFE_PP0P__1244  (.L_HI(net1244));
 sg13g2_tiehi \synth.voice.accs[0][6]$_SDFFE_PP0P__1245  (.L_HI(net1245));
 sg13g2_tiehi \synth.voice.accs[0][7]$_SDFFE_PP0P__1246  (.L_HI(net1246));
 sg13g2_tiehi \synth.voice.accs[0][8]$_SDFFE_PP0P__1247  (.L_HI(net1247));
 sg13g2_tiehi \synth.voice.accs[0][9]$_SDFFE_PP0P__1248  (.L_HI(net1248));
 sg13g2_tiehi \synth.voice.accs[1][0]$_SDFFE_PP0P__1249  (.L_HI(net1249));
 sg13g2_tiehi \synth.voice.accs[1][10]$_SDFFE_PP0P__1250  (.L_HI(net1250));
 sg13g2_tiehi \synth.voice.accs[1][11]$_SDFFE_PP0P__1251  (.L_HI(net1251));
 sg13g2_tiehi \synth.voice.accs[1][12]$_SDFFE_PP0P__1252  (.L_HI(net1252));
 sg13g2_tiehi \synth.voice.accs[1][13]$_SDFFE_PP0P__1253  (.L_HI(net1253));
 sg13g2_tiehi \synth.voice.accs[1][14]$_SDFFE_PP0P__1254  (.L_HI(net1254));
 sg13g2_tiehi \synth.voice.accs[1][15]$_SDFFE_PP0P__1255  (.L_HI(net1255));
 sg13g2_tiehi \synth.voice.accs[1][16]$_SDFFE_PP0P__1256  (.L_HI(net1256));
 sg13g2_tiehi \synth.voice.accs[1][17]$_SDFFE_PP0P__1257  (.L_HI(net1257));
 sg13g2_tiehi \synth.voice.accs[1][18]$_SDFFE_PP0P__1258  (.L_HI(net1258));
 sg13g2_tiehi \synth.voice.accs[1][19]$_SDFFE_PP0P__1259  (.L_HI(net1259));
 sg13g2_tiehi \synth.voice.accs[1][1]$_SDFFE_PP0P__1260  (.L_HI(net1260));
 sg13g2_tiehi \synth.voice.accs[1][2]$_SDFFE_PP0P__1261  (.L_HI(net1261));
 sg13g2_tiehi \synth.voice.accs[1][3]$_SDFFE_PP0P__1262  (.L_HI(net1262));
 sg13g2_tiehi \synth.voice.accs[1][4]$_SDFFE_PP0P__1263  (.L_HI(net1263));
 sg13g2_tiehi \synth.voice.accs[1][5]$_SDFFE_PP0P__1264  (.L_HI(net1264));
 sg13g2_tiehi \synth.voice.accs[1][6]$_SDFFE_PP0P__1265  (.L_HI(net1265));
 sg13g2_tiehi \synth.voice.accs[1][7]$_SDFFE_PP0P__1266  (.L_HI(net1266));
 sg13g2_tiehi \synth.voice.accs[1][8]$_SDFFE_PP0P__1267  (.L_HI(net1267));
 sg13g2_tiehi \synth.voice.accs[1][9]$_SDFFE_PP0P__1268  (.L_HI(net1268));
 sg13g2_tiehi \synth.voice.accs[2][0]$_SDFFE_PP0P__1269  (.L_HI(net1269));
 sg13g2_tiehi \synth.voice.accs[2][10]$_SDFFE_PP0P__1270  (.L_HI(net1270));
 sg13g2_tiehi \synth.voice.accs[2][11]$_SDFFE_PP0P__1271  (.L_HI(net1271));
 sg13g2_tiehi \synth.voice.accs[2][12]$_SDFFE_PP0P__1272  (.L_HI(net1272));
 sg13g2_tiehi \synth.voice.accs[2][13]$_SDFFE_PP0P__1273  (.L_HI(net1273));
 sg13g2_tiehi \synth.voice.accs[2][14]$_SDFFE_PP0P__1274  (.L_HI(net1274));
 sg13g2_tiehi \synth.voice.accs[2][15]$_SDFFE_PP0P__1275  (.L_HI(net1275));
 sg13g2_tiehi \synth.voice.accs[2][16]$_SDFFE_PP0P__1276  (.L_HI(net1276));
 sg13g2_tiehi \synth.voice.accs[2][17]$_SDFFE_PP0P__1277  (.L_HI(net1277));
 sg13g2_tiehi \synth.voice.accs[2][18]$_SDFFE_PP0P__1278  (.L_HI(net1278));
 sg13g2_tiehi \synth.voice.accs[2][19]$_SDFFE_PP0P__1279  (.L_HI(net1279));
 sg13g2_tiehi \synth.voice.accs[2][1]$_SDFFE_PP0P__1280  (.L_HI(net1280));
 sg13g2_tiehi \synth.voice.accs[2][2]$_SDFFE_PP0P__1281  (.L_HI(net1281));
 sg13g2_tiehi \synth.voice.accs[2][3]$_SDFFE_PP0P__1282  (.L_HI(net1282));
 sg13g2_tiehi \synth.voice.accs[2][4]$_SDFFE_PP0P__1283  (.L_HI(net1283));
 sg13g2_tiehi \synth.voice.accs[2][5]$_SDFFE_PP0P__1284  (.L_HI(net1284));
 sg13g2_tiehi \synth.voice.accs[2][6]$_SDFFE_PP0P__1285  (.L_HI(net1285));
 sg13g2_tiehi \synth.voice.accs[2][7]$_SDFFE_PP0P__1286  (.L_HI(net1286));
 sg13g2_tiehi \synth.voice.accs[2][8]$_SDFFE_PP0P__1287  (.L_HI(net1287));
 sg13g2_tiehi \synth.voice.accs[2][9]$_SDFFE_PP0P__1288  (.L_HI(net1288));
 sg13g2_tiehi \synth.voice.accs[3][0]$_SDFFE_PP0P__1289  (.L_HI(net1289));
 sg13g2_tiehi \synth.voice.accs[3][10]$_SDFFE_PP0P__1290  (.L_HI(net1290));
 sg13g2_tiehi \synth.voice.accs[3][11]$_SDFFE_PP0P__1291  (.L_HI(net1291));
 sg13g2_tiehi \synth.voice.accs[3][12]$_SDFFE_PP0P__1292  (.L_HI(net1292));
 sg13g2_tiehi \synth.voice.accs[3][13]$_SDFFE_PP0P__1293  (.L_HI(net1293));
 sg13g2_tiehi \synth.voice.accs[3][14]$_SDFFE_PP0P__1294  (.L_HI(net1294));
 sg13g2_tiehi \synth.voice.accs[3][15]$_SDFFE_PP0P__1295  (.L_HI(net1295));
 sg13g2_tiehi \synth.voice.accs[3][16]$_SDFFE_PP0P__1296  (.L_HI(net1296));
 sg13g2_tiehi \synth.voice.accs[3][17]$_SDFFE_PP0P__1297  (.L_HI(net1297));
 sg13g2_tiehi \synth.voice.accs[3][18]$_SDFFE_PP0P__1298  (.L_HI(net1298));
 sg13g2_tiehi \synth.voice.accs[3][19]$_SDFFE_PP0P__1299  (.L_HI(net1299));
 sg13g2_tiehi \synth.voice.accs[3][1]$_SDFFE_PP0P__1300  (.L_HI(net1300));
 sg13g2_tiehi \synth.voice.accs[3][2]$_SDFFE_PP0P__1301  (.L_HI(net1301));
 sg13g2_tiehi \synth.voice.accs[3][3]$_SDFFE_PP0P__1302  (.L_HI(net1302));
 sg13g2_tiehi \synth.voice.accs[3][4]$_SDFFE_PP0P__1303  (.L_HI(net1303));
 sg13g2_tiehi \synth.voice.accs[3][5]$_SDFFE_PP0P__1304  (.L_HI(net1304));
 sg13g2_tiehi \synth.voice.accs[3][6]$_SDFFE_PP0P__1305  (.L_HI(net1305));
 sg13g2_tiehi \synth.voice.accs[3][7]$_SDFFE_PP0P__1306  (.L_HI(net1306));
 sg13g2_tiehi \synth.voice.accs[3][8]$_SDFFE_PP0P__1307  (.L_HI(net1307));
 sg13g2_tiehi \synth.voice.accs[3][9]$_SDFFE_PP0P__1308  (.L_HI(net1308));
 sg13g2_tiehi \synth.voice.accs[4][0]$_SDFFE_PP0P__1309  (.L_HI(net1309));
 sg13g2_tiehi \synth.voice.accs[4][10]$_SDFFE_PP0P__1310  (.L_HI(net1310));
 sg13g2_tiehi \synth.voice.accs[4][11]$_SDFFE_PP0P__1311  (.L_HI(net1311));
 sg13g2_tiehi \synth.voice.accs[4][12]$_SDFFE_PP0P__1312  (.L_HI(net1312));
 sg13g2_tiehi \synth.voice.accs[4][13]$_SDFFE_PP0P__1313  (.L_HI(net1313));
 sg13g2_tiehi \synth.voice.accs[4][14]$_SDFFE_PP0P__1314  (.L_HI(net1314));
 sg13g2_tiehi \synth.voice.accs[4][15]$_SDFFE_PP0P__1315  (.L_HI(net1315));
 sg13g2_tiehi \synth.voice.accs[4][16]$_SDFFE_PP0P__1316  (.L_HI(net1316));
 sg13g2_tiehi \synth.voice.accs[4][17]$_SDFFE_PP0P__1317  (.L_HI(net1317));
 sg13g2_tiehi \synth.voice.accs[4][18]$_SDFFE_PP0P__1318  (.L_HI(net1318));
 sg13g2_tiehi \synth.voice.accs[4][19]$_SDFFE_PP0P__1319  (.L_HI(net1319));
 sg13g2_tiehi \synth.voice.accs[4][1]$_SDFFE_PP0P__1320  (.L_HI(net1320));
 sg13g2_tiehi \synth.voice.accs[4][2]$_SDFFE_PP0P__1321  (.L_HI(net1321));
 sg13g2_tiehi \synth.voice.accs[4][3]$_SDFFE_PP0P__1322  (.L_HI(net1322));
 sg13g2_tiehi \synth.voice.accs[4][4]$_SDFFE_PP0P__1323  (.L_HI(net1323));
 sg13g2_tiehi \synth.voice.accs[4][5]$_SDFFE_PP0P__1324  (.L_HI(net1324));
 sg13g2_tiehi \synth.voice.accs[4][6]$_SDFFE_PP0P__1325  (.L_HI(net1325));
 sg13g2_tiehi \synth.voice.accs[4][7]$_SDFFE_PP0P__1326  (.L_HI(net1326));
 sg13g2_tiehi \synth.voice.accs[4][8]$_SDFFE_PP0P__1327  (.L_HI(net1327));
 sg13g2_tiehi \synth.voice.accs[4][9]$_SDFFE_PP0P__1328  (.L_HI(net1328));
 sg13g2_tiehi \synth.voice.accs[5][0]$_SDFFE_PP0P__1329  (.L_HI(net1329));
 sg13g2_tiehi \synth.voice.accs[5][10]$_SDFFE_PP0P__1330  (.L_HI(net1330));
 sg13g2_tiehi \synth.voice.accs[5][11]$_SDFFE_PP0P__1331  (.L_HI(net1331));
 sg13g2_tiehi \synth.voice.accs[5][12]$_SDFFE_PP0P__1332  (.L_HI(net1332));
 sg13g2_tiehi \synth.voice.accs[5][13]$_SDFFE_PP0P__1333  (.L_HI(net1333));
 sg13g2_tiehi \synth.voice.accs[5][14]$_SDFFE_PP0P__1334  (.L_HI(net1334));
 sg13g2_tiehi \synth.voice.accs[5][15]$_SDFFE_PP0P__1335  (.L_HI(net1335));
 sg13g2_tiehi \synth.voice.accs[5][16]$_SDFFE_PP0P__1336  (.L_HI(net1336));
 sg13g2_tiehi \synth.voice.accs[5][17]$_SDFFE_PP0P__1337  (.L_HI(net1337));
 sg13g2_tiehi \synth.voice.accs[5][18]$_SDFFE_PP0P__1338  (.L_HI(net1338));
 sg13g2_tiehi \synth.voice.accs[5][19]$_SDFFE_PP0P__1339  (.L_HI(net1339));
 sg13g2_tiehi \synth.voice.accs[5][1]$_SDFFE_PP0P__1340  (.L_HI(net1340));
 sg13g2_tiehi \synth.voice.accs[5][2]$_SDFFE_PP0P__1341  (.L_HI(net1341));
 sg13g2_tiehi \synth.voice.accs[5][3]$_SDFFE_PP0P__1342  (.L_HI(net1342));
 sg13g2_tiehi \synth.voice.accs[5][4]$_SDFFE_PP0P__1343  (.L_HI(net1343));
 sg13g2_tiehi \synth.voice.accs[5][5]$_SDFFE_PP0P__1344  (.L_HI(net1344));
 sg13g2_tiehi \synth.voice.accs[5][6]$_SDFFE_PP0P__1345  (.L_HI(net1345));
 sg13g2_tiehi \synth.voice.accs[5][7]$_SDFFE_PP0P__1346  (.L_HI(net1346));
 sg13g2_tiehi \synth.voice.accs[5][8]$_SDFFE_PP0P__1347  (.L_HI(net1347));
 sg13g2_tiehi \synth.voice.accs[5][9]$_SDFFE_PP0P__1348  (.L_HI(net1348));
 sg13g2_tiehi \synth.voice.b_sel_reg[0]$_DFF_P__1349  (.L_HI(net1349));
 sg13g2_tiehi \synth.voice.b_sel_reg[2]$_DFF_P__1350  (.L_HI(net1350));
 sg13g2_tiehi \synth.voice.fir_offset_msbs[0]$_SDFF_PN0__1351  (.L_HI(net1351));
 sg13g2_tiehi \synth.voice.fir_offset_msbs[1]$_SDFF_PN0__1352  (.L_HI(net1352));
 sg13g2_tiehi \synth.voice.flip_sign_fir$_DFF_P__1353  (.L_HI(net1353));
 sg13g2_tiehi \synth.voice.flip_sign_reg$_DFF_P__1354  (.L_HI(net1354));
 sg13g2_tiehi \synth.voice.oct_counter[0]$_SDFFE_PP0P__1355  (.L_HI(net1355));
 sg13g2_tiehi \synth.voice.oct_counter[10]$_SDFFE_PP0P__1356  (.L_HI(net1356));
 sg13g2_tiehi \synth.voice.oct_counter[1]$_SDFFE_PP0P__1357  (.L_HI(net1357));
 sg13g2_tiehi \synth.voice.oct_counter[2]$_SDFFE_PP0P__1358  (.L_HI(net1358));
 sg13g2_tiehi \synth.voice.oct_counter[3]$_SDFFE_PP0P__1359  (.L_HI(net1359));
 sg13g2_tiehi \synth.voice.oct_counter[4]$_SDFFE_PP0P__1360  (.L_HI(net1360));
 sg13g2_tiehi \synth.voice.oct_counter[5]$_SDFFE_PP0P__1361  (.L_HI(net1361));
 sg13g2_tiehi \synth.voice.oct_counter[6]$_SDFFE_PP0P__1362  (.L_HI(net1362));
 sg13g2_tiehi \synth.voice.oct_counter[7]$_SDFFE_PP0P__1363  (.L_HI(net1363));
 sg13g2_tiehi \synth.voice.oct_counter[8]$_SDFFE_PP0P__1364  (.L_HI(net1364));
 sg13g2_tiehi \synth.voice.oct_counter[9]$_SDFFE_PP0P__1365  (.L_HI(net1365));
 sg13g2_tiehi \synth.voice.restart_acc_reg$_DFF_P__1366  (.L_HI(net1366));
 sg13g2_tiehi \synth.voice.rshift_reg0[0]$_DFF_P__1367  (.L_HI(net1367));
 sg13g2_tiehi \synth.voice.rshift_reg0[1]$_DFF_P__1368  (.L_HI(net1368));
 sg13g2_tiehi \synth.voice.rshift_reg0[2]$_DFF_P__1369  (.L_HI(net1369));
 sg13g2_tiehi \synth.voice.rshift_reg0[3]$_DFF_P__1370  (.L_HI(net1370));
 sg13g2_tiehi \synth.voice.rshift_reg[0]$_DFF_P__1371  (.L_HI(net1371));
 sg13g2_tiehi \synth.voice.rshift_reg[1]$_DFF_P__1372  (.L_HI(net1372));
 sg13g2_tiehi \synth.voice.rshift_reg[2]$_DFF_P__1373  (.L_HI(net1373));
 sg13g2_tiehi \synth.voice.rshift_reg[3]$_DFF_P__1374  (.L_HI(net1374));
 sg13g2_tiehi \synth.voice.scan_accs_reg$_DFF_P__1375  (.L_HI(net1375));
 sg13g2_tiehi \synth.voice.state[0]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \synth.voice.state[100]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \synth.voice.state[101]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \synth.voice.state[102]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \synth.voice.state[103]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \synth.voice.state[104]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \synth.voice.state[105]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \synth.voice.state[106]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \synth.voice.state[107]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \synth.voice.state[108]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \synth.voice.state[109]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \synth.voice.state[10]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \synth.voice.state[110]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \synth.voice.state[111]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \synth.voice.state[112]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \synth.voice.state[113]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \synth.voice.state[114]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \synth.voice.state[115]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \synth.voice.state[116]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \synth.voice.state[117]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \synth.voice.state[118]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \synth.voice.state[119]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \synth.voice.state[11]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \synth.voice.state[120]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \synth.voice.state[121]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \synth.voice.state[122]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \synth.voice.state[123]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \synth.voice.state[124]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \synth.voice.state[125]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \synth.voice.state[126]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \synth.voice.state[127]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \synth.voice.state[128]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \synth.voice.state[129]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \synth.voice.state[12]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \synth.voice.state[130]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \synth.voice.state[131]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \synth.voice.state[132]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \synth.voice.state[133]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \synth.voice.state[134]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \synth.voice.state[135]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \synth.voice.state[136]$_DFFE_PN__1416  (.L_HI(net1416));
 sg13g2_tiehi \synth.voice.state[137]$_DFFE_PN__1417  (.L_HI(net1417));
 sg13g2_tiehi \synth.voice.state[138]$_DFFE_PN__1418  (.L_HI(net1418));
 sg13g2_tiehi \synth.voice.state[139]$_DFFE_PN__1419  (.L_HI(net1419));
 sg13g2_tiehi \synth.voice.state[13]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \synth.voice.state[140]$_DFFE_PN__1421  (.L_HI(net1421));
 sg13g2_tiehi \synth.voice.state[141]$_DFFE_PN__1422  (.L_HI(net1422));
 sg13g2_tiehi \synth.voice.state[142]$_DFFE_PN__1423  (.L_HI(net1423));
 sg13g2_tiehi \synth.voice.state[143]$_DFFE_PN__1424  (.L_HI(net1424));
 sg13g2_tiehi \synth.voice.state[144]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \synth.voice.state[145]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \synth.voice.state[146]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \synth.voice.state[147]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \synth.voice.state[148]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \synth.voice.state[149]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \synth.voice.state[14]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \synth.voice.state[150]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \synth.voice.state[151]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \synth.voice.state[152]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \synth.voice.state[153]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \synth.voice.state[154]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \synth.voice.state[155]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \synth.voice.state[156]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \synth.voice.state[157]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \synth.voice.state[158]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \synth.voice.state[159]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \synth.voice.state[15]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \synth.voice.state[160]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \synth.voice.state[161]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \synth.voice.state[162]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \synth.voice.state[163]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \synth.voice.state[164]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \synth.voice.state[165]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \synth.voice.state[166]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \synth.voice.state[167]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \synth.voice.state[168]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \synth.voice.state[169]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \synth.voice.state[16]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \synth.voice.state[170]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \synth.voice.state[171]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \synth.voice.state[172]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \synth.voice.state[173]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \synth.voice.state[174]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \synth.voice.state[175]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \synth.voice.state[176]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \synth.voice.state[177]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \synth.voice.state[178]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \synth.voice.state[179]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \synth.voice.state[17]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \synth.voice.state[180]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \synth.voice.state[181]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \synth.voice.state[182]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \synth.voice.state[183]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \synth.voice.state[184]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \synth.voice.state[185]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \synth.voice.state[186]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \synth.voice.state[187]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \synth.voice.state[188]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \synth.voice.state[189]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \synth.voice.state[18]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \synth.voice.state[190]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \synth.voice.state[191]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \synth.voice.state[19]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \synth.voice.state[1]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \synth.voice.state[20]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \synth.voice.state[21]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \synth.voice.state[22]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \synth.voice.state[23]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \synth.voice.state[24]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \synth.voice.state[25]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \synth.voice.state[26]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \synth.voice.state[27]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \synth.voice.state[28]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \synth.voice.state[29]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \synth.voice.state[2]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \synth.voice.state[30]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \synth.voice.state[31]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \synth.voice.state[32]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \synth.voice.state[33]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \synth.voice.state[34]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \synth.voice.state[35]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \synth.voice.state[36]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \synth.voice.state[37]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \synth.voice.state[38]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \synth.voice.state[39]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \synth.voice.state[3]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \synth.voice.state[40]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \synth.voice.state[41]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \synth.voice.state[42]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \synth.voice.state[43]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \synth.voice.state[44]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \synth.voice.state[45]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \synth.voice.state[46]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \synth.voice.state[47]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \synth.voice.state[48]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \synth.voice.state[49]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \synth.voice.state[4]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \synth.voice.state[50]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \synth.voice.state[51]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \synth.voice.state[52]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \synth.voice.state[53]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \synth.voice.state[54]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \synth.voice.state[55]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \synth.voice.state[56]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \synth.voice.state[57]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \synth.voice.state[58]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \synth.voice.state[59]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \synth.voice.state[5]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \synth.voice.state[60]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \synth.voice.state[61]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \synth.voice.state[62]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \synth.voice.state[63]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \synth.voice.state[64]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \synth.voice.state[65]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \synth.voice.state[66]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \synth.voice.state[67]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \synth.voice.state[68]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \synth.voice.state[69]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \synth.voice.state[6]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \synth.voice.state[70]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \synth.voice.state[71]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \synth.voice.state[72]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \synth.voice.state[73]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \synth.voice.state[74]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \synth.voice.state[75]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \synth.voice.state[76]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \synth.voice.state[77]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \synth.voice.state[78]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \synth.voice.state[79]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \synth.voice.state[7]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \synth.voice.state[80]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \synth.voice.state[81]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \synth.voice.state[82]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \synth.voice.state[83]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \synth.voice.state[84]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \synth.voice.state[85]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \synth.voice.state[86]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \synth.voice.state[87]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \synth.voice.state[88]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \synth.voice.state[89]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \synth.voice.state[8]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \synth.voice.state[90]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \synth.voice.state[91]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \synth.voice.state[92]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \synth.voice.state[93]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \synth.voice.state[94]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \synth.voice.state[95]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \synth.voice.state[96]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \synth.voice.state[97]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \synth.voice.state[98]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \synth.voice.state[99]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \synth.voice.state[9]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[0]$_SDFFE_PP0P__1568  (.L_HI(net1568));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[10]$_SDFFE_PP0P__1569  (.L_HI(net1569));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[11]$_SDFFE_PP0P__1570  (.L_HI(net1570));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[12]$_SDFFE_PP0P__1571  (.L_HI(net1571));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[13]$_SDFFE_PP0P__1572  (.L_HI(net1572));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[1]$_SDFFE_PP0P__1573  (.L_HI(net1573));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[2]$_SDFFE_PP0P__1574  (.L_HI(net1574));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[3]$_SDFFE_PP0P__1575  (.L_HI(net1575));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[4]$_SDFFE_PP0P__1576  (.L_HI(net1576));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[5]$_SDFFE_PP0P__1577  (.L_HI(net1577));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[6]$_SDFFE_PP0P__1578  (.L_HI(net1578));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[7]$_SDFFE_PP0P__1579  (.L_HI(net1579));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[8]$_SDFFE_PP0P__1580  (.L_HI(net1580));
 sg13g2_tiehi \synth.voice.sweep_oct_counter[9]$_SDFFE_PP0P__1581  (.L_HI(net1581));
 sg13g2_tiehi \synth.voice.tap[0]$_SDFF_PP0__1582  (.L_HI(net1582));
 sg13g2_tiehi \synth.voice.tap[1]$_SDFF_PP0__1583  (.L_HI(net1583));
 sg13g2_tiehi \synth.voice.target_reg[1]$_DFF_P__1584  (.L_HI(net1584));
 sg13g2_tiehi \synth.voice.target_reg[2]$_DFF_P__1585  (.L_HI(net1585));
 sg13g2_tiehi \synth.voice.target_reg[3]$_DFF_P__1586  (.L_HI(net1586));
 sg13g2_tiehi \synth.voice.term_index[0]$_SDFF_PP0__1587  (.L_HI(net1587));
 sg13g2_tiehi \synth.voice.term_index[1]$_SDFF_PP0__1588  (.L_HI(net1588));
 sg13g2_tiehi \synth.voice.term_index[2]$_SDFF_PP0__1589  (.L_HI(net1589));
 sg13g2_tiehi \synth.voice.wave_reg[0]$_SDFFCE_PP0P__1590  (.L_HI(net1590));
 sg13g2_tiehi \synth.voice.wave_reg[1]$_SDFFCE_PP0P__1591  (.L_HI(net1591));
 sg13g2_tiehi \synth.voice.wave_reg[2]$_SDFFCE_PP0P__1592  (.L_HI(net1592));
 sg13g2_tiehi \synth.voice.wave_reg[3]$_SDFFCE_PP0P__1593  (.L_HI(net1593));
 sg13g2_tiehi \synth.voice.wave_reg[4]$_SDFFCE_PP0P__1594  (.L_HI(net1594));
 sg13g2_tiehi \synth.voice.wave_reg[5]$_SDFFCE_PP0P__1595  (.L_HI(net1595));
 sg13g2_tiehi \synth.voice.wave_reg[6]$_SDFFCE_PP0P__1596  (.L_HI(net1596));
 sg13g2_tiehi \synth.voice.wave_reg[7]$_SDFFCE_PP1P__1597  (.L_HI(net1597));
 sg13g2_tiehi \synth.voice.wave_reg[8]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \synth.voice.wave_reg[9]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \synth.voice.zero_shifter_out_reg$_DFF_P__1600  (.L_HI(net1600));
 sg13g2_tiehi \ui_in_reg[0]$_DFF_P__1601  (.L_HI(net1601));
 sg13g2_tiehi \ui_in_reg[1]$_DFF_P__1602  (.L_HI(net1602));
 sg13g2_tiehi \ui_in_reg[2]$_DFF_P__1603  (.L_HI(net1603));
 sg13g2_tiehi \ui_in_reg[3]$_DFF_P__1604  (.L_HI(net1604));
 sg13g2_tiehi \uio_out_reg[0]$_DFF_P__1605  (.L_HI(net1605));
 sg13g2_tiehi \uio_out_reg[1]$_DFF_P__1606  (.L_HI(net1606));
 sg13g2_tiehi \uio_out_reg[2]$_DFF_P__1607  (.L_HI(net1607));
 sg13g2_tiehi \uio_out_reg[3]$_DFF_P__1608  (.L_HI(net1608));
 sg13g2_tiehi \uio_out_reg[4]$_DFF_P__1609  (.L_HI(net1609));
 sg13g2_tiehi \uio_out_reg[5]$_SDFF_PP0__1610  (.L_HI(net1610));
 sg13g2_tiehi \uio_out_reg[6]$_DFF_P__1611  (.L_HI(net1611));
 sg13g2_tiehi \uio_out_reg[7]$_DFF_P__1612  (.L_HI(net1612));
 sg13g2_tiehi \uo_out_reg[0]$_DFF_P__1613  (.L_HI(net1613));
 sg13g2_tiehi \uo_out_reg[1]$_DFF_P__1614  (.L_HI(net1614));
 sg13g2_tiehi \uo_out_reg[2]$_DFF_P__1615  (.L_HI(net1615));
 sg13g2_tiehi \uo_out_reg[3]$_DFF_P__1616  (.L_HI(net1616));
 sg13g2_tiehi \uo_out_reg[4]$_DFF_P__1617  (.L_HI(net1617));
 sg13g2_tiehi \uo_out_reg[5]$_DFF_P__1618  (.L_HI(net1618));
 sg13g2_tiehi \uo_out_reg[6]$_DFF_P__1619  (.L_HI(net1619));
 sg13g2_tiehi \uo_out_reg[7]$_DFF_P__1620  (.L_HI(net1620));
 sg13g2_tiehi \vblank_pending$_SDFF_PP0__1621  (.L_HI(net1621));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_62_clk (.X(clknet_leaf_62_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_63_clk (.X(clknet_leaf_63_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_64_clk (.X(clknet_leaf_64_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_65_clk (.X(clknet_leaf_65_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_66_clk (.X(clknet_leaf_66_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_67_clk (.X(clknet_leaf_67_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_68_clk (.X(clknet_leaf_68_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_69_clk (.X(clknet_leaf_69_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_70_clk (.X(clknet_leaf_70_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_71_clk (.X(clknet_leaf_71_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_72_clk (.X(clknet_leaf_72_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_73_clk (.X(clknet_leaf_73_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_74_clk (.X(clknet_leaf_74_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_75_clk (.X(clknet_leaf_75_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_76_clk (.X(clknet_leaf_76_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_77_clk (.X(clknet_leaf_77_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_78_clk (.X(clknet_leaf_78_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_79_clk (.X(clknet_leaf_79_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_80_clk (.X(clknet_leaf_80_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_81_clk (.X(clknet_leaf_81_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_82_clk (.X(clknet_leaf_82_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_83_clk (.X(clknet_leaf_83_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_84_clk (.X(clknet_leaf_84_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_85_clk (.X(clknet_leaf_85_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_86_clk (.X(clknet_leaf_86_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_87_clk (.X(clknet_leaf_87_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_88_clk (.X(clknet_leaf_88_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_89_clk (.X(clknet_leaf_89_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_90_clk (.X(clknet_leaf_90_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_91_clk (.X(clknet_leaf_91_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_92_clk (.X(clknet_leaf_92_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_93_clk (.X(clknet_leaf_93_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_94_clk (.X(clknet_leaf_94_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_95_clk (.X(clknet_leaf_95_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_96_clk (.X(clknet_leaf_96_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_97_clk (.X(clknet_leaf_97_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_98_clk (.X(clknet_leaf_98_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_99_clk (.X(clknet_leaf_99_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_100_clk (.X(clknet_leaf_100_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_101_clk (.X(clknet_leaf_101_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_102_clk (.X(clknet_leaf_102_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_103_clk (.X(clknet_leaf_103_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_104_clk (.X(clknet_leaf_104_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_105_clk (.X(clknet_leaf_105_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_106_clk (.X(clknet_leaf_106_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_107_clk (.X(clknet_leaf_107_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_108_clk (.X(clknet_leaf_108_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_109_clk (.X(clknet_leaf_109_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_110_clk (.X(clknet_leaf_110_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_111_clk (.X(clknet_leaf_111_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_112_clk (.X(clknet_leaf_112_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_113_clk (.X(clknet_leaf_113_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_114_clk (.X(clknet_leaf_114_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_115_clk (.X(clknet_leaf_115_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_116_clk (.X(clknet_leaf_116_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_117_clk (.X(clknet_leaf_117_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_118_clk (.X(clknet_leaf_118_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_119_clk (.X(clknet_leaf_119_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_120_clk (.X(clknet_leaf_120_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_121_clk (.X(clknet_leaf_121_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_122_clk (.X(clknet_leaf_122_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_123_clk (.X(clknet_leaf_123_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_124_clk (.X(clknet_leaf_124_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_125_clk (.X(clknet_leaf_125_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_126_clk (.X(clknet_leaf_126_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_127_clk (.X(clknet_leaf_127_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_128_clk (.X(clknet_leaf_128_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_129_clk (.X(clknet_leaf_129_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_130_clk (.X(clknet_leaf_130_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_131_clk (.X(clknet_leaf_131_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_132_clk (.X(clknet_leaf_132_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_133_clk (.X(clknet_leaf_133_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_134_clk (.X(clknet_leaf_134_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_135_clk (.X(clknet_leaf_135_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_136_clk (.X(clknet_leaf_136_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_137_clk (.X(clknet_leaf_137_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_138_clk (.X(clknet_leaf_138_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_139_clk (.X(clknet_leaf_139_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_140_clk (.X(clknet_leaf_140_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_141_clk (.X(clknet_leaf_141_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_142_clk (.X(clknet_leaf_142_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_143_clk (.X(clknet_leaf_143_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_144_clk (.X(clknet_leaf_144_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_145_clk (.X(clknet_leaf_145_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_146_clk (.X(clknet_leaf_146_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_147_clk (.X(clknet_leaf_147_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_148_clk (.X(clknet_leaf_148_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_149_clk (.X(clknet_leaf_149_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_150_clk (.X(clknet_leaf_150_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkload3 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkload4 (.A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkload5 (.A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkload6 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkload7 (.A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkload8 (.A(clknet_5_31__leaf_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_150_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_02686_));
 sg13g2_antennanp ANTENNA_2 (.A(_02686_));
 sg13g2_antennanp ANTENNA_3 (.A(_02686_));
 sg13g2_antennanp ANTENNA_4 (.A(_07677_));
 sg13g2_antennanp ANTENNA_5 (.A(_07677_));
 sg13g2_antennanp ANTENNA_6 (.A(\addr_pins_out[1] ));
 sg13g2_antennanp ANTENNA_7 (.A(\addr_pins_out[2] ));
 sg13g2_antennanp ANTENNA_8 (.A(clk));
 sg13g2_antennanp ANTENNA_9 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_10 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_11 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_12 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_13 (.A(hsync));
 sg13g2_antennanp ANTENNA_14 (.A(hsync));
 sg13g2_antennanp ANTENNA_15 (.A(hsync));
 sg13g2_antennanp ANTENNA_16 (.A(hsync));
 sg13g2_antennanp ANTENNA_17 (.A(hsync));
 sg13g2_antennanp ANTENNA_18 (.A(\ppu.pal_data_out[2] ));
 sg13g2_antennanp ANTENNA_19 (.A(\ppu.pal_data_out[2] ));
 sg13g2_antennanp ANTENNA_20 (.A(_02686_));
 sg13g2_antennanp ANTENNA_21 (.A(_02686_));
 sg13g2_antennanp ANTENNA_22 (.A(_02686_));
 sg13g2_antennanp ANTENNA_23 (.A(_07677_));
 sg13g2_antennanp ANTENNA_24 (.A(_07677_));
 sg13g2_antennanp ANTENNA_25 (.A(\addr_pins_out[0] ));
 sg13g2_antennanp ANTENNA_26 (.A(\addr_pins_out[2] ));
 sg13g2_antennanp ANTENNA_27 (.A(clk));
 sg13g2_antennanp ANTENNA_28 (.A(clk));
 sg13g2_antennanp ANTENNA_29 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_30 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_31 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_32 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_33 (.A(hsync));
 sg13g2_antennanp ANTENNA_34 (.A(hsync));
 sg13g2_antennanp ANTENNA_35 (.A(hsync));
 sg13g2_antennanp ANTENNA_36 (.A(hsync));
 sg13g2_antennanp ANTENNA_37 (.A(hsync));
 sg13g2_antennanp ANTENNA_38 (.A(\ppu.pal_data_out[2] ));
 sg13g2_antennanp ANTENNA_39 (.A(\ppu.pal_data_out[2] ));
 sg13g2_antennanp ANTENNA_40 (.A(_02686_));
 sg13g2_antennanp ANTENNA_41 (.A(_02686_));
 sg13g2_antennanp ANTENNA_42 (.A(_02686_));
 sg13g2_antennanp ANTENNA_43 (.A(_07677_));
 sg13g2_antennanp ANTENNA_44 (.A(_07677_));
 sg13g2_antennanp ANTENNA_45 (.A(\addr_pins_out[0] ));
 sg13g2_antennanp ANTENNA_46 (.A(clk));
 sg13g2_antennanp ANTENNA_47 (.A(clk));
 sg13g2_antennanp ANTENNA_48 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_49 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_50 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_51 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_52 (.A(\ppu.pal_data_out[2] ));
 sg13g2_antennanp ANTENNA_53 (.A(\ppu.pal_data_out[2] ));
 sg13g2_antennanp ANTENNA_54 (.A(_02686_));
 sg13g2_antennanp ANTENNA_55 (.A(_02686_));
 sg13g2_antennanp ANTENNA_56 (.A(_02686_));
 sg13g2_antennanp ANTENNA_57 (.A(_07677_));
 sg13g2_antennanp ANTENNA_58 (.A(_07677_));
 sg13g2_antennanp ANTENNA_59 (.A(\addr_pins_out[0] ));
 sg13g2_antennanp ANTENNA_60 (.A(\addr_pins_out[0] ));
 sg13g2_antennanp ANTENNA_61 (.A(clk));
 sg13g2_antennanp ANTENNA_62 (.A(clk));
 sg13g2_antennanp ANTENNA_63 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_64 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_65 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_66 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_67 (.A(_02686_));
 sg13g2_antennanp ANTENNA_68 (.A(_02686_));
 sg13g2_antennanp ANTENNA_69 (.A(_02686_));
 sg13g2_antennanp ANTENNA_70 (.A(_07677_));
 sg13g2_antennanp ANTENNA_71 (.A(_07677_));
 sg13g2_antennanp ANTENNA_72 (.A(\addr_pins_out[0] ));
 sg13g2_antennanp ANTENNA_73 (.A(\addr_pins_out[0] ));
 sg13g2_antennanp ANTENNA_74 (.A(clk));
 sg13g2_antennanp ANTENNA_75 (.A(clk));
 sg13g2_antennanp ANTENNA_76 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_77 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_78 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_79 (.A(\data_pins[2] ));
 sg13g2_antennanp ANTENNA_80 (.A(hsync));
 sg13g2_antennanp ANTENNA_81 (.A(hsync));
 sg13g2_antennanp ANTENNA_82 (.A(hsync));
 sg13g2_antennanp ANTENNA_83 (.A(hsync));
 sg13g2_antennanp ANTENNA_84 (.A(hsync));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_4 FILLER_0_42 ();
 sg13g2_fill_2 FILLER_0_46 ();
 sg13g2_decap_8 FILLER_0_52 ();
 sg13g2_fill_2 FILLER_0_59 ();
 sg13g2_fill_1 FILLER_0_61 ();
 sg13g2_decap_8 FILLER_0_65 ();
 sg13g2_decap_8 FILLER_0_72 ();
 sg13g2_decap_4 FILLER_0_79 ();
 sg13g2_fill_2 FILLER_0_87 ();
 sg13g2_decap_8 FILLER_0_101 ();
 sg13g2_fill_2 FILLER_0_112 ();
 sg13g2_fill_1 FILLER_0_114 ();
 sg13g2_decap_8 FILLER_0_120 ();
 sg13g2_decap_4 FILLER_0_127 ();
 sg13g2_fill_2 FILLER_0_138 ();
 sg13g2_fill_2 FILLER_0_145 ();
 sg13g2_fill_1 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_178 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_fill_2 FILLER_0_213 ();
 sg13g2_fill_1 FILLER_0_215 ();
 sg13g2_decap_4 FILLER_0_246 ();
 sg13g2_fill_1 FILLER_0_250 ();
 sg13g2_decap_4 FILLER_0_277 ();
 sg13g2_fill_1 FILLER_0_281 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_decap_4 FILLER_0_333 ();
 sg13g2_fill_2 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_fill_2 FILLER_0_376 ();
 sg13g2_fill_2 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_436 ();
 sg13g2_fill_1 FILLER_0_440 ();
 sg13g2_decap_8 FILLER_0_467 ();
 sg13g2_decap_8 FILLER_0_474 ();
 sg13g2_fill_1 FILLER_0_481 ();
 sg13g2_fill_1 FILLER_0_512 ();
 sg13g2_decap_8 FILLER_0_517 ();
 sg13g2_decap_8 FILLER_0_524 ();
 sg13g2_fill_1 FILLER_0_531 ();
 sg13g2_decap_8 FILLER_0_544 ();
 sg13g2_decap_4 FILLER_0_551 ();
 sg13g2_decap_8 FILLER_0_565 ();
 sg13g2_decap_8 FILLER_0_572 ();
 sg13g2_fill_2 FILLER_0_579 ();
 sg13g2_fill_1 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_608 ();
 sg13g2_fill_1 FILLER_0_615 ();
 sg13g2_decap_8 FILLER_0_646 ();
 sg13g2_fill_2 FILLER_0_653 ();
 sg13g2_decap_8 FILLER_0_659 ();
 sg13g2_decap_8 FILLER_0_666 ();
 sg13g2_decap_8 FILLER_0_673 ();
 sg13g2_decap_8 FILLER_0_680 ();
 sg13g2_decap_8 FILLER_0_687 ();
 sg13g2_decap_4 FILLER_0_694 ();
 sg13g2_fill_2 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_726 ();
 sg13g2_fill_1 FILLER_0_763 ();
 sg13g2_fill_2 FILLER_0_808 ();
 sg13g2_fill_1 FILLER_0_810 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_fill_1 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_827 ();
 sg13g2_decap_8 FILLER_0_860 ();
 sg13g2_fill_1 FILLER_0_867 ();
 sg13g2_decap_8 FILLER_0_894 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_4 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_1020 ();
 sg13g2_decap_8 FILLER_0_1027 ();
 sg13g2_fill_1 FILLER_0_1034 ();
 sg13g2_decap_8 FILLER_0_1039 ();
 sg13g2_decap_8 FILLER_0_1046 ();
 sg13g2_decap_8 FILLER_0_1053 ();
 sg13g2_decap_8 FILLER_0_1060 ();
 sg13g2_decap_8 FILLER_0_1067 ();
 sg13g2_decap_4 FILLER_0_1074 ();
 sg13g2_fill_2 FILLER_0_1078 ();
 sg13g2_decap_8 FILLER_0_1084 ();
 sg13g2_fill_2 FILLER_0_1091 ();
 sg13g2_fill_1 FILLER_0_1093 ();
 sg13g2_decap_8 FILLER_0_1114 ();
 sg13g2_decap_8 FILLER_0_1121 ();
 sg13g2_fill_1 FILLER_0_1128 ();
 sg13g2_fill_2 FILLER_0_1139 ();
 sg13g2_fill_1 FILLER_0_1141 ();
 sg13g2_fill_1 FILLER_0_1146 ();
 sg13g2_decap_8 FILLER_0_1157 ();
 sg13g2_decap_8 FILLER_0_1168 ();
 sg13g2_decap_8 FILLER_0_1175 ();
 sg13g2_decap_8 FILLER_0_1182 ();
 sg13g2_decap_8 FILLER_0_1189 ();
 sg13g2_decap_8 FILLER_0_1196 ();
 sg13g2_decap_8 FILLER_0_1203 ();
 sg13g2_decap_8 FILLER_0_1210 ();
 sg13g2_decap_8 FILLER_0_1217 ();
 sg13g2_decap_8 FILLER_0_1224 ();
 sg13g2_decap_8 FILLER_0_1231 ();
 sg13g2_decap_8 FILLER_0_1238 ();
 sg13g2_decap_8 FILLER_0_1245 ();
 sg13g2_decap_8 FILLER_0_1252 ();
 sg13g2_decap_8 FILLER_0_1259 ();
 sg13g2_decap_8 FILLER_0_1266 ();
 sg13g2_decap_8 FILLER_0_1273 ();
 sg13g2_decap_8 FILLER_0_1280 ();
 sg13g2_decap_8 FILLER_0_1287 ();
 sg13g2_decap_8 FILLER_0_1294 ();
 sg13g2_decap_8 FILLER_0_1301 ();
 sg13g2_decap_8 FILLER_0_1308 ();
 sg13g2_decap_8 FILLER_0_1315 ();
 sg13g2_decap_4 FILLER_0_1322 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_4 FILLER_1_28 ();
 sg13g2_decap_4 FILLER_1_35 ();
 sg13g2_fill_2 FILLER_1_39 ();
 sg13g2_fill_2 FILLER_1_49 ();
 sg13g2_fill_1 FILLER_1_51 ();
 sg13g2_fill_2 FILLER_1_60 ();
 sg13g2_fill_1 FILLER_1_94 ();
 sg13g2_decap_4 FILLER_1_101 ();
 sg13g2_fill_1 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_117 ();
 sg13g2_fill_2 FILLER_1_124 ();
 sg13g2_fill_1 FILLER_1_129 ();
 sg13g2_fill_2 FILLER_1_142 ();
 sg13g2_fill_2 FILLER_1_149 ();
 sg13g2_decap_8 FILLER_1_155 ();
 sg13g2_decap_8 FILLER_1_162 ();
 sg13g2_fill_2 FILLER_1_169 ();
 sg13g2_fill_1 FILLER_1_171 ();
 sg13g2_decap_8 FILLER_1_177 ();
 sg13g2_decap_4 FILLER_1_184 ();
 sg13g2_fill_2 FILLER_1_188 ();
 sg13g2_decap_8 FILLER_1_194 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_decap_8 FILLER_1_212 ();
 sg13g2_decap_4 FILLER_1_219 ();
 sg13g2_fill_2 FILLER_1_223 ();
 sg13g2_fill_1 FILLER_1_230 ();
 sg13g2_decap_4 FILLER_1_236 ();
 sg13g2_fill_2 FILLER_1_240 ();
 sg13g2_fill_1 FILLER_1_247 ();
 sg13g2_decap_8 FILLER_1_253 ();
 sg13g2_fill_1 FILLER_1_260 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_fill_2 FILLER_1_277 ();
 sg13g2_fill_1 FILLER_1_279 ();
 sg13g2_fill_2 FILLER_1_283 ();
 sg13g2_fill_2 FILLER_1_295 ();
 sg13g2_fill_1 FILLER_1_297 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_decap_8 FILLER_1_327 ();
 sg13g2_decap_8 FILLER_1_334 ();
 sg13g2_decap_4 FILLER_1_341 ();
 sg13g2_decap_4 FILLER_1_350 ();
 sg13g2_decap_4 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_fill_1 FILLER_1_381 ();
 sg13g2_fill_2 FILLER_1_391 ();
 sg13g2_fill_1 FILLER_1_393 ();
 sg13g2_fill_1 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_424 ();
 sg13g2_fill_1 FILLER_1_431 ();
 sg13g2_fill_1 FILLER_1_472 ();
 sg13g2_fill_2 FILLER_1_478 ();
 sg13g2_decap_4 FILLER_1_501 ();
 sg13g2_fill_1 FILLER_1_505 ();
 sg13g2_fill_1 FILLER_1_593 ();
 sg13g2_fill_2 FILLER_1_599 ();
 sg13g2_fill_1 FILLER_1_601 ();
 sg13g2_fill_2 FILLER_1_633 ();
 sg13g2_decap_8 FILLER_1_674 ();
 sg13g2_decap_8 FILLER_1_681 ();
 sg13g2_decap_8 FILLER_1_688 ();
 sg13g2_fill_2 FILLER_1_695 ();
 sg13g2_fill_1 FILLER_1_697 ();
 sg13g2_fill_2 FILLER_1_719 ();
 sg13g2_fill_2 FILLER_1_725 ();
 sg13g2_decap_4 FILLER_1_731 ();
 sg13g2_fill_2 FILLER_1_735 ();
 sg13g2_fill_2 FILLER_1_741 ();
 sg13g2_fill_1 FILLER_1_743 ();
 sg13g2_fill_1 FILLER_1_748 ();
 sg13g2_decap_8 FILLER_1_775 ();
 sg13g2_decap_4 FILLER_1_782 ();
 sg13g2_fill_2 FILLER_1_786 ();
 sg13g2_decap_8 FILLER_1_792 ();
 sg13g2_fill_2 FILLER_1_840 ();
 sg13g2_fill_1 FILLER_1_842 ();
 sg13g2_decap_4 FILLER_1_855 ();
 sg13g2_fill_1 FILLER_1_864 ();
 sg13g2_fill_1 FILLER_1_869 ();
 sg13g2_fill_1 FILLER_1_874 ();
 sg13g2_decap_4 FILLER_1_879 ();
 sg13g2_fill_2 FILLER_1_883 ();
 sg13g2_decap_4 FILLER_1_902 ();
 sg13g2_fill_2 FILLER_1_906 ();
 sg13g2_decap_8 FILLER_1_912 ();
 sg13g2_decap_8 FILLER_1_919 ();
 sg13g2_decap_8 FILLER_1_926 ();
 sg13g2_decap_8 FILLER_1_933 ();
 sg13g2_decap_8 FILLER_1_940 ();
 sg13g2_decap_8 FILLER_1_947 ();
 sg13g2_decap_8 FILLER_1_954 ();
 sg13g2_decap_8 FILLER_1_961 ();
 sg13g2_decap_8 FILLER_1_968 ();
 sg13g2_decap_8 FILLER_1_975 ();
 sg13g2_decap_8 FILLER_1_982 ();
 sg13g2_decap_8 FILLER_1_989 ();
 sg13g2_decap_4 FILLER_1_996 ();
 sg13g2_fill_1 FILLER_1_1000 ();
 sg13g2_fill_1 FILLER_1_1005 ();
 sg13g2_fill_1 FILLER_1_1026 ();
 sg13g2_decap_8 FILLER_1_1053 ();
 sg13g2_decap_8 FILLER_1_1060 ();
 sg13g2_decap_4 FILLER_1_1067 ();
 sg13g2_fill_2 FILLER_1_1071 ();
 sg13g2_fill_2 FILLER_1_1099 ();
 sg13g2_fill_1 FILLER_1_1101 ();
 sg13g2_fill_2 FILLER_1_1128 ();
 sg13g2_fill_1 FILLER_1_1130 ();
 sg13g2_decap_8 FILLER_1_1183 ();
 sg13g2_decap_8 FILLER_1_1190 ();
 sg13g2_decap_8 FILLER_1_1197 ();
 sg13g2_decap_8 FILLER_1_1204 ();
 sg13g2_decap_8 FILLER_1_1211 ();
 sg13g2_decap_8 FILLER_1_1218 ();
 sg13g2_decap_8 FILLER_1_1225 ();
 sg13g2_decap_8 FILLER_1_1232 ();
 sg13g2_decap_8 FILLER_1_1239 ();
 sg13g2_decap_8 FILLER_1_1246 ();
 sg13g2_decap_8 FILLER_1_1253 ();
 sg13g2_decap_8 FILLER_1_1260 ();
 sg13g2_decap_8 FILLER_1_1267 ();
 sg13g2_decap_8 FILLER_1_1274 ();
 sg13g2_decap_8 FILLER_1_1281 ();
 sg13g2_decap_8 FILLER_1_1288 ();
 sg13g2_decap_8 FILLER_1_1295 ();
 sg13g2_decap_8 FILLER_1_1302 ();
 sg13g2_decap_8 FILLER_1_1309 ();
 sg13g2_decap_8 FILLER_1_1316 ();
 sg13g2_fill_2 FILLER_1_1323 ();
 sg13g2_fill_1 FILLER_1_1325 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_4 FILLER_2_28 ();
 sg13g2_fill_2 FILLER_2_32 ();
 sg13g2_decap_4 FILLER_2_42 ();
 sg13g2_fill_2 FILLER_2_46 ();
 sg13g2_fill_2 FILLER_2_56 ();
 sg13g2_fill_1 FILLER_2_62 ();
 sg13g2_fill_1 FILLER_2_69 ();
 sg13g2_fill_1 FILLER_2_75 ();
 sg13g2_decap_4 FILLER_2_100 ();
 sg13g2_fill_2 FILLER_2_104 ();
 sg13g2_fill_2 FILLER_2_114 ();
 sg13g2_decap_4 FILLER_2_120 ();
 sg13g2_fill_1 FILLER_2_128 ();
 sg13g2_decap_8 FILLER_2_135 ();
 sg13g2_fill_1 FILLER_2_142 ();
 sg13g2_fill_2 FILLER_2_151 ();
 sg13g2_decap_4 FILLER_2_164 ();
 sg13g2_fill_1 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_174 ();
 sg13g2_fill_2 FILLER_2_181 ();
 sg13g2_fill_1 FILLER_2_183 ();
 sg13g2_fill_1 FILLER_2_210 ();
 sg13g2_fill_1 FILLER_2_241 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_fill_2 FILLER_2_265 ();
 sg13g2_fill_1 FILLER_2_285 ();
 sg13g2_decap_4 FILLER_2_294 ();
 sg13g2_decap_4 FILLER_2_311 ();
 sg13g2_fill_1 FILLER_2_315 ();
 sg13g2_fill_2 FILLER_2_342 ();
 sg13g2_fill_1 FILLER_2_373 ();
 sg13g2_decap_4 FILLER_2_383 ();
 sg13g2_fill_1 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_fill_2 FILLER_2_398 ();
 sg13g2_fill_1 FILLER_2_400 ();
 sg13g2_fill_1 FILLER_2_405 ();
 sg13g2_fill_1 FILLER_2_458 ();
 sg13g2_fill_1 FILLER_2_490 ();
 sg13g2_decap_4 FILLER_2_517 ();
 sg13g2_fill_2 FILLER_2_521 ();
 sg13g2_decap_4 FILLER_2_541 ();
 sg13g2_fill_1 FILLER_2_545 ();
 sg13g2_fill_2 FILLER_2_551 ();
 sg13g2_fill_2 FILLER_2_561 ();
 sg13g2_fill_1 FILLER_2_567 ();
 sg13g2_fill_2 FILLER_2_573 ();
 sg13g2_fill_2 FILLER_2_583 ();
 sg13g2_fill_1 FILLER_2_585 ();
 sg13g2_fill_2 FILLER_2_589 ();
 sg13g2_fill_1 FILLER_2_591 ();
 sg13g2_fill_2 FILLER_2_597 ();
 sg13g2_fill_1 FILLER_2_599 ();
 sg13g2_decap_4 FILLER_2_603 ();
 sg13g2_fill_1 FILLER_2_607 ();
 sg13g2_decap_4 FILLER_2_612 ();
 sg13g2_fill_1 FILLER_2_616 ();
 sg13g2_fill_1 FILLER_2_620 ();
 sg13g2_fill_2 FILLER_2_626 ();
 sg13g2_decap_4 FILLER_2_633 ();
 sg13g2_fill_2 FILLER_2_637 ();
 sg13g2_fill_2 FILLER_2_642 ();
 sg13g2_fill_2 FILLER_2_703 ();
 sg13g2_fill_2 FILLER_2_751 ();
 sg13g2_fill_2 FILLER_2_766 ();
 sg13g2_decap_8 FILLER_2_804 ();
 sg13g2_fill_2 FILLER_2_811 ();
 sg13g2_fill_1 FILLER_2_813 ();
 sg13g2_fill_1 FILLER_2_818 ();
 sg13g2_decap_8 FILLER_2_822 ();
 sg13g2_fill_1 FILLER_2_829 ();
 sg13g2_decap_4 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_848 ();
 sg13g2_decap_8 FILLER_2_855 ();
 sg13g2_fill_2 FILLER_2_896 ();
 sg13g2_fill_1 FILLER_2_898 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_fill_2 FILLER_2_970 ();
 sg13g2_fill_1 FILLER_2_972 ();
 sg13g2_decap_8 FILLER_2_983 ();
 sg13g2_decap_8 FILLER_2_990 ();
 sg13g2_fill_2 FILLER_2_997 ();
 sg13g2_fill_1 FILLER_2_999 ();
 sg13g2_decap_8 FILLER_2_1010 ();
 sg13g2_decap_8 FILLER_2_1017 ();
 sg13g2_decap_8 FILLER_2_1024 ();
 sg13g2_decap_4 FILLER_2_1031 ();
 sg13g2_fill_1 FILLER_2_1035 ();
 sg13g2_decap_4 FILLER_2_1072 ();
 sg13g2_fill_2 FILLER_2_1076 ();
 sg13g2_decap_4 FILLER_2_1104 ();
 sg13g2_fill_2 FILLER_2_1108 ();
 sg13g2_decap_8 FILLER_2_1114 ();
 sg13g2_decap_8 FILLER_2_1121 ();
 sg13g2_decap_4 FILLER_2_1128 ();
 sg13g2_fill_2 FILLER_2_1132 ();
 sg13g2_fill_1 FILLER_2_1144 ();
 sg13g2_decap_8 FILLER_2_1155 ();
 sg13g2_decap_8 FILLER_2_1162 ();
 sg13g2_decap_4 FILLER_2_1169 ();
 sg13g2_fill_2 FILLER_2_1173 ();
 sg13g2_decap_8 FILLER_2_1185 ();
 sg13g2_decap_8 FILLER_2_1192 ();
 sg13g2_decap_8 FILLER_2_1199 ();
 sg13g2_decap_8 FILLER_2_1206 ();
 sg13g2_decap_8 FILLER_2_1213 ();
 sg13g2_decap_8 FILLER_2_1220 ();
 sg13g2_decap_8 FILLER_2_1227 ();
 sg13g2_decap_8 FILLER_2_1234 ();
 sg13g2_decap_8 FILLER_2_1241 ();
 sg13g2_decap_8 FILLER_2_1248 ();
 sg13g2_decap_8 FILLER_2_1255 ();
 sg13g2_decap_8 FILLER_2_1262 ();
 sg13g2_decap_8 FILLER_2_1269 ();
 sg13g2_decap_8 FILLER_2_1276 ();
 sg13g2_decap_8 FILLER_2_1283 ();
 sg13g2_decap_8 FILLER_2_1290 ();
 sg13g2_decap_8 FILLER_2_1297 ();
 sg13g2_decap_8 FILLER_2_1304 ();
 sg13g2_decap_8 FILLER_2_1311 ();
 sg13g2_decap_8 FILLER_2_1318 ();
 sg13g2_fill_1 FILLER_2_1325 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_1 FILLER_3_28 ();
 sg13g2_decap_4 FILLER_3_36 ();
 sg13g2_fill_2 FILLER_3_40 ();
 sg13g2_fill_1 FILLER_3_46 ();
 sg13g2_decap_4 FILLER_3_50 ();
 sg13g2_fill_2 FILLER_3_78 ();
 sg13g2_fill_2 FILLER_3_91 ();
 sg13g2_fill_2 FILLER_3_97 ();
 sg13g2_fill_1 FILLER_3_99 ();
 sg13g2_fill_2 FILLER_3_113 ();
 sg13g2_decap_4 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_136 ();
 sg13g2_fill_1 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_158 ();
 sg13g2_fill_1 FILLER_3_160 ();
 sg13g2_fill_2 FILLER_3_169 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_decap_8 FILLER_3_198 ();
 sg13g2_decap_8 FILLER_3_205 ();
 sg13g2_fill_2 FILLER_3_212 ();
 sg13g2_fill_1 FILLER_3_214 ();
 sg13g2_fill_2 FILLER_3_223 ();
 sg13g2_decap_4 FILLER_3_234 ();
 sg13g2_fill_2 FILLER_3_290 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_fill_2 FILLER_3_315 ();
 sg13g2_fill_1 FILLER_3_317 ();
 sg13g2_decap_8 FILLER_3_352 ();
 sg13g2_decap_4 FILLER_3_359 ();
 sg13g2_fill_1 FILLER_3_363 ();
 sg13g2_fill_1 FILLER_3_372 ();
 sg13g2_fill_1 FILLER_3_404 ();
 sg13g2_decap_8 FILLER_3_425 ();
 sg13g2_decap_8 FILLER_3_432 ();
 sg13g2_fill_2 FILLER_3_439 ();
 sg13g2_decap_4 FILLER_3_445 ();
 sg13g2_fill_1 FILLER_3_449 ();
 sg13g2_decap_4 FILLER_3_456 ();
 sg13g2_fill_1 FILLER_3_460 ();
 sg13g2_fill_1 FILLER_3_469 ();
 sg13g2_decap_4 FILLER_3_474 ();
 sg13g2_fill_1 FILLER_3_481 ();
 sg13g2_fill_2 FILLER_3_509 ();
 sg13g2_fill_1 FILLER_3_511 ();
 sg13g2_fill_2 FILLER_3_516 ();
 sg13g2_fill_2 FILLER_3_544 ();
 sg13g2_fill_2 FILLER_3_572 ();
 sg13g2_fill_2 FILLER_3_613 ();
 sg13g2_fill_1 FILLER_3_615 ();
 sg13g2_decap_8 FILLER_3_668 ();
 sg13g2_decap_8 FILLER_3_675 ();
 sg13g2_fill_2 FILLER_3_682 ();
 sg13g2_decap_8 FILLER_3_688 ();
 sg13g2_fill_2 FILLER_3_708 ();
 sg13g2_fill_1 FILLER_3_710 ();
 sg13g2_fill_2 FILLER_3_716 ();
 sg13g2_fill_1 FILLER_3_718 ();
 sg13g2_fill_2 FILLER_3_723 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_4 FILLER_3_742 ();
 sg13g2_fill_2 FILLER_3_746 ();
 sg13g2_fill_1 FILLER_3_755 ();
 sg13g2_fill_1 FILLER_3_765 ();
 sg13g2_fill_1 FILLER_3_774 ();
 sg13g2_fill_2 FILLER_3_785 ();
 sg13g2_fill_1 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_792 ();
 sg13g2_decap_4 FILLER_3_799 ();
 sg13g2_decap_8 FILLER_3_863 ();
 sg13g2_fill_1 FILLER_3_870 ();
 sg13g2_decap_4 FILLER_3_883 ();
 sg13g2_fill_1 FILLER_3_887 ();
 sg13g2_fill_2 FILLER_3_892 ();
 sg13g2_decap_8 FILLER_3_898 ();
 sg13g2_fill_2 FILLER_3_905 ();
 sg13g2_fill_2 FILLER_3_917 ();
 sg13g2_fill_1 FILLER_3_919 ();
 sg13g2_fill_2 FILLER_3_924 ();
 sg13g2_fill_1 FILLER_3_926 ();
 sg13g2_decap_8 FILLER_3_931 ();
 sg13g2_decap_8 FILLER_3_938 ();
 sg13g2_decap_8 FILLER_3_945 ();
 sg13g2_decap_8 FILLER_3_952 ();
 sg13g2_fill_2 FILLER_3_1037 ();
 sg13g2_decap_8 FILLER_3_1069 ();
 sg13g2_decap_8 FILLER_3_1076 ();
 sg13g2_fill_1 FILLER_3_1083 ();
 sg13g2_decap_8 FILLER_3_1088 ();
 sg13g2_fill_1 FILLER_3_1095 ();
 sg13g2_decap_8 FILLER_3_1106 ();
 sg13g2_fill_2 FILLER_3_1149 ();
 sg13g2_fill_1 FILLER_3_1151 ();
 sg13g2_fill_2 FILLER_3_1178 ();
 sg13g2_fill_1 FILLER_3_1180 ();
 sg13g2_decap_8 FILLER_3_1207 ();
 sg13g2_decap_8 FILLER_3_1214 ();
 sg13g2_decap_8 FILLER_3_1221 ();
 sg13g2_decap_8 FILLER_3_1228 ();
 sg13g2_decap_8 FILLER_3_1235 ();
 sg13g2_decap_8 FILLER_3_1242 ();
 sg13g2_decap_8 FILLER_3_1249 ();
 sg13g2_decap_8 FILLER_3_1256 ();
 sg13g2_decap_8 FILLER_3_1263 ();
 sg13g2_decap_8 FILLER_3_1270 ();
 sg13g2_decap_8 FILLER_3_1277 ();
 sg13g2_decap_8 FILLER_3_1284 ();
 sg13g2_decap_8 FILLER_3_1291 ();
 sg13g2_decap_8 FILLER_3_1298 ();
 sg13g2_decap_8 FILLER_3_1305 ();
 sg13g2_decap_8 FILLER_3_1312 ();
 sg13g2_decap_8 FILLER_3_1319 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_21 ();
 sg13g2_fill_2 FILLER_4_31 ();
 sg13g2_fill_1 FILLER_4_44 ();
 sg13g2_fill_2 FILLER_4_49 ();
 sg13g2_fill_1 FILLER_4_51 ();
 sg13g2_fill_2 FILLER_4_58 ();
 sg13g2_fill_1 FILLER_4_65 ();
 sg13g2_fill_2 FILLER_4_81 ();
 sg13g2_fill_1 FILLER_4_92 ();
 sg13g2_decap_4 FILLER_4_97 ();
 sg13g2_fill_1 FILLER_4_101 ();
 sg13g2_fill_1 FILLER_4_105 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_fill_1 FILLER_4_128 ();
 sg13g2_decap_4 FILLER_4_133 ();
 sg13g2_fill_2 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_fill_1 FILLER_4_158 ();
 sg13g2_fill_2 FILLER_4_164 ();
 sg13g2_fill_1 FILLER_4_170 ();
 sg13g2_fill_1 FILLER_4_176 ();
 sg13g2_fill_1 FILLER_4_181 ();
 sg13g2_fill_2 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_4 FILLER_4_200 ();
 sg13g2_fill_1 FILLER_4_204 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_fill_2 FILLER_4_217 ();
 sg13g2_fill_2 FILLER_4_227 ();
 sg13g2_fill_1 FILLER_4_246 ();
 sg13g2_fill_2 FILLER_4_252 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_258 ();
 sg13g2_decap_4 FILLER_4_301 ();
 sg13g2_fill_2 FILLER_4_310 ();
 sg13g2_fill_2 FILLER_4_316 ();
 sg13g2_fill_1 FILLER_4_318 ();
 sg13g2_fill_2 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_325 ();
 sg13g2_decap_4 FILLER_4_330 ();
 sg13g2_fill_2 FILLER_4_334 ();
 sg13g2_fill_1 FILLER_4_341 ();
 sg13g2_fill_1 FILLER_4_347 ();
 sg13g2_fill_1 FILLER_4_374 ();
 sg13g2_fill_2 FILLER_4_380 ();
 sg13g2_fill_1 FILLER_4_411 ();
 sg13g2_fill_1 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_517 ();
 sg13g2_fill_2 FILLER_4_524 ();
 sg13g2_fill_1 FILLER_4_526 ();
 sg13g2_fill_2 FILLER_4_532 ();
 sg13g2_fill_1 FILLER_4_534 ();
 sg13g2_decap_8 FILLER_4_538 ();
 sg13g2_fill_2 FILLER_4_545 ();
 sg13g2_decap_4 FILLER_4_550 ();
 sg13g2_fill_1 FILLER_4_554 ();
 sg13g2_fill_1 FILLER_4_559 ();
 sg13g2_fill_2 FILLER_4_563 ();
 sg13g2_fill_1 FILLER_4_565 ();
 sg13g2_fill_2 FILLER_4_571 ();
 sg13g2_decap_4 FILLER_4_576 ();
 sg13g2_fill_2 FILLER_4_585 ();
 sg13g2_decap_8 FILLER_4_591 ();
 sg13g2_decap_4 FILLER_4_598 ();
 sg13g2_fill_2 FILLER_4_602 ();
 sg13g2_fill_2 FILLER_4_608 ();
 sg13g2_fill_1 FILLER_4_615 ();
 sg13g2_decap_8 FILLER_4_621 ();
 sg13g2_fill_2 FILLER_4_628 ();
 sg13g2_fill_2 FILLER_4_642 ();
 sg13g2_fill_1 FILLER_4_678 ();
 sg13g2_fill_1 FILLER_4_705 ();
 sg13g2_fill_1 FILLER_4_810 ();
 sg13g2_fill_2 FILLER_4_816 ();
 sg13g2_fill_2 FILLER_4_831 ();
 sg13g2_fill_1 FILLER_4_842 ();
 sg13g2_decap_8 FILLER_4_848 ();
 sg13g2_decap_8 FILLER_4_869 ();
 sg13g2_decap_8 FILLER_4_876 ();
 sg13g2_fill_2 FILLER_4_913 ();
 sg13g2_fill_1 FILLER_4_915 ();
 sg13g2_decap_8 FILLER_4_942 ();
 sg13g2_decap_4 FILLER_4_949 ();
 sg13g2_fill_2 FILLER_4_953 ();
 sg13g2_decap_8 FILLER_4_971 ();
 sg13g2_fill_2 FILLER_4_978 ();
 sg13g2_fill_1 FILLER_4_980 ();
 sg13g2_decap_8 FILLER_4_995 ();
 sg13g2_decap_8 FILLER_4_1002 ();
 sg13g2_decap_4 FILLER_4_1009 ();
 sg13g2_fill_1 FILLER_4_1053 ();
 sg13g2_decap_8 FILLER_4_1080 ();
 sg13g2_decap_8 FILLER_4_1087 ();
 sg13g2_fill_2 FILLER_4_1094 ();
 sg13g2_fill_1 FILLER_4_1096 ();
 sg13g2_fill_2 FILLER_4_1127 ();
 sg13g2_fill_1 FILLER_4_1129 ();
 sg13g2_decap_8 FILLER_4_1134 ();
 sg13g2_decap_8 FILLER_4_1141 ();
 sg13g2_decap_4 FILLER_4_1148 ();
 sg13g2_fill_2 FILLER_4_1162 ();
 sg13g2_decap_4 FILLER_4_1168 ();
 sg13g2_fill_2 FILLER_4_1176 ();
 sg13g2_decap_8 FILLER_4_1192 ();
 sg13g2_decap_8 FILLER_4_1199 ();
 sg13g2_decap_8 FILLER_4_1206 ();
 sg13g2_decap_8 FILLER_4_1213 ();
 sg13g2_decap_8 FILLER_4_1220 ();
 sg13g2_decap_8 FILLER_4_1227 ();
 sg13g2_decap_8 FILLER_4_1234 ();
 sg13g2_decap_8 FILLER_4_1241 ();
 sg13g2_decap_8 FILLER_4_1248 ();
 sg13g2_decap_8 FILLER_4_1255 ();
 sg13g2_decap_8 FILLER_4_1262 ();
 sg13g2_decap_8 FILLER_4_1269 ();
 sg13g2_decap_8 FILLER_4_1276 ();
 sg13g2_decap_8 FILLER_4_1283 ();
 sg13g2_decap_8 FILLER_4_1290 ();
 sg13g2_decap_8 FILLER_4_1297 ();
 sg13g2_decap_8 FILLER_4_1304 ();
 sg13g2_decap_8 FILLER_4_1311 ();
 sg13g2_decap_8 FILLER_4_1318 ();
 sg13g2_fill_1 FILLER_4_1325 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_4 FILLER_5_14 ();
 sg13g2_fill_1 FILLER_5_18 ();
 sg13g2_fill_1 FILLER_5_22 ();
 sg13g2_fill_1 FILLER_5_27 ();
 sg13g2_fill_1 FILLER_5_32 ();
 sg13g2_fill_1 FILLER_5_41 ();
 sg13g2_fill_2 FILLER_5_66 ();
 sg13g2_fill_1 FILLER_5_104 ();
 sg13g2_fill_2 FILLER_5_113 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_131 ();
 sg13g2_fill_2 FILLER_5_140 ();
 sg13g2_fill_2 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_fill_1 FILLER_5_193 ();
 sg13g2_decap_4 FILLER_5_197 ();
 sg13g2_fill_2 FILLER_5_201 ();
 sg13g2_fill_1 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_226 ();
 sg13g2_fill_1 FILLER_5_233 ();
 sg13g2_fill_2 FILLER_5_252 ();
 sg13g2_fill_2 FILLER_5_298 ();
 sg13g2_fill_1 FILLER_5_304 ();
 sg13g2_decap_4 FILLER_5_331 ();
 sg13g2_fill_1 FILLER_5_335 ();
 sg13g2_fill_2 FILLER_5_346 ();
 sg13g2_fill_1 FILLER_5_356 ();
 sg13g2_fill_1 FILLER_5_361 ();
 sg13g2_fill_1 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_fill_2 FILLER_5_397 ();
 sg13g2_fill_1 FILLER_5_409 ();
 sg13g2_fill_2 FILLER_5_415 ();
 sg13g2_fill_1 FILLER_5_417 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_decap_8 FILLER_5_429 ();
 sg13g2_fill_1 FILLER_5_436 ();
 sg13g2_fill_2 FILLER_5_442 ();
 sg13g2_fill_1 FILLER_5_444 ();
 sg13g2_fill_2 FILLER_5_449 ();
 sg13g2_fill_1 FILLER_5_451 ();
 sg13g2_decap_8 FILLER_5_482 ();
 sg13g2_decap_4 FILLER_5_489 ();
 sg13g2_fill_2 FILLER_5_493 ();
 sg13g2_fill_2 FILLER_5_499 ();
 sg13g2_fill_1 FILLER_5_501 ();
 sg13g2_decap_8 FILLER_5_505 ();
 sg13g2_decap_8 FILLER_5_512 ();
 sg13g2_decap_4 FILLER_5_519 ();
 sg13g2_fill_2 FILLER_5_523 ();
 sg13g2_decap_4 FILLER_5_530 ();
 sg13g2_fill_2 FILLER_5_547 ();
 sg13g2_fill_1 FILLER_5_549 ();
 sg13g2_fill_1 FILLER_5_554 ();
 sg13g2_fill_2 FILLER_5_560 ();
 sg13g2_decap_4 FILLER_5_622 ();
 sg13g2_fill_1 FILLER_5_626 ();
 sg13g2_fill_2 FILLER_5_632 ();
 sg13g2_decap_8 FILLER_5_638 ();
 sg13g2_fill_2 FILLER_5_645 ();
 sg13g2_fill_2 FILLER_5_658 ();
 sg13g2_fill_1 FILLER_5_660 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_fill_1 FILLER_5_686 ();
 sg13g2_fill_1 FILLER_5_691 ();
 sg13g2_fill_1 FILLER_5_696 ();
 sg13g2_decap_8 FILLER_5_701 ();
 sg13g2_fill_2 FILLER_5_708 ();
 sg13g2_fill_1 FILLER_5_719 ();
 sg13g2_decap_8 FILLER_5_724 ();
 sg13g2_decap_8 FILLER_5_731 ();
 sg13g2_fill_1 FILLER_5_742 ();
 sg13g2_fill_1 FILLER_5_747 ();
 sg13g2_fill_1 FILLER_5_753 ();
 sg13g2_fill_1 FILLER_5_758 ();
 sg13g2_fill_2 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_775 ();
 sg13g2_decap_8 FILLER_5_782 ();
 sg13g2_decap_4 FILLER_5_789 ();
 sg13g2_decap_4 FILLER_5_797 ();
 sg13g2_fill_1 FILLER_5_801 ();
 sg13g2_fill_2 FILLER_5_810 ();
 sg13g2_fill_2 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_fill_2 FILLER_5_851 ();
 sg13g2_fill_2 FILLER_5_879 ();
 sg13g2_fill_1 FILLER_5_881 ();
 sg13g2_fill_2 FILLER_5_918 ();
 sg13g2_fill_1 FILLER_5_920 ();
 sg13g2_decap_8 FILLER_5_925 ();
 sg13g2_decap_8 FILLER_5_932 ();
 sg13g2_decap_8 FILLER_5_939 ();
 sg13g2_fill_2 FILLER_5_946 ();
 sg13g2_fill_1 FILLER_5_948 ();
 sg13g2_fill_1 FILLER_5_979 ();
 sg13g2_fill_2 FILLER_5_985 ();
 sg13g2_fill_1 FILLER_5_987 ();
 sg13g2_fill_2 FILLER_5_1001 ();
 sg13g2_decap_4 FILLER_5_1013 ();
 sg13g2_fill_1 FILLER_5_1017 ();
 sg13g2_decap_8 FILLER_5_1022 ();
 sg13g2_fill_2 FILLER_5_1029 ();
 sg13g2_fill_1 FILLER_5_1061 ();
 sg13g2_decap_4 FILLER_5_1066 ();
 sg13g2_fill_1 FILLER_5_1070 ();
 sg13g2_fill_1 FILLER_5_1075 ();
 sg13g2_decap_8 FILLER_5_1110 ();
 sg13g2_fill_1 FILLER_5_1153 ();
 sg13g2_decap_4 FILLER_5_1180 ();
 sg13g2_fill_2 FILLER_5_1184 ();
 sg13g2_decap_8 FILLER_5_1212 ();
 sg13g2_decap_8 FILLER_5_1219 ();
 sg13g2_decap_8 FILLER_5_1226 ();
 sg13g2_decap_8 FILLER_5_1233 ();
 sg13g2_decap_8 FILLER_5_1240 ();
 sg13g2_decap_8 FILLER_5_1247 ();
 sg13g2_decap_8 FILLER_5_1254 ();
 sg13g2_decap_8 FILLER_5_1261 ();
 sg13g2_decap_8 FILLER_5_1268 ();
 sg13g2_decap_8 FILLER_5_1275 ();
 sg13g2_decap_8 FILLER_5_1282 ();
 sg13g2_decap_8 FILLER_5_1289 ();
 sg13g2_decap_8 FILLER_5_1296 ();
 sg13g2_decap_8 FILLER_5_1303 ();
 sg13g2_decap_8 FILLER_5_1310 ();
 sg13g2_decap_8 FILLER_5_1317 ();
 sg13g2_fill_2 FILLER_5_1324 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_17 ();
 sg13g2_fill_1 FILLER_6_27 ();
 sg13g2_fill_2 FILLER_6_32 ();
 sg13g2_decap_4 FILLER_6_43 ();
 sg13g2_fill_1 FILLER_6_51 ();
 sg13g2_fill_1 FILLER_6_56 ();
 sg13g2_fill_2 FILLER_6_62 ();
 sg13g2_fill_2 FILLER_6_68 ();
 sg13g2_fill_2 FILLER_6_91 ();
 sg13g2_fill_1 FILLER_6_93 ();
 sg13g2_fill_2 FILLER_6_97 ();
 sg13g2_fill_2 FILLER_6_104 ();
 sg13g2_fill_1 FILLER_6_116 ();
 sg13g2_fill_2 FILLER_6_122 ();
 sg13g2_fill_1 FILLER_6_124 ();
 sg13g2_decap_8 FILLER_6_134 ();
 sg13g2_decap_8 FILLER_6_141 ();
 sg13g2_decap_4 FILLER_6_148 ();
 sg13g2_fill_1 FILLER_6_152 ();
 sg13g2_decap_4 FILLER_6_156 ();
 sg13g2_fill_2 FILLER_6_164 ();
 sg13g2_fill_1 FILLER_6_166 ();
 sg13g2_fill_2 FILLER_6_205 ();
 sg13g2_fill_1 FILLER_6_207 ();
 sg13g2_fill_2 FILLER_6_226 ();
 sg13g2_fill_2 FILLER_6_239 ();
 sg13g2_fill_1 FILLER_6_241 ();
 sg13g2_decap_4 FILLER_6_252 ();
 sg13g2_fill_1 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_fill_2 FILLER_6_312 ();
 sg13g2_fill_1 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_4 FILLER_6_365 ();
 sg13g2_fill_1 FILLER_6_369 ();
 sg13g2_decap_4 FILLER_6_377 ();
 sg13g2_fill_2 FILLER_6_391 ();
 sg13g2_fill_1 FILLER_6_397 ();
 sg13g2_fill_1 FILLER_6_440 ();
 sg13g2_decap_4 FILLER_6_445 ();
 sg13g2_fill_2 FILLER_6_449 ();
 sg13g2_decap_4 FILLER_6_456 ();
 sg13g2_fill_1 FILLER_6_460 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_4 FILLER_6_473 ();
 sg13g2_decap_4 FILLER_6_481 ();
 sg13g2_decap_4 FILLER_6_489 ();
 sg13g2_fill_2 FILLER_6_493 ();
 sg13g2_fill_1 FILLER_6_512 ();
 sg13g2_fill_2 FILLER_6_539 ();
 sg13g2_fill_2 FILLER_6_575 ();
 sg13g2_fill_2 FILLER_6_580 ();
 sg13g2_decap_8 FILLER_6_613 ();
 sg13g2_fill_2 FILLER_6_620 ();
 sg13g2_fill_2 FILLER_6_684 ();
 sg13g2_fill_2 FILLER_6_698 ();
 sg13g2_fill_1 FILLER_6_700 ();
 sg13g2_fill_1 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_fill_1 FILLER_6_768 ();
 sg13g2_fill_2 FILLER_6_830 ();
 sg13g2_decap_4 FILLER_6_841 ();
 sg13g2_decap_8 FILLER_6_850 ();
 sg13g2_decap_4 FILLER_6_857 ();
 sg13g2_fill_2 FILLER_6_874 ();
 sg13g2_fill_1 FILLER_6_876 ();
 sg13g2_fill_1 FILLER_6_882 ();
 sg13g2_fill_2 FILLER_6_895 ();
 sg13g2_decap_8 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_940 ();
 sg13g2_decap_8 FILLER_6_947 ();
 sg13g2_fill_1 FILLER_6_954 ();
 sg13g2_decap_8 FILLER_6_959 ();
 sg13g2_decap_8 FILLER_6_966 ();
 sg13g2_decap_8 FILLER_6_973 ();
 sg13g2_decap_4 FILLER_6_980 ();
 sg13g2_fill_1 FILLER_6_984 ();
 sg13g2_fill_2 FILLER_6_1037 ();
 sg13g2_fill_1 FILLER_6_1039 ();
 sg13g2_decap_4 FILLER_6_1052 ();
 sg13g2_fill_1 FILLER_6_1056 ();
 sg13g2_decap_8 FILLER_6_1096 ();
 sg13g2_fill_1 FILLER_6_1103 ();
 sg13g2_decap_8 FILLER_6_1109 ();
 sg13g2_fill_1 FILLER_6_1116 ();
 sg13g2_fill_2 FILLER_6_1121 ();
 sg13g2_fill_1 FILLER_6_1131 ();
 sg13g2_decap_8 FILLER_6_1136 ();
 sg13g2_decap_8 FILLER_6_1143 ();
 sg13g2_decap_4 FILLER_6_1150 ();
 sg13g2_decap_8 FILLER_6_1164 ();
 sg13g2_decap_4 FILLER_6_1171 ();
 sg13g2_fill_2 FILLER_6_1175 ();
 sg13g2_decap_8 FILLER_6_1186 ();
 sg13g2_decap_8 FILLER_6_1231 ();
 sg13g2_fill_2 FILLER_6_1238 ();
 sg13g2_fill_1 FILLER_6_1240 ();
 sg13g2_decap_8 FILLER_6_1245 ();
 sg13g2_decap_8 FILLER_6_1252 ();
 sg13g2_decap_8 FILLER_6_1259 ();
 sg13g2_decap_8 FILLER_6_1266 ();
 sg13g2_decap_8 FILLER_6_1273 ();
 sg13g2_decap_8 FILLER_6_1280 ();
 sg13g2_decap_8 FILLER_6_1287 ();
 sg13g2_decap_8 FILLER_6_1294 ();
 sg13g2_decap_8 FILLER_6_1301 ();
 sg13g2_decap_8 FILLER_6_1308 ();
 sg13g2_decap_8 FILLER_6_1315 ();
 sg13g2_decap_4 FILLER_6_1322 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_19 ();
 sg13g2_fill_2 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_33 ();
 sg13g2_fill_2 FILLER_7_39 ();
 sg13g2_fill_2 FILLER_7_54 ();
 sg13g2_fill_2 FILLER_7_80 ();
 sg13g2_fill_2 FILLER_7_86 ();
 sg13g2_fill_1 FILLER_7_88 ();
 sg13g2_decap_8 FILLER_7_92 ();
 sg13g2_fill_1 FILLER_7_99 ();
 sg13g2_fill_1 FILLER_7_136 ();
 sg13g2_decap_8 FILLER_7_141 ();
 sg13g2_fill_1 FILLER_7_148 ();
 sg13g2_fill_2 FILLER_7_154 ();
 sg13g2_fill_1 FILLER_7_165 ();
 sg13g2_decap_8 FILLER_7_179 ();
 sg13g2_fill_2 FILLER_7_190 ();
 sg13g2_fill_2 FILLER_7_195 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_209 ();
 sg13g2_fill_1 FILLER_7_215 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_decap_8 FILLER_7_234 ();
 sg13g2_fill_2 FILLER_7_241 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_4 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_276 ();
 sg13g2_decap_4 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_fill_1 FILLER_7_334 ();
 sg13g2_decap_4 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_fill_1 FILLER_7_409 ();
 sg13g2_fill_1 FILLER_7_414 ();
 sg13g2_fill_2 FILLER_7_419 ();
 sg13g2_fill_2 FILLER_7_425 ();
 sg13g2_fill_1 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_433 ();
 sg13g2_fill_2 FILLER_7_460 ();
 sg13g2_decap_4 FILLER_7_488 ();
 sg13g2_fill_1 FILLER_7_492 ();
 sg13g2_decap_4 FILLER_7_523 ();
 sg13g2_fill_2 FILLER_7_530 ();
 sg13g2_decap_4 FILLER_7_537 ();
 sg13g2_decap_4 FILLER_7_546 ();
 sg13g2_fill_2 FILLER_7_550 ();
 sg13g2_fill_1 FILLER_7_575 ();
 sg13g2_fill_1 FILLER_7_581 ();
 sg13g2_fill_1 FILLER_7_586 ();
 sg13g2_fill_2 FILLER_7_603 ();
 sg13g2_decap_8 FILLER_7_634 ();
 sg13g2_decap_8 FILLER_7_641 ();
 sg13g2_fill_1 FILLER_7_648 ();
 sg13g2_decap_8 FILLER_7_657 ();
 sg13g2_fill_1 FILLER_7_664 ();
 sg13g2_decap_8 FILLER_7_669 ();
 sg13g2_fill_1 FILLER_7_702 ();
 sg13g2_fill_2 FILLER_7_708 ();
 sg13g2_fill_1 FILLER_7_710 ();
 sg13g2_decap_8 FILLER_7_741 ();
 sg13g2_decap_4 FILLER_7_752 ();
 sg13g2_fill_1 FILLER_7_756 ();
 sg13g2_fill_2 FILLER_7_776 ();
 sg13g2_decap_8 FILLER_7_782 ();
 sg13g2_decap_8 FILLER_7_789 ();
 sg13g2_decap_8 FILLER_7_796 ();
 sg13g2_decap_4 FILLER_7_803 ();
 sg13g2_fill_2 FILLER_7_871 ();
 sg13g2_fill_1 FILLER_7_873 ();
 sg13g2_fill_1 FILLER_7_879 ();
 sg13g2_fill_1 FILLER_7_906 ();
 sg13g2_fill_2 FILLER_7_933 ();
 sg13g2_decap_8 FILLER_7_939 ();
 sg13g2_fill_2 FILLER_7_946 ();
 sg13g2_fill_1 FILLER_7_978 ();
 sg13g2_decap_8 FILLER_7_988 ();
 sg13g2_decap_8 FILLER_7_995 ();
 sg13g2_fill_2 FILLER_7_1002 ();
 sg13g2_fill_1 FILLER_7_1004 ();
 sg13g2_decap_4 FILLER_7_1051 ();
 sg13g2_decap_8 FILLER_7_1059 ();
 sg13g2_decap_4 FILLER_7_1066 ();
 sg13g2_fill_1 FILLER_7_1070 ();
 sg13g2_decap_4 FILLER_7_1080 ();
 sg13g2_decap_8 FILLER_7_1088 ();
 sg13g2_fill_2 FILLER_7_1095 ();
 sg13g2_fill_2 FILLER_7_1132 ();
 sg13g2_fill_1 FILLER_7_1134 ();
 sg13g2_decap_8 FILLER_7_1143 ();
 sg13g2_fill_1 FILLER_7_1150 ();
 sg13g2_decap_8 FILLER_7_1206 ();
 sg13g2_fill_1 FILLER_7_1213 ();
 sg13g2_decap_4 FILLER_7_1228 ();
 sg13g2_fill_2 FILLER_7_1232 ();
 sg13g2_decap_8 FILLER_7_1260 ();
 sg13g2_decap_8 FILLER_7_1267 ();
 sg13g2_decap_8 FILLER_7_1274 ();
 sg13g2_decap_8 FILLER_7_1281 ();
 sg13g2_decap_8 FILLER_7_1288 ();
 sg13g2_decap_8 FILLER_7_1295 ();
 sg13g2_decap_8 FILLER_7_1302 ();
 sg13g2_decap_8 FILLER_7_1309 ();
 sg13g2_decap_8 FILLER_7_1316 ();
 sg13g2_fill_2 FILLER_7_1323 ();
 sg13g2_fill_1 FILLER_7_1325 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_4 FILLER_8_14 ();
 sg13g2_fill_1 FILLER_8_18 ();
 sg13g2_fill_1 FILLER_8_23 ();
 sg13g2_fill_2 FILLER_8_28 ();
 sg13g2_fill_2 FILLER_8_40 ();
 sg13g2_fill_1 FILLER_8_42 ();
 sg13g2_fill_2 FILLER_8_50 ();
 sg13g2_fill_2 FILLER_8_64 ();
 sg13g2_fill_1 FILLER_8_66 ();
 sg13g2_decap_8 FILLER_8_71 ();
 sg13g2_fill_1 FILLER_8_78 ();
 sg13g2_fill_1 FILLER_8_90 ();
 sg13g2_decap_8 FILLER_8_96 ();
 sg13g2_fill_1 FILLER_8_103 ();
 sg13g2_decap_4 FILLER_8_118 ();
 sg13g2_fill_2 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_131 ();
 sg13g2_decap_4 FILLER_8_136 ();
 sg13g2_fill_2 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_fill_2 FILLER_8_158 ();
 sg13g2_fill_1 FILLER_8_160 ();
 sg13g2_decap_8 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_195 ();
 sg13g2_fill_2 FILLER_8_204 ();
 sg13g2_fill_2 FILLER_8_211 ();
 sg13g2_fill_1 FILLER_8_213 ();
 sg13g2_decap_8 FILLER_8_219 ();
 sg13g2_fill_2 FILLER_8_226 ();
 sg13g2_fill_1 FILLER_8_246 ();
 sg13g2_fill_1 FILLER_8_263 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_297 ();
 sg13g2_fill_1 FILLER_8_299 ();
 sg13g2_decap_8 FILLER_8_304 ();
 sg13g2_decap_8 FILLER_8_311 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_320 ();
 sg13g2_decap_8 FILLER_8_325 ();
 sg13g2_decap_4 FILLER_8_332 ();
 sg13g2_fill_2 FILLER_8_339 ();
 sg13g2_decap_8 FILLER_8_353 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_fill_2 FILLER_8_381 ();
 sg13g2_fill_1 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_456 ();
 sg13g2_fill_1 FILLER_8_463 ();
 sg13g2_decap_4 FILLER_8_472 ();
 sg13g2_fill_1 FILLER_8_476 ();
 sg13g2_fill_2 FILLER_8_482 ();
 sg13g2_fill_1 FILLER_8_484 ();
 sg13g2_fill_1 FILLER_8_494 ();
 sg13g2_fill_2 FILLER_8_535 ();
 sg13g2_fill_1 FILLER_8_537 ();
 sg13g2_fill_2 FILLER_8_576 ();
 sg13g2_fill_2 FILLER_8_583 ();
 sg13g2_fill_1 FILLER_8_590 ();
 sg13g2_fill_1 FILLER_8_615 ();
 sg13g2_fill_1 FILLER_8_621 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_4 FILLER_8_704 ();
 sg13g2_fill_2 FILLER_8_708 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_fill_2 FILLER_8_735 ();
 sg13g2_fill_1 FILLER_8_737 ();
 sg13g2_decap_8 FILLER_8_765 ();
 sg13g2_fill_1 FILLER_8_777 ();
 sg13g2_decap_4 FILLER_8_783 ();
 sg13g2_decap_8 FILLER_8_813 ();
 sg13g2_fill_2 FILLER_8_820 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_fill_1 FILLER_8_833 ();
 sg13g2_decap_4 FILLER_8_839 ();
 sg13g2_fill_1 FILLER_8_843 ();
 sg13g2_decap_8 FILLER_8_848 ();
 sg13g2_fill_2 FILLER_8_855 ();
 sg13g2_fill_1 FILLER_8_857 ();
 sg13g2_fill_2 FILLER_8_887 ();
 sg13g2_decap_8 FILLER_8_919 ();
 sg13g2_fill_2 FILLER_8_926 ();
 sg13g2_fill_2 FILLER_8_958 ();
 sg13g2_fill_1 FILLER_8_960 ();
 sg13g2_fill_2 FILLER_8_965 ();
 sg13g2_fill_1 FILLER_8_977 ();
 sg13g2_fill_1 FILLER_8_1004 ();
 sg13g2_fill_1 FILLER_8_1031 ();
 sg13g2_fill_2 FILLER_8_1036 ();
 sg13g2_fill_2 FILLER_8_1074 ();
 sg13g2_fill_1 FILLER_8_1076 ();
 sg13g2_fill_1 FILLER_8_1115 ();
 sg13g2_fill_2 FILLER_8_1119 ();
 sg13g2_fill_1 FILLER_8_1121 ();
 sg13g2_fill_2 FILLER_8_1126 ();
 sg13g2_fill_1 FILLER_8_1154 ();
 sg13g2_fill_2 FILLER_8_1164 ();
 sg13g2_fill_1 FILLER_8_1166 ();
 sg13g2_decap_4 FILLER_8_1171 ();
 sg13g2_decap_4 FILLER_8_1180 ();
 sg13g2_decap_8 FILLER_8_1188 ();
 sg13g2_fill_1 FILLER_8_1195 ();
 sg13g2_fill_2 FILLER_8_1236 ();
 sg13g2_fill_1 FILLER_8_1238 ();
 sg13g2_decap_4 FILLER_8_1248 ();
 sg13g2_fill_1 FILLER_8_1252 ();
 sg13g2_fill_1 FILLER_8_1263 ();
 sg13g2_decap_8 FILLER_8_1300 ();
 sg13g2_decap_8 FILLER_8_1307 ();
 sg13g2_decap_8 FILLER_8_1314 ();
 sg13g2_decap_4 FILLER_8_1321 ();
 sg13g2_fill_1 FILLER_8_1325 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_29 ();
 sg13g2_fill_1 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_41 ();
 sg13g2_fill_1 FILLER_9_47 ();
 sg13g2_fill_2 FILLER_9_57 ();
 sg13g2_fill_1 FILLER_9_59 ();
 sg13g2_fill_2 FILLER_9_84 ();
 sg13g2_fill_2 FILLER_9_92 ();
 sg13g2_fill_2 FILLER_9_98 ();
 sg13g2_fill_1 FILLER_9_100 ();
 sg13g2_fill_2 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_107 ();
 sg13g2_fill_2 FILLER_9_113 ();
 sg13g2_fill_2 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_153 ();
 sg13g2_fill_1 FILLER_9_160 ();
 sg13g2_fill_1 FILLER_9_165 ();
 sg13g2_fill_1 FILLER_9_192 ();
 sg13g2_fill_2 FILLER_9_219 ();
 sg13g2_fill_1 FILLER_9_226 ();
 sg13g2_fill_2 FILLER_9_235 ();
 sg13g2_fill_1 FILLER_9_313 ();
 sg13g2_fill_2 FILLER_9_340 ();
 sg13g2_fill_1 FILLER_9_342 ();
 sg13g2_fill_2 FILLER_9_403 ();
 sg13g2_decap_4 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_431 ();
 sg13g2_decap_8 FILLER_9_436 ();
 sg13g2_fill_1 FILLER_9_443 ();
 sg13g2_fill_1 FILLER_9_449 ();
 sg13g2_fill_1 FILLER_9_476 ();
 sg13g2_fill_1 FILLER_9_482 ();
 sg13g2_fill_2 FILLER_9_488 ();
 sg13g2_decap_4 FILLER_9_495 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_515 ();
 sg13g2_fill_2 FILLER_9_535 ();
 sg13g2_fill_1 FILLER_9_537 ();
 sg13g2_fill_2 FILLER_9_561 ();
 sg13g2_fill_1 FILLER_9_563 ();
 sg13g2_fill_1 FILLER_9_590 ();
 sg13g2_fill_2 FILLER_9_599 ();
 sg13g2_fill_2 FILLER_9_621 ();
 sg13g2_fill_1 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_627 ();
 sg13g2_fill_2 FILLER_9_634 ();
 sg13g2_decap_8 FILLER_9_640 ();
 sg13g2_fill_2 FILLER_9_647 ();
 sg13g2_fill_2 FILLER_9_657 ();
 sg13g2_fill_1 FILLER_9_659 ();
 sg13g2_decap_8 FILLER_9_664 ();
 sg13g2_decap_4 FILLER_9_671 ();
 sg13g2_decap_4 FILLER_9_679 ();
 sg13g2_fill_1 FILLER_9_683 ();
 sg13g2_fill_2 FILLER_9_746 ();
 sg13g2_decap_4 FILLER_9_769 ();
 sg13g2_fill_2 FILLER_9_773 ();
 sg13g2_fill_2 FILLER_9_784 ();
 sg13g2_fill_1 FILLER_9_790 ();
 sg13g2_fill_1 FILLER_9_796 ();
 sg13g2_fill_2 FILLER_9_801 ();
 sg13g2_decap_4 FILLER_9_848 ();
 sg13g2_fill_2 FILLER_9_852 ();
 sg13g2_fill_2 FILLER_9_863 ();
 sg13g2_fill_1 FILLER_9_865 ();
 sg13g2_fill_2 FILLER_9_870 ();
 sg13g2_fill_2 FILLER_9_898 ();
 sg13g2_decap_4 FILLER_9_926 ();
 sg13g2_fill_2 FILLER_9_930 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_1018 ();
 sg13g2_fill_2 FILLER_9_1025 ();
 sg13g2_decap_8 FILLER_9_1045 ();
 sg13g2_decap_4 FILLER_9_1052 ();
 sg13g2_fill_2 FILLER_9_1056 ();
 sg13g2_decap_8 FILLER_9_1067 ();
 sg13g2_fill_2 FILLER_9_1074 ();
 sg13g2_decap_4 FILLER_9_1084 ();
 sg13g2_fill_2 FILLER_9_1088 ();
 sg13g2_fill_2 FILLER_9_1131 ();
 sg13g2_fill_1 FILLER_9_1133 ();
 sg13g2_fill_2 FILLER_9_1151 ();
 sg13g2_fill_1 FILLER_9_1153 ();
 sg13g2_decap_8 FILLER_9_1184 ();
 sg13g2_decap_8 FILLER_9_1191 ();
 sg13g2_decap_4 FILLER_9_1198 ();
 sg13g2_fill_1 FILLER_9_1202 ();
 sg13g2_decap_4 FILLER_9_1207 ();
 sg13g2_fill_1 FILLER_9_1234 ();
 sg13g2_decap_8 FILLER_9_1291 ();
 sg13g2_decap_8 FILLER_9_1298 ();
 sg13g2_decap_8 FILLER_9_1305 ();
 sg13g2_decap_8 FILLER_9_1312 ();
 sg13g2_decap_8 FILLER_9_1319 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_14 ();
 sg13g2_fill_1 FILLER_10_27 ();
 sg13g2_fill_2 FILLER_10_39 ();
 sg13g2_fill_1 FILLER_10_45 ();
 sg13g2_fill_1 FILLER_10_50 ();
 sg13g2_fill_2 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_84 ();
 sg13g2_fill_1 FILLER_10_86 ();
 sg13g2_fill_2 FILLER_10_138 ();
 sg13g2_decap_8 FILLER_10_170 ();
 sg13g2_decap_8 FILLER_10_177 ();
 sg13g2_decap_8 FILLER_10_184 ();
 sg13g2_fill_2 FILLER_10_191 ();
 sg13g2_decap_4 FILLER_10_197 ();
 sg13g2_fill_1 FILLER_10_201 ();
 sg13g2_decap_8 FILLER_10_206 ();
 sg13g2_decap_4 FILLER_10_218 ();
 sg13g2_fill_1 FILLER_10_222 ();
 sg13g2_fill_2 FILLER_10_228 ();
 sg13g2_fill_1 FILLER_10_230 ();
 sg13g2_fill_2 FILLER_10_239 ();
 sg13g2_fill_1 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_246 ();
 sg13g2_fill_1 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_273 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_fill_1 FILLER_10_312 ();
 sg13g2_fill_2 FILLER_10_343 ();
 sg13g2_fill_2 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_fill_2 FILLER_10_363 ();
 sg13g2_fill_2 FILLER_10_370 ();
 sg13g2_decap_4 FILLER_10_379 ();
 sg13g2_fill_1 FILLER_10_383 ();
 sg13g2_decap_4 FILLER_10_392 ();
 sg13g2_fill_1 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_432 ();
 sg13g2_decap_8 FILLER_10_439 ();
 sg13g2_fill_2 FILLER_10_457 ();
 sg13g2_decap_4 FILLER_10_463 ();
 sg13g2_fill_2 FILLER_10_467 ();
 sg13g2_fill_1 FILLER_10_524 ();
 sg13g2_fill_2 FILLER_10_529 ();
 sg13g2_fill_1 FILLER_10_531 ();
 sg13g2_fill_1 FILLER_10_548 ();
 sg13g2_fill_1 FILLER_10_575 ();
 sg13g2_fill_1 FILLER_10_581 ();
 sg13g2_fill_1 FILLER_10_608 ();
 sg13g2_fill_1 FILLER_10_614 ();
 sg13g2_fill_2 FILLER_10_641 ();
 sg13g2_fill_2 FILLER_10_648 ();
 sg13g2_fill_2 FILLER_10_653 ();
 sg13g2_decap_8 FILLER_10_659 ();
 sg13g2_fill_1 FILLER_10_692 ();
 sg13g2_fill_2 FILLER_10_697 ();
 sg13g2_fill_2 FILLER_10_703 ();
 sg13g2_fill_2 FILLER_10_710 ();
 sg13g2_fill_1 FILLER_10_712 ();
 sg13g2_fill_2 FILLER_10_716 ();
 sg13g2_fill_1 FILLER_10_727 ();
 sg13g2_decap_4 FILLER_10_732 ();
 sg13g2_fill_1 FILLER_10_781 ();
 sg13g2_fill_1 FILLER_10_787 ();
 sg13g2_fill_1 FILLER_10_795 ();
 sg13g2_decap_4 FILLER_10_804 ();
 sg13g2_fill_1 FILLER_10_808 ();
 sg13g2_decap_4 FILLER_10_854 ();
 sg13g2_fill_2 FILLER_10_862 ();
 sg13g2_fill_1 FILLER_10_864 ();
 sg13g2_decap_8 FILLER_10_869 ();
 sg13g2_fill_1 FILLER_10_876 ();
 sg13g2_decap_8 FILLER_10_881 ();
 sg13g2_fill_2 FILLER_10_888 ();
 sg13g2_decap_8 FILLER_10_893 ();
 sg13g2_decap_4 FILLER_10_900 ();
 sg13g2_fill_1 FILLER_10_904 ();
 sg13g2_decap_8 FILLER_10_944 ();
 sg13g2_decap_4 FILLER_10_951 ();
 sg13g2_decap_4 FILLER_10_960 ();
 sg13g2_fill_2 FILLER_10_964 ();
 sg13g2_decap_4 FILLER_10_975 ();
 sg13g2_fill_1 FILLER_10_1005 ();
 sg13g2_fill_2 FILLER_10_1110 ();
 sg13g2_fill_1 FILLER_10_1169 ();
 sg13g2_fill_1 FILLER_10_1174 ();
 sg13g2_fill_1 FILLER_10_1237 ();
 sg13g2_decap_8 FILLER_10_1251 ();
 sg13g2_decap_8 FILLER_10_1258 ();
 sg13g2_fill_2 FILLER_10_1265 ();
 sg13g2_decap_8 FILLER_10_1271 ();
 sg13g2_decap_8 FILLER_10_1278 ();
 sg13g2_fill_1 FILLER_10_1285 ();
 sg13g2_decap_4 FILLER_10_1322 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_25 ();
 sg13g2_fill_1 FILLER_11_27 ();
 sg13g2_fill_2 FILLER_11_41 ();
 sg13g2_fill_1 FILLER_11_43 ();
 sg13g2_fill_1 FILLER_11_52 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_fill_2 FILLER_11_76 ();
 sg13g2_fill_1 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_96 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_fill_1 FILLER_11_117 ();
 sg13g2_fill_1 FILLER_11_137 ();
 sg13g2_decap_4 FILLER_11_143 ();
 sg13g2_fill_2 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_153 ();
 sg13g2_decap_8 FILLER_11_160 ();
 sg13g2_decap_8 FILLER_11_167 ();
 sg13g2_decap_8 FILLER_11_174 ();
 sg13g2_decap_4 FILLER_11_181 ();
 sg13g2_fill_1 FILLER_11_185 ();
 sg13g2_decap_8 FILLER_11_201 ();
 sg13g2_fill_2 FILLER_11_208 ();
 sg13g2_fill_1 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_216 ();
 sg13g2_fill_1 FILLER_11_223 ();
 sg13g2_fill_2 FILLER_11_243 ();
 sg13g2_fill_1 FILLER_11_245 ();
 sg13g2_decap_4 FILLER_11_264 ();
 sg13g2_fill_2 FILLER_11_268 ();
 sg13g2_fill_1 FILLER_11_307 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_4 FILLER_11_319 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_decap_8 FILLER_11_332 ();
 sg13g2_fill_2 FILLER_11_355 ();
 sg13g2_decap_4 FILLER_11_362 ();
 sg13g2_fill_2 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_372 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_4 FILLER_11_393 ();
 sg13g2_fill_1 FILLER_11_397 ();
 sg13g2_fill_2 FILLER_11_405 ();
 sg13g2_fill_1 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_11_412 ();
 sg13g2_fill_2 FILLER_11_419 ();
 sg13g2_fill_1 FILLER_11_421 ();
 sg13g2_decap_8 FILLER_11_468 ();
 sg13g2_fill_1 FILLER_11_475 ();
 sg13g2_fill_2 FILLER_11_485 ();
 sg13g2_fill_1 FILLER_11_506 ();
 sg13g2_fill_2 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_544 ();
 sg13g2_fill_1 FILLER_11_592 ();
 sg13g2_decap_8 FILLER_11_601 ();
 sg13g2_decap_4 FILLER_11_608 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_fill_1 FILLER_11_637 ();
 sg13g2_decap_4 FILLER_11_674 ();
 sg13g2_fill_2 FILLER_11_678 ();
 sg13g2_decap_8 FILLER_11_684 ();
 sg13g2_fill_2 FILLER_11_691 ();
 sg13g2_fill_1 FILLER_11_693 ();
 sg13g2_decap_4 FILLER_11_708 ();
 sg13g2_decap_4 FILLER_11_717 ();
 sg13g2_decap_8 FILLER_11_726 ();
 sg13g2_decap_8 FILLER_11_733 ();
 sg13g2_fill_2 FILLER_11_753 ();
 sg13g2_fill_1 FILLER_11_759 ();
 sg13g2_decap_8 FILLER_11_764 ();
 sg13g2_fill_2 FILLER_11_771 ();
 sg13g2_fill_1 FILLER_11_773 ();
 sg13g2_decap_8 FILLER_11_778 ();
 sg13g2_decap_4 FILLER_11_785 ();
 sg13g2_decap_4 FILLER_11_815 ();
 sg13g2_fill_1 FILLER_11_829 ();
 sg13g2_decap_8 FILLER_11_834 ();
 sg13g2_decap_8 FILLER_11_841 ();
 sg13g2_fill_1 FILLER_11_848 ();
 sg13g2_decap_8 FILLER_11_896 ();
 sg13g2_fill_1 FILLER_11_915 ();
 sg13g2_decap_4 FILLER_11_920 ();
 sg13g2_decap_4 FILLER_11_993 ();
 sg13g2_fill_2 FILLER_11_997 ();
 sg13g2_decap_8 FILLER_11_1003 ();
 sg13g2_fill_2 FILLER_11_1010 ();
 sg13g2_decap_4 FILLER_11_1016 ();
 sg13g2_fill_2 FILLER_11_1020 ();
 sg13g2_decap_4 FILLER_11_1026 ();
 sg13g2_decap_4 FILLER_11_1034 ();
 sg13g2_fill_1 FILLER_11_1038 ();
 sg13g2_fill_2 FILLER_11_1043 ();
 sg13g2_decap_8 FILLER_11_1058 ();
 sg13g2_fill_1 FILLER_11_1065 ();
 sg13g2_decap_8 FILLER_11_1070 ();
 sg13g2_fill_1 FILLER_11_1077 ();
 sg13g2_decap_8 FILLER_11_1082 ();
 sg13g2_decap_4 FILLER_11_1089 ();
 sg13g2_decap_8 FILLER_11_1137 ();
 sg13g2_fill_2 FILLER_11_1148 ();
 sg13g2_fill_2 FILLER_11_1160 ();
 sg13g2_fill_1 FILLER_11_1175 ();
 sg13g2_decap_8 FILLER_11_1179 ();
 sg13g2_decap_4 FILLER_11_1186 ();
 sg13g2_fill_1 FILLER_11_1190 ();
 sg13g2_decap_8 FILLER_11_1195 ();
 sg13g2_decap_8 FILLER_11_1202 ();
 sg13g2_decap_8 FILLER_11_1209 ();
 sg13g2_fill_1 FILLER_11_1216 ();
 sg13g2_fill_2 FILLER_11_1221 ();
 sg13g2_fill_1 FILLER_11_1223 ();
 sg13g2_decap_4 FILLER_11_1234 ();
 sg13g2_fill_1 FILLER_11_1238 ();
 sg13g2_decap_4 FILLER_11_1265 ();
 sg13g2_fill_2 FILLER_11_1269 ();
 sg13g2_decap_8 FILLER_11_1275 ();
 sg13g2_decap_8 FILLER_11_1282 ();
 sg13g2_decap_8 FILLER_11_1289 ();
 sg13g2_decap_8 FILLER_11_1296 ();
 sg13g2_decap_8 FILLER_11_1311 ();
 sg13g2_decap_8 FILLER_11_1318 ();
 sg13g2_fill_1 FILLER_11_1325 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_11 ();
 sg13g2_fill_1 FILLER_12_32 ();
 sg13g2_fill_1 FILLER_12_50 ();
 sg13g2_decap_4 FILLER_12_55 ();
 sg13g2_fill_2 FILLER_12_92 ();
 sg13g2_fill_1 FILLER_12_102 ();
 sg13g2_fill_2 FILLER_12_108 ();
 sg13g2_decap_4 FILLER_12_114 ();
 sg13g2_fill_2 FILLER_12_118 ();
 sg13g2_decap_8 FILLER_12_125 ();
 sg13g2_decap_8 FILLER_12_132 ();
 sg13g2_fill_2 FILLER_12_139 ();
 sg13g2_fill_1 FILLER_12_141 ();
 sg13g2_fill_2 FILLER_12_168 ();
 sg13g2_fill_1 FILLER_12_170 ();
 sg13g2_fill_1 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_fill_1 FILLER_12_205 ();
 sg13g2_fill_2 FILLER_12_211 ();
 sg13g2_fill_2 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_258 ();
 sg13g2_decap_8 FILLER_12_265 ();
 sg13g2_decap_8 FILLER_12_272 ();
 sg13g2_decap_4 FILLER_12_279 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_4 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_319 ();
 sg13g2_fill_1 FILLER_12_360 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_decap_4 FILLER_12_453 ();
 sg13g2_fill_2 FILLER_12_457 ();
 sg13g2_fill_2 FILLER_12_488 ();
 sg13g2_decap_8 FILLER_12_521 ();
 sg13g2_decap_4 FILLER_12_528 ();
 sg13g2_decap_8 FILLER_12_535 ();
 sg13g2_decap_8 FILLER_12_542 ();
 sg13g2_fill_2 FILLER_12_549 ();
 sg13g2_fill_1 FILLER_12_551 ();
 sg13g2_decap_4 FILLER_12_559 ();
 sg13g2_fill_1 FILLER_12_563 ();
 sg13g2_fill_2 FILLER_12_568 ();
 sg13g2_decap_4 FILLER_12_574 ();
 sg13g2_fill_2 FILLER_12_583 ();
 sg13g2_fill_1 FILLER_12_585 ();
 sg13g2_decap_4 FILLER_12_594 ();
 sg13g2_decap_8 FILLER_12_603 ();
 sg13g2_fill_2 FILLER_12_610 ();
 sg13g2_fill_1 FILLER_12_672 ();
 sg13g2_fill_2 FILLER_12_699 ();
 sg13g2_fill_1 FILLER_12_701 ();
 sg13g2_fill_2 FILLER_12_754 ();
 sg13g2_fill_2 FILLER_12_761 ();
 sg13g2_fill_1 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_768 ();
 sg13g2_fill_1 FILLER_12_775 ();
 sg13g2_decap_4 FILLER_12_780 ();
 sg13g2_fill_2 FILLER_12_789 ();
 sg13g2_fill_2 FILLER_12_822 ();
 sg13g2_fill_1 FILLER_12_824 ();
 sg13g2_fill_1 FILLER_12_864 ();
 sg13g2_fill_2 FILLER_12_881 ();
 sg13g2_fill_1 FILLER_12_923 ();
 sg13g2_fill_2 FILLER_12_939 ();
 sg13g2_decap_8 FILLER_12_945 ();
 sg13g2_decap_4 FILLER_12_952 ();
 sg13g2_fill_1 FILLER_12_956 ();
 sg13g2_fill_2 FILLER_12_966 ();
 sg13g2_fill_1 FILLER_12_968 ();
 sg13g2_decap_8 FILLER_12_973 ();
 sg13g2_decap_4 FILLER_12_1016 ();
 sg13g2_fill_1 FILLER_12_1020 ();
 sg13g2_fill_2 FILLER_12_1075 ();
 sg13g2_fill_1 FILLER_12_1077 ();
 sg13g2_decap_4 FILLER_12_1114 ();
 sg13g2_fill_1 FILLER_12_1118 ();
 sg13g2_fill_2 FILLER_12_1129 ();
 sg13g2_decap_8 FILLER_12_1187 ();
 sg13g2_decap_8 FILLER_12_1194 ();
 sg13g2_fill_2 FILLER_12_1205 ();
 sg13g2_fill_2 FILLER_12_1233 ();
 sg13g2_fill_1 FILLER_12_1235 ();
 sg13g2_fill_2 FILLER_12_1244 ();
 sg13g2_fill_1 FILLER_12_1246 ();
 sg13g2_fill_2 FILLER_12_1251 ();
 sg13g2_fill_1 FILLER_12_1253 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_38 ();
 sg13g2_fill_2 FILLER_13_44 ();
 sg13g2_decap_4 FILLER_13_69 ();
 sg13g2_fill_2 FILLER_13_73 ();
 sg13g2_fill_2 FILLER_13_88 ();
 sg13g2_fill_1 FILLER_13_90 ();
 sg13g2_decap_4 FILLER_13_95 ();
 sg13g2_fill_2 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_127 ();
 sg13g2_fill_1 FILLER_13_132 ();
 sg13g2_decap_4 FILLER_13_137 ();
 sg13g2_fill_2 FILLER_13_141 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_fill_2 FILLER_13_154 ();
 sg13g2_fill_1 FILLER_13_156 ();
 sg13g2_decap_8 FILLER_13_170 ();
 sg13g2_decap_4 FILLER_13_177 ();
 sg13g2_fill_1 FILLER_13_192 ();
 sg13g2_decap_4 FILLER_13_199 ();
 sg13g2_fill_2 FILLER_13_203 ();
 sg13g2_fill_1 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_233 ();
 sg13g2_fill_1 FILLER_13_240 ();
 sg13g2_decap_8 FILLER_13_244 ();
 sg13g2_fill_2 FILLER_13_251 ();
 sg13g2_fill_1 FILLER_13_253 ();
 sg13g2_fill_2 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_270 ();
 sg13g2_fill_2 FILLER_13_290 ();
 sg13g2_fill_2 FILLER_13_297 ();
 sg13g2_fill_1 FILLER_13_299 ();
 sg13g2_decap_4 FILLER_13_326 ();
 sg13g2_decap_4 FILLER_13_366 ();
 sg13g2_fill_1 FILLER_13_370 ();
 sg13g2_fill_2 FILLER_13_375 ();
 sg13g2_fill_1 FILLER_13_377 ();
 sg13g2_decap_4 FILLER_13_382 ();
 sg13g2_fill_1 FILLER_13_430 ();
 sg13g2_decap_8 FILLER_13_435 ();
 sg13g2_fill_1 FILLER_13_442 ();
 sg13g2_decap_8 FILLER_13_446 ();
 sg13g2_decap_8 FILLER_13_453 ();
 sg13g2_decap_8 FILLER_13_460 ();
 sg13g2_fill_2 FILLER_13_467 ();
 sg13g2_fill_1 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_474 ();
 sg13g2_decap_8 FILLER_13_481 ();
 sg13g2_fill_1 FILLER_13_488 ();
 sg13g2_fill_2 FILLER_13_513 ();
 sg13g2_fill_1 FILLER_13_515 ();
 sg13g2_fill_1 FILLER_13_546 ();
 sg13g2_fill_2 FILLER_13_573 ();
 sg13g2_fill_2 FILLER_13_584 ();
 sg13g2_fill_1 FILLER_13_586 ();
 sg13g2_fill_2 FILLER_13_624 ();
 sg13g2_fill_1 FILLER_13_626 ();
 sg13g2_fill_1 FILLER_13_637 ();
 sg13g2_fill_1 FILLER_13_643 ();
 sg13g2_fill_1 FILLER_13_653 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_4 FILLER_13_693 ();
 sg13g2_fill_2 FILLER_13_697 ();
 sg13g2_decap_8 FILLER_13_703 ();
 sg13g2_fill_1 FILLER_13_710 ();
 sg13g2_decap_8 FILLER_13_715 ();
 sg13g2_decap_4 FILLER_13_722 ();
 sg13g2_decap_4 FILLER_13_730 ();
 sg13g2_fill_1 FILLER_13_734 ();
 sg13g2_fill_1 FILLER_13_739 ();
 sg13g2_fill_2 FILLER_13_745 ();
 sg13g2_fill_1 FILLER_13_757 ();
 sg13g2_decap_4 FILLER_13_788 ();
 sg13g2_fill_1 FILLER_13_792 ();
 sg13g2_fill_1 FILLER_13_797 ();
 sg13g2_fill_2 FILLER_13_802 ();
 sg13g2_fill_2 FILLER_13_808 ();
 sg13g2_fill_2 FILLER_13_814 ();
 sg13g2_decap_4 FILLER_13_826 ();
 sg13g2_fill_2 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_836 ();
 sg13g2_fill_2 FILLER_13_843 ();
 sg13g2_fill_1 FILLER_13_845 ();
 sg13g2_fill_2 FILLER_13_868 ();
 sg13g2_fill_1 FILLER_13_870 ();
 sg13g2_fill_2 FILLER_13_876 ();
 sg13g2_decap_4 FILLER_13_888 ();
 sg13g2_fill_2 FILLER_13_892 ();
 sg13g2_decap_4 FILLER_13_898 ();
 sg13g2_fill_1 FILLER_13_902 ();
 sg13g2_fill_1 FILLER_13_929 ();
 sg13g2_fill_2 FILLER_13_956 ();
 sg13g2_fill_1 FILLER_13_958 ();
 sg13g2_fill_1 FILLER_13_989 ();
 sg13g2_decap_8 FILLER_13_1025 ();
 sg13g2_fill_2 FILLER_13_1032 ();
 sg13g2_fill_2 FILLER_13_1056 ();
 sg13g2_fill_1 FILLER_13_1058 ();
 sg13g2_decap_4 FILLER_13_1088 ();
 sg13g2_fill_1 FILLER_13_1092 ();
 sg13g2_decap_8 FILLER_13_1097 ();
 sg13g2_decap_8 FILLER_13_1104 ();
 sg13g2_decap_8 FILLER_13_1111 ();
 sg13g2_fill_1 FILLER_13_1118 ();
 sg13g2_decap_4 FILLER_13_1129 ();
 sg13g2_fill_2 FILLER_13_1133 ();
 sg13g2_decap_4 FILLER_13_1155 ();
 sg13g2_fill_2 FILLER_13_1163 ();
 sg13g2_fill_2 FILLER_13_1191 ();
 sg13g2_fill_1 FILLER_13_1193 ();
 sg13g2_fill_1 FILLER_13_1220 ();
 sg13g2_decap_4 FILLER_13_1225 ();
 sg13g2_fill_1 FILLER_13_1229 ();
 sg13g2_fill_2 FILLER_13_1239 ();
 sg13g2_fill_1 FILLER_13_1246 ();
 sg13g2_decap_4 FILLER_13_1251 ();
 sg13g2_fill_2 FILLER_13_1259 ();
 sg13g2_fill_1 FILLER_13_1264 ();
 sg13g2_fill_1 FILLER_13_1287 ();
 sg13g2_fill_2 FILLER_13_1324 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_fill_2 FILLER_14_40 ();
 sg13g2_decap_8 FILLER_14_48 ();
 sg13g2_decap_4 FILLER_14_55 ();
 sg13g2_fill_2 FILLER_14_69 ();
 sg13g2_fill_1 FILLER_14_71 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_88 ();
 sg13g2_decap_8 FILLER_14_93 ();
 sg13g2_decap_8 FILLER_14_100 ();
 sg13g2_decap_4 FILLER_14_107 ();
 sg13g2_fill_2 FILLER_14_111 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_decap_4 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_decap_8 FILLER_14_145 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_215 ();
 sg13g2_fill_2 FILLER_14_280 ();
 sg13g2_fill_1 FILLER_14_287 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_304 ();
 sg13g2_fill_1 FILLER_14_306 ();
 sg13g2_decap_4 FILLER_14_333 ();
 sg13g2_fill_1 FILLER_14_349 ();
 sg13g2_decap_8 FILLER_14_353 ();
 sg13g2_decap_4 FILLER_14_360 ();
 sg13g2_fill_2 FILLER_14_413 ();
 sg13g2_fill_1 FILLER_14_415 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_1 FILLER_14_433 ();
 sg13g2_fill_2 FILLER_14_492 ();
 sg13g2_fill_1 FILLER_14_523 ();
 sg13g2_decap_4 FILLER_14_529 ();
 sg13g2_decap_8 FILLER_14_542 ();
 sg13g2_fill_1 FILLER_14_549 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_fill_2 FILLER_14_560 ();
 sg13g2_fill_1 FILLER_14_562 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_fill_1 FILLER_14_574 ();
 sg13g2_fill_2 FILLER_14_579 ();
 sg13g2_fill_1 FILLER_14_594 ();
 sg13g2_fill_1 FILLER_14_599 ();
 sg13g2_fill_2 FILLER_14_671 ();
 sg13g2_fill_1 FILLER_14_673 ();
 sg13g2_decap_8 FILLER_14_678 ();
 sg13g2_fill_1 FILLER_14_685 ();
 sg13g2_fill_1 FILLER_14_726 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_746 ();
 sg13g2_fill_2 FILLER_14_753 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_fill_1 FILLER_14_784 ();
 sg13g2_fill_2 FILLER_14_816 ();
 sg13g2_fill_1 FILLER_14_822 ();
 sg13g2_fill_2 FILLER_14_857 ();
 sg13g2_fill_1 FILLER_14_859 ();
 sg13g2_fill_1 FILLER_14_912 ();
 sg13g2_decap_4 FILLER_14_917 ();
 sg13g2_fill_1 FILLER_14_921 ();
 sg13g2_decap_4 FILLER_14_931 ();
 sg13g2_fill_2 FILLER_14_935 ();
 sg13g2_decap_8 FILLER_14_941 ();
 sg13g2_decap_8 FILLER_14_948 ();
 sg13g2_decap_4 FILLER_14_955 ();
 sg13g2_fill_1 FILLER_14_959 ();
 sg13g2_decap_8 FILLER_14_996 ();
 sg13g2_decap_8 FILLER_14_1003 ();
 sg13g2_decap_4 FILLER_14_1013 ();
 sg13g2_decap_8 FILLER_14_1030 ();
 sg13g2_fill_2 FILLER_14_1037 ();
 sg13g2_fill_1 FILLER_14_1039 ();
 sg13g2_fill_2 FILLER_14_1066 ();
 sg13g2_fill_1 FILLER_14_1068 ();
 sg13g2_fill_2 FILLER_14_1073 ();
 sg13g2_fill_2 FILLER_14_1084 ();
 sg13g2_fill_1 FILLER_14_1086 ();
 sg13g2_fill_2 FILLER_14_1092 ();
 sg13g2_fill_1 FILLER_14_1094 ();
 sg13g2_decap_8 FILLER_14_1151 ();
 sg13g2_fill_1 FILLER_14_1158 ();
 sg13g2_fill_1 FILLER_14_1180 ();
 sg13g2_decap_8 FILLER_14_1191 ();
 sg13g2_fill_2 FILLER_14_1198 ();
 sg13g2_decap_4 FILLER_14_1203 ();
 sg13g2_fill_2 FILLER_14_1207 ();
 sg13g2_decap_4 FILLER_14_1213 ();
 sg13g2_fill_1 FILLER_14_1221 ();
 sg13g2_fill_1 FILLER_14_1227 ();
 sg13g2_fill_2 FILLER_14_1233 ();
 sg13g2_fill_1 FILLER_14_1239 ();
 sg13g2_fill_2 FILLER_14_1266 ();
 sg13g2_decap_8 FILLER_14_1294 ();
 sg13g2_fill_2 FILLER_14_1301 ();
 sg13g2_fill_1 FILLER_14_1303 ();
 sg13g2_decap_8 FILLER_14_1312 ();
 sg13g2_decap_8 FILLER_14_1319 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_23 ();
 sg13g2_fill_1 FILLER_15_25 ();
 sg13g2_decap_4 FILLER_15_31 ();
 sg13g2_decap_8 FILLER_15_43 ();
 sg13g2_decap_8 FILLER_15_50 ();
 sg13g2_decap_8 FILLER_15_65 ();
 sg13g2_decap_8 FILLER_15_72 ();
 sg13g2_fill_2 FILLER_15_79 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_108 ();
 sg13g2_decap_8 FILLER_15_115 ();
 sg13g2_decap_8 FILLER_15_122 ();
 sg13g2_decap_4 FILLER_15_129 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_fill_2 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_197 ();
 sg13g2_fill_1 FILLER_15_199 ();
 sg13g2_decap_4 FILLER_15_216 ();
 sg13g2_fill_2 FILLER_15_220 ();
 sg13g2_decap_8 FILLER_15_226 ();
 sg13g2_decap_8 FILLER_15_233 ();
 sg13g2_decap_4 FILLER_15_240 ();
 sg13g2_fill_2 FILLER_15_254 ();
 sg13g2_fill_1 FILLER_15_256 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_268 ();
 sg13g2_decap_8 FILLER_15_275 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_301 ();
 sg13g2_fill_1 FILLER_15_307 ();
 sg13g2_decap_4 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_4 FILLER_15_362 ();
 sg13g2_fill_1 FILLER_15_366 ();
 sg13g2_decap_4 FILLER_15_372 ();
 sg13g2_fill_2 FILLER_15_386 ();
 sg13g2_decap_4 FILLER_15_444 ();
 sg13g2_fill_2 FILLER_15_453 ();
 sg13g2_fill_1 FILLER_15_477 ();
 sg13g2_fill_1 FILLER_15_483 ();
 sg13g2_fill_2 FILLER_15_488 ();
 sg13g2_fill_1 FILLER_15_490 ();
 sg13g2_fill_1 FILLER_15_495 ();
 sg13g2_decap_8 FILLER_15_505 ();
 sg13g2_fill_2 FILLER_15_512 ();
 sg13g2_fill_2 FILLER_15_527 ();
 sg13g2_fill_1 FILLER_15_529 ();
 sg13g2_fill_1 FILLER_15_556 ();
 sg13g2_fill_1 FILLER_15_588 ();
 sg13g2_fill_1 FILLER_15_593 ();
 sg13g2_fill_2 FILLER_15_629 ();
 sg13g2_fill_1 FILLER_15_631 ();
 sg13g2_fill_2 FILLER_15_643 ();
 sg13g2_decap_4 FILLER_15_650 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_fill_2 FILLER_15_665 ();
 sg13g2_decap_4 FILLER_15_705 ();
 sg13g2_fill_1 FILLER_15_709 ();
 sg13g2_fill_1 FILLER_15_721 ();
 sg13g2_decap_4 FILLER_15_757 ();
 sg13g2_fill_1 FILLER_15_761 ();
 sg13g2_decap_8 FILLER_15_771 ();
 sg13g2_decap_8 FILLER_15_778 ();
 sg13g2_decap_4 FILLER_15_785 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_4 FILLER_15_805 ();
 sg13g2_fill_2 FILLER_15_809 ();
 sg13g2_decap_4 FILLER_15_815 ();
 sg13g2_decap_8 FILLER_15_823 ();
 sg13g2_fill_1 FILLER_15_830 ();
 sg13g2_decap_8 FILLER_15_835 ();
 sg13g2_fill_1 FILLER_15_842 ();
 sg13g2_decap_8 FILLER_15_869 ();
 sg13g2_decap_8 FILLER_15_876 ();
 sg13g2_decap_8 FILLER_15_883 ();
 sg13g2_decap_4 FILLER_15_890 ();
 sg13g2_fill_2 FILLER_15_894 ();
 sg13g2_decap_8 FILLER_15_925 ();
 sg13g2_fill_1 FILLER_15_961 ();
 sg13g2_decap_8 FILLER_15_966 ();
 sg13g2_fill_1 FILLER_15_973 ();
 sg13g2_fill_2 FILLER_15_981 ();
 sg13g2_decap_8 FILLER_15_1039 ();
 sg13g2_decap_4 FILLER_15_1046 ();
 sg13g2_decap_8 FILLER_15_1112 ();
 sg13g2_fill_2 FILLER_15_1119 ();
 sg13g2_fill_2 FILLER_15_1130 ();
 sg13g2_fill_1 FILLER_15_1132 ();
 sg13g2_decap_4 FILLER_15_1258 ();
 sg13g2_fill_2 FILLER_15_1262 ();
 sg13g2_decap_8 FILLER_15_1268 ();
 sg13g2_decap_8 FILLER_15_1275 ();
 sg13g2_decap_4 FILLER_15_1282 ();
 sg13g2_fill_1 FILLER_15_1286 ();
 sg13g2_fill_2 FILLER_15_1323 ();
 sg13g2_fill_1 FILLER_15_1325 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_17 ();
 sg13g2_fill_1 FILLER_16_25 ();
 sg13g2_decap_4 FILLER_16_31 ();
 sg13g2_decap_8 FILLER_16_43 ();
 sg13g2_fill_1 FILLER_16_50 ();
 sg13g2_decap_4 FILLER_16_59 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_fill_2 FILLER_16_98 ();
 sg13g2_fill_1 FILLER_16_134 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_194 ();
 sg13g2_decap_8 FILLER_16_225 ();
 sg13g2_decap_8 FILLER_16_232 ();
 sg13g2_decap_8 FILLER_16_239 ();
 sg13g2_decap_4 FILLER_16_246 ();
 sg13g2_decap_4 FILLER_16_276 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_fill_1 FILLER_16_299 ();
 sg13g2_decap_8 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_fill_2 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_351 ();
 sg13g2_fill_2 FILLER_16_396 ();
 sg13g2_fill_1 FILLER_16_403 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_16_419 ();
 sg13g2_fill_1 FILLER_16_421 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_decap_4 FILLER_16_439 ();
 sg13g2_decap_4 FILLER_16_447 ();
 sg13g2_fill_1 FILLER_16_455 ();
 sg13g2_fill_1 FILLER_16_464 ();
 sg13g2_fill_1 FILLER_16_470 ();
 sg13g2_fill_1 FILLER_16_475 ();
 sg13g2_fill_1 FILLER_16_493 ();
 sg13g2_fill_2 FILLER_16_499 ();
 sg13g2_decap_8 FILLER_16_505 ();
 sg13g2_decap_4 FILLER_16_512 ();
 sg13g2_fill_1 FILLER_16_516 ();
 sg13g2_fill_1 FILLER_16_520 ();
 sg13g2_fill_2 FILLER_16_530 ();
 sg13g2_decap_8 FILLER_16_545 ();
 sg13g2_decap_8 FILLER_16_552 ();
 sg13g2_decap_8 FILLER_16_559 ();
 sg13g2_decap_4 FILLER_16_566 ();
 sg13g2_decap_8 FILLER_16_589 ();
 sg13g2_fill_1 FILLER_16_596 ();
 sg13g2_decap_4 FILLER_16_605 ();
 sg13g2_fill_2 FILLER_16_613 ();
 sg13g2_decap_4 FILLER_16_630 ();
 sg13g2_fill_1 FILLER_16_634 ();
 sg13g2_fill_1 FILLER_16_638 ();
 sg13g2_fill_2 FILLER_16_705 ();
 sg13g2_fill_1 FILLER_16_707 ();
 sg13g2_decap_4 FILLER_16_717 ();
 sg13g2_fill_1 FILLER_16_721 ();
 sg13g2_fill_2 FILLER_16_735 ();
 sg13g2_fill_1 FILLER_16_737 ();
 sg13g2_fill_2 FILLER_16_779 ();
 sg13g2_fill_1 FILLER_16_795 ();
 sg13g2_decap_8 FILLER_16_822 ();
 sg13g2_fill_2 FILLER_16_829 ();
 sg13g2_decap_4 FILLER_16_835 ();
 sg13g2_fill_2 FILLER_16_843 ();
 sg13g2_fill_1 FILLER_16_849 ();
 sg13g2_decap_4 FILLER_16_859 ();
 sg13g2_fill_2 FILLER_16_863 ();
 sg13g2_decap_4 FILLER_16_879 ();
 sg13g2_decap_8 FILLER_16_887 ();
 sg13g2_decap_8 FILLER_16_894 ();
 sg13g2_fill_2 FILLER_16_901 ();
 sg13g2_decap_8 FILLER_16_907 ();
 sg13g2_decap_8 FILLER_16_914 ();
 sg13g2_fill_1 FILLER_16_932 ();
 sg13g2_fill_1 FILLER_16_943 ();
 sg13g2_fill_2 FILLER_16_989 ();
 sg13g2_decap_8 FILLER_16_1002 ();
 sg13g2_decap_4 FILLER_16_1009 ();
 sg13g2_fill_1 FILLER_16_1018 ();
 sg13g2_fill_2 FILLER_16_1063 ();
 sg13g2_fill_1 FILLER_16_1065 ();
 sg13g2_decap_8 FILLER_16_1070 ();
 sg13g2_decap_8 FILLER_16_1077 ();
 sg13g2_decap_8 FILLER_16_1084 ();
 sg13g2_decap_8 FILLER_16_1124 ();
 sg13g2_decap_8 FILLER_16_1131 ();
 sg13g2_decap_8 FILLER_16_1138 ();
 sg13g2_decap_8 FILLER_16_1145 ();
 sg13g2_fill_2 FILLER_16_1152 ();
 sg13g2_fill_1 FILLER_16_1154 ();
 sg13g2_decap_4 FILLER_16_1176 ();
 sg13g2_decap_8 FILLER_16_1188 ();
 sg13g2_decap_8 FILLER_16_1195 ();
 sg13g2_fill_2 FILLER_16_1202 ();
 sg13g2_decap_8 FILLER_16_1208 ();
 sg13g2_decap_4 FILLER_16_1215 ();
 sg13g2_fill_2 FILLER_16_1219 ();
 sg13g2_fill_2 FILLER_16_1231 ();
 sg13g2_fill_1 FILLER_16_1233 ();
 sg13g2_fill_1 FILLER_16_1247 ();
 sg13g2_decap_4 FILLER_16_1284 ();
 sg13g2_fill_2 FILLER_16_1324 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_50 ();
 sg13g2_fill_2 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_58 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_2 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_72 ();
 sg13g2_fill_1 FILLER_17_76 ();
 sg13g2_fill_2 FILLER_17_110 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_134 ();
 sg13g2_fill_1 FILLER_17_166 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_fill_2 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_184 ();
 sg13g2_fill_1 FILLER_17_190 ();
 sg13g2_fill_2 FILLER_17_247 ();
 sg13g2_fill_1 FILLER_17_249 ();
 sg13g2_decap_4 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_fill_2 FILLER_17_298 ();
 sg13g2_fill_1 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_fill_2 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_fill_1 FILLER_17_341 ();
 sg13g2_fill_1 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_4 FILLER_17_371 ();
 sg13g2_fill_2 FILLER_17_409 ();
 sg13g2_fill_1 FILLER_17_411 ();
 sg13g2_fill_1 FILLER_17_428 ();
 sg13g2_fill_1 FILLER_17_434 ();
 sg13g2_fill_2 FILLER_17_448 ();
 sg13g2_fill_1 FILLER_17_460 ();
 sg13g2_decap_8 FILLER_17_465 ();
 sg13g2_fill_2 FILLER_17_472 ();
 sg13g2_fill_1 FILLER_17_474 ();
 sg13g2_fill_1 FILLER_17_488 ();
 sg13g2_fill_2 FILLER_17_520 ();
 sg13g2_fill_1 FILLER_17_522 ();
 sg13g2_fill_2 FILLER_17_532 ();
 sg13g2_fill_2 FILLER_17_543 ();
 sg13g2_fill_1 FILLER_17_545 ();
 sg13g2_fill_2 FILLER_17_550 ();
 sg13g2_fill_1 FILLER_17_552 ();
 sg13g2_fill_1 FILLER_17_579 ();
 sg13g2_fill_1 FILLER_17_585 ();
 sg13g2_fill_1 FILLER_17_612 ();
 sg13g2_fill_1 FILLER_17_639 ();
 sg13g2_decap_8 FILLER_17_666 ();
 sg13g2_decap_4 FILLER_17_673 ();
 sg13g2_decap_8 FILLER_17_681 ();
 sg13g2_decap_8 FILLER_17_688 ();
 sg13g2_decap_8 FILLER_17_699 ();
 sg13g2_decap_4 FILLER_17_706 ();
 sg13g2_fill_1 FILLER_17_710 ();
 sg13g2_decap_4 FILLER_17_742 ();
 sg13g2_fill_1 FILLER_17_746 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_fill_2 FILLER_17_763 ();
 sg13g2_fill_2 FILLER_17_811 ();
 sg13g2_fill_1 FILLER_17_813 ();
 sg13g2_fill_1 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_859 ();
 sg13g2_decap_4 FILLER_17_866 ();
 sg13g2_fill_2 FILLER_17_870 ();
 sg13g2_decap_8 FILLER_17_902 ();
 sg13g2_decap_8 FILLER_17_909 ();
 sg13g2_fill_2 FILLER_17_916 ();
 sg13g2_fill_1 FILLER_17_935 ();
 sg13g2_fill_2 FILLER_17_948 ();
 sg13g2_decap_8 FILLER_17_955 ();
 sg13g2_decap_4 FILLER_17_962 ();
 sg13g2_fill_2 FILLER_17_966 ();
 sg13g2_fill_2 FILLER_17_998 ();
 sg13g2_decap_8 FILLER_17_1032 ();
 sg13g2_fill_2 FILLER_17_1039 ();
 sg13g2_fill_1 FILLER_17_1041 ();
 sg13g2_decap_8 FILLER_17_1050 ();
 sg13g2_fill_2 FILLER_17_1057 ();
 sg13g2_fill_1 FILLER_17_1059 ();
 sg13g2_fill_1 FILLER_17_1090 ();
 sg13g2_fill_1 FILLER_17_1101 ();
 sg13g2_decap_8 FILLER_17_1106 ();
 sg13g2_fill_2 FILLER_17_1117 ();
 sg13g2_fill_2 FILLER_17_1164 ();
 sg13g2_fill_1 FILLER_17_1166 ();
 sg13g2_fill_1 FILLER_17_1171 ();
 sg13g2_fill_2 FILLER_17_1263 ();
 sg13g2_decap_8 FILLER_17_1295 ();
 sg13g2_fill_2 FILLER_17_1302 ();
 sg13g2_fill_1 FILLER_17_1304 ();
 sg13g2_decap_8 FILLER_17_1309 ();
 sg13g2_decap_8 FILLER_17_1316 ();
 sg13g2_fill_2 FILLER_17_1323 ();
 sg13g2_fill_1 FILLER_17_1325 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_fill_2 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_37 ();
 sg13g2_decap_4 FILLER_18_52 ();
 sg13g2_fill_1 FILLER_18_66 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_4 FILLER_18_108 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_fill_1 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_131 ();
 sg13g2_fill_2 FILLER_18_164 ();
 sg13g2_fill_1 FILLER_18_166 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_fill_2 FILLER_18_189 ();
 sg13g2_fill_1 FILLER_18_201 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_227 ();
 sg13g2_fill_2 FILLER_18_234 ();
 sg13g2_decap_8 FILLER_18_241 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_fill_1 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_260 ();
 sg13g2_decap_4 FILLER_18_267 ();
 sg13g2_decap_4 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_279 ();
 sg13g2_fill_2 FILLER_18_292 ();
 sg13g2_decap_4 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_344 ();
 sg13g2_decap_4 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_374 ();
 sg13g2_fill_1 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_fill_2 FILLER_18_400 ();
 sg13g2_fill_1 FILLER_18_402 ();
 sg13g2_fill_2 FILLER_18_436 ();
 sg13g2_fill_2 FILLER_18_484 ();
 sg13g2_fill_2 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_501 ();
 sg13g2_decap_8 FILLER_18_508 ();
 sg13g2_decap_4 FILLER_18_515 ();
 sg13g2_fill_2 FILLER_18_519 ();
 sg13g2_fill_1 FILLER_18_563 ();
 sg13g2_fill_2 FILLER_18_568 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_fill_2 FILLER_18_581 ();
 sg13g2_fill_1 FILLER_18_583 ();
 sg13g2_decap_8 FILLER_18_610 ();
 sg13g2_fill_1 FILLER_18_617 ();
 sg13g2_fill_2 FILLER_18_627 ();
 sg13g2_fill_1 FILLER_18_629 ();
 sg13g2_fill_2 FILLER_18_635 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_fill_2 FILLER_18_693 ();
 sg13g2_fill_1 FILLER_18_695 ();
 sg13g2_decap_4 FILLER_18_722 ();
 sg13g2_fill_1 FILLER_18_726 ();
 sg13g2_decap_4 FILLER_18_771 ();
 sg13g2_fill_1 FILLER_18_775 ();
 sg13g2_fill_2 FILLER_18_796 ();
 sg13g2_decap_8 FILLER_18_802 ();
 sg13g2_fill_2 FILLER_18_809 ();
 sg13g2_fill_1 FILLER_18_811 ();
 sg13g2_fill_2 FILLER_18_822 ();
 sg13g2_fill_1 FILLER_18_824 ();
 sg13g2_fill_2 FILLER_18_829 ();
 sg13g2_fill_1 FILLER_18_831 ();
 sg13g2_fill_1 FILLER_18_842 ();
 sg13g2_fill_1 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_852 ();
 sg13g2_fill_1 FILLER_18_859 ();
 sg13g2_decap_8 FILLER_18_865 ();
 sg13g2_fill_2 FILLER_18_872 ();
 sg13g2_decap_4 FILLER_18_891 ();
 sg13g2_fill_1 FILLER_18_899 ();
 sg13g2_fill_1 FILLER_18_926 ();
 sg13g2_fill_1 FILLER_18_944 ();
 sg13g2_fill_2 FILLER_18_949 ();
 sg13g2_decap_8 FILLER_18_956 ();
 sg13g2_fill_2 FILLER_18_963 ();
 sg13g2_fill_1 FILLER_18_965 ();
 sg13g2_fill_1 FILLER_18_975 ();
 sg13g2_decap_8 FILLER_18_980 ();
 sg13g2_fill_1 FILLER_18_987 ();
 sg13g2_decap_4 FILLER_18_993 ();
 sg13g2_fill_2 FILLER_18_1007 ();
 sg13g2_decap_8 FILLER_18_1013 ();
 sg13g2_decap_4 FILLER_18_1020 ();
 sg13g2_fill_2 FILLER_18_1024 ();
 sg13g2_decap_8 FILLER_18_1061 ();
 sg13g2_decap_8 FILLER_18_1068 ();
 sg13g2_decap_8 FILLER_18_1079 ();
 sg13g2_decap_4 FILLER_18_1086 ();
 sg13g2_decap_8 FILLER_18_1094 ();
 sg13g2_decap_8 FILLER_18_1101 ();
 sg13g2_decap_8 FILLER_18_1108 ();
 sg13g2_fill_2 FILLER_18_1115 ();
 sg13g2_fill_1 FILLER_18_1117 ();
 sg13g2_fill_1 FILLER_18_1132 ();
 sg13g2_decap_4 FILLER_18_1169 ();
 sg13g2_fill_2 FILLER_18_1178 ();
 sg13g2_fill_2 FILLER_18_1185 ();
 sg13g2_fill_1 FILLER_18_1187 ();
 sg13g2_fill_2 FILLER_18_1214 ();
 sg13g2_fill_1 FILLER_18_1216 ();
 sg13g2_fill_1 FILLER_18_1232 ();
 sg13g2_fill_2 FILLER_18_1237 ();
 sg13g2_fill_1 FILLER_18_1239 ();
 sg13g2_fill_2 FILLER_18_1244 ();
 sg13g2_decap_4 FILLER_18_1251 ();
 sg13g2_decap_8 FILLER_18_1268 ();
 sg13g2_decap_4 FILLER_18_1275 ();
 sg13g2_fill_2 FILLER_18_1323 ();
 sg13g2_fill_1 FILLER_18_1325 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_2 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_57 ();
 sg13g2_fill_1 FILLER_19_62 ();
 sg13g2_fill_2 FILLER_19_77 ();
 sg13g2_fill_1 FILLER_19_79 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_fill_1 FILLER_19_91 ();
 sg13g2_decap_4 FILLER_19_96 ();
 sg13g2_fill_1 FILLER_19_100 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_decap_4 FILLER_19_117 ();
 sg13g2_fill_2 FILLER_19_121 ();
 sg13g2_decap_8 FILLER_19_128 ();
 sg13g2_decap_8 FILLER_19_135 ();
 sg13g2_decap_8 FILLER_19_142 ();
 sg13g2_fill_2 FILLER_19_149 ();
 sg13g2_fill_1 FILLER_19_151 ();
 sg13g2_fill_1 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_165 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_fill_2 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_fill_2 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_fill_2 FILLER_19_298 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_309 ();
 sg13g2_fill_2 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_317 ();
 sg13g2_fill_1 FILLER_19_338 ();
 sg13g2_fill_1 FILLER_19_353 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_4 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_fill_2 FILLER_19_398 ();
 sg13g2_decap_8 FILLER_19_431 ();
 sg13g2_fill_2 FILLER_19_441 ();
 sg13g2_fill_1 FILLER_19_452 ();
 sg13g2_fill_1 FILLER_19_458 ();
 sg13g2_decap_4 FILLER_19_485 ();
 sg13g2_fill_2 FILLER_19_489 ();
 sg13g2_decap_4 FILLER_19_527 ();
 sg13g2_fill_1 FILLER_19_531 ();
 sg13g2_decap_8 FILLER_19_537 ();
 sg13g2_fill_1 FILLER_19_544 ();
 sg13g2_fill_1 FILLER_19_549 ();
 sg13g2_fill_1 FILLER_19_576 ();
 sg13g2_fill_1 FILLER_19_587 ();
 sg13g2_fill_2 FILLER_19_600 ();
 sg13g2_fill_1 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_613 ();
 sg13g2_decap_8 FILLER_19_620 ();
 sg13g2_decap_4 FILLER_19_627 ();
 sg13g2_fill_1 FILLER_19_636 ();
 sg13g2_fill_2 FILLER_19_642 ();
 sg13g2_fill_1 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_671 ();
 sg13g2_fill_1 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_718 ();
 sg13g2_decap_8 FILLER_19_725 ();
 sg13g2_fill_2 FILLER_19_732 ();
 sg13g2_decap_4 FILLER_19_743 ();
 sg13g2_fill_2 FILLER_19_759 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_4 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_2 FILLER_19_938 ();
 sg13g2_fill_1 FILLER_19_940 ();
 sg13g2_fill_1 FILLER_19_946 ();
 sg13g2_fill_2 FILLER_19_973 ();
 sg13g2_fill_1 FILLER_19_980 ();
 sg13g2_fill_2 FILLER_19_985 ();
 sg13g2_decap_8 FILLER_19_991 ();
 sg13g2_fill_1 FILLER_19_1003 ();
 sg13g2_fill_2 FILLER_19_1030 ();
 sg13g2_fill_1 FILLER_19_1032 ();
 sg13g2_fill_1 FILLER_19_1126 ();
 sg13g2_decap_4 FILLER_19_1149 ();
 sg13g2_decap_8 FILLER_19_1157 ();
 sg13g2_fill_2 FILLER_19_1164 ();
 sg13g2_decap_4 FILLER_19_1192 ();
 sg13g2_fill_1 FILLER_19_1196 ();
 sg13g2_fill_1 FILLER_19_1209 ();
 sg13g2_decap_8 FILLER_19_1214 ();
 sg13g2_fill_1 FILLER_19_1221 ();
 sg13g2_fill_1 FILLER_19_1240 ();
 sg13g2_fill_1 FILLER_19_1267 ();
 sg13g2_fill_1 FILLER_19_1272 ();
 sg13g2_fill_1 FILLER_19_1283 ();
 sg13g2_fill_2 FILLER_19_1294 ();
 sg13g2_fill_1 FILLER_19_1296 ();
 sg13g2_fill_2 FILLER_19_1301 ();
 sg13g2_decap_8 FILLER_19_1307 ();
 sg13g2_decap_8 FILLER_19_1314 ();
 sg13g2_decap_4 FILLER_19_1321 ();
 sg13g2_fill_1 FILLER_19_1325 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_18 ();
 sg13g2_fill_2 FILLER_20_38 ();
 sg13g2_fill_1 FILLER_20_48 ();
 sg13g2_decap_4 FILLER_20_54 ();
 sg13g2_fill_2 FILLER_20_58 ();
 sg13g2_fill_2 FILLER_20_69 ();
 sg13g2_fill_2 FILLER_20_86 ();
 sg13g2_decap_8 FILLER_20_92 ();
 sg13g2_decap_4 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_103 ();
 sg13g2_decap_4 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_fill_2 FILLER_20_140 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_decap_4 FILLER_20_154 ();
 sg13g2_fill_1 FILLER_20_176 ();
 sg13g2_decap_4 FILLER_20_185 ();
 sg13g2_decap_4 FILLER_20_225 ();
 sg13g2_fill_2 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_decap_4 FILLER_20_286 ();
 sg13g2_decap_4 FILLER_20_302 ();
 sg13g2_decap_8 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_328 ();
 sg13g2_fill_1 FILLER_20_330 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_344 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_356 ();
 sg13g2_fill_1 FILLER_20_360 ();
 sg13g2_fill_1 FILLER_20_366 ();
 sg13g2_decap_4 FILLER_20_440 ();
 sg13g2_fill_2 FILLER_20_462 ();
 sg13g2_fill_1 FILLER_20_464 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_4 FILLER_20_476 ();
 sg13g2_fill_2 FILLER_20_480 ();
 sg13g2_decap_8 FILLER_20_488 ();
 sg13g2_decap_4 FILLER_20_495 ();
 sg13g2_fill_1 FILLER_20_499 ();
 sg13g2_fill_2 FILLER_20_510 ();
 sg13g2_fill_1 FILLER_20_551 ();
 sg13g2_fill_2 FILLER_20_560 ();
 sg13g2_fill_1 FILLER_20_572 ();
 sg13g2_fill_1 FILLER_20_578 ();
 sg13g2_fill_1 FILLER_20_584 ();
 sg13g2_decap_8 FILLER_20_611 ();
 sg13g2_fill_2 FILLER_20_618 ();
 sg13g2_decap_4 FILLER_20_630 ();
 sg13g2_fill_2 FILLER_20_664 ();
 sg13g2_decap_8 FILLER_20_692 ();
 sg13g2_decap_8 FILLER_20_699 ();
 sg13g2_fill_1 FILLER_20_706 ();
 sg13g2_decap_8 FILLER_20_716 ();
 sg13g2_fill_2 FILLER_20_723 ();
 sg13g2_fill_1 FILLER_20_725 ();
 sg13g2_fill_1 FILLER_20_730 ();
 sg13g2_fill_1 FILLER_20_745 ();
 sg13g2_fill_1 FILLER_20_750 ();
 sg13g2_fill_2 FILLER_20_764 ();
 sg13g2_fill_2 FILLER_20_803 ();
 sg13g2_fill_1 FILLER_20_805 ();
 sg13g2_fill_1 FILLER_20_811 ();
 sg13g2_decap_8 FILLER_20_820 ();
 sg13g2_decap_4 FILLER_20_827 ();
 sg13g2_fill_1 FILLER_20_835 ();
 sg13g2_decap_8 FILLER_20_867 ();
 sg13g2_fill_1 FILLER_20_883 ();
 sg13g2_decap_8 FILLER_20_888 ();
 sg13g2_decap_8 FILLER_20_895 ();
 sg13g2_decap_4 FILLER_20_902 ();
 sg13g2_fill_1 FILLER_20_906 ();
 sg13g2_decap_4 FILLER_20_919 ();
 sg13g2_fill_1 FILLER_20_923 ();
 sg13g2_fill_2 FILLER_20_937 ();
 sg13g2_fill_1 FILLER_20_948 ();
 sg13g2_fill_2 FILLER_20_960 ();
 sg13g2_fill_1 FILLER_20_962 ();
 sg13g2_fill_2 FILLER_20_1013 ();
 sg13g2_decap_4 FILLER_20_1019 ();
 sg13g2_fill_1 FILLER_20_1023 ();
 sg13g2_fill_2 FILLER_20_1032 ();
 sg13g2_decap_8 FILLER_20_1038 ();
 sg13g2_fill_2 FILLER_20_1045 ();
 sg13g2_decap_4 FILLER_20_1051 ();
 sg13g2_fill_1 FILLER_20_1055 ();
 sg13g2_fill_1 FILLER_20_1088 ();
 sg13g2_fill_2 FILLER_20_1132 ();
 sg13g2_decap_4 FILLER_20_1176 ();
 sg13g2_decap_8 FILLER_20_1184 ();
 sg13g2_decap_8 FILLER_20_1191 ();
 sg13g2_decap_4 FILLER_20_1198 ();
 sg13g2_fill_1 FILLER_20_1202 ();
 sg13g2_fill_1 FILLER_20_1229 ();
 sg13g2_fill_2 FILLER_20_1237 ();
 sg13g2_fill_1 FILLER_20_1244 ();
 sg13g2_decap_8 FILLER_20_1253 ();
 sg13g2_decap_4 FILLER_20_1260 ();
 sg13g2_fill_1 FILLER_20_1264 ();
 sg13g2_decap_8 FILLER_20_1317 ();
 sg13g2_fill_2 FILLER_20_1324 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_36 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_decap_4 FILLER_21_72 ();
 sg13g2_decap_4 FILLER_21_94 ();
 sg13g2_fill_2 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_111 ();
 sg13g2_fill_2 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_174 ();
 sg13g2_decap_4 FILLER_21_181 ();
 sg13g2_fill_2 FILLER_21_185 ();
 sg13g2_decap_4 FILLER_21_196 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_241 ();
 sg13g2_decap_8 FILLER_21_250 ();
 sg13g2_decap_4 FILLER_21_257 ();
 sg13g2_fill_1 FILLER_21_270 ();
 sg13g2_decap_4 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_fill_1 FILLER_21_284 ();
 sg13g2_fill_2 FILLER_21_293 ();
 sg13g2_fill_1 FILLER_21_295 ();
 sg13g2_fill_2 FILLER_21_311 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_fill_2 FILLER_21_328 ();
 sg13g2_fill_1 FILLER_21_330 ();
 sg13g2_decap_4 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_4 FILLER_21_383 ();
 sg13g2_fill_1 FILLER_21_387 ();
 sg13g2_decap_4 FILLER_21_393 ();
 sg13g2_fill_2 FILLER_21_397 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_450 ();
 sg13g2_decap_8 FILLER_21_457 ();
 sg13g2_decap_8 FILLER_21_464 ();
 sg13g2_fill_1 FILLER_21_471 ();
 sg13g2_decap_4 FILLER_21_519 ();
 sg13g2_fill_1 FILLER_21_523 ();
 sg13g2_decap_8 FILLER_21_528 ();
 sg13g2_fill_2 FILLER_21_535 ();
 sg13g2_fill_2 FILLER_21_541 ();
 sg13g2_fill_2 FILLER_21_549 ();
 sg13g2_decap_8 FILLER_21_605 ();
 sg13g2_decap_4 FILLER_21_624 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_fill_1 FILLER_21_689 ();
 sg13g2_decap_4 FILLER_21_726 ();
 sg13g2_decap_8 FILLER_21_744 ();
 sg13g2_decap_8 FILLER_21_751 ();
 sg13g2_fill_2 FILLER_21_766 ();
 sg13g2_fill_2 FILLER_21_798 ();
 sg13g2_decap_4 FILLER_21_834 ();
 sg13g2_fill_2 FILLER_21_838 ();
 sg13g2_decap_4 FILLER_21_852 ();
 sg13g2_fill_2 FILLER_21_860 ();
 sg13g2_fill_1 FILLER_21_862 ();
 sg13g2_fill_2 FILLER_21_871 ();
 sg13g2_fill_1 FILLER_21_873 ();
 sg13g2_fill_1 FILLER_21_935 ();
 sg13g2_fill_2 FILLER_21_944 ();
 sg13g2_decap_8 FILLER_21_956 ();
 sg13g2_decap_8 FILLER_21_963 ();
 sg13g2_decap_4 FILLER_21_970 ();
 sg13g2_fill_2 FILLER_21_978 ();
 sg13g2_fill_2 FILLER_21_985 ();
 sg13g2_fill_1 FILLER_21_987 ();
 sg13g2_fill_2 FILLER_21_993 ();
 sg13g2_fill_1 FILLER_21_995 ();
 sg13g2_fill_2 FILLER_21_1002 ();
 sg13g2_fill_1 FILLER_21_1004 ();
 sg13g2_fill_1 FILLER_21_1026 ();
 sg13g2_decap_8 FILLER_21_1053 ();
 sg13g2_decap_4 FILLER_21_1060 ();
 sg13g2_fill_1 FILLER_21_1064 ();
 sg13g2_decap_4 FILLER_21_1077 ();
 sg13g2_fill_1 FILLER_21_1081 ();
 sg13g2_decap_4 FILLER_21_1092 ();
 sg13g2_fill_2 FILLER_21_1096 ();
 sg13g2_fill_2 FILLER_21_1102 ();
 sg13g2_fill_2 FILLER_21_1108 ();
 sg13g2_fill_2 FILLER_21_1114 ();
 sg13g2_fill_1 FILLER_21_1116 ();
 sg13g2_fill_2 FILLER_21_1127 ();
 sg13g2_fill_1 FILLER_21_1129 ();
 sg13g2_decap_4 FILLER_21_1134 ();
 sg13g2_fill_2 FILLER_21_1142 ();
 sg13g2_fill_1 FILLER_21_1144 ();
 sg13g2_decap_8 FILLER_21_1154 ();
 sg13g2_fill_2 FILLER_21_1161 ();
 sg13g2_decap_4 FILLER_21_1230 ();
 sg13g2_fill_1 FILLER_21_1234 ();
 sg13g2_decap_4 FILLER_21_1265 ();
 sg13g2_fill_1 FILLER_21_1269 ();
 sg13g2_decap_8 FILLER_21_1280 ();
 sg13g2_fill_2 FILLER_21_1287 ();
 sg13g2_fill_1 FILLER_21_1289 ();
 sg13g2_decap_8 FILLER_21_1300 ();
 sg13g2_decap_8 FILLER_21_1307 ();
 sg13g2_decap_8 FILLER_21_1314 ();
 sg13g2_decap_4 FILLER_21_1321 ();
 sg13g2_fill_1 FILLER_21_1325 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_fill_2 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_2 FILLER_22_51 ();
 sg13g2_fill_1 FILLER_22_75 ();
 sg13g2_fill_2 FILLER_22_81 ();
 sg13g2_fill_2 FILLER_22_88 ();
 sg13g2_fill_2 FILLER_22_94 ();
 sg13g2_fill_1 FILLER_22_104 ();
 sg13g2_fill_1 FILLER_22_116 ();
 sg13g2_fill_1 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_2 FILLER_22_156 ();
 sg13g2_fill_2 FILLER_22_176 ();
 sg13g2_decap_4 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_fill_2 FILLER_22_213 ();
 sg13g2_fill_1 FILLER_22_215 ();
 sg13g2_fill_2 FILLER_22_221 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_229 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_fill_2 FILLER_22_240 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_decap_8 FILLER_22_293 ();
 sg13g2_decap_4 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_304 ();
 sg13g2_decap_4 FILLER_22_311 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_fill_2 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_337 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_4 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_decap_8 FILLER_22_418 ();
 sg13g2_decap_8 FILLER_22_425 ();
 sg13g2_decap_4 FILLER_22_432 ();
 sg13g2_decap_4 FILLER_22_441 ();
 sg13g2_decap_4 FILLER_22_475 ();
 sg13g2_fill_1 FILLER_22_490 ();
 sg13g2_fill_2 FILLER_22_495 ();
 sg13g2_decap_8 FILLER_22_502 ();
 sg13g2_decap_4 FILLER_22_509 ();
 sg13g2_fill_2 FILLER_22_554 ();
 sg13g2_decap_4 FILLER_22_582 ();
 sg13g2_fill_2 FILLER_22_586 ();
 sg13g2_decap_4 FILLER_22_606 ();
 sg13g2_decap_8 FILLER_22_621 ();
 sg13g2_decap_4 FILLER_22_628 ();
 sg13g2_fill_1 FILLER_22_632 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_fill_2 FILLER_22_644 ();
 sg13g2_fill_1 FILLER_22_646 ();
 sg13g2_decap_4 FILLER_22_684 ();
 sg13g2_fill_1 FILLER_22_693 ();
 sg13g2_fill_1 FILLER_22_702 ();
 sg13g2_decap_8 FILLER_22_729 ();
 sg13g2_fill_2 FILLER_22_736 ();
 sg13g2_decap_8 FILLER_22_743 ();
 sg13g2_decap_8 FILLER_22_750 ();
 sg13g2_decap_4 FILLER_22_757 ();
 sg13g2_fill_2 FILLER_22_761 ();
 sg13g2_fill_2 FILLER_22_779 ();
 sg13g2_fill_1 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_800 ();
 sg13g2_fill_2 FILLER_22_807 ();
 sg13g2_decap_4 FILLER_22_818 ();
 sg13g2_decap_4 FILLER_22_834 ();
 sg13g2_fill_2 FILLER_22_838 ();
 sg13g2_fill_1 FILLER_22_848 ();
 sg13g2_fill_2 FILLER_22_875 ();
 sg13g2_fill_2 FILLER_22_913 ();
 sg13g2_fill_2 FILLER_22_919 ();
 sg13g2_fill_1 FILLER_22_921 ();
 sg13g2_fill_1 FILLER_22_932 ();
 sg13g2_fill_1 FILLER_22_938 ();
 sg13g2_fill_1 FILLER_22_1003 ();
 sg13g2_fill_1 FILLER_22_1030 ();
 sg13g2_fill_1 FILLER_22_1041 ();
 sg13g2_fill_1 FILLER_22_1068 ();
 sg13g2_fill_1 FILLER_22_1173 ();
 sg13g2_decap_8 FILLER_22_1200 ();
 sg13g2_fill_2 FILLER_22_1207 ();
 sg13g2_fill_2 FILLER_22_1213 ();
 sg13g2_decap_4 FILLER_22_1220 ();
 sg13g2_fill_1 FILLER_22_1224 ();
 sg13g2_fill_1 FILLER_22_1229 ();
 sg13g2_decap_4 FILLER_22_1240 ();
 sg13g2_decap_4 FILLER_22_1270 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_34 ();
 sg13g2_decap_4 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_44 ();
 sg13g2_decap_8 FILLER_23_50 ();
 sg13g2_fill_2 FILLER_23_57 ();
 sg13g2_decap_4 FILLER_23_71 ();
 sg13g2_fill_1 FILLER_23_75 ();
 sg13g2_decap_4 FILLER_23_79 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_96 ();
 sg13g2_fill_2 FILLER_23_103 ();
 sg13g2_decap_4 FILLER_23_117 ();
 sg13g2_fill_1 FILLER_23_130 ();
 sg13g2_fill_1 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_146 ();
 sg13g2_fill_1 FILLER_23_150 ();
 sg13g2_decap_8 FILLER_23_155 ();
 sg13g2_decap_8 FILLER_23_162 ();
 sg13g2_decap_8 FILLER_23_169 ();
 sg13g2_decap_8 FILLER_23_176 ();
 sg13g2_decap_8 FILLER_23_183 ();
 sg13g2_decap_4 FILLER_23_190 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_decap_8 FILLER_23_209 ();
 sg13g2_decap_4 FILLER_23_216 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_251 ();
 sg13g2_decap_8 FILLER_23_257 ();
 sg13g2_fill_2 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_270 ();
 sg13g2_fill_1 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_fill_2 FILLER_23_390 ();
 sg13g2_fill_1 FILLER_23_392 ();
 sg13g2_fill_1 FILLER_23_401 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_fill_2 FILLER_23_413 ();
 sg13g2_fill_1 FILLER_23_441 ();
 sg13g2_fill_2 FILLER_23_463 ();
 sg13g2_fill_1 FILLER_23_474 ();
 sg13g2_decap_4 FILLER_23_479 ();
 sg13g2_decap_4 FILLER_23_487 ();
 sg13g2_fill_2 FILLER_23_491 ();
 sg13g2_decap_4 FILLER_23_528 ();
 sg13g2_decap_8 FILLER_23_541 ();
 sg13g2_decap_8 FILLER_23_548 ();
 sg13g2_decap_4 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_568 ();
 sg13g2_fill_1 FILLER_23_575 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_4 FILLER_23_644 ();
 sg13g2_fill_2 FILLER_23_648 ();
 sg13g2_decap_8 FILLER_23_654 ();
 sg13g2_decap_4 FILLER_23_661 ();
 sg13g2_decap_4 FILLER_23_675 ();
 sg13g2_fill_2 FILLER_23_720 ();
 sg13g2_fill_1 FILLER_23_722 ();
 sg13g2_fill_1 FILLER_23_759 ();
 sg13g2_fill_1 FILLER_23_786 ();
 sg13g2_fill_1 FILLER_23_813 ();
 sg13g2_fill_1 FILLER_23_819 ();
 sg13g2_fill_1 FILLER_23_829 ();
 sg13g2_decap_8 FILLER_23_834 ();
 sg13g2_fill_2 FILLER_23_841 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_fill_2 FILLER_23_854 ();
 sg13g2_decap_8 FILLER_23_901 ();
 sg13g2_decap_8 FILLER_23_912 ();
 sg13g2_decap_4 FILLER_23_919 ();
 sg13g2_fill_1 FILLER_23_923 ();
 sg13g2_decap_4 FILLER_23_940 ();
 sg13g2_fill_2 FILLER_23_944 ();
 sg13g2_decap_4 FILLER_23_958 ();
 sg13g2_fill_2 FILLER_23_962 ();
 sg13g2_fill_1 FILLER_23_968 ();
 sg13g2_fill_1 FILLER_23_974 ();
 sg13g2_fill_1 FILLER_23_984 ();
 sg13g2_fill_1 FILLER_23_989 ();
 sg13g2_fill_2 FILLER_23_995 ();
 sg13g2_decap_8 FILLER_23_1001 ();
 sg13g2_decap_4 FILLER_23_1008 ();
 sg13g2_fill_1 FILLER_23_1012 ();
 sg13g2_decap_8 FILLER_23_1027 ();
 sg13g2_fill_1 FILLER_23_1034 ();
 sg13g2_decap_4 FILLER_23_1045 ();
 sg13g2_decap_8 FILLER_23_1057 ();
 sg13g2_decap_8 FILLER_23_1064 ();
 sg13g2_fill_2 FILLER_23_1071 ();
 sg13g2_fill_1 FILLER_23_1073 ();
 sg13g2_decap_8 FILLER_23_1078 ();
 sg13g2_fill_2 FILLER_23_1085 ();
 sg13g2_fill_2 FILLER_23_1109 ();
 sg13g2_fill_1 FILLER_23_1111 ();
 sg13g2_decap_8 FILLER_23_1138 ();
 sg13g2_decap_4 FILLER_23_1145 ();
 sg13g2_fill_1 FILLER_23_1149 ();
 sg13g2_decap_8 FILLER_23_1159 ();
 sg13g2_fill_1 FILLER_23_1166 ();
 sg13g2_decap_4 FILLER_23_1177 ();
 sg13g2_fill_2 FILLER_23_1181 ();
 sg13g2_fill_2 FILLER_23_1187 ();
 sg13g2_decap_4 FILLER_23_1193 ();
 sg13g2_fill_1 FILLER_23_1219 ();
 sg13g2_fill_2 FILLER_23_1246 ();
 sg13g2_fill_1 FILLER_23_1248 ();
 sg13g2_decap_8 FILLER_23_1263 ();
 sg13g2_decap_8 FILLER_23_1270 ();
 sg13g2_decap_4 FILLER_23_1277 ();
 sg13g2_decap_8 FILLER_23_1285 ();
 sg13g2_decap_8 FILLER_23_1292 ();
 sg13g2_decap_8 FILLER_23_1299 ();
 sg13g2_fill_2 FILLER_23_1310 ();
 sg13g2_decap_8 FILLER_23_1316 ();
 sg13g2_fill_2 FILLER_23_1323 ();
 sg13g2_fill_1 FILLER_23_1325 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_27 ();
 sg13g2_fill_1 FILLER_24_32 ();
 sg13g2_fill_2 FILLER_24_38 ();
 sg13g2_fill_1 FILLER_24_45 ();
 sg13g2_decap_8 FILLER_24_50 ();
 sg13g2_fill_1 FILLER_24_62 ();
 sg13g2_decap_8 FILLER_24_72 ();
 sg13g2_fill_1 FILLER_24_79 ();
 sg13g2_fill_1 FILLER_24_89 ();
 sg13g2_fill_2 FILLER_24_95 ();
 sg13g2_fill_2 FILLER_24_102 ();
 sg13g2_fill_2 FILLER_24_109 ();
 sg13g2_fill_1 FILLER_24_111 ();
 sg13g2_decap_4 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_151 ();
 sg13g2_decap_4 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_fill_2 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_181 ();
 sg13g2_fill_1 FILLER_24_227 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_fill_2 FILLER_24_252 ();
 sg13g2_decap_4 FILLER_24_293 ();
 sg13g2_decap_4 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_318 ();
 sg13g2_fill_2 FILLER_24_323 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_fill_2 FILLER_24_340 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_decap_4 FILLER_24_351 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_425 ();
 sg13g2_fill_2 FILLER_24_463 ();
 sg13g2_fill_1 FILLER_24_495 ();
 sg13g2_fill_1 FILLER_24_500 ();
 sg13g2_fill_1 FILLER_24_505 ();
 sg13g2_fill_2 FILLER_24_510 ();
 sg13g2_fill_1 FILLER_24_598 ();
 sg13g2_decap_8 FILLER_24_603 ();
 sg13g2_fill_2 FILLER_24_610 ();
 sg13g2_fill_1 FILLER_24_643 ();
 sg13g2_fill_1 FILLER_24_670 ();
 sg13g2_fill_1 FILLER_24_675 ();
 sg13g2_decap_4 FILLER_24_702 ();
 sg13g2_fill_2 FILLER_24_706 ();
 sg13g2_fill_1 FILLER_24_738 ();
 sg13g2_decap_8 FILLER_24_743 ();
 sg13g2_decap_8 FILLER_24_750 ();
 sg13g2_fill_2 FILLER_24_757 ();
 sg13g2_fill_1 FILLER_24_768 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_4 FILLER_24_784 ();
 sg13g2_fill_1 FILLER_24_788 ();
 sg13g2_fill_2 FILLER_24_797 ();
 sg13g2_fill_2 FILLER_24_830 ();
 sg13g2_fill_2 FILLER_24_836 ();
 sg13g2_fill_2 FILLER_24_848 ();
 sg13g2_fill_1 FILLER_24_863 ();
 sg13g2_decap_8 FILLER_24_884 ();
 sg13g2_decap_4 FILLER_24_891 ();
 sg13g2_fill_2 FILLER_24_895 ();
 sg13g2_fill_2 FILLER_24_927 ();
 sg13g2_fill_2 FILLER_24_952 ();
 sg13g2_fill_1 FILLER_24_954 ();
 sg13g2_decap_4 FILLER_24_972 ();
 sg13g2_fill_2 FILLER_24_976 ();
 sg13g2_decap_4 FILLER_24_1013 ();
 sg13g2_fill_2 FILLER_24_1069 ();
 sg13g2_decap_4 FILLER_24_1075 ();
 sg13g2_fill_2 FILLER_24_1079 ();
 sg13g2_fill_2 FILLER_24_1085 ();
 sg13g2_fill_2 FILLER_24_1097 ();
 sg13g2_fill_1 FILLER_24_1099 ();
 sg13g2_fill_2 FILLER_24_1104 ();
 sg13g2_fill_1 FILLER_24_1106 ();
 sg13g2_fill_2 FILLER_24_1111 ();
 sg13g2_fill_1 FILLER_24_1113 ();
 sg13g2_fill_2 FILLER_24_1118 ();
 sg13g2_decap_8 FILLER_24_1124 ();
 sg13g2_decap_8 FILLER_24_1139 ();
 sg13g2_fill_1 FILLER_24_1146 ();
 sg13g2_decap_8 FILLER_24_1152 ();
 sg13g2_decap_4 FILLER_24_1159 ();
 sg13g2_fill_1 FILLER_24_1163 ();
 sg13g2_decap_4 FILLER_24_1229 ();
 sg13g2_fill_2 FILLER_24_1233 ();
 sg13g2_decap_8 FILLER_24_1261 ();
 sg13g2_decap_8 FILLER_24_1268 ();
 sg13g2_fill_2 FILLER_24_1279 ();
 sg13g2_fill_1 FILLER_24_1325 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_15 ();
 sg13g2_decap_8 FILLER_25_22 ();
 sg13g2_fill_2 FILLER_25_29 ();
 sg13g2_fill_1 FILLER_25_34 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_fill_1 FILLER_25_50 ();
 sg13g2_decap_8 FILLER_25_59 ();
 sg13g2_fill_1 FILLER_25_66 ();
 sg13g2_fill_2 FILLER_25_77 ();
 sg13g2_fill_1 FILLER_25_89 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_fill_2 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_decap_4 FILLER_25_230 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_285 ();
 sg13g2_decap_4 FILLER_25_293 ();
 sg13g2_decap_4 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_371 ();
 sg13g2_fill_1 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_411 ();
 sg13g2_decap_8 FILLER_25_418 ();
 sg13g2_fill_2 FILLER_25_425 ();
 sg13g2_decap_8 FILLER_25_440 ();
 sg13g2_fill_2 FILLER_25_451 ();
 sg13g2_fill_1 FILLER_25_457 ();
 sg13g2_fill_2 FILLER_25_462 ();
 sg13g2_fill_2 FILLER_25_468 ();
 sg13g2_fill_2 FILLER_25_474 ();
 sg13g2_fill_1 FILLER_25_486 ();
 sg13g2_fill_2 FILLER_25_492 ();
 sg13g2_fill_2 FILLER_25_498 ();
 sg13g2_fill_1 FILLER_25_500 ();
 sg13g2_fill_1 FILLER_25_506 ();
 sg13g2_decap_4 FILLER_25_528 ();
 sg13g2_fill_1 FILLER_25_532 ();
 sg13g2_fill_2 FILLER_25_546 ();
 sg13g2_fill_1 FILLER_25_548 ();
 sg13g2_fill_1 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_558 ();
 sg13g2_decap_8 FILLER_25_565 ();
 sg13g2_fill_1 FILLER_25_577 ();
 sg13g2_decap_4 FILLER_25_582 ();
 sg13g2_fill_2 FILLER_25_586 ();
 sg13g2_fill_1 FILLER_25_593 ();
 sg13g2_decap_8 FILLER_25_598 ();
 sg13g2_decap_8 FILLER_25_605 ();
 sg13g2_fill_2 FILLER_25_625 ();
 sg13g2_fill_2 FILLER_25_631 ();
 sg13g2_fill_1 FILLER_25_633 ();
 sg13g2_fill_2 FILLER_25_638 ();
 sg13g2_fill_1 FILLER_25_640 ();
 sg13g2_fill_2 FILLER_25_667 ();
 sg13g2_decap_8 FILLER_25_677 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_fill_1 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_719 ();
 sg13g2_decap_8 FILLER_25_726 ();
 sg13g2_fill_2 FILLER_25_733 ();
 sg13g2_fill_2 FILLER_25_739 ();
 sg13g2_fill_1 FILLER_25_746 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_fill_2 FILLER_25_768 ();
 sg13g2_fill_1 FILLER_25_770 ();
 sg13g2_decap_4 FILLER_25_807 ();
 sg13g2_decap_4 FILLER_25_815 ();
 sg13g2_fill_2 FILLER_25_838 ();
 sg13g2_fill_2 FILLER_25_858 ();
 sg13g2_decap_4 FILLER_25_866 ();
 sg13g2_fill_2 FILLER_25_870 ();
 sg13g2_fill_1 FILLER_25_907 ();
 sg13g2_decap_8 FILLER_25_913 ();
 sg13g2_decap_4 FILLER_25_920 ();
 sg13g2_fill_1 FILLER_25_936 ();
 sg13g2_fill_1 FILLER_25_942 ();
 sg13g2_decap_4 FILLER_25_951 ();
 sg13g2_fill_2 FILLER_25_955 ();
 sg13g2_decap_8 FILLER_25_962 ();
 sg13g2_decap_4 FILLER_25_969 ();
 sg13g2_fill_2 FILLER_25_973 ();
 sg13g2_decap_8 FILLER_25_997 ();
 sg13g2_decap_8 FILLER_25_1004 ();
 sg13g2_decap_4 FILLER_25_1015 ();
 sg13g2_fill_1 FILLER_25_1019 ();
 sg13g2_decap_8 FILLER_25_1032 ();
 sg13g2_decap_8 FILLER_25_1039 ();
 sg13g2_fill_2 FILLER_25_1046 ();
 sg13g2_fill_1 FILLER_25_1048 ();
 sg13g2_fill_1 FILLER_25_1058 ();
 sg13g2_fill_1 FILLER_25_1173 ();
 sg13g2_fill_2 FILLER_25_1189 ();
 sg13g2_fill_2 FILLER_25_1204 ();
 sg13g2_fill_1 FILLER_25_1206 ();
 sg13g2_decap_4 FILLER_25_1233 ();
 sg13g2_decap_4 FILLER_25_1250 ();
 sg13g2_fill_2 FILLER_25_1294 ();
 sg13g2_decap_4 FILLER_26_30 ();
 sg13g2_fill_1 FILLER_26_34 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_64 ();
 sg13g2_decap_8 FILLER_26_73 ();
 sg13g2_decap_4 FILLER_26_99 ();
 sg13g2_decap_8 FILLER_26_107 ();
 sg13g2_fill_2 FILLER_26_114 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_decap_4 FILLER_26_138 ();
 sg13g2_fill_2 FILLER_26_142 ();
 sg13g2_decap_4 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_152 ();
 sg13g2_decap_8 FILLER_26_166 ();
 sg13g2_decap_4 FILLER_26_188 ();
 sg13g2_fill_2 FILLER_26_210 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_302 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_323 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_fill_2 FILLER_26_352 ();
 sg13g2_fill_1 FILLER_26_354 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_decap_4 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_fill_2 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_391 ();
 sg13g2_fill_1 FILLER_26_452 ();
 sg13g2_decap_8 FILLER_26_566 ();
 sg13g2_fill_1 FILLER_26_573 ();
 sg13g2_decap_8 FILLER_26_578 ();
 sg13g2_fill_2 FILLER_26_585 ();
 sg13g2_fill_2 FILLER_26_613 ();
 sg13g2_decap_4 FILLER_26_641 ();
 sg13g2_decap_8 FILLER_26_649 ();
 sg13g2_decap_4 FILLER_26_656 ();
 sg13g2_fill_1 FILLER_26_660 ();
 sg13g2_fill_2 FILLER_26_671 ();
 sg13g2_fill_2 FILLER_26_704 ();
 sg13g2_fill_1 FILLER_26_706 ();
 sg13g2_fill_1 FILLER_26_741 ();
 sg13g2_fill_1 FILLER_26_746 ();
 sg13g2_fill_1 FILLER_26_751 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_fill_2 FILLER_26_763 ();
 sg13g2_fill_1 FILLER_26_770 ();
 sg13g2_fill_2 FILLER_26_774 ();
 sg13g2_fill_1 FILLER_26_776 ();
 sg13g2_decap_8 FILLER_26_785 ();
 sg13g2_fill_2 FILLER_26_792 ();
 sg13g2_fill_1 FILLER_26_794 ();
 sg13g2_fill_2 FILLER_26_844 ();
 sg13g2_fill_2 FILLER_26_863 ();
 sg13g2_decap_8 FILLER_26_869 ();
 sg13g2_decap_8 FILLER_26_876 ();
 sg13g2_decap_8 FILLER_26_883 ();
 sg13g2_fill_2 FILLER_26_890 ();
 sg13g2_fill_2 FILLER_26_901 ();
 sg13g2_fill_1 FILLER_26_903 ();
 sg13g2_fill_2 FILLER_26_933 ();
 sg13g2_fill_1 FILLER_26_935 ();
 sg13g2_fill_1 FILLER_26_941 ();
 sg13g2_fill_1 FILLER_26_946 ();
 sg13g2_fill_2 FILLER_26_955 ();
 sg13g2_fill_2 FILLER_26_993 ();
 sg13g2_decap_4 FILLER_26_1030 ();
 sg13g2_fill_2 FILLER_26_1034 ();
 sg13g2_fill_2 FILLER_26_1071 ();
 sg13g2_fill_1 FILLER_26_1073 ();
 sg13g2_decap_4 FILLER_26_1077 ();
 sg13g2_decap_8 FILLER_26_1096 ();
 sg13g2_fill_2 FILLER_26_1103 ();
 sg13g2_fill_1 FILLER_26_1105 ();
 sg13g2_fill_2 FILLER_26_1116 ();
 sg13g2_fill_1 FILLER_26_1118 ();
 sg13g2_decap_8 FILLER_26_1123 ();
 sg13g2_fill_2 FILLER_26_1130 ();
 sg13g2_fill_2 FILLER_26_1148 ();
 sg13g2_fill_1 FILLER_26_1150 ();
 sg13g2_fill_2 FILLER_26_1160 ();
 sg13g2_fill_1 FILLER_26_1172 ();
 sg13g2_fill_2 FILLER_26_1187 ();
 sg13g2_fill_2 FILLER_26_1199 ();
 sg13g2_decap_8 FILLER_26_1219 ();
 sg13g2_decap_8 FILLER_26_1226 ();
 sg13g2_fill_1 FILLER_26_1233 ();
 sg13g2_decap_8 FILLER_26_1269 ();
 sg13g2_decap_4 FILLER_26_1276 ();
 sg13g2_fill_2 FILLER_26_1280 ();
 sg13g2_fill_2 FILLER_26_1285 ();
 sg13g2_fill_1 FILLER_26_1291 ();
 sg13g2_decap_4 FILLER_26_1302 ();
 sg13g2_fill_1 FILLER_26_1306 ();
 sg13g2_decap_8 FILLER_26_1311 ();
 sg13g2_decap_8 FILLER_26_1318 ();
 sg13g2_fill_1 FILLER_26_1325 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_17 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_35 ();
 sg13g2_decap_4 FILLER_27_72 ();
 sg13g2_decap_8 FILLER_27_80 ();
 sg13g2_decap_8 FILLER_27_129 ();
 sg13g2_decap_4 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_fill_2 FILLER_27_158 ();
 sg13g2_fill_1 FILLER_27_160 ();
 sg13g2_decap_8 FILLER_27_166 ();
 sg13g2_fill_2 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_4 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_232 ();
 sg13g2_fill_2 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_1 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_303 ();
 sg13g2_fill_1 FILLER_27_305 ();
 sg13g2_fill_2 FILLER_27_365 ();
 sg13g2_fill_2 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_4 FILLER_27_413 ();
 sg13g2_fill_1 FILLER_27_417 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_decap_8 FILLER_27_442 ();
 sg13g2_fill_1 FILLER_27_449 ();
 sg13g2_decap_8 FILLER_27_454 ();
 sg13g2_decap_8 FILLER_27_461 ();
 sg13g2_fill_1 FILLER_27_468 ();
 sg13g2_decap_4 FILLER_27_478 ();
 sg13g2_fill_2 FILLER_27_486 ();
 sg13g2_decap_8 FILLER_27_492 ();
 sg13g2_decap_4 FILLER_27_499 ();
 sg13g2_fill_1 FILLER_27_503 ();
 sg13g2_fill_1 FILLER_27_508 ();
 sg13g2_fill_2 FILLER_27_513 ();
 sg13g2_fill_1 FILLER_27_520 ();
 sg13g2_fill_2 FILLER_27_527 ();
 sg13g2_decap_4 FILLER_27_533 ();
 sg13g2_fill_1 FILLER_27_537 ();
 sg13g2_decap_8 FILLER_27_542 ();
 sg13g2_decap_4 FILLER_27_549 ();
 sg13g2_fill_2 FILLER_27_553 ();
 sg13g2_fill_1 FILLER_27_589 ();
 sg13g2_decap_4 FILLER_27_606 ();
 sg13g2_fill_2 FILLER_27_610 ();
 sg13g2_decap_4 FILLER_27_616 ();
 sg13g2_fill_1 FILLER_27_624 ();
 sg13g2_fill_2 FILLER_27_629 ();
 sg13g2_fill_2 FILLER_27_665 ();
 sg13g2_fill_1 FILLER_27_667 ();
 sg13g2_decap_4 FILLER_27_676 ();
 sg13g2_fill_1 FILLER_27_680 ();
 sg13g2_fill_1 FILLER_27_688 ();
 sg13g2_decap_4 FILLER_27_693 ();
 sg13g2_fill_2 FILLER_27_697 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_fill_1 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_719 ();
 sg13g2_fill_2 FILLER_27_726 ();
 sg13g2_fill_1 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_737 ();
 sg13g2_decap_4 FILLER_27_744 ();
 sg13g2_fill_2 FILLER_27_752 ();
 sg13g2_fill_2 FILLER_27_758 ();
 sg13g2_fill_1 FILLER_27_760 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_860 ();
 sg13g2_decap_8 FILLER_27_867 ();
 sg13g2_fill_2 FILLER_27_874 ();
 sg13g2_decap_8 FILLER_27_915 ();
 sg13g2_decap_8 FILLER_27_922 ();
 sg13g2_fill_2 FILLER_27_929 ();
 sg13g2_fill_1 FILLER_27_936 ();
 sg13g2_decap_4 FILLER_27_946 ();
 sg13g2_decap_8 FILLER_27_959 ();
 sg13g2_decap_8 FILLER_27_966 ();
 sg13g2_fill_2 FILLER_27_973 ();
 sg13g2_fill_1 FILLER_27_975 ();
 sg13g2_decap_8 FILLER_27_980 ();
 sg13g2_decap_4 FILLER_27_987 ();
 sg13g2_fill_2 FILLER_27_991 ();
 sg13g2_decap_8 FILLER_27_997 ();
 sg13g2_fill_2 FILLER_27_1044 ();
 sg13g2_fill_1 FILLER_27_1046 ();
 sg13g2_decap_4 FILLER_27_1051 ();
 sg13g2_fill_2 FILLER_27_1058 ();
 sg13g2_fill_2 FILLER_27_1168 ();
 sg13g2_decap_4 FILLER_27_1200 ();
 sg13g2_fill_1 FILLER_27_1204 ();
 sg13g2_fill_1 FILLER_27_1231 ();
 sg13g2_decap_8 FILLER_27_1249 ();
 sg13g2_fill_2 FILLER_27_1256 ();
 sg13g2_fill_1 FILLER_27_1289 ();
 sg13g2_fill_1 FILLER_28_26 ();
 sg13g2_fill_1 FILLER_28_36 ();
 sg13g2_decap_4 FILLER_28_41 ();
 sg13g2_fill_2 FILLER_28_45 ();
 sg13g2_decap_4 FILLER_28_51 ();
 sg13g2_fill_1 FILLER_28_55 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_fill_2 FILLER_28_67 ();
 sg13g2_decap_4 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_decap_4 FILLER_28_110 ();
 sg13g2_fill_1 FILLER_28_114 ();
 sg13g2_fill_1 FILLER_28_141 ();
 sg13g2_decap_4 FILLER_28_180 ();
 sg13g2_fill_1 FILLER_28_184 ();
 sg13g2_fill_1 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_198 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_218 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_fill_2 FILLER_28_259 ();
 sg13g2_fill_2 FILLER_28_265 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_decap_8 FILLER_28_310 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_fill_2 FILLER_28_379 ();
 sg13g2_fill_1 FILLER_28_467 ();
 sg13g2_fill_2 FILLER_28_498 ();
 sg13g2_fill_1 FILLER_28_526 ();
 sg13g2_fill_2 FILLER_28_571 ();
 sg13g2_fill_1 FILLER_28_573 ();
 sg13g2_fill_1 FILLER_28_580 ();
 sg13g2_fill_2 FILLER_28_611 ();
 sg13g2_decap_4 FILLER_28_643 ();
 sg13g2_fill_2 FILLER_28_647 ();
 sg13g2_decap_8 FILLER_28_653 ();
 sg13g2_fill_1 FILLER_28_660 ();
 sg13g2_fill_2 FILLER_28_675 ();
 sg13g2_fill_1 FILLER_28_677 ();
 sg13g2_decap_4 FILLER_28_682 ();
 sg13g2_fill_1 FILLER_28_686 ();
 sg13g2_decap_4 FILLER_28_692 ();
 sg13g2_decap_4 FILLER_28_755 ();
 sg13g2_fill_2 FILLER_28_759 ();
 sg13g2_fill_1 FILLER_28_787 ();
 sg13g2_fill_2 FILLER_28_832 ();
 sg13g2_decap_4 FILLER_28_844 ();
 sg13g2_fill_2 FILLER_28_864 ();
 sg13g2_fill_1 FILLER_28_866 ();
 sg13g2_decap_8 FILLER_28_871 ();
 sg13g2_decap_4 FILLER_28_878 ();
 sg13g2_fill_2 FILLER_28_882 ();
 sg13g2_decap_8 FILLER_28_901 ();
 sg13g2_fill_2 FILLER_28_913 ();
 sg13g2_fill_2 FILLER_28_919 ();
 sg13g2_decap_8 FILLER_28_927 ();
 sg13g2_decap_8 FILLER_28_957 ();
 sg13g2_fill_1 FILLER_28_964 ();
 sg13g2_decap_8 FILLER_28_1012 ();
 sg13g2_fill_2 FILLER_28_1019 ();
 sg13g2_decap_8 FILLER_28_1029 ();
 sg13g2_decap_8 FILLER_28_1036 ();
 sg13g2_decap_4 FILLER_28_1043 ();
 sg13g2_fill_2 FILLER_28_1047 ();
 sg13g2_fill_2 FILLER_28_1053 ();
 sg13g2_fill_2 FILLER_28_1060 ();
 sg13g2_fill_1 FILLER_28_1062 ();
 sg13g2_fill_2 FILLER_28_1066 ();
 sg13g2_decap_4 FILLER_28_1072 ();
 sg13g2_fill_1 FILLER_28_1081 ();
 sg13g2_fill_2 FILLER_28_1091 ();
 sg13g2_fill_1 FILLER_28_1093 ();
 sg13g2_fill_1 FILLER_28_1107 ();
 sg13g2_fill_2 FILLER_28_1113 ();
 sg13g2_fill_1 FILLER_28_1115 ();
 sg13g2_fill_2 FILLER_28_1121 ();
 sg13g2_fill_1 FILLER_28_1123 ();
 sg13g2_fill_2 FILLER_28_1129 ();
 sg13g2_fill_1 FILLER_28_1131 ();
 sg13g2_decap_4 FILLER_28_1160 ();
 sg13g2_fill_2 FILLER_28_1164 ();
 sg13g2_fill_1 FILLER_28_1169 ();
 sg13g2_fill_2 FILLER_28_1179 ();
 sg13g2_decap_8 FILLER_28_1189 ();
 sg13g2_fill_2 FILLER_28_1196 ();
 sg13g2_decap_8 FILLER_28_1202 ();
 sg13g2_decap_4 FILLER_28_1209 ();
 sg13g2_fill_1 FILLER_28_1213 ();
 sg13g2_decap_8 FILLER_28_1250 ();
 sg13g2_fill_2 FILLER_28_1265 ();
 sg13g2_fill_1 FILLER_28_1267 ();
 sg13g2_fill_2 FILLER_28_1276 ();
 sg13g2_fill_1 FILLER_28_1278 ();
 sg13g2_fill_2 FILLER_28_1284 ();
 sg13g2_fill_1 FILLER_28_1286 ();
 sg13g2_fill_2 FILLER_28_1323 ();
 sg13g2_fill_1 FILLER_28_1325 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_11 ();
 sg13g2_fill_2 FILLER_29_15 ();
 sg13g2_fill_2 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_27 ();
 sg13g2_fill_1 FILLER_29_31 ();
 sg13g2_fill_1 FILLER_29_37 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_fill_2 FILLER_29_48 ();
 sg13g2_fill_2 FILLER_29_54 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_decap_4 FILLER_29_62 ();
 sg13g2_decap_4 FILLER_29_75 ();
 sg13g2_fill_2 FILLER_29_83 ();
 sg13g2_fill_2 FILLER_29_90 ();
 sg13g2_decap_4 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_116 ();
 sg13g2_fill_2 FILLER_29_122 ();
 sg13g2_fill_2 FILLER_29_131 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_147 ();
 sg13g2_decap_4 FILLER_29_153 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_168 ();
 sg13g2_fill_1 FILLER_29_170 ();
 sg13g2_decap_8 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_226 ();
 sg13g2_decap_8 FILLER_29_233 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_decap_4 FILLER_29_263 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_decap_4 FILLER_29_288 ();
 sg13g2_fill_1 FILLER_29_292 ();
 sg13g2_decap_4 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_311 ();
 sg13g2_fill_2 FILLER_29_317 ();
 sg13g2_decap_4 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_fill_2 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_8 FILLER_29_404 ();
 sg13g2_fill_2 FILLER_29_411 ();
 sg13g2_decap_4 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_453 ();
 sg13g2_fill_2 FILLER_29_460 ();
 sg13g2_fill_1 FILLER_29_462 ();
 sg13g2_fill_2 FILLER_29_469 ();
 sg13g2_fill_1 FILLER_29_479 ();
 sg13g2_decap_8 FILLER_29_484 ();
 sg13g2_decap_4 FILLER_29_491 ();
 sg13g2_fill_1 FILLER_29_495 ();
 sg13g2_fill_1 FILLER_29_504 ();
 sg13g2_fill_2 FILLER_29_509 ();
 sg13g2_fill_1 FILLER_29_511 ();
 sg13g2_fill_2 FILLER_29_517 ();
 sg13g2_fill_1 FILLER_29_519 ();
 sg13g2_fill_2 FILLER_29_530 ();
 sg13g2_fill_1 FILLER_29_532 ();
 sg13g2_fill_2 FILLER_29_537 ();
 sg13g2_decap_8 FILLER_29_548 ();
 sg13g2_fill_2 FILLER_29_555 ();
 sg13g2_fill_1 FILLER_29_557 ();
 sg13g2_fill_2 FILLER_29_578 ();
 sg13g2_decap_4 FILLER_29_586 ();
 sg13g2_fill_2 FILLER_29_590 ();
 sg13g2_fill_2 FILLER_29_600 ();
 sg13g2_fill_1 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_613 ();
 sg13g2_fill_1 FILLER_29_624 ();
 sg13g2_decap_8 FILLER_29_629 ();
 sg13g2_decap_4 FILLER_29_636 ();
 sg13g2_fill_2 FILLER_29_640 ();
 sg13g2_fill_1 FILLER_29_698 ();
 sg13g2_decap_4 FILLER_29_725 ();
 sg13g2_fill_1 FILLER_29_729 ();
 sg13g2_decap_8 FILLER_29_734 ();
 sg13g2_decap_8 FILLER_29_741 ();
 sg13g2_decap_4 FILLER_29_748 ();
 sg13g2_fill_1 FILLER_29_756 ();
 sg13g2_fill_1 FILLER_29_762 ();
 sg13g2_fill_1 FILLER_29_767 ();
 sg13g2_fill_2 FILLER_29_772 ();
 sg13g2_fill_1 FILLER_29_774 ();
 sg13g2_fill_2 FILLER_29_779 ();
 sg13g2_fill_1 FILLER_29_781 ();
 sg13g2_decap_4 FILLER_29_796 ();
 sg13g2_decap_8 FILLER_29_804 ();
 sg13g2_decap_8 FILLER_29_811 ();
 sg13g2_decap_8 FILLER_29_818 ();
 sg13g2_decap_8 FILLER_29_825 ();
 sg13g2_decap_4 FILLER_29_832 ();
 sg13g2_fill_2 FILLER_29_848 ();
 sg13g2_fill_1 FILLER_29_950 ();
 sg13g2_fill_2 FILLER_29_960 ();
 sg13g2_fill_2 FILLER_29_973 ();
 sg13g2_fill_1 FILLER_29_975 ();
 sg13g2_decap_4 FILLER_29_990 ();
 sg13g2_decap_4 FILLER_29_998 ();
 sg13g2_fill_2 FILLER_29_1002 ();
 sg13g2_decap_4 FILLER_29_1097 ();
 sg13g2_fill_2 FILLER_29_1101 ();
 sg13g2_fill_1 FILLER_29_1108 ();
 sg13g2_decap_4 FILLER_29_1119 ();
 sg13g2_fill_1 FILLER_29_1123 ();
 sg13g2_decap_4 FILLER_29_1129 ();
 sg13g2_fill_2 FILLER_29_1148 ();
 sg13g2_fill_1 FILLER_29_1150 ();
 sg13g2_fill_2 FILLER_29_1156 ();
 sg13g2_fill_2 FILLER_29_1180 ();
 sg13g2_fill_2 FILLER_29_1284 ();
 sg13g2_fill_2 FILLER_29_1295 ();
 sg13g2_fill_2 FILLER_29_1323 ();
 sg13g2_fill_1 FILLER_29_1325 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_11 ();
 sg13g2_fill_1 FILLER_30_17 ();
 sg13g2_fill_2 FILLER_30_22 ();
 sg13g2_decap_4 FILLER_30_29 ();
 sg13g2_fill_2 FILLER_30_33 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_fill_1 FILLER_30_41 ();
 sg13g2_fill_1 FILLER_30_81 ();
 sg13g2_fill_1 FILLER_30_85 ();
 sg13g2_fill_1 FILLER_30_90 ();
 sg13g2_fill_2 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_121 ();
 sg13g2_fill_2 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_187 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_fill_2 FILLER_30_194 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_fill_2 FILLER_30_281 ();
 sg13g2_decap_4 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_295 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_decap_4 FILLER_30_363 ();
 sg13g2_fill_1 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_decap_4 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_381 ();
 sg13g2_fill_1 FILLER_30_386 ();
 sg13g2_fill_2 FILLER_30_468 ();
 sg13g2_fill_1 FILLER_30_470 ();
 sg13g2_decap_8 FILLER_30_501 ();
 sg13g2_fill_1 FILLER_30_508 ();
 sg13g2_decap_4 FILLER_30_513 ();
 sg13g2_fill_2 FILLER_30_527 ();
 sg13g2_fill_1 FILLER_30_529 ();
 sg13g2_decap_4 FILLER_30_588 ();
 sg13g2_fill_1 FILLER_30_618 ();
 sg13g2_decap_8 FILLER_30_653 ();
 sg13g2_decap_8 FILLER_30_660 ();
 sg13g2_decap_8 FILLER_30_667 ();
 sg13g2_decap_8 FILLER_30_674 ();
 sg13g2_fill_1 FILLER_30_699 ();
 sg13g2_fill_2 FILLER_30_708 ();
 sg13g2_fill_1 FILLER_30_753 ();
 sg13g2_fill_2 FILLER_30_758 ();
 sg13g2_fill_2 FILLER_30_777 ();
 sg13g2_fill_2 FILLER_30_820 ();
 sg13g2_fill_1 FILLER_30_822 ();
 sg13g2_decap_8 FILLER_30_827 ();
 sg13g2_decap_4 FILLER_30_838 ();
 sg13g2_fill_1 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_decap_4 FILLER_30_861 ();
 sg13g2_fill_1 FILLER_30_865 ();
 sg13g2_decap_4 FILLER_30_882 ();
 sg13g2_fill_2 FILLER_30_886 ();
 sg13g2_fill_2 FILLER_30_893 ();
 sg13g2_decap_4 FILLER_30_899 ();
 sg13g2_fill_1 FILLER_30_903 ();
 sg13g2_fill_2 FILLER_30_908 ();
 sg13g2_fill_1 FILLER_30_910 ();
 sg13g2_decap_8 FILLER_30_916 ();
 sg13g2_decap_8 FILLER_30_931 ();
 sg13g2_fill_2 FILLER_30_967 ();
 sg13g2_fill_2 FILLER_30_995 ();
 sg13g2_decap_8 FILLER_30_1006 ();
 sg13g2_decap_8 FILLER_30_1013 ();
 sg13g2_decap_8 FILLER_30_1020 ();
 sg13g2_decap_8 FILLER_30_1027 ();
 sg13g2_decap_4 FILLER_30_1034 ();
 sg13g2_fill_2 FILLER_30_1053 ();
 sg13g2_fill_1 FILLER_30_1055 ();
 sg13g2_fill_1 FILLER_30_1060 ();
 sg13g2_decap_4 FILLER_30_1069 ();
 sg13g2_fill_2 FILLER_30_1073 ();
 sg13g2_decap_8 FILLER_30_1100 ();
 sg13g2_fill_2 FILLER_30_1112 ();
 sg13g2_fill_1 FILLER_30_1114 ();
 sg13g2_decap_4 FILLER_30_1127 ();
 sg13g2_fill_2 FILLER_30_1131 ();
 sg13g2_fill_2 FILLER_30_1145 ();
 sg13g2_fill_1 FILLER_30_1156 ();
 sg13g2_fill_2 FILLER_30_1164 ();
 sg13g2_decap_8 FILLER_30_1190 ();
 sg13g2_fill_2 FILLER_30_1197 ();
 sg13g2_decap_4 FILLER_30_1204 ();
 sg13g2_fill_2 FILLER_30_1208 ();
 sg13g2_decap_4 FILLER_30_1220 ();
 sg13g2_fill_1 FILLER_30_1224 ();
 sg13g2_fill_1 FILLER_30_1229 ();
 sg13g2_decap_8 FILLER_30_1242 ();
 sg13g2_fill_2 FILLER_30_1249 ();
 sg13g2_fill_1 FILLER_30_1251 ();
 sg13g2_decap_4 FILLER_30_1256 ();
 sg13g2_fill_1 FILLER_30_1260 ();
 sg13g2_fill_2 FILLER_30_1271 ();
 sg13g2_fill_1 FILLER_30_1273 ();
 sg13g2_fill_2 FILLER_30_1283 ();
 sg13g2_fill_1 FILLER_30_1289 ();
 sg13g2_fill_1 FILLER_31_26 ();
 sg13g2_fill_2 FILLER_31_48 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_fill_1 FILLER_31_60 ();
 sg13g2_decap_4 FILLER_31_74 ();
 sg13g2_fill_2 FILLER_31_86 ();
 sg13g2_fill_1 FILLER_31_88 ();
 sg13g2_decap_8 FILLER_31_100 ();
 sg13g2_decap_4 FILLER_31_107 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_127 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_decap_4 FILLER_31_154 ();
 sg13g2_decap_4 FILLER_31_162 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_decap_4 FILLER_31_173 ();
 sg13g2_decap_8 FILLER_31_186 ();
 sg13g2_decap_4 FILLER_31_193 ();
 sg13g2_fill_2 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_decap_8 FILLER_31_263 ();
 sg13g2_fill_2 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_277 ();
 sg13g2_decap_4 FILLER_31_284 ();
 sg13g2_fill_2 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_4 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_fill_1 FILLER_31_394 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_425 ();
 sg13g2_decap_4 FILLER_31_431 ();
 sg13g2_fill_2 FILLER_31_435 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_fill_2 FILLER_31_455 ();
 sg13g2_fill_1 FILLER_31_457 ();
 sg13g2_decap_4 FILLER_31_466 ();
 sg13g2_fill_1 FILLER_31_504 ();
 sg13g2_fill_2 FILLER_31_516 ();
 sg13g2_fill_1 FILLER_31_518 ();
 sg13g2_decap_4 FILLER_31_523 ();
 sg13g2_fill_1 FILLER_31_527 ();
 sg13g2_decap_8 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_fill_2 FILLER_31_546 ();
 sg13g2_fill_1 FILLER_31_556 ();
 sg13g2_fill_2 FILLER_31_568 ();
 sg13g2_fill_1 FILLER_31_570 ();
 sg13g2_decap_4 FILLER_31_575 ();
 sg13g2_fill_1 FILLER_31_579 ();
 sg13g2_decap_8 FILLER_31_584 ();
 sg13g2_decap_8 FILLER_31_591 ();
 sg13g2_fill_1 FILLER_31_598 ();
 sg13g2_fill_2 FILLER_31_603 ();
 sg13g2_fill_1 FILLER_31_605 ();
 sg13g2_fill_2 FILLER_31_618 ();
 sg13g2_decap_4 FILLER_31_628 ();
 sg13g2_fill_2 FILLER_31_632 ();
 sg13g2_fill_1 FILLER_31_687 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_4 FILLER_31_735 ();
 sg13g2_fill_2 FILLER_31_739 ();
 sg13g2_decap_4 FILLER_31_755 ();
 sg13g2_fill_1 FILLER_31_759 ();
 sg13g2_decap_4 FILLER_31_790 ();
 sg13g2_decap_4 FILLER_31_798 ();
 sg13g2_fill_1 FILLER_31_802 ();
 sg13g2_decap_4 FILLER_31_818 ();
 sg13g2_fill_2 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_31_828 ();
 sg13g2_decap_8 FILLER_31_839 ();
 sg13g2_fill_2 FILLER_31_846 ();
 sg13g2_decap_8 FILLER_31_852 ();
 sg13g2_decap_8 FILLER_31_859 ();
 sg13g2_fill_2 FILLER_31_866 ();
 sg13g2_decap_4 FILLER_31_881 ();
 sg13g2_fill_1 FILLER_31_944 ();
 sg13g2_fill_2 FILLER_31_950 ();
 sg13g2_fill_1 FILLER_31_952 ();
 sg13g2_fill_2 FILLER_31_958 ();
 sg13g2_decap_4 FILLER_31_972 ();
 sg13g2_fill_2 FILLER_31_976 ();
 sg13g2_fill_1 FILLER_31_991 ();
 sg13g2_decap_4 FILLER_31_1018 ();
 sg13g2_decap_4 FILLER_31_1056 ();
 sg13g2_fill_1 FILLER_31_1060 ();
 sg13g2_fill_2 FILLER_31_1065 ();
 sg13g2_fill_1 FILLER_31_1067 ();
 sg13g2_decap_8 FILLER_31_1073 ();
 sg13g2_decap_4 FILLER_31_1080 ();
 sg13g2_fill_2 FILLER_31_1084 ();
 sg13g2_decap_8 FILLER_31_1090 ();
 sg13g2_decap_8 FILLER_31_1097 ();
 sg13g2_decap_4 FILLER_31_1104 ();
 sg13g2_fill_1 FILLER_31_1108 ();
 sg13g2_decap_8 FILLER_31_1117 ();
 sg13g2_decap_8 FILLER_31_1124 ();
 sg13g2_decap_4 FILLER_31_1131 ();
 sg13g2_fill_2 FILLER_31_1135 ();
 sg13g2_fill_2 FILLER_31_1141 ();
 sg13g2_decap_8 FILLER_31_1151 ();
 sg13g2_decap_4 FILLER_31_1162 ();
 sg13g2_fill_2 FILLER_31_1166 ();
 sg13g2_fill_1 FILLER_31_1174 ();
 sg13g2_fill_2 FILLER_31_1183 ();
 sg13g2_fill_2 FILLER_31_1189 ();
 sg13g2_fill_1 FILLER_31_1217 ();
 sg13g2_fill_1 FILLER_31_1244 ();
 sg13g2_decap_4 FILLER_31_1271 ();
 sg13g2_fill_1 FILLER_31_1301 ();
 sg13g2_fill_1 FILLER_31_1310 ();
 sg13g2_decap_4 FILLER_31_1315 ();
 sg13g2_decap_4 FILLER_31_1322 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_15 ();
 sg13g2_fill_2 FILLER_32_22 ();
 sg13g2_fill_1 FILLER_32_24 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_41 ();
 sg13g2_fill_1 FILLER_32_48 ();
 sg13g2_fill_2 FILLER_32_66 ();
 sg13g2_fill_2 FILLER_32_90 ();
 sg13g2_fill_2 FILLER_32_97 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_151 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_decap_4 FILLER_32_170 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_decap_4 FILLER_32_274 ();
 sg13g2_fill_2 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_284 ();
 sg13g2_fill_2 FILLER_32_289 ();
 sg13g2_fill_1 FILLER_32_291 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_333 ();
 sg13g2_fill_2 FILLER_32_360 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_fill_2 FILLER_32_402 ();
 sg13g2_fill_2 FILLER_32_408 ();
 sg13g2_fill_1 FILLER_32_410 ();
 sg13g2_fill_2 FILLER_32_416 ();
 sg13g2_fill_2 FILLER_32_423 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_fill_1 FILLER_32_435 ();
 sg13g2_fill_2 FILLER_32_440 ();
 sg13g2_fill_1 FILLER_32_446 ();
 sg13g2_fill_1 FILLER_32_456 ();
 sg13g2_fill_1 FILLER_32_460 ();
 sg13g2_fill_2 FILLER_32_484 ();
 sg13g2_fill_1 FILLER_32_486 ();
 sg13g2_fill_2 FILLER_32_491 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_fill_1 FILLER_32_504 ();
 sg13g2_fill_2 FILLER_32_509 ();
 sg13g2_fill_1 FILLER_32_511 ();
 sg13g2_fill_1 FILLER_32_564 ();
 sg13g2_fill_2 FILLER_32_599 ();
 sg13g2_decap_8 FILLER_32_613 ();
 sg13g2_decap_8 FILLER_32_620 ();
 sg13g2_decap_4 FILLER_32_653 ();
 sg13g2_fill_1 FILLER_32_657 ();
 sg13g2_decap_8 FILLER_32_662 ();
 sg13g2_decap_8 FILLER_32_669 ();
 sg13g2_decap_4 FILLER_32_676 ();
 sg13g2_decap_4 FILLER_32_685 ();
 sg13g2_fill_1 FILLER_32_689 ();
 sg13g2_decap_8 FILLER_32_699 ();
 sg13g2_decap_8 FILLER_32_706 ();
 sg13g2_decap_4 FILLER_32_713 ();
 sg13g2_fill_1 FILLER_32_717 ();
 sg13g2_decap_4 FILLER_32_722 ();
 sg13g2_fill_2 FILLER_32_735 ();
 sg13g2_fill_2 FILLER_32_741 ();
 sg13g2_decap_8 FILLER_32_757 ();
 sg13g2_decap_4 FILLER_32_764 ();
 sg13g2_decap_4 FILLER_32_773 ();
 sg13g2_fill_1 FILLER_32_777 ();
 sg13g2_fill_2 FILLER_32_812 ();
 sg13g2_fill_1 FILLER_32_875 ();
 sg13g2_decap_8 FILLER_32_880 ();
 sg13g2_decap_4 FILLER_32_887 ();
 sg13g2_decap_4 FILLER_32_900 ();
 sg13g2_fill_2 FILLER_32_917 ();
 sg13g2_fill_1 FILLER_32_919 ();
 sg13g2_decap_8 FILLER_32_924 ();
 sg13g2_decap_4 FILLER_32_931 ();
 sg13g2_fill_2 FILLER_32_935 ();
 sg13g2_fill_1 FILLER_32_970 ();
 sg13g2_decap_4 FILLER_32_975 ();
 sg13g2_fill_2 FILLER_32_979 ();
 sg13g2_fill_1 FILLER_32_1007 ();
 sg13g2_decap_8 FILLER_32_1012 ();
 sg13g2_decap_8 FILLER_32_1019 ();
 sg13g2_fill_2 FILLER_32_1026 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_decap_8 FILLER_32_1033 ();
 sg13g2_fill_2 FILLER_32_1084 ();
 sg13g2_fill_1 FILLER_32_1135 ();
 sg13g2_decap_8 FILLER_32_1141 ();
 sg13g2_fill_1 FILLER_32_1148 ();
 sg13g2_decap_4 FILLER_32_1154 ();
 sg13g2_fill_1 FILLER_32_1158 ();
 sg13g2_fill_2 FILLER_32_1163 ();
 sg13g2_fill_2 FILLER_32_1174 ();
 sg13g2_decap_4 FILLER_32_1184 ();
 sg13g2_fill_2 FILLER_32_1198 ();
 sg13g2_fill_1 FILLER_32_1200 ();
 sg13g2_decap_8 FILLER_32_1205 ();
 sg13g2_decap_4 FILLER_32_1212 ();
 sg13g2_fill_1 FILLER_32_1216 ();
 sg13g2_decap_8 FILLER_32_1253 ();
 sg13g2_decap_4 FILLER_32_1260 ();
 sg13g2_fill_2 FILLER_32_1264 ();
 sg13g2_fill_1 FILLER_32_1271 ();
 sg13g2_fill_1 FILLER_32_1277 ();
 sg13g2_decap_4 FILLER_32_1282 ();
 sg13g2_fill_2 FILLER_32_1289 ();
 sg13g2_fill_1 FILLER_32_1291 ();
 sg13g2_decap_8 FILLER_32_1302 ();
 sg13g2_decap_8 FILLER_32_1309 ();
 sg13g2_decap_8 FILLER_32_1316 ();
 sg13g2_fill_2 FILLER_32_1323 ();
 sg13g2_fill_1 FILLER_32_1325 ();
 sg13g2_decap_4 FILLER_33_37 ();
 sg13g2_fill_1 FILLER_33_57 ();
 sg13g2_fill_2 FILLER_33_62 ();
 sg13g2_decap_8 FILLER_33_68 ();
 sg13g2_fill_2 FILLER_33_79 ();
 sg13g2_fill_2 FILLER_33_100 ();
 sg13g2_fill_1 FILLER_33_102 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_fill_1 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_4 FILLER_33_154 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_178 ();
 sg13g2_decap_4 FILLER_33_190 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_decap_4 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_212 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_258 ();
 sg13g2_decap_4 FILLER_33_264 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_361 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_decap_4 FILLER_33_406 ();
 sg13g2_decap_4 FILLER_33_456 ();
 sg13g2_fill_1 FILLER_33_460 ();
 sg13g2_fill_2 FILLER_33_468 ();
 sg13g2_fill_1 FILLER_33_470 ();
 sg13g2_fill_1 FILLER_33_474 ();
 sg13g2_decap_4 FILLER_33_483 ();
 sg13g2_fill_1 FILLER_33_487 ();
 sg13g2_decap_8 FILLER_33_492 ();
 sg13g2_fill_1 FILLER_33_499 ();
 sg13g2_fill_2 FILLER_33_504 ();
 sg13g2_fill_2 FILLER_33_518 ();
 sg13g2_decap_4 FILLER_33_524 ();
 sg13g2_fill_1 FILLER_33_537 ();
 sg13g2_fill_1 FILLER_33_551 ();
 sg13g2_fill_1 FILLER_33_570 ();
 sg13g2_fill_2 FILLER_33_575 ();
 sg13g2_fill_2 FILLER_33_584 ();
 sg13g2_decap_4 FILLER_33_589 ();
 sg13g2_fill_2 FILLER_33_593 ();
 sg13g2_fill_2 FILLER_33_617 ();
 sg13g2_decap_8 FILLER_33_645 ();
 sg13g2_fill_1 FILLER_33_652 ();
 sg13g2_fill_2 FILLER_33_691 ();
 sg13g2_fill_1 FILLER_33_753 ();
 sg13g2_fill_2 FILLER_33_780 ();
 sg13g2_fill_1 FILLER_33_782 ();
 sg13g2_decap_4 FILLER_33_787 ();
 sg13g2_fill_2 FILLER_33_791 ();
 sg13g2_fill_2 FILLER_33_797 ();
 sg13g2_fill_1 FILLER_33_799 ();
 sg13g2_fill_2 FILLER_33_810 ();
 sg13g2_decap_4 FILLER_33_816 ();
 sg13g2_fill_1 FILLER_33_820 ();
 sg13g2_decap_8 FILLER_33_825 ();
 sg13g2_decap_8 FILLER_33_832 ();
 sg13g2_decap_8 FILLER_33_839 ();
 sg13g2_fill_1 FILLER_33_846 ();
 sg13g2_fill_2 FILLER_33_855 ();
 sg13g2_fill_2 FILLER_33_872 ();
 sg13g2_fill_1 FILLER_33_874 ();
 sg13g2_fill_2 FILLER_33_885 ();
 sg13g2_fill_2 FILLER_33_892 ();
 sg13g2_fill_1 FILLER_33_894 ();
 sg13g2_fill_1 FILLER_33_935 ();
 sg13g2_fill_1 FILLER_33_941 ();
 sg13g2_fill_1 FILLER_33_955 ();
 sg13g2_fill_1 FILLER_33_964 ();
 sg13g2_fill_1 FILLER_33_970 ();
 sg13g2_fill_1 FILLER_33_979 ();
 sg13g2_fill_2 FILLER_33_985 ();
 sg13g2_fill_1 FILLER_33_1053 ();
 sg13g2_fill_2 FILLER_33_1059 ();
 sg13g2_decap_8 FILLER_33_1065 ();
 sg13g2_decap_4 FILLER_33_1072 ();
 sg13g2_fill_1 FILLER_33_1076 ();
 sg13g2_decap_4 FILLER_33_1107 ();
 sg13g2_fill_1 FILLER_33_1111 ();
 sg13g2_decap_4 FILLER_33_1117 ();
 sg13g2_fill_1 FILLER_33_1121 ();
 sg13g2_fill_2 FILLER_33_1134 ();
 sg13g2_fill_2 FILLER_33_1167 ();
 sg13g2_decap_8 FILLER_33_1175 ();
 sg13g2_decap_8 FILLER_33_1182 ();
 sg13g2_fill_1 FILLER_33_1189 ();
 sg13g2_decap_4 FILLER_33_1199 ();
 sg13g2_fill_1 FILLER_33_1208 ();
 sg13g2_decap_8 FILLER_33_1291 ();
 sg13g2_fill_2 FILLER_33_1298 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_16 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_4 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_37 ();
 sg13g2_fill_1 FILLER_34_42 ();
 sg13g2_fill_1 FILLER_34_51 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_decap_4 FILLER_34_80 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_89 ();
 sg13g2_decap_4 FILLER_34_96 ();
 sg13g2_fill_2 FILLER_34_100 ();
 sg13g2_fill_1 FILLER_34_111 ();
 sg13g2_decap_4 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_4 FILLER_34_137 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_172 ();
 sg13g2_fill_1 FILLER_34_174 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_187 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_decap_8 FILLER_34_211 ();
 sg13g2_fill_2 FILLER_34_218 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_251 ();
 sg13g2_fill_2 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_1 FILLER_34_305 ();
 sg13g2_decap_4 FILLER_34_310 ();
 sg13g2_fill_2 FILLER_34_314 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_fill_2 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_338 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_4 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_358 ();
 sg13g2_fill_1 FILLER_34_360 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_4 FILLER_34_406 ();
 sg13g2_decap_4 FILLER_34_427 ();
 sg13g2_decap_8 FILLER_34_436 ();
 sg13g2_fill_2 FILLER_34_443 ();
 sg13g2_fill_1 FILLER_34_453 ();
 sg13g2_decap_8 FILLER_34_458 ();
 sg13g2_fill_1 FILLER_34_469 ();
 sg13g2_fill_1 FILLER_34_476 ();
 sg13g2_fill_1 FILLER_34_521 ();
 sg13g2_fill_2 FILLER_34_526 ();
 sg13g2_fill_2 FILLER_34_554 ();
 sg13g2_fill_2 FILLER_34_564 ();
 sg13g2_fill_1 FILLER_34_569 ();
 sg13g2_fill_2 FILLER_34_583 ();
 sg13g2_decap_4 FILLER_34_592 ();
 sg13g2_fill_1 FILLER_34_605 ();
 sg13g2_fill_2 FILLER_34_610 ();
 sg13g2_fill_1 FILLER_34_616 ();
 sg13g2_fill_1 FILLER_34_623 ();
 sg13g2_fill_1 FILLER_34_628 ();
 sg13g2_fill_1 FILLER_34_633 ();
 sg13g2_fill_1 FILLER_34_646 ();
 sg13g2_decap_4 FILLER_34_673 ();
 sg13g2_fill_2 FILLER_34_685 ();
 sg13g2_decap_4 FILLER_34_696 ();
 sg13g2_decap_8 FILLER_34_704 ();
 sg13g2_decap_8 FILLER_34_711 ();
 sg13g2_fill_1 FILLER_34_718 ();
 sg13g2_fill_1 FILLER_34_724 ();
 sg13g2_fill_2 FILLER_34_734 ();
 sg13g2_fill_2 FILLER_34_744 ();
 sg13g2_decap_4 FILLER_34_750 ();
 sg13g2_fill_2 FILLER_34_754 ();
 sg13g2_fill_2 FILLER_34_760 ();
 sg13g2_fill_1 FILLER_34_762 ();
 sg13g2_decap_4 FILLER_34_768 ();
 sg13g2_fill_1 FILLER_34_772 ();
 sg13g2_fill_2 FILLER_34_803 ();
 sg13g2_fill_1 FILLER_34_831 ();
 sg13g2_fill_2 FILLER_34_858 ();
 sg13g2_fill_2 FILLER_34_874 ();
 sg13g2_fill_1 FILLER_34_876 ();
 sg13g2_fill_1 FILLER_34_907 ();
 sg13g2_decap_8 FILLER_34_913 ();
 sg13g2_fill_2 FILLER_34_924 ();
 sg13g2_fill_2 FILLER_34_931 ();
 sg13g2_fill_1 FILLER_34_933 ();
 sg13g2_decap_4 FILLER_34_975 ();
 sg13g2_fill_1 FILLER_34_979 ();
 sg13g2_fill_2 FILLER_34_985 ();
 sg13g2_fill_2 FILLER_34_996 ();
 sg13g2_fill_1 FILLER_34_998 ();
 sg13g2_decap_8 FILLER_34_1003 ();
 sg13g2_decap_8 FILLER_34_1010 ();
 sg13g2_decap_8 FILLER_34_1017 ();
 sg13g2_fill_1 FILLER_34_1024 ();
 sg13g2_fill_2 FILLER_34_1033 ();
 sg13g2_fill_1 FILLER_34_1035 ();
 sg13g2_fill_2 FILLER_34_1040 ();
 sg13g2_fill_1 FILLER_34_1042 ();
 sg13g2_fill_1 FILLER_34_1047 ();
 sg13g2_decap_4 FILLER_34_1087 ();
 sg13g2_fill_1 FILLER_34_1107 ();
 sg13g2_fill_2 FILLER_34_1143 ();
 sg13g2_decap_8 FILLER_34_1149 ();
 sg13g2_decap_8 FILLER_34_1156 ();
 sg13g2_fill_1 FILLER_34_1174 ();
 sg13g2_fill_2 FILLER_34_1213 ();
 sg13g2_decap_8 FILLER_34_1219 ();
 sg13g2_decap_8 FILLER_34_1226 ();
 sg13g2_decap_8 FILLER_34_1233 ();
 sg13g2_decap_4 FILLER_34_1240 ();
 sg13g2_fill_2 FILLER_34_1244 ();
 sg13g2_decap_4 FILLER_34_1250 ();
 sg13g2_fill_2 FILLER_34_1254 ();
 sg13g2_fill_2 FILLER_34_1269 ();
 sg13g2_decap_4 FILLER_34_1284 ();
 sg13g2_fill_2 FILLER_34_1288 ();
 sg13g2_decap_4 FILLER_34_1320 ();
 sg13g2_fill_2 FILLER_34_1324 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_33 ();
 sg13g2_fill_2 FILLER_35_39 ();
 sg13g2_fill_1 FILLER_35_41 ();
 sg13g2_fill_1 FILLER_35_50 ();
 sg13g2_fill_1 FILLER_35_55 ();
 sg13g2_decap_4 FILLER_35_86 ();
 sg13g2_fill_2 FILLER_35_90 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_2 FILLER_35_111 ();
 sg13g2_decap_4 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_150 ();
 sg13g2_decap_4 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_160 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_decap_4 FILLER_35_181 ();
 sg13g2_fill_2 FILLER_35_185 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_decap_4 FILLER_35_198 ();
 sg13g2_fill_1 FILLER_35_202 ();
 sg13g2_decap_8 FILLER_35_206 ();
 sg13g2_decap_4 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_217 ();
 sg13g2_fill_2 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_254 ();
 sg13g2_decap_4 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_decap_4 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_fill_2 FILLER_35_287 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_fill_2 FILLER_35_352 ();
 sg13g2_fill_1 FILLER_35_354 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_fill_1 FILLER_35_407 ();
 sg13g2_fill_1 FILLER_35_413 ();
 sg13g2_fill_1 FILLER_35_418 ();
 sg13g2_fill_2 FILLER_35_424 ();
 sg13g2_fill_2 FILLER_35_450 ();
 sg13g2_decap_4 FILLER_35_487 ();
 sg13g2_fill_2 FILLER_35_491 ();
 sg13g2_decap_8 FILLER_35_498 ();
 sg13g2_decap_8 FILLER_35_505 ();
 sg13g2_decap_4 FILLER_35_512 ();
 sg13g2_fill_2 FILLER_35_516 ();
 sg13g2_decap_4 FILLER_35_525 ();
 sg13g2_fill_2 FILLER_35_533 ();
 sg13g2_fill_2 FILLER_35_551 ();
 sg13g2_fill_1 FILLER_35_553 ();
 sg13g2_fill_2 FILLER_35_660 ();
 sg13g2_decap_4 FILLER_35_666 ();
 sg13g2_fill_2 FILLER_35_670 ();
 sg13g2_fill_1 FILLER_35_680 ();
 sg13g2_fill_2 FILLER_35_693 ();
 sg13g2_fill_1 FILLER_35_695 ();
 sg13g2_decap_8 FILLER_35_705 ();
 sg13g2_decap_4 FILLER_35_712 ();
 sg13g2_fill_2 FILLER_35_716 ();
 sg13g2_decap_8 FILLER_35_753 ();
 sg13g2_decap_8 FILLER_35_760 ();
 sg13g2_fill_2 FILLER_35_767 ();
 sg13g2_fill_1 FILLER_35_769 ();
 sg13g2_fill_1 FILLER_35_782 ();
 sg13g2_decap_4 FILLER_35_791 ();
 sg13g2_fill_2 FILLER_35_795 ();
 sg13g2_decap_8 FILLER_35_815 ();
 sg13g2_fill_2 FILLER_35_822 ();
 sg13g2_decap_8 FILLER_35_828 ();
 sg13g2_fill_2 FILLER_35_835 ();
 sg13g2_fill_1 FILLER_35_837 ();
 sg13g2_decap_4 FILLER_35_842 ();
 sg13g2_fill_2 FILLER_35_857 ();
 sg13g2_decap_8 FILLER_35_872 ();
 sg13g2_decap_8 FILLER_35_879 ();
 sg13g2_decap_4 FILLER_35_886 ();
 sg13g2_fill_1 FILLER_35_933 ();
 sg13g2_decap_4 FILLER_35_939 ();
 sg13g2_fill_1 FILLER_35_953 ();
 sg13g2_fill_1 FILLER_35_964 ();
 sg13g2_decap_8 FILLER_35_968 ();
 sg13g2_decap_8 FILLER_35_975 ();
 sg13g2_fill_1 FILLER_35_987 ();
 sg13g2_decap_4 FILLER_35_1014 ();
 sg13g2_fill_2 FILLER_35_1018 ();
 sg13g2_decap_4 FILLER_35_1024 ();
 sg13g2_decap_4 FILLER_35_1032 ();
 sg13g2_fill_1 FILLER_35_1036 ();
 sg13g2_decap_8 FILLER_35_1051 ();
 sg13g2_decap_4 FILLER_35_1058 ();
 sg13g2_fill_1 FILLER_35_1062 ();
 sg13g2_decap_8 FILLER_35_1067 ();
 sg13g2_decap_4 FILLER_35_1074 ();
 sg13g2_fill_1 FILLER_35_1078 ();
 sg13g2_decap_4 FILLER_35_1087 ();
 sg13g2_fill_2 FILLER_35_1091 ();
 sg13g2_fill_2 FILLER_35_1103 ();
 sg13g2_decap_4 FILLER_35_1115 ();
 sg13g2_decap_4 FILLER_35_1129 ();
 sg13g2_fill_2 FILLER_35_1136 ();
 sg13g2_decap_8 FILLER_35_1159 ();
 sg13g2_decap_8 FILLER_35_1166 ();
 sg13g2_fill_2 FILLER_35_1173 ();
 sg13g2_fill_1 FILLER_35_1188 ();
 sg13g2_decap_4 FILLER_35_1196 ();
 sg13g2_decap_4 FILLER_35_1204 ();
 sg13g2_fill_2 FILLER_35_1208 ();
 sg13g2_fill_1 FILLER_35_1214 ();
 sg13g2_fill_1 FILLER_35_1219 ();
 sg13g2_fill_1 FILLER_35_1225 ();
 sg13g2_decap_4 FILLER_35_1252 ();
 sg13g2_fill_2 FILLER_35_1256 ();
 sg13g2_decap_4 FILLER_35_1284 ();
 sg13g2_fill_1 FILLER_35_1288 ();
 sg13g2_decap_8 FILLER_35_1315 ();
 sg13g2_decap_4 FILLER_35_1322 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_15 ();
 sg13g2_fill_2 FILLER_36_22 ();
 sg13g2_fill_1 FILLER_36_24 ();
 sg13g2_fill_1 FILLER_36_34 ();
 sg13g2_fill_1 FILLER_36_40 ();
 sg13g2_fill_1 FILLER_36_51 ();
 sg13g2_decap_4 FILLER_36_57 ();
 sg13g2_decap_4 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_78 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_fill_2 FILLER_36_101 ();
 sg13g2_fill_2 FILLER_36_116 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_fill_1 FILLER_36_129 ();
 sg13g2_fill_2 FILLER_36_137 ();
 sg13g2_fill_2 FILLER_36_144 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_decap_4 FILLER_36_177 ();
 sg13g2_fill_1 FILLER_36_181 ();
 sg13g2_fill_2 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_290 ();
 sg13g2_decap_8 FILLER_36_297 ();
 sg13g2_decap_8 FILLER_36_304 ();
 sg13g2_fill_2 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_decap_4 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_fill_2 FILLER_36_349 ();
 sg13g2_decap_8 FILLER_36_377 ();
 sg13g2_fill_2 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_8 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_410 ();
 sg13g2_fill_2 FILLER_36_415 ();
 sg13g2_fill_1 FILLER_36_421 ();
 sg13g2_decap_8 FILLER_36_430 ();
 sg13g2_decap_4 FILLER_36_437 ();
 sg13g2_fill_1 FILLER_36_441 ();
 sg13g2_fill_2 FILLER_36_450 ();
 sg13g2_fill_1 FILLER_36_452 ();
 sg13g2_fill_2 FILLER_36_464 ();
 sg13g2_fill_1 FILLER_36_466 ();
 sg13g2_fill_1 FILLER_36_493 ();
 sg13g2_decap_4 FILLER_36_533 ();
 sg13g2_fill_1 FILLER_36_537 ();
 sg13g2_fill_2 FILLER_36_544 ();
 sg13g2_decap_4 FILLER_36_554 ();
 sg13g2_fill_2 FILLER_36_558 ();
 sg13g2_fill_2 FILLER_36_568 ();
 sg13g2_fill_1 FILLER_36_585 ();
 sg13g2_fill_2 FILLER_36_590 ();
 sg13g2_fill_2 FILLER_36_597 ();
 sg13g2_fill_1 FILLER_36_599 ();
 sg13g2_decap_4 FILLER_36_614 ();
 sg13g2_fill_1 FILLER_36_618 ();
 sg13g2_decap_8 FILLER_36_623 ();
 sg13g2_decap_4 FILLER_36_630 ();
 sg13g2_fill_2 FILLER_36_634 ();
 sg13g2_decap_8 FILLER_36_640 ();
 sg13g2_decap_8 FILLER_36_647 ();
 sg13g2_fill_1 FILLER_36_654 ();
 sg13g2_fill_2 FILLER_36_681 ();
 sg13g2_fill_1 FILLER_36_683 ();
 sg13g2_decap_4 FILLER_36_738 ();
 sg13g2_fill_1 FILLER_36_865 ();
 sg13g2_fill_2 FILLER_36_870 ();
 sg13g2_fill_1 FILLER_36_872 ();
 sg13g2_decap_4 FILLER_36_902 ();
 sg13g2_fill_1 FILLER_36_906 ();
 sg13g2_decap_4 FILLER_36_912 ();
 sg13g2_fill_1 FILLER_36_916 ();
 sg13g2_decap_8 FILLER_36_925 ();
 sg13g2_decap_8 FILLER_36_932 ();
 sg13g2_fill_1 FILLER_36_943 ();
 sg13g2_decap_4 FILLER_36_949 ();
 sg13g2_decap_4 FILLER_36_957 ();
 sg13g2_fill_2 FILLER_36_961 ();
 sg13g2_decap_8 FILLER_36_981 ();
 sg13g2_decap_8 FILLER_36_988 ();
 sg13g2_fill_2 FILLER_36_995 ();
 sg13g2_decap_4 FILLER_36_1002 ();
 sg13g2_fill_2 FILLER_36_1006 ();
 sg13g2_decap_4 FILLER_36_1012 ();
 sg13g2_fill_2 FILLER_36_1148 ();
 sg13g2_fill_1 FILLER_36_1150 ();
 sg13g2_fill_1 FILLER_36_1158 ();
 sg13g2_fill_1 FILLER_36_1162 ();
 sg13g2_decap_4 FILLER_36_1175 ();
 sg13g2_fill_1 FILLER_36_1179 ();
 sg13g2_decap_4 FILLER_36_1188 ();
 sg13g2_fill_2 FILLER_36_1227 ();
 sg13g2_decap_8 FILLER_36_1255 ();
 sg13g2_fill_1 FILLER_36_1271 ();
 sg13g2_decap_8 FILLER_36_1275 ();
 sg13g2_decap_4 FILLER_36_1282 ();
 sg13g2_fill_1 FILLER_36_1286 ();
 sg13g2_fill_2 FILLER_36_1323 ();
 sg13g2_fill_1 FILLER_36_1325 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_27 ();
 sg13g2_fill_2 FILLER_37_37 ();
 sg13g2_fill_2 FILLER_37_43 ();
 sg13g2_fill_1 FILLER_37_45 ();
 sg13g2_fill_2 FILLER_37_50 ();
 sg13g2_fill_1 FILLER_37_52 ();
 sg13g2_fill_1 FILLER_37_57 ();
 sg13g2_fill_2 FILLER_37_63 ();
 sg13g2_decap_4 FILLER_37_74 ();
 sg13g2_fill_1 FILLER_37_78 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_decap_8 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_fill_1 FILLER_37_161 ();
 sg13g2_fill_1 FILLER_37_170 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_fill_1 FILLER_37_193 ();
 sg13g2_decap_4 FILLER_37_209 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_218 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_decap_4 FILLER_37_235 ();
 sg13g2_fill_1 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_281 ();
 sg13g2_fill_2 FILLER_37_309 ();
 sg13g2_decap_4 FILLER_37_315 ();
 sg13g2_fill_2 FILLER_37_319 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_decap_8 FILLER_37_338 ();
 sg13g2_decap_8 FILLER_37_345 ();
 sg13g2_decap_4 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_356 ();
 sg13g2_decap_4 FILLER_37_362 ();
 sg13g2_fill_2 FILLER_37_392 ();
 sg13g2_fill_1 FILLER_37_411 ();
 sg13g2_decap_8 FILLER_37_419 ();
 sg13g2_fill_2 FILLER_37_426 ();
 sg13g2_fill_2 FILLER_37_438 ();
 sg13g2_fill_2 FILLER_37_445 ();
 sg13g2_fill_2 FILLER_37_451 ();
 sg13g2_decap_8 FILLER_37_467 ();
 sg13g2_fill_2 FILLER_37_474 ();
 sg13g2_fill_1 FILLER_37_476 ();
 sg13g2_fill_2 FILLER_37_499 ();
 sg13g2_decap_4 FILLER_37_505 ();
 sg13g2_fill_2 FILLER_37_535 ();
 sg13g2_decap_4 FILLER_37_542 ();
 sg13g2_fill_1 FILLER_37_546 ();
 sg13g2_decap_4 FILLER_37_555 ();
 sg13g2_decap_8 FILLER_37_565 ();
 sg13g2_decap_4 FILLER_37_572 ();
 sg13g2_decap_8 FILLER_37_605 ();
 sg13g2_fill_2 FILLER_37_612 ();
 sg13g2_fill_1 FILLER_37_614 ();
 sg13g2_fill_1 FILLER_37_631 ();
 sg13g2_fill_2 FILLER_37_658 ();
 sg13g2_decap_4 FILLER_37_664 ();
 sg13g2_fill_1 FILLER_37_672 ();
 sg13g2_decap_4 FILLER_37_687 ();
 sg13g2_decap_8 FILLER_37_695 ();
 sg13g2_decap_4 FILLER_37_702 ();
 sg13g2_fill_1 FILLER_37_706 ();
 sg13g2_decap_8 FILLER_37_766 ();
 sg13g2_decap_8 FILLER_37_773 ();
 sg13g2_decap_8 FILLER_37_792 ();
 sg13g2_decap_8 FILLER_37_799 ();
 sg13g2_decap_4 FILLER_37_806 ();
 sg13g2_fill_2 FILLER_37_810 ();
 sg13g2_decap_4 FILLER_37_820 ();
 sg13g2_fill_1 FILLER_37_824 ();
 sg13g2_fill_2 FILLER_37_828 ();
 sg13g2_fill_1 FILLER_37_830 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_4 FILLER_37_847 ();
 sg13g2_fill_1 FILLER_37_851 ();
 sg13g2_decap_8 FILLER_37_863 ();
 sg13g2_decap_8 FILLER_37_870 ();
 sg13g2_fill_2 FILLER_37_877 ();
 sg13g2_fill_1 FILLER_37_879 ();
 sg13g2_fill_1 FILLER_37_884 ();
 sg13g2_decap_8 FILLER_37_893 ();
 sg13g2_fill_2 FILLER_37_911 ();
 sg13g2_fill_1 FILLER_37_913 ();
 sg13g2_fill_2 FILLER_37_951 ();
 sg13g2_decap_8 FILLER_37_957 ();
 sg13g2_fill_1 FILLER_37_964 ();
 sg13g2_fill_1 FILLER_37_970 ();
 sg13g2_decap_4 FILLER_37_986 ();
 sg13g2_fill_1 FILLER_37_990 ();
 sg13g2_fill_2 FILLER_37_1027 ();
 sg13g2_fill_1 FILLER_37_1029 ();
 sg13g2_decap_4 FILLER_37_1034 ();
 sg13g2_fill_2 FILLER_37_1038 ();
 sg13g2_fill_1 FILLER_37_1059 ();
 sg13g2_fill_2 FILLER_37_1064 ();
 sg13g2_fill_1 FILLER_37_1066 ();
 sg13g2_decap_4 FILLER_37_1071 ();
 sg13g2_fill_2 FILLER_37_1075 ();
 sg13g2_decap_8 FILLER_37_1081 ();
 sg13g2_fill_1 FILLER_37_1088 ();
 sg13g2_decap_4 FILLER_37_1096 ();
 sg13g2_fill_1 FILLER_37_1100 ();
 sg13g2_fill_1 FILLER_37_1107 ();
 sg13g2_fill_2 FILLER_37_1118 ();
 sg13g2_fill_2 FILLER_37_1129 ();
 sg13g2_fill_1 FILLER_37_1134 ();
 sg13g2_decap_8 FILLER_37_1138 ();
 sg13g2_decap_8 FILLER_37_1145 ();
 sg13g2_fill_1 FILLER_37_1156 ();
 sg13g2_fill_2 FILLER_37_1161 ();
 sg13g2_decap_4 FILLER_37_1167 ();
 sg13g2_fill_2 FILLER_37_1171 ();
 sg13g2_decap_4 FILLER_37_1176 ();
 sg13g2_fill_2 FILLER_37_1180 ();
 sg13g2_decap_4 FILLER_37_1198 ();
 sg13g2_decap_4 FILLER_37_1215 ();
 sg13g2_fill_2 FILLER_37_1219 ();
 sg13g2_decap_8 FILLER_37_1226 ();
 sg13g2_decap_8 FILLER_37_1241 ();
 sg13g2_decap_4 FILLER_37_1248 ();
 sg13g2_fill_1 FILLER_37_1252 ();
 sg13g2_fill_1 FILLER_37_1283 ();
 sg13g2_decap_4 FILLER_37_1320 ();
 sg13g2_fill_2 FILLER_37_1324 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_11 ();
 sg13g2_fill_2 FILLER_38_15 ();
 sg13g2_decap_8 FILLER_38_43 ();
 sg13g2_decap_4 FILLER_38_75 ();
 sg13g2_fill_2 FILLER_38_88 ();
 sg13g2_decap_4 FILLER_38_94 ();
 sg13g2_fill_1 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_110 ();
 sg13g2_decap_8 FILLER_38_117 ();
 sg13g2_decap_8 FILLER_38_124 ();
 sg13g2_decap_8 FILLER_38_136 ();
 sg13g2_fill_2 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_145 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_fill_2 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_183 ();
 sg13g2_fill_2 FILLER_38_195 ();
 sg13g2_fill_2 FILLER_38_202 ();
 sg13g2_fill_1 FILLER_38_204 ();
 sg13g2_fill_2 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_211 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_fill_2 FILLER_38_226 ();
 sg13g2_fill_1 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_234 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_fill_2 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_271 ();
 sg13g2_fill_2 FILLER_38_284 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_303 ();
 sg13g2_fill_2 FILLER_38_330 ();
 sg13g2_fill_1 FILLER_38_332 ();
 sg13g2_decap_8 FILLER_38_359 ();
 sg13g2_decap_4 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_4 FILLER_38_382 ();
 sg13g2_fill_2 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_fill_1 FILLER_38_435 ();
 sg13g2_fill_2 FILLER_38_466 ();
 sg13g2_fill_1 FILLER_38_491 ();
 sg13g2_fill_1 FILLER_38_497 ();
 sg13g2_fill_1 FILLER_38_502 ();
 sg13g2_fill_1 FILLER_38_510 ();
 sg13g2_fill_2 FILLER_38_527 ();
 sg13g2_fill_1 FILLER_38_529 ();
 sg13g2_fill_2 FILLER_38_533 ();
 sg13g2_fill_1 FILLER_38_535 ();
 sg13g2_decap_4 FILLER_38_540 ();
 sg13g2_decap_8 FILLER_38_583 ();
 sg13g2_decap_4 FILLER_38_590 ();
 sg13g2_fill_2 FILLER_38_594 ();
 sg13g2_decap_4 FILLER_38_605 ();
 sg13g2_decap_8 FILLER_38_613 ();
 sg13g2_decap_4 FILLER_38_620 ();
 sg13g2_decap_4 FILLER_38_632 ();
 sg13g2_fill_2 FILLER_38_636 ();
 sg13g2_decap_8 FILLER_38_646 ();
 sg13g2_fill_1 FILLER_38_653 ();
 sg13g2_decap_4 FILLER_38_680 ();
 sg13g2_fill_2 FILLER_38_710 ();
 sg13g2_fill_1 FILLER_38_712 ();
 sg13g2_fill_1 FILLER_38_722 ();
 sg13g2_fill_2 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_fill_1 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_747 ();
 sg13g2_decap_4 FILLER_38_754 ();
 sg13g2_fill_2 FILLER_38_758 ();
 sg13g2_decap_8 FILLER_38_769 ();
 sg13g2_fill_2 FILLER_38_832 ();
 sg13g2_fill_1 FILLER_38_834 ();
 sg13g2_decap_8 FILLER_38_843 ();
 sg13g2_decap_4 FILLER_38_850 ();
 sg13g2_fill_1 FILLER_38_871 ();
 sg13g2_fill_1 FILLER_38_906 ();
 sg13g2_fill_1 FILLER_38_912 ();
 sg13g2_fill_1 FILLER_38_942 ();
 sg13g2_decap_4 FILLER_38_969 ();
 sg13g2_fill_2 FILLER_38_1003 ();
 sg13g2_fill_1 FILLER_38_1005 ();
 sg13g2_decap_8 FILLER_38_1010 ();
 sg13g2_decap_8 FILLER_38_1017 ();
 sg13g2_decap_4 FILLER_38_1076 ();
 sg13g2_fill_2 FILLER_38_1080 ();
 sg13g2_fill_2 FILLER_38_1087 ();
 sg13g2_fill_2 FILLER_38_1093 ();
 sg13g2_fill_2 FILLER_38_1099 ();
 sg13g2_decap_4 FILLER_38_1111 ();
 sg13g2_fill_1 FILLER_38_1119 ();
 sg13g2_fill_2 FILLER_38_1126 ();
 sg13g2_fill_1 FILLER_38_1128 ();
 sg13g2_fill_2 FILLER_38_1155 ();
 sg13g2_fill_1 FILLER_38_1165 ();
 sg13g2_fill_1 FILLER_38_1170 ();
 sg13g2_decap_8 FILLER_38_1176 ();
 sg13g2_fill_2 FILLER_38_1209 ();
 sg13g2_fill_2 FILLER_38_1242 ();
 sg13g2_decap_4 FILLER_38_1256 ();
 sg13g2_fill_1 FILLER_38_1260 ();
 sg13g2_fill_1 FILLER_38_1271 ();
 sg13g2_decap_4 FILLER_38_1276 ();
 sg13g2_fill_2 FILLER_38_1293 ();
 sg13g2_fill_1 FILLER_38_1295 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_27 ();
 sg13g2_decap_4 FILLER_39_33 ();
 sg13g2_fill_2 FILLER_39_45 ();
 sg13g2_fill_2 FILLER_39_53 ();
 sg13g2_fill_2 FILLER_39_59 ();
 sg13g2_fill_1 FILLER_39_99 ();
 sg13g2_fill_1 FILLER_39_107 ();
 sg13g2_decap_8 FILLER_39_114 ();
 sg13g2_fill_2 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_132 ();
 sg13g2_fill_1 FILLER_39_138 ();
 sg13g2_fill_1 FILLER_39_145 ();
 sg13g2_fill_1 FILLER_39_151 ();
 sg13g2_fill_1 FILLER_39_167 ();
 sg13g2_fill_2 FILLER_39_182 ();
 sg13g2_fill_2 FILLER_39_193 ();
 sg13g2_fill_1 FILLER_39_200 ();
 sg13g2_fill_2 FILLER_39_227 ();
 sg13g2_fill_1 FILLER_39_229 ();
 sg13g2_fill_1 FILLER_39_256 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_fill_1 FILLER_39_292 ();
 sg13g2_fill_2 FILLER_39_309 ();
 sg13g2_decap_4 FILLER_39_320 ();
 sg13g2_fill_1 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_330 ();
 sg13g2_fill_2 FILLER_39_337 ();
 sg13g2_decap_4 FILLER_39_343 ();
 sg13g2_fill_2 FILLER_39_367 ();
 sg13g2_decap_4 FILLER_39_373 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_decap_8 FILLER_39_383 ();
 sg13g2_decap_4 FILLER_39_390 ();
 sg13g2_fill_1 FILLER_39_394 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_4 FILLER_39_406 ();
 sg13g2_fill_2 FILLER_39_410 ();
 sg13g2_fill_2 FILLER_39_416 ();
 sg13g2_fill_1 FILLER_39_418 ();
 sg13g2_decap_8 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_39_439 ();
 sg13g2_decap_8 FILLER_39_446 ();
 sg13g2_decap_8 FILLER_39_453 ();
 sg13g2_decap_4 FILLER_39_460 ();
 sg13g2_fill_1 FILLER_39_464 ();
 sg13g2_decap_4 FILLER_39_469 ();
 sg13g2_fill_2 FILLER_39_473 ();
 sg13g2_decap_8 FILLER_39_517 ();
 sg13g2_decap_8 FILLER_39_524 ();
 sg13g2_decap_8 FILLER_39_536 ();
 sg13g2_decap_8 FILLER_39_543 ();
 sg13g2_decap_8 FILLER_39_550 ();
 sg13g2_decap_8 FILLER_39_557 ();
 sg13g2_fill_2 FILLER_39_564 ();
 sg13g2_fill_1 FILLER_39_566 ();
 sg13g2_decap_8 FILLER_39_571 ();
 sg13g2_fill_2 FILLER_39_578 ();
 sg13g2_fill_1 FILLER_39_580 ();
 sg13g2_fill_2 FILLER_39_589 ();
 sg13g2_fill_1 FILLER_39_600 ();
 sg13g2_decap_4 FILLER_39_605 ();
 sg13g2_decap_4 FILLER_39_613 ();
 sg13g2_fill_2 FILLER_39_621 ();
 sg13g2_fill_1 FILLER_39_627 ();
 sg13g2_decap_8 FILLER_39_658 ();
 sg13g2_decap_4 FILLER_39_665 ();
 sg13g2_fill_2 FILLER_39_669 ();
 sg13g2_decap_4 FILLER_39_675 ();
 sg13g2_fill_1 FILLER_39_679 ();
 sg13g2_decap_4 FILLER_39_685 ();
 sg13g2_fill_1 FILLER_39_689 ();
 sg13g2_fill_2 FILLER_39_695 ();
 sg13g2_fill_1 FILLER_39_697 ();
 sg13g2_decap_4 FILLER_39_702 ();
 sg13g2_fill_1 FILLER_39_706 ();
 sg13g2_decap_8 FILLER_39_712 ();
 sg13g2_decap_4 FILLER_39_723 ();
 sg13g2_fill_1 FILLER_39_731 ();
 sg13g2_decap_4 FILLER_39_736 ();
 sg13g2_fill_1 FILLER_39_740 ();
 sg13g2_decap_8 FILLER_39_746 ();
 sg13g2_decap_8 FILLER_39_783 ();
 sg13g2_decap_8 FILLER_39_790 ();
 sg13g2_decap_4 FILLER_39_797 ();
 sg13g2_fill_1 FILLER_39_801 ();
 sg13g2_fill_1 FILLER_39_811 ();
 sg13g2_decap_8 FILLER_39_820 ();
 sg13g2_decap_4 FILLER_39_827 ();
 sg13g2_fill_2 FILLER_39_831 ();
 sg13g2_fill_1 FILLER_39_854 ();
 sg13g2_fill_1 FILLER_39_859 ();
 sg13g2_decap_8 FILLER_39_864 ();
 sg13g2_decap_4 FILLER_39_871 ();
 sg13g2_decap_4 FILLER_39_880 ();
 sg13g2_decap_4 FILLER_39_888 ();
 sg13g2_decap_8 FILLER_39_901 ();
 sg13g2_fill_1 FILLER_39_908 ();
 sg13g2_fill_1 FILLER_39_920 ();
 sg13g2_fill_2 FILLER_39_931 ();
 sg13g2_fill_1 FILLER_39_937 ();
 sg13g2_fill_2 FILLER_39_951 ();
 sg13g2_fill_2 FILLER_39_962 ();
 sg13g2_decap_8 FILLER_39_967 ();
 sg13g2_decap_4 FILLER_39_974 ();
 sg13g2_fill_2 FILLER_39_978 ();
 sg13g2_decap_4 FILLER_39_984 ();
 sg13g2_fill_1 FILLER_39_988 ();
 sg13g2_fill_1 FILLER_39_993 ();
 sg13g2_fill_1 FILLER_39_1030 ();
 sg13g2_decap_8 FILLER_39_1035 ();
 sg13g2_fill_2 FILLER_39_1042 ();
 sg13g2_fill_1 FILLER_39_1044 ();
 sg13g2_fill_2 FILLER_39_1054 ();
 sg13g2_fill_1 FILLER_39_1056 ();
 sg13g2_fill_2 FILLER_39_1156 ();
 sg13g2_fill_1 FILLER_39_1158 ();
 sg13g2_fill_1 FILLER_39_1174 ();
 sg13g2_fill_2 FILLER_39_1178 ();
 sg13g2_fill_1 FILLER_39_1180 ();
 sg13g2_fill_2 FILLER_39_1185 ();
 sg13g2_fill_2 FILLER_39_1213 ();
 sg13g2_decap_4 FILLER_39_1219 ();
 sg13g2_fill_2 FILLER_39_1223 ();
 sg13g2_decap_4 FILLER_39_1229 ();
 sg13g2_fill_2 FILLER_39_1233 ();
 sg13g2_decap_4 FILLER_39_1302 ();
 sg13g2_fill_1 FILLER_39_1306 ();
 sg13g2_decap_8 FILLER_39_1315 ();
 sg13g2_decap_4 FILLER_39_1322 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_15 ();
 sg13g2_fill_1 FILLER_40_22 ();
 sg13g2_decap_4 FILLER_40_28 ();
 sg13g2_fill_2 FILLER_40_54 ();
 sg13g2_fill_1 FILLER_40_56 ();
 sg13g2_decap_4 FILLER_40_62 ();
 sg13g2_fill_1 FILLER_40_66 ();
 sg13g2_decap_4 FILLER_40_71 ();
 sg13g2_fill_1 FILLER_40_75 ();
 sg13g2_fill_2 FILLER_40_80 ();
 sg13g2_fill_1 FILLER_40_82 ();
 sg13g2_fill_1 FILLER_40_93 ();
 sg13g2_decap_4 FILLER_40_126 ();
 sg13g2_fill_2 FILLER_40_130 ();
 sg13g2_fill_2 FILLER_40_138 ();
 sg13g2_fill_1 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_4 FILLER_40_154 ();
 sg13g2_fill_1 FILLER_40_158 ();
 sg13g2_decap_4 FILLER_40_169 ();
 sg13g2_fill_1 FILLER_40_178 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_4 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_211 ();
 sg13g2_fill_2 FILLER_40_218 ();
 sg13g2_decap_4 FILLER_40_229 ();
 sg13g2_fill_2 FILLER_40_233 ();
 sg13g2_decap_8 FILLER_40_239 ();
 sg13g2_fill_1 FILLER_40_246 ();
 sg13g2_decap_4 FILLER_40_260 ();
 sg13g2_fill_1 FILLER_40_264 ();
 sg13g2_fill_1 FILLER_40_269 ();
 sg13g2_decap_4 FILLER_40_284 ();
 sg13g2_fill_2 FILLER_40_288 ();
 sg13g2_fill_1 FILLER_40_312 ();
 sg13g2_fill_1 FILLER_40_322 ();
 sg13g2_fill_1 FILLER_40_418 ();
 sg13g2_fill_2 FILLER_40_425 ();
 sg13g2_fill_1 FILLER_40_433 ();
 sg13g2_fill_1 FILLER_40_438 ();
 sg13g2_fill_1 FILLER_40_445 ();
 sg13g2_fill_1 FILLER_40_450 ();
 sg13g2_decap_8 FILLER_40_459 ();
 sg13g2_decap_4 FILLER_40_470 ();
 sg13g2_fill_2 FILLER_40_477 ();
 sg13g2_fill_2 FILLER_40_492 ();
 sg13g2_decap_8 FILLER_40_498 ();
 sg13g2_decap_8 FILLER_40_505 ();
 sg13g2_decap_4 FILLER_40_512 ();
 sg13g2_fill_2 FILLER_40_520 ();
 sg13g2_decap_8 FILLER_40_548 ();
 sg13g2_fill_2 FILLER_40_563 ();
 sg13g2_fill_1 FILLER_40_565 ();
 sg13g2_decap_8 FILLER_40_578 ();
 sg13g2_decap_8 FILLER_40_585 ();
 sg13g2_fill_1 FILLER_40_596 ();
 sg13g2_fill_2 FILLER_40_622 ();
 sg13g2_fill_2 FILLER_40_632 ();
 sg13g2_decap_8 FILLER_40_638 ();
 sg13g2_decap_4 FILLER_40_645 ();
 sg13g2_fill_2 FILLER_40_733 ();
 sg13g2_decap_4 FILLER_40_791 ();
 sg13g2_fill_1 FILLER_40_795 ();
 sg13g2_decap_8 FILLER_40_822 ();
 sg13g2_decap_4 FILLER_40_829 ();
 sg13g2_fill_1 FILLER_40_833 ();
 sg13g2_fill_2 FILLER_40_864 ();
 sg13g2_fill_2 FILLER_40_874 ();
 sg13g2_fill_1 FILLER_40_876 ();
 sg13g2_decap_8 FILLER_40_887 ();
 sg13g2_decap_8 FILLER_40_894 ();
 sg13g2_decap_8 FILLER_40_901 ();
 sg13g2_decap_8 FILLER_40_908 ();
 sg13g2_decap_8 FILLER_40_915 ();
 sg13g2_decap_8 FILLER_40_922 ();
 sg13g2_fill_2 FILLER_40_929 ();
 sg13g2_fill_2 FILLER_40_936 ();
 sg13g2_fill_2 FILLER_40_1000 ();
 sg13g2_fill_1 FILLER_40_1002 ();
 sg13g2_decap_8 FILLER_40_1007 ();
 sg13g2_decap_8 FILLER_40_1014 ();
 sg13g2_decap_8 FILLER_40_1056 ();
 sg13g2_fill_2 FILLER_40_1063 ();
 sg13g2_fill_1 FILLER_40_1065 ();
 sg13g2_decap_8 FILLER_40_1070 ();
 sg13g2_decap_4 FILLER_40_1077 ();
 sg13g2_fill_2 FILLER_40_1081 ();
 sg13g2_fill_1 FILLER_40_1087 ();
 sg13g2_fill_1 FILLER_40_1098 ();
 sg13g2_decap_8 FILLER_40_1103 ();
 sg13g2_decap_8 FILLER_40_1110 ();
 sg13g2_decap_8 FILLER_40_1117 ();
 sg13g2_decap_4 FILLER_40_1124 ();
 sg13g2_fill_1 FILLER_40_1138 ();
 sg13g2_fill_2 FILLER_40_1145 ();
 sg13g2_fill_2 FILLER_40_1151 ();
 sg13g2_fill_1 FILLER_40_1156 ();
 sg13g2_fill_1 FILLER_40_1161 ();
 sg13g2_fill_1 FILLER_40_1173 ();
 sg13g2_decap_4 FILLER_40_1177 ();
 sg13g2_fill_1 FILLER_40_1181 ();
 sg13g2_fill_2 FILLER_40_1191 ();
 sg13g2_fill_2 FILLER_40_1204 ();
 sg13g2_fill_1 FILLER_40_1206 ();
 sg13g2_fill_2 FILLER_40_1212 ();
 sg13g2_fill_1 FILLER_40_1214 ();
 sg13g2_decap_4 FILLER_40_1249 ();
 sg13g2_fill_2 FILLER_40_1253 ();
 sg13g2_decap_8 FILLER_40_1263 ();
 sg13g2_fill_2 FILLER_40_1270 ();
 sg13g2_fill_1 FILLER_40_1272 ();
 sg13g2_decap_4 FILLER_40_1277 ();
 sg13g2_fill_1 FILLER_41_34 ();
 sg13g2_fill_2 FILLER_41_40 ();
 sg13g2_fill_1 FILLER_41_46 ();
 sg13g2_decap_8 FILLER_41_52 ();
 sg13g2_decap_8 FILLER_41_59 ();
 sg13g2_decap_4 FILLER_41_66 ();
 sg13g2_fill_2 FILLER_41_76 ();
 sg13g2_decap_8 FILLER_41_88 ();
 sg13g2_decap_8 FILLER_41_95 ();
 sg13g2_decap_4 FILLER_41_106 ();
 sg13g2_fill_1 FILLER_41_110 ();
 sg13g2_decap_8 FILLER_41_116 ();
 sg13g2_decap_8 FILLER_41_123 ();
 sg13g2_fill_2 FILLER_41_130 ();
 sg13g2_decap_8 FILLER_41_144 ();
 sg13g2_fill_1 FILLER_41_178 ();
 sg13g2_fill_1 FILLER_41_193 ();
 sg13g2_decap_8 FILLER_41_198 ();
 sg13g2_fill_1 FILLER_41_205 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_fill_1 FILLER_41_217 ();
 sg13g2_fill_2 FILLER_41_236 ();
 sg13g2_decap_4 FILLER_41_243 ();
 sg13g2_decap_4 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_260 ();
 sg13g2_decap_4 FILLER_41_267 ();
 sg13g2_fill_2 FILLER_41_280 ();
 sg13g2_fill_1 FILLER_41_282 ();
 sg13g2_fill_2 FILLER_41_287 ();
 sg13g2_fill_1 FILLER_41_298 ();
 sg13g2_fill_2 FILLER_41_315 ();
 sg13g2_fill_1 FILLER_41_317 ();
 sg13g2_decap_8 FILLER_41_323 ();
 sg13g2_decap_8 FILLER_41_334 ();
 sg13g2_fill_2 FILLER_41_341 ();
 sg13g2_fill_2 FILLER_41_348 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_382 ();
 sg13g2_decap_4 FILLER_41_389 ();
 sg13g2_fill_1 FILLER_41_402 ();
 sg13g2_decap_4 FILLER_41_423 ();
 sg13g2_fill_2 FILLER_41_427 ();
 sg13g2_decap_4 FILLER_41_433 ();
 sg13g2_fill_2 FILLER_41_437 ();
 sg13g2_fill_2 FILLER_41_445 ();
 sg13g2_fill_1 FILLER_41_473 ();
 sg13g2_fill_2 FILLER_41_513 ();
 sg13g2_fill_2 FILLER_41_524 ();
 sg13g2_fill_1 FILLER_41_534 ();
 sg13g2_fill_2 FILLER_41_547 ();
 sg13g2_fill_1 FILLER_41_549 ();
 sg13g2_decap_4 FILLER_41_562 ();
 sg13g2_fill_2 FILLER_41_566 ();
 sg13g2_fill_2 FILLER_41_589 ();
 sg13g2_fill_1 FILLER_41_595 ();
 sg13g2_fill_2 FILLER_41_607 ();
 sg13g2_decap_8 FILLER_41_613 ();
 sg13g2_decap_4 FILLER_41_620 ();
 sg13g2_fill_2 FILLER_41_624 ();
 sg13g2_fill_2 FILLER_41_634 ();
 sg13g2_fill_1 FILLER_41_636 ();
 sg13g2_fill_2 FILLER_41_679 ();
 sg13g2_fill_1 FILLER_41_681 ();
 sg13g2_fill_1 FILLER_41_694 ();
 sg13g2_decap_4 FILLER_41_700 ();
 sg13g2_decap_4 FILLER_41_712 ();
 sg13g2_fill_1 FILLER_41_716 ();
 sg13g2_decap_4 FILLER_41_722 ();
 sg13g2_fill_1 FILLER_41_726 ();
 sg13g2_decap_8 FILLER_41_732 ();
 sg13g2_decap_4 FILLER_41_739 ();
 sg13g2_fill_1 FILLER_41_743 ();
 sg13g2_fill_1 FILLER_41_748 ();
 sg13g2_fill_1 FILLER_41_754 ();
 sg13g2_fill_2 FILLER_41_760 ();
 sg13g2_fill_1 FILLER_41_762 ();
 sg13g2_fill_1 FILLER_41_767 ();
 sg13g2_fill_2 FILLER_41_773 ();
 sg13g2_fill_1 FILLER_41_810 ();
 sg13g2_fill_2 FILLER_41_823 ();
 sg13g2_fill_1 FILLER_41_833 ();
 sg13g2_fill_2 FILLER_41_838 ();
 sg13g2_fill_2 FILLER_41_848 ();
 sg13g2_fill_1 FILLER_41_854 ();
 sg13g2_fill_2 FILLER_41_858 ();
 sg13g2_fill_1 FILLER_41_860 ();
 sg13g2_decap_4 FILLER_41_865 ();
 sg13g2_fill_1 FILLER_41_895 ();
 sg13g2_decap_8 FILLER_41_909 ();
 sg13g2_fill_1 FILLER_41_916 ();
 sg13g2_decap_4 FILLER_41_952 ();
 sg13g2_fill_2 FILLER_41_956 ();
 sg13g2_decap_8 FILLER_41_966 ();
 sg13g2_decap_4 FILLER_41_973 ();
 sg13g2_fill_1 FILLER_41_977 ();
 sg13g2_fill_1 FILLER_41_996 ();
 sg13g2_decap_4 FILLER_41_1032 ();
 sg13g2_decap_8 FILLER_41_1040 ();
 sg13g2_fill_1 FILLER_41_1059 ();
 sg13g2_fill_1 FILLER_41_1096 ();
 sg13g2_decap_4 FILLER_41_1105 ();
 sg13g2_decap_8 FILLER_41_1113 ();
 sg13g2_decap_8 FILLER_41_1120 ();
 sg13g2_fill_2 FILLER_41_1127 ();
 sg13g2_fill_2 FILLER_41_1147 ();
 sg13g2_decap_4 FILLER_41_1152 ();
 sg13g2_fill_1 FILLER_41_1175 ();
 sg13g2_decap_8 FILLER_41_1181 ();
 sg13g2_decap_4 FILLER_41_1188 ();
 sg13g2_fill_2 FILLER_41_1192 ();
 sg13g2_fill_2 FILLER_41_1225 ();
 sg13g2_fill_1 FILLER_41_1227 ();
 sg13g2_decap_4 FILLER_41_1232 ();
 sg13g2_fill_1 FILLER_41_1236 ();
 sg13g2_fill_2 FILLER_41_1242 ();
 sg13g2_decap_4 FILLER_41_1248 ();
 sg13g2_fill_2 FILLER_41_1252 ();
 sg13g2_decap_4 FILLER_41_1268 ();
 sg13g2_decap_8 FILLER_41_1276 ();
 sg13g2_fill_2 FILLER_41_1283 ();
 sg13g2_decap_4 FILLER_41_1295 ();
 sg13g2_fill_1 FILLER_41_1299 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_11 ();
 sg13g2_decap_4 FILLER_42_18 ();
 sg13g2_fill_1 FILLER_42_22 ();
 sg13g2_decap_4 FILLER_42_34 ();
 sg13g2_fill_1 FILLER_42_38 ();
 sg13g2_decap_4 FILLER_42_74 ();
 sg13g2_fill_2 FILLER_42_91 ();
 sg13g2_decap_4 FILLER_42_123 ();
 sg13g2_fill_1 FILLER_42_135 ();
 sg13g2_fill_2 FILLER_42_144 ();
 sg13g2_fill_1 FILLER_42_146 ();
 sg13g2_decap_8 FILLER_42_151 ();
 sg13g2_decap_8 FILLER_42_158 ();
 sg13g2_decap_8 FILLER_42_165 ();
 sg13g2_fill_1 FILLER_42_172 ();
 sg13g2_decap_8 FILLER_42_185 ();
 sg13g2_fill_2 FILLER_42_192 ();
 sg13g2_fill_2 FILLER_42_251 ();
 sg13g2_fill_1 FILLER_42_258 ();
 sg13g2_fill_1 FILLER_42_308 ();
 sg13g2_fill_1 FILLER_42_316 ();
 sg13g2_fill_2 FILLER_42_321 ();
 sg13g2_fill_1 FILLER_42_328 ();
 sg13g2_fill_2 FILLER_42_355 ();
 sg13g2_fill_2 FILLER_42_360 ();
 sg13g2_fill_1 FILLER_42_362 ();
 sg13g2_decap_8 FILLER_42_367 ();
 sg13g2_decap_8 FILLER_42_374 ();
 sg13g2_fill_2 FILLER_42_381 ();
 sg13g2_fill_1 FILLER_42_383 ();
 sg13g2_fill_2 FILLER_42_414 ();
 sg13g2_fill_2 FILLER_42_426 ();
 sg13g2_decap_4 FILLER_42_432 ();
 sg13g2_fill_1 FILLER_42_436 ();
 sg13g2_decap_8 FILLER_42_443 ();
 sg13g2_fill_2 FILLER_42_450 ();
 sg13g2_decap_8 FILLER_42_456 ();
 sg13g2_fill_1 FILLER_42_463 ();
 sg13g2_decap_4 FILLER_42_502 ();
 sg13g2_fill_1 FILLER_42_506 ();
 sg13g2_decap_8 FILLER_42_510 ();
 sg13g2_decap_8 FILLER_42_517 ();
 sg13g2_fill_2 FILLER_42_524 ();
 sg13g2_decap_4 FILLER_42_530 ();
 sg13g2_decap_8 FILLER_42_538 ();
 sg13g2_decap_4 FILLER_42_545 ();
 sg13g2_fill_2 FILLER_42_549 ();
 sg13g2_fill_1 FILLER_42_567 ();
 sg13g2_fill_2 FILLER_42_579 ();
 sg13g2_fill_1 FILLER_42_581 ();
 sg13g2_fill_1 FILLER_42_586 ();
 sg13g2_fill_2 FILLER_42_592 ();
 sg13g2_decap_8 FILLER_42_603 ();
 sg13g2_decap_8 FILLER_42_610 ();
 sg13g2_decap_4 FILLER_42_617 ();
 sg13g2_decap_8 FILLER_42_639 ();
 sg13g2_decap_4 FILLER_42_646 ();
 sg13g2_decap_4 FILLER_42_655 ();
 sg13g2_fill_1 FILLER_42_659 ();
 sg13g2_fill_2 FILLER_42_665 ();
 sg13g2_fill_1 FILLER_42_667 ();
 sg13g2_fill_1 FILLER_42_676 ();
 sg13g2_decap_8 FILLER_42_686 ();
 sg13g2_fill_2 FILLER_42_693 ();
 sg13g2_fill_1 FILLER_42_695 ();
 sg13g2_fill_2 FILLER_42_699 ();
 sg13g2_decap_8 FILLER_42_779 ();
 sg13g2_fill_2 FILLER_42_786 ();
 sg13g2_decap_4 FILLER_42_792 ();
 sg13g2_fill_2 FILLER_42_796 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_4 FILLER_42_825 ();
 sg13g2_decap_4 FILLER_42_837 ();
 sg13g2_fill_2 FILLER_42_841 ();
 sg13g2_decap_4 FILLER_42_874 ();
 sg13g2_decap_4 FILLER_42_882 ();
 sg13g2_fill_1 FILLER_42_925 ();
 sg13g2_decap_8 FILLER_42_933 ();
 sg13g2_fill_1 FILLER_42_980 ();
 sg13g2_decap_8 FILLER_42_1007 ();
 sg13g2_fill_2 FILLER_42_1014 ();
 sg13g2_fill_1 FILLER_42_1016 ();
 sg13g2_decap_8 FILLER_42_1029 ();
 sg13g2_fill_1 FILLER_42_1036 ();
 sg13g2_decap_4 FILLER_42_1049 ();
 sg13g2_fill_2 FILLER_42_1053 ();
 sg13g2_decap_4 FILLER_42_1064 ();
 sg13g2_decap_8 FILLER_42_1072 ();
 sg13g2_decap_4 FILLER_42_1079 ();
 sg13g2_fill_1 FILLER_42_1083 ();
 sg13g2_fill_2 FILLER_42_1089 ();
 sg13g2_decap_4 FILLER_42_1095 ();
 sg13g2_decap_8 FILLER_42_1104 ();
 sg13g2_fill_2 FILLER_42_1111 ();
 sg13g2_fill_2 FILLER_42_1121 ();
 sg13g2_fill_1 FILLER_42_1123 ();
 sg13g2_fill_2 FILLER_42_1132 ();
 sg13g2_fill_2 FILLER_42_1139 ();
 sg13g2_fill_1 FILLER_42_1141 ();
 sg13g2_fill_2 FILLER_42_1147 ();
 sg13g2_fill_1 FILLER_42_1149 ();
 sg13g2_fill_1 FILLER_42_1159 ();
 sg13g2_fill_2 FILLER_42_1165 ();
 sg13g2_decap_8 FILLER_42_1179 ();
 sg13g2_decap_8 FILLER_42_1186 ();
 sg13g2_decap_8 FILLER_42_1193 ();
 sg13g2_decap_8 FILLER_42_1209 ();
 sg13g2_fill_2 FILLER_42_1216 ();
 sg13g2_decap_8 FILLER_42_1223 ();
 sg13g2_decap_4 FILLER_42_1230 ();
 sg13g2_fill_2 FILLER_42_1234 ();
 sg13g2_fill_2 FILLER_42_1262 ();
 sg13g2_decap_4 FILLER_42_1290 ();
 sg13g2_fill_1 FILLER_42_1294 ();
 sg13g2_decap_4 FILLER_42_1321 ();
 sg13g2_fill_1 FILLER_42_1325 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_32 ();
 sg13g2_fill_1 FILLER_43_34 ();
 sg13g2_decap_4 FILLER_43_47 ();
 sg13g2_fill_2 FILLER_43_60 ();
 sg13g2_fill_1 FILLER_43_62 ();
 sg13g2_decap_4 FILLER_43_67 ();
 sg13g2_decap_8 FILLER_43_74 ();
 sg13g2_fill_1 FILLER_43_81 ();
 sg13g2_decap_8 FILLER_43_87 ();
 sg13g2_decap_4 FILLER_43_94 ();
 sg13g2_fill_2 FILLER_43_98 ();
 sg13g2_decap_4 FILLER_43_104 ();
 sg13g2_fill_1 FILLER_43_108 ();
 sg13g2_decap_8 FILLER_43_166 ();
 sg13g2_fill_2 FILLER_43_173 ();
 sg13g2_fill_1 FILLER_43_175 ();
 sg13g2_fill_1 FILLER_43_181 ();
 sg13g2_fill_2 FILLER_43_190 ();
 sg13g2_fill_1 FILLER_43_192 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_4 FILLER_43_206 ();
 sg13g2_fill_1 FILLER_43_210 ();
 sg13g2_fill_2 FILLER_43_215 ();
 sg13g2_fill_1 FILLER_43_217 ();
 sg13g2_fill_1 FILLER_43_222 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_fill_1 FILLER_43_239 ();
 sg13g2_fill_2 FILLER_43_244 ();
 sg13g2_fill_1 FILLER_43_254 ();
 sg13g2_fill_2 FILLER_43_262 ();
 sg13g2_fill_2 FILLER_43_268 ();
 sg13g2_decap_8 FILLER_43_274 ();
 sg13g2_decap_8 FILLER_43_281 ();
 sg13g2_fill_2 FILLER_43_288 ();
 sg13g2_fill_1 FILLER_43_290 ();
 sg13g2_decap_4 FILLER_43_298 ();
 sg13g2_fill_2 FILLER_43_302 ();
 sg13g2_fill_1 FILLER_43_324 ();
 sg13g2_fill_1 FILLER_43_329 ();
 sg13g2_fill_1 FILLER_43_334 ();
 sg13g2_decap_8 FILLER_43_339 ();
 sg13g2_fill_2 FILLER_43_346 ();
 sg13g2_fill_1 FILLER_43_348 ();
 sg13g2_decap_4 FILLER_43_358 ();
 sg13g2_decap_8 FILLER_43_379 ();
 sg13g2_decap_8 FILLER_43_386 ();
 sg13g2_fill_1 FILLER_43_393 ();
 sg13g2_fill_2 FILLER_43_399 ();
 sg13g2_fill_1 FILLER_43_401 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_fill_2 FILLER_43_420 ();
 sg13g2_fill_1 FILLER_43_422 ();
 sg13g2_fill_2 FILLER_43_471 ();
 sg13g2_fill_1 FILLER_43_473 ();
 sg13g2_decap_8 FILLER_43_478 ();
 sg13g2_decap_8 FILLER_43_485 ();
 sg13g2_decap_4 FILLER_43_492 ();
 sg13g2_fill_2 FILLER_43_549 ();
 sg13g2_fill_1 FILLER_43_580 ();
 sg13g2_fill_2 FILLER_43_593 ();
 sg13g2_decap_4 FILLER_43_616 ();
 sg13g2_fill_1 FILLER_43_620 ();
 sg13g2_decap_8 FILLER_43_633 ();
 sg13g2_fill_2 FILLER_43_640 ();
 sg13g2_fill_2 FILLER_43_672 ();
 sg13g2_decap_8 FILLER_43_700 ();
 sg13g2_fill_2 FILLER_43_707 ();
 sg13g2_fill_1 FILLER_43_709 ();
 sg13g2_fill_2 FILLER_43_719 ();
 sg13g2_fill_2 FILLER_43_724 ();
 sg13g2_fill_2 FILLER_43_731 ();
 sg13g2_fill_1 FILLER_43_733 ();
 sg13g2_decap_8 FILLER_43_738 ();
 sg13g2_fill_1 FILLER_43_749 ();
 sg13g2_fill_1 FILLER_43_754 ();
 sg13g2_fill_1 FILLER_43_760 ();
 sg13g2_decap_4 FILLER_43_766 ();
 sg13g2_fill_1 FILLER_43_770 ();
 sg13g2_fill_2 FILLER_43_780 ();
 sg13g2_decap_4 FILLER_43_786 ();
 sg13g2_fill_1 FILLER_43_798 ();
 sg13g2_fill_1 FILLER_43_809 ();
 sg13g2_fill_2 FILLER_43_843 ();
 sg13g2_decap_8 FILLER_43_855 ();
 sg13g2_fill_1 FILLER_43_862 ();
 sg13g2_fill_2 FILLER_43_868 ();
 sg13g2_fill_1 FILLER_43_870 ();
 sg13g2_fill_1 FILLER_43_900 ();
 sg13g2_decap_8 FILLER_43_905 ();
 sg13g2_decap_4 FILLER_43_912 ();
 sg13g2_fill_1 FILLER_43_916 ();
 sg13g2_decap_4 FILLER_43_921 ();
 sg13g2_decap_8 FILLER_43_955 ();
 sg13g2_decap_8 FILLER_43_962 ();
 sg13g2_decap_4 FILLER_43_969 ();
 sg13g2_decap_4 FILLER_43_980 ();
 sg13g2_fill_2 FILLER_43_984 ();
 sg13g2_fill_1 FILLER_43_993 ();
 sg13g2_fill_2 FILLER_43_997 ();
 sg13g2_decap_8 FILLER_43_1013 ();
 sg13g2_fill_2 FILLER_43_1020 ();
 sg13g2_fill_1 FILLER_43_1022 ();
 sg13g2_fill_1 FILLER_43_1026 ();
 sg13g2_fill_1 FILLER_43_1033 ();
 sg13g2_fill_1 FILLER_43_1038 ();
 sg13g2_fill_2 FILLER_43_1042 ();
 sg13g2_fill_2 FILLER_43_1051 ();
 sg13g2_fill_1 FILLER_43_1053 ();
 sg13g2_decap_4 FILLER_43_1062 ();
 sg13g2_decap_4 FILLER_43_1069 ();
 sg13g2_fill_1 FILLER_43_1073 ();
 sg13g2_fill_2 FILLER_43_1083 ();
 sg13g2_fill_1 FILLER_43_1085 ();
 sg13g2_decap_8 FILLER_43_1147 ();
 sg13g2_fill_1 FILLER_43_1154 ();
 sg13g2_decap_4 FILLER_43_1159 ();
 sg13g2_fill_2 FILLER_43_1163 ();
 sg13g2_fill_1 FILLER_43_1168 ();
 sg13g2_decap_4 FILLER_43_1174 ();
 sg13g2_decap_4 FILLER_43_1242 ();
 sg13g2_fill_1 FILLER_43_1246 ();
 sg13g2_fill_2 FILLER_43_1252 ();
 sg13g2_fill_1 FILLER_43_1254 ();
 sg13g2_decap_8 FILLER_43_1260 ();
 sg13g2_fill_2 FILLER_43_1267 ();
 sg13g2_decap_8 FILLER_43_1282 ();
 sg13g2_fill_1 FILLER_43_1289 ();
 sg13g2_fill_2 FILLER_43_1304 ();
 sg13g2_fill_1 FILLER_43_1306 ();
 sg13g2_decap_8 FILLER_43_1311 ();
 sg13g2_decap_8 FILLER_43_1318 ();
 sg13g2_fill_1 FILLER_43_1325 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_11 ();
 sg13g2_fill_2 FILLER_44_18 ();
 sg13g2_fill_1 FILLER_44_25 ();
 sg13g2_decap_4 FILLER_44_34 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_75 ();
 sg13g2_fill_1 FILLER_44_85 ();
 sg13g2_decap_8 FILLER_44_100 ();
 sg13g2_fill_1 FILLER_44_107 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_fill_2 FILLER_44_119 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_decap_4 FILLER_44_126 ();
 sg13g2_fill_2 FILLER_44_130 ();
 sg13g2_decap_4 FILLER_44_136 ();
 sg13g2_fill_2 FILLER_44_143 ();
 sg13g2_fill_2 FILLER_44_201 ();
 sg13g2_fill_1 FILLER_44_203 ();
 sg13g2_fill_2 FILLER_44_287 ();
 sg13g2_fill_1 FILLER_44_289 ();
 sg13g2_decap_4 FILLER_44_300 ();
 sg13g2_fill_1 FILLER_44_304 ();
 sg13g2_decap_8 FILLER_44_309 ();
 sg13g2_decap_8 FILLER_44_316 ();
 sg13g2_decap_8 FILLER_44_327 ();
 sg13g2_fill_1 FILLER_44_334 ();
 sg13g2_fill_2 FILLER_44_338 ();
 sg13g2_fill_1 FILLER_44_349 ();
 sg13g2_fill_2 FILLER_44_355 ();
 sg13g2_decap_8 FILLER_44_388 ();
 sg13g2_decap_4 FILLER_44_425 ();
 sg13g2_decap_8 FILLER_44_433 ();
 sg13g2_fill_1 FILLER_44_440 ();
 sg13g2_fill_2 FILLER_44_445 ();
 sg13g2_fill_1 FILLER_44_447 ();
 sg13g2_decap_8 FILLER_44_452 ();
 sg13g2_decap_4 FILLER_44_459 ();
 sg13g2_fill_2 FILLER_44_463 ();
 sg13g2_fill_2 FILLER_44_473 ();
 sg13g2_fill_1 FILLER_44_475 ();
 sg13g2_decap_8 FILLER_44_492 ();
 sg13g2_decap_4 FILLER_44_499 ();
 sg13g2_fill_1 FILLER_44_515 ();
 sg13g2_fill_2 FILLER_44_520 ();
 sg13g2_fill_2 FILLER_44_527 ();
 sg13g2_decap_8 FILLER_44_536 ();
 sg13g2_decap_8 FILLER_44_543 ();
 sg13g2_decap_4 FILLER_44_550 ();
 sg13g2_fill_1 FILLER_44_554 ();
 sg13g2_fill_2 FILLER_44_563 ();
 sg13g2_fill_2 FILLER_44_573 ();
 sg13g2_fill_1 FILLER_44_578 ();
 sg13g2_fill_1 FILLER_44_586 ();
 sg13g2_decap_4 FILLER_44_591 ();
 sg13g2_fill_2 FILLER_44_595 ();
 sg13g2_fill_2 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_643 ();
 sg13g2_fill_2 FILLER_44_650 ();
 sg13g2_fill_1 FILLER_44_652 ();
 sg13g2_decap_4 FILLER_44_662 ();
 sg13g2_fill_2 FILLER_44_666 ();
 sg13g2_decap_4 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_688 ();
 sg13g2_decap_8 FILLER_44_704 ();
 sg13g2_fill_2 FILLER_44_724 ();
 sg13g2_fill_1 FILLER_44_726 ();
 sg13g2_fill_2 FILLER_44_737 ();
 sg13g2_fill_2 FILLER_44_798 ();
 sg13g2_fill_1 FILLER_44_800 ();
 sg13g2_decap_8 FILLER_44_827 ();
 sg13g2_fill_2 FILLER_44_890 ();
 sg13g2_decap_8 FILLER_44_936 ();
 sg13g2_fill_2 FILLER_44_943 ();
 sg13g2_fill_1 FILLER_44_945 ();
 sg13g2_fill_2 FILLER_44_950 ();
 sg13g2_decap_4 FILLER_44_963 ();
 sg13g2_fill_1 FILLER_44_967 ();
 sg13g2_fill_1 FILLER_44_976 ();
 sg13g2_decap_8 FILLER_44_981 ();
 sg13g2_fill_1 FILLER_44_988 ();
 sg13g2_fill_1 FILLER_44_1005 ();
 sg13g2_fill_1 FILLER_44_1010 ();
 sg13g2_decap_4 FILLER_44_1016 ();
 sg13g2_fill_1 FILLER_44_1020 ();
 sg13g2_fill_2 FILLER_44_1029 ();
 sg13g2_fill_1 FILLER_44_1031 ();
 sg13g2_fill_1 FILLER_44_1036 ();
 sg13g2_fill_2 FILLER_44_1065 ();
 sg13g2_fill_1 FILLER_44_1084 ();
 sg13g2_decap_8 FILLER_44_1093 ();
 sg13g2_decap_8 FILLER_44_1104 ();
 sg13g2_decap_4 FILLER_44_1111 ();
 sg13g2_fill_1 FILLER_44_1115 ();
 sg13g2_decap_4 FILLER_44_1121 ();
 sg13g2_fill_2 FILLER_44_1130 ();
 sg13g2_fill_1 FILLER_44_1132 ();
 sg13g2_fill_1 FILLER_44_1147 ();
 sg13g2_decap_8 FILLER_44_1160 ();
 sg13g2_fill_1 FILLER_44_1175 ();
 sg13g2_fill_2 FILLER_44_1180 ();
 sg13g2_fill_1 FILLER_44_1182 ();
 sg13g2_fill_1 FILLER_44_1222 ();
 sg13g2_decap_8 FILLER_44_1227 ();
 sg13g2_fill_2 FILLER_44_1282 ();
 sg13g2_decap_8 FILLER_44_1310 ();
 sg13g2_decap_8 FILLER_44_1317 ();
 sg13g2_fill_2 FILLER_44_1324 ();
 sg13g2_fill_1 FILLER_45_35 ();
 sg13g2_fill_1 FILLER_45_41 ();
 sg13g2_fill_1 FILLER_45_45 ();
 sg13g2_fill_1 FILLER_45_50 ();
 sg13g2_fill_2 FILLER_45_55 ();
 sg13g2_fill_2 FILLER_45_61 ();
 sg13g2_fill_2 FILLER_45_66 ();
 sg13g2_fill_1 FILLER_45_97 ();
 sg13g2_fill_2 FILLER_45_102 ();
 sg13g2_fill_1 FILLER_45_104 ();
 sg13g2_fill_2 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_165 ();
 sg13g2_decap_4 FILLER_45_169 ();
 sg13g2_decap_8 FILLER_45_176 ();
 sg13g2_decap_8 FILLER_45_183 ();
 sg13g2_fill_2 FILLER_45_190 ();
 sg13g2_decap_4 FILLER_45_196 ();
 sg13g2_fill_2 FILLER_45_213 ();
 sg13g2_fill_2 FILLER_45_220 ();
 sg13g2_fill_1 FILLER_45_222 ();
 sg13g2_fill_1 FILLER_45_232 ();
 sg13g2_decap_8 FILLER_45_242 ();
 sg13g2_decap_4 FILLER_45_261 ();
 sg13g2_fill_2 FILLER_45_265 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_decap_4 FILLER_45_278 ();
 sg13g2_fill_2 FILLER_45_295 ();
 sg13g2_decap_8 FILLER_45_300 ();
 sg13g2_decap_4 FILLER_45_307 ();
 sg13g2_fill_1 FILLER_45_321 ();
 sg13g2_fill_2 FILLER_45_330 ();
 sg13g2_fill_1 FILLER_45_332 ();
 sg13g2_fill_2 FILLER_45_348 ();
 sg13g2_fill_1 FILLER_45_350 ();
 sg13g2_fill_2 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_fill_2 FILLER_45_375 ();
 sg13g2_decap_4 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_415 ();
 sg13g2_decap_4 FILLER_45_452 ();
 sg13g2_decap_8 FILLER_45_464 ();
 sg13g2_fill_1 FILLER_45_471 ();
 sg13g2_decap_4 FILLER_45_496 ();
 sg13g2_fill_2 FILLER_45_500 ();
 sg13g2_fill_1 FILLER_45_509 ();
 sg13g2_fill_1 FILLER_45_513 ();
 sg13g2_fill_1 FILLER_45_518 ();
 sg13g2_decap_8 FILLER_45_531 ();
 sg13g2_fill_2 FILLER_45_538 ();
 sg13g2_fill_1 FILLER_45_560 ();
 sg13g2_fill_1 FILLER_45_568 ();
 sg13g2_fill_1 FILLER_45_573 ();
 sg13g2_fill_1 FILLER_45_579 ();
 sg13g2_fill_1 FILLER_45_586 ();
 sg13g2_decap_4 FILLER_45_592 ();
 sg13g2_fill_1 FILLER_45_596 ();
 sg13g2_decap_4 FILLER_45_618 ();
 sg13g2_fill_2 FILLER_45_622 ();
 sg13g2_fill_1 FILLER_45_633 ();
 sg13g2_decap_8 FILLER_45_643 ();
 sg13g2_fill_1 FILLER_45_689 ();
 sg13g2_decap_8 FILLER_45_698 ();
 sg13g2_fill_2 FILLER_45_705 ();
 sg13g2_fill_1 FILLER_45_717 ();
 sg13g2_fill_2 FILLER_45_723 ();
 sg13g2_fill_2 FILLER_45_729 ();
 sg13g2_fill_1 FILLER_45_731 ();
 sg13g2_decap_4 FILLER_45_740 ();
 sg13g2_fill_1 FILLER_45_744 ();
 sg13g2_fill_1 FILLER_45_748 ();
 sg13g2_fill_2 FILLER_45_753 ();
 sg13g2_fill_1 FILLER_45_755 ();
 sg13g2_fill_2 FILLER_45_768 ();
 sg13g2_decap_4 FILLER_45_773 ();
 sg13g2_fill_1 FILLER_45_777 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_decap_4 FILLER_45_805 ();
 sg13g2_fill_1 FILLER_45_809 ();
 sg13g2_fill_2 FILLER_45_814 ();
 sg13g2_fill_2 FILLER_45_828 ();
 sg13g2_decap_4 FILLER_45_834 ();
 sg13g2_fill_1 FILLER_45_838 ();
 sg13g2_fill_2 FILLER_45_844 ();
 sg13g2_decap_8 FILLER_45_851 ();
 sg13g2_decap_8 FILLER_45_858 ();
 sg13g2_fill_2 FILLER_45_865 ();
 sg13g2_fill_1 FILLER_45_867 ();
 sg13g2_fill_2 FILLER_45_882 ();
 sg13g2_fill_2 FILLER_45_893 ();
 sg13g2_fill_1 FILLER_45_895 ();
 sg13g2_decap_4 FILLER_45_900 ();
 sg13g2_fill_2 FILLER_45_904 ();
 sg13g2_fill_2 FILLER_45_910 ();
 sg13g2_decap_4 FILLER_45_916 ();
 sg13g2_fill_1 FILLER_45_963 ();
 sg13g2_decap_8 FILLER_45_968 ();
 sg13g2_fill_2 FILLER_45_975 ();
 sg13g2_fill_1 FILLER_45_977 ();
 sg13g2_fill_2 FILLER_45_982 ();
 sg13g2_decap_4 FILLER_45_999 ();
 sg13g2_fill_1 FILLER_45_1003 ();
 sg13g2_fill_1 FILLER_45_1025 ();
 sg13g2_decap_8 FILLER_45_1030 ();
 sg13g2_fill_2 FILLER_45_1045 ();
 sg13g2_fill_1 FILLER_45_1057 ();
 sg13g2_fill_2 FILLER_45_1065 ();
 sg13g2_decap_4 FILLER_45_1087 ();
 sg13g2_decap_4 FILLER_45_1108 ();
 sg13g2_fill_1 FILLER_45_1112 ();
 sg13g2_fill_1 FILLER_45_1153 ();
 sg13g2_fill_1 FILLER_45_1199 ();
 sg13g2_fill_1 FILLER_45_1203 ();
 sg13g2_fill_1 FILLER_45_1209 ();
 sg13g2_fill_1 FILLER_45_1218 ();
 sg13g2_fill_1 FILLER_45_1245 ();
 sg13g2_decap_4 FILLER_45_1286 ();
 sg13g2_fill_1 FILLER_45_1290 ();
 sg13g2_decap_8 FILLER_45_1295 ();
 sg13g2_decap_8 FILLER_45_1302 ();
 sg13g2_decap_8 FILLER_45_1309 ();
 sg13g2_decap_8 FILLER_45_1316 ();
 sg13g2_fill_2 FILLER_45_1323 ();
 sg13g2_fill_1 FILLER_45_1325 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_fill_1 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_23 ();
 sg13g2_fill_2 FILLER_46_36 ();
 sg13g2_fill_1 FILLER_46_49 ();
 sg13g2_fill_2 FILLER_46_85 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_decap_8 FILLER_46_97 ();
 sg13g2_decap_8 FILLER_46_104 ();
 sg13g2_decap_4 FILLER_46_111 ();
 sg13g2_fill_2 FILLER_46_133 ();
 sg13g2_fill_1 FILLER_46_145 ();
 sg13g2_fill_2 FILLER_46_154 ();
 sg13g2_fill_2 FILLER_46_208 ();
 sg13g2_decap_8 FILLER_46_225 ();
 sg13g2_decap_4 FILLER_46_232 ();
 sg13g2_decap_4 FILLER_46_266 ();
 sg13g2_fill_1 FILLER_46_270 ();
 sg13g2_fill_2 FILLER_46_275 ();
 sg13g2_fill_1 FILLER_46_277 ();
 sg13g2_decap_8 FILLER_46_286 ();
 sg13g2_decap_4 FILLER_46_293 ();
 sg13g2_fill_1 FILLER_46_297 ();
 sg13g2_fill_1 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_321 ();
 sg13g2_fill_2 FILLER_46_335 ();
 sg13g2_fill_2 FILLER_46_340 ();
 sg13g2_fill_1 FILLER_46_342 ();
 sg13g2_decap_8 FILLER_46_386 ();
 sg13g2_decap_4 FILLER_46_393 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_decap_8 FILLER_46_414 ();
 sg13g2_decap_8 FILLER_46_421 ();
 sg13g2_decap_8 FILLER_46_428 ();
 sg13g2_fill_1 FILLER_46_435 ();
 sg13g2_fill_1 FILLER_46_455 ();
 sg13g2_decap_4 FILLER_46_472 ();
 sg13g2_fill_2 FILLER_46_476 ();
 sg13g2_fill_1 FILLER_46_486 ();
 sg13g2_decap_8 FILLER_46_495 ();
 sg13g2_fill_2 FILLER_46_502 ();
 sg13g2_fill_2 FILLER_46_525 ();
 sg13g2_fill_1 FILLER_46_527 ();
 sg13g2_decap_4 FILLER_46_533 ();
 sg13g2_fill_2 FILLER_46_537 ();
 sg13g2_fill_2 FILLER_46_550 ();
 sg13g2_fill_1 FILLER_46_552 ();
 sg13g2_fill_1 FILLER_46_569 ();
 sg13g2_decap_8 FILLER_46_579 ();
 sg13g2_decap_4 FILLER_46_600 ();
 sg13g2_fill_2 FILLER_46_604 ();
 sg13g2_fill_1 FILLER_46_614 ();
 sg13g2_fill_1 FILLER_46_619 ();
 sg13g2_decap_8 FILLER_46_628 ();
 sg13g2_decap_4 FILLER_46_635 ();
 sg13g2_fill_2 FILLER_46_668 ();
 sg13g2_decap_8 FILLER_46_703 ();
 sg13g2_fill_1 FILLER_46_710 ();
 sg13g2_decap_4 FILLER_46_749 ();
 sg13g2_fill_1 FILLER_46_773 ();
 sg13g2_fill_2 FILLER_46_782 ();
 sg13g2_fill_1 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_797 ();
 sg13g2_decap_8 FILLER_46_804 ();
 sg13g2_fill_2 FILLER_46_811 ();
 sg13g2_fill_1 FILLER_46_817 ();
 sg13g2_fill_1 FILLER_46_913 ();
 sg13g2_fill_2 FILLER_46_919 ();
 sg13g2_fill_1 FILLER_46_921 ();
 sg13g2_fill_1 FILLER_46_929 ();
 sg13g2_decap_8 FILLER_46_937 ();
 sg13g2_decap_8 FILLER_46_944 ();
 sg13g2_decap_8 FILLER_46_951 ();
 sg13g2_decap_8 FILLER_46_958 ();
 sg13g2_fill_2 FILLER_46_965 ();
 sg13g2_decap_8 FILLER_46_970 ();
 sg13g2_decap_8 FILLER_46_977 ();
 sg13g2_fill_1 FILLER_46_992 ();
 sg13g2_fill_2 FILLER_46_1015 ();
 sg13g2_decap_8 FILLER_46_1041 ();
 sg13g2_fill_2 FILLER_46_1048 ();
 sg13g2_fill_1 FILLER_46_1050 ();
 sg13g2_decap_8 FILLER_46_1054 ();
 sg13g2_decap_8 FILLER_46_1061 ();
 sg13g2_decap_4 FILLER_46_1068 ();
 sg13g2_fill_2 FILLER_46_1072 ();
 sg13g2_fill_1 FILLER_46_1088 ();
 sg13g2_fill_2 FILLER_46_1094 ();
 sg13g2_decap_4 FILLER_46_1130 ();
 sg13g2_fill_1 FILLER_46_1134 ();
 sg13g2_decap_8 FILLER_46_1148 ();
 sg13g2_decap_8 FILLER_46_1155 ();
 sg13g2_fill_1 FILLER_46_1170 ();
 sg13g2_fill_1 FILLER_46_1185 ();
 sg13g2_fill_1 FILLER_46_1195 ();
 sg13g2_fill_1 FILLER_46_1200 ();
 sg13g2_decap_8 FILLER_46_1206 ();
 sg13g2_fill_1 FILLER_46_1222 ();
 sg13g2_decap_8 FILLER_46_1231 ();
 sg13g2_decap_8 FILLER_46_1238 ();
 sg13g2_decap_8 FILLER_46_1245 ();
 sg13g2_fill_2 FILLER_46_1252 ();
 sg13g2_decap_8 FILLER_46_1264 ();
 sg13g2_decap_4 FILLER_46_1271 ();
 sg13g2_fill_1 FILLER_46_1275 ();
 sg13g2_decap_8 FILLER_46_1307 ();
 sg13g2_decap_8 FILLER_46_1314 ();
 sg13g2_decap_4 FILLER_46_1321 ();
 sg13g2_fill_1 FILLER_46_1325 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_26 ();
 sg13g2_decap_8 FILLER_47_34 ();
 sg13g2_fill_2 FILLER_47_41 ();
 sg13g2_fill_1 FILLER_47_51 ();
 sg13g2_fill_1 FILLER_47_60 ();
 sg13g2_decap_4 FILLER_47_65 ();
 sg13g2_fill_2 FILLER_47_69 ();
 sg13g2_fill_1 FILLER_47_81 ();
 sg13g2_fill_1 FILLER_47_112 ();
 sg13g2_fill_1 FILLER_47_139 ();
 sg13g2_fill_2 FILLER_47_166 ();
 sg13g2_fill_1 FILLER_47_173 ();
 sg13g2_fill_1 FILLER_47_178 ();
 sg13g2_fill_2 FILLER_47_183 ();
 sg13g2_fill_1 FILLER_47_185 ();
 sg13g2_fill_1 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_209 ();
 sg13g2_fill_1 FILLER_47_214 ();
 sg13g2_fill_2 FILLER_47_226 ();
 sg13g2_decap_4 FILLER_47_232 ();
 sg13g2_decap_8 FILLER_47_253 ();
 sg13g2_decap_8 FILLER_47_260 ();
 sg13g2_fill_1 FILLER_47_267 ();
 sg13g2_decap_4 FILLER_47_289 ();
 sg13g2_fill_1 FILLER_47_293 ();
 sg13g2_fill_1 FILLER_47_305 ();
 sg13g2_fill_1 FILLER_47_326 ();
 sg13g2_fill_2 FILLER_47_342 ();
 sg13g2_fill_1 FILLER_47_344 ();
 sg13g2_fill_1 FILLER_47_431 ();
 sg13g2_fill_1 FILLER_47_440 ();
 sg13g2_fill_1 FILLER_47_449 ();
 sg13g2_decap_4 FILLER_47_454 ();
 sg13g2_fill_1 FILLER_47_458 ();
 sg13g2_fill_1 FILLER_47_463 ();
 sg13g2_fill_1 FILLER_47_468 ();
 sg13g2_fill_1 FILLER_47_473 ();
 sg13g2_fill_1 FILLER_47_486 ();
 sg13g2_decap_8 FILLER_47_492 ();
 sg13g2_decap_8 FILLER_47_499 ();
 sg13g2_fill_1 FILLER_47_510 ();
 sg13g2_fill_1 FILLER_47_515 ();
 sg13g2_fill_1 FILLER_47_524 ();
 sg13g2_fill_1 FILLER_47_534 ();
 sg13g2_decap_4 FILLER_47_540 ();
 sg13g2_fill_2 FILLER_47_544 ();
 sg13g2_fill_2 FILLER_47_551 ();
 sg13g2_fill_1 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_558 ();
 sg13g2_fill_1 FILLER_47_565 ();
 sg13g2_fill_2 FILLER_47_569 ();
 sg13g2_fill_1 FILLER_47_571 ();
 sg13g2_decap_8 FILLER_47_576 ();
 sg13g2_fill_2 FILLER_47_598 ();
 sg13g2_fill_1 FILLER_47_600 ();
 sg13g2_fill_1 FILLER_47_625 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_fill_1 FILLER_47_644 ();
 sg13g2_fill_1 FILLER_47_663 ();
 sg13g2_fill_1 FILLER_47_680 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_fill_1 FILLER_47_693 ();
 sg13g2_fill_1 FILLER_47_734 ();
 sg13g2_fill_2 FILLER_47_739 ();
 sg13g2_fill_2 FILLER_47_749 ();
 sg13g2_fill_2 FILLER_47_759 ();
 sg13g2_fill_1 FILLER_47_761 ();
 sg13g2_fill_1 FILLER_47_770 ();
 sg13g2_fill_2 FILLER_47_776 ();
 sg13g2_fill_1 FILLER_47_783 ();
 sg13g2_fill_2 FILLER_47_788 ();
 sg13g2_fill_2 FILLER_47_798 ();
 sg13g2_fill_1 FILLER_47_800 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_832 ();
 sg13g2_decap_8 FILLER_47_843 ();
 sg13g2_fill_2 FILLER_47_850 ();
 sg13g2_decap_8 FILLER_47_857 ();
 sg13g2_fill_1 FILLER_47_864 ();
 sg13g2_decap_8 FILLER_47_869 ();
 sg13g2_decap_8 FILLER_47_876 ();
 sg13g2_fill_2 FILLER_47_883 ();
 sg13g2_fill_1 FILLER_47_890 ();
 sg13g2_fill_2 FILLER_47_895 ();
 sg13g2_fill_1 FILLER_47_897 ();
 sg13g2_fill_1 FILLER_47_903 ();
 sg13g2_fill_1 FILLER_47_930 ();
 sg13g2_decap_4 FILLER_47_961 ();
 sg13g2_fill_1 FILLER_47_965 ();
 sg13g2_decap_8 FILLER_47_970 ();
 sg13g2_decap_8 FILLER_47_977 ();
 sg13g2_decap_8 FILLER_47_984 ();
 sg13g2_fill_2 FILLER_47_991 ();
 sg13g2_fill_1 FILLER_47_993 ();
 sg13g2_fill_2 FILLER_47_997 ();
 sg13g2_fill_1 FILLER_47_1008 ();
 sg13g2_fill_2 FILLER_47_1013 ();
 sg13g2_fill_1 FILLER_47_1015 ();
 sg13g2_fill_1 FILLER_47_1030 ();
 sg13g2_fill_1 FILLER_47_1036 ();
 sg13g2_decap_4 FILLER_47_1050 ();
 sg13g2_fill_2 FILLER_47_1054 ();
 sg13g2_fill_2 FILLER_47_1062 ();
 sg13g2_fill_2 FILLER_47_1090 ();
 sg13g2_decap_8 FILLER_47_1108 ();
 sg13g2_decap_4 FILLER_47_1115 ();
 sg13g2_fill_1 FILLER_47_1123 ();
 sg13g2_fill_2 FILLER_47_1150 ();
 sg13g2_fill_1 FILLER_47_1152 ();
 sg13g2_fill_1 FILLER_47_1157 ();
 sg13g2_fill_2 FILLER_47_1162 ();
 sg13g2_fill_2 FILLER_47_1168 ();
 sg13g2_fill_2 FILLER_47_1175 ();
 sg13g2_fill_1 FILLER_47_1177 ();
 sg13g2_fill_1 FILLER_47_1182 ();
 sg13g2_decap_8 FILLER_47_1190 ();
 sg13g2_decap_8 FILLER_47_1202 ();
 sg13g2_decap_4 FILLER_47_1209 ();
 sg13g2_fill_1 FILLER_47_1213 ();
 sg13g2_fill_2 FILLER_47_1221 ();
 sg13g2_decap_8 FILLER_47_1236 ();
 sg13g2_fill_1 FILLER_47_1269 ();
 sg13g2_fill_2 FILLER_47_1275 ();
 sg13g2_fill_1 FILLER_47_1281 ();
 sg13g2_fill_1 FILLER_47_1285 ();
 sg13g2_fill_2 FILLER_47_1290 ();
 sg13g2_decap_8 FILLER_47_1296 ();
 sg13g2_decap_8 FILLER_47_1303 ();
 sg13g2_decap_8 FILLER_47_1310 ();
 sg13g2_decap_8 FILLER_47_1317 ();
 sg13g2_fill_2 FILLER_47_1324 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_32 ();
 sg13g2_fill_1 FILLER_48_36 ();
 sg13g2_fill_2 FILLER_48_45 ();
 sg13g2_fill_1 FILLER_48_47 ();
 sg13g2_decap_8 FILLER_48_67 ();
 sg13g2_decap_4 FILLER_48_74 ();
 sg13g2_fill_2 FILLER_48_82 ();
 sg13g2_fill_1 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_108 ();
 sg13g2_decap_8 FILLER_48_115 ();
 sg13g2_fill_2 FILLER_48_122 ();
 sg13g2_decap_8 FILLER_48_137 ();
 sg13g2_fill_2 FILLER_48_144 ();
 sg13g2_decap_8 FILLER_48_177 ();
 sg13g2_decap_8 FILLER_48_184 ();
 sg13g2_fill_1 FILLER_48_191 ();
 sg13g2_fill_1 FILLER_48_199 ();
 sg13g2_fill_2 FILLER_48_215 ();
 sg13g2_fill_1 FILLER_48_217 ();
 sg13g2_decap_4 FILLER_48_228 ();
 sg13g2_decap_4 FILLER_48_244 ();
 sg13g2_fill_2 FILLER_48_248 ();
 sg13g2_fill_2 FILLER_48_255 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_fill_2 FILLER_48_280 ();
 sg13g2_fill_1 FILLER_48_288 ();
 sg13g2_fill_1 FILLER_48_294 ();
 sg13g2_fill_2 FILLER_48_299 ();
 sg13g2_fill_1 FILLER_48_306 ();
 sg13g2_fill_2 FILLER_48_310 ();
 sg13g2_fill_1 FILLER_48_316 ();
 sg13g2_decap_8 FILLER_48_330 ();
 sg13g2_decap_8 FILLER_48_337 ();
 sg13g2_decap_8 FILLER_48_344 ();
 sg13g2_decap_8 FILLER_48_351 ();
 sg13g2_fill_2 FILLER_48_363 ();
 sg13g2_fill_2 FILLER_48_369 ();
 sg13g2_fill_1 FILLER_48_371 ();
 sg13g2_decap_4 FILLER_48_376 ();
 sg13g2_fill_1 FILLER_48_380 ();
 sg13g2_decap_8 FILLER_48_389 ();
 sg13g2_fill_1 FILLER_48_396 ();
 sg13g2_fill_2 FILLER_48_401 ();
 sg13g2_decap_4 FILLER_48_407 ();
 sg13g2_fill_1 FILLER_48_411 ();
 sg13g2_fill_1 FILLER_48_432 ();
 sg13g2_fill_2 FILLER_48_437 ();
 sg13g2_fill_2 FILLER_48_451 ();
 sg13g2_decap_8 FILLER_48_485 ();
 sg13g2_decap_8 FILLER_48_492 ();
 sg13g2_decap_8 FILLER_48_499 ();
 sg13g2_decap_8 FILLER_48_506 ();
 sg13g2_fill_2 FILLER_48_513 ();
 sg13g2_fill_1 FILLER_48_515 ();
 sg13g2_decap_4 FILLER_48_524 ();
 sg13g2_fill_1 FILLER_48_575 ();
 sg13g2_fill_1 FILLER_48_580 ();
 sg13g2_fill_1 FILLER_48_589 ();
 sg13g2_fill_1 FILLER_48_594 ();
 sg13g2_decap_8 FILLER_48_599 ();
 sg13g2_fill_2 FILLER_48_606 ();
 sg13g2_fill_2 FILLER_48_631 ();
 sg13g2_decap_8 FILLER_48_638 ();
 sg13g2_fill_2 FILLER_48_645 ();
 sg13g2_fill_1 FILLER_48_647 ();
 sg13g2_fill_2 FILLER_48_674 ();
 sg13g2_fill_1 FILLER_48_676 ();
 sg13g2_fill_1 FILLER_48_682 ();
 sg13g2_fill_2 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_739 ();
 sg13g2_decap_4 FILLER_48_746 ();
 sg13g2_fill_2 FILLER_48_750 ();
 sg13g2_decap_4 FILLER_48_760 ();
 sg13g2_fill_2 FILLER_48_770 ();
 sg13g2_fill_1 FILLER_48_772 ();
 sg13g2_fill_1 FILLER_48_823 ();
 sg13g2_fill_2 FILLER_48_842 ();
 sg13g2_fill_1 FILLER_48_844 ();
 sg13g2_fill_1 FILLER_48_876 ();
 sg13g2_decap_4 FILLER_48_908 ();
 sg13g2_decap_4 FILLER_48_938 ();
 sg13g2_decap_8 FILLER_48_946 ();
 sg13g2_decap_4 FILLER_48_953 ();
 sg13g2_decap_4 FILLER_48_991 ();
 sg13g2_fill_2 FILLER_48_995 ();
 sg13g2_decap_8 FILLER_48_1005 ();
 sg13g2_fill_1 FILLER_48_1012 ();
 sg13g2_fill_2 FILLER_48_1037 ();
 sg13g2_fill_2 FILLER_48_1056 ();
 sg13g2_decap_4 FILLER_48_1064 ();
 sg13g2_fill_2 FILLER_48_1072 ();
 sg13g2_fill_1 FILLER_48_1074 ();
 sg13g2_decap_4 FILLER_48_1086 ();
 sg13g2_fill_1 FILLER_48_1090 ();
 sg13g2_decap_8 FILLER_48_1131 ();
 sg13g2_decap_8 FILLER_48_1138 ();
 sg13g2_fill_2 FILLER_48_1145 ();
 sg13g2_fill_1 FILLER_48_1155 ();
 sg13g2_fill_2 FILLER_48_1164 ();
 sg13g2_fill_1 FILLER_48_1166 ();
 sg13g2_decap_8 FILLER_48_1172 ();
 sg13g2_fill_2 FILLER_48_1191 ();
 sg13g2_fill_2 FILLER_48_1206 ();
 sg13g2_fill_2 FILLER_48_1213 ();
 sg13g2_fill_1 FILLER_48_1236 ();
 sg13g2_fill_2 FILLER_48_1246 ();
 sg13g2_fill_2 FILLER_48_1252 ();
 sg13g2_decap_8 FILLER_48_1259 ();
 sg13g2_fill_2 FILLER_48_1266 ();
 sg13g2_fill_1 FILLER_48_1285 ();
 sg13g2_decap_8 FILLER_48_1312 ();
 sg13g2_decap_8 FILLER_48_1319 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_7 ();
 sg13g2_fill_2 FILLER_49_21 ();
 sg13g2_fill_1 FILLER_49_33 ();
 sg13g2_fill_2 FILLER_49_39 ();
 sg13g2_fill_2 FILLER_49_54 ();
 sg13g2_decap_8 FILLER_49_64 ();
 sg13g2_decap_4 FILLER_49_71 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_4 FILLER_49_88 ();
 sg13g2_decap_4 FILLER_49_97 ();
 sg13g2_fill_2 FILLER_49_101 ();
 sg13g2_decap_4 FILLER_49_139 ();
 sg13g2_decap_8 FILLER_49_157 ();
 sg13g2_decap_8 FILLER_49_164 ();
 sg13g2_decap_8 FILLER_49_171 ();
 sg13g2_decap_8 FILLER_49_178 ();
 sg13g2_fill_1 FILLER_49_194 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_246 ();
 sg13g2_fill_2 FILLER_49_253 ();
 sg13g2_fill_1 FILLER_49_255 ();
 sg13g2_fill_1 FILLER_49_265 ();
 sg13g2_decap_8 FILLER_49_274 ();
 sg13g2_fill_2 FILLER_49_281 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_331 ();
 sg13g2_decap_8 FILLER_49_340 ();
 sg13g2_fill_2 FILLER_49_363 ();
 sg13g2_fill_2 FILLER_49_391 ();
 sg13g2_fill_1 FILLER_49_393 ();
 sg13g2_fill_2 FILLER_49_428 ();
 sg13g2_fill_1 FILLER_49_438 ();
 sg13g2_fill_2 FILLER_49_447 ();
 sg13g2_fill_1 FILLER_49_458 ();
 sg13g2_fill_2 FILLER_49_476 ();
 sg13g2_fill_1 FILLER_49_482 ();
 sg13g2_decap_8 FILLER_49_493 ();
 sg13g2_decap_8 FILLER_49_500 ();
 sg13g2_decap_4 FILLER_49_511 ();
 sg13g2_fill_2 FILLER_49_522 ();
 sg13g2_fill_1 FILLER_49_528 ();
 sg13g2_decap_8 FILLER_49_533 ();
 sg13g2_fill_2 FILLER_49_540 ();
 sg13g2_fill_1 FILLER_49_542 ();
 sg13g2_decap_4 FILLER_49_551 ();
 sg13g2_fill_2 FILLER_49_555 ();
 sg13g2_fill_1 FILLER_49_561 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_4 FILLER_49_574 ();
 sg13g2_decap_4 FILLER_49_582 ();
 sg13g2_fill_2 FILLER_49_590 ();
 sg13g2_fill_1 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_640 ();
 sg13g2_decap_8 FILLER_49_647 ();
 sg13g2_fill_1 FILLER_49_654 ();
 sg13g2_decap_4 FILLER_49_659 ();
 sg13g2_fill_2 FILLER_49_663 ();
 sg13g2_fill_1 FILLER_49_676 ();
 sg13g2_decap_4 FILLER_49_705 ();
 sg13g2_fill_2 FILLER_49_709 ();
 sg13g2_decap_8 FILLER_49_737 ();
 sg13g2_decap_4 FILLER_49_744 ();
 sg13g2_fill_1 FILLER_49_748 ();
 sg13g2_decap_8 FILLER_49_757 ();
 sg13g2_fill_2 FILLER_49_764 ();
 sg13g2_decap_4 FILLER_49_774 ();
 sg13g2_fill_1 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_789 ();
 sg13g2_decap_8 FILLER_49_796 ();
 sg13g2_fill_1 FILLER_49_803 ();
 sg13g2_fill_1 FILLER_49_821 ();
 sg13g2_fill_2 FILLER_49_834 ();
 sg13g2_fill_1 FILLER_49_836 ();
 sg13g2_decap_4 FILLER_49_841 ();
 sg13g2_fill_1 FILLER_49_845 ();
 sg13g2_decap_4 FILLER_49_893 ();
 sg13g2_fill_1 FILLER_49_905 ();
 sg13g2_fill_1 FILLER_49_915 ();
 sg13g2_decap_8 FILLER_49_923 ();
 sg13g2_decap_4 FILLER_49_930 ();
 sg13g2_fill_2 FILLER_49_934 ();
 sg13g2_fill_2 FILLER_49_940 ();
 sg13g2_fill_1 FILLER_49_942 ();
 sg13g2_decap_8 FILLER_49_947 ();
 sg13g2_decap_4 FILLER_49_954 ();
 sg13g2_fill_2 FILLER_49_958 ();
 sg13g2_fill_2 FILLER_49_963 ();
 sg13g2_decap_8 FILLER_49_1013 ();
 sg13g2_decap_8 FILLER_49_1024 ();
 sg13g2_decap_4 FILLER_49_1031 ();
 sg13g2_decap_4 FILLER_49_1057 ();
 sg13g2_fill_1 FILLER_49_1061 ();
 sg13g2_fill_1 FILLER_49_1066 ();
 sg13g2_decap_4 FILLER_49_1072 ();
 sg13g2_fill_1 FILLER_49_1076 ();
 sg13g2_fill_1 FILLER_49_1102 ();
 sg13g2_fill_1 FILLER_49_1113 ();
 sg13g2_decap_8 FILLER_49_1117 ();
 sg13g2_decap_8 FILLER_49_1124 ();
 sg13g2_decap_4 FILLER_49_1131 ();
 sg13g2_fill_2 FILLER_49_1161 ();
 sg13g2_fill_2 FILLER_49_1166 ();
 sg13g2_decap_4 FILLER_49_1181 ();
 sg13g2_fill_2 FILLER_49_1194 ();
 sg13g2_fill_1 FILLER_49_1196 ();
 sg13g2_fill_2 FILLER_49_1202 ();
 sg13g2_fill_1 FILLER_49_1213 ();
 sg13g2_decap_4 FILLER_49_1260 ();
 sg13g2_fill_1 FILLER_49_1269 ();
 sg13g2_decap_8 FILLER_49_1284 ();
 sg13g2_decap_8 FILLER_49_1291 ();
 sg13g2_decap_8 FILLER_49_1298 ();
 sg13g2_decap_8 FILLER_49_1305 ();
 sg13g2_decap_8 FILLER_49_1312 ();
 sg13g2_decap_8 FILLER_49_1319 ();
 sg13g2_fill_2 FILLER_50_47 ();
 sg13g2_fill_2 FILLER_50_53 ();
 sg13g2_fill_2 FILLER_50_59 ();
 sg13g2_decap_4 FILLER_50_65 ();
 sg13g2_fill_1 FILLER_50_69 ();
 sg13g2_fill_1 FILLER_50_96 ();
 sg13g2_decap_8 FILLER_50_101 ();
 sg13g2_fill_1 FILLER_50_108 ();
 sg13g2_fill_2 FILLER_50_211 ();
 sg13g2_decap_4 FILLER_50_222 ();
 sg13g2_decap_8 FILLER_50_230 ();
 sg13g2_fill_2 FILLER_50_237 ();
 sg13g2_fill_1 FILLER_50_239 ();
 sg13g2_fill_2 FILLER_50_249 ();
 sg13g2_decap_8 FILLER_50_256 ();
 sg13g2_decap_8 FILLER_50_263 ();
 sg13g2_decap_4 FILLER_50_270 ();
 sg13g2_fill_2 FILLER_50_274 ();
 sg13g2_decap_4 FILLER_50_284 ();
 sg13g2_fill_1 FILLER_50_298 ();
 sg13g2_fill_2 FILLER_50_310 ();
 sg13g2_fill_2 FILLER_50_316 ();
 sg13g2_fill_1 FILLER_50_318 ();
 sg13g2_decap_8 FILLER_50_329 ();
 sg13g2_fill_2 FILLER_50_379 ();
 sg13g2_decap_8 FILLER_50_411 ();
 sg13g2_fill_1 FILLER_50_418 ();
 sg13g2_decap_8 FILLER_50_423 ();
 sg13g2_decap_4 FILLER_50_430 ();
 sg13g2_fill_1 FILLER_50_434 ();
 sg13g2_decap_4 FILLER_50_468 ();
 sg13g2_fill_1 FILLER_50_479 ();
 sg13g2_fill_2 FILLER_50_485 ();
 sg13g2_fill_1 FILLER_50_487 ();
 sg13g2_fill_2 FILLER_50_510 ();
 sg13g2_fill_1 FILLER_50_512 ();
 sg13g2_decap_4 FILLER_50_519 ();
 sg13g2_decap_8 FILLER_50_535 ();
 sg13g2_decap_4 FILLER_50_542 ();
 sg13g2_fill_1 FILLER_50_551 ();
 sg13g2_fill_1 FILLER_50_556 ();
 sg13g2_fill_1 FILLER_50_561 ();
 sg13g2_fill_1 FILLER_50_566 ();
 sg13g2_fill_1 FILLER_50_596 ();
 sg13g2_fill_2 FILLER_50_607 ();
 sg13g2_decap_8 FILLER_50_612 ();
 sg13g2_decap_4 FILLER_50_619 ();
 sg13g2_fill_1 FILLER_50_623 ();
 sg13g2_fill_1 FILLER_50_628 ();
 sg13g2_fill_2 FILLER_50_640 ();
 sg13g2_fill_1 FILLER_50_642 ();
 sg13g2_fill_1 FILLER_50_647 ();
 sg13g2_fill_2 FILLER_50_674 ();
 sg13g2_fill_1 FILLER_50_702 ();
 sg13g2_fill_2 FILLER_50_708 ();
 sg13g2_fill_2 FILLER_50_715 ();
 sg13g2_decap_4 FILLER_50_726 ();
 sg13g2_fill_2 FILLER_50_735 ();
 sg13g2_fill_1 FILLER_50_737 ();
 sg13g2_decap_4 FILLER_50_763 ();
 sg13g2_fill_2 FILLER_50_801 ();
 sg13g2_fill_1 FILLER_50_803 ();
 sg13g2_fill_2 FILLER_50_808 ();
 sg13g2_decap_8 FILLER_50_818 ();
 sg13g2_fill_1 FILLER_50_829 ();
 sg13g2_decap_8 FILLER_50_836 ();
 sg13g2_fill_2 FILLER_50_843 ();
 sg13g2_fill_2 FILLER_50_849 ();
 sg13g2_fill_2 FILLER_50_855 ();
 sg13g2_fill_2 FILLER_50_861 ();
 sg13g2_fill_1 FILLER_50_863 ();
 sg13g2_fill_2 FILLER_50_899 ();
 sg13g2_fill_1 FILLER_50_901 ();
 sg13g2_fill_1 FILLER_50_990 ();
 sg13g2_fill_2 FILLER_50_996 ();
 sg13g2_fill_1 FILLER_50_1003 ();
 sg13g2_decap_8 FILLER_50_1034 ();
 sg13g2_decap_8 FILLER_50_1041 ();
 sg13g2_decap_8 FILLER_50_1048 ();
 sg13g2_fill_1 FILLER_50_1055 ();
 sg13g2_decap_4 FILLER_50_1063 ();
 sg13g2_decap_8 FILLER_50_1071 ();
 sg13g2_decap_8 FILLER_50_1078 ();
 sg13g2_decap_4 FILLER_50_1085 ();
 sg13g2_fill_1 FILLER_50_1089 ();
 sg13g2_decap_8 FILLER_50_1103 ();
 sg13g2_fill_2 FILLER_50_1110 ();
 sg13g2_fill_1 FILLER_50_1112 ();
 sg13g2_decap_8 FILLER_50_1134 ();
 sg13g2_fill_2 FILLER_50_1141 ();
 sg13g2_fill_1 FILLER_50_1143 ();
 sg13g2_decap_4 FILLER_50_1148 ();
 sg13g2_fill_1 FILLER_50_1161 ();
 sg13g2_decap_4 FILLER_50_1166 ();
 sg13g2_decap_4 FILLER_50_1178 ();
 sg13g2_decap_4 FILLER_50_1212 ();
 sg13g2_fill_2 FILLER_50_1230 ();
 sg13g2_decap_4 FILLER_50_1258 ();
 sg13g2_fill_1 FILLER_50_1262 ();
 sg13g2_decap_8 FILLER_50_1289 ();
 sg13g2_decap_8 FILLER_50_1296 ();
 sg13g2_decap_8 FILLER_50_1303 ();
 sg13g2_decap_8 FILLER_50_1310 ();
 sg13g2_decap_8 FILLER_50_1317 ();
 sg13g2_fill_2 FILLER_50_1324 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_4 ();
 sg13g2_decap_8 FILLER_51_10 ();
 sg13g2_decap_4 FILLER_51_17 ();
 sg13g2_fill_2 FILLER_51_25 ();
 sg13g2_decap_4 FILLER_51_33 ();
 sg13g2_fill_2 FILLER_51_42 ();
 sg13g2_fill_1 FILLER_51_44 ();
 sg13g2_decap_4 FILLER_51_50 ();
 sg13g2_decap_4 FILLER_51_58 ();
 sg13g2_fill_1 FILLER_51_62 ();
 sg13g2_decap_4 FILLER_51_80 ();
 sg13g2_fill_1 FILLER_51_92 ();
 sg13g2_decap_4 FILLER_51_100 ();
 sg13g2_fill_1 FILLER_51_104 ();
 sg13g2_decap_4 FILLER_51_109 ();
 sg13g2_fill_2 FILLER_51_119 ();
 sg13g2_fill_1 FILLER_51_121 ();
 sg13g2_fill_2 FILLER_51_132 ();
 sg13g2_fill_1 FILLER_51_134 ();
 sg13g2_decap_8 FILLER_51_139 ();
 sg13g2_decap_8 FILLER_51_146 ();
 sg13g2_decap_4 FILLER_51_153 ();
 sg13g2_fill_2 FILLER_51_157 ();
 sg13g2_decap_8 FILLER_51_171 ();
 sg13g2_fill_2 FILLER_51_178 ();
 sg13g2_decap_8 FILLER_51_187 ();
 sg13g2_decap_8 FILLER_51_194 ();
 sg13g2_decap_4 FILLER_51_201 ();
 sg13g2_decap_4 FILLER_51_245 ();
 sg13g2_decap_4 FILLER_51_254 ();
 sg13g2_decap_8 FILLER_51_284 ();
 sg13g2_fill_2 FILLER_51_291 ();
 sg13g2_fill_2 FILLER_51_297 ();
 sg13g2_fill_2 FILLER_51_309 ();
 sg13g2_fill_1 FILLER_51_311 ();
 sg13g2_fill_2 FILLER_51_316 ();
 sg13g2_fill_1 FILLER_51_318 ();
 sg13g2_fill_1 FILLER_51_323 ();
 sg13g2_fill_1 FILLER_51_328 ();
 sg13g2_decap_4 FILLER_51_333 ();
 sg13g2_fill_1 FILLER_51_340 ();
 sg13g2_decap_8 FILLER_51_348 ();
 sg13g2_fill_1 FILLER_51_355 ();
 sg13g2_fill_1 FILLER_51_368 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_decap_4 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_410 ();
 sg13g2_decap_4 FILLER_51_415 ();
 sg13g2_fill_1 FILLER_51_435 ();
 sg13g2_decap_4 FILLER_51_453 ();
 sg13g2_fill_1 FILLER_51_457 ();
 sg13g2_fill_1 FILLER_51_463 ();
 sg13g2_decap_4 FILLER_51_490 ();
 sg13g2_decap_4 FILLER_51_508 ();
 sg13g2_fill_1 FILLER_51_512 ();
 sg13g2_fill_2 FILLER_51_526 ();
 sg13g2_decap_4 FILLER_51_542 ();
 sg13g2_fill_2 FILLER_51_546 ();
 sg13g2_decap_8 FILLER_51_556 ();
 sg13g2_fill_2 FILLER_51_563 ();
 sg13g2_fill_2 FILLER_51_572 ();
 sg13g2_decap_4 FILLER_51_578 ();
 sg13g2_fill_2 FILLER_51_582 ();
 sg13g2_decap_4 FILLER_51_592 ();
 sg13g2_decap_4 FILLER_51_600 ();
 sg13g2_decap_8 FILLER_51_612 ();
 sg13g2_decap_4 FILLER_51_619 ();
 sg13g2_decap_8 FILLER_51_639 ();
 sg13g2_fill_2 FILLER_51_646 ();
 sg13g2_fill_1 FILLER_51_648 ();
 sg13g2_decap_4 FILLER_51_661 ();
 sg13g2_fill_1 FILLER_51_665 ();
 sg13g2_decap_8 FILLER_51_671 ();
 sg13g2_decap_4 FILLER_51_678 ();
 sg13g2_fill_2 FILLER_51_682 ();
 sg13g2_decap_8 FILLER_51_688 ();
 sg13g2_fill_2 FILLER_51_695 ();
 sg13g2_decap_8 FILLER_51_737 ();
 sg13g2_decap_4 FILLER_51_744 ();
 sg13g2_fill_1 FILLER_51_753 ();
 sg13g2_fill_2 FILLER_51_762 ();
 sg13g2_fill_1 FILLER_51_767 ();
 sg13g2_decap_8 FILLER_51_774 ();
 sg13g2_decap_8 FILLER_51_781 ();
 sg13g2_decap_4 FILLER_51_788 ();
 sg13g2_fill_1 FILLER_51_792 ();
 sg13g2_decap_8 FILLER_51_798 ();
 sg13g2_decap_8 FILLER_51_805 ();
 sg13g2_fill_1 FILLER_51_812 ();
 sg13g2_fill_2 FILLER_51_864 ();
 sg13g2_decap_8 FILLER_51_875 ();
 sg13g2_fill_2 FILLER_51_882 ();
 sg13g2_decap_4 FILLER_51_893 ();
 sg13g2_fill_2 FILLER_51_902 ();
 sg13g2_fill_2 FILLER_51_908 ();
 sg13g2_fill_2 FILLER_51_915 ();
 sg13g2_fill_1 FILLER_51_917 ();
 sg13g2_decap_8 FILLER_51_922 ();
 sg13g2_fill_2 FILLER_51_929 ();
 sg13g2_fill_1 FILLER_51_931 ();
 sg13g2_decap_4 FILLER_51_946 ();
 sg13g2_fill_2 FILLER_51_954 ();
 sg13g2_decap_4 FILLER_51_973 ();
 sg13g2_fill_1 FILLER_51_977 ();
 sg13g2_fill_1 FILLER_51_982 ();
 sg13g2_fill_1 FILLER_51_997 ();
 sg13g2_fill_1 FILLER_51_1009 ();
 sg13g2_decap_8 FILLER_51_1017 ();
 sg13g2_fill_2 FILLER_51_1024 ();
 sg13g2_fill_1 FILLER_51_1026 ();
 sg13g2_decap_8 FILLER_51_1035 ();
 sg13g2_fill_2 FILLER_51_1042 ();
 sg13g2_decap_8 FILLER_51_1048 ();
 sg13g2_fill_2 FILLER_51_1055 ();
 sg13g2_fill_1 FILLER_51_1057 ();
 sg13g2_decap_4 FILLER_51_1089 ();
 sg13g2_fill_2 FILLER_51_1119 ();
 sg13g2_fill_1 FILLER_51_1121 ();
 sg13g2_decap_8 FILLER_51_1126 ();
 sg13g2_fill_2 FILLER_51_1133 ();
 sg13g2_fill_1 FILLER_51_1140 ();
 sg13g2_fill_1 FILLER_51_1145 ();
 sg13g2_fill_1 FILLER_51_1152 ();
 sg13g2_fill_1 FILLER_51_1157 ();
 sg13g2_decap_8 FILLER_51_1167 ();
 sg13g2_decap_4 FILLER_51_1174 ();
 sg13g2_fill_1 FILLER_51_1178 ();
 sg13g2_decap_8 FILLER_51_1196 ();
 sg13g2_decap_8 FILLER_51_1203 ();
 sg13g2_fill_2 FILLER_51_1210 ();
 sg13g2_fill_1 FILLER_51_1212 ();
 sg13g2_decap_4 FILLER_51_1223 ();
 sg13g2_fill_1 FILLER_51_1227 ();
 sg13g2_decap_4 FILLER_51_1232 ();
 sg13g2_fill_2 FILLER_51_1236 ();
 sg13g2_decap_4 FILLER_51_1246 ();
 sg13g2_fill_1 FILLER_51_1250 ();
 sg13g2_decap_8 FILLER_51_1255 ();
 sg13g2_decap_8 FILLER_51_1262 ();
 sg13g2_decap_8 FILLER_51_1273 ();
 sg13g2_decap_8 FILLER_51_1280 ();
 sg13g2_decap_8 FILLER_51_1287 ();
 sg13g2_decap_8 FILLER_51_1294 ();
 sg13g2_decap_8 FILLER_51_1301 ();
 sg13g2_decap_8 FILLER_51_1308 ();
 sg13g2_decap_8 FILLER_51_1315 ();
 sg13g2_decap_4 FILLER_51_1322 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_27 ();
 sg13g2_fill_2 FILLER_52_34 ();
 sg13g2_fill_2 FILLER_52_42 ();
 sg13g2_fill_2 FILLER_52_52 ();
 sg13g2_fill_1 FILLER_52_54 ();
 sg13g2_decap_8 FILLER_52_60 ();
 sg13g2_decap_8 FILLER_52_67 ();
 sg13g2_decap_4 FILLER_52_74 ();
 sg13g2_fill_2 FILLER_52_78 ();
 sg13g2_fill_1 FILLER_52_93 ();
 sg13g2_fill_2 FILLER_52_124 ();
 sg13g2_fill_2 FILLER_52_130 ();
 sg13g2_fill_1 FILLER_52_132 ();
 sg13g2_decap_4 FILLER_52_159 ();
 sg13g2_fill_2 FILLER_52_166 ();
 sg13g2_fill_1 FILLER_52_168 ();
 sg13g2_fill_1 FILLER_52_178 ();
 sg13g2_fill_1 FILLER_52_183 ();
 sg13g2_decap_8 FILLER_52_220 ();
 sg13g2_fill_1 FILLER_52_227 ();
 sg13g2_fill_2 FILLER_52_259 ();
 sg13g2_fill_1 FILLER_52_261 ();
 sg13g2_fill_2 FILLER_52_278 ();
 sg13g2_fill_1 FILLER_52_280 ();
 sg13g2_decap_4 FILLER_52_284 ();
 sg13g2_fill_1 FILLER_52_288 ();
 sg13g2_decap_8 FILLER_52_302 ();
 sg13g2_decap_8 FILLER_52_309 ();
 sg13g2_decap_8 FILLER_52_316 ();
 sg13g2_fill_1 FILLER_52_323 ();
 sg13g2_fill_1 FILLER_52_331 ();
 sg13g2_fill_2 FILLER_52_335 ();
 sg13g2_fill_1 FILLER_52_337 ();
 sg13g2_fill_2 FILLER_52_381 ();
 sg13g2_decap_8 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_398 ();
 sg13g2_decap_8 FILLER_52_409 ();
 sg13g2_decap_4 FILLER_52_416 ();
 sg13g2_fill_1 FILLER_52_420 ();
 sg13g2_fill_2 FILLER_52_429 ();
 sg13g2_decap_4 FILLER_52_436 ();
 sg13g2_fill_2 FILLER_52_462 ();
 sg13g2_fill_1 FILLER_52_464 ();
 sg13g2_fill_1 FILLER_52_469 ();
 sg13g2_fill_1 FILLER_52_485 ();
 sg13g2_fill_2 FILLER_52_537 ();
 sg13g2_fill_2 FILLER_52_563 ();
 sg13g2_fill_1 FILLER_52_565 ();
 sg13g2_decap_4 FILLER_52_578 ();
 sg13g2_fill_2 FILLER_52_582 ();
 sg13g2_decap_8 FILLER_52_632 ();
 sg13g2_decap_8 FILLER_52_639 ();
 sg13g2_fill_1 FILLER_52_646 ();
 sg13g2_decap_8 FILLER_52_673 ();
 sg13g2_fill_2 FILLER_52_680 ();
 sg13g2_fill_1 FILLER_52_682 ();
 sg13g2_fill_1 FILLER_52_697 ();
 sg13g2_fill_1 FILLER_52_702 ();
 sg13g2_fill_1 FILLER_52_708 ();
 sg13g2_fill_2 FILLER_52_714 ();
 sg13g2_fill_2 FILLER_52_721 ();
 sg13g2_fill_2 FILLER_52_726 ();
 sg13g2_fill_1 FILLER_52_737 ();
 sg13g2_fill_2 FILLER_52_746 ();
 sg13g2_fill_1 FILLER_52_768 ();
 sg13g2_fill_1 FILLER_52_774 ();
 sg13g2_decap_8 FILLER_52_781 ();
 sg13g2_fill_1 FILLER_52_788 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_fill_2 FILLER_52_819 ();
 sg13g2_fill_2 FILLER_52_825 ();
 sg13g2_decap_8 FILLER_52_849 ();
 sg13g2_fill_1 FILLER_52_856 ();
 sg13g2_decap_8 FILLER_52_863 ();
 sg13g2_fill_1 FILLER_52_870 ();
 sg13g2_fill_1 FILLER_52_875 ();
 sg13g2_fill_2 FILLER_52_905 ();
 sg13g2_fill_1 FILLER_52_907 ();
 sg13g2_fill_2 FILLER_52_985 ();
 sg13g2_fill_1 FILLER_52_987 ();
 sg13g2_fill_1 FILLER_52_997 ();
 sg13g2_fill_1 FILLER_52_1014 ();
 sg13g2_decap_8 FILLER_52_1048 ();
 sg13g2_fill_2 FILLER_52_1055 ();
 sg13g2_fill_1 FILLER_52_1057 ();
 sg13g2_decap_4 FILLER_52_1071 ();
 sg13g2_fill_1 FILLER_52_1075 ();
 sg13g2_fill_2 FILLER_52_1096 ();
 sg13g2_fill_1 FILLER_52_1098 ();
 sg13g2_decap_8 FILLER_52_1103 ();
 sg13g2_decap_4 FILLER_52_1110 ();
 sg13g2_fill_1 FILLER_52_1114 ();
 sg13g2_fill_2 FILLER_52_1145 ();
 sg13g2_fill_1 FILLER_52_1147 ();
 sg13g2_fill_1 FILLER_52_1160 ();
 sg13g2_fill_2 FILLER_52_1165 ();
 sg13g2_fill_2 FILLER_52_1177 ();
 sg13g2_fill_2 FILLER_52_1187 ();
 sg13g2_fill_1 FILLER_52_1189 ();
 sg13g2_decap_8 FILLER_52_1194 ();
 sg13g2_decap_4 FILLER_52_1201 ();
 sg13g2_fill_2 FILLER_52_1205 ();
 sg13g2_decap_4 FILLER_52_1211 ();
 sg13g2_fill_2 FILLER_52_1215 ();
 sg13g2_fill_1 FILLER_52_1227 ();
 sg13g2_fill_2 FILLER_52_1232 ();
 sg13g2_fill_2 FILLER_52_1242 ();
 sg13g2_decap_8 FILLER_52_1274 ();
 sg13g2_decap_8 FILLER_52_1281 ();
 sg13g2_decap_8 FILLER_52_1288 ();
 sg13g2_decap_8 FILLER_52_1295 ();
 sg13g2_decap_8 FILLER_52_1302 ();
 sg13g2_decap_8 FILLER_52_1309 ();
 sg13g2_decap_8 FILLER_52_1316 ();
 sg13g2_fill_2 FILLER_52_1323 ();
 sg13g2_fill_1 FILLER_52_1325 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_8 ();
 sg13g2_fill_1 FILLER_53_10 ();
 sg13g2_fill_1 FILLER_53_15 ();
 sg13g2_fill_2 FILLER_53_35 ();
 sg13g2_fill_1 FILLER_53_37 ();
 sg13g2_fill_1 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_51 ();
 sg13g2_decap_8 FILLER_53_58 ();
 sg13g2_fill_2 FILLER_53_65 ();
 sg13g2_fill_1 FILLER_53_67 ();
 sg13g2_fill_2 FILLER_53_81 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_fill_1 FILLER_53_93 ();
 sg13g2_fill_1 FILLER_53_104 ();
 sg13g2_fill_1 FILLER_53_110 ();
 sg13g2_decap_8 FILLER_53_203 ();
 sg13g2_fill_2 FILLER_53_210 ();
 sg13g2_fill_1 FILLER_53_217 ();
 sg13g2_decap_4 FILLER_53_231 ();
 sg13g2_decap_4 FILLER_53_239 ();
 sg13g2_fill_1 FILLER_53_243 ();
 sg13g2_decap_8 FILLER_53_248 ();
 sg13g2_fill_2 FILLER_53_268 ();
 sg13g2_fill_1 FILLER_53_270 ();
 sg13g2_decap_4 FILLER_53_280 ();
 sg13g2_fill_1 FILLER_53_284 ();
 sg13g2_decap_8 FILLER_53_289 ();
 sg13g2_decap_4 FILLER_53_296 ();
 sg13g2_fill_2 FILLER_53_300 ();
 sg13g2_decap_8 FILLER_53_306 ();
 sg13g2_decap_8 FILLER_53_313 ();
 sg13g2_decap_4 FILLER_53_327 ();
 sg13g2_decap_8 FILLER_53_335 ();
 sg13g2_fill_2 FILLER_53_346 ();
 sg13g2_fill_2 FILLER_53_352 ();
 sg13g2_fill_2 FILLER_53_359 ();
 sg13g2_decap_8 FILLER_53_395 ();
 sg13g2_decap_8 FILLER_53_402 ();
 sg13g2_decap_8 FILLER_53_409 ();
 sg13g2_decap_4 FILLER_53_416 ();
 sg13g2_fill_2 FILLER_53_420 ();
 sg13g2_fill_2 FILLER_53_447 ();
 sg13g2_fill_1 FILLER_53_453 ();
 sg13g2_fill_1 FILLER_53_468 ();
 sg13g2_fill_1 FILLER_53_474 ();
 sg13g2_fill_1 FILLER_53_480 ();
 sg13g2_fill_1 FILLER_53_490 ();
 sg13g2_decap_4 FILLER_53_497 ();
 sg13g2_decap_8 FILLER_53_505 ();
 sg13g2_decap_8 FILLER_53_512 ();
 sg13g2_fill_2 FILLER_53_519 ();
 sg13g2_decap_4 FILLER_53_539 ();
 sg13g2_decap_8 FILLER_53_547 ();
 sg13g2_fill_2 FILLER_53_554 ();
 sg13g2_fill_1 FILLER_53_556 ();
 sg13g2_fill_1 FILLER_53_561 ();
 sg13g2_fill_1 FILLER_53_572 ();
 sg13g2_fill_1 FILLER_53_578 ();
 sg13g2_fill_2 FILLER_53_583 ();
 sg13g2_fill_1 FILLER_53_585 ();
 sg13g2_decap_8 FILLER_53_591 ();
 sg13g2_fill_1 FILLER_53_602 ();
 sg13g2_fill_2 FILLER_53_607 ();
 sg13g2_fill_1 FILLER_53_613 ();
 sg13g2_fill_2 FILLER_53_623 ();
 sg13g2_decap_8 FILLER_53_630 ();
 sg13g2_decap_8 FILLER_53_637 ();
 sg13g2_decap_8 FILLER_53_644 ();
 sg13g2_decap_4 FILLER_53_651 ();
 sg13g2_fill_1 FILLER_53_659 ();
 sg13g2_fill_2 FILLER_53_663 ();
 sg13g2_fill_1 FILLER_53_665 ();
 sg13g2_fill_2 FILLER_53_718 ();
 sg13g2_fill_1 FILLER_53_720 ();
 sg13g2_decap_4 FILLER_53_726 ();
 sg13g2_fill_2 FILLER_53_734 ();
 sg13g2_fill_1 FILLER_53_736 ();
 sg13g2_fill_1 FILLER_53_741 ();
 sg13g2_fill_2 FILLER_53_747 ();
 sg13g2_fill_1 FILLER_53_749 ();
 sg13g2_fill_2 FILLER_53_802 ();
 sg13g2_fill_2 FILLER_53_814 ();
 sg13g2_decap_4 FILLER_53_824 ();
 sg13g2_fill_1 FILLER_53_865 ();
 sg13g2_decap_8 FILLER_53_871 ();
 sg13g2_fill_1 FILLER_53_878 ();
 sg13g2_fill_1 FILLER_53_918 ();
 sg13g2_fill_2 FILLER_53_922 ();
 sg13g2_fill_1 FILLER_53_924 ();
 sg13g2_decap_8 FILLER_53_933 ();
 sg13g2_decap_8 FILLER_53_940 ();
 sg13g2_decap_8 FILLER_53_952 ();
 sg13g2_fill_1 FILLER_53_959 ();
 sg13g2_fill_1 FILLER_53_1019 ();
 sg13g2_decap_4 FILLER_53_1024 ();
 sg13g2_fill_2 FILLER_53_1028 ();
 sg13g2_decap_8 FILLER_53_1065 ();
 sg13g2_fill_2 FILLER_53_1076 ();
 sg13g2_decap_8 FILLER_53_1116 ();
 sg13g2_decap_8 FILLER_53_1123 ();
 sg13g2_decap_8 FILLER_53_1130 ();
 sg13g2_fill_2 FILLER_53_1137 ();
 sg13g2_fill_1 FILLER_53_1139 ();
 sg13g2_decap_8 FILLER_53_1145 ();
 sg13g2_decap_4 FILLER_53_1152 ();
 sg13g2_fill_1 FILLER_53_1161 ();
 sg13g2_fill_1 FILLER_53_1171 ();
 sg13g2_fill_1 FILLER_53_1177 ();
 sg13g2_fill_1 FILLER_53_1183 ();
 sg13g2_fill_1 FILLER_53_1210 ();
 sg13g2_fill_1 FILLER_53_1219 ();
 sg13g2_fill_1 FILLER_53_1229 ();
 sg13g2_decap_4 FILLER_53_1233 ();
 sg13g2_decap_8 FILLER_53_1279 ();
 sg13g2_decap_8 FILLER_53_1286 ();
 sg13g2_decap_8 FILLER_53_1293 ();
 sg13g2_decap_8 FILLER_53_1300 ();
 sg13g2_decap_8 FILLER_53_1307 ();
 sg13g2_decap_8 FILLER_53_1314 ();
 sg13g2_decap_4 FILLER_53_1321 ();
 sg13g2_fill_1 FILLER_53_1325 ();
 sg13g2_decap_4 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_4 ();
 sg13g2_fill_2 FILLER_54_10 ();
 sg13g2_fill_2 FILLER_54_17 ();
 sg13g2_fill_1 FILLER_54_19 ();
 sg13g2_fill_1 FILLER_54_28 ();
 sg13g2_fill_2 FILLER_54_47 ();
 sg13g2_decap_4 FILLER_54_62 ();
 sg13g2_fill_1 FILLER_54_71 ();
 sg13g2_fill_2 FILLER_54_106 ();
 sg13g2_fill_1 FILLER_54_113 ();
 sg13g2_fill_1 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_124 ();
 sg13g2_decap_8 FILLER_54_131 ();
 sg13g2_fill_1 FILLER_54_138 ();
 sg13g2_fill_1 FILLER_54_143 ();
 sg13g2_fill_1 FILLER_54_148 ();
 sg13g2_fill_1 FILLER_54_153 ();
 sg13g2_fill_2 FILLER_54_159 ();
 sg13g2_fill_1 FILLER_54_170 ();
 sg13g2_fill_2 FILLER_54_175 ();
 sg13g2_fill_1 FILLER_54_177 ();
 sg13g2_fill_2 FILLER_54_183 ();
 sg13g2_fill_2 FILLER_54_188 ();
 sg13g2_fill_1 FILLER_54_190 ();
 sg13g2_decap_8 FILLER_54_194 ();
 sg13g2_fill_2 FILLER_54_201 ();
 sg13g2_fill_1 FILLER_54_216 ();
 sg13g2_fill_1 FILLER_54_221 ();
 sg13g2_decap_4 FILLER_54_305 ();
 sg13g2_fill_2 FILLER_54_320 ();
 sg13g2_decap_4 FILLER_54_330 ();
 sg13g2_fill_2 FILLER_54_334 ();
 sg13g2_fill_2 FILLER_54_367 ();
 sg13g2_fill_1 FILLER_54_379 ();
 sg13g2_fill_2 FILLER_54_410 ();
 sg13g2_decap_4 FILLER_54_417 ();
 sg13g2_fill_2 FILLER_54_421 ();
 sg13g2_fill_1 FILLER_54_426 ();
 sg13g2_decap_4 FILLER_54_435 ();
 sg13g2_fill_1 FILLER_54_439 ();
 sg13g2_fill_1 FILLER_54_468 ();
 sg13g2_fill_1 FILLER_54_489 ();
 sg13g2_fill_1 FILLER_54_499 ();
 sg13g2_fill_1 FILLER_54_505 ();
 sg13g2_decap_4 FILLER_54_516 ();
 sg13g2_decap_8 FILLER_54_525 ();
 sg13g2_decap_4 FILLER_54_540 ();
 sg13g2_fill_1 FILLER_54_544 ();
 sg13g2_fill_2 FILLER_54_554 ();
 sg13g2_fill_1 FILLER_54_560 ();
 sg13g2_fill_2 FILLER_54_565 ();
 sg13g2_fill_1 FILLER_54_575 ();
 sg13g2_fill_2 FILLER_54_580 ();
 sg13g2_decap_8 FILLER_54_591 ();
 sg13g2_fill_1 FILLER_54_598 ();
 sg13g2_fill_1 FILLER_54_602 ();
 sg13g2_fill_1 FILLER_54_607 ();
 sg13g2_fill_1 FILLER_54_612 ();
 sg13g2_fill_2 FILLER_54_617 ();
 sg13g2_fill_1 FILLER_54_626 ();
 sg13g2_decap_8 FILLER_54_631 ();
 sg13g2_decap_8 FILLER_54_638 ();
 sg13g2_fill_2 FILLER_54_645 ();
 sg13g2_decap_4 FILLER_54_656 ();
 sg13g2_decap_4 FILLER_54_664 ();
 sg13g2_fill_2 FILLER_54_668 ();
 sg13g2_fill_2 FILLER_54_674 ();
 sg13g2_fill_1 FILLER_54_676 ();
 sg13g2_decap_4 FILLER_54_681 ();
 sg13g2_fill_1 FILLER_54_685 ();
 sg13g2_fill_1 FILLER_54_696 ();
 sg13g2_fill_2 FILLER_54_702 ();
 sg13g2_decap_8 FILLER_54_709 ();
 sg13g2_fill_2 FILLER_54_716 ();
 sg13g2_decap_4 FILLER_54_731 ();
 sg13g2_fill_1 FILLER_54_735 ();
 sg13g2_fill_1 FILLER_54_752 ();
 sg13g2_fill_2 FILLER_54_769 ();
 sg13g2_fill_2 FILLER_54_776 ();
 sg13g2_fill_1 FILLER_54_778 ();
 sg13g2_fill_2 FILLER_54_786 ();
 sg13g2_fill_1 FILLER_54_792 ();
 sg13g2_decap_8 FILLER_54_803 ();
 sg13g2_decap_8 FILLER_54_810 ();
 sg13g2_fill_2 FILLER_54_817 ();
 sg13g2_fill_1 FILLER_54_819 ();
 sg13g2_fill_1 FILLER_54_825 ();
 sg13g2_fill_2 FILLER_54_838 ();
 sg13g2_fill_1 FILLER_54_840 ();
 sg13g2_fill_2 FILLER_54_854 ();
 sg13g2_decap_8 FILLER_54_869 ();
 sg13g2_decap_8 FILLER_54_876 ();
 sg13g2_fill_1 FILLER_54_883 ();
 sg13g2_decap_8 FILLER_54_899 ();
 sg13g2_decap_4 FILLER_54_906 ();
 sg13g2_fill_1 FILLER_54_978 ();
 sg13g2_fill_2 FILLER_54_984 ();
 sg13g2_fill_2 FILLER_54_990 ();
 sg13g2_fill_2 FILLER_54_997 ();
 sg13g2_fill_1 FILLER_54_999 ();
 sg13g2_decap_8 FILLER_54_1004 ();
 sg13g2_decap_4 FILLER_54_1011 ();
 sg13g2_decap_8 FILLER_54_1066 ();
 sg13g2_decap_4 FILLER_54_1073 ();
 sg13g2_fill_2 FILLER_54_1090 ();
 sg13g2_fill_1 FILLER_54_1092 ();
 sg13g2_decap_8 FILLER_54_1101 ();
 sg13g2_decap_4 FILLER_54_1108 ();
 sg13g2_fill_2 FILLER_54_1116 ();
 sg13g2_fill_2 FILLER_54_1153 ();
 sg13g2_fill_1 FILLER_54_1196 ();
 sg13g2_fill_1 FILLER_54_1206 ();
 sg13g2_fill_1 FILLER_54_1211 ();
 sg13g2_fill_2 FILLER_54_1238 ();
 sg13g2_fill_1 FILLER_54_1240 ();
 sg13g2_fill_1 FILLER_54_1249 ();
 sg13g2_decap_4 FILLER_54_1254 ();
 sg13g2_fill_2 FILLER_54_1262 ();
 sg13g2_decap_8 FILLER_54_1268 ();
 sg13g2_decap_8 FILLER_54_1280 ();
 sg13g2_decap_8 FILLER_54_1287 ();
 sg13g2_decap_8 FILLER_54_1294 ();
 sg13g2_decap_8 FILLER_54_1301 ();
 sg13g2_decap_8 FILLER_54_1308 ();
 sg13g2_decap_8 FILLER_54_1315 ();
 sg13g2_decap_4 FILLER_54_1322 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_26 ();
 sg13g2_fill_1 FILLER_55_35 ();
 sg13g2_fill_1 FILLER_55_50 ();
 sg13g2_decap_8 FILLER_55_62 ();
 sg13g2_decap_8 FILLER_55_69 ();
 sg13g2_fill_2 FILLER_55_76 ();
 sg13g2_decap_8 FILLER_55_83 ();
 sg13g2_fill_2 FILLER_55_90 ();
 sg13g2_fill_2 FILLER_55_100 ();
 sg13g2_decap_4 FILLER_55_106 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_fill_2 FILLER_55_142 ();
 sg13g2_fill_1 FILLER_55_144 ();
 sg13g2_fill_2 FILLER_55_158 ();
 sg13g2_fill_1 FILLER_55_160 ();
 sg13g2_fill_1 FILLER_55_183 ();
 sg13g2_decap_4 FILLER_55_204 ();
 sg13g2_decap_8 FILLER_55_242 ();
 sg13g2_decap_8 FILLER_55_249 ();
 sg13g2_fill_2 FILLER_55_256 ();
 sg13g2_fill_2 FILLER_55_263 ();
 sg13g2_fill_1 FILLER_55_269 ();
 sg13g2_fill_1 FILLER_55_283 ();
 sg13g2_fill_1 FILLER_55_289 ();
 sg13g2_decap_4 FILLER_55_297 ();
 sg13g2_decap_4 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_318 ();
 sg13g2_decap_4 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_330 ();
 sg13g2_fill_1 FILLER_55_332 ();
 sg13g2_decap_4 FILLER_55_336 ();
 sg13g2_fill_1 FILLER_55_340 ();
 sg13g2_decap_8 FILLER_55_379 ();
 sg13g2_fill_2 FILLER_55_390 ();
 sg13g2_fill_1 FILLER_55_392 ();
 sg13g2_decap_4 FILLER_55_423 ();
 sg13g2_decap_8 FILLER_55_432 ();
 sg13g2_fill_2 FILLER_55_439 ();
 sg13g2_fill_1 FILLER_55_441 ();
 sg13g2_fill_2 FILLER_55_454 ();
 sg13g2_fill_1 FILLER_55_475 ();
 sg13g2_fill_1 FILLER_55_486 ();
 sg13g2_fill_1 FILLER_55_501 ();
 sg13g2_decap_4 FILLER_55_507 ();
 sg13g2_fill_1 FILLER_55_521 ();
 sg13g2_fill_2 FILLER_55_527 ();
 sg13g2_decap_8 FILLER_55_534 ();
 sg13g2_decap_8 FILLER_55_541 ();
 sg13g2_fill_2 FILLER_55_548 ();
 sg13g2_fill_2 FILLER_55_554 ();
 sg13g2_fill_1 FILLER_55_556 ();
 sg13g2_decap_4 FILLER_55_569 ();
 sg13g2_fill_1 FILLER_55_607 ();
 sg13g2_decap_8 FILLER_55_631 ();
 sg13g2_decap_4 FILLER_55_638 ();
 sg13g2_fill_2 FILLER_55_668 ();
 sg13g2_fill_2 FILLER_55_696 ();
 sg13g2_fill_1 FILLER_55_698 ();
 sg13g2_fill_1 FILLER_55_725 ();
 sg13g2_fill_2 FILLER_55_731 ();
 sg13g2_fill_1 FILLER_55_733 ();
 sg13g2_fill_1 FILLER_55_753 ();
 sg13g2_decap_8 FILLER_55_758 ();
 sg13g2_decap_8 FILLER_55_769 ();
 sg13g2_fill_1 FILLER_55_780 ();
 sg13g2_fill_1 FILLER_55_829 ();
 sg13g2_fill_2 FILLER_55_891 ();
 sg13g2_fill_1 FILLER_55_902 ();
 sg13g2_fill_2 FILLER_55_923 ();
 sg13g2_decap_8 FILLER_55_929 ();
 sg13g2_decap_4 FILLER_55_936 ();
 sg13g2_fill_2 FILLER_55_940 ();
 sg13g2_fill_1 FILLER_55_950 ();
 sg13g2_decap_4 FILLER_55_955 ();
 sg13g2_fill_1 FILLER_55_959 ();
 sg13g2_fill_2 FILLER_55_987 ();
 sg13g2_fill_1 FILLER_55_1045 ();
 sg13g2_decap_4 FILLER_55_1051 ();
 sg13g2_decap_4 FILLER_55_1081 ();
 sg13g2_fill_2 FILLER_55_1085 ();
 sg13g2_decap_8 FILLER_55_1125 ();
 sg13g2_decap_4 FILLER_55_1132 ();
 sg13g2_fill_2 FILLER_55_1140 ();
 sg13g2_decap_8 FILLER_55_1147 ();
 sg13g2_decap_4 FILLER_55_1154 ();
 sg13g2_fill_1 FILLER_55_1158 ();
 sg13g2_fill_2 FILLER_55_1163 ();
 sg13g2_fill_1 FILLER_55_1165 ();
 sg13g2_fill_1 FILLER_55_1170 ();
 sg13g2_fill_1 FILLER_55_1187 ();
 sg13g2_fill_1 FILLER_55_1219 ();
 sg13g2_decap_8 FILLER_55_1225 ();
 sg13g2_decap_8 FILLER_55_1232 ();
 sg13g2_fill_2 FILLER_55_1239 ();
 sg13g2_fill_1 FILLER_55_1241 ();
 sg13g2_decap_4 FILLER_55_1247 ();
 sg13g2_decap_8 FILLER_55_1282 ();
 sg13g2_decap_8 FILLER_55_1289 ();
 sg13g2_decap_8 FILLER_55_1296 ();
 sg13g2_decap_8 FILLER_55_1303 ();
 sg13g2_decap_8 FILLER_55_1310 ();
 sg13g2_decap_8 FILLER_55_1317 ();
 sg13g2_fill_2 FILLER_55_1324 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_27 ();
 sg13g2_fill_1 FILLER_56_34 ();
 sg13g2_fill_2 FILLER_56_39 ();
 sg13g2_fill_1 FILLER_56_41 ();
 sg13g2_fill_2 FILLER_56_51 ();
 sg13g2_decap_8 FILLER_56_57 ();
 sg13g2_fill_1 FILLER_56_64 ();
 sg13g2_fill_1 FILLER_56_95 ();
 sg13g2_decap_8 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_116 ();
 sg13g2_fill_1 FILLER_56_118 ();
 sg13g2_decap_4 FILLER_56_123 ();
 sg13g2_fill_1 FILLER_56_127 ();
 sg13g2_fill_1 FILLER_56_136 ();
 sg13g2_fill_2 FILLER_56_141 ();
 sg13g2_decap_4 FILLER_56_151 ();
 sg13g2_fill_2 FILLER_56_155 ();
 sg13g2_fill_1 FILLER_56_162 ();
 sg13g2_fill_2 FILLER_56_167 ();
 sg13g2_fill_1 FILLER_56_169 ();
 sg13g2_fill_1 FILLER_56_174 ();
 sg13g2_fill_1 FILLER_56_179 ();
 sg13g2_decap_4 FILLER_56_184 ();
 sg13g2_fill_1 FILLER_56_214 ();
 sg13g2_fill_1 FILLER_56_228 ();
 sg13g2_decap_8 FILLER_56_243 ();
 sg13g2_decap_8 FILLER_56_250 ();
 sg13g2_fill_2 FILLER_56_279 ();
 sg13g2_fill_2 FILLER_56_291 ();
 sg13g2_decap_4 FILLER_56_323 ();
 sg13g2_fill_1 FILLER_56_327 ();
 sg13g2_fill_2 FILLER_56_331 ();
 sg13g2_fill_1 FILLER_56_337 ();
 sg13g2_decap_8 FILLER_56_382 ();
 sg13g2_decap_8 FILLER_56_389 ();
 sg13g2_fill_2 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_403 ();
 sg13g2_decap_8 FILLER_56_408 ();
 sg13g2_fill_1 FILLER_56_424 ();
 sg13g2_decap_8 FILLER_56_431 ();
 sg13g2_decap_8 FILLER_56_438 ();
 sg13g2_decap_8 FILLER_56_445 ();
 sg13g2_fill_1 FILLER_56_470 ();
 sg13g2_fill_2 FILLER_56_484 ();
 sg13g2_fill_1 FILLER_56_486 ();
 sg13g2_decap_4 FILLER_56_511 ();
 sg13g2_fill_1 FILLER_56_515 ();
 sg13g2_fill_1 FILLER_56_537 ();
 sg13g2_decap_8 FILLER_56_543 ();
 sg13g2_decap_8 FILLER_56_550 ();
 sg13g2_fill_2 FILLER_56_557 ();
 sg13g2_fill_1 FILLER_56_559 ();
 sg13g2_decap_8 FILLER_56_568 ();
 sg13g2_decap_8 FILLER_56_584 ();
 sg13g2_decap_8 FILLER_56_591 ();
 sg13g2_fill_1 FILLER_56_606 ();
 sg13g2_fill_2 FILLER_56_611 ();
 sg13g2_fill_2 FILLER_56_616 ();
 sg13g2_decap_8 FILLER_56_622 ();
 sg13g2_decap_8 FILLER_56_629 ();
 sg13g2_decap_8 FILLER_56_636 ();
 sg13g2_fill_1 FILLER_56_643 ();
 sg13g2_decap_4 FILLER_56_648 ();
 sg13g2_fill_2 FILLER_56_652 ();
 sg13g2_decap_4 FILLER_56_659 ();
 sg13g2_fill_2 FILLER_56_663 ();
 sg13g2_fill_2 FILLER_56_668 ();
 sg13g2_fill_1 FILLER_56_670 ();
 sg13g2_fill_1 FILLER_56_676 ();
 sg13g2_decap_8 FILLER_56_684 ();
 sg13g2_fill_1 FILLER_56_691 ();
 sg13g2_fill_2 FILLER_56_704 ();
 sg13g2_decap_4 FILLER_56_742 ();
 sg13g2_fill_2 FILLER_56_746 ();
 sg13g2_fill_1 FILLER_56_751 ();
 sg13g2_fill_2 FILLER_56_791 ();
 sg13g2_fill_2 FILLER_56_798 ();
 sg13g2_decap_8 FILLER_56_803 ();
 sg13g2_fill_1 FILLER_56_810 ();
 sg13g2_decap_8 FILLER_56_815 ();
 sg13g2_fill_2 FILLER_56_822 ();
 sg13g2_decap_4 FILLER_56_832 ();
 sg13g2_decap_8 FILLER_56_840 ();
 sg13g2_fill_2 FILLER_56_847 ();
 sg13g2_fill_2 FILLER_56_853 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_fill_1 FILLER_56_862 ();
 sg13g2_fill_2 FILLER_56_867 ();
 sg13g2_fill_1 FILLER_56_869 ();
 sg13g2_fill_2 FILLER_56_874 ();
 sg13g2_fill_1 FILLER_56_876 ();
 sg13g2_fill_1 FILLER_56_882 ();
 sg13g2_fill_1 FILLER_56_917 ();
 sg13g2_decap_8 FILLER_56_923 ();
 sg13g2_decap_4 FILLER_56_930 ();
 sg13g2_fill_2 FILLER_56_934 ();
 sg13g2_fill_1 FILLER_56_939 ();
 sg13g2_decap_8 FILLER_56_949 ();
 sg13g2_fill_2 FILLER_56_961 ();
 sg13g2_fill_2 FILLER_56_968 ();
 sg13g2_decap_4 FILLER_56_974 ();
 sg13g2_fill_1 FILLER_56_991 ();
 sg13g2_fill_1 FILLER_56_996 ();
 sg13g2_decap_8 FILLER_56_1003 ();
 sg13g2_fill_2 FILLER_56_1010 ();
 sg13g2_decap_8 FILLER_56_1028 ();
 sg13g2_fill_2 FILLER_56_1035 ();
 sg13g2_fill_2 FILLER_56_1041 ();
 sg13g2_fill_1 FILLER_56_1043 ();
 sg13g2_decap_4 FILLER_56_1067 ();
 sg13g2_decap_8 FILLER_56_1106 ();
 sg13g2_fill_2 FILLER_56_1117 ();
 sg13g2_fill_2 FILLER_56_1154 ();
 sg13g2_fill_2 FILLER_56_1170 ();
 sg13g2_fill_1 FILLER_56_1181 ();
 sg13g2_fill_2 FILLER_56_1189 ();
 sg13g2_fill_1 FILLER_56_1196 ();
 sg13g2_decap_8 FILLER_56_1208 ();
 sg13g2_decap_8 FILLER_56_1215 ();
 sg13g2_fill_2 FILLER_56_1222 ();
 sg13g2_decap_4 FILLER_56_1228 ();
 sg13g2_fill_2 FILLER_56_1253 ();
 sg13g2_decap_8 FILLER_56_1293 ();
 sg13g2_decap_8 FILLER_56_1300 ();
 sg13g2_decap_8 FILLER_56_1307 ();
 sg13g2_decap_8 FILLER_56_1314 ();
 sg13g2_decap_4 FILLER_56_1321 ();
 sg13g2_fill_1 FILLER_56_1325 ();
 sg13g2_decap_4 FILLER_57_51 ();
 sg13g2_fill_2 FILLER_57_64 ();
 sg13g2_fill_2 FILLER_57_70 ();
 sg13g2_fill_1 FILLER_57_72 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_fill_2 FILLER_57_84 ();
 sg13g2_fill_1 FILLER_57_86 ();
 sg13g2_fill_1 FILLER_57_90 ();
 sg13g2_fill_1 FILLER_57_96 ();
 sg13g2_fill_1 FILLER_57_103 ();
 sg13g2_decap_8 FILLER_57_110 ();
 sg13g2_decap_8 FILLER_57_117 ();
 sg13g2_decap_4 FILLER_57_124 ();
 sg13g2_fill_2 FILLER_57_128 ();
 sg13g2_fill_1 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_228 ();
 sg13g2_fill_1 FILLER_57_230 ();
 sg13g2_decap_8 FILLER_57_236 ();
 sg13g2_fill_2 FILLER_57_243 ();
 sg13g2_fill_2 FILLER_57_250 ();
 sg13g2_decap_4 FILLER_57_256 ();
 sg13g2_fill_2 FILLER_57_264 ();
 sg13g2_fill_1 FILLER_57_283 ();
 sg13g2_fill_1 FILLER_57_288 ();
 sg13g2_decap_8 FILLER_57_293 ();
 sg13g2_decap_8 FILLER_57_300 ();
 sg13g2_decap_4 FILLER_57_307 ();
 sg13g2_fill_1 FILLER_57_311 ();
 sg13g2_decap_8 FILLER_57_350 ();
 sg13g2_fill_1 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_362 ();
 sg13g2_decap_4 FILLER_57_369 ();
 sg13g2_fill_1 FILLER_57_380 ();
 sg13g2_fill_2 FILLER_57_396 ();
 sg13g2_decap_8 FILLER_57_402 ();
 sg13g2_fill_1 FILLER_57_409 ();
 sg13g2_fill_2 FILLER_57_458 ();
 sg13g2_fill_1 FILLER_57_464 ();
 sg13g2_fill_2 FILLER_57_473 ();
 sg13g2_fill_1 FILLER_57_475 ();
 sg13g2_fill_1 FILLER_57_480 ();
 sg13g2_fill_2 FILLER_57_486 ();
 sg13g2_fill_1 FILLER_57_488 ();
 sg13g2_fill_2 FILLER_57_504 ();
 sg13g2_decap_4 FILLER_57_511 ();
 sg13g2_fill_1 FILLER_57_515 ();
 sg13g2_fill_1 FILLER_57_529 ();
 sg13g2_decap_4 FILLER_57_545 ();
 sg13g2_fill_1 FILLER_57_549 ();
 sg13g2_decap_8 FILLER_57_554 ();
 sg13g2_fill_1 FILLER_57_585 ();
 sg13g2_fill_2 FILLER_57_590 ();
 sg13g2_fill_1 FILLER_57_607 ();
 sg13g2_decap_4 FILLER_57_613 ();
 sg13g2_fill_1 FILLER_57_617 ();
 sg13g2_decap_4 FILLER_57_626 ();
 sg13g2_decap_8 FILLER_57_683 ();
 sg13g2_decap_8 FILLER_57_690 ();
 sg13g2_fill_2 FILLER_57_704 ();
 sg13g2_fill_1 FILLER_57_716 ();
 sg13g2_fill_2 FILLER_57_721 ();
 sg13g2_fill_1 FILLER_57_723 ();
 sg13g2_decap_8 FILLER_57_759 ();
 sg13g2_fill_1 FILLER_57_770 ();
 sg13g2_fill_1 FILLER_57_779 ();
 sg13g2_fill_2 FILLER_57_790 ();
 sg13g2_fill_2 FILLER_57_823 ();
 sg13g2_fill_1 FILLER_57_845 ();
 sg13g2_fill_1 FILLER_57_860 ();
 sg13g2_decap_4 FILLER_57_873 ();
 sg13g2_fill_2 FILLER_57_884 ();
 sg13g2_fill_1 FILLER_57_886 ();
 sg13g2_fill_2 FILLER_57_896 ();
 sg13g2_fill_1 FILLER_57_898 ();
 sg13g2_decap_4 FILLER_57_903 ();
 sg13g2_fill_1 FILLER_57_921 ();
 sg13g2_decap_4 FILLER_57_983 ();
 sg13g2_fill_1 FILLER_57_987 ();
 sg13g2_fill_1 FILLER_57_991 ();
 sg13g2_fill_2 FILLER_57_1023 ();
 sg13g2_fill_1 FILLER_57_1025 ();
 sg13g2_fill_2 FILLER_57_1030 ();
 sg13g2_fill_1 FILLER_57_1044 ();
 sg13g2_decap_4 FILLER_57_1058 ();
 sg13g2_decap_8 FILLER_57_1070 ();
 sg13g2_decap_8 FILLER_57_1077 ();
 sg13g2_decap_8 FILLER_57_1092 ();
 sg13g2_fill_2 FILLER_57_1099 ();
 sg13g2_fill_1 FILLER_57_1106 ();
 sg13g2_fill_2 FILLER_57_1115 ();
 sg13g2_fill_1 FILLER_57_1117 ();
 sg13g2_decap_8 FILLER_57_1137 ();
 sg13g2_fill_1 FILLER_57_1144 ();
 sg13g2_fill_1 FILLER_57_1157 ();
 sg13g2_decap_8 FILLER_57_1162 ();
 sg13g2_decap_8 FILLER_57_1169 ();
 sg13g2_decap_4 FILLER_57_1176 ();
 sg13g2_fill_2 FILLER_57_1192 ();
 sg13g2_fill_1 FILLER_57_1206 ();
 sg13g2_decap_4 FILLER_57_1215 ();
 sg13g2_fill_1 FILLER_57_1219 ();
 sg13g2_decap_4 FILLER_57_1228 ();
 sg13g2_fill_2 FILLER_57_1232 ();
 sg13g2_decap_4 FILLER_57_1239 ();
 sg13g2_fill_2 FILLER_57_1243 ();
 sg13g2_fill_2 FILLER_57_1253 ();
 sg13g2_fill_1 FILLER_57_1261 ();
 sg13g2_decap_8 FILLER_57_1318 ();
 sg13g2_fill_1 FILLER_57_1325 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_11 ();
 sg13g2_decap_8 FILLER_58_18 ();
 sg13g2_decap_8 FILLER_58_30 ();
 sg13g2_decap_4 FILLER_58_37 ();
 sg13g2_fill_2 FILLER_58_41 ();
 sg13g2_fill_2 FILLER_58_53 ();
 sg13g2_fill_1 FILLER_58_55 ();
 sg13g2_fill_1 FILLER_58_116 ();
 sg13g2_fill_2 FILLER_58_148 ();
 sg13g2_fill_1 FILLER_58_150 ();
 sg13g2_fill_2 FILLER_58_155 ();
 sg13g2_fill_1 FILLER_58_157 ();
 sg13g2_fill_2 FILLER_58_167 ();
 sg13g2_fill_1 FILLER_58_169 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_fill_2 FILLER_58_195 ();
 sg13g2_fill_2 FILLER_58_206 ();
 sg13g2_fill_1 FILLER_58_260 ();
 sg13g2_fill_1 FILLER_58_273 ();
 sg13g2_fill_2 FILLER_58_283 ();
 sg13g2_decap_8 FILLER_58_323 ();
 sg13g2_decap_8 FILLER_58_330 ();
 sg13g2_decap_4 FILLER_58_337 ();
 sg13g2_fill_2 FILLER_58_344 ();
 sg13g2_fill_1 FILLER_58_385 ();
 sg13g2_fill_1 FILLER_58_394 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_fill_1 FILLER_58_412 ();
 sg13g2_fill_1 FILLER_58_432 ();
 sg13g2_decap_8 FILLER_58_443 ();
 sg13g2_decap_8 FILLER_58_450 ();
 sg13g2_decap_8 FILLER_58_457 ();
 sg13g2_fill_1 FILLER_58_472 ();
 sg13g2_fill_1 FILLER_58_497 ();
 sg13g2_fill_1 FILLER_58_520 ();
 sg13g2_fill_1 FILLER_58_530 ();
 sg13g2_decap_4 FILLER_58_540 ();
 sg13g2_decap_8 FILLER_58_555 ();
 sg13g2_decap_8 FILLER_58_562 ();
 sg13g2_fill_2 FILLER_58_594 ();
 sg13g2_decap_4 FILLER_58_613 ();
 sg13g2_fill_1 FILLER_58_617 ();
 sg13g2_fill_2 FILLER_58_647 ();
 sg13g2_fill_1 FILLER_58_668 ();
 sg13g2_fill_1 FILLER_58_673 ();
 sg13g2_fill_2 FILLER_58_736 ();
 sg13g2_decap_8 FILLER_58_742 ();
 sg13g2_decap_8 FILLER_58_749 ();
 sg13g2_decap_4 FILLER_58_756 ();
 sg13g2_decap_4 FILLER_58_800 ();
 sg13g2_fill_2 FILLER_58_804 ();
 sg13g2_decap_8 FILLER_58_810 ();
 sg13g2_decap_8 FILLER_58_817 ();
 sg13g2_fill_2 FILLER_58_824 ();
 sg13g2_fill_1 FILLER_58_826 ();
 sg13g2_fill_2 FILLER_58_831 ();
 sg13g2_fill_1 FILLER_58_833 ();
 sg13g2_decap_4 FILLER_58_844 ();
 sg13g2_fill_2 FILLER_58_848 ();
 sg13g2_fill_2 FILLER_58_862 ();
 sg13g2_fill_1 FILLER_58_917 ();
 sg13g2_decap_4 FILLER_58_923 ();
 sg13g2_fill_1 FILLER_58_927 ();
 sg13g2_decap_8 FILLER_58_932 ();
 sg13g2_fill_2 FILLER_58_939 ();
 sg13g2_fill_2 FILLER_58_950 ();
 sg13g2_decap_4 FILLER_58_956 ();
 sg13g2_decap_8 FILLER_58_964 ();
 sg13g2_fill_1 FILLER_58_971 ();
 sg13g2_fill_1 FILLER_58_1007 ();
 sg13g2_decap_8 FILLER_58_1012 ();
 sg13g2_decap_4 FILLER_58_1019 ();
 sg13g2_fill_2 FILLER_58_1030 ();
 sg13g2_fill_1 FILLER_58_1032 ();
 sg13g2_fill_2 FILLER_58_1046 ();
 sg13g2_decap_4 FILLER_58_1057 ();
 sg13g2_fill_1 FILLER_58_1061 ();
 sg13g2_fill_2 FILLER_58_1078 ();
 sg13g2_fill_1 FILLER_58_1080 ();
 sg13g2_fill_2 FILLER_58_1095 ();
 sg13g2_fill_1 FILLER_58_1107 ();
 sg13g2_fill_1 FILLER_58_1116 ();
 sg13g2_fill_1 FILLER_58_1120 ();
 sg13g2_fill_1 FILLER_58_1125 ();
 sg13g2_fill_1 FILLER_58_1130 ();
 sg13g2_decap_4 FILLER_58_1136 ();
 sg13g2_fill_1 FILLER_58_1140 ();
 sg13g2_decap_8 FILLER_58_1145 ();
 sg13g2_fill_1 FILLER_58_1152 ();
 sg13g2_fill_1 FILLER_58_1179 ();
 sg13g2_fill_2 FILLER_58_1183 ();
 sg13g2_fill_1 FILLER_58_1185 ();
 sg13g2_fill_1 FILLER_58_1238 ();
 sg13g2_decap_8 FILLER_58_1248 ();
 sg13g2_fill_2 FILLER_58_1255 ();
 sg13g2_fill_1 FILLER_58_1257 ();
 sg13g2_decap_8 FILLER_58_1310 ();
 sg13g2_decap_8 FILLER_58_1317 ();
 sg13g2_fill_2 FILLER_58_1324 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_4 FILLER_59_14 ();
 sg13g2_fill_1 FILLER_59_18 ();
 sg13g2_fill_1 FILLER_59_54 ();
 sg13g2_fill_2 FILLER_59_67 ();
 sg13g2_fill_1 FILLER_59_74 ();
 sg13g2_fill_1 FILLER_59_80 ();
 sg13g2_decap_8 FILLER_59_93 ();
 sg13g2_decap_4 FILLER_59_100 ();
 sg13g2_fill_2 FILLER_59_104 ();
 sg13g2_fill_2 FILLER_59_110 ();
 sg13g2_decap_4 FILLER_59_116 ();
 sg13g2_decap_4 FILLER_59_124 ();
 sg13g2_decap_8 FILLER_59_132 ();
 sg13g2_fill_2 FILLER_59_139 ();
 sg13g2_decap_8 FILLER_59_144 ();
 sg13g2_fill_2 FILLER_59_151 ();
 sg13g2_fill_2 FILLER_59_157 ();
 sg13g2_fill_1 FILLER_59_163 ();
 sg13g2_fill_1 FILLER_59_169 ();
 sg13g2_decap_4 FILLER_59_180 ();
 sg13g2_fill_2 FILLER_59_184 ();
 sg13g2_decap_4 FILLER_59_220 ();
 sg13g2_fill_2 FILLER_59_228 ();
 sg13g2_decap_8 FILLER_59_239 ();
 sg13g2_decap_4 FILLER_59_246 ();
 sg13g2_fill_2 FILLER_59_250 ();
 sg13g2_decap_8 FILLER_59_255 ();
 sg13g2_fill_2 FILLER_59_262 ();
 sg13g2_decap_4 FILLER_59_273 ();
 sg13g2_decap_4 FILLER_59_282 ();
 sg13g2_decap_4 FILLER_59_295 ();
 sg13g2_fill_2 FILLER_59_303 ();
 sg13g2_decap_8 FILLER_59_309 ();
 sg13g2_decap_8 FILLER_59_316 ();
 sg13g2_decap_8 FILLER_59_323 ();
 sg13g2_fill_1 FILLER_59_330 ();
 sg13g2_fill_2 FILLER_59_361 ();
 sg13g2_fill_1 FILLER_59_363 ();
 sg13g2_decap_8 FILLER_59_368 ();
 sg13g2_fill_2 FILLER_59_375 ();
 sg13g2_fill_1 FILLER_59_377 ();
 sg13g2_fill_2 FILLER_59_382 ();
 sg13g2_fill_1 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_402 ();
 sg13g2_fill_2 FILLER_59_409 ();
 sg13g2_fill_2 FILLER_59_416 ();
 sg13g2_fill_1 FILLER_59_435 ();
 sg13g2_decap_4 FILLER_59_466 ();
 sg13g2_fill_1 FILLER_59_470 ();
 sg13g2_fill_1 FILLER_59_498 ();
 sg13g2_fill_1 FILLER_59_516 ();
 sg13g2_fill_2 FILLER_59_521 ();
 sg13g2_fill_2 FILLER_59_527 ();
 sg13g2_fill_1 FILLER_59_529 ();
 sg13g2_fill_2 FILLER_59_535 ();
 sg13g2_decap_8 FILLER_59_541 ();
 sg13g2_fill_1 FILLER_59_548 ();
 sg13g2_decap_8 FILLER_59_553 ();
 sg13g2_decap_8 FILLER_59_560 ();
 sg13g2_decap_8 FILLER_59_567 ();
 sg13g2_decap_8 FILLER_59_574 ();
 sg13g2_decap_4 FILLER_59_581 ();
 sg13g2_fill_2 FILLER_59_585 ();
 sg13g2_decap_4 FILLER_59_621 ();
 sg13g2_decap_4 FILLER_59_637 ();
 sg13g2_fill_1 FILLER_59_641 ();
 sg13g2_fill_2 FILLER_59_646 ();
 sg13g2_fill_2 FILLER_59_651 ();
 sg13g2_fill_1 FILLER_59_653 ();
 sg13g2_fill_1 FILLER_59_659 ();
 sg13g2_fill_2 FILLER_59_669 ();
 sg13g2_fill_1 FILLER_59_671 ();
 sg13g2_decap_8 FILLER_59_676 ();
 sg13g2_decap_4 FILLER_59_683 ();
 sg13g2_fill_1 FILLER_59_687 ();
 sg13g2_decap_4 FILLER_59_693 ();
 sg13g2_fill_2 FILLER_59_701 ();
 sg13g2_fill_1 FILLER_59_703 ();
 sg13g2_fill_1 FILLER_59_708 ();
 sg13g2_fill_1 FILLER_59_713 ();
 sg13g2_fill_2 FILLER_59_728 ();
 sg13g2_fill_2 FILLER_59_788 ();
 sg13g2_decap_4 FILLER_59_821 ();
 sg13g2_fill_1 FILLER_59_825 ();
 sg13g2_fill_2 FILLER_59_834 ();
 sg13g2_fill_1 FILLER_59_840 ();
 sg13g2_fill_2 FILLER_59_852 ();
 sg13g2_fill_1 FILLER_59_854 ();
 sg13g2_fill_2 FILLER_59_875 ();
 sg13g2_decap_4 FILLER_59_889 ();
 sg13g2_decap_4 FILLER_59_897 ();
 sg13g2_fill_1 FILLER_59_901 ();
 sg13g2_decap_8 FILLER_59_906 ();
 sg13g2_fill_2 FILLER_59_913 ();
 sg13g2_fill_1 FILLER_59_915 ();
 sg13g2_fill_1 FILLER_59_947 ();
 sg13g2_decap_4 FILLER_59_982 ();
 sg13g2_fill_1 FILLER_59_986 ();
 sg13g2_decap_8 FILLER_59_991 ();
 sg13g2_decap_8 FILLER_59_998 ();
 sg13g2_fill_1 FILLER_59_1005 ();
 sg13g2_decap_8 FILLER_59_1010 ();
 sg13g2_decap_4 FILLER_59_1017 ();
 sg13g2_fill_2 FILLER_59_1021 ();
 sg13g2_decap_8 FILLER_59_1032 ();
 sg13g2_fill_2 FILLER_59_1039 ();
 sg13g2_fill_1 FILLER_59_1041 ();
 sg13g2_fill_2 FILLER_59_1068 ();
 sg13g2_fill_1 FILLER_59_1070 ();
 sg13g2_fill_2 FILLER_59_1133 ();
 sg13g2_decap_8 FILLER_59_1165 ();
 sg13g2_decap_4 FILLER_59_1172 ();
 sg13g2_fill_1 FILLER_59_1176 ();
 sg13g2_decap_8 FILLER_59_1185 ();
 sg13g2_fill_1 FILLER_59_1192 ();
 sg13g2_decap_8 FILLER_59_1197 ();
 sg13g2_decap_4 FILLER_59_1204 ();
 sg13g2_fill_1 FILLER_59_1208 ();
 sg13g2_decap_8 FILLER_59_1213 ();
 sg13g2_fill_1 FILLER_59_1220 ();
 sg13g2_decap_8 FILLER_59_1226 ();
 sg13g2_fill_1 FILLER_59_1233 ();
 sg13g2_decap_4 FILLER_59_1264 ();
 sg13g2_fill_1 FILLER_59_1268 ();
 sg13g2_fill_2 FILLER_59_1277 ();
 sg13g2_fill_2 FILLER_59_1284 ();
 sg13g2_fill_1 FILLER_59_1286 ();
 sg13g2_fill_1 FILLER_59_1291 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_decap_8 FILLER_60_46 ();
 sg13g2_decap_4 FILLER_60_53 ();
 sg13g2_fill_1 FILLER_60_57 ();
 sg13g2_fill_1 FILLER_60_71 ();
 sg13g2_fill_2 FILLER_60_77 ();
 sg13g2_fill_2 FILLER_60_83 ();
 sg13g2_fill_2 FILLER_60_111 ();
 sg13g2_fill_1 FILLER_60_113 ();
 sg13g2_fill_2 FILLER_60_126 ();
 sg13g2_fill_1 FILLER_60_154 ();
 sg13g2_fill_1 FILLER_60_159 ();
 sg13g2_fill_1 FILLER_60_164 ();
 sg13g2_fill_1 FILLER_60_173 ();
 sg13g2_decap_8 FILLER_60_178 ();
 sg13g2_fill_1 FILLER_60_190 ();
 sg13g2_fill_1 FILLER_60_203 ();
 sg13g2_fill_1 FILLER_60_209 ();
 sg13g2_fill_2 FILLER_60_219 ();
 sg13g2_fill_2 FILLER_60_255 ();
 sg13g2_fill_2 FILLER_60_276 ();
 sg13g2_fill_1 FILLER_60_278 ();
 sg13g2_fill_2 FILLER_60_289 ();
 sg13g2_fill_2 FILLER_60_295 ();
 sg13g2_fill_1 FILLER_60_297 ();
 sg13g2_decap_8 FILLER_60_324 ();
 sg13g2_fill_1 FILLER_60_331 ();
 sg13g2_decap_4 FILLER_60_347 ();
 sg13g2_fill_2 FILLER_60_351 ();
 sg13g2_fill_2 FILLER_60_403 ();
 sg13g2_fill_2 FILLER_60_434 ();
 sg13g2_fill_2 FILLER_60_441 ();
 sg13g2_decap_8 FILLER_60_451 ();
 sg13g2_decap_8 FILLER_60_471 ();
 sg13g2_fill_1 FILLER_60_478 ();
 sg13g2_fill_2 FILLER_60_483 ();
 sg13g2_fill_1 FILLER_60_485 ();
 sg13g2_fill_2 FILLER_60_519 ();
 sg13g2_fill_2 FILLER_60_526 ();
 sg13g2_decap_4 FILLER_60_532 ();
 sg13g2_fill_2 FILLER_60_536 ();
 sg13g2_fill_1 FILLER_60_542 ();
 sg13g2_fill_1 FILLER_60_569 ();
 sg13g2_fill_1 FILLER_60_596 ();
 sg13g2_fill_2 FILLER_60_607 ();
 sg13g2_decap_4 FILLER_60_666 ();
 sg13g2_fill_1 FILLER_60_670 ();
 sg13g2_fill_1 FILLER_60_675 ();
 sg13g2_fill_1 FILLER_60_705 ();
 sg13g2_fill_2 FILLER_60_710 ();
 sg13g2_fill_2 FILLER_60_717 ();
 sg13g2_fill_2 FILLER_60_745 ();
 sg13g2_fill_1 FILLER_60_747 ();
 sg13g2_decap_8 FILLER_60_752 ();
 sg13g2_decap_8 FILLER_60_794 ();
 sg13g2_fill_2 FILLER_60_801 ();
 sg13g2_fill_1 FILLER_60_803 ();
 sg13g2_decap_8 FILLER_60_808 ();
 sg13g2_decap_8 FILLER_60_815 ();
 sg13g2_decap_4 FILLER_60_822 ();
 sg13g2_fill_1 FILLER_60_835 ();
 sg13g2_decap_8 FILLER_60_840 ();
 sg13g2_decap_8 FILLER_60_847 ();
 sg13g2_fill_2 FILLER_60_854 ();
 sg13g2_fill_1 FILLER_60_856 ();
 sg13g2_fill_2 FILLER_60_874 ();
 sg13g2_fill_1 FILLER_60_876 ();
 sg13g2_decap_8 FILLER_60_888 ();
 sg13g2_decap_4 FILLER_60_895 ();
 sg13g2_fill_1 FILLER_60_899 ();
 sg13g2_fill_2 FILLER_60_930 ();
 sg13g2_decap_8 FILLER_60_936 ();
 sg13g2_decap_8 FILLER_60_943 ();
 sg13g2_decap_8 FILLER_60_950 ();
 sg13g2_fill_2 FILLER_60_957 ();
 sg13g2_decap_8 FILLER_60_964 ();
 sg13g2_decap_4 FILLER_60_971 ();
 sg13g2_fill_1 FILLER_60_975 ();
 sg13g2_decap_4 FILLER_60_994 ();
 sg13g2_fill_2 FILLER_60_998 ();
 sg13g2_fill_1 FILLER_60_1038 ();
 sg13g2_fill_1 FILLER_60_1056 ();
 sg13g2_fill_2 FILLER_60_1061 ();
 sg13g2_fill_2 FILLER_60_1067 ();
 sg13g2_fill_2 FILLER_60_1074 ();
 sg13g2_fill_1 FILLER_60_1076 ();
 sg13g2_fill_2 FILLER_60_1086 ();
 sg13g2_fill_1 FILLER_60_1093 ();
 sg13g2_decap_8 FILLER_60_1098 ();
 sg13g2_fill_2 FILLER_60_1109 ();
 sg13g2_fill_1 FILLER_60_1111 ();
 sg13g2_fill_1 FILLER_60_1125 ();
 sg13g2_decap_8 FILLER_60_1129 ();
 sg13g2_decap_4 FILLER_60_1136 ();
 sg13g2_fill_2 FILLER_60_1140 ();
 sg13g2_decap_8 FILLER_60_1146 ();
 sg13g2_decap_8 FILLER_60_1153 ();
 sg13g2_decap_4 FILLER_60_1160 ();
 sg13g2_fill_1 FILLER_60_1164 ();
 sg13g2_fill_2 FILLER_60_1191 ();
 sg13g2_fill_1 FILLER_60_1193 ();
 sg13g2_decap_4 FILLER_60_1198 ();
 sg13g2_fill_1 FILLER_60_1202 ();
 sg13g2_fill_1 FILLER_60_1242 ();
 sg13g2_fill_2 FILLER_60_1247 ();
 sg13g2_fill_2 FILLER_60_1288 ();
 sg13g2_fill_1 FILLER_60_1290 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_31 ();
 sg13g2_decap_4 FILLER_61_38 ();
 sg13g2_decap_8 FILLER_61_46 ();
 sg13g2_fill_2 FILLER_61_53 ();
 sg13g2_fill_1 FILLER_61_55 ();
 sg13g2_fill_1 FILLER_61_60 ();
 sg13g2_fill_1 FILLER_61_65 ();
 sg13g2_decap_4 FILLER_61_75 ();
 sg13g2_fill_2 FILLER_61_93 ();
 sg13g2_decap_4 FILLER_61_100 ();
 sg13g2_decap_4 FILLER_61_108 ();
 sg13g2_fill_2 FILLER_61_124 ();
 sg13g2_decap_4 FILLER_61_130 ();
 sg13g2_decap_4 FILLER_61_138 ();
 sg13g2_fill_2 FILLER_61_147 ();
 sg13g2_fill_1 FILLER_61_149 ();
 sg13g2_decap_8 FILLER_61_172 ();
 sg13g2_decap_8 FILLER_61_179 ();
 sg13g2_fill_2 FILLER_61_186 ();
 sg13g2_fill_1 FILLER_61_188 ();
 sg13g2_fill_2 FILLER_61_194 ();
 sg13g2_fill_2 FILLER_61_200 ();
 sg13g2_fill_1 FILLER_61_202 ();
 sg13g2_fill_1 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_212 ();
 sg13g2_fill_2 FILLER_61_217 ();
 sg13g2_decap_8 FILLER_61_223 ();
 sg13g2_fill_2 FILLER_61_230 ();
 sg13g2_fill_2 FILLER_61_244 ();
 sg13g2_decap_4 FILLER_61_250 ();
 sg13g2_decap_4 FILLER_61_257 ();
 sg13g2_fill_1 FILLER_61_261 ();
 sg13g2_fill_2 FILLER_61_266 ();
 sg13g2_fill_1 FILLER_61_268 ();
 sg13g2_decap_4 FILLER_61_273 ();
 sg13g2_fill_2 FILLER_61_277 ();
 sg13g2_fill_2 FILLER_61_283 ();
 sg13g2_fill_1 FILLER_61_285 ();
 sg13g2_decap_4 FILLER_61_312 ();
 sg13g2_fill_2 FILLER_61_316 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_fill_1 FILLER_61_324 ();
 sg13g2_decap_4 FILLER_61_329 ();
 sg13g2_fill_1 FILLER_61_333 ();
 sg13g2_fill_2 FILLER_61_343 ();
 sg13g2_fill_2 FILLER_61_349 ();
 sg13g2_fill_1 FILLER_61_351 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_fill_1 FILLER_61_386 ();
 sg13g2_fill_2 FILLER_61_411 ();
 sg13g2_fill_1 FILLER_61_450 ();
 sg13g2_decap_4 FILLER_61_455 ();
 sg13g2_fill_1 FILLER_61_459 ();
 sg13g2_fill_2 FILLER_61_464 ();
 sg13g2_fill_1 FILLER_61_466 ();
 sg13g2_decap_8 FILLER_61_502 ();
 sg13g2_decap_8 FILLER_61_509 ();
 sg13g2_decap_8 FILLER_61_516 ();
 sg13g2_decap_8 FILLER_61_523 ();
 sg13g2_fill_1 FILLER_61_530 ();
 sg13g2_fill_2 FILLER_61_565 ();
 sg13g2_fill_1 FILLER_61_567 ();
 sg13g2_decap_4 FILLER_61_572 ();
 sg13g2_fill_2 FILLER_61_576 ();
 sg13g2_decap_8 FILLER_61_582 ();
 sg13g2_fill_2 FILLER_61_589 ();
 sg13g2_fill_1 FILLER_61_604 ();
 sg13g2_fill_1 FILLER_61_631 ();
 sg13g2_fill_2 FILLER_61_641 ();
 sg13g2_fill_1 FILLER_61_652 ();
 sg13g2_fill_1 FILLER_61_657 ();
 sg13g2_fill_1 FILLER_61_663 ();
 sg13g2_fill_1 FILLER_61_668 ();
 sg13g2_fill_2 FILLER_61_673 ();
 sg13g2_fill_2 FILLER_61_680 ();
 sg13g2_fill_1 FILLER_61_682 ();
 sg13g2_decap_4 FILLER_61_687 ();
 sg13g2_decap_4 FILLER_61_696 ();
 sg13g2_fill_1 FILLER_61_700 ();
 sg13g2_fill_1 FILLER_61_710 ();
 sg13g2_fill_2 FILLER_61_721 ();
 sg13g2_fill_1 FILLER_61_728 ();
 sg13g2_decap_8 FILLER_61_737 ();
 sg13g2_decap_8 FILLER_61_744 ();
 sg13g2_fill_2 FILLER_61_751 ();
 sg13g2_decap_4 FILLER_61_757 ();
 sg13g2_decap_8 FILLER_61_765 ();
 sg13g2_decap_8 FILLER_61_772 ();
 sg13g2_decap_8 FILLER_61_779 ();
 sg13g2_decap_8 FILLER_61_786 ();
 sg13g2_fill_1 FILLER_61_793 ();
 sg13g2_decap_4 FILLER_61_820 ();
 sg13g2_fill_2 FILLER_61_824 ();
 sg13g2_fill_1 FILLER_61_864 ();
 sg13g2_fill_1 FILLER_61_899 ();
 sg13g2_fill_2 FILLER_61_917 ();
 sg13g2_fill_1 FILLER_61_919 ();
 sg13g2_fill_2 FILLER_61_930 ();
 sg13g2_fill_1 FILLER_61_932 ();
 sg13g2_decap_8 FILLER_61_937 ();
 sg13g2_fill_1 FILLER_61_951 ();
 sg13g2_fill_1 FILLER_61_970 ();
 sg13g2_fill_2 FILLER_61_981 ();
 sg13g2_decap_8 FILLER_61_1016 ();
 sg13g2_fill_2 FILLER_61_1023 ();
 sg13g2_fill_1 FILLER_61_1029 ();
 sg13g2_fill_1 FILLER_61_1038 ();
 sg13g2_fill_1 FILLER_61_1043 ();
 sg13g2_decap_8 FILLER_61_1049 ();
 sg13g2_fill_2 FILLER_61_1056 ();
 sg13g2_fill_2 FILLER_61_1084 ();
 sg13g2_fill_1 FILLER_61_1086 ();
 sg13g2_decap_4 FILLER_61_1113 ();
 sg13g2_fill_1 FILLER_61_1125 ();
 sg13g2_fill_2 FILLER_61_1160 ();
 sg13g2_fill_1 FILLER_61_1162 ();
 sg13g2_fill_2 FILLER_61_1168 ();
 sg13g2_fill_1 FILLER_61_1170 ();
 sg13g2_decap_4 FILLER_61_1213 ();
 sg13g2_fill_1 FILLER_61_1217 ();
 sg13g2_decap_8 FILLER_61_1222 ();
 sg13g2_fill_1 FILLER_61_1229 ();
 sg13g2_fill_1 FILLER_61_1272 ();
 sg13g2_fill_1 FILLER_61_1277 ();
 sg13g2_decap_8 FILLER_61_1282 ();
 sg13g2_decap_4 FILLER_61_1289 ();
 sg13g2_fill_1 FILLER_61_1293 ();
 sg13g2_fill_1 FILLER_61_1299 ();
 sg13g2_fill_1 FILLER_62_74 ();
 sg13g2_fill_2 FILLER_62_79 ();
 sg13g2_fill_1 FILLER_62_81 ();
 sg13g2_fill_1 FILLER_62_87 ();
 sg13g2_fill_2 FILLER_62_92 ();
 sg13g2_decap_4 FILLER_62_99 ();
 sg13g2_fill_1 FILLER_62_103 ();
 sg13g2_fill_1 FILLER_62_143 ();
 sg13g2_decap_4 FILLER_62_152 ();
 sg13g2_fill_1 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_179 ();
 sg13g2_fill_1 FILLER_62_186 ();
 sg13g2_decap_8 FILLER_62_191 ();
 sg13g2_decap_8 FILLER_62_198 ();
 sg13g2_decap_4 FILLER_62_205 ();
 sg13g2_fill_2 FILLER_62_209 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_4 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_258 ();
 sg13g2_decap_8 FILLER_62_265 ();
 sg13g2_decap_8 FILLER_62_276 ();
 sg13g2_decap_8 FILLER_62_287 ();
 sg13g2_fill_1 FILLER_62_294 ();
 sg13g2_fill_1 FILLER_62_299 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_fill_2 FILLER_62_331 ();
 sg13g2_fill_2 FILLER_62_389 ();
 sg13g2_decap_4 FILLER_62_417 ();
 sg13g2_fill_2 FILLER_62_421 ();
 sg13g2_decap_4 FILLER_62_428 ();
 sg13g2_fill_2 FILLER_62_432 ();
 sg13g2_decap_8 FILLER_62_467 ();
 sg13g2_decap_4 FILLER_62_474 ();
 sg13g2_fill_2 FILLER_62_478 ();
 sg13g2_fill_2 FILLER_62_487 ();
 sg13g2_fill_1 FILLER_62_489 ();
 sg13g2_decap_4 FILLER_62_494 ();
 sg13g2_fill_2 FILLER_62_498 ();
 sg13g2_decap_8 FILLER_62_504 ();
 sg13g2_decap_8 FILLER_62_511 ();
 sg13g2_decap_4 FILLER_62_522 ();
 sg13g2_fill_2 FILLER_62_552 ();
 sg13g2_fill_2 FILLER_62_558 ();
 sg13g2_fill_2 FILLER_62_564 ();
 sg13g2_fill_1 FILLER_62_566 ();
 sg13g2_fill_1 FILLER_62_572 ();
 sg13g2_decap_8 FILLER_62_577 ();
 sg13g2_decap_8 FILLER_62_584 ();
 sg13g2_fill_1 FILLER_62_591 ();
 sg13g2_decap_4 FILLER_62_604 ();
 sg13g2_decap_8 FILLER_62_621 ();
 sg13g2_fill_2 FILLER_62_628 ();
 sg13g2_decap_8 FILLER_62_635 ();
 sg13g2_decap_4 FILLER_62_642 ();
 sg13g2_fill_1 FILLER_62_646 ();
 sg13g2_fill_2 FILLER_62_651 ();
 sg13g2_fill_1 FILLER_62_653 ();
 sg13g2_fill_2 FILLER_62_661 ();
 sg13g2_fill_1 FILLER_62_663 ();
 sg13g2_decap_4 FILLER_62_693 ();
 sg13g2_fill_2 FILLER_62_697 ();
 sg13g2_fill_1 FILLER_62_703 ();
 sg13g2_fill_2 FILLER_62_709 ();
 sg13g2_fill_2 FILLER_62_718 ();
 sg13g2_fill_2 FILLER_62_727 ();
 sg13g2_fill_2 FILLER_62_747 ();
 sg13g2_fill_2 FILLER_62_759 ();
 sg13g2_fill_1 FILLER_62_761 ();
 sg13g2_fill_2 FILLER_62_767 ();
 sg13g2_fill_2 FILLER_62_783 ();
 sg13g2_fill_1 FILLER_62_785 ();
 sg13g2_decap_8 FILLER_62_804 ();
 sg13g2_decap_4 FILLER_62_811 ();
 sg13g2_fill_2 FILLER_62_815 ();
 sg13g2_fill_1 FILLER_62_831 ();
 sg13g2_decap_8 FILLER_62_845 ();
 sg13g2_fill_2 FILLER_62_864 ();
 sg13g2_fill_1 FILLER_62_866 ();
 sg13g2_fill_2 FILLER_62_872 ();
 sg13g2_fill_1 FILLER_62_874 ();
 sg13g2_fill_2 FILLER_62_884 ();
 sg13g2_fill_1 FILLER_62_886 ();
 sg13g2_decap_4 FILLER_62_891 ();
 sg13g2_decap_8 FILLER_62_904 ();
 sg13g2_fill_2 FILLER_62_911 ();
 sg13g2_fill_2 FILLER_62_917 ();
 sg13g2_fill_1 FILLER_62_919 ();
 sg13g2_decap_4 FILLER_62_956 ();
 sg13g2_decap_8 FILLER_62_965 ();
 sg13g2_fill_1 FILLER_62_972 ();
 sg13g2_fill_1 FILLER_62_991 ();
 sg13g2_fill_1 FILLER_62_997 ();
 sg13g2_fill_1 FILLER_62_1007 ();
 sg13g2_fill_1 FILLER_62_1012 ();
 sg13g2_fill_1 FILLER_62_1019 ();
 sg13g2_fill_2 FILLER_62_1051 ();
 sg13g2_fill_2 FILLER_62_1060 ();
 sg13g2_fill_2 FILLER_62_1088 ();
 sg13g2_fill_1 FILLER_62_1090 ();
 sg13g2_fill_2 FILLER_62_1104 ();
 sg13g2_fill_2 FILLER_62_1116 ();
 sg13g2_fill_1 FILLER_62_1118 ();
 sg13g2_fill_2 FILLER_62_1131 ();
 sg13g2_fill_1 FILLER_62_1133 ();
 sg13g2_fill_2 FILLER_62_1139 ();
 sg13g2_fill_1 FILLER_62_1141 ();
 sg13g2_decap_4 FILLER_62_1189 ();
 sg13g2_decap_8 FILLER_62_1197 ();
 sg13g2_decap_8 FILLER_62_1204 ();
 sg13g2_decap_8 FILLER_62_1211 ();
 sg13g2_decap_4 FILLER_62_1235 ();
 sg13g2_fill_2 FILLER_62_1243 ();
 sg13g2_decap_8 FILLER_62_1252 ();
 sg13g2_decap_8 FILLER_62_1259 ();
 sg13g2_fill_2 FILLER_62_1266 ();
 sg13g2_fill_1 FILLER_62_1268 ();
 sg13g2_decap_8 FILLER_62_1315 ();
 sg13g2_decap_4 FILLER_62_1322 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_8 ();
 sg13g2_fill_1 FILLER_63_13 ();
 sg13g2_decap_8 FILLER_63_44 ();
 sg13g2_decap_8 FILLER_63_51 ();
 sg13g2_fill_2 FILLER_63_58 ();
 sg13g2_fill_2 FILLER_63_73 ();
 sg13g2_fill_1 FILLER_63_75 ();
 sg13g2_fill_1 FILLER_63_100 ();
 sg13g2_decap_8 FILLER_63_127 ();
 sg13g2_decap_8 FILLER_63_134 ();
 sg13g2_decap_4 FILLER_63_141 ();
 sg13g2_decap_8 FILLER_63_150 ();
 sg13g2_decap_4 FILLER_63_157 ();
 sg13g2_fill_2 FILLER_63_166 ();
 sg13g2_decap_4 FILLER_63_221 ();
 sg13g2_fill_1 FILLER_63_229 ();
 sg13g2_fill_2 FILLER_63_235 ();
 sg13g2_fill_1 FILLER_63_247 ();
 sg13g2_fill_1 FILLER_63_262 ();
 sg13g2_fill_2 FILLER_63_289 ();
 sg13g2_decap_4 FILLER_63_296 ();
 sg13g2_decap_8 FILLER_63_311 ();
 sg13g2_fill_1 FILLER_63_318 ();
 sg13g2_decap_8 FILLER_63_327 ();
 sg13g2_decap_8 FILLER_63_334 ();
 sg13g2_decap_8 FILLER_63_341 ();
 sg13g2_decap_4 FILLER_63_348 ();
 sg13g2_fill_2 FILLER_63_352 ();
 sg13g2_decap_8 FILLER_63_361 ();
 sg13g2_fill_2 FILLER_63_368 ();
 sg13g2_decap_8 FILLER_63_374 ();
 sg13g2_decap_8 FILLER_63_381 ();
 sg13g2_decap_8 FILLER_63_388 ();
 sg13g2_fill_2 FILLER_63_395 ();
 sg13g2_fill_1 FILLER_63_397 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_decap_8 FILLER_63_409 ();
 sg13g2_fill_1 FILLER_63_416 ();
 sg13g2_decap_8 FILLER_63_430 ();
 sg13g2_decap_8 FILLER_63_437 ();
 sg13g2_decap_8 FILLER_63_444 ();
 sg13g2_fill_1 FILLER_63_451 ();
 sg13g2_fill_1 FILLER_63_456 ();
 sg13g2_decap_8 FILLER_63_461 ();
 sg13g2_fill_2 FILLER_63_468 ();
 sg13g2_fill_1 FILLER_63_470 ();
 sg13g2_fill_1 FILLER_63_502 ();
 sg13g2_decap_8 FILLER_63_538 ();
 sg13g2_fill_2 FILLER_63_545 ();
 sg13g2_fill_1 FILLER_63_547 ();
 sg13g2_decap_4 FILLER_63_552 ();
 sg13g2_fill_2 FILLER_63_556 ();
 sg13g2_fill_2 FILLER_63_563 ();
 sg13g2_fill_1 FILLER_63_565 ();
 sg13g2_decap_4 FILLER_63_600 ();
 sg13g2_fill_1 FILLER_63_604 ();
 sg13g2_fill_1 FILLER_63_635 ();
 sg13g2_decap_8 FILLER_63_645 ();
 sg13g2_fill_1 FILLER_63_652 ();
 sg13g2_fill_2 FILLER_63_663 ();
 sg13g2_fill_1 FILLER_63_670 ();
 sg13g2_fill_2 FILLER_63_705 ();
 sg13g2_fill_1 FILLER_63_707 ();
 sg13g2_decap_8 FILLER_63_729 ();
 sg13g2_decap_8 FILLER_63_736 ();
 sg13g2_decap_4 FILLER_63_743 ();
 sg13g2_fill_2 FILLER_63_773 ();
 sg13g2_fill_1 FILLER_63_775 ();
 sg13g2_decap_4 FILLER_63_781 ();
 sg13g2_fill_2 FILLER_63_785 ();
 sg13g2_fill_1 FILLER_63_792 ();
 sg13g2_fill_1 FILLER_63_822 ();
 sg13g2_decap_8 FILLER_63_849 ();
 sg13g2_decap_4 FILLER_63_856 ();
 sg13g2_fill_2 FILLER_63_864 ();
 sg13g2_fill_1 FILLER_63_866 ();
 sg13g2_decap_4 FILLER_63_876 ();
 sg13g2_decap_4 FILLER_63_887 ();
 sg13g2_fill_1 FILLER_63_891 ();
 sg13g2_decap_8 FILLER_63_922 ();
 sg13g2_decap_8 FILLER_63_929 ();
 sg13g2_decap_8 FILLER_63_936 ();
 sg13g2_fill_1 FILLER_63_943 ();
 sg13g2_decap_8 FILLER_63_948 ();
 sg13g2_decap_4 FILLER_63_955 ();
 sg13g2_decap_4 FILLER_63_963 ();
 sg13g2_fill_1 FILLER_63_967 ();
 sg13g2_fill_2 FILLER_63_992 ();
 sg13g2_fill_2 FILLER_63_1020 ();
 sg13g2_fill_2 FILLER_63_1033 ();
 sg13g2_fill_1 FILLER_63_1035 ();
 sg13g2_fill_2 FILLER_63_1041 ();
 sg13g2_fill_1 FILLER_63_1043 ();
 sg13g2_decap_8 FILLER_63_1049 ();
 sg13g2_decap_4 FILLER_63_1056 ();
 sg13g2_decap_4 FILLER_63_1064 ();
 sg13g2_decap_4 FILLER_63_1077 ();
 sg13g2_fill_1 FILLER_63_1092 ();
 sg13g2_fill_2 FILLER_63_1119 ();
 sg13g2_decap_4 FILLER_63_1125 ();
 sg13g2_decap_8 FILLER_63_1143 ();
 sg13g2_fill_2 FILLER_63_1150 ();
 sg13g2_fill_1 FILLER_63_1152 ();
 sg13g2_fill_2 FILLER_63_1160 ();
 sg13g2_fill_1 FILLER_63_1174 ();
 sg13g2_fill_1 FILLER_63_1180 ();
 sg13g2_fill_1 FILLER_63_1185 ();
 sg13g2_decap_4 FILLER_63_1212 ();
 sg13g2_fill_2 FILLER_63_1216 ();
 sg13g2_decap_8 FILLER_63_1263 ();
 sg13g2_decap_4 FILLER_63_1270 ();
 sg13g2_fill_1 FILLER_63_1274 ();
 sg13g2_fill_1 FILLER_63_1280 ();
 sg13g2_decap_8 FILLER_63_1300 ();
 sg13g2_decap_8 FILLER_63_1307 ();
 sg13g2_decap_8 FILLER_63_1314 ();
 sg13g2_decap_4 FILLER_63_1321 ();
 sg13g2_fill_1 FILLER_63_1325 ();
 sg13g2_fill_1 FILLER_64_35 ();
 sg13g2_fill_1 FILLER_64_44 ();
 sg13g2_fill_1 FILLER_64_49 ();
 sg13g2_fill_1 FILLER_64_55 ();
 sg13g2_fill_1 FILLER_64_68 ();
 sg13g2_fill_1 FILLER_64_73 ();
 sg13g2_decap_8 FILLER_64_87 ();
 sg13g2_fill_2 FILLER_64_94 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_1 FILLER_64_105 ();
 sg13g2_fill_2 FILLER_64_110 ();
 sg13g2_fill_1 FILLER_64_142 ();
 sg13g2_decap_4 FILLER_64_148 ();
 sg13g2_decap_4 FILLER_64_155 ();
 sg13g2_fill_2 FILLER_64_194 ();
 sg13g2_fill_1 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_202 ();
 sg13g2_decap_8 FILLER_64_213 ();
 sg13g2_fill_2 FILLER_64_245 ();
 sg13g2_fill_1 FILLER_64_251 ();
 sg13g2_fill_2 FILLER_64_266 ();
 sg13g2_fill_1 FILLER_64_268 ();
 sg13g2_decap_4 FILLER_64_273 ();
 sg13g2_fill_1 FILLER_64_303 ();
 sg13g2_fill_1 FILLER_64_312 ();
 sg13g2_decap_4 FILLER_64_317 ();
 sg13g2_fill_1 FILLER_64_321 ();
 sg13g2_fill_1 FILLER_64_334 ();
 sg13g2_fill_1 FILLER_64_344 ();
 sg13g2_fill_2 FILLER_64_371 ();
 sg13g2_fill_2 FILLER_64_404 ();
 sg13g2_fill_1 FILLER_64_411 ();
 sg13g2_fill_2 FILLER_64_416 ();
 sg13g2_fill_1 FILLER_64_444 ();
 sg13g2_decap_8 FILLER_64_476 ();
 sg13g2_fill_2 FILLER_64_483 ();
 sg13g2_fill_1 FILLER_64_485 ();
 sg13g2_fill_1 FILLER_64_498 ();
 sg13g2_fill_1 FILLER_64_503 ();
 sg13g2_decap_4 FILLER_64_511 ();
 sg13g2_fill_2 FILLER_64_515 ();
 sg13g2_fill_1 FILLER_64_521 ();
 sg13g2_decap_4 FILLER_64_525 ();
 sg13g2_fill_1 FILLER_64_529 ();
 sg13g2_fill_1 FILLER_64_564 ();
 sg13g2_fill_1 FILLER_64_580 ();
 sg13g2_fill_2 FILLER_64_642 ();
 sg13g2_decap_8 FILLER_64_649 ();
 sg13g2_decap_8 FILLER_64_656 ();
 sg13g2_decap_4 FILLER_64_663 ();
 sg13g2_fill_2 FILLER_64_667 ();
 sg13g2_decap_8 FILLER_64_674 ();
 sg13g2_fill_1 FILLER_64_681 ();
 sg13g2_fill_2 FILLER_64_690 ();
 sg13g2_fill_1 FILLER_64_692 ();
 sg13g2_fill_1 FILLER_64_698 ();
 sg13g2_fill_2 FILLER_64_707 ();
 sg13g2_fill_1 FILLER_64_747 ();
 sg13g2_fill_2 FILLER_64_753 ();
 sg13g2_fill_2 FILLER_64_763 ();
 sg13g2_fill_1 FILLER_64_765 ();
 sg13g2_fill_2 FILLER_64_799 ();
 sg13g2_fill_1 FILLER_64_801 ();
 sg13g2_fill_2 FILLER_64_814 ();
 sg13g2_fill_2 FILLER_64_820 ();
 sg13g2_fill_2 FILLER_64_827 ();
 sg13g2_fill_1 FILLER_64_842 ();
 sg13g2_fill_1 FILLER_64_848 ();
 sg13g2_decap_8 FILLER_64_853 ();
 sg13g2_decap_4 FILLER_64_860 ();
 sg13g2_fill_2 FILLER_64_864 ();
 sg13g2_decap_4 FILLER_64_892 ();
 sg13g2_fill_1 FILLER_64_896 ();
 sg13g2_fill_2 FILLER_64_901 ();
 sg13g2_fill_1 FILLER_64_903 ();
 sg13g2_decap_8 FILLER_64_911 ();
 sg13g2_fill_1 FILLER_64_918 ();
 sg13g2_fill_2 FILLER_64_967 ();
 sg13g2_fill_1 FILLER_64_975 ();
 sg13g2_decap_8 FILLER_64_981 ();
 sg13g2_decap_4 FILLER_64_988 ();
 sg13g2_decap_4 FILLER_64_997 ();
 sg13g2_fill_2 FILLER_64_1009 ();
 sg13g2_decap_8 FILLER_64_1021 ();
 sg13g2_fill_2 FILLER_64_1028 ();
 sg13g2_fill_1 FILLER_64_1030 ();
 sg13g2_decap_8 FILLER_64_1039 ();
 sg13g2_decap_8 FILLER_64_1046 ();
 sg13g2_fill_2 FILLER_64_1053 ();
 sg13g2_decap_4 FILLER_64_1060 ();
 sg13g2_fill_1 FILLER_64_1064 ();
 sg13g2_fill_2 FILLER_64_1091 ();
 sg13g2_fill_1 FILLER_64_1093 ();
 sg13g2_fill_2 FILLER_64_1103 ();
 sg13g2_fill_2 FILLER_64_1112 ();
 sg13g2_decap_4 FILLER_64_1118 ();
 sg13g2_fill_1 FILLER_64_1182 ();
 sg13g2_fill_2 FILLER_64_1187 ();
 sg13g2_fill_1 FILLER_64_1189 ();
 sg13g2_fill_2 FILLER_64_1216 ();
 sg13g2_fill_2 FILLER_64_1231 ();
 sg13g2_fill_1 FILLER_64_1233 ();
 sg13g2_fill_2 FILLER_64_1272 ();
 sg13g2_fill_1 FILLER_64_1274 ();
 sg13g2_fill_2 FILLER_64_1292 ();
 sg13g2_fill_1 FILLER_64_1294 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_11 ();
 sg13g2_fill_1 FILLER_65_15 ();
 sg13g2_fill_2 FILLER_65_20 ();
 sg13g2_fill_1 FILLER_65_22 ();
 sg13g2_fill_2 FILLER_65_27 ();
 sg13g2_decap_4 FILLER_65_39 ();
 sg13g2_fill_1 FILLER_65_66 ();
 sg13g2_fill_1 FILLER_65_79 ();
 sg13g2_fill_2 FILLER_65_88 ();
 sg13g2_decap_8 FILLER_65_100 ();
 sg13g2_fill_1 FILLER_65_107 ();
 sg13g2_fill_2 FILLER_65_114 ();
 sg13g2_fill_1 FILLER_65_116 ();
 sg13g2_fill_2 FILLER_65_126 ();
 sg13g2_fill_1 FILLER_65_128 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_fill_2 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_171 ();
 sg13g2_decap_8 FILLER_65_178 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_fill_2 FILLER_65_195 ();
 sg13g2_fill_1 FILLER_65_197 ();
 sg13g2_fill_2 FILLER_65_213 ();
 sg13g2_fill_1 FILLER_65_215 ();
 sg13g2_decap_8 FILLER_65_220 ();
 sg13g2_decap_4 FILLER_65_227 ();
 sg13g2_fill_1 FILLER_65_231 ();
 sg13g2_fill_2 FILLER_65_255 ();
 sg13g2_fill_1 FILLER_65_257 ();
 sg13g2_decap_8 FILLER_65_263 ();
 sg13g2_fill_1 FILLER_65_270 ();
 sg13g2_decap_4 FILLER_65_280 ();
 sg13g2_fill_1 FILLER_65_284 ();
 sg13g2_decap_8 FILLER_65_289 ();
 sg13g2_decap_8 FILLER_65_296 ();
 sg13g2_fill_2 FILLER_65_303 ();
 sg13g2_decap_4 FILLER_65_314 ();
 sg13g2_fill_2 FILLER_65_318 ();
 sg13g2_fill_2 FILLER_65_325 ();
 sg13g2_fill_2 FILLER_65_332 ();
 sg13g2_fill_2 FILLER_65_352 ();
 sg13g2_fill_1 FILLER_65_354 ();
 sg13g2_fill_1 FILLER_65_359 ();
 sg13g2_fill_1 FILLER_65_365 ();
 sg13g2_decap_4 FILLER_65_371 ();
 sg13g2_fill_1 FILLER_65_375 ();
 sg13g2_fill_1 FILLER_65_386 ();
 sg13g2_decap_4 FILLER_65_391 ();
 sg13g2_fill_2 FILLER_65_411 ();
 sg13g2_fill_2 FILLER_65_429 ();
 sg13g2_fill_1 FILLER_65_431 ();
 sg13g2_fill_1 FILLER_65_437 ();
 sg13g2_fill_2 FILLER_65_443 ();
 sg13g2_fill_2 FILLER_65_450 ();
 sg13g2_fill_2 FILLER_65_475 ();
 sg13g2_fill_1 FILLER_65_477 ();
 sg13g2_fill_1 FILLER_65_485 ();
 sg13g2_fill_2 FILLER_65_509 ();
 sg13g2_decap_4 FILLER_65_537 ();
 sg13g2_fill_2 FILLER_65_541 ();
 sg13g2_decap_8 FILLER_65_547 ();
 sg13g2_fill_2 FILLER_65_554 ();
 sg13g2_fill_1 FILLER_65_574 ();
 sg13g2_fill_1 FILLER_65_580 ();
 sg13g2_fill_1 FILLER_65_600 ();
 sg13g2_decap_8 FILLER_65_605 ();
 sg13g2_decap_4 FILLER_65_612 ();
 sg13g2_fill_1 FILLER_65_616 ();
 sg13g2_decap_8 FILLER_65_629 ();
 sg13g2_decap_8 FILLER_65_645 ();
 sg13g2_fill_2 FILLER_65_652 ();
 sg13g2_fill_1 FILLER_65_661 ();
 sg13g2_decap_8 FILLER_65_677 ();
 sg13g2_fill_1 FILLER_65_684 ();
 sg13g2_fill_1 FILLER_65_689 ();
 sg13g2_fill_2 FILLER_65_724 ();
 sg13g2_fill_1 FILLER_65_726 ();
 sg13g2_decap_8 FILLER_65_735 ();
 sg13g2_decap_4 FILLER_65_742 ();
 sg13g2_fill_1 FILLER_65_746 ();
 sg13g2_fill_2 FILLER_65_751 ();
 sg13g2_fill_1 FILLER_65_753 ();
 sg13g2_decap_8 FILLER_65_759 ();
 sg13g2_decap_8 FILLER_65_766 ();
 sg13g2_decap_4 FILLER_65_773 ();
 sg13g2_fill_1 FILLER_65_781 ();
 sg13g2_decap_8 FILLER_65_802 ();
 sg13g2_fill_1 FILLER_65_809 ();
 sg13g2_fill_2 FILLER_65_818 ();
 sg13g2_fill_1 FILLER_65_820 ();
 sg13g2_decap_4 FILLER_65_868 ();
 sg13g2_fill_2 FILLER_65_877 ();
 sg13g2_fill_1 FILLER_65_879 ();
 sg13g2_fill_1 FILLER_65_889 ();
 sg13g2_decap_4 FILLER_65_916 ();
 sg13g2_fill_2 FILLER_65_920 ();
 sg13g2_decap_4 FILLER_65_948 ();
 sg13g2_fill_1 FILLER_65_987 ();
 sg13g2_fill_1 FILLER_65_1022 ();
 sg13g2_fill_2 FILLER_65_1060 ();
 sg13g2_fill_1 FILLER_65_1065 ();
 sg13g2_fill_1 FILLER_65_1070 ();
 sg13g2_fill_1 FILLER_65_1075 ();
 sg13g2_fill_1 FILLER_65_1081 ();
 sg13g2_fill_2 FILLER_65_1088 ();
 sg13g2_decap_8 FILLER_65_1093 ();
 sg13g2_fill_2 FILLER_65_1100 ();
 sg13g2_fill_1 FILLER_65_1102 ();
 sg13g2_decap_4 FILLER_65_1120 ();
 sg13g2_fill_1 FILLER_65_1124 ();
 sg13g2_fill_2 FILLER_65_1130 ();
 sg13g2_decap_8 FILLER_65_1136 ();
 sg13g2_decap_8 FILLER_65_1143 ();
 sg13g2_fill_2 FILLER_65_1150 ();
 sg13g2_fill_2 FILLER_65_1155 ();
 sg13g2_fill_1 FILLER_65_1160 ();
 sg13g2_decap_8 FILLER_65_1165 ();
 sg13g2_fill_2 FILLER_65_1172 ();
 sg13g2_fill_2 FILLER_65_1178 ();
 sg13g2_fill_2 FILLER_65_1250 ();
 sg13g2_fill_2 FILLER_65_1256 ();
 sg13g2_fill_1 FILLER_65_1258 ();
 sg13g2_fill_2 FILLER_65_1308 ();
 sg13g2_fill_1 FILLER_65_1310 ();
 sg13g2_decap_8 FILLER_65_1315 ();
 sg13g2_decap_4 FILLER_65_1322 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_11 ();
 sg13g2_fill_1 FILLER_66_15 ();
 sg13g2_decap_4 FILLER_66_20 ();
 sg13g2_decap_8 FILLER_66_36 ();
 sg13g2_fill_2 FILLER_66_43 ();
 sg13g2_fill_1 FILLER_66_65 ();
 sg13g2_fill_2 FILLER_66_72 ();
 sg13g2_decap_4 FILLER_66_77 ();
 sg13g2_fill_2 FILLER_66_86 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_fill_1 FILLER_66_93 ();
 sg13g2_fill_2 FILLER_66_105 ();
 sg13g2_fill_2 FILLER_66_126 ();
 sg13g2_fill_1 FILLER_66_132 ();
 sg13g2_fill_2 FILLER_66_143 ();
 sg13g2_fill_2 FILLER_66_158 ();
 sg13g2_fill_2 FILLER_66_168 ();
 sg13g2_fill_1 FILLER_66_170 ();
 sg13g2_decap_4 FILLER_66_191 ();
 sg13g2_decap_8 FILLER_66_199 ();
 sg13g2_decap_8 FILLER_66_206 ();
 sg13g2_fill_2 FILLER_66_213 ();
 sg13g2_decap_4 FILLER_66_224 ();
 sg13g2_fill_2 FILLER_66_228 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_242 ();
 sg13g2_decap_4 FILLER_66_251 ();
 sg13g2_fill_2 FILLER_66_255 ();
 sg13g2_fill_2 FILLER_66_262 ();
 sg13g2_fill_1 FILLER_66_264 ();
 sg13g2_decap_4 FILLER_66_273 ();
 sg13g2_fill_2 FILLER_66_277 ();
 sg13g2_decap_4 FILLER_66_292 ();
 sg13g2_fill_2 FILLER_66_327 ();
 sg13g2_fill_1 FILLER_66_337 ();
 sg13g2_fill_1 FILLER_66_372 ();
 sg13g2_fill_2 FILLER_66_404 ();
 sg13g2_fill_2 FILLER_66_411 ();
 sg13g2_fill_1 FILLER_66_413 ();
 sg13g2_fill_2 FILLER_66_418 ();
 sg13g2_fill_1 FILLER_66_420 ();
 sg13g2_fill_2 FILLER_66_463 ();
 sg13g2_decap_4 FILLER_66_491 ();
 sg13g2_fill_2 FILLER_66_495 ();
 sg13g2_decap_8 FILLER_66_531 ();
 sg13g2_decap_4 FILLER_66_538 ();
 sg13g2_decap_8 FILLER_66_551 ();
 sg13g2_decap_4 FILLER_66_571 ();
 sg13g2_fill_2 FILLER_66_575 ();
 sg13g2_fill_2 FILLER_66_586 ();
 sg13g2_fill_1 FILLER_66_588 ();
 sg13g2_decap_8 FILLER_66_597 ();
 sg13g2_decap_8 FILLER_66_604 ();
 sg13g2_decap_8 FILLER_66_650 ();
 sg13g2_fill_1 FILLER_66_657 ();
 sg13g2_fill_2 FILLER_66_668 ();
 sg13g2_fill_1 FILLER_66_714 ();
 sg13g2_fill_1 FILLER_66_745 ();
 sg13g2_fill_1 FILLER_66_751 ();
 sg13g2_fill_1 FILLER_66_760 ();
 sg13g2_fill_2 FILLER_66_788 ();
 sg13g2_decap_8 FILLER_66_804 ();
 sg13g2_decap_4 FILLER_66_811 ();
 sg13g2_fill_2 FILLER_66_829 ();
 sg13g2_fill_1 FILLER_66_831 ();
 sg13g2_decap_8 FILLER_66_840 ();
 sg13g2_decap_4 FILLER_66_847 ();
 sg13g2_fill_2 FILLER_66_851 ();
 sg13g2_decap_4 FILLER_66_867 ();
 sg13g2_fill_1 FILLER_66_871 ();
 sg13g2_fill_1 FILLER_66_877 ();
 sg13g2_fill_1 FILLER_66_888 ();
 sg13g2_fill_1 FILLER_66_910 ();
 sg13g2_fill_1 FILLER_66_919 ();
 sg13g2_fill_2 FILLER_66_928 ();
 sg13g2_fill_1 FILLER_66_930 ();
 sg13g2_decap_8 FILLER_66_935 ();
 sg13g2_decap_4 FILLER_66_942 ();
 sg13g2_fill_2 FILLER_66_946 ();
 sg13g2_fill_1 FILLER_66_953 ();
 sg13g2_fill_1 FILLER_66_962 ();
 sg13g2_decap_8 FILLER_66_977 ();
 sg13g2_fill_2 FILLER_66_984 ();
 sg13g2_fill_1 FILLER_66_986 ();
 sg13g2_fill_1 FILLER_66_1013 ();
 sg13g2_fill_2 FILLER_66_1019 ();
 sg13g2_fill_1 FILLER_66_1021 ();
 sg13g2_decap_8 FILLER_66_1026 ();
 sg13g2_decap_8 FILLER_66_1033 ();
 sg13g2_decap_4 FILLER_66_1040 ();
 sg13g2_fill_1 FILLER_66_1044 ();
 sg13g2_fill_1 FILLER_66_1067 ();
 sg13g2_decap_8 FILLER_66_1098 ();
 sg13g2_fill_2 FILLER_66_1105 ();
 sg13g2_decap_4 FILLER_66_1116 ();
 sg13g2_fill_2 FILLER_66_1120 ();
 sg13g2_fill_1 FILLER_66_1158 ();
 sg13g2_fill_2 FILLER_66_1175 ();
 sg13g2_fill_1 FILLER_66_1177 ();
 sg13g2_decap_4 FILLER_66_1213 ();
 sg13g2_fill_1 FILLER_66_1217 ();
 sg13g2_decap_8 FILLER_66_1227 ();
 sg13g2_fill_1 FILLER_66_1234 ();
 sg13g2_fill_1 FILLER_66_1247 ();
 sg13g2_fill_1 FILLER_66_1256 ();
 sg13g2_fill_2 FILLER_66_1261 ();
 sg13g2_decap_4 FILLER_66_1267 ();
 sg13g2_fill_1 FILLER_66_1280 ();
 sg13g2_decap_4 FILLER_66_1284 ();
 sg13g2_fill_2 FILLER_66_1288 ();
 sg13g2_decap_8 FILLER_67_30 ();
 sg13g2_fill_1 FILLER_67_37 ();
 sg13g2_fill_1 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_62 ();
 sg13g2_fill_2 FILLER_67_69 ();
 sg13g2_fill_1 FILLER_67_76 ();
 sg13g2_fill_2 FILLER_67_100 ();
 sg13g2_fill_1 FILLER_67_102 ();
 sg13g2_decap_8 FILLER_67_125 ();
 sg13g2_fill_1 FILLER_67_132 ();
 sg13g2_fill_2 FILLER_67_155 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_decap_8 FILLER_67_163 ();
 sg13g2_decap_8 FILLER_67_170 ();
 sg13g2_decap_4 FILLER_67_177 ();
 sg13g2_fill_1 FILLER_67_186 ();
 sg13g2_decap_4 FILLER_67_191 ();
 sg13g2_decap_8 FILLER_67_207 ();
 sg13g2_decap_8 FILLER_67_214 ();
 sg13g2_decap_8 FILLER_67_221 ();
 sg13g2_fill_1 FILLER_67_235 ();
 sg13g2_fill_2 FILLER_67_260 ();
 sg13g2_decap_8 FILLER_67_271 ();
 sg13g2_fill_2 FILLER_67_286 ();
 sg13g2_decap_8 FILLER_67_297 ();
 sg13g2_fill_2 FILLER_67_304 ();
 sg13g2_fill_1 FILLER_67_306 ();
 sg13g2_decap_8 FILLER_67_311 ();
 sg13g2_decap_4 FILLER_67_318 ();
 sg13g2_decap_4 FILLER_67_326 ();
 sg13g2_decap_8 FILLER_67_337 ();
 sg13g2_decap_8 FILLER_67_344 ();
 sg13g2_fill_2 FILLER_67_359 ();
 sg13g2_fill_1 FILLER_67_361 ();
 sg13g2_decap_8 FILLER_67_373 ();
 sg13g2_decap_4 FILLER_67_380 ();
 sg13g2_decap_8 FILLER_67_388 ();
 sg13g2_decap_8 FILLER_67_395 ();
 sg13g2_fill_1 FILLER_67_440 ();
 sg13g2_fill_1 FILLER_67_446 ();
 sg13g2_fill_1 FILLER_67_452 ();
 sg13g2_fill_2 FILLER_67_456 ();
 sg13g2_fill_1 FILLER_67_475 ();
 sg13g2_decap_8 FILLER_67_484 ();
 sg13g2_fill_2 FILLER_67_491 ();
 sg13g2_fill_1 FILLER_67_493 ();
 sg13g2_decap_8 FILLER_67_504 ();
 sg13g2_fill_1 FILLER_67_511 ();
 sg13g2_fill_1 FILLER_67_516 ();
 sg13g2_fill_2 FILLER_67_547 ();
 sg13g2_decap_4 FILLER_67_559 ();
 sg13g2_fill_2 FILLER_67_563 ();
 sg13g2_decap_8 FILLER_67_573 ();
 sg13g2_decap_4 FILLER_67_580 ();
 sg13g2_fill_2 FILLER_67_584 ();
 sg13g2_decap_8 FILLER_67_592 ();
 sg13g2_decap_8 FILLER_67_599 ();
 sg13g2_decap_4 FILLER_67_606 ();
 sg13g2_fill_1 FILLER_67_610 ();
 sg13g2_fill_1 FILLER_67_650 ();
 sg13g2_fill_1 FILLER_67_678 ();
 sg13g2_decap_8 FILLER_67_684 ();
 sg13g2_fill_1 FILLER_67_691 ();
 sg13g2_decap_8 FILLER_67_699 ();
 sg13g2_fill_1 FILLER_67_706 ();
 sg13g2_decap_8 FILLER_67_730 ();
 sg13g2_fill_1 FILLER_67_737 ();
 sg13g2_fill_1 FILLER_67_757 ();
 sg13g2_decap_8 FILLER_67_770 ();
 sg13g2_decap_8 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_784 ();
 sg13g2_decap_4 FILLER_67_791 ();
 sg13g2_fill_2 FILLER_67_804 ();
 sg13g2_fill_1 FILLER_67_827 ();
 sg13g2_decap_8 FILLER_67_862 ();
 sg13g2_fill_2 FILLER_67_869 ();
 sg13g2_fill_1 FILLER_67_871 ();
 sg13g2_fill_2 FILLER_67_880 ();
 sg13g2_fill_1 FILLER_67_913 ();
 sg13g2_fill_2 FILLER_67_920 ();
 sg13g2_fill_1 FILLER_67_922 ();
 sg13g2_fill_2 FILLER_67_963 ();
 sg13g2_fill_1 FILLER_67_970 ();
 sg13g2_decap_8 FILLER_67_1006 ();
 sg13g2_fill_2 FILLER_67_1013 ();
 sg13g2_decap_8 FILLER_67_1045 ();
 sg13g2_decap_8 FILLER_67_1052 ();
 sg13g2_decap_8 FILLER_67_1059 ();
 sg13g2_decap_4 FILLER_67_1066 ();
 sg13g2_fill_1 FILLER_67_1070 ();
 sg13g2_fill_2 FILLER_67_1075 ();
 sg13g2_fill_2 FILLER_67_1082 ();
 sg13g2_fill_1 FILLER_67_1084 ();
 sg13g2_fill_2 FILLER_67_1098 ();
 sg13g2_fill_2 FILLER_67_1105 ();
 sg13g2_fill_1 FILLER_67_1107 ();
 sg13g2_decap_4 FILLER_67_1112 ();
 sg13g2_fill_2 FILLER_67_1116 ();
 sg13g2_fill_2 FILLER_67_1130 ();
 sg13g2_decap_4 FILLER_67_1137 ();
 sg13g2_fill_2 FILLER_67_1141 ();
 sg13g2_decap_8 FILLER_67_1153 ();
 sg13g2_decap_8 FILLER_67_1160 ();
 sg13g2_fill_2 FILLER_67_1167 ();
 sg13g2_fill_1 FILLER_67_1169 ();
 sg13g2_fill_2 FILLER_67_1174 ();
 sg13g2_fill_1 FILLER_67_1176 ();
 sg13g2_fill_1 FILLER_67_1200 ();
 sg13g2_fill_1 FILLER_67_1232 ();
 sg13g2_fill_2 FILLER_67_1237 ();
 sg13g2_fill_1 FILLER_67_1239 ();
 sg13g2_fill_2 FILLER_67_1292 ();
 sg13g2_fill_1 FILLER_67_1294 ();
 sg13g2_decap_8 FILLER_67_1299 ();
 sg13g2_fill_1 FILLER_67_1306 ();
 sg13g2_decap_8 FILLER_67_1311 ();
 sg13g2_decap_8 FILLER_67_1318 ();
 sg13g2_fill_1 FILLER_67_1325 ();
 sg13g2_fill_2 FILLER_68_26 ();
 sg13g2_fill_1 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_33 ();
 sg13g2_decap_4 FILLER_68_40 ();
 sg13g2_fill_1 FILLER_68_49 ();
 sg13g2_fill_1 FILLER_68_55 ();
 sg13g2_fill_1 FILLER_68_61 ();
 sg13g2_decap_8 FILLER_68_67 ();
 sg13g2_decap_8 FILLER_68_74 ();
 sg13g2_fill_1 FILLER_68_81 ();
 sg13g2_fill_2 FILLER_68_100 ();
 sg13g2_fill_1 FILLER_68_102 ();
 sg13g2_decap_4 FILLER_68_115 ();
 sg13g2_fill_1 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_125 ();
 sg13g2_decap_8 FILLER_68_132 ();
 sg13g2_fill_1 FILLER_68_139 ();
 sg13g2_fill_2 FILLER_68_144 ();
 sg13g2_fill_1 FILLER_68_146 ();
 sg13g2_fill_2 FILLER_68_192 ();
 sg13g2_fill_2 FILLER_68_219 ();
 sg13g2_fill_2 FILLER_68_237 ();
 sg13g2_fill_2 FILLER_68_246 ();
 sg13g2_fill_1 FILLER_68_280 ();
 sg13g2_fill_1 FILLER_68_285 ();
 sg13g2_decap_8 FILLER_68_299 ();
 sg13g2_fill_2 FILLER_68_341 ();
 sg13g2_fill_1 FILLER_68_343 ();
 sg13g2_decap_8 FILLER_68_370 ();
 sg13g2_fill_2 FILLER_68_377 ();
 sg13g2_decap_8 FILLER_68_383 ();
 sg13g2_decap_8 FILLER_68_390 ();
 sg13g2_decap_4 FILLER_68_397 ();
 sg13g2_decap_8 FILLER_68_406 ();
 sg13g2_decap_8 FILLER_68_413 ();
 sg13g2_decap_4 FILLER_68_420 ();
 sg13g2_fill_1 FILLER_68_424 ();
 sg13g2_decap_8 FILLER_68_431 ();
 sg13g2_decap_4 FILLER_68_438 ();
 sg13g2_fill_1 FILLER_68_442 ();
 sg13g2_decap_4 FILLER_68_474 ();
 sg13g2_fill_2 FILLER_68_478 ();
 sg13g2_decap_8 FILLER_68_510 ();
 sg13g2_decap_8 FILLER_68_517 ();
 sg13g2_decap_4 FILLER_68_524 ();
 sg13g2_decap_8 FILLER_68_532 ();
 sg13g2_decap_4 FILLER_68_539 ();
 sg13g2_fill_1 FILLER_68_543 ();
 sg13g2_fill_2 FILLER_68_559 ();
 sg13g2_fill_1 FILLER_68_564 ();
 sg13g2_fill_1 FILLER_68_570 ();
 sg13g2_fill_2 FILLER_68_580 ();
 sg13g2_fill_1 FILLER_68_582 ();
 sg13g2_decap_4 FILLER_68_595 ();
 sg13g2_fill_2 FILLER_68_599 ();
 sg13g2_decap_4 FILLER_68_627 ();
 sg13g2_fill_1 FILLER_68_631 ();
 sg13g2_fill_1 FILLER_68_640 ();
 sg13g2_decap_8 FILLER_68_650 ();
 sg13g2_decap_4 FILLER_68_657 ();
 sg13g2_fill_2 FILLER_68_661 ();
 sg13g2_fill_1 FILLER_68_666 ();
 sg13g2_fill_1 FILLER_68_671 ();
 sg13g2_fill_1 FILLER_68_701 ();
 sg13g2_decap_8 FILLER_68_706 ();
 sg13g2_decap_4 FILLER_68_713 ();
 sg13g2_fill_2 FILLER_68_717 ();
 sg13g2_decap_8 FILLER_68_724 ();
 sg13g2_decap_8 FILLER_68_731 ();
 sg13g2_fill_1 FILLER_68_738 ();
 sg13g2_decap_4 FILLER_68_753 ();
 sg13g2_fill_1 FILLER_68_765 ();
 sg13g2_fill_1 FILLER_68_771 ();
 sg13g2_decap_4 FILLER_68_794 ();
 sg13g2_fill_1 FILLER_68_798 ();
 sg13g2_fill_1 FILLER_68_813 ();
 sg13g2_fill_2 FILLER_68_831 ();
 sg13g2_fill_1 FILLER_68_833 ();
 sg13g2_decap_8 FILLER_68_847 ();
 sg13g2_fill_2 FILLER_68_854 ();
 sg13g2_decap_4 FILLER_68_865 ();
 sg13g2_decap_4 FILLER_68_872 ();
 sg13g2_fill_1 FILLER_68_876 ();
 sg13g2_decap_4 FILLER_68_881 ();
 sg13g2_fill_2 FILLER_68_885 ();
 sg13g2_fill_1 FILLER_68_900 ();
 sg13g2_fill_2 FILLER_68_905 ();
 sg13g2_fill_2 FILLER_68_911 ();
 sg13g2_decap_4 FILLER_68_918 ();
 sg13g2_fill_2 FILLER_68_935 ();
 sg13g2_fill_1 FILLER_68_937 ();
 sg13g2_decap_8 FILLER_68_942 ();
 sg13g2_fill_2 FILLER_68_949 ();
 sg13g2_fill_1 FILLER_68_951 ();
 sg13g2_decap_8 FILLER_68_965 ();
 sg13g2_fill_1 FILLER_68_972 ();
 sg13g2_fill_2 FILLER_68_977 ();
 sg13g2_decap_8 FILLER_68_988 ();
 sg13g2_fill_2 FILLER_68_995 ();
 sg13g2_fill_1 FILLER_68_1010 ();
 sg13g2_decap_4 FILLER_68_1034 ();
 sg13g2_fill_1 FILLER_68_1038 ();
 sg13g2_fill_1 FILLER_68_1065 ();
 sg13g2_fill_2 FILLER_68_1072 ();
 sg13g2_fill_1 FILLER_68_1100 ();
 sg13g2_fill_2 FILLER_68_1132 ();
 sg13g2_fill_1 FILLER_68_1134 ();
 sg13g2_fill_2 FILLER_68_1174 ();
 sg13g2_fill_1 FILLER_68_1180 ();
 sg13g2_fill_1 FILLER_68_1185 ();
 sg13g2_decap_8 FILLER_68_1216 ();
 sg13g2_fill_1 FILLER_68_1223 ();
 sg13g2_fill_1 FILLER_68_1241 ();
 sg13g2_fill_1 FILLER_68_1247 ();
 sg13g2_fill_2 FILLER_68_1252 ();
 sg13g2_fill_1 FILLER_68_1264 ();
 sg13g2_fill_2 FILLER_68_1274 ();
 sg13g2_decap_4 FILLER_68_1281 ();
 sg13g2_fill_1 FILLER_68_1289 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_11 ();
 sg13g2_fill_1 FILLER_69_18 ();
 sg13g2_fill_1 FILLER_69_45 ();
 sg13g2_fill_1 FILLER_69_55 ();
 sg13g2_fill_2 FILLER_69_60 ();
 sg13g2_decap_4 FILLER_69_70 ();
 sg13g2_fill_1 FILLER_69_74 ();
 sg13g2_fill_2 FILLER_69_80 ();
 sg13g2_decap_8 FILLER_69_86 ();
 sg13g2_decap_8 FILLER_69_103 ();
 sg13g2_decap_8 FILLER_69_110 ();
 sg13g2_decap_8 FILLER_69_117 ();
 sg13g2_decap_8 FILLER_69_124 ();
 sg13g2_fill_2 FILLER_69_131 ();
 sg13g2_fill_1 FILLER_69_133 ();
 sg13g2_fill_2 FILLER_69_139 ();
 sg13g2_fill_1 FILLER_69_141 ();
 sg13g2_decap_4 FILLER_69_157 ();
 sg13g2_decap_8 FILLER_69_165 ();
 sg13g2_decap_4 FILLER_69_172 ();
 sg13g2_fill_2 FILLER_69_176 ();
 sg13g2_fill_2 FILLER_69_187 ();
 sg13g2_fill_1 FILLER_69_192 ();
 sg13g2_fill_1 FILLER_69_197 ();
 sg13g2_fill_1 FILLER_69_203 ();
 sg13g2_fill_1 FILLER_69_223 ();
 sg13g2_fill_1 FILLER_69_228 ();
 sg13g2_fill_1 FILLER_69_234 ();
 sg13g2_fill_1 FILLER_69_239 ();
 sg13g2_decap_4 FILLER_69_244 ();
 sg13g2_fill_1 FILLER_69_248 ();
 sg13g2_fill_2 FILLER_69_271 ();
 sg13g2_fill_2 FILLER_69_320 ();
 sg13g2_decap_8 FILLER_69_327 ();
 sg13g2_decap_4 FILLER_69_334 ();
 sg13g2_fill_2 FILLER_69_338 ();
 sg13g2_decap_4 FILLER_69_345 ();
 sg13g2_fill_1 FILLER_69_349 ();
 sg13g2_decap_8 FILLER_69_354 ();
 sg13g2_decap_4 FILLER_69_361 ();
 sg13g2_fill_2 FILLER_69_365 ();
 sg13g2_decap_4 FILLER_69_402 ();
 sg13g2_fill_1 FILLER_69_414 ();
 sg13g2_fill_2 FILLER_69_418 ();
 sg13g2_fill_1 FILLER_69_425 ();
 sg13g2_fill_1 FILLER_69_430 ();
 sg13g2_decap_8 FILLER_69_444 ();
 sg13g2_decap_8 FILLER_69_455 ();
 sg13g2_fill_1 FILLER_69_462 ();
 sg13g2_fill_2 FILLER_69_473 ();
 sg13g2_fill_1 FILLER_69_478 ();
 sg13g2_fill_1 FILLER_69_482 ();
 sg13g2_fill_1 FILLER_69_488 ();
 sg13g2_fill_1 FILLER_69_493 ();
 sg13g2_fill_2 FILLER_69_498 ();
 sg13g2_decap_8 FILLER_69_504 ();
 sg13g2_decap_4 FILLER_69_511 ();
 sg13g2_fill_2 FILLER_69_523 ();
 sg13g2_fill_1 FILLER_69_525 ();
 sg13g2_decap_8 FILLER_69_530 ();
 sg13g2_decap_8 FILLER_69_537 ();
 sg13g2_fill_2 FILLER_69_544 ();
 sg13g2_fill_2 FILLER_69_551 ();
 sg13g2_fill_1 FILLER_69_558 ();
 sg13g2_fill_2 FILLER_69_594 ();
 sg13g2_fill_1 FILLER_69_638 ();
 sg13g2_decap_4 FILLER_69_670 ();
 sg13g2_decap_8 FILLER_69_678 ();
 sg13g2_fill_1 FILLER_69_768 ();
 sg13g2_decap_8 FILLER_69_778 ();
 sg13g2_fill_1 FILLER_69_800 ();
 sg13g2_decap_4 FILLER_69_807 ();
 sg13g2_fill_2 FILLER_69_811 ();
 sg13g2_decap_8 FILLER_69_821 ();
 sg13g2_fill_1 FILLER_69_828 ();
 sg13g2_fill_2 FILLER_69_847 ();
 sg13g2_fill_1 FILLER_69_849 ();
 sg13g2_fill_1 FILLER_69_930 ();
 sg13g2_fill_2 FILLER_69_957 ();
 sg13g2_fill_2 FILLER_69_963 ();
 sg13g2_fill_2 FILLER_69_979 ();
 sg13g2_fill_1 FILLER_69_995 ();
 sg13g2_fill_1 FILLER_69_1005 ();
 sg13g2_decap_8 FILLER_69_1017 ();
 sg13g2_fill_1 FILLER_69_1024 ();
 sg13g2_decap_8 FILLER_69_1029 ();
 sg13g2_decap_8 FILLER_69_1036 ();
 sg13g2_fill_2 FILLER_69_1043 ();
 sg13g2_fill_1 FILLER_69_1045 ();
 sg13g2_fill_1 FILLER_69_1050 ();
 sg13g2_fill_1 FILLER_69_1055 ();
 sg13g2_fill_1 FILLER_69_1060 ();
 sg13g2_fill_1 FILLER_69_1065 ();
 sg13g2_decap_4 FILLER_69_1070 ();
 sg13g2_decap_4 FILLER_69_1087 ();
 sg13g2_decap_8 FILLER_69_1108 ();
 sg13g2_fill_2 FILLER_69_1115 ();
 sg13g2_fill_2 FILLER_69_1122 ();
 sg13g2_fill_1 FILLER_69_1124 ();
 sg13g2_fill_1 FILLER_69_1130 ();
 sg13g2_fill_2 FILLER_69_1137 ();
 sg13g2_fill_2 FILLER_69_1142 ();
 sg13g2_fill_2 FILLER_69_1149 ();
 sg13g2_decap_8 FILLER_69_1155 ();
 sg13g2_decap_4 FILLER_69_1162 ();
 sg13g2_fill_2 FILLER_69_1166 ();
 sg13g2_fill_1 FILLER_69_1177 ();
 sg13g2_fill_2 FILLER_69_1182 ();
 sg13g2_fill_1 FILLER_69_1188 ();
 sg13g2_decap_8 FILLER_69_1198 ();
 sg13g2_decap_8 FILLER_69_1205 ();
 sg13g2_decap_8 FILLER_69_1212 ();
 sg13g2_fill_2 FILLER_69_1219 ();
 sg13g2_fill_2 FILLER_69_1247 ();
 sg13g2_decap_8 FILLER_69_1292 ();
 sg13g2_decap_8 FILLER_69_1299 ();
 sg13g2_fill_1 FILLER_69_1310 ();
 sg13g2_decap_8 FILLER_69_1315 ();
 sg13g2_decap_4 FILLER_69_1322 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_7 ();
 sg13g2_fill_2 FILLER_70_11 ();
 sg13g2_fill_2 FILLER_70_39 ();
 sg13g2_fill_2 FILLER_70_46 ();
 sg13g2_decap_8 FILLER_70_55 ();
 sg13g2_decap_4 FILLER_70_62 ();
 sg13g2_fill_2 FILLER_70_66 ();
 sg13g2_decap_4 FILLER_70_72 ();
 sg13g2_fill_1 FILLER_70_76 ();
 sg13g2_fill_2 FILLER_70_86 ();
 sg13g2_fill_2 FILLER_70_92 ();
 sg13g2_fill_1 FILLER_70_94 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_4 FILLER_70_140 ();
 sg13g2_fill_2 FILLER_70_144 ();
 sg13g2_fill_2 FILLER_70_160 ();
 sg13g2_decap_4 FILLER_70_171 ();
 sg13g2_fill_1 FILLER_70_175 ();
 sg13g2_fill_1 FILLER_70_190 ();
 sg13g2_fill_2 FILLER_70_203 ();
 sg13g2_fill_1 FILLER_70_205 ();
 sg13g2_decap_8 FILLER_70_215 ();
 sg13g2_fill_2 FILLER_70_222 ();
 sg13g2_fill_1 FILLER_70_224 ();
 sg13g2_fill_1 FILLER_70_236 ();
 sg13g2_fill_1 FILLER_70_241 ();
 sg13g2_decap_8 FILLER_70_247 ();
 sg13g2_fill_1 FILLER_70_258 ();
 sg13g2_fill_2 FILLER_70_278 ();
 sg13g2_fill_1 FILLER_70_280 ();
 sg13g2_fill_1 FILLER_70_285 ();
 sg13g2_decap_8 FILLER_70_290 ();
 sg13g2_fill_1 FILLER_70_297 ();
 sg13g2_decap_8 FILLER_70_305 ();
 sg13g2_decap_4 FILLER_70_312 ();
 sg13g2_fill_2 FILLER_70_350 ();
 sg13g2_decap_4 FILLER_70_357 ();
 sg13g2_fill_2 FILLER_70_365 ();
 sg13g2_decap_4 FILLER_70_375 ();
 sg13g2_fill_2 FILLER_70_379 ();
 sg13g2_fill_2 FILLER_70_419 ();
 sg13g2_fill_2 FILLER_70_429 ();
 sg13g2_decap_4 FILLER_70_435 ();
 sg13g2_fill_1 FILLER_70_439 ();
 sg13g2_fill_1 FILLER_70_445 ();
 sg13g2_fill_1 FILLER_70_449 ();
 sg13g2_fill_2 FILLER_70_458 ();
 sg13g2_fill_1 FILLER_70_473 ();
 sg13g2_fill_2 FILLER_70_517 ();
 sg13g2_fill_1 FILLER_70_606 ();
 sg13g2_decap_8 FILLER_70_611 ();
 sg13g2_decap_8 FILLER_70_618 ();
 sg13g2_decap_8 FILLER_70_625 ();
 sg13g2_decap_8 FILLER_70_641 ();
 sg13g2_fill_2 FILLER_70_648 ();
 sg13g2_decap_8 FILLER_70_654 ();
 sg13g2_decap_8 FILLER_70_661 ();
 sg13g2_decap_8 FILLER_70_668 ();
 sg13g2_decap_8 FILLER_70_675 ();
 sg13g2_decap_4 FILLER_70_682 ();
 sg13g2_decap_4 FILLER_70_718 ();
 sg13g2_decap_8 FILLER_70_726 ();
 sg13g2_decap_4 FILLER_70_733 ();
 sg13g2_fill_1 FILLER_70_737 ();
 sg13g2_decap_4 FILLER_70_741 ();
 sg13g2_decap_4 FILLER_70_754 ();
 sg13g2_fill_2 FILLER_70_758 ();
 sg13g2_decap_8 FILLER_70_767 ();
 sg13g2_decap_4 FILLER_70_774 ();
 sg13g2_fill_2 FILLER_70_778 ();
 sg13g2_fill_1 FILLER_70_786 ();
 sg13g2_fill_1 FILLER_70_814 ();
 sg13g2_fill_2 FILLER_70_823 ();
 sg13g2_fill_1 FILLER_70_825 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_fill_2 FILLER_70_847 ();
 sg13g2_decap_4 FILLER_70_852 ();
 sg13g2_fill_2 FILLER_70_885 ();
 sg13g2_decap_8 FILLER_70_913 ();
 sg13g2_fill_2 FILLER_70_920 ();
 sg13g2_fill_1 FILLER_70_955 ();
 sg13g2_decap_4 FILLER_70_964 ();
 sg13g2_fill_2 FILLER_70_977 ();
 sg13g2_fill_2 FILLER_70_994 ();
 sg13g2_fill_1 FILLER_70_996 ();
 sg13g2_fill_2 FILLER_70_1007 ();
 sg13g2_fill_2 FILLER_70_1049 ();
 sg13g2_fill_2 FILLER_70_1056 ();
 sg13g2_fill_1 FILLER_70_1071 ();
 sg13g2_decap_8 FILLER_70_1076 ();
 sg13g2_fill_1 FILLER_70_1083 ();
 sg13g2_fill_1 FILLER_70_1088 ();
 sg13g2_fill_1 FILLER_70_1115 ();
 sg13g2_fill_1 FILLER_70_1142 ();
 sg13g2_fill_1 FILLER_70_1195 ();
 sg13g2_fill_2 FILLER_70_1222 ();
 sg13g2_fill_1 FILLER_70_1224 ();
 sg13g2_decap_4 FILLER_70_1234 ();
 sg13g2_fill_1 FILLER_70_1246 ();
 sg13g2_fill_2 FILLER_70_1255 ();
 sg13g2_fill_1 FILLER_70_1257 ();
 sg13g2_decap_8 FILLER_70_1262 ();
 sg13g2_fill_1 FILLER_70_1269 ();
 sg13g2_fill_2 FILLER_70_1274 ();
 sg13g2_fill_1 FILLER_70_1276 ();
 sg13g2_decap_4 FILLER_70_1287 ();
 sg13g2_fill_1 FILLER_70_1291 ();
 sg13g2_fill_2 FILLER_70_1297 ();
 sg13g2_fill_1 FILLER_70_1325 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_fill_1 FILLER_71_21 ();
 sg13g2_fill_1 FILLER_71_26 ();
 sg13g2_fill_2 FILLER_71_52 ();
 sg13g2_fill_1 FILLER_71_66 ();
 sg13g2_decap_8 FILLER_71_72 ();
 sg13g2_fill_2 FILLER_71_79 ();
 sg13g2_fill_1 FILLER_71_81 ();
 sg13g2_fill_1 FILLER_71_85 ();
 sg13g2_fill_1 FILLER_71_103 ();
 sg13g2_fill_2 FILLER_71_117 ();
 sg13g2_decap_8 FILLER_71_124 ();
 sg13g2_decap_4 FILLER_71_131 ();
 sg13g2_fill_1 FILLER_71_148 ();
 sg13g2_fill_2 FILLER_71_157 ();
 sg13g2_fill_2 FILLER_71_179 ();
 sg13g2_fill_1 FILLER_71_181 ();
 sg13g2_decap_8 FILLER_71_190 ();
 sg13g2_fill_2 FILLER_71_197 ();
 sg13g2_fill_2 FILLER_71_214 ();
 sg13g2_fill_1 FILLER_71_224 ();
 sg13g2_fill_1 FILLER_71_230 ();
 sg13g2_fill_2 FILLER_71_236 ();
 sg13g2_fill_1 FILLER_71_266 ();
 sg13g2_decap_4 FILLER_71_277 ();
 sg13g2_fill_1 FILLER_71_290 ();
 sg13g2_fill_1 FILLER_71_317 ();
 sg13g2_fill_1 FILLER_71_323 ();
 sg13g2_fill_1 FILLER_71_328 ();
 sg13g2_fill_1 FILLER_71_333 ();
 sg13g2_fill_1 FILLER_71_389 ();
 sg13g2_fill_2 FILLER_71_408 ();
 sg13g2_fill_1 FILLER_71_410 ();
 sg13g2_fill_1 FILLER_71_456 ();
 sg13g2_fill_2 FILLER_71_462 ();
 sg13g2_fill_1 FILLER_71_469 ();
 sg13g2_fill_1 FILLER_71_475 ();
 sg13g2_fill_1 FILLER_71_495 ();
 sg13g2_decap_8 FILLER_71_500 ();
 sg13g2_fill_1 FILLER_71_507 ();
 sg13g2_decap_8 FILLER_71_512 ();
 sg13g2_decap_8 FILLER_71_519 ();
 sg13g2_decap_8 FILLER_71_526 ();
 sg13g2_fill_2 FILLER_71_533 ();
 sg13g2_fill_1 FILLER_71_535 ();
 sg13g2_fill_2 FILLER_71_541 ();
 sg13g2_fill_1 FILLER_71_543 ();
 sg13g2_decap_8 FILLER_71_558 ();
 sg13g2_fill_2 FILLER_71_565 ();
 sg13g2_fill_1 FILLER_71_567 ();
 sg13g2_decap_8 FILLER_71_575 ();
 sg13g2_fill_1 FILLER_71_627 ();
 sg13g2_fill_2 FILLER_71_635 ();
 sg13g2_fill_1 FILLER_71_672 ();
 sg13g2_fill_1 FILLER_71_678 ();
 sg13g2_fill_2 FILLER_71_684 ();
 sg13g2_fill_2 FILLER_71_689 ();
 sg13g2_decap_8 FILLER_71_715 ();
 sg13g2_decap_8 FILLER_71_722 ();
 sg13g2_decap_8 FILLER_71_734 ();
 sg13g2_fill_1 FILLER_71_741 ();
 sg13g2_fill_2 FILLER_71_747 ();
 sg13g2_fill_1 FILLER_71_785 ();
 sg13g2_fill_1 FILLER_71_789 ();
 sg13g2_fill_2 FILLER_71_795 ();
 sg13g2_fill_1 FILLER_71_802 ();
 sg13g2_fill_2 FILLER_71_811 ();
 sg13g2_fill_1 FILLER_71_827 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_decap_4 FILLER_71_867 ();
 sg13g2_fill_2 FILLER_71_871 ();
 sg13g2_decap_8 FILLER_71_883 ();
 sg13g2_decap_4 FILLER_71_899 ();
 sg13g2_fill_1 FILLER_71_939 ();
 sg13g2_fill_2 FILLER_71_948 ();
 sg13g2_fill_1 FILLER_71_950 ();
 sg13g2_decap_8 FILLER_71_956 ();
 sg13g2_fill_2 FILLER_71_963 ();
 sg13g2_decap_8 FILLER_71_974 ();
 sg13g2_decap_4 FILLER_71_981 ();
 sg13g2_fill_1 FILLER_71_985 ();
 sg13g2_decap_8 FILLER_71_991 ();
 sg13g2_fill_2 FILLER_71_1003 ();
 sg13g2_decap_4 FILLER_71_1021 ();
 sg13g2_fill_1 FILLER_71_1025 ();
 sg13g2_decap_8 FILLER_71_1031 ();
 sg13g2_decap_8 FILLER_71_1048 ();
 sg13g2_fill_2 FILLER_71_1055 ();
 sg13g2_fill_1 FILLER_71_1057 ();
 sg13g2_decap_8 FILLER_71_1095 ();
 sg13g2_fill_1 FILLER_71_1102 ();
 sg13g2_fill_1 FILLER_71_1115 ();
 sg13g2_fill_2 FILLER_71_1120 ();
 sg13g2_fill_2 FILLER_71_1126 ();
 sg13g2_fill_2 FILLER_71_1137 ();
 sg13g2_fill_1 FILLER_71_1139 ();
 sg13g2_decap_4 FILLER_71_1146 ();
 sg13g2_decap_8 FILLER_71_1154 ();
 sg13g2_fill_2 FILLER_71_1161 ();
 sg13g2_decap_8 FILLER_71_1166 ();
 sg13g2_decap_8 FILLER_71_1173 ();
 sg13g2_fill_2 FILLER_71_1180 ();
 sg13g2_fill_2 FILLER_71_1198 ();
 sg13g2_fill_1 FILLER_71_1200 ();
 sg13g2_fill_2 FILLER_71_1205 ();
 sg13g2_decap_8 FILLER_71_1211 ();
 sg13g2_fill_2 FILLER_71_1218 ();
 sg13g2_fill_1 FILLER_71_1220 ();
 sg13g2_fill_1 FILLER_71_1247 ();
 sg13g2_fill_2 FILLER_71_1253 ();
 sg13g2_decap_4 FILLER_71_1262 ();
 sg13g2_fill_1 FILLER_71_1266 ();
 sg13g2_decap_4 FILLER_71_1271 ();
 sg13g2_decap_4 FILLER_71_1284 ();
 sg13g2_fill_1 FILLER_71_1288 ();
 sg13g2_fill_2 FILLER_71_1323 ();
 sg13g2_fill_1 FILLER_71_1325 ();
 sg13g2_decap_4 FILLER_72_26 ();
 sg13g2_fill_1 FILLER_72_30 ();
 sg13g2_fill_2 FILLER_72_40 ();
 sg13g2_decap_4 FILLER_72_50 ();
 sg13g2_decap_8 FILLER_72_58 ();
 sg13g2_fill_2 FILLER_72_65 ();
 sg13g2_fill_1 FILLER_72_72 ();
 sg13g2_fill_1 FILLER_72_78 ();
 sg13g2_fill_2 FILLER_72_101 ();
 sg13g2_decap_8 FILLER_72_107 ();
 sg13g2_decap_4 FILLER_72_114 ();
 sg13g2_fill_1 FILLER_72_118 ();
 sg13g2_decap_8 FILLER_72_124 ();
 sg13g2_decap_8 FILLER_72_131 ();
 sg13g2_fill_1 FILLER_72_138 ();
 sg13g2_fill_2 FILLER_72_160 ();
 sg13g2_fill_1 FILLER_72_167 ();
 sg13g2_fill_2 FILLER_72_175 ();
 sg13g2_decap_4 FILLER_72_185 ();
 sg13g2_fill_1 FILLER_72_189 ();
 sg13g2_decap_4 FILLER_72_193 ();
 sg13g2_fill_1 FILLER_72_197 ();
 sg13g2_decap_4 FILLER_72_204 ();
 sg13g2_fill_2 FILLER_72_212 ();
 sg13g2_fill_1 FILLER_72_231 ();
 sg13g2_fill_2 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_254 ();
 sg13g2_decap_8 FILLER_72_261 ();
 sg13g2_fill_2 FILLER_72_296 ();
 sg13g2_fill_1 FILLER_72_318 ();
 sg13g2_fill_1 FILLER_72_345 ();
 sg13g2_fill_2 FILLER_72_349 ();
 sg13g2_decap_4 FILLER_72_355 ();
 sg13g2_fill_1 FILLER_72_371 ();
 sg13g2_fill_1 FILLER_72_402 ();
 sg13g2_decap_8 FILLER_72_412 ();
 sg13g2_decap_8 FILLER_72_419 ();
 sg13g2_fill_1 FILLER_72_426 ();
 sg13g2_fill_2 FILLER_72_432 ();
 sg13g2_fill_2 FILLER_72_451 ();
 sg13g2_decap_8 FILLER_72_468 ();
 sg13g2_fill_2 FILLER_72_475 ();
 sg13g2_fill_2 FILLER_72_484 ();
 sg13g2_fill_1 FILLER_72_494 ();
 sg13g2_fill_2 FILLER_72_498 ();
 sg13g2_decap_4 FILLER_72_530 ();
 sg13g2_fill_2 FILLER_72_534 ();
 sg13g2_fill_2 FILLER_72_560 ();
 sg13g2_fill_1 FILLER_72_562 ();
 sg13g2_fill_1 FILLER_72_581 ();
 sg13g2_fill_2 FILLER_72_605 ();
 sg13g2_decap_8 FILLER_72_611 ();
 sg13g2_decap_8 FILLER_72_618 ();
 sg13g2_decap_4 FILLER_72_633 ();
 sg13g2_fill_2 FILLER_72_637 ();
 sg13g2_decap_4 FILLER_72_648 ();
 sg13g2_fill_2 FILLER_72_652 ();
 sg13g2_fill_2 FILLER_72_657 ();
 sg13g2_decap_4 FILLER_72_665 ();
 sg13g2_fill_1 FILLER_72_678 ();
 sg13g2_fill_2 FILLER_72_690 ();
 sg13g2_fill_1 FILLER_72_692 ();
 sg13g2_fill_2 FILLER_72_697 ();
 sg13g2_fill_2 FILLER_72_702 ();
 sg13g2_fill_2 FILLER_72_744 ();
 sg13g2_decap_8 FILLER_72_768 ();
 sg13g2_decap_4 FILLER_72_779 ();
 sg13g2_decap_8 FILLER_72_788 ();
 sg13g2_decap_4 FILLER_72_799 ();
 sg13g2_fill_1 FILLER_72_803 ();
 sg13g2_fill_2 FILLER_72_809 ();
 sg13g2_fill_2 FILLER_72_816 ();
 sg13g2_fill_1 FILLER_72_824 ();
 sg13g2_fill_1 FILLER_72_834 ();
 sg13g2_fill_2 FILLER_72_840 ();
 sg13g2_fill_2 FILLER_72_852 ();
 sg13g2_decap_8 FILLER_72_878 ();
 sg13g2_decap_8 FILLER_72_885 ();
 sg13g2_fill_2 FILLER_72_906 ();
 sg13g2_fill_1 FILLER_72_908 ();
 sg13g2_fill_2 FILLER_72_921 ();
 sg13g2_fill_1 FILLER_72_926 ();
 sg13g2_fill_1 FILLER_72_931 ();
 sg13g2_fill_2 FILLER_72_951 ();
 sg13g2_fill_1 FILLER_72_953 ();
 sg13g2_fill_1 FILLER_72_959 ();
 sg13g2_fill_1 FILLER_72_965 ();
 sg13g2_fill_1 FILLER_72_984 ();
 sg13g2_fill_1 FILLER_72_989 ();
 sg13g2_fill_1 FILLER_72_996 ();
 sg13g2_fill_2 FILLER_72_1002 ();
 sg13g2_fill_1 FILLER_72_1017 ();
 sg13g2_decap_4 FILLER_72_1040 ();
 sg13g2_fill_2 FILLER_72_1071 ();
 sg13g2_fill_1 FILLER_72_1073 ();
 sg13g2_decap_8 FILLER_72_1079 ();
 sg13g2_fill_2 FILLER_72_1086 ();
 sg13g2_fill_1 FILLER_72_1088 ();
 sg13g2_decap_8 FILLER_72_1095 ();
 sg13g2_fill_2 FILLER_72_1102 ();
 sg13g2_fill_2 FILLER_72_1109 ();
 sg13g2_decap_4 FILLER_72_1149 ();
 sg13g2_fill_1 FILLER_72_1153 ();
 sg13g2_fill_1 FILLER_72_1159 ();
 sg13g2_decap_8 FILLER_72_1170 ();
 sg13g2_decap_8 FILLER_72_1177 ();
 sg13g2_fill_1 FILLER_72_1184 ();
 sg13g2_fill_2 FILLER_72_1220 ();
 sg13g2_fill_1 FILLER_72_1222 ();
 sg13g2_fill_2 FILLER_72_1231 ();
 sg13g2_fill_1 FILLER_72_1241 ();
 sg13g2_decap_4 FILLER_72_1277 ();
 sg13g2_fill_2 FILLER_72_1284 ();
 sg13g2_fill_1 FILLER_72_1286 ();
 sg13g2_fill_1 FILLER_72_1291 ();
 sg13g2_decap_8 FILLER_72_1305 ();
 sg13g2_decap_8 FILLER_72_1312 ();
 sg13g2_decap_8 FILLER_72_1319 ();
 sg13g2_decap_4 FILLER_73_0 ();
 sg13g2_decap_4 FILLER_73_34 ();
 sg13g2_fill_2 FILLER_73_38 ();
 sg13g2_fill_2 FILLER_73_49 ();
 sg13g2_fill_2 FILLER_73_59 ();
 sg13g2_fill_1 FILLER_73_61 ();
 sg13g2_fill_1 FILLER_73_70 ();
 sg13g2_fill_2 FILLER_73_88 ();
 sg13g2_fill_2 FILLER_73_99 ();
 sg13g2_fill_2 FILLER_73_105 ();
 sg13g2_fill_1 FILLER_73_107 ();
 sg13g2_decap_4 FILLER_73_134 ();
 sg13g2_fill_1 FILLER_73_155 ();
 sg13g2_fill_2 FILLER_73_183 ();
 sg13g2_fill_1 FILLER_73_189 ();
 sg13g2_fill_2 FILLER_73_208 ();
 sg13g2_fill_1 FILLER_73_210 ();
 sg13g2_fill_1 FILLER_73_220 ();
 sg13g2_fill_1 FILLER_73_229 ();
 sg13g2_fill_1 FILLER_73_235 ();
 sg13g2_fill_1 FILLER_73_245 ();
 sg13g2_decap_8 FILLER_73_250 ();
 sg13g2_fill_1 FILLER_73_257 ();
 sg13g2_fill_2 FILLER_73_264 ();
 sg13g2_fill_1 FILLER_73_266 ();
 sg13g2_decap_4 FILLER_73_271 ();
 sg13g2_fill_1 FILLER_73_275 ();
 sg13g2_fill_1 FILLER_73_319 ();
 sg13g2_fill_1 FILLER_73_324 ();
 sg13g2_fill_1 FILLER_73_329 ();
 sg13g2_fill_1 FILLER_73_334 ();
 sg13g2_fill_2 FILLER_73_345 ();
 sg13g2_decap_8 FILLER_73_360 ();
 sg13g2_fill_1 FILLER_73_367 ();
 sg13g2_fill_1 FILLER_73_381 ();
 sg13g2_decap_8 FILLER_73_386 ();
 sg13g2_decap_8 FILLER_73_393 ();
 sg13g2_decap_8 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_fill_1 FILLER_73_441 ();
 sg13g2_decap_8 FILLER_73_455 ();
 sg13g2_decap_8 FILLER_73_462 ();
 sg13g2_decap_4 FILLER_73_469 ();
 sg13g2_fill_1 FILLER_73_478 ();
 sg13g2_fill_2 FILLER_73_492 ();
 sg13g2_decap_8 FILLER_73_498 ();
 sg13g2_fill_2 FILLER_73_505 ();
 sg13g2_fill_2 FILLER_73_512 ();
 sg13g2_fill_1 FILLER_73_545 ();
 sg13g2_decap_4 FILLER_73_556 ();
 sg13g2_fill_1 FILLER_73_560 ();
 sg13g2_decap_8 FILLER_73_570 ();
 sg13g2_fill_1 FILLER_73_590 ();
 sg13g2_decap_4 FILLER_73_594 ();
 sg13g2_fill_2 FILLER_73_598 ();
 sg13g2_fill_2 FILLER_73_626 ();
 sg13g2_fill_1 FILLER_73_628 ();
 sg13g2_decap_4 FILLER_73_634 ();
 sg13g2_fill_1 FILLER_73_638 ();
 sg13g2_decap_4 FILLER_73_644 ();
 sg13g2_fill_1 FILLER_73_658 ();
 sg13g2_fill_2 FILLER_73_664 ();
 sg13g2_fill_1 FILLER_73_666 ();
 sg13g2_decap_4 FILLER_73_678 ();
 sg13g2_fill_1 FILLER_73_685 ();
 sg13g2_fill_1 FILLER_73_690 ();
 sg13g2_fill_2 FILLER_73_695 ();
 sg13g2_fill_1 FILLER_73_702 ();
 sg13g2_fill_1 FILLER_73_708 ();
 sg13g2_fill_2 FILLER_73_714 ();
 sg13g2_decap_8 FILLER_73_720 ();
 sg13g2_fill_2 FILLER_73_727 ();
 sg13g2_fill_2 FILLER_73_742 ();
 sg13g2_fill_2 FILLER_73_753 ();
 sg13g2_fill_1 FILLER_73_794 ();
 sg13g2_fill_1 FILLER_73_803 ();
 sg13g2_decap_4 FILLER_73_812 ();
 sg13g2_fill_2 FILLER_73_816 ();
 sg13g2_fill_2 FILLER_73_822 ();
 sg13g2_fill_1 FILLER_73_824 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_73_915 ();
 sg13g2_decap_8 FILLER_73_929 ();
 sg13g2_fill_1 FILLER_73_936 ();
 sg13g2_fill_1 FILLER_73_943 ();
 sg13g2_fill_1 FILLER_73_950 ();
 sg13g2_fill_1 FILLER_73_955 ();
 sg13g2_decap_4 FILLER_73_961 ();
 sg13g2_fill_2 FILLER_73_965 ();
 sg13g2_fill_2 FILLER_73_972 ();
 sg13g2_fill_1 FILLER_73_974 ();
 sg13g2_decap_4 FILLER_73_979 ();
 sg13g2_fill_2 FILLER_73_983 ();
 sg13g2_decap_8 FILLER_73_990 ();
 sg13g2_fill_2 FILLER_73_997 ();
 sg13g2_decap_8 FILLER_73_1009 ();
 sg13g2_decap_4 FILLER_73_1016 ();
 sg13g2_fill_1 FILLER_73_1024 ();
 sg13g2_decap_8 FILLER_73_1029 ();
 sg13g2_decap_8 FILLER_73_1036 ();
 sg13g2_decap_4 FILLER_73_1055 ();
 sg13g2_fill_2 FILLER_73_1059 ();
 sg13g2_fill_1 FILLER_73_1069 ();
 sg13g2_decap_4 FILLER_73_1075 ();
 sg13g2_decap_8 FILLER_73_1118 ();
 sg13g2_fill_2 FILLER_73_1129 ();
 sg13g2_fill_1 FILLER_73_1131 ();
 sg13g2_decap_8 FILLER_73_1136 ();
 sg13g2_fill_1 FILLER_73_1143 ();
 sg13g2_fill_1 FILLER_73_1178 ();
 sg13g2_decap_4 FILLER_73_1193 ();
 sg13g2_decap_8 FILLER_73_1223 ();
 sg13g2_fill_1 FILLER_73_1230 ();
 sg13g2_decap_8 FILLER_73_1236 ();
 sg13g2_decap_4 FILLER_73_1243 ();
 sg13g2_fill_2 FILLER_73_1247 ();
 sg13g2_fill_1 FILLER_73_1252 ();
 sg13g2_decap_8 FILLER_73_1257 ();
 sg13g2_fill_2 FILLER_73_1264 ();
 sg13g2_fill_1 FILLER_73_1266 ();
 sg13g2_fill_1 FILLER_73_1298 ();
 sg13g2_fill_1 FILLER_73_1303 ();
 sg13g2_decap_8 FILLER_73_1307 ();
 sg13g2_decap_8 FILLER_73_1314 ();
 sg13g2_decap_4 FILLER_73_1321 ();
 sg13g2_fill_1 FILLER_73_1325 ();
 sg13g2_fill_1 FILLER_74_4 ();
 sg13g2_fill_1 FILLER_74_44 ();
 sg13g2_fill_1 FILLER_74_49 ();
 sg13g2_decap_4 FILLER_74_96 ();
 sg13g2_fill_1 FILLER_74_100 ();
 sg13g2_fill_2 FILLER_74_105 ();
 sg13g2_fill_1 FILLER_74_107 ();
 sg13g2_fill_2 FILLER_74_134 ();
 sg13g2_fill_2 FILLER_74_146 ();
 sg13g2_fill_2 FILLER_74_161 ();
 sg13g2_fill_1 FILLER_74_163 ();
 sg13g2_fill_2 FILLER_74_175 ();
 sg13g2_fill_2 FILLER_74_191 ();
 sg13g2_decap_8 FILLER_74_205 ();
 sg13g2_decap_8 FILLER_74_216 ();
 sg13g2_fill_2 FILLER_74_223 ();
 sg13g2_fill_1 FILLER_74_225 ();
 sg13g2_decap_4 FILLER_74_231 ();
 sg13g2_fill_2 FILLER_74_267 ();
 sg13g2_decap_8 FILLER_74_273 ();
 sg13g2_fill_1 FILLER_74_280 ();
 sg13g2_fill_2 FILLER_74_286 ();
 sg13g2_fill_1 FILLER_74_295 ();
 sg13g2_decap_4 FILLER_74_300 ();
 sg13g2_fill_2 FILLER_74_304 ();
 sg13g2_decap_8 FILLER_74_310 ();
 sg13g2_fill_2 FILLER_74_317 ();
 sg13g2_fill_1 FILLER_74_319 ();
 sg13g2_decap_8 FILLER_74_324 ();
 sg13g2_decap_4 FILLER_74_331 ();
 sg13g2_fill_2 FILLER_74_335 ();
 sg13g2_fill_2 FILLER_74_377 ();
 sg13g2_fill_1 FILLER_74_379 ();
 sg13g2_decap_8 FILLER_74_423 ();
 sg13g2_fill_1 FILLER_74_445 ();
 sg13g2_decap_4 FILLER_74_450 ();
 sg13g2_decap_4 FILLER_74_458 ();
 sg13g2_fill_2 FILLER_74_467 ();
 sg13g2_fill_1 FILLER_74_469 ();
 sg13g2_fill_2 FILLER_74_475 ();
 sg13g2_fill_2 FILLER_74_482 ();
 sg13g2_decap_8 FILLER_74_515 ();
 sg13g2_fill_1 FILLER_74_522 ();
 sg13g2_decap_8 FILLER_74_527 ();
 sg13g2_decap_8 FILLER_74_534 ();
 sg13g2_fill_2 FILLER_74_541 ();
 sg13g2_fill_1 FILLER_74_543 ();
 sg13g2_fill_2 FILLER_74_547 ();
 sg13g2_decap_4 FILLER_74_554 ();
 sg13g2_fill_1 FILLER_74_572 ();
 sg13g2_fill_2 FILLER_74_577 ();
 sg13g2_fill_2 FILLER_74_584 ();
 sg13g2_fill_2 FILLER_74_589 ();
 sg13g2_decap_8 FILLER_74_636 ();
 sg13g2_decap_4 FILLER_74_643 ();
 sg13g2_fill_1 FILLER_74_665 ();
 sg13g2_fill_1 FILLER_74_675 ();
 sg13g2_fill_1 FILLER_74_681 ();
 sg13g2_fill_1 FILLER_74_687 ();
 sg13g2_fill_1 FILLER_74_692 ();
 sg13g2_fill_2 FILLER_74_698 ();
 sg13g2_fill_1 FILLER_74_709 ();
 sg13g2_decap_8 FILLER_74_714 ();
 sg13g2_fill_2 FILLER_74_721 ();
 sg13g2_decap_4 FILLER_74_728 ();
 sg13g2_fill_1 FILLER_74_741 ();
 sg13g2_decap_8 FILLER_74_751 ();
 sg13g2_decap_4 FILLER_74_758 ();
 sg13g2_fill_2 FILLER_74_766 ();
 sg13g2_fill_1 FILLER_74_768 ();
 sg13g2_decap_4 FILLER_74_774 ();
 sg13g2_fill_1 FILLER_74_778 ();
 sg13g2_fill_1 FILLER_74_795 ();
 sg13g2_decap_8 FILLER_74_813 ();
 sg13g2_decap_8 FILLER_74_820 ();
 sg13g2_fill_1 FILLER_74_827 ();
 sg13g2_decap_8 FILLER_74_854 ();
 sg13g2_fill_2 FILLER_74_861 ();
 sg13g2_fill_1 FILLER_74_863 ();
 sg13g2_decap_8 FILLER_74_869 ();
 sg13g2_fill_2 FILLER_74_876 ();
 sg13g2_decap_4 FILLER_74_883 ();
 sg13g2_fill_1 FILLER_74_887 ();
 sg13g2_fill_1 FILLER_74_923 ();
 sg13g2_fill_2 FILLER_74_938 ();
 sg13g2_fill_2 FILLER_74_1011 ();
 sg13g2_decap_8 FILLER_74_1044 ();
 sg13g2_decap_8 FILLER_74_1051 ();
 sg13g2_fill_1 FILLER_74_1058 ();
 sg13g2_fill_2 FILLER_74_1085 ();
 sg13g2_fill_1 FILLER_74_1087 ();
 sg13g2_decap_4 FILLER_74_1093 ();
 sg13g2_fill_2 FILLER_74_1097 ();
 sg13g2_fill_2 FILLER_74_1103 ();
 sg13g2_fill_1 FILLER_74_1105 ();
 sg13g2_decap_8 FILLER_74_1110 ();
 sg13g2_decap_8 FILLER_74_1146 ();
 sg13g2_decap_8 FILLER_74_1167 ();
 sg13g2_fill_1 FILLER_74_1174 ();
 sg13g2_fill_1 FILLER_74_1179 ();
 sg13g2_fill_2 FILLER_74_1184 ();
 sg13g2_fill_1 FILLER_74_1186 ();
 sg13g2_fill_1 FILLER_74_1192 ();
 sg13g2_fill_2 FILLER_74_1197 ();
 sg13g2_fill_1 FILLER_74_1260 ();
 sg13g2_decap_8 FILLER_74_1265 ();
 sg13g2_fill_2 FILLER_74_1272 ();
 sg13g2_decap_8 FILLER_74_1281 ();
 sg13g2_fill_1 FILLER_74_1288 ();
 sg13g2_decap_8 FILLER_74_1315 ();
 sg13g2_decap_4 FILLER_74_1322 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_4 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_15 ();
 sg13g2_decap_8 FILLER_75_22 ();
 sg13g2_decap_8 FILLER_75_29 ();
 sg13g2_decap_8 FILLER_75_36 ();
 sg13g2_fill_1 FILLER_75_52 ();
 sg13g2_decap_4 FILLER_75_57 ();
 sg13g2_fill_2 FILLER_75_65 ();
 sg13g2_fill_1 FILLER_75_67 ();
 sg13g2_decap_4 FILLER_75_72 ();
 sg13g2_fill_2 FILLER_75_76 ();
 sg13g2_fill_1 FILLER_75_125 ();
 sg13g2_decap_8 FILLER_75_130 ();
 sg13g2_decap_4 FILLER_75_137 ();
 sg13g2_fill_1 FILLER_75_141 ();
 sg13g2_fill_2 FILLER_75_147 ();
 sg13g2_decap_4 FILLER_75_154 ();
 sg13g2_fill_1 FILLER_75_214 ();
 sg13g2_fill_2 FILLER_75_223 ();
 sg13g2_fill_1 FILLER_75_234 ();
 sg13g2_fill_2 FILLER_75_248 ();
 sg13g2_fill_1 FILLER_75_250 ();
 sg13g2_fill_2 FILLER_75_259 ();
 sg13g2_fill_2 FILLER_75_269 ();
 sg13g2_decap_4 FILLER_75_308 ();
 sg13g2_fill_1 FILLER_75_312 ();
 sg13g2_fill_1 FILLER_75_339 ();
 sg13g2_fill_2 FILLER_75_348 ();
 sg13g2_fill_1 FILLER_75_350 ();
 sg13g2_fill_1 FILLER_75_355 ();
 sg13g2_fill_2 FILLER_75_361 ();
 sg13g2_fill_2 FILLER_75_368 ();
 sg13g2_decap_4 FILLER_75_388 ();
 sg13g2_fill_1 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_397 ();
 sg13g2_decap_8 FILLER_75_404 ();
 sg13g2_decap_8 FILLER_75_411 ();
 sg13g2_fill_2 FILLER_75_418 ();
 sg13g2_fill_1 FILLER_75_420 ();
 sg13g2_decap_4 FILLER_75_426 ();
 sg13g2_fill_2 FILLER_75_430 ();
 sg13g2_fill_1 FILLER_75_440 ();
 sg13g2_fill_2 FILLER_75_446 ();
 sg13g2_fill_1 FILLER_75_448 ();
 sg13g2_fill_1 FILLER_75_473 ();
 sg13g2_fill_1 FILLER_75_501 ();
 sg13g2_decap_8 FILLER_75_507 ();
 sg13g2_fill_2 FILLER_75_514 ();
 sg13g2_fill_1 FILLER_75_516 ();
 sg13g2_fill_1 FILLER_75_543 ();
 sg13g2_fill_2 FILLER_75_555 ();
 sg13g2_fill_2 FILLER_75_589 ();
 sg13g2_fill_2 FILLER_75_605 ();
 sg13g2_decap_8 FILLER_75_611 ();
 sg13g2_decap_8 FILLER_75_618 ();
 sg13g2_fill_2 FILLER_75_625 ();
 sg13g2_fill_1 FILLER_75_627 ();
 sg13g2_fill_2 FILLER_75_637 ();
 sg13g2_fill_1 FILLER_75_644 ();
 sg13g2_fill_1 FILLER_75_649 ();
 sg13g2_fill_1 FILLER_75_656 ();
 sg13g2_fill_1 FILLER_75_670 ();
 sg13g2_fill_1 FILLER_75_689 ();
 sg13g2_decap_4 FILLER_75_693 ();
 sg13g2_fill_2 FILLER_75_697 ();
 sg13g2_fill_1 FILLER_75_746 ();
 sg13g2_fill_1 FILLER_75_773 ();
 sg13g2_fill_2 FILLER_75_779 ();
 sg13g2_fill_1 FILLER_75_786 ();
 sg13g2_fill_1 FILLER_75_792 ();
 sg13g2_fill_2 FILLER_75_798 ();
 sg13g2_fill_2 FILLER_75_804 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_fill_2 FILLER_75_822 ();
 sg13g2_fill_1 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_828 ();
 sg13g2_decap_8 FILLER_75_848 ();
 sg13g2_fill_2 FILLER_75_855 ();
 sg13g2_fill_1 FILLER_75_888 ();
 sg13g2_fill_2 FILLER_75_893 ();
 sg13g2_fill_1 FILLER_75_895 ();
 sg13g2_decap_4 FILLER_75_901 ();
 sg13g2_fill_1 FILLER_75_905 ();
 sg13g2_fill_1 FILLER_75_914 ();
 sg13g2_fill_2 FILLER_75_925 ();
 sg13g2_fill_2 FILLER_75_938 ();
 sg13g2_fill_2 FILLER_75_943 ();
 sg13g2_fill_1 FILLER_75_959 ();
 sg13g2_fill_1 FILLER_75_963 ();
 sg13g2_decap_8 FILLER_75_972 ();
 sg13g2_fill_2 FILLER_75_996 ();
 sg13g2_fill_2 FILLER_75_1002 ();
 sg13g2_fill_1 FILLER_75_1004 ();
 sg13g2_decap_4 FILLER_75_1013 ();
 sg13g2_fill_2 FILLER_75_1017 ();
 sg13g2_fill_1 FILLER_75_1024 ();
 sg13g2_fill_2 FILLER_75_1064 ();
 sg13g2_decap_8 FILLER_75_1079 ();
 sg13g2_decap_8 FILLER_75_1086 ();
 sg13g2_decap_8 FILLER_75_1105 ();
 sg13g2_fill_1 FILLER_75_1125 ();
 sg13g2_fill_1 FILLER_75_1130 ();
 sg13g2_fill_1 FILLER_75_1170 ();
 sg13g2_fill_2 FILLER_75_1174 ();
 sg13g2_decap_4 FILLER_75_1188 ();
 sg13g2_fill_1 FILLER_75_1192 ();
 sg13g2_fill_2 FILLER_75_1198 ();
 sg13g2_decap_8 FILLER_75_1204 ();
 sg13g2_decap_8 FILLER_75_1215 ();
 sg13g2_decap_8 FILLER_75_1222 ();
 sg13g2_decap_8 FILLER_75_1229 ();
 sg13g2_decap_8 FILLER_75_1240 ();
 sg13g2_decap_8 FILLER_75_1247 ();
 sg13g2_decap_8 FILLER_75_1280 ();
 sg13g2_decap_8 FILLER_75_1287 ();
 sg13g2_decap_8 FILLER_75_1294 ();
 sg13g2_decap_8 FILLER_75_1301 ();
 sg13g2_decap_8 FILLER_75_1308 ();
 sg13g2_decap_8 FILLER_75_1315 ();
 sg13g2_decap_4 FILLER_75_1322 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_decap_4 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_32 ();
 sg13g2_fill_2 FILLER_76_89 ();
 sg13g2_decap_4 FILLER_76_100 ();
 sg13g2_fill_2 FILLER_76_108 ();
 sg13g2_fill_1 FILLER_76_110 ();
 sg13g2_fill_2 FILLER_76_137 ();
 sg13g2_fill_1 FILLER_76_139 ();
 sg13g2_decap_4 FILLER_76_144 ();
 sg13g2_fill_2 FILLER_76_148 ();
 sg13g2_fill_2 FILLER_76_167 ();
 sg13g2_fill_2 FILLER_76_173 ();
 sg13g2_decap_4 FILLER_76_181 ();
 sg13g2_fill_2 FILLER_76_185 ();
 sg13g2_fill_2 FILLER_76_193 ();
 sg13g2_fill_1 FILLER_76_195 ();
 sg13g2_decap_8 FILLER_76_201 ();
 sg13g2_decap_8 FILLER_76_208 ();
 sg13g2_decap_4 FILLER_76_215 ();
 sg13g2_fill_1 FILLER_76_219 ();
 sg13g2_fill_1 FILLER_76_224 ();
 sg13g2_fill_1 FILLER_76_230 ();
 sg13g2_fill_1 FILLER_76_261 ();
 sg13g2_decap_4 FILLER_76_266 ();
 sg13g2_fill_2 FILLER_76_270 ();
 sg13g2_fill_1 FILLER_76_277 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_fill_2 FILLER_76_294 ();
 sg13g2_fill_2 FILLER_76_301 ();
 sg13g2_decap_4 FILLER_76_329 ();
 sg13g2_fill_1 FILLER_76_333 ();
 sg13g2_decap_8 FILLER_76_355 ();
 sg13g2_fill_2 FILLER_76_362 ();
 sg13g2_fill_2 FILLER_76_428 ();
 sg13g2_decap_8 FILLER_76_448 ();
 sg13g2_decap_4 FILLER_76_455 ();
 sg13g2_decap_4 FILLER_76_466 ();
 sg13g2_fill_1 FILLER_76_470 ();
 sg13g2_fill_1 FILLER_76_475 ();
 sg13g2_decap_4 FILLER_76_485 ();
 sg13g2_fill_2 FILLER_76_489 ();
 sg13g2_fill_2 FILLER_76_506 ();
 sg13g2_fill_2 FILLER_76_534 ();
 sg13g2_fill_1 FILLER_76_551 ();
 sg13g2_decap_4 FILLER_76_573 ();
 sg13g2_fill_2 FILLER_76_601 ();
 sg13g2_fill_2 FILLER_76_629 ();
 sg13g2_fill_1 FILLER_76_631 ();
 sg13g2_fill_1 FILLER_76_637 ();
 sg13g2_fill_1 FILLER_76_671 ();
 sg13g2_decap_8 FILLER_76_683 ();
 sg13g2_decap_4 FILLER_76_690 ();
 sg13g2_fill_2 FILLER_76_694 ();
 sg13g2_decap_4 FILLER_76_700 ();
 sg13g2_fill_1 FILLER_76_704 ();
 sg13g2_decap_8 FILLER_76_710 ();
 sg13g2_decap_8 FILLER_76_717 ();
 sg13g2_decap_4 FILLER_76_724 ();
 sg13g2_fill_2 FILLER_76_728 ();
 sg13g2_fill_2 FILLER_76_746 ();
 sg13g2_decap_4 FILLER_76_778 ();
 sg13g2_fill_2 FILLER_76_787 ();
 sg13g2_fill_1 FILLER_76_789 ();
 sg13g2_fill_2 FILLER_76_809 ();
 sg13g2_fill_1 FILLER_76_811 ();
 sg13g2_fill_2 FILLER_76_838 ();
 sg13g2_fill_1 FILLER_76_840 ();
 sg13g2_fill_2 FILLER_76_871 ();
 sg13g2_fill_1 FILLER_76_878 ();
 sg13g2_fill_2 FILLER_76_884 ();
 sg13g2_fill_2 FILLER_76_890 ();
 sg13g2_fill_1 FILLER_76_892 ();
 sg13g2_fill_1 FILLER_76_898 ();
 sg13g2_fill_2 FILLER_76_904 ();
 sg13g2_fill_1 FILLER_76_906 ();
 sg13g2_fill_1 FILLER_76_915 ();
 sg13g2_fill_2 FILLER_76_924 ();
 sg13g2_fill_2 FILLER_76_948 ();
 sg13g2_fill_1 FILLER_76_950 ();
 sg13g2_decap_4 FILLER_76_962 ();
 sg13g2_fill_2 FILLER_76_966 ();
 sg13g2_decap_8 FILLER_76_975 ();
 sg13g2_decap_8 FILLER_76_982 ();
 sg13g2_decap_8 FILLER_76_989 ();
 sg13g2_fill_2 FILLER_76_996 ();
 sg13g2_fill_1 FILLER_76_998 ();
 sg13g2_fill_2 FILLER_76_1030 ();
 sg13g2_fill_1 FILLER_76_1032 ();
 sg13g2_decap_8 FILLER_76_1053 ();
 sg13g2_fill_1 FILLER_76_1060 ();
 sg13g2_fill_1 FILLER_76_1065 ();
 sg13g2_fill_1 FILLER_76_1092 ();
 sg13g2_fill_1 FILLER_76_1119 ();
 sg13g2_fill_2 FILLER_76_1125 ();
 sg13g2_fill_2 FILLER_76_1131 ();
 sg13g2_fill_1 FILLER_76_1133 ();
 sg13g2_fill_1 FILLER_76_1146 ();
 sg13g2_decap_8 FILLER_76_1185 ();
 sg13g2_fill_1 FILLER_76_1192 ();
 sg13g2_decap_8 FILLER_76_1219 ();
 sg13g2_decap_8 FILLER_76_1226 ();
 sg13g2_decap_8 FILLER_76_1233 ();
 sg13g2_decap_8 FILLER_76_1240 ();
 sg13g2_decap_8 FILLER_76_1247 ();
 sg13g2_decap_8 FILLER_76_1254 ();
 sg13g2_decap_8 FILLER_76_1261 ();
 sg13g2_decap_8 FILLER_76_1268 ();
 sg13g2_decap_8 FILLER_76_1275 ();
 sg13g2_decap_8 FILLER_76_1282 ();
 sg13g2_decap_8 FILLER_76_1289 ();
 sg13g2_decap_8 FILLER_76_1296 ();
 sg13g2_decap_8 FILLER_76_1303 ();
 sg13g2_decap_8 FILLER_76_1310 ();
 sg13g2_decap_8 FILLER_76_1317 ();
 sg13g2_fill_2 FILLER_76_1324 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_6 ();
 sg13g2_fill_1 FILLER_77_8 ();
 sg13g2_fill_2 FILLER_77_35 ();
 sg13g2_fill_1 FILLER_77_37 ();
 sg13g2_fill_2 FILLER_77_42 ();
 sg13g2_fill_2 FILLER_77_49 ();
 sg13g2_fill_2 FILLER_77_55 ();
 sg13g2_fill_1 FILLER_77_57 ();
 sg13g2_decap_4 FILLER_77_75 ();
 sg13g2_fill_2 FILLER_77_79 ();
 sg13g2_decap_8 FILLER_77_85 ();
 sg13g2_fill_2 FILLER_77_92 ();
 sg13g2_decap_8 FILLER_77_102 ();
 sg13g2_decap_8 FILLER_77_109 ();
 sg13g2_fill_1 FILLER_77_116 ();
 sg13g2_decap_4 FILLER_77_121 ();
 sg13g2_fill_1 FILLER_77_213 ();
 sg13g2_fill_1 FILLER_77_240 ();
 sg13g2_decap_4 FILLER_77_245 ();
 sg13g2_fill_2 FILLER_77_249 ();
 sg13g2_fill_2 FILLER_77_277 ();
 sg13g2_fill_2 FILLER_77_313 ();
 sg13g2_decap_4 FILLER_77_341 ();
 sg13g2_decap_8 FILLER_77_375 ();
 sg13g2_decap_8 FILLER_77_382 ();
 sg13g2_decap_8 FILLER_77_389 ();
 sg13g2_decap_4 FILLER_77_396 ();
 sg13g2_decap_8 FILLER_77_404 ();
 sg13g2_decap_8 FILLER_77_411 ();
 sg13g2_decap_8 FILLER_77_418 ();
 sg13g2_fill_2 FILLER_77_429 ();
 sg13g2_fill_2 FILLER_77_440 ();
 sg13g2_decap_8 FILLER_77_446 ();
 sg13g2_fill_2 FILLER_77_453 ();
 sg13g2_fill_1 FILLER_77_455 ();
 sg13g2_fill_1 FILLER_77_474 ();
 sg13g2_decap_8 FILLER_77_479 ();
 sg13g2_decap_8 FILLER_77_486 ();
 sg13g2_decap_8 FILLER_77_493 ();
 sg13g2_fill_1 FILLER_77_500 ();
 sg13g2_decap_4 FILLER_77_508 ();
 sg13g2_fill_2 FILLER_77_512 ();
 sg13g2_fill_2 FILLER_77_529 ();
 sg13g2_decap_8 FILLER_77_535 ();
 sg13g2_decap_8 FILLER_77_542 ();
 sg13g2_fill_1 FILLER_77_549 ();
 sg13g2_decap_8 FILLER_77_555 ();
 sg13g2_fill_2 FILLER_77_598 ();
 sg13g2_fill_1 FILLER_77_600 ();
 sg13g2_fill_1 FILLER_77_606 ();
 sg13g2_decap_8 FILLER_77_611 ();
 sg13g2_decap_8 FILLER_77_618 ();
 sg13g2_decap_8 FILLER_77_625 ();
 sg13g2_decap_8 FILLER_77_632 ();
 sg13g2_decap_4 FILLER_77_639 ();
 sg13g2_fill_2 FILLER_77_643 ();
 sg13g2_fill_2 FILLER_77_666 ();
 sg13g2_fill_1 FILLER_77_698 ();
 sg13g2_fill_1 FILLER_77_722 ();
 sg13g2_fill_2 FILLER_77_737 ();
 sg13g2_fill_1 FILLER_77_748 ();
 sg13g2_decap_8 FILLER_77_757 ();
 sg13g2_decap_8 FILLER_77_764 ();
 sg13g2_fill_2 FILLER_77_771 ();
 sg13g2_fill_1 FILLER_77_773 ();
 sg13g2_fill_1 FILLER_77_805 ();
 sg13g2_fill_2 FILLER_77_811 ();
 sg13g2_fill_1 FILLER_77_813 ();
 sg13g2_decap_8 FILLER_77_823 ();
 sg13g2_fill_1 FILLER_77_830 ();
 sg13g2_decap_4 FILLER_77_843 ();
 sg13g2_fill_2 FILLER_77_847 ();
 sg13g2_fill_2 FILLER_77_857 ();
 sg13g2_fill_1 FILLER_77_859 ();
 sg13g2_fill_2 FILLER_77_868 ();
 sg13g2_decap_8 FILLER_77_875 ();
 sg13g2_fill_2 FILLER_77_882 ();
 sg13g2_decap_4 FILLER_77_889 ();
 sg13g2_fill_1 FILLER_77_893 ();
 sg13g2_fill_2 FILLER_77_899 ();
 sg13g2_fill_2 FILLER_77_909 ();
 sg13g2_fill_1 FILLER_77_911 ();
 sg13g2_fill_2 FILLER_77_920 ();
 sg13g2_fill_2 FILLER_77_925 ();
 sg13g2_fill_2 FILLER_77_932 ();
 sg13g2_decap_8 FILLER_77_939 ();
 sg13g2_fill_2 FILLER_77_1024 ();
 sg13g2_decap_4 FILLER_77_1095 ();
 sg13g2_fill_1 FILLER_77_1099 ();
 sg13g2_decap_8 FILLER_77_1107 ();
 sg13g2_decap_8 FILLER_77_1149 ();
 sg13g2_fill_1 FILLER_77_1156 ();
 sg13g2_decap_4 FILLER_77_1161 ();
 sg13g2_fill_2 FILLER_77_1165 ();
 sg13g2_fill_2 FILLER_77_1170 ();
 sg13g2_decap_8 FILLER_77_1222 ();
 sg13g2_decap_8 FILLER_77_1229 ();
 sg13g2_decap_8 FILLER_77_1236 ();
 sg13g2_decap_8 FILLER_77_1243 ();
 sg13g2_decap_8 FILLER_77_1250 ();
 sg13g2_decap_8 FILLER_77_1257 ();
 sg13g2_decap_8 FILLER_77_1264 ();
 sg13g2_decap_8 FILLER_77_1271 ();
 sg13g2_decap_8 FILLER_77_1278 ();
 sg13g2_decap_8 FILLER_77_1285 ();
 sg13g2_decap_8 FILLER_77_1292 ();
 sg13g2_decap_8 FILLER_77_1299 ();
 sg13g2_decap_8 FILLER_77_1306 ();
 sg13g2_decap_8 FILLER_77_1313 ();
 sg13g2_decap_4 FILLER_77_1320 ();
 sg13g2_fill_2 FILLER_77_1324 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_4 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_11 ();
 sg13g2_fill_1 FILLER_78_16 ();
 sg13g2_fill_1 FILLER_78_64 ();
 sg13g2_fill_1 FILLER_78_69 ();
 sg13g2_decap_8 FILLER_78_74 ();
 sg13g2_decap_4 FILLER_78_81 ();
 sg13g2_fill_1 FILLER_78_85 ();
 sg13g2_fill_2 FILLER_78_99 ();
 sg13g2_fill_1 FILLER_78_101 ();
 sg13g2_decap_4 FILLER_78_106 ();
 sg13g2_fill_1 FILLER_78_110 ();
 sg13g2_fill_2 FILLER_78_115 ();
 sg13g2_fill_1 FILLER_78_117 ();
 sg13g2_decap_8 FILLER_78_122 ();
 sg13g2_decap_4 FILLER_78_129 ();
 sg13g2_fill_1 FILLER_78_191 ();
 sg13g2_fill_2 FILLER_78_207 ();
 sg13g2_fill_1 FILLER_78_209 ();
 sg13g2_decap_8 FILLER_78_236 ();
 sg13g2_fill_1 FILLER_78_243 ();
 sg13g2_decap_8 FILLER_78_270 ();
 sg13g2_decap_8 FILLER_78_277 ();
 sg13g2_decap_8 FILLER_78_296 ();
 sg13g2_decap_8 FILLER_78_303 ();
 sg13g2_decap_4 FILLER_78_310 ();
 sg13g2_fill_2 FILLER_78_314 ();
 sg13g2_decap_4 FILLER_78_355 ();
 sg13g2_decap_8 FILLER_78_363 ();
 sg13g2_decap_8 FILLER_78_370 ();
 sg13g2_decap_8 FILLER_78_377 ();
 sg13g2_fill_2 FILLER_78_388 ();
 sg13g2_fill_1 FILLER_78_395 ();
 sg13g2_fill_2 FILLER_78_422 ();
 sg13g2_fill_1 FILLER_78_428 ();
 sg13g2_fill_2 FILLER_78_433 ();
 sg13g2_fill_2 FILLER_78_439 ();
 sg13g2_decap_8 FILLER_78_450 ();
 sg13g2_decap_4 FILLER_78_457 ();
 sg13g2_fill_1 FILLER_78_461 ();
 sg13g2_fill_1 FILLER_78_476 ();
 sg13g2_fill_1 FILLER_78_481 ();
 sg13g2_fill_2 FILLER_78_500 ();
 sg13g2_fill_2 FILLER_78_507 ();
 sg13g2_fill_1 FILLER_78_509 ();
 sg13g2_decap_8 FILLER_78_536 ();
 sg13g2_decap_8 FILLER_78_547 ();
 sg13g2_decap_8 FILLER_78_554 ();
 sg13g2_fill_1 FILLER_78_561 ();
 sg13g2_fill_2 FILLER_78_570 ();
 sg13g2_decap_4 FILLER_78_582 ();
 sg13g2_fill_2 FILLER_78_591 ();
 sg13g2_fill_2 FILLER_78_619 ();
 sg13g2_fill_1 FILLER_78_621 ();
 sg13g2_fill_1 FILLER_78_648 ();
 sg13g2_fill_1 FILLER_78_653 ();
 sg13g2_fill_1 FILLER_78_658 ();
 sg13g2_fill_1 FILLER_78_670 ();
 sg13g2_decap_8 FILLER_78_684 ();
 sg13g2_decap_4 FILLER_78_691 ();
 sg13g2_fill_2 FILLER_78_709 ();
 sg13g2_decap_8 FILLER_78_718 ();
 sg13g2_decap_8 FILLER_78_730 ();
 sg13g2_fill_1 FILLER_78_742 ();
 sg13g2_fill_2 FILLER_78_772 ();
 sg13g2_fill_2 FILLER_78_803 ();
 sg13g2_fill_1 FILLER_78_835 ();
 sg13g2_decap_8 FILLER_78_845 ();
 sg13g2_fill_2 FILLER_78_856 ();
 sg13g2_decap_4 FILLER_78_862 ();
 sg13g2_fill_2 FILLER_78_866 ();
 sg13g2_decap_8 FILLER_78_872 ();
 sg13g2_fill_2 FILLER_78_879 ();
 sg13g2_fill_1 FILLER_78_881 ();
 sg13g2_fill_1 FILLER_78_908 ();
 sg13g2_fill_1 FILLER_78_935 ();
 sg13g2_fill_1 FILLER_78_983 ();
 sg13g2_fill_2 FILLER_78_989 ();
 sg13g2_fill_2 FILLER_78_995 ();
 sg13g2_fill_2 FILLER_78_1001 ();
 sg13g2_decap_8 FILLER_78_1008 ();
 sg13g2_decap_8 FILLER_78_1015 ();
 sg13g2_fill_2 FILLER_78_1022 ();
 sg13g2_decap_4 FILLER_78_1029 ();
 sg13g2_fill_1 FILLER_78_1033 ();
 sg13g2_decap_8 FILLER_78_1038 ();
 sg13g2_decap_8 FILLER_78_1045 ();
 sg13g2_decap_8 FILLER_78_1052 ();
 sg13g2_fill_2 FILLER_78_1059 ();
 sg13g2_fill_1 FILLER_78_1061 ();
 sg13g2_decap_8 FILLER_78_1071 ();
 sg13g2_fill_1 FILLER_78_1078 ();
 sg13g2_fill_2 FILLER_78_1082 ();
 sg13g2_decap_8 FILLER_78_1115 ();
 sg13g2_fill_2 FILLER_78_1122 ();
 sg13g2_fill_1 FILLER_78_1124 ();
 sg13g2_decap_4 FILLER_78_1129 ();
 sg13g2_fill_1 FILLER_78_1133 ();
 sg13g2_fill_2 FILLER_78_1141 ();
 sg13g2_fill_1 FILLER_78_1143 ();
 sg13g2_fill_1 FILLER_78_1170 ();
 sg13g2_decap_4 FILLER_78_1183 ();
 sg13g2_fill_1 FILLER_78_1187 ();
 sg13g2_fill_2 FILLER_78_1192 ();
 sg13g2_decap_8 FILLER_78_1198 ();
 sg13g2_decap_8 FILLER_78_1205 ();
 sg13g2_decap_8 FILLER_78_1212 ();
 sg13g2_decap_8 FILLER_78_1219 ();
 sg13g2_decap_8 FILLER_78_1226 ();
 sg13g2_decap_8 FILLER_78_1233 ();
 sg13g2_decap_8 FILLER_78_1240 ();
 sg13g2_decap_8 FILLER_78_1247 ();
 sg13g2_decap_8 FILLER_78_1254 ();
 sg13g2_decap_8 FILLER_78_1261 ();
 sg13g2_decap_8 FILLER_78_1268 ();
 sg13g2_decap_8 FILLER_78_1275 ();
 sg13g2_decap_8 FILLER_78_1282 ();
 sg13g2_decap_8 FILLER_78_1289 ();
 sg13g2_decap_8 FILLER_78_1296 ();
 sg13g2_decap_8 FILLER_78_1303 ();
 sg13g2_decap_8 FILLER_78_1310 ();
 sg13g2_decap_8 FILLER_78_1317 ();
 sg13g2_fill_2 FILLER_78_1324 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_fill_2 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_27 ();
 sg13g2_decap_4 FILLER_79_34 ();
 sg13g2_fill_1 FILLER_79_42 ();
 sg13g2_fill_2 FILLER_79_47 ();
 sg13g2_fill_2 FILLER_79_53 ();
 sg13g2_fill_2 FILLER_79_59 ();
 sg13g2_fill_2 FILLER_79_117 ();
 sg13g2_fill_1 FILLER_79_119 ();
 sg13g2_fill_2 FILLER_79_158 ();
 sg13g2_fill_1 FILLER_79_174 ();
 sg13g2_fill_2 FILLER_79_185 ();
 sg13g2_fill_2 FILLER_79_225 ();
 sg13g2_fill_1 FILLER_79_227 ();
 sg13g2_fill_2 FILLER_79_254 ();
 sg13g2_fill_1 FILLER_79_256 ();
 sg13g2_decap_4 FILLER_79_287 ();
 sg13g2_fill_1 FILLER_79_291 ();
 sg13g2_decap_4 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_330 ();
 sg13g2_fill_1 FILLER_79_363 ();
 sg13g2_fill_1 FILLER_79_390 ();
 sg13g2_decap_4 FILLER_79_419 ();
 sg13g2_decap_4 FILLER_79_449 ();
 sg13g2_decap_8 FILLER_79_457 ();
 sg13g2_fill_2 FILLER_79_464 ();
 sg13g2_fill_1 FILLER_79_466 ();
 sg13g2_fill_1 FILLER_79_474 ();
 sg13g2_fill_2 FILLER_79_480 ();
 sg13g2_decap_8 FILLER_79_486 ();
 sg13g2_fill_2 FILLER_79_519 ();
 sg13g2_decap_8 FILLER_79_525 ();
 sg13g2_fill_2 FILLER_79_532 ();
 sg13g2_fill_2 FILLER_79_569 ();
 sg13g2_decap_4 FILLER_79_576 ();
 sg13g2_fill_2 FILLER_79_585 ();
 sg13g2_fill_1 FILLER_79_590 ();
 sg13g2_decap_8 FILLER_79_618 ();
 sg13g2_fill_2 FILLER_79_625 ();
 sg13g2_fill_1 FILLER_79_627 ();
 sg13g2_fill_2 FILLER_79_632 ();
 sg13g2_fill_1 FILLER_79_634 ();
 sg13g2_decap_8 FILLER_79_639 ();
 sg13g2_fill_2 FILLER_79_646 ();
 sg13g2_fill_1 FILLER_79_648 ();
 sg13g2_fill_2 FILLER_79_653 ();
 sg13g2_decap_8 FILLER_79_665 ();
 sg13g2_decap_4 FILLER_79_672 ();
 sg13g2_fill_1 FILLER_79_676 ();
 sg13g2_decap_4 FILLER_79_681 ();
 sg13g2_fill_2 FILLER_79_685 ();
 sg13g2_decap_8 FILLER_79_692 ();
 sg13g2_fill_1 FILLER_79_699 ();
 sg13g2_fill_1 FILLER_79_752 ();
 sg13g2_fill_1 FILLER_79_761 ();
 sg13g2_fill_1 FILLER_79_800 ();
 sg13g2_decap_8 FILLER_79_817 ();
 sg13g2_fill_2 FILLER_79_824 ();
 sg13g2_decap_4 FILLER_79_836 ();
 sg13g2_decap_4 FILLER_79_870 ();
 sg13g2_fill_1 FILLER_79_874 ();
 sg13g2_decap_8 FILLER_79_879 ();
 sg13g2_decap_4 FILLER_79_886 ();
 sg13g2_fill_1 FILLER_79_890 ();
 sg13g2_fill_2 FILLER_79_921 ();
 sg13g2_fill_1 FILLER_79_923 ();
 sg13g2_decap_4 FILLER_79_928 ();
 sg13g2_fill_2 FILLER_79_932 ();
 sg13g2_fill_2 FILLER_79_938 ();
 sg13g2_fill_1 FILLER_79_940 ();
 sg13g2_decap_4 FILLER_79_944 ();
 sg13g2_fill_2 FILLER_79_948 ();
 sg13g2_decap_8 FILLER_79_954 ();
 sg13g2_fill_2 FILLER_79_961 ();
 sg13g2_decap_8 FILLER_79_971 ();
 sg13g2_fill_2 FILLER_79_1056 ();
 sg13g2_fill_1 FILLER_79_1105 ();
 sg13g2_fill_1 FILLER_79_1145 ();
 sg13g2_decap_8 FILLER_79_1150 ();
 sg13g2_fill_2 FILLER_79_1157 ();
 sg13g2_decap_8 FILLER_79_1219 ();
 sg13g2_decap_8 FILLER_79_1226 ();
 sg13g2_decap_8 FILLER_79_1233 ();
 sg13g2_decap_8 FILLER_79_1240 ();
 sg13g2_decap_8 FILLER_79_1247 ();
 sg13g2_decap_8 FILLER_79_1254 ();
 sg13g2_decap_8 FILLER_79_1261 ();
 sg13g2_decap_8 FILLER_79_1268 ();
 sg13g2_decap_8 FILLER_79_1275 ();
 sg13g2_decap_8 FILLER_79_1282 ();
 sg13g2_decap_8 FILLER_79_1289 ();
 sg13g2_decap_8 FILLER_79_1296 ();
 sg13g2_decap_8 FILLER_79_1303 ();
 sg13g2_decap_8 FILLER_79_1310 ();
 sg13g2_decap_8 FILLER_79_1317 ();
 sg13g2_fill_2 FILLER_79_1324 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_4 FILLER_80_28 ();
 sg13g2_fill_2 FILLER_80_62 ();
 sg13g2_fill_1 FILLER_80_64 ();
 sg13g2_fill_1 FILLER_80_113 ();
 sg13g2_fill_1 FILLER_80_170 ();
 sg13g2_fill_1 FILLER_80_224 ();
 sg13g2_fill_1 FILLER_80_229 ();
 sg13g2_fill_2 FILLER_80_234 ();
 sg13g2_decap_4 FILLER_80_244 ();
 sg13g2_fill_1 FILLER_80_248 ();
 sg13g2_decap_8 FILLER_80_253 ();
 sg13g2_decap_4 FILLER_80_260 ();
 sg13g2_fill_1 FILLER_80_264 ();
 sg13g2_decap_4 FILLER_80_273 ();
 sg13g2_fill_2 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_283 ();
 sg13g2_decap_4 FILLER_80_290 ();
 sg13g2_fill_2 FILLER_80_294 ();
 sg13g2_decap_4 FILLER_80_304 ();
 sg13g2_fill_1 FILLER_80_312 ();
 sg13g2_fill_2 FILLER_80_323 ();
 sg13g2_fill_1 FILLER_80_325 ();
 sg13g2_decap_4 FILLER_80_336 ();
 sg13g2_fill_2 FILLER_80_340 ();
 sg13g2_decap_4 FILLER_80_354 ();
 sg13g2_fill_2 FILLER_80_358 ();
 sg13g2_decap_4 FILLER_80_428 ();
 sg13g2_decap_8 FILLER_80_436 ();
 sg13g2_fill_2 FILLER_80_443 ();
 sg13g2_fill_1 FILLER_80_445 ();
 sg13g2_fill_2 FILLER_80_472 ();
 sg13g2_fill_1 FILLER_80_474 ();
 sg13g2_decap_8 FILLER_80_505 ();
 sg13g2_decap_8 FILLER_80_512 ();
 sg13g2_decap_8 FILLER_80_519 ();
 sg13g2_decap_8 FILLER_80_526 ();
 sg13g2_decap_8 FILLER_80_533 ();
 sg13g2_decap_8 FILLER_80_540 ();
 sg13g2_decap_8 FILLER_80_547 ();
 sg13g2_decap_8 FILLER_80_554 ();
 sg13g2_fill_1 FILLER_80_561 ();
 sg13g2_decap_4 FILLER_80_592 ();
 sg13g2_fill_2 FILLER_80_596 ();
 sg13g2_decap_4 FILLER_80_624 ();
 sg13g2_decap_8 FILLER_80_654 ();
 sg13g2_decap_8 FILLER_80_661 ();
 sg13g2_decap_8 FILLER_80_694 ();
 sg13g2_decap_8 FILLER_80_701 ();
 sg13g2_decap_8 FILLER_80_712 ();
 sg13g2_fill_1 FILLER_80_719 ();
 sg13g2_decap_8 FILLER_80_725 ();
 sg13g2_fill_2 FILLER_80_732 ();
 sg13g2_decap_8 FILLER_80_738 ();
 sg13g2_fill_1 FILLER_80_745 ();
 sg13g2_fill_1 FILLER_80_796 ();
 sg13g2_decap_4 FILLER_80_828 ();
 sg13g2_fill_2 FILLER_80_832 ();
 sg13g2_decap_8 FILLER_80_860 ();
 sg13g2_fill_1 FILLER_80_867 ();
 sg13g2_fill_2 FILLER_80_898 ();
 sg13g2_fill_1 FILLER_80_900 ();
 sg13g2_decap_8 FILLER_80_905 ();
 sg13g2_decap_8 FILLER_80_912 ();
 sg13g2_decap_8 FILLER_80_919 ();
 sg13g2_decap_8 FILLER_80_926 ();
 sg13g2_decap_8 FILLER_80_933 ();
 sg13g2_fill_2 FILLER_80_940 ();
 sg13g2_fill_1 FILLER_80_942 ();
 sg13g2_decap_8 FILLER_80_969 ();
 sg13g2_decap_8 FILLER_80_976 ();
 sg13g2_fill_1 FILLER_80_983 ();
 sg13g2_decap_4 FILLER_80_988 ();
 sg13g2_decap_4 FILLER_80_1005 ();
 sg13g2_fill_2 FILLER_80_1009 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_fill_2 FILLER_80_1022 ();
 sg13g2_decap_8 FILLER_80_1028 ();
 sg13g2_decap_4 FILLER_80_1035 ();
 sg13g2_decap_8 FILLER_80_1043 ();
 sg13g2_decap_8 FILLER_80_1050 ();
 sg13g2_fill_1 FILLER_80_1057 ();
 sg13g2_decap_8 FILLER_80_1071 ();
 sg13g2_decap_4 FILLER_80_1078 ();
 sg13g2_fill_2 FILLER_80_1085 ();
 sg13g2_fill_1 FILLER_80_1087 ();
 sg13g2_fill_2 FILLER_80_1114 ();
 sg13g2_fill_1 FILLER_80_1116 ();
 sg13g2_decap_8 FILLER_80_1121 ();
 sg13g2_decap_8 FILLER_80_1128 ();
 sg13g2_fill_2 FILLER_80_1135 ();
 sg13g2_fill_1 FILLER_80_1137 ();
 sg13g2_decap_8 FILLER_80_1164 ();
 sg13g2_decap_4 FILLER_80_1171 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_fill_2 FILLER_80_1186 ();
 sg13g2_fill_1 FILLER_80_1188 ();
 sg13g2_decap_8 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1205 ();
 sg13g2_decap_8 FILLER_80_1212 ();
 sg13g2_decap_8 FILLER_80_1219 ();
 sg13g2_decap_8 FILLER_80_1226 ();
 sg13g2_decap_8 FILLER_80_1233 ();
 sg13g2_decap_8 FILLER_80_1240 ();
 sg13g2_decap_8 FILLER_80_1247 ();
 sg13g2_decap_8 FILLER_80_1254 ();
 sg13g2_decap_8 FILLER_80_1261 ();
 sg13g2_decap_8 FILLER_80_1268 ();
 sg13g2_decap_8 FILLER_80_1275 ();
 sg13g2_decap_8 FILLER_80_1282 ();
 sg13g2_decap_8 FILLER_80_1289 ();
 sg13g2_decap_8 FILLER_80_1296 ();
 sg13g2_decap_8 FILLER_80_1303 ();
 sg13g2_decap_8 FILLER_80_1310 ();
 sg13g2_decap_8 FILLER_80_1317 ();
 sg13g2_fill_2 FILLER_80_1324 ();
endmodule
