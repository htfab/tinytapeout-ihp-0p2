module tt_um_rebeccargb_intercal_alu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire clknet_0_clk;
 wire \a[0] ;
 wire \a[10] ;
 wire \a[11] ;
 wire \a[12] ;
 wire \a[13] ;
 wire \a[14] ;
 wire \a[15] ;
 wire \a[16] ;
 wire \a[17] ;
 wire \a[18] ;
 wire \a[19] ;
 wire \a[1] ;
 wire \a[20] ;
 wire \a[21] ;
 wire \a[22] ;
 wire \a[23] ;
 wire \a[24] ;
 wire \a[25] ;
 wire \a[26] ;
 wire \a[27] ;
 wire \a[28] ;
 wire \a[29] ;
 wire \a[2] ;
 wire \a[30] ;
 wire \a[31] ;
 wire \a[3] ;
 wire \a[4] ;
 wire \a[5] ;
 wire \a[6] ;
 wire \a[7] ;
 wire \a[8] ;
 wire \a[9] ;
 wire \ayayayayayaya.b[0] ;
 wire \ayayayayayaya.b[10] ;
 wire \ayayayayayaya.b[11] ;
 wire \ayayayayayaya.b[12] ;
 wire \ayayayayayaya.b[13] ;
 wire \ayayayayayaya.b[14] ;
 wire \ayayayayayaya.b[15] ;
 wire \ayayayayayaya.b[16] ;
 wire \ayayayayayaya.b[17] ;
 wire \ayayayayayaya.b[18] ;
 wire \ayayayayayaya.b[19] ;
 wire \ayayayayayaya.b[1] ;
 wire \ayayayayayaya.b[20] ;
 wire \ayayayayayaya.b[21] ;
 wire \ayayayayayaya.b[22] ;
 wire \ayayayayayaya.b[23] ;
 wire \ayayayayayaya.b[24] ;
 wire \ayayayayayaya.b[25] ;
 wire \ayayayayayaya.b[26] ;
 wire \ayayayayayaya.b[27] ;
 wire \ayayayayayaya.b[28] ;
 wire \ayayayayayaya.b[29] ;
 wire \ayayayayayaya.b[2] ;
 wire \ayayayayayaya.b[30] ;
 wire \ayayayayayaya.b[31] ;
 wire \ayayayayayaya.b[3] ;
 wire \ayayayayayaya.b[4] ;
 wire \ayayayayayaya.b[5] ;
 wire \ayayayayayaya.b[6] ;
 wire \ayayayayayaya.b[7] ;
 wire \ayayayayayaya.b[8] ;
 wire \ayayayayayaya.b[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_2 _2262_ (.A(uio_in[0]),
    .X(_1260_));
 sg13g2_inv_1 _2263_ (.Y(_1271_),
    .A(_1260_));
 sg13g2_nor2_1 _2264_ (.A(net1),
    .B(net2),
    .Y(_1282_));
 sg13g2_buf_1 _2265_ (.A(_1282_),
    .X(_1293_));
 sg13g2_inv_1 _2266_ (.Y(_1304_),
    .A(net188));
 sg13g2_buf_1 _2267_ (.A(ui_in[3]),
    .X(_1315_));
 sg13g2_buf_1 _2268_ (.A(ui_in[2]),
    .X(_1325_));
 sg13g2_nor2_1 _2269_ (.A(net189),
    .B(_1325_),
    .Y(_1336_));
 sg13g2_inv_1 _2270_ (.Y(_1347_),
    .A(_1336_));
 sg13g2_nor2_1 _2271_ (.A(_1304_),
    .B(_1347_),
    .Y(_1358_));
 sg13g2_buf_2 _2272_ (.A(_1358_),
    .X(_1369_));
 sg13g2_inv_1 _2273_ (.Y(_1380_),
    .A(_1369_));
 sg13g2_buf_1 _2274_ (.A(ui_in[1]),
    .X(_1391_));
 sg13g2_buf_1 _2275_ (.A(ui_in[0]),
    .X(_1402_));
 sg13g2_nor2_1 _2276_ (.A(_1391_),
    .B(_1402_),
    .Y(_1412_));
 sg13g2_inv_1 _2277_ (.Y(_1423_),
    .A(_1412_));
 sg13g2_nor2_1 _2278_ (.A(net4),
    .B(_1423_),
    .Y(_1434_));
 sg13g2_nor2b_1 _2279_ (.A(net56),
    .B_N(_1434_),
    .Y(_1445_));
 sg13g2_buf_1 _2280_ (.A(_1445_),
    .X(_1456_));
 sg13g2_buf_1 _2281_ (.A(_1456_),
    .X(_1467_));
 sg13g2_buf_1 _2282_ (.A(\a[0] ),
    .X(_1478_));
 sg13g2_nor2_1 _2283_ (.A(net187),
    .B(net36),
    .Y(_1488_));
 sg13g2_a21oi_1 _2284_ (.A1(_1271_),
    .A2(net36),
    .Y(_0060_),
    .B1(_1488_));
 sg13g2_buf_2 _2285_ (.A(uio_in[2]),
    .X(_1509_));
 sg13g2_inv_1 _2286_ (.Y(_1520_),
    .A(_1509_));
 sg13g2_inv_1 _2287_ (.Y(_1531_),
    .A(_1402_));
 sg13g2_nor2_2 _2288_ (.A(_1391_),
    .B(_1531_),
    .Y(_1542_));
 sg13g2_inv_1 _2289_ (.Y(_1553_),
    .A(_1542_));
 sg13g2_nor2_1 _2290_ (.A(net4),
    .B(_1553_),
    .Y(_1563_));
 sg13g2_buf_1 _2291_ (.A(_1369_),
    .X(_1564_));
 sg13g2_nand2_1 _2292_ (.Y(_1565_),
    .A(_1563_),
    .B(net55));
 sg13g2_buf_1 _2293_ (.A(_1565_),
    .X(_1566_));
 sg13g2_buf_1 _2294_ (.A(_1566_),
    .X(_1567_));
 sg13g2_buf_1 _2295_ (.A(\a[10] ),
    .X(_1568_));
 sg13g2_nand2_1 _2296_ (.Y(_1569_),
    .A(_1567_),
    .B(_1568_));
 sg13g2_o21ai_1 _2297_ (.B1(_1569_),
    .Y(_0061_),
    .A1(_1520_),
    .A2(_1567_));
 sg13g2_buf_2 _2298_ (.A(uio_in[3]),
    .X(_1570_));
 sg13g2_inv_1 _2299_ (.Y(_1571_),
    .A(_1570_));
 sg13g2_nand2_1 _2300_ (.Y(_1572_),
    .A(net35),
    .B(\a[11] ));
 sg13g2_o21ai_1 _2301_ (.B1(_1572_),
    .Y(_0062_),
    .A1(_1571_),
    .A2(net35));
 sg13g2_buf_2 _2302_ (.A(uio_in[4]),
    .X(_1573_));
 sg13g2_inv_1 _2303_ (.Y(_1574_),
    .A(_1573_));
 sg13g2_nand2_1 _2304_ (.Y(_1575_),
    .A(_1566_),
    .B(\a[12] ));
 sg13g2_o21ai_1 _2305_ (.B1(_1575_),
    .Y(_0063_),
    .A1(_1574_),
    .A2(net35));
 sg13g2_buf_2 _2306_ (.A(uio_in[5]),
    .X(_1576_));
 sg13g2_inv_1 _2307_ (.Y(_1577_),
    .A(_1576_));
 sg13g2_buf_1 _2308_ (.A(\a[13] ),
    .X(_1578_));
 sg13g2_nand2_1 _2309_ (.Y(_1579_),
    .A(_1566_),
    .B(_1578_));
 sg13g2_o21ai_1 _2310_ (.B1(_1579_),
    .Y(_0064_),
    .A1(_1577_),
    .A2(net35));
 sg13g2_buf_2 _2311_ (.A(uio_in[6]),
    .X(_1580_));
 sg13g2_inv_1 _2312_ (.Y(_1581_),
    .A(_1580_));
 sg13g2_buf_1 _2313_ (.A(\a[14] ),
    .X(_1582_));
 sg13g2_nand2_1 _2314_ (.Y(_1583_),
    .A(_1566_),
    .B(_1582_));
 sg13g2_o21ai_1 _2315_ (.B1(_1583_),
    .Y(_0065_),
    .A1(_1581_),
    .A2(net35));
 sg13g2_buf_2 _2316_ (.A(uio_in[7]),
    .X(_1584_));
 sg13g2_inv_1 _2317_ (.Y(_1585_),
    .A(_1584_));
 sg13g2_buf_1 _2318_ (.A(\a[15] ),
    .X(_1586_));
 sg13g2_nand2_1 _2319_ (.Y(_1587_),
    .A(_1566_),
    .B(net186));
 sg13g2_o21ai_1 _2320_ (.B1(_1587_),
    .Y(_0066_),
    .A1(_1585_),
    .A2(net35));
 sg13g2_buf_2 _2321_ (.A(\a[16] ),
    .X(_1588_));
 sg13g2_inv_1 _2322_ (.Y(_1589_),
    .A(_1588_));
 sg13g2_nand2_1 _2323_ (.Y(_1590_),
    .A(_1531_),
    .B(_1391_));
 sg13g2_buf_2 _2324_ (.A(_1590_),
    .X(_1591_));
 sg13g2_nor2_1 _2325_ (.A(net4),
    .B(_1591_),
    .Y(_1592_));
 sg13g2_nand2_1 _2326_ (.Y(_1593_),
    .A(net55),
    .B(_1592_));
 sg13g2_buf_1 _2327_ (.A(_1593_),
    .X(_1594_));
 sg13g2_buf_1 _2328_ (.A(_1594_),
    .X(_1595_));
 sg13g2_nor2_1 _2329_ (.A(_1260_),
    .B(net34),
    .Y(_1596_));
 sg13g2_a21oi_1 _2330_ (.A1(_1589_),
    .A2(net34),
    .Y(_0067_),
    .B1(_1596_));
 sg13g2_buf_1 _2331_ (.A(\a[17] ),
    .X(_1597_));
 sg13g2_inv_1 _2332_ (.Y(_1598_),
    .A(_1597_));
 sg13g2_buf_2 _2333_ (.A(uio_in[1]),
    .X(_1599_));
 sg13g2_nor2_1 _2334_ (.A(_1599_),
    .B(net34),
    .Y(_1600_));
 sg13g2_a21oi_1 _2335_ (.A1(_1598_),
    .A2(net34),
    .Y(_0068_),
    .B1(_1600_));
 sg13g2_inv_1 _2336_ (.Y(_1601_),
    .A(\a[18] ));
 sg13g2_nor2_1 _2337_ (.A(_1509_),
    .B(_1594_),
    .Y(_1602_));
 sg13g2_a21oi_1 _2338_ (.A1(_1601_),
    .A2(net34),
    .Y(_0069_),
    .B1(_1602_));
 sg13g2_inv_1 _2339_ (.Y(_1603_),
    .A(\a[19] ));
 sg13g2_nor2_1 _2340_ (.A(_1570_),
    .B(_1594_),
    .Y(_1604_));
 sg13g2_a21oi_1 _2341_ (.A1(_1603_),
    .A2(_1595_),
    .Y(_0070_),
    .B1(_1604_));
 sg13g2_inv_1 _2342_ (.Y(_1605_),
    .A(_1599_));
 sg13g2_buf_2 _2343_ (.A(\a[1] ),
    .X(_1606_));
 sg13g2_nor2_1 _2344_ (.A(_1606_),
    .B(_1467_),
    .Y(_1607_));
 sg13g2_a21oi_1 _2345_ (.A1(_1605_),
    .A2(_1467_),
    .Y(_0071_),
    .B1(_1607_));
 sg13g2_inv_1 _2346_ (.Y(_1608_),
    .A(\a[20] ));
 sg13g2_nor2_1 _2347_ (.A(_1573_),
    .B(_1594_),
    .Y(_1609_));
 sg13g2_a21oi_1 _2348_ (.A1(_1608_),
    .A2(net34),
    .Y(_0072_),
    .B1(_1609_));
 sg13g2_buf_1 _2349_ (.A(\a[21] ),
    .X(_1610_));
 sg13g2_inv_1 _2350_ (.Y(_1611_),
    .A(_1610_));
 sg13g2_nor2_1 _2351_ (.A(_1576_),
    .B(_1594_),
    .Y(_1612_));
 sg13g2_a21oi_1 _2352_ (.A1(_1611_),
    .A2(net34),
    .Y(_0073_),
    .B1(_1612_));
 sg13g2_inv_1 _2353_ (.Y(_1613_),
    .A(\a[22] ));
 sg13g2_nor2_1 _2354_ (.A(_1580_),
    .B(_1594_),
    .Y(_1614_));
 sg13g2_a21oi_1 _2355_ (.A1(_1613_),
    .A2(net34),
    .Y(_0074_),
    .B1(_1614_));
 sg13g2_inv_1 _2356_ (.Y(_1615_),
    .A(\a[23] ));
 sg13g2_nor2_1 _2357_ (.A(_1584_),
    .B(_1594_),
    .Y(_1616_));
 sg13g2_a21oi_1 _2358_ (.A1(_1615_),
    .A2(_1595_),
    .Y(_0075_),
    .B1(_1616_));
 sg13g2_buf_1 _2359_ (.A(\a[24] ),
    .X(_1617_));
 sg13g2_inv_1 _2360_ (.Y(_1618_),
    .A(_1617_));
 sg13g2_nand2_1 _2361_ (.Y(_1619_),
    .A(_1391_),
    .B(_1402_));
 sg13g2_buf_8 _2362_ (.A(_1619_),
    .X(_1620_));
 sg13g2_nor2_1 _2363_ (.A(net4),
    .B(_1620_),
    .Y(_1621_));
 sg13g2_nand2_1 _2364_ (.Y(_1622_),
    .A(net55),
    .B(_1621_));
 sg13g2_buf_1 _2365_ (.A(_1622_),
    .X(_1623_));
 sg13g2_buf_1 _2366_ (.A(_1623_),
    .X(_1624_));
 sg13g2_nor2_1 _2367_ (.A(_1260_),
    .B(net33),
    .Y(_1625_));
 sg13g2_a21oi_1 _2368_ (.A1(_1618_),
    .A2(net33),
    .Y(_0076_),
    .B1(_1625_));
 sg13g2_buf_1 _2369_ (.A(\a[25] ),
    .X(_1626_));
 sg13g2_inv_1 _2370_ (.Y(_1627_),
    .A(_1626_));
 sg13g2_nor2_1 _2371_ (.A(_1599_),
    .B(net33),
    .Y(_1628_));
 sg13g2_a21oi_1 _2372_ (.A1(_1627_),
    .A2(_1624_),
    .Y(_0077_),
    .B1(_1628_));
 sg13g2_inv_1 _2373_ (.Y(_1629_),
    .A(\a[26] ));
 sg13g2_nor2_1 _2374_ (.A(_1509_),
    .B(_1623_),
    .Y(_1630_));
 sg13g2_a21oi_1 _2375_ (.A1(_1629_),
    .A2(_1624_),
    .Y(_0078_),
    .B1(_1630_));
 sg13g2_inv_1 _2376_ (.Y(_1631_),
    .A(\a[27] ));
 sg13g2_nor2_1 _2377_ (.A(_1570_),
    .B(_1623_),
    .Y(_1632_));
 sg13g2_a21oi_1 _2378_ (.A1(_1631_),
    .A2(net33),
    .Y(_0079_),
    .B1(_1632_));
 sg13g2_inv_1 _2379_ (.Y(_1633_),
    .A(\a[28] ));
 sg13g2_nor2_1 _2380_ (.A(_1573_),
    .B(_1623_),
    .Y(_1634_));
 sg13g2_a21oi_1 _2381_ (.A1(_1633_),
    .A2(net33),
    .Y(_0080_),
    .B1(_1634_));
 sg13g2_inv_1 _2382_ (.Y(_1635_),
    .A(\a[29] ));
 sg13g2_nor2_1 _2383_ (.A(_1576_),
    .B(_1623_),
    .Y(_1636_));
 sg13g2_a21oi_1 _2384_ (.A1(_1635_),
    .A2(net33),
    .Y(_0081_),
    .B1(_1636_));
 sg13g2_buf_1 _2385_ (.A(\a[2] ),
    .X(_1637_));
 sg13g2_nor2_1 _2386_ (.A(_1637_),
    .B(_1456_),
    .Y(_1638_));
 sg13g2_a21oi_1 _2387_ (.A1(_1520_),
    .A2(net36),
    .Y(_0082_),
    .B1(_1638_));
 sg13g2_buf_1 _2388_ (.A(\a[30] ),
    .X(_1639_));
 sg13g2_inv_1 _2389_ (.Y(_1640_),
    .A(_1639_));
 sg13g2_nor2_1 _2390_ (.A(_1580_),
    .B(_1623_),
    .Y(_1641_));
 sg13g2_a21oi_1 _2391_ (.A1(_1640_),
    .A2(net33),
    .Y(_0083_),
    .B1(_1641_));
 sg13g2_buf_8 _2392_ (.A(\a[31] ),
    .X(_1642_));
 sg13g2_inv_1 _2393_ (.Y(_1643_),
    .A(_1642_));
 sg13g2_nor2_1 _2394_ (.A(_1584_),
    .B(_1623_),
    .Y(_1644_));
 sg13g2_a21oi_1 _2395_ (.A1(_1643_),
    .A2(net33),
    .Y(_0084_),
    .B1(_1644_));
 sg13g2_buf_1 _2396_ (.A(\a[3] ),
    .X(_1645_));
 sg13g2_nor2_1 _2397_ (.A(_1645_),
    .B(_1456_),
    .Y(_1646_));
 sg13g2_a21oi_1 _2398_ (.A1(_1571_),
    .A2(net36),
    .Y(_0085_),
    .B1(_1646_));
 sg13g2_nor2_1 _2399_ (.A(\a[4] ),
    .B(_1456_),
    .Y(_1647_));
 sg13g2_a21oi_1 _2400_ (.A1(_1574_),
    .A2(net36),
    .Y(_0086_),
    .B1(_1647_));
 sg13g2_nor2_1 _2401_ (.A(\a[5] ),
    .B(_1456_),
    .Y(_1648_));
 sg13g2_a21oi_1 _2402_ (.A1(_1577_),
    .A2(net36),
    .Y(_0087_),
    .B1(_1648_));
 sg13g2_nor2_1 _2403_ (.A(\a[6] ),
    .B(_1456_),
    .Y(_1649_));
 sg13g2_a21oi_1 _2404_ (.A1(_1581_),
    .A2(net36),
    .Y(_0088_),
    .B1(_1649_));
 sg13g2_buf_1 _2405_ (.A(\a[7] ),
    .X(_1650_));
 sg13g2_nor2_1 _2406_ (.A(_1650_),
    .B(_1456_),
    .Y(_1651_));
 sg13g2_a21oi_1 _2407_ (.A1(_1585_),
    .A2(net36),
    .Y(_0089_),
    .B1(_1651_));
 sg13g2_buf_1 _2408_ (.A(\a[8] ),
    .X(_1652_));
 sg13g2_nand2_1 _2409_ (.Y(_1653_),
    .A(_1566_),
    .B(_1652_));
 sg13g2_o21ai_1 _2410_ (.B1(_1653_),
    .Y(_0090_),
    .A1(_1271_),
    .A2(net35));
 sg13g2_nand2_1 _2411_ (.Y(_1654_),
    .A(_1566_),
    .B(\a[9] ));
 sg13g2_o21ai_1 _2412_ (.B1(_1654_),
    .Y(_0091_),
    .A1(_1605_),
    .A2(net35));
 sg13g2_buf_1 _2413_ (.A(\ayayayayayaya.b[0] ),
    .X(_1655_));
 sg13g2_inv_2 _2414_ (.Y(_1656_),
    .A(_1655_));
 sg13g2_buf_1 _2415_ (.A(_1656_),
    .X(_1657_));
 sg13g2_buf_1 _2416_ (.A(_1304_),
    .X(_1658_));
 sg13g2_inv_1 _2417_ (.Y(_1659_),
    .A(_1325_));
 sg13g2_nor2_1 _2418_ (.A(net189),
    .B(_1659_),
    .Y(_1660_));
 sg13g2_buf_2 _2419_ (.A(_1660_),
    .X(_1661_));
 sg13g2_inv_1 _2420_ (.Y(_1662_),
    .A(_1661_));
 sg13g2_nor2_1 _2421_ (.A(net138),
    .B(_1662_),
    .Y(_1663_));
 sg13g2_buf_1 _2422_ (.A(_1663_),
    .X(_1664_));
 sg13g2_nand2_1 _2423_ (.Y(_1665_),
    .A(net42),
    .B(_1434_));
 sg13g2_buf_1 _2424_ (.A(_1665_),
    .X(_1666_));
 sg13g2_buf_1 _2425_ (.A(_1666_),
    .X(_1667_));
 sg13g2_nor2_1 _2426_ (.A(_1260_),
    .B(_1667_),
    .Y(_1668_));
 sg13g2_a21oi_1 _2427_ (.A1(net139),
    .A2(_1667_),
    .Y(_0092_),
    .B1(_1668_));
 sg13g2_buf_1 _2428_ (.A(\ayayayayayaya.b[10] ),
    .X(_1669_));
 sg13g2_inv_1 _2429_ (.Y(_1670_),
    .A(net185));
 sg13g2_buf_1 _2430_ (.A(_1670_),
    .X(_1671_));
 sg13g2_buf_1 _2431_ (.A(net137),
    .X(_1672_));
 sg13g2_buf_1 _2432_ (.A(net91),
    .X(_1673_));
 sg13g2_nand2_1 _2433_ (.Y(_1674_),
    .A(_1664_),
    .B(_1563_));
 sg13g2_buf_2 _2434_ (.A(_1674_),
    .X(_1675_));
 sg13g2_buf_1 _2435_ (.A(_1675_),
    .X(_1676_));
 sg13g2_nor2_1 _2436_ (.A(_1509_),
    .B(net31),
    .Y(_1677_));
 sg13g2_a21oi_1 _2437_ (.A1(net54),
    .A2(net31),
    .Y(_0093_),
    .B1(_1677_));
 sg13g2_buf_1 _2438_ (.A(\ayayayayayaya.b[11] ),
    .X(_1678_));
 sg13g2_inv_2 _2439_ (.Y(_1679_),
    .A(net184));
 sg13g2_buf_1 _2440_ (.A(_1679_),
    .X(_1680_));
 sg13g2_buf_1 _2441_ (.A(net136),
    .X(_1681_));
 sg13g2_nor2_1 _2442_ (.A(_1570_),
    .B(net31),
    .Y(_1682_));
 sg13g2_a21oi_1 _2443_ (.A1(net90),
    .A2(net31),
    .Y(_0094_),
    .B1(_1682_));
 sg13g2_buf_1 _2444_ (.A(\ayayayayayaya.b[12] ),
    .X(_1683_));
 sg13g2_inv_1 _2445_ (.Y(_1684_),
    .A(net183));
 sg13g2_buf_1 _2446_ (.A(_1684_),
    .X(_1685_));
 sg13g2_buf_1 _2447_ (.A(net135),
    .X(_1686_));
 sg13g2_nor2_1 _2448_ (.A(_1573_),
    .B(_1675_),
    .Y(_1687_));
 sg13g2_a21oi_1 _2449_ (.A1(net89),
    .A2(net31),
    .Y(_0095_),
    .B1(_1687_));
 sg13g2_buf_2 _2450_ (.A(\ayayayayayaya.b[13] ),
    .X(_1688_));
 sg13g2_inv_1 _2451_ (.Y(_1689_),
    .A(_1688_));
 sg13g2_buf_1 _2452_ (.A(_1689_),
    .X(_1690_));
 sg13g2_buf_1 _2453_ (.A(net134),
    .X(_1691_));
 sg13g2_nor2_1 _2454_ (.A(_1576_),
    .B(_1675_),
    .Y(_1692_));
 sg13g2_a21oi_1 _2455_ (.A1(_1691_),
    .A2(net31),
    .Y(_0096_),
    .B1(_1692_));
 sg13g2_buf_8 _2456_ (.A(\ayayayayayaya.b[14] ),
    .X(_1693_));
 sg13g2_inv_1 _2457_ (.Y(_1694_),
    .A(net182));
 sg13g2_buf_8 _2458_ (.A(_1694_),
    .X(_1695_));
 sg13g2_buf_1 _2459_ (.A(net133),
    .X(_1696_));
 sg13g2_nor2_1 _2460_ (.A(_1580_),
    .B(_1675_),
    .Y(_1697_));
 sg13g2_a21oi_1 _2461_ (.A1(net87),
    .A2(_1676_),
    .Y(_0097_),
    .B1(_1697_));
 sg13g2_buf_8 _2462_ (.A(\ayayayayayaya.b[15] ),
    .X(_1698_));
 sg13g2_inv_2 _2463_ (.Y(_1699_),
    .A(net181));
 sg13g2_buf_1 _2464_ (.A(_1699_),
    .X(_1700_));
 sg13g2_nor2_1 _2465_ (.A(_1584_),
    .B(_1675_),
    .Y(_1701_));
 sg13g2_a21oi_1 _2466_ (.A1(net132),
    .A2(_1676_),
    .Y(_0098_),
    .B1(_1701_));
 sg13g2_buf_1 _2467_ (.A(\ayayayayayaya.b[16] ),
    .X(_1702_));
 sg13g2_inv_2 _2468_ (.Y(_1703_),
    .A(net180));
 sg13g2_buf_1 _2469_ (.A(_1703_),
    .X(_1704_));
 sg13g2_nand2_1 _2470_ (.Y(_1705_),
    .A(net42),
    .B(_1592_));
 sg13g2_buf_1 _2471_ (.A(_1705_),
    .X(_1706_));
 sg13g2_buf_1 _2472_ (.A(_1706_),
    .X(_1707_));
 sg13g2_nor2_1 _2473_ (.A(_1260_),
    .B(net30),
    .Y(_1708_));
 sg13g2_a21oi_1 _2474_ (.A1(net131),
    .A2(net30),
    .Y(_0099_),
    .B1(_1708_));
 sg13g2_buf_2 _2475_ (.A(\ayayayayayaya.b[17] ),
    .X(_1709_));
 sg13g2_inv_2 _2476_ (.Y(_1710_),
    .A(_1709_));
 sg13g2_buf_1 _2477_ (.A(_1710_),
    .X(_1711_));
 sg13g2_nor2_1 _2478_ (.A(_1599_),
    .B(net30),
    .Y(_1712_));
 sg13g2_a21oi_1 _2479_ (.A1(net130),
    .A2(net30),
    .Y(_0100_),
    .B1(_1712_));
 sg13g2_buf_2 _2480_ (.A(\ayayayayayaya.b[18] ),
    .X(_1713_));
 sg13g2_inv_2 _2481_ (.Y(_1714_),
    .A(_1713_));
 sg13g2_buf_1 _2482_ (.A(_1714_),
    .X(_1715_));
 sg13g2_nor2_1 _2483_ (.A(_1509_),
    .B(_1706_),
    .Y(_1716_));
 sg13g2_a21oi_1 _2484_ (.A1(net129),
    .A2(net30),
    .Y(_0101_),
    .B1(_1716_));
 sg13g2_buf_2 _2485_ (.A(\ayayayayayaya.b[19] ),
    .X(_1717_));
 sg13g2_inv_1 _2486_ (.Y(_1718_),
    .A(_1717_));
 sg13g2_buf_1 _2487_ (.A(_1718_),
    .X(_1719_));
 sg13g2_nor2_1 _2488_ (.A(_1570_),
    .B(_1706_),
    .Y(_1720_));
 sg13g2_a21oi_1 _2489_ (.A1(_1719_),
    .A2(_1707_),
    .Y(_0102_),
    .B1(_1720_));
 sg13g2_buf_1 _2490_ (.A(\ayayayayayaya.b[1] ),
    .X(_1721_));
 sg13g2_inv_1 _2491_ (.Y(_1722_),
    .A(_1721_));
 sg13g2_buf_1 _2492_ (.A(net170),
    .X(_1723_));
 sg13g2_buf_1 _2493_ (.A(net127),
    .X(_1724_));
 sg13g2_nor2_1 _2494_ (.A(_1599_),
    .B(net32),
    .Y(_1725_));
 sg13g2_a21oi_1 _2495_ (.A1(net86),
    .A2(net32),
    .Y(_0103_),
    .B1(_1725_));
 sg13g2_buf_1 _2496_ (.A(\ayayayayayaya.b[20] ),
    .X(_1726_));
 sg13g2_inv_1 _2497_ (.Y(_1727_),
    .A(_1726_));
 sg13g2_buf_1 _2498_ (.A(_1727_),
    .X(_1728_));
 sg13g2_nor2_1 _2499_ (.A(_1573_),
    .B(_1706_),
    .Y(_1729_));
 sg13g2_a21oi_1 _2500_ (.A1(net126),
    .A2(net30),
    .Y(_0104_),
    .B1(_1729_));
 sg13g2_buf_1 _2501_ (.A(\ayayayayayaya.b[21] ),
    .X(_1730_));
 sg13g2_inv_1 _2502_ (.Y(_1731_),
    .A(_1730_));
 sg13g2_buf_1 _2503_ (.A(_1731_),
    .X(_1732_));
 sg13g2_nor2_1 _2504_ (.A(_1576_),
    .B(_1706_),
    .Y(_1733_));
 sg13g2_a21oi_1 _2505_ (.A1(net125),
    .A2(net30),
    .Y(_0105_),
    .B1(_1733_));
 sg13g2_buf_1 _2506_ (.A(\ayayayayayaya.b[22] ),
    .X(_1734_));
 sg13g2_inv_2 _2507_ (.Y(_1735_),
    .A(_1734_));
 sg13g2_nor2_1 _2508_ (.A(_1580_),
    .B(_1706_),
    .Y(_1736_));
 sg13g2_a21oi_1 _2509_ (.A1(net169),
    .A2(_1707_),
    .Y(_0106_),
    .B1(_1736_));
 sg13g2_inv_2 _2510_ (.Y(_1737_),
    .A(\ayayayayayaya.b[23] ));
 sg13g2_nor2_1 _2511_ (.A(_1584_),
    .B(_1706_),
    .Y(_1738_));
 sg13g2_a21oi_1 _2512_ (.A1(net179),
    .A2(net30),
    .Y(_0107_),
    .B1(_1738_));
 sg13g2_nand2_1 _2513_ (.Y(_1739_),
    .A(net42),
    .B(_1621_));
 sg13g2_buf_2 _2514_ (.A(_1739_),
    .X(_1740_));
 sg13g2_buf_1 _2515_ (.A(_1740_),
    .X(_1741_));
 sg13g2_buf_1 _2516_ (.A(\ayayayayayaya.b[24] ),
    .X(_1742_));
 sg13g2_nand2_1 _2517_ (.Y(_1743_),
    .A(net29),
    .B(net178));
 sg13g2_o21ai_1 _2518_ (.B1(_1743_),
    .Y(_0108_),
    .A1(_1271_),
    .A2(net29));
 sg13g2_buf_1 _2519_ (.A(\ayayayayayaya.b[25] ),
    .X(_1744_));
 sg13g2_nand2_1 _2520_ (.Y(_1745_),
    .A(_1741_),
    .B(net177));
 sg13g2_o21ai_1 _2521_ (.B1(_1745_),
    .Y(_0109_),
    .A1(_1605_),
    .A2(net29));
 sg13g2_buf_1 _2522_ (.A(\ayayayayayaya.b[26] ),
    .X(_1746_));
 sg13g2_nand2_1 _2523_ (.Y(_1747_),
    .A(_1740_),
    .B(net176));
 sg13g2_o21ai_1 _2524_ (.B1(_1747_),
    .Y(_0110_),
    .A1(_1520_),
    .A2(_1741_));
 sg13g2_buf_2 _2525_ (.A(\ayayayayayaya.b[27] ),
    .X(_1748_));
 sg13g2_nand2_1 _2526_ (.Y(_1749_),
    .A(_1740_),
    .B(_1748_));
 sg13g2_o21ai_1 _2527_ (.B1(_1749_),
    .Y(_0111_),
    .A1(_1571_),
    .A2(net29));
 sg13g2_buf_2 _2528_ (.A(\ayayayayayaya.b[28] ),
    .X(_1750_));
 sg13g2_nand2_1 _2529_ (.Y(_1751_),
    .A(_1740_),
    .B(_1750_));
 sg13g2_o21ai_1 _2530_ (.B1(_1751_),
    .Y(_0112_),
    .A1(_1574_),
    .A2(net29));
 sg13g2_buf_8 _2531_ (.A(\ayayayayayaya.b[29] ),
    .X(_1752_));
 sg13g2_nand2_1 _2532_ (.Y(_1753_),
    .A(_1740_),
    .B(_1752_));
 sg13g2_o21ai_1 _2533_ (.B1(_1753_),
    .Y(_0113_),
    .A1(_1577_),
    .A2(net29));
 sg13g2_buf_2 _2534_ (.A(\ayayayayayaya.b[2] ),
    .X(_1754_));
 sg13g2_inv_2 _2535_ (.Y(_1755_),
    .A(_1754_));
 sg13g2_buf_1 _2536_ (.A(_1755_),
    .X(_1756_));
 sg13g2_buf_1 _2537_ (.A(net124),
    .X(_1757_));
 sg13g2_nor2_1 _2538_ (.A(_1509_),
    .B(_1666_),
    .Y(_1758_));
 sg13g2_a21oi_1 _2539_ (.A1(net85),
    .A2(net32),
    .Y(_0114_),
    .B1(_1758_));
 sg13g2_buf_8 _2540_ (.A(\ayayayayayaya.b[30] ),
    .X(_1759_));
 sg13g2_nand2_1 _2541_ (.Y(_1760_),
    .A(_1740_),
    .B(_1759_));
 sg13g2_o21ai_1 _2542_ (.B1(_1760_),
    .Y(_0115_),
    .A1(_1581_),
    .A2(net29));
 sg13g2_nand2_1 _2543_ (.Y(_1761_),
    .A(_1740_),
    .B(\ayayayayayaya.b[31] ));
 sg13g2_o21ai_1 _2544_ (.B1(_1761_),
    .Y(_0116_),
    .A1(_1585_),
    .A2(net29));
 sg13g2_buf_1 _2545_ (.A(\ayayayayayaya.b[3] ),
    .X(_1762_));
 sg13g2_inv_2 _2546_ (.Y(_1763_),
    .A(_1762_));
 sg13g2_buf_1 _2547_ (.A(net168),
    .X(_1764_));
 sg13g2_buf_1 _2548_ (.A(net123),
    .X(_1765_));
 sg13g2_nor2_1 _2549_ (.A(_1570_),
    .B(_1666_),
    .Y(_1766_));
 sg13g2_a21oi_1 _2550_ (.A1(net84),
    .A2(net32),
    .Y(_0117_),
    .B1(_1766_));
 sg13g2_buf_1 _2551_ (.A(\ayayayayayaya.b[4] ),
    .X(_1767_));
 sg13g2_inv_1 _2552_ (.Y(_1768_),
    .A(_1767_));
 sg13g2_buf_1 _2553_ (.A(_1768_),
    .X(_1769_));
 sg13g2_buf_1 _2554_ (.A(_1769_),
    .X(_1770_));
 sg13g2_buf_1 _2555_ (.A(net83),
    .X(_1771_));
 sg13g2_nor2_1 _2556_ (.A(_1573_),
    .B(_1666_),
    .Y(_1772_));
 sg13g2_a21oi_1 _2557_ (.A1(net53),
    .A2(net32),
    .Y(_0118_),
    .B1(_1772_));
 sg13g2_buf_1 _2558_ (.A(\ayayayayayaya.b[5] ),
    .X(_1773_));
 sg13g2_inv_1 _2559_ (.Y(_1774_),
    .A(_1773_));
 sg13g2_buf_1 _2560_ (.A(net167),
    .X(_1775_));
 sg13g2_buf_1 _2561_ (.A(net121),
    .X(_1776_));
 sg13g2_nor2_1 _2562_ (.A(_1576_),
    .B(_1666_),
    .Y(_1777_));
 sg13g2_a21oi_1 _2563_ (.A1(net82),
    .A2(net32),
    .Y(_0119_),
    .B1(_1777_));
 sg13g2_buf_1 _2564_ (.A(\ayayayayayaya.b[6] ),
    .X(_1778_));
 sg13g2_inv_2 _2565_ (.Y(_1779_),
    .A(_1778_));
 sg13g2_buf_1 _2566_ (.A(_1779_),
    .X(_1780_));
 sg13g2_buf_1 _2567_ (.A(net120),
    .X(_1781_));
 sg13g2_nor2_1 _2568_ (.A(_1580_),
    .B(_1666_),
    .Y(_1782_));
 sg13g2_a21oi_1 _2569_ (.A1(net81),
    .A2(net32),
    .Y(_0120_),
    .B1(_1782_));
 sg13g2_buf_1 _2570_ (.A(\ayayayayayaya.b[7] ),
    .X(_1783_));
 sg13g2_inv_2 _2571_ (.Y(_1784_),
    .A(net174));
 sg13g2_buf_8 _2572_ (.A(_1784_),
    .X(_1785_));
 sg13g2_buf_1 _2573_ (.A(net119),
    .X(_1786_));
 sg13g2_nor2_1 _2574_ (.A(_1584_),
    .B(_1666_),
    .Y(_1787_));
 sg13g2_a21oi_1 _2575_ (.A1(net80),
    .A2(net32),
    .Y(_0121_),
    .B1(_1787_));
 sg13g2_buf_2 _2576_ (.A(\ayayayayayaya.b[8] ),
    .X(_1788_));
 sg13g2_inv_1 _2577_ (.Y(_1789_),
    .A(_1788_));
 sg13g2_buf_1 _2578_ (.A(_1789_),
    .X(_1790_));
 sg13g2_buf_1 _2579_ (.A(net118),
    .X(_1791_));
 sg13g2_buf_1 _2580_ (.A(net79),
    .X(_1792_));
 sg13g2_nor2_1 _2581_ (.A(_1260_),
    .B(_1675_),
    .Y(_1793_));
 sg13g2_a21oi_1 _2582_ (.A1(_1792_),
    .A2(net31),
    .Y(_0122_),
    .B1(_1793_));
 sg13g2_buf_2 _2583_ (.A(\ayayayayayaya.b[9] ),
    .X(_1794_));
 sg13g2_inv_1 _2584_ (.Y(_1795_),
    .A(_1794_));
 sg13g2_buf_8 _2585_ (.A(_1795_),
    .X(_1796_));
 sg13g2_buf_1 _2586_ (.A(_1796_),
    .X(_1797_));
 sg13g2_buf_1 _2587_ (.A(net78),
    .X(_1798_));
 sg13g2_nor2_1 _2588_ (.A(_1599_),
    .B(_1675_),
    .Y(_1799_));
 sg13g2_a21oi_1 _2589_ (.A1(net51),
    .A2(net31),
    .Y(_0123_),
    .B1(_1799_));
 sg13g2_inv_1 _2590_ (.Y(net12),
    .A(net3));
 sg13g2_nand2_1 _2591_ (.Y(_1800_),
    .A(_1642_),
    .B(\ayayayayayaya.b[31] ));
 sg13g2_inv_2 _2592_ (.Y(_1801_),
    .A(_1759_));
 sg13g2_nand2_1 _2593_ (.Y(_1802_),
    .A(_1800_),
    .B(_1801_));
 sg13g2_inv_1 _2594_ (.Y(_1803_),
    .A(_1752_));
 sg13g2_nand2_1 _2595_ (.Y(_1804_),
    .A(_0030_),
    .B(_1759_));
 sg13g2_nand3_1 _2596_ (.B(_1803_),
    .C(_1804_),
    .A(_1802_),
    .Y(_1805_));
 sg13g2_nand2b_1 _2597_ (.Y(_1806_),
    .B(_1752_),
    .A_N(_0029_));
 sg13g2_nand3_1 _2598_ (.B(_1750_),
    .C(_1806_),
    .A(_1805_),
    .Y(_1807_));
 sg13g2_nand3_1 _2599_ (.B(_1752_),
    .C(_1804_),
    .A(_1802_),
    .Y(_1808_));
 sg13g2_inv_1 _2600_ (.Y(_1809_),
    .A(_1750_));
 sg13g2_nor2_1 _2601_ (.A(_1801_),
    .B(_1800_),
    .Y(_1810_));
 sg13g2_nand2_1 _2602_ (.Y(_1811_),
    .A(_1810_),
    .B(_1803_));
 sg13g2_nand3_1 _2603_ (.B(_1809_),
    .C(_1811_),
    .A(_1808_),
    .Y(_1812_));
 sg13g2_nand3_1 _2604_ (.B(_1812_),
    .C(_1748_),
    .A(_1807_),
    .Y(_1813_));
 sg13g2_nand3_1 _2605_ (.B(_1750_),
    .C(_1811_),
    .A(_1808_),
    .Y(_1814_));
 sg13g2_inv_1 _2606_ (.Y(_1815_),
    .A(_1748_));
 sg13g2_nand2_1 _2607_ (.Y(_1816_),
    .A(_1810_),
    .B(_1752_));
 sg13g2_nand2_1 _2608_ (.Y(_1817_),
    .A(_1816_),
    .B(_1809_));
 sg13g2_nand3_1 _2609_ (.B(_1815_),
    .C(_1817_),
    .A(_1814_),
    .Y(_1818_));
 sg13g2_nand3_1 _2610_ (.B(_1818_),
    .C(net176),
    .A(_1813_),
    .Y(_1819_));
 sg13g2_nand3_1 _2611_ (.B(_1748_),
    .C(_1817_),
    .A(_1814_),
    .Y(_1820_));
 sg13g2_inv_1 _2612_ (.Y(_1821_),
    .A(net176));
 sg13g2_nor2_1 _2613_ (.A(_0059_),
    .B(_1816_),
    .Y(_1822_));
 sg13g2_nand2_1 _2614_ (.Y(_1823_),
    .A(_1822_),
    .B(_1815_));
 sg13g2_nand3_1 _2615_ (.B(_1821_),
    .C(_1823_),
    .A(_1820_),
    .Y(_1824_));
 sg13g2_nand3_1 _2616_ (.B(_1824_),
    .C(net177),
    .A(_1819_),
    .Y(_1825_));
 sg13g2_nand3_1 _2617_ (.B(net176),
    .C(_1823_),
    .A(_1820_),
    .Y(_1826_));
 sg13g2_inv_2 _2618_ (.Y(_1827_),
    .A(net177));
 sg13g2_nor3_1 _2619_ (.A(_0059_),
    .B(_0058_),
    .C(_1816_),
    .Y(_1828_));
 sg13g2_inv_1 _2620_ (.Y(_1829_),
    .A(_1828_));
 sg13g2_nand2_1 _2621_ (.Y(_1830_),
    .A(_1829_),
    .B(_1821_));
 sg13g2_nand3_1 _2622_ (.B(_1827_),
    .C(_1830_),
    .A(_1826_),
    .Y(_1831_));
 sg13g2_nand3_1 _2623_ (.B(_1831_),
    .C(net178),
    .A(_1825_),
    .Y(_1832_));
 sg13g2_nand3_1 _2624_ (.B(net177),
    .C(_1830_),
    .A(_1826_),
    .Y(_1833_));
 sg13g2_inv_2 _2625_ (.Y(_1834_),
    .A(\ayayayayayaya.b[24] ));
 sg13g2_nor2_1 _2626_ (.A(_0057_),
    .B(_1829_),
    .Y(_1835_));
 sg13g2_nand2_1 _2627_ (.Y(_1836_),
    .A(_1835_),
    .B(_1827_));
 sg13g2_nand3_1 _2628_ (.B(_1834_),
    .C(_1836_),
    .A(_1833_),
    .Y(_1837_));
 sg13g2_buf_1 _2629_ (.A(\ayayayayayaya.b[23] ),
    .X(_1838_));
 sg13g2_nand3_1 _2630_ (.B(_1837_),
    .C(net173),
    .A(_1832_),
    .Y(_1839_));
 sg13g2_nand3_1 _2631_ (.B(net178),
    .C(_1836_),
    .A(_1833_),
    .Y(_1840_));
 sg13g2_nor3_1 _2632_ (.A(_0057_),
    .B(_0056_),
    .C(_1829_),
    .Y(_1841_));
 sg13g2_inv_1 _2633_ (.Y(_1842_),
    .A(_1841_));
 sg13g2_nand2_1 _2634_ (.Y(_1843_),
    .A(_1842_),
    .B(_1834_));
 sg13g2_nand3_1 _2635_ (.B(net179),
    .C(_1843_),
    .A(_1840_),
    .Y(_1844_));
 sg13g2_buf_1 _2636_ (.A(_1734_),
    .X(_1845_));
 sg13g2_nand3_1 _2637_ (.B(_1844_),
    .C(net166),
    .A(_1839_),
    .Y(_1846_));
 sg13g2_nand3_1 _2638_ (.B(net173),
    .C(_1843_),
    .A(_1840_),
    .Y(_1847_));
 sg13g2_nor2_1 _2639_ (.A(_0055_),
    .B(_1842_),
    .Y(_1848_));
 sg13g2_nand2_1 _2640_ (.Y(_1849_),
    .A(_1848_),
    .B(net179));
 sg13g2_nand3_1 _2641_ (.B(_1735_),
    .C(_1849_),
    .A(_1847_),
    .Y(_1850_));
 sg13g2_nand3_1 _2642_ (.B(_1850_),
    .C(_1730_),
    .A(_1846_),
    .Y(_1851_));
 sg13g2_nand3_1 _2643_ (.B(_1734_),
    .C(_1849_),
    .A(_1847_),
    .Y(_1852_));
 sg13g2_nor3_1 _2644_ (.A(_0055_),
    .B(_0054_),
    .C(_1842_),
    .Y(_1853_));
 sg13g2_inv_1 _2645_ (.Y(_1854_),
    .A(_1853_));
 sg13g2_nand2_1 _2646_ (.Y(_1855_),
    .A(_1854_),
    .B(net169));
 sg13g2_nand3_1 _2647_ (.B(net125),
    .C(_1855_),
    .A(_1852_),
    .Y(_1856_));
 sg13g2_nand3_1 _2648_ (.B(_1856_),
    .C(_1726_),
    .A(_1851_),
    .Y(_1857_));
 sg13g2_nand3_1 _2649_ (.B(_1730_),
    .C(_1855_),
    .A(_1852_),
    .Y(_1858_));
 sg13g2_nor2_1 _2650_ (.A(_0053_),
    .B(_1854_),
    .Y(_1859_));
 sg13g2_nand2_1 _2651_ (.Y(_1860_),
    .A(_1859_),
    .B(_1731_));
 sg13g2_nand3_1 _2652_ (.B(_1727_),
    .C(_1860_),
    .A(_1858_),
    .Y(_1861_));
 sg13g2_nand3_1 _2653_ (.B(_1861_),
    .C(_1717_),
    .A(_1857_),
    .Y(_1862_));
 sg13g2_nand3_1 _2654_ (.B(_1726_),
    .C(_1860_),
    .A(_1858_),
    .Y(_1863_));
 sg13g2_nor3_1 _2655_ (.A(_0053_),
    .B(_0052_),
    .C(_1854_),
    .Y(_1864_));
 sg13g2_inv_1 _2656_ (.Y(_1865_),
    .A(_1864_));
 sg13g2_nand2_1 _2657_ (.Y(_1866_),
    .A(_1865_),
    .B(_1727_));
 sg13g2_nand3_1 _2658_ (.B(_1718_),
    .C(_1866_),
    .A(_1863_),
    .Y(_1867_));
 sg13g2_nand3_1 _2659_ (.B(_1867_),
    .C(_1713_),
    .A(_1862_),
    .Y(_1868_));
 sg13g2_nand3_1 _2660_ (.B(_1717_),
    .C(_1866_),
    .A(_1863_),
    .Y(_1869_));
 sg13g2_nor2_1 _2661_ (.A(_0051_),
    .B(_1865_),
    .Y(_1870_));
 sg13g2_nand2_1 _2662_ (.Y(_1871_),
    .A(_1870_),
    .B(_1718_));
 sg13g2_nand3_1 _2663_ (.B(_1714_),
    .C(_1871_),
    .A(_1869_),
    .Y(_1872_));
 sg13g2_nand3_1 _2664_ (.B(_1872_),
    .C(_1709_),
    .A(_1868_),
    .Y(_1873_));
 sg13g2_nand3_1 _2665_ (.B(_1713_),
    .C(_1871_),
    .A(_1869_),
    .Y(_1874_));
 sg13g2_nor3_1 _2666_ (.A(_0051_),
    .B(_0050_),
    .C(_1865_),
    .Y(_1875_));
 sg13g2_inv_1 _2667_ (.Y(_1876_),
    .A(_1875_));
 sg13g2_nand2_1 _2668_ (.Y(_1877_),
    .A(_1876_),
    .B(_1714_));
 sg13g2_nand3_1 _2669_ (.B(_1710_),
    .C(_1877_),
    .A(_1874_),
    .Y(_1878_));
 sg13g2_nand3_1 _2670_ (.B(_1878_),
    .C(net180),
    .A(_1873_),
    .Y(_1879_));
 sg13g2_nand3_1 _2671_ (.B(_1709_),
    .C(_1877_),
    .A(_1874_),
    .Y(_1880_));
 sg13g2_nor2_1 _2672_ (.A(_0049_),
    .B(_1876_),
    .Y(_1881_));
 sg13g2_nand2_1 _2673_ (.Y(_1882_),
    .A(_1881_),
    .B(_1710_));
 sg13g2_nand3_1 _2674_ (.B(_1703_),
    .C(_1882_),
    .A(_1880_),
    .Y(_1883_));
 sg13g2_nand3_1 _2675_ (.B(_1883_),
    .C(net181),
    .A(_1879_),
    .Y(_1884_));
 sg13g2_nand3_1 _2676_ (.B(net180),
    .C(_1882_),
    .A(_1880_),
    .Y(_1885_));
 sg13g2_nor3_1 _2677_ (.A(_0049_),
    .B(_0048_),
    .C(_1876_),
    .Y(_1886_));
 sg13g2_inv_1 _2678_ (.Y(_1887_),
    .A(_1886_));
 sg13g2_nand2_1 _2679_ (.Y(_1888_),
    .A(_1887_),
    .B(_1703_));
 sg13g2_nand3_1 _2680_ (.B(_1699_),
    .C(_1888_),
    .A(_1885_),
    .Y(_1889_));
 sg13g2_nand3_1 _2681_ (.B(_1889_),
    .C(net182),
    .A(_1884_),
    .Y(_1890_));
 sg13g2_nand3_1 _2682_ (.B(net181),
    .C(_1888_),
    .A(_1885_),
    .Y(_1891_));
 sg13g2_nor2_1 _2683_ (.A(_0047_),
    .B(_1887_),
    .Y(_1892_));
 sg13g2_nand2_1 _2684_ (.Y(_1893_),
    .A(_1892_),
    .B(_1699_));
 sg13g2_nand3_1 _2685_ (.B(net133),
    .C(_1893_),
    .A(_1891_),
    .Y(_1894_));
 sg13g2_nand3_1 _2686_ (.B(_1894_),
    .C(_1688_),
    .A(_1890_),
    .Y(_1895_));
 sg13g2_nand3_1 _2687_ (.B(net182),
    .C(_1893_),
    .A(_1891_),
    .Y(_1896_));
 sg13g2_inv_1 _2688_ (.Y(_1897_),
    .A(_1892_));
 sg13g2_nor2_1 _2689_ (.A(_0046_),
    .B(_1897_),
    .Y(_1898_));
 sg13g2_inv_1 _2690_ (.Y(_1899_),
    .A(_1898_));
 sg13g2_nand2_1 _2691_ (.Y(_1900_),
    .A(_1899_),
    .B(net133));
 sg13g2_nand3_1 _2692_ (.B(_1689_),
    .C(_1900_),
    .A(_1896_),
    .Y(_1901_));
 sg13g2_nand2_1 _2693_ (.Y(_1902_),
    .A(_1895_),
    .B(_1901_));
 sg13g2_nand2_1 _2694_ (.Y(_1903_),
    .A(_1902_),
    .B(net183));
 sg13g2_nand2_1 _2695_ (.Y(_1904_),
    .A(_1896_),
    .B(_1900_));
 sg13g2_buf_1 _2696_ (.A(_1688_),
    .X(_1905_));
 sg13g2_nand2_1 _2697_ (.Y(_1906_),
    .A(_1904_),
    .B(net165));
 sg13g2_nor2_1 _2698_ (.A(_0045_),
    .B(_1899_),
    .Y(_1907_));
 sg13g2_inv_1 _2699_ (.Y(_1908_),
    .A(_1907_));
 sg13g2_nand2_1 _2700_ (.Y(_1909_),
    .A(_1908_),
    .B(net134));
 sg13g2_nand3_1 _2701_ (.B(_1684_),
    .C(_1909_),
    .A(_1906_),
    .Y(_1910_));
 sg13g2_nand2_1 _2702_ (.Y(_1911_),
    .A(_1903_),
    .B(_1910_));
 sg13g2_nand2_1 _2703_ (.Y(_1912_),
    .A(_1911_),
    .B(net136));
 sg13g2_nand3_1 _2704_ (.B(_1812_),
    .C(_1815_),
    .A(_1807_),
    .Y(_1913_));
 sg13g2_nand3_1 _2705_ (.B(_1809_),
    .C(_1806_),
    .A(_1805_),
    .Y(_1914_));
 sg13g2_nand2_1 _2706_ (.Y(_1915_),
    .A(_0028_),
    .B(_1750_));
 sg13g2_nand3_1 _2707_ (.B(_1748_),
    .C(_1915_),
    .A(_1914_),
    .Y(_1916_));
 sg13g2_nand3_1 _2708_ (.B(_1916_),
    .C(net176),
    .A(_1913_),
    .Y(_1917_));
 sg13g2_nand3_1 _2709_ (.B(_1818_),
    .C(_1821_),
    .A(_1813_),
    .Y(_1918_));
 sg13g2_nand3_1 _2710_ (.B(_1918_),
    .C(net177),
    .A(_1917_),
    .Y(_1919_));
 sg13g2_nand3_1 _2711_ (.B(_1824_),
    .C(_1827_),
    .A(_1819_),
    .Y(_1920_));
 sg13g2_nand3_1 _2712_ (.B(_1920_),
    .C(net178),
    .A(_1919_),
    .Y(_1921_));
 sg13g2_nand3_1 _2713_ (.B(_1831_),
    .C(_1834_),
    .A(_1825_),
    .Y(_1922_));
 sg13g2_nand3_1 _2714_ (.B(_1922_),
    .C(net173),
    .A(_1921_),
    .Y(_1923_));
 sg13g2_nand3_1 _2715_ (.B(_1837_),
    .C(_1737_),
    .A(_1832_),
    .Y(_1924_));
 sg13g2_nand3_1 _2716_ (.B(_1924_),
    .C(net166),
    .A(_1923_),
    .Y(_1925_));
 sg13g2_nand3_1 _2717_ (.B(_1844_),
    .C(net169),
    .A(_1839_),
    .Y(_1926_));
 sg13g2_buf_1 _2718_ (.A(_1730_),
    .X(_1927_));
 sg13g2_nand3_1 _2719_ (.B(_1926_),
    .C(net164),
    .A(_1925_),
    .Y(_1928_));
 sg13g2_nand3_1 _2720_ (.B(_1850_),
    .C(_1732_),
    .A(_1846_),
    .Y(_1929_));
 sg13g2_buf_1 _2721_ (.A(_1726_),
    .X(_1930_));
 sg13g2_nand3_1 _2722_ (.B(_1929_),
    .C(net163),
    .A(_1928_),
    .Y(_1931_));
 sg13g2_nand3_1 _2723_ (.B(_1856_),
    .C(net126),
    .A(_1851_),
    .Y(_1932_));
 sg13g2_nand3_1 _2724_ (.B(_1932_),
    .C(_1717_),
    .A(_1931_),
    .Y(_1933_));
 sg13g2_nand3_1 _2725_ (.B(_1861_),
    .C(net128),
    .A(_1857_),
    .Y(_1934_));
 sg13g2_nand3_1 _2726_ (.B(_1934_),
    .C(_1713_),
    .A(_1933_),
    .Y(_1935_));
 sg13g2_nand3_1 _2727_ (.B(_1867_),
    .C(_1714_),
    .A(_1862_),
    .Y(_1936_));
 sg13g2_nand3_1 _2728_ (.B(_1936_),
    .C(_1709_),
    .A(_1935_),
    .Y(_1937_));
 sg13g2_nand3_1 _2729_ (.B(_1872_),
    .C(_1710_),
    .A(_1868_),
    .Y(_1938_));
 sg13g2_nand3_1 _2730_ (.B(_1938_),
    .C(net180),
    .A(_1937_),
    .Y(_1939_));
 sg13g2_nand3_1 _2731_ (.B(_1878_),
    .C(_1703_),
    .A(_1873_),
    .Y(_1940_));
 sg13g2_nand3_1 _2732_ (.B(_1940_),
    .C(_1698_),
    .A(_1939_),
    .Y(_1941_));
 sg13g2_nand3_1 _2733_ (.B(_1883_),
    .C(_1699_),
    .A(_1879_),
    .Y(_1942_));
 sg13g2_nand3_1 _2734_ (.B(_1942_),
    .C(net182),
    .A(_1941_),
    .Y(_1943_));
 sg13g2_nand3_1 _2735_ (.B(_1889_),
    .C(net133),
    .A(_1884_),
    .Y(_1944_));
 sg13g2_nand3_1 _2736_ (.B(_1944_),
    .C(net165),
    .A(_1943_),
    .Y(_1945_));
 sg13g2_nand3_1 _2737_ (.B(_1894_),
    .C(net134),
    .A(_1890_),
    .Y(_1946_));
 sg13g2_nand3_1 _2738_ (.B(_1946_),
    .C(_1683_),
    .A(_1945_),
    .Y(_1947_));
 sg13g2_nand3_1 _2739_ (.B(_1901_),
    .C(_1684_),
    .A(_1895_),
    .Y(_1948_));
 sg13g2_nand3_1 _2740_ (.B(_1948_),
    .C(net184),
    .A(_1947_),
    .Y(_1949_));
 sg13g2_nand2_1 _2741_ (.Y(_1950_),
    .A(_1912_),
    .B(_1949_));
 sg13g2_nand2_1 _2742_ (.Y(_1951_),
    .A(_1950_),
    .B(net185));
 sg13g2_nand2_1 _2743_ (.Y(_1952_),
    .A(_1911_),
    .B(net184));
 sg13g2_nand3_1 _2744_ (.B(net165),
    .C(_1900_),
    .A(_1896_),
    .Y(_1953_));
 sg13g2_buf_1 _2745_ (.A(net183),
    .X(_1954_));
 sg13g2_nand2_1 _2746_ (.Y(_1955_),
    .A(_1907_),
    .B(net134));
 sg13g2_nand3_1 _2747_ (.B(net162),
    .C(_1955_),
    .A(_1953_),
    .Y(_1956_));
 sg13g2_nor2_1 _2748_ (.A(_0044_),
    .B(_1908_),
    .Y(_1957_));
 sg13g2_inv_1 _2749_ (.Y(_1958_),
    .A(_1957_));
 sg13g2_nand2_1 _2750_ (.Y(_1959_),
    .A(_1958_),
    .B(net135));
 sg13g2_nand3_1 _2751_ (.B(_1679_),
    .C(_1959_),
    .A(_1956_),
    .Y(_1960_));
 sg13g2_nand2_1 _2752_ (.Y(_1961_),
    .A(_1952_),
    .B(_1960_));
 sg13g2_nand2_1 _2753_ (.Y(_1962_),
    .A(_1961_),
    .B(net137));
 sg13g2_nand2_1 _2754_ (.Y(_1963_),
    .A(_1951_),
    .B(_1962_));
 sg13g2_buf_1 _2755_ (.A(_1794_),
    .X(_1964_));
 sg13g2_nand2_1 _2756_ (.Y(_1965_),
    .A(_1963_),
    .B(_1964_));
 sg13g2_nand3_1 _2757_ (.B(_1901_),
    .C(_1683_),
    .A(_1895_),
    .Y(_1966_));
 sg13g2_nand3_1 _2758_ (.B(_1684_),
    .C(_1955_),
    .A(_1953_),
    .Y(_1967_));
 sg13g2_nand2_1 _2759_ (.Y(_1968_),
    .A(_1966_),
    .B(_1967_));
 sg13g2_nand2_1 _2760_ (.Y(_1969_),
    .A(_1968_),
    .B(_1678_));
 sg13g2_nand3_1 _2761_ (.B(net162),
    .C(_1909_),
    .A(_1906_),
    .Y(_1970_));
 sg13g2_nand2_1 _2762_ (.Y(_1971_),
    .A(_1957_),
    .B(net135));
 sg13g2_nand3_1 _2763_ (.B(_1679_),
    .C(_1971_),
    .A(_1970_),
    .Y(_1972_));
 sg13g2_nand2_1 _2764_ (.Y(_1973_),
    .A(_1969_),
    .B(_1972_));
 sg13g2_buf_1 _2765_ (.A(net185),
    .X(_1974_));
 sg13g2_nand2_1 _2766_ (.Y(_1975_),
    .A(_1973_),
    .B(net160));
 sg13g2_nand3_1 _2767_ (.B(_1678_),
    .C(_1959_),
    .A(_1956_),
    .Y(_1976_));
 sg13g2_nor2_1 _2768_ (.A(_0043_),
    .B(_1958_),
    .Y(_1977_));
 sg13g2_nand2_1 _2769_ (.Y(_1978_),
    .A(_1977_),
    .B(_1679_));
 sg13g2_nand3_1 _2770_ (.B(net137),
    .C(_1978_),
    .A(_1976_),
    .Y(_1979_));
 sg13g2_nand3_1 _2771_ (.B(net117),
    .C(_1979_),
    .A(_1975_),
    .Y(_1980_));
 sg13g2_nand2_1 _2772_ (.Y(_1981_),
    .A(_1965_),
    .B(_1980_));
 sg13g2_nand2_1 _2773_ (.Y(_1982_),
    .A(_1981_),
    .B(net118));
 sg13g2_nand2_1 _2774_ (.Y(_1983_),
    .A(_1963_),
    .B(net117));
 sg13g2_nand2_1 _2775_ (.Y(_1984_),
    .A(_1947_),
    .B(_1948_));
 sg13g2_buf_1 _2776_ (.A(net184),
    .X(_1985_));
 sg13g2_nand2_1 _2777_ (.Y(_1986_),
    .A(_1984_),
    .B(net159));
 sg13g2_nand2_1 _2778_ (.Y(_1987_),
    .A(_1968_),
    .B(_1679_));
 sg13g2_nand2_1 _2779_ (.Y(_1988_),
    .A(_1986_),
    .B(_1987_));
 sg13g2_nand2_1 _2780_ (.Y(_1989_),
    .A(_1988_),
    .B(net91));
 sg13g2_nand3_1 _2781_ (.B(_1918_),
    .C(_1827_),
    .A(_1917_),
    .Y(_1990_));
 sg13g2_nand3_1 _2782_ (.B(_1916_),
    .C(_1821_),
    .A(_1913_),
    .Y(_1991_));
 sg13g2_nand3_1 _2783_ (.B(_1815_),
    .C(_1915_),
    .A(_1914_),
    .Y(_1992_));
 sg13g2_nand2b_1 _2784_ (.Y(_1993_),
    .B(_1748_),
    .A_N(_0027_));
 sg13g2_nand3_1 _2785_ (.B(net176),
    .C(_1993_),
    .A(_1992_),
    .Y(_1994_));
 sg13g2_nand3_1 _2786_ (.B(_1994_),
    .C(net177),
    .A(_1991_),
    .Y(_1995_));
 sg13g2_nand3_1 _2787_ (.B(_1995_),
    .C(net178),
    .A(_1990_),
    .Y(_1996_));
 sg13g2_nand3_1 _2788_ (.B(_1920_),
    .C(_1834_),
    .A(_1919_),
    .Y(_1997_));
 sg13g2_nand3_1 _2789_ (.B(_1997_),
    .C(net173),
    .A(_1996_),
    .Y(_1998_));
 sg13g2_nand3_1 _2790_ (.B(_1922_),
    .C(net179),
    .A(_1921_),
    .Y(_1999_));
 sg13g2_nand3_1 _2791_ (.B(_1999_),
    .C(net166),
    .A(_1998_),
    .Y(_2000_));
 sg13g2_nand3_1 _2792_ (.B(_1924_),
    .C(_1735_),
    .A(_1923_),
    .Y(_2001_));
 sg13g2_nand3_1 _2793_ (.B(_2001_),
    .C(net164),
    .A(_2000_),
    .Y(_2002_));
 sg13g2_nand3_1 _2794_ (.B(_1926_),
    .C(net125),
    .A(_1925_),
    .Y(_2003_));
 sg13g2_nand3_1 _2795_ (.B(_2003_),
    .C(net163),
    .A(_2002_),
    .Y(_2004_));
 sg13g2_nand3_1 _2796_ (.B(_1929_),
    .C(_1728_),
    .A(_1928_),
    .Y(_2005_));
 sg13g2_buf_1 _2797_ (.A(_1717_),
    .X(_2006_));
 sg13g2_nand3_1 _2798_ (.B(_2005_),
    .C(net158),
    .A(_2004_),
    .Y(_2007_));
 sg13g2_nand3_1 _2799_ (.B(_1932_),
    .C(net128),
    .A(_1931_),
    .Y(_2008_));
 sg13g2_buf_1 _2800_ (.A(_1713_),
    .X(_2009_));
 sg13g2_nand3_1 _2801_ (.B(_2008_),
    .C(net157),
    .A(_2007_),
    .Y(_2010_));
 sg13g2_nand3_1 _2802_ (.B(_1934_),
    .C(_1714_),
    .A(_1933_),
    .Y(_2011_));
 sg13g2_nand3_1 _2803_ (.B(_2011_),
    .C(_1709_),
    .A(_2010_),
    .Y(_2012_));
 sg13g2_nand3_1 _2804_ (.B(_1936_),
    .C(_1710_),
    .A(_1935_),
    .Y(_2013_));
 sg13g2_nand3_1 _2805_ (.B(_2013_),
    .C(_1702_),
    .A(_2012_),
    .Y(_2014_));
 sg13g2_nand3_1 _2806_ (.B(_1938_),
    .C(_1703_),
    .A(_1937_),
    .Y(_2015_));
 sg13g2_nand3_1 _2807_ (.B(_2015_),
    .C(_1698_),
    .A(_2014_),
    .Y(_2016_));
 sg13g2_nand3_1 _2808_ (.B(_1940_),
    .C(_1699_),
    .A(_1939_),
    .Y(_2017_));
 sg13g2_nand3_1 _2809_ (.B(_2017_),
    .C(_1693_),
    .A(_2016_),
    .Y(_2018_));
 sg13g2_nand3_1 _2810_ (.B(_1942_),
    .C(net133),
    .A(_1941_),
    .Y(_2019_));
 sg13g2_nand3_1 _2811_ (.B(_2019_),
    .C(net165),
    .A(_2018_),
    .Y(_2020_));
 sg13g2_nand3_1 _2812_ (.B(_1944_),
    .C(_1690_),
    .A(_1943_),
    .Y(_2021_));
 sg13g2_nand3_1 _2813_ (.B(_2021_),
    .C(_1954_),
    .A(_2020_),
    .Y(_2022_));
 sg13g2_nand3_1 _2814_ (.B(_1946_),
    .C(net135),
    .A(_1945_),
    .Y(_2023_));
 sg13g2_nand3_1 _2815_ (.B(_2023_),
    .C(net159),
    .A(_2022_),
    .Y(_2024_));
 sg13g2_nand3_1 _2816_ (.B(_1948_),
    .C(net136),
    .A(_1947_),
    .Y(_2025_));
 sg13g2_nand3_1 _2817_ (.B(_2025_),
    .C(net160),
    .A(_2024_),
    .Y(_2026_));
 sg13g2_nand3_1 _2818_ (.B(_2026_),
    .C(net161),
    .A(_1989_),
    .Y(_2027_));
 sg13g2_nand2_1 _2819_ (.Y(_2028_),
    .A(_1983_),
    .B(_2027_));
 sg13g2_buf_8 _2820_ (.A(_1788_),
    .X(_2029_));
 sg13g2_nand2_1 _2821_ (.Y(_2030_),
    .A(_2028_),
    .B(_2029_));
 sg13g2_nand2_1 _2822_ (.Y(_2031_),
    .A(_1982_),
    .B(_2030_));
 sg13g2_buf_8 _2823_ (.A(net174),
    .X(_2032_));
 sg13g2_nand2_1 _2824_ (.Y(_2033_),
    .A(_2031_),
    .B(_2032_));
 sg13g2_nand2_1 _2825_ (.Y(_2034_),
    .A(_1981_),
    .B(net156));
 sg13g2_nand2_1 _2826_ (.Y(_2035_),
    .A(_1961_),
    .B(_1669_));
 sg13g2_nand2_1 _2827_ (.Y(_2036_),
    .A(_1976_),
    .B(_1978_));
 sg13g2_nand2_1 _2828_ (.Y(_2037_),
    .A(_2036_),
    .B(net137));
 sg13g2_nand3_1 _2829_ (.B(net161),
    .C(_2037_),
    .A(_2035_),
    .Y(_2038_));
 sg13g2_nand3_1 _2830_ (.B(net185),
    .C(_1978_),
    .A(_1976_),
    .Y(_2039_));
 sg13g2_nor3_1 _2831_ (.A(_0043_),
    .B(_0042_),
    .C(_1958_),
    .Y(_2040_));
 sg13g2_inv_1 _2832_ (.Y(_2041_),
    .A(_2040_));
 sg13g2_nand2_1 _2833_ (.Y(_2042_),
    .A(_2041_),
    .B(net137));
 sg13g2_nand2_1 _2834_ (.Y(_2043_),
    .A(_2039_),
    .B(_2042_));
 sg13g2_nand2_1 _2835_ (.Y(_2044_),
    .A(_2043_),
    .B(net78));
 sg13g2_nand3_1 _2836_ (.B(net118),
    .C(_2044_),
    .A(_2038_),
    .Y(_2045_));
 sg13g2_nand2_1 _2837_ (.Y(_2046_),
    .A(_2034_),
    .B(_2045_));
 sg13g2_nand2_1 _2838_ (.Y(_2047_),
    .A(_2046_),
    .B(net119));
 sg13g2_nand2_1 _2839_ (.Y(_2048_),
    .A(_2033_),
    .B(_2047_));
 sg13g2_nand2_1 _2840_ (.Y(_2049_),
    .A(_2048_),
    .B(net120));
 sg13g2_nand2_1 _2841_ (.Y(_2050_),
    .A(_2031_),
    .B(net119));
 sg13g2_nand3_1 _2842_ (.B(_2026_),
    .C(net78),
    .A(_1989_),
    .Y(_2051_));
 sg13g2_nand3_1 _2843_ (.B(_1997_),
    .C(net179),
    .A(_1996_),
    .Y(_2052_));
 sg13g2_nand3_1 _2844_ (.B(_1995_),
    .C(_1834_),
    .A(_1990_),
    .Y(_2053_));
 sg13g2_nand3_1 _2845_ (.B(_1994_),
    .C(_1827_),
    .A(_1991_),
    .Y(_2054_));
 sg13g2_nand3_1 _2846_ (.B(_1821_),
    .C(_1993_),
    .A(_1992_),
    .Y(_2055_));
 sg13g2_nand2_1 _2847_ (.Y(_2056_),
    .A(_0026_),
    .B(_1746_));
 sg13g2_nand3_1 _2848_ (.B(net177),
    .C(_2056_),
    .A(_2055_),
    .Y(_2057_));
 sg13g2_nand3_1 _2849_ (.B(_2057_),
    .C(_1742_),
    .A(_2054_),
    .Y(_2058_));
 sg13g2_nand3_1 _2850_ (.B(_2058_),
    .C(net173),
    .A(_2053_),
    .Y(_2059_));
 sg13g2_nand3_1 _2851_ (.B(_2059_),
    .C(net166),
    .A(_2052_),
    .Y(_2060_));
 sg13g2_nand3_1 _2852_ (.B(_1999_),
    .C(net169),
    .A(_1998_),
    .Y(_2061_));
 sg13g2_nand3_1 _2853_ (.B(_2061_),
    .C(net164),
    .A(_2060_),
    .Y(_2062_));
 sg13g2_nand3_1 _2854_ (.B(_2001_),
    .C(_1732_),
    .A(_2000_),
    .Y(_2063_));
 sg13g2_nand3_1 _2855_ (.B(_2063_),
    .C(_1930_),
    .A(_2062_),
    .Y(_2064_));
 sg13g2_nand3_1 _2856_ (.B(_2003_),
    .C(net126),
    .A(_2002_),
    .Y(_2065_));
 sg13g2_nand3_1 _2857_ (.B(_2065_),
    .C(net158),
    .A(_2064_),
    .Y(_2066_));
 sg13g2_nand3_1 _2858_ (.B(_2005_),
    .C(net128),
    .A(_2004_),
    .Y(_2067_));
 sg13g2_nand3_1 _2859_ (.B(_2067_),
    .C(_2009_),
    .A(_2066_),
    .Y(_2068_));
 sg13g2_nand3_1 _2860_ (.B(_2008_),
    .C(net129),
    .A(_2007_),
    .Y(_2069_));
 sg13g2_nand3_1 _2861_ (.B(_2069_),
    .C(_1709_),
    .A(_2068_),
    .Y(_2070_));
 sg13g2_nand3_1 _2862_ (.B(_2011_),
    .C(_1711_),
    .A(_2010_),
    .Y(_2071_));
 sg13g2_nand3_1 _2863_ (.B(_2071_),
    .C(net180),
    .A(_2070_),
    .Y(_2072_));
 sg13g2_nand3_1 _2864_ (.B(_2013_),
    .C(_1703_),
    .A(_2012_),
    .Y(_2073_));
 sg13g2_nand3_1 _2865_ (.B(_2073_),
    .C(net181),
    .A(_2072_),
    .Y(_2074_));
 sg13g2_nand3_1 _2866_ (.B(_2015_),
    .C(_1699_),
    .A(_2014_),
    .Y(_2075_));
 sg13g2_nand3_1 _2867_ (.B(_2075_),
    .C(net182),
    .A(_2074_),
    .Y(_2076_));
 sg13g2_nand3_1 _2868_ (.B(_2017_),
    .C(net133),
    .A(_2016_),
    .Y(_2077_));
 sg13g2_nand3_1 _2869_ (.B(_2077_),
    .C(net165),
    .A(_2076_),
    .Y(_2078_));
 sg13g2_nand3_1 _2870_ (.B(_2019_),
    .C(net134),
    .A(_2018_),
    .Y(_2079_));
 sg13g2_nand3_1 _2871_ (.B(_2079_),
    .C(net162),
    .A(_2078_),
    .Y(_2080_));
 sg13g2_nand3_1 _2872_ (.B(_2021_),
    .C(net135),
    .A(_2020_),
    .Y(_2081_));
 sg13g2_nand3_1 _2873_ (.B(_2081_),
    .C(_1985_),
    .A(_2080_),
    .Y(_2082_));
 sg13g2_nand3_1 _2874_ (.B(_2023_),
    .C(net136),
    .A(_2022_),
    .Y(_2083_));
 sg13g2_nand3_1 _2875_ (.B(_2083_),
    .C(_1974_),
    .A(_2082_),
    .Y(_2084_));
 sg13g2_nand3_1 _2876_ (.B(_2025_),
    .C(net91),
    .A(_2024_),
    .Y(_2085_));
 sg13g2_buf_1 _2877_ (.A(_1964_),
    .X(_2086_));
 sg13g2_nand3_1 _2878_ (.B(_2085_),
    .C(_2086_),
    .A(_2084_),
    .Y(_2087_));
 sg13g2_nand3_1 _2879_ (.B(_2087_),
    .C(net156),
    .A(_2051_),
    .Y(_2088_));
 sg13g2_nand3_1 _2880_ (.B(_2027_),
    .C(net79),
    .A(_1983_),
    .Y(_2089_));
 sg13g2_nand3_1 _2881_ (.B(_2089_),
    .C(net155),
    .A(_2088_),
    .Y(_2090_));
 sg13g2_nand2_1 _2882_ (.Y(_2091_),
    .A(_2050_),
    .B(_2090_));
 sg13g2_buf_1 _2883_ (.A(_1778_),
    .X(_2092_));
 sg13g2_buf_1 _2884_ (.A(_2092_),
    .X(_2093_));
 sg13g2_nand2_1 _2885_ (.Y(_2094_),
    .A(_2091_),
    .B(net115));
 sg13g2_nand2_1 _2886_ (.Y(_2095_),
    .A(_2049_),
    .B(_2094_));
 sg13g2_buf_1 _2887_ (.A(_1773_),
    .X(_2096_));
 sg13g2_buf_1 _2888_ (.A(net153),
    .X(_2097_));
 sg13g2_buf_1 _2889_ (.A(_2097_),
    .X(_2098_));
 sg13g2_nand2_1 _2890_ (.Y(_2099_),
    .A(_2095_),
    .B(net77));
 sg13g2_nand2_1 _2891_ (.Y(_2100_),
    .A(_2048_),
    .B(net115));
 sg13g2_nand2_1 _2892_ (.Y(_2101_),
    .A(_1988_),
    .B(net185));
 sg13g2_nand2_1 _2893_ (.Y(_2102_),
    .A(_1973_),
    .B(_1671_));
 sg13g2_nand2_1 _2894_ (.Y(_2103_),
    .A(_2101_),
    .B(_2102_));
 sg13g2_nand2_1 _2895_ (.Y(_2104_),
    .A(_2103_),
    .B(net161));
 sg13g2_nand3_1 _2896_ (.B(net117),
    .C(_2037_),
    .A(_2035_),
    .Y(_2105_));
 sg13g2_nand2_1 _2897_ (.Y(_2106_),
    .A(_2104_),
    .B(_2105_));
 sg13g2_nand2_1 _2898_ (.Y(_2107_),
    .A(_2106_),
    .B(net156));
 sg13g2_nand3_1 _2899_ (.B(net161),
    .C(_1979_),
    .A(_1975_),
    .Y(_2108_));
 sg13g2_nand3_1 _2900_ (.B(net117),
    .C(_2042_),
    .A(_2039_),
    .Y(_2109_));
 sg13g2_nand3_1 _2901_ (.B(_1790_),
    .C(_2109_),
    .A(_2108_),
    .Y(_2110_));
 sg13g2_nand2_1 _2902_ (.Y(_2111_),
    .A(_2107_),
    .B(_2110_));
 sg13g2_buf_1 _2903_ (.A(net155),
    .X(_2112_));
 sg13g2_nand2_1 _2904_ (.Y(_2113_),
    .A(_2111_),
    .B(net113));
 sg13g2_nand3_1 _2905_ (.B(net156),
    .C(_2109_),
    .A(_2108_),
    .Y(_2114_));
 sg13g2_nand3_1 _2906_ (.B(net161),
    .C(_2042_),
    .A(_2039_),
    .Y(_2115_));
 sg13g2_nor2_1 _2907_ (.A(_0041_),
    .B(_2041_),
    .Y(_2116_));
 sg13g2_nand2_1 _2908_ (.Y(_2117_),
    .A(_2116_),
    .B(net117));
 sg13g2_nand3_1 _2909_ (.B(net118),
    .C(_2117_),
    .A(_2115_),
    .Y(_2118_));
 sg13g2_nand2_1 _2910_ (.Y(_2119_),
    .A(_2114_),
    .B(_2118_));
 sg13g2_nand2_1 _2911_ (.Y(_2120_),
    .A(_2119_),
    .B(_1785_));
 sg13g2_nand3_1 _2912_ (.B(_2120_),
    .C(net120),
    .A(_2113_),
    .Y(_2121_));
 sg13g2_nand2_1 _2913_ (.Y(_2122_),
    .A(_2100_),
    .B(_2121_));
 sg13g2_nand2_1 _2914_ (.Y(_2123_),
    .A(_2122_),
    .B(net121));
 sg13g2_nand2_1 _2915_ (.Y(_2124_),
    .A(_2099_),
    .B(_2123_));
 sg13g2_buf_1 _2916_ (.A(_1767_),
    .X(_2125_));
 sg13g2_buf_1 _2917_ (.A(_2125_),
    .X(_2126_));
 sg13g2_buf_1 _2918_ (.A(net112),
    .X(_2127_));
 sg13g2_nand2_1 _2919_ (.Y(_2128_),
    .A(_2124_),
    .B(net76));
 sg13g2_nand2_1 _2920_ (.Y(_2129_),
    .A(_2122_),
    .B(net77));
 sg13g2_nand2_1 _2921_ (.Y(_2130_),
    .A(_2046_),
    .B(net155));
 sg13g2_nand3_1 _2922_ (.B(net119),
    .C(_2118_),
    .A(_2114_),
    .Y(_2131_));
 sg13g2_nand3_1 _2923_ (.B(_2093_),
    .C(_2131_),
    .A(_2130_),
    .Y(_2132_));
 sg13g2_nand3_1 _2924_ (.B(net155),
    .C(_2118_),
    .A(_2114_),
    .Y(_2133_));
 sg13g2_nand3_1 _2925_ (.B(net156),
    .C(_2117_),
    .A(_2115_),
    .Y(_2134_));
 sg13g2_nor3_1 _2926_ (.A(_0041_),
    .B(_0040_),
    .C(_2041_),
    .Y(_2135_));
 sg13g2_inv_1 _2927_ (.Y(_2136_),
    .A(_2135_));
 sg13g2_nand2_1 _2928_ (.Y(_2137_),
    .A(_2136_),
    .B(net118));
 sg13g2_nand3_1 _2929_ (.B(net119),
    .C(_2137_),
    .A(_2134_),
    .Y(_2138_));
 sg13g2_nand3_1 _2930_ (.B(net120),
    .C(_2138_),
    .A(_2133_),
    .Y(_2139_));
 sg13g2_nand3_1 _2931_ (.B(net121),
    .C(_2139_),
    .A(_2132_),
    .Y(_2140_));
 sg13g2_nand2_1 _2932_ (.Y(_2141_),
    .A(_2129_),
    .B(_2140_));
 sg13g2_nand2_1 _2933_ (.Y(_2142_),
    .A(_2141_),
    .B(net53));
 sg13g2_nand2_1 _2934_ (.Y(_2143_),
    .A(_2128_),
    .B(_2142_));
 sg13g2_nand2_1 _2935_ (.Y(_2144_),
    .A(_2143_),
    .B(net84));
 sg13g2_nand2_1 _2936_ (.Y(_2145_),
    .A(_2106_),
    .B(_1790_));
 sg13g2_nand3_1 _2937_ (.B(_2027_),
    .C(_2029_),
    .A(_1983_),
    .Y(_2146_));
 sg13g2_nand2_1 _2938_ (.Y(_2147_),
    .A(_2145_),
    .B(_2146_));
 sg13g2_nand2_1 _2939_ (.Y(_2148_),
    .A(_2147_),
    .B(_2032_));
 sg13g2_nand2_1 _2940_ (.Y(_2149_),
    .A(_2111_),
    .B(_1785_));
 sg13g2_nand2_1 _2941_ (.Y(_2150_),
    .A(_2148_),
    .B(_2149_));
 sg13g2_nand2_1 _2942_ (.Y(_2151_),
    .A(_2150_),
    .B(net120));
 sg13g2_nand3_1 _2943_ (.B(_2090_),
    .C(_2093_),
    .A(_2050_),
    .Y(_2152_));
 sg13g2_nand2_1 _2944_ (.Y(_2153_),
    .A(_2151_),
    .B(_2152_));
 sg13g2_nand2_1 _2945_ (.Y(_2154_),
    .A(_2153_),
    .B(_2097_));
 sg13g2_nand2_1 _2946_ (.Y(_2155_),
    .A(_2150_),
    .B(net115));
 sg13g2_nand3_1 _2947_ (.B(_1780_),
    .C(_2131_),
    .A(_2130_),
    .Y(_2156_));
 sg13g2_nand2_1 _2948_ (.Y(_2157_),
    .A(_2155_),
    .B(_2156_));
 sg13g2_nand2_1 _2949_ (.Y(_2158_),
    .A(_2157_),
    .B(_1775_));
 sg13g2_nand2_1 _2950_ (.Y(_2159_),
    .A(_2154_),
    .B(_2158_));
 sg13g2_nand2_1 _2951_ (.Y(_2160_),
    .A(_2159_),
    .B(net53));
 sg13g2_nand2_1 _2952_ (.Y(_2161_),
    .A(_2095_),
    .B(net82));
 sg13g2_nand3_1 _2953_ (.B(_2090_),
    .C(net81),
    .A(_2050_),
    .Y(_2162_));
 sg13g2_nand3_1 _2954_ (.B(_2061_),
    .C(net125),
    .A(_2060_),
    .Y(_2163_));
 sg13g2_nand3_1 _2955_ (.B(_2059_),
    .C(net169),
    .A(_2052_),
    .Y(_2164_));
 sg13g2_nand3_1 _2956_ (.B(_2058_),
    .C(net179),
    .A(_2053_),
    .Y(_2165_));
 sg13g2_nand3_1 _2957_ (.B(_2057_),
    .C(_1834_),
    .A(_2054_),
    .Y(_2166_));
 sg13g2_nand3_1 _2958_ (.B(_1827_),
    .C(_2056_),
    .A(_2055_),
    .Y(_2167_));
 sg13g2_nand2b_1 _2959_ (.Y(_2168_),
    .B(_1744_),
    .A_N(_0025_));
 sg13g2_nand3_1 _2960_ (.B(_1742_),
    .C(_2168_),
    .A(_2167_),
    .Y(_2169_));
 sg13g2_nand3_1 _2961_ (.B(_2169_),
    .C(net173),
    .A(_2166_),
    .Y(_2170_));
 sg13g2_nand3_1 _2962_ (.B(_2170_),
    .C(net166),
    .A(_2165_),
    .Y(_2171_));
 sg13g2_nand3_1 _2963_ (.B(_2171_),
    .C(net164),
    .A(_2164_),
    .Y(_2172_));
 sg13g2_nand3_1 _2964_ (.B(_2172_),
    .C(_1930_),
    .A(_2163_),
    .Y(_2173_));
 sg13g2_nand3_1 _2965_ (.B(_2063_),
    .C(net126),
    .A(_2062_),
    .Y(_2174_));
 sg13g2_nand3_1 _2966_ (.B(_2174_),
    .C(net158),
    .A(_2173_),
    .Y(_2175_));
 sg13g2_nand3_1 _2967_ (.B(_2065_),
    .C(_1719_),
    .A(_2064_),
    .Y(_2176_));
 sg13g2_nand3_1 _2968_ (.B(_2176_),
    .C(net157),
    .A(_2175_),
    .Y(_2177_));
 sg13g2_nand3_1 _2969_ (.B(_2067_),
    .C(net129),
    .A(_2066_),
    .Y(_2178_));
 sg13g2_buf_1 _2970_ (.A(_1709_),
    .X(_2179_));
 sg13g2_nand3_1 _2971_ (.B(_2178_),
    .C(net151),
    .A(_2177_),
    .Y(_2180_));
 sg13g2_nand3_1 _2972_ (.B(_2069_),
    .C(net130),
    .A(_2068_),
    .Y(_2181_));
 sg13g2_nand3_1 _2973_ (.B(_2181_),
    .C(net180),
    .A(_2180_),
    .Y(_2182_));
 sg13g2_nand3_1 _2974_ (.B(_2071_),
    .C(_1704_),
    .A(_2070_),
    .Y(_2183_));
 sg13g2_nand3_1 _2975_ (.B(_2183_),
    .C(net181),
    .A(_2182_),
    .Y(_2184_));
 sg13g2_nand3_1 _2976_ (.B(_2073_),
    .C(_1699_),
    .A(_2072_),
    .Y(_2185_));
 sg13g2_nand3_1 _2977_ (.B(_2185_),
    .C(net182),
    .A(_2184_),
    .Y(_2186_));
 sg13g2_nand3_1 _2978_ (.B(_2075_),
    .C(_1695_),
    .A(_2074_),
    .Y(_2187_));
 sg13g2_nand3_1 _2979_ (.B(_2187_),
    .C(net165),
    .A(_2186_),
    .Y(_2188_));
 sg13g2_nand3_1 _2980_ (.B(_2077_),
    .C(net134),
    .A(_2076_),
    .Y(_2189_));
 sg13g2_nand3_1 _2981_ (.B(_2189_),
    .C(net162),
    .A(_2188_),
    .Y(_2190_));
 sg13g2_nand3_1 _2982_ (.B(_2079_),
    .C(net135),
    .A(_2078_),
    .Y(_2191_));
 sg13g2_nand3_1 _2983_ (.B(_2191_),
    .C(net159),
    .A(_2190_),
    .Y(_2192_));
 sg13g2_nand3_1 _2984_ (.B(_2081_),
    .C(net136),
    .A(_2080_),
    .Y(_2193_));
 sg13g2_nand3_1 _2985_ (.B(_2193_),
    .C(net160),
    .A(_2192_),
    .Y(_2194_));
 sg13g2_nand3_1 _2986_ (.B(_2083_),
    .C(net91),
    .A(_2082_),
    .Y(_2195_));
 sg13g2_nand2_1 _2987_ (.Y(_2196_),
    .A(_2194_),
    .B(_2195_));
 sg13g2_nand2_1 _2988_ (.Y(_2197_),
    .A(_2196_),
    .B(_2086_));
 sg13g2_nand2_1 _2989_ (.Y(_2198_),
    .A(_2084_),
    .B(_2085_));
 sg13g2_nand2_1 _2990_ (.Y(_2199_),
    .A(_2198_),
    .B(net78));
 sg13g2_nand2_1 _2991_ (.Y(_2200_),
    .A(_2197_),
    .B(_2199_));
 sg13g2_buf_1 _2992_ (.A(net156),
    .X(_2201_));
 sg13g2_buf_1 _2993_ (.A(net111),
    .X(_2202_));
 sg13g2_nand2_1 _2994_ (.Y(_2203_),
    .A(_2200_),
    .B(net75));
 sg13g2_nand3_1 _2995_ (.B(_2087_),
    .C(net79),
    .A(_2051_),
    .Y(_2204_));
 sg13g2_buf_1 _2996_ (.A(net155),
    .X(_2205_));
 sg13g2_nand3_1 _2997_ (.B(_2204_),
    .C(net110),
    .A(_2203_),
    .Y(_2206_));
 sg13g2_buf_1 _2998_ (.A(net119),
    .X(_2207_));
 sg13g2_nand3_1 _2999_ (.B(_2089_),
    .C(net74),
    .A(_2088_),
    .Y(_2208_));
 sg13g2_buf_1 _3000_ (.A(net115),
    .X(_2209_));
 sg13g2_nand3_1 _3001_ (.B(_2208_),
    .C(net73),
    .A(_2206_),
    .Y(_2210_));
 sg13g2_buf_1 _3002_ (.A(net114),
    .X(_2211_));
 sg13g2_nand3_1 _3003_ (.B(_2210_),
    .C(net72),
    .A(_2162_),
    .Y(_2212_));
 sg13g2_nand3_1 _3004_ (.B(_2212_),
    .C(net76),
    .A(_2161_),
    .Y(_2213_));
 sg13g2_buf_1 _3005_ (.A(net175),
    .X(_2214_));
 sg13g2_buf_1 _3006_ (.A(net150),
    .X(_2215_));
 sg13g2_buf_1 _3007_ (.A(net109),
    .X(_2216_));
 sg13g2_nand3_1 _3008_ (.B(_2213_),
    .C(net71),
    .A(_2160_),
    .Y(_2217_));
 sg13g2_buf_8 _3009_ (.A(_1754_),
    .X(_2218_));
 sg13g2_buf_1 _3010_ (.A(_2218_),
    .X(_2219_));
 sg13g2_buf_1 _3011_ (.A(net108),
    .X(_2220_));
 sg13g2_nand3_1 _3012_ (.B(_2217_),
    .C(net70),
    .A(_2144_),
    .Y(_2221_));
 sg13g2_nand2_1 _3013_ (.Y(_2222_),
    .A(_2159_),
    .B(net112));
 sg13g2_nand2_1 _3014_ (.Y(_2223_),
    .A(_2157_),
    .B(net114));
 sg13g2_nand2_1 _3015_ (.Y(_2224_),
    .A(_2132_),
    .B(_2139_));
 sg13g2_nand2_1 _3016_ (.Y(_2225_),
    .A(_2224_),
    .B(_1774_));
 sg13g2_nand2_1 _3017_ (.Y(_2226_),
    .A(_2223_),
    .B(_2225_));
 sg13g2_nand2_1 _3018_ (.Y(_2227_),
    .A(_2226_),
    .B(net83));
 sg13g2_nand2_1 _3019_ (.Y(_2228_),
    .A(_2222_),
    .B(_2227_));
 sg13g2_nand2_1 _3020_ (.Y(_2229_),
    .A(_2228_),
    .B(net109));
 sg13g2_nand2_1 _3021_ (.Y(_2230_),
    .A(_2226_),
    .B(_2125_));
 sg13g2_nand3_1 _3022_ (.B(net114),
    .C(_2139_),
    .A(_2132_),
    .Y(_2231_));
 sg13g2_nand3_1 _3023_ (.B(net115),
    .C(_2138_),
    .A(_2133_),
    .Y(_2232_));
 sg13g2_nand3_1 _3024_ (.B(net155),
    .C(_2137_),
    .A(_2134_),
    .Y(_2233_));
 sg13g2_nor2_1 _3025_ (.A(_0039_),
    .B(_2136_),
    .Y(_2234_));
 sg13g2_nand2_1 _3026_ (.Y(_2235_),
    .A(_2234_),
    .B(net119));
 sg13g2_nand3_1 _3027_ (.B(net120),
    .C(_2235_),
    .A(_2233_),
    .Y(_2236_));
 sg13g2_nand3_1 _3028_ (.B(_1774_),
    .C(_2236_),
    .A(_2232_),
    .Y(_2237_));
 sg13g2_nand3_1 _3029_ (.B(net83),
    .C(_2237_),
    .A(_2231_),
    .Y(_2238_));
 sg13g2_nand2_1 _3030_ (.Y(_2239_),
    .A(_2230_),
    .B(_2238_));
 sg13g2_nand2_1 _3031_ (.Y(_2240_),
    .A(_2239_),
    .B(net123));
 sg13g2_nand2_1 _3032_ (.Y(_2241_),
    .A(_2229_),
    .B(_2240_));
 sg13g2_nand2_1 _3033_ (.Y(_2242_),
    .A(_2241_),
    .B(net85));
 sg13g2_nand3_1 _3034_ (.B(_2242_),
    .C(net86),
    .A(_2221_),
    .Y(_2243_));
 sg13g2_nand3_1 _3035_ (.B(_2217_),
    .C(net85),
    .A(_2144_),
    .Y(_2244_));
 sg13g2_nand3_1 _3036_ (.B(_2213_),
    .C(net84),
    .A(_2160_),
    .Y(_2245_));
 sg13g2_nand3_1 _3037_ (.B(_2212_),
    .C(net53),
    .A(_2161_),
    .Y(_2246_));
 sg13g2_buf_1 _3038_ (.A(net121),
    .X(_2247_));
 sg13g2_nand3_1 _3039_ (.B(_2210_),
    .C(net69),
    .A(_2162_),
    .Y(_2248_));
 sg13g2_nand3_1 _3040_ (.B(_2174_),
    .C(net128),
    .A(_2173_),
    .Y(_2249_));
 sg13g2_nand3_1 _3041_ (.B(_2172_),
    .C(net126),
    .A(_2163_),
    .Y(_2250_));
 sg13g2_nand3_1 _3042_ (.B(_2171_),
    .C(net125),
    .A(_2164_),
    .Y(_2251_));
 sg13g2_nand3_1 _3043_ (.B(_2170_),
    .C(net169),
    .A(_2165_),
    .Y(_2252_));
 sg13g2_nand3_1 _3044_ (.B(_2169_),
    .C(net179),
    .A(_2166_),
    .Y(_2253_));
 sg13g2_nand3_1 _3045_ (.B(_1834_),
    .C(_2168_),
    .A(_2167_),
    .Y(_2254_));
 sg13g2_nand2_1 _3046_ (.Y(_2255_),
    .A(_0024_),
    .B(net178));
 sg13g2_nand3_1 _3047_ (.B(_1838_),
    .C(_2255_),
    .A(_2254_),
    .Y(_2256_));
 sg13g2_nand3_1 _3048_ (.B(_2256_),
    .C(net166),
    .A(_2253_),
    .Y(_0124_));
 sg13g2_nand3_1 _3049_ (.B(_0124_),
    .C(net164),
    .A(_2252_),
    .Y(_0125_));
 sg13g2_nand3_1 _3050_ (.B(_0125_),
    .C(net163),
    .A(_2251_),
    .Y(_0126_));
 sg13g2_nand3_1 _3051_ (.B(_0126_),
    .C(net158),
    .A(_2250_),
    .Y(_0127_));
 sg13g2_nand3_1 _3052_ (.B(_0127_),
    .C(net157),
    .A(_2249_),
    .Y(_0128_));
 sg13g2_nand3_1 _3053_ (.B(_2176_),
    .C(_1715_),
    .A(_2175_),
    .Y(_0129_));
 sg13g2_nand3_1 _3054_ (.B(_0129_),
    .C(net151),
    .A(_0128_),
    .Y(_0130_));
 sg13g2_nand3_1 _3055_ (.B(_2178_),
    .C(_1711_),
    .A(_2177_),
    .Y(_0131_));
 sg13g2_buf_1 _3056_ (.A(net180),
    .X(_0132_));
 sg13g2_nand3_1 _3057_ (.B(_0131_),
    .C(net148),
    .A(_0130_),
    .Y(_0133_));
 sg13g2_nand3_1 _3058_ (.B(_2181_),
    .C(_1704_),
    .A(_2180_),
    .Y(_0134_));
 sg13g2_nand3_1 _3059_ (.B(_0134_),
    .C(net181),
    .A(_0133_),
    .Y(_0135_));
 sg13g2_nand3_1 _3060_ (.B(_2183_),
    .C(net132),
    .A(_2182_),
    .Y(_0136_));
 sg13g2_nand3_1 _3061_ (.B(_0136_),
    .C(net182),
    .A(_0135_),
    .Y(_0137_));
 sg13g2_nand3_1 _3062_ (.B(_2185_),
    .C(_1695_),
    .A(_2184_),
    .Y(_0138_));
 sg13g2_nand3_1 _3063_ (.B(_0138_),
    .C(net165),
    .A(_0137_),
    .Y(_0139_));
 sg13g2_nand3_1 _3064_ (.B(_2187_),
    .C(_1690_),
    .A(_2186_),
    .Y(_0140_));
 sg13g2_nand3_1 _3065_ (.B(_0140_),
    .C(net162),
    .A(_0139_),
    .Y(_0141_));
 sg13g2_nand3_1 _3066_ (.B(_2189_),
    .C(net135),
    .A(_2188_),
    .Y(_0142_));
 sg13g2_nand3_1 _3067_ (.B(_0142_),
    .C(net159),
    .A(_0141_),
    .Y(_0143_));
 sg13g2_nand3_1 _3068_ (.B(_2191_),
    .C(net136),
    .A(_2190_),
    .Y(_0144_));
 sg13g2_nand3_1 _3069_ (.B(_0144_),
    .C(net160),
    .A(_0143_),
    .Y(_0145_));
 sg13g2_nand3_1 _3070_ (.B(_2193_),
    .C(net91),
    .A(_2192_),
    .Y(_0146_));
 sg13g2_nand3_1 _3071_ (.B(_0146_),
    .C(net116),
    .A(_0145_),
    .Y(_0147_));
 sg13g2_nand3_1 _3072_ (.B(_2195_),
    .C(net78),
    .A(_2194_),
    .Y(_0148_));
 sg13g2_nand2_1 _3073_ (.Y(_0149_),
    .A(_0147_),
    .B(_0148_));
 sg13g2_nand2_1 _3074_ (.Y(_0150_),
    .A(_0149_),
    .B(_2201_));
 sg13g2_nand3_1 _3075_ (.B(_2199_),
    .C(net79),
    .A(_2197_),
    .Y(_0151_));
 sg13g2_nand2_1 _3076_ (.Y(_0152_),
    .A(_0150_),
    .B(_0151_));
 sg13g2_nand2_1 _3077_ (.Y(_0153_),
    .A(_0152_),
    .B(net110));
 sg13g2_nand3_1 _3078_ (.B(_2204_),
    .C(net74),
    .A(_2203_),
    .Y(_0154_));
 sg13g2_nand3_1 _3079_ (.B(_0154_),
    .C(net73),
    .A(_0153_),
    .Y(_0155_));
 sg13g2_buf_1 _3080_ (.A(_1780_),
    .X(_0156_));
 sg13g2_nand3_1 _3081_ (.B(_2208_),
    .C(_0156_),
    .A(_2206_),
    .Y(_0157_));
 sg13g2_nand3_1 _3082_ (.B(_0157_),
    .C(net77),
    .A(_0155_),
    .Y(_0158_));
 sg13g2_buf_1 _3083_ (.A(net112),
    .X(_0159_));
 sg13g2_nand3_1 _3084_ (.B(_0158_),
    .C(net67),
    .A(_2248_),
    .Y(_0160_));
 sg13g2_buf_1 _3085_ (.A(net109),
    .X(_0161_));
 sg13g2_nand3_1 _3086_ (.B(_0160_),
    .C(net66),
    .A(_2246_),
    .Y(_0162_));
 sg13g2_buf_1 _3087_ (.A(net149),
    .X(_0163_));
 sg13g2_nand3_1 _3088_ (.B(_0162_),
    .C(net107),
    .A(_2245_),
    .Y(_0164_));
 sg13g2_buf_1 _3089_ (.A(_1721_),
    .X(_0165_));
 sg13g2_buf_1 _3090_ (.A(_0165_),
    .X(_0166_));
 sg13g2_nand3_1 _3091_ (.B(_0164_),
    .C(net106),
    .A(_2244_),
    .Y(_0167_));
 sg13g2_buf_1 _3092_ (.A(_1655_),
    .X(_0168_));
 sg13g2_buf_1 _3093_ (.A(net146),
    .X(_0169_));
 sg13g2_nand3_1 _3094_ (.B(_0167_),
    .C(net105),
    .A(_2243_),
    .Y(_0170_));
 sg13g2_buf_1 _3095_ (.A(_0165_),
    .X(_0171_));
 sg13g2_nand3_1 _3096_ (.B(_2242_),
    .C(net104),
    .A(_2221_),
    .Y(_0172_));
 sg13g2_nand2_1 _3097_ (.Y(_0173_),
    .A(_2241_),
    .B(net108));
 sg13g2_buf_1 _3098_ (.A(net170),
    .X(_0174_));
 sg13g2_nand3_1 _3099_ (.B(net109),
    .C(_2238_),
    .A(_2230_),
    .Y(_0175_));
 sg13g2_nand3_1 _3100_ (.B(net112),
    .C(_2237_),
    .A(_2231_),
    .Y(_0176_));
 sg13g2_nand3_1 _3101_ (.B(net114),
    .C(_2236_),
    .A(_2232_),
    .Y(_0177_));
 sg13g2_nand3_1 _3102_ (.B(net115),
    .C(_2235_),
    .A(_2233_),
    .Y(_0178_));
 sg13g2_inv_1 _3103_ (.Y(_0179_),
    .A(_0038_));
 sg13g2_nand2_1 _3104_ (.Y(_0180_),
    .A(_2234_),
    .B(_0179_));
 sg13g2_nand2_1 _3105_ (.Y(_0181_),
    .A(_0180_),
    .B(net120));
 sg13g2_nand3_1 _3106_ (.B(net121),
    .C(_0181_),
    .A(_0178_),
    .Y(_0182_));
 sg13g2_nand3_1 _3107_ (.B(net83),
    .C(_0182_),
    .A(_0177_),
    .Y(_0183_));
 sg13g2_nand3_1 _3108_ (.B(net123),
    .C(_0183_),
    .A(_0176_),
    .Y(_0184_));
 sg13g2_nand3_1 _3109_ (.B(net124),
    .C(_0184_),
    .A(_0175_),
    .Y(_0185_));
 sg13g2_nand3_1 _3110_ (.B(net103),
    .C(_0185_),
    .A(_0173_),
    .Y(_0186_));
 sg13g2_buf_1 _3111_ (.A(net171),
    .X(_0187_));
 sg13g2_nand3_1 _3112_ (.B(_0186_),
    .C(net102),
    .A(_0172_),
    .Y(_0188_));
 sg13g2_inv_1 _3113_ (.Y(_0189_),
    .A(net189));
 sg13g2_inv_1 _3114_ (.Y(_0190_),
    .A(net2));
 sg13g2_nor2_1 _3115_ (.A(net1),
    .B(_0190_),
    .Y(_0191_));
 sg13g2_inv_1 _3116_ (.Y(_0192_),
    .A(_0191_));
 sg13g2_nor3_1 _3117_ (.A(_0189_),
    .B(_1659_),
    .C(_0192_),
    .Y(_0193_));
 sg13g2_buf_1 _3118_ (.A(_0193_),
    .X(_0194_));
 sg13g2_buf_1 _3119_ (.A(_0194_),
    .X(_0195_));
 sg13g2_nand3_1 _3120_ (.B(_0188_),
    .C(net50),
    .A(_0170_),
    .Y(_0196_));
 sg13g2_buf_1 _3121_ (.A(net162),
    .X(_0197_));
 sg13g2_nor2_1 _3122_ (.A(_1347_),
    .B(_0192_),
    .Y(_0198_));
 sg13g2_buf_1 _3123_ (.A(_0198_),
    .X(_0199_));
 sg13g2_buf_1 _3124_ (.A(_0199_),
    .X(_0200_));
 sg13g2_a22oi_1 _3125_ (.Y(_0201_),
    .B1(net101),
    .B2(net49),
    .A2(_1617_),
    .A1(net55));
 sg13g2_nand2_1 _3126_ (.Y(_0202_),
    .A(_0190_),
    .B(net1));
 sg13g2_buf_1 _3127_ (.A(_0202_),
    .X(_0203_));
 sg13g2_inv_2 _3128_ (.Y(_0204_),
    .A(net145));
 sg13g2_buf_1 _3129_ (.A(_0204_),
    .X(_0205_));
 sg13g2_nand3_1 _3130_ (.B(_1627_),
    .C(_1617_),
    .A(net64),
    .Y(_0206_));
 sg13g2_nand2_1 _3131_ (.Y(_0207_),
    .A(_0201_),
    .B(_0206_));
 sg13g2_buf_1 _3132_ (.A(_0204_),
    .X(_0208_));
 sg13g2_buf_1 _3133_ (.A(net189),
    .X(_0209_));
 sg13g2_nand2_1 _3134_ (.Y(_0210_),
    .A(net172),
    .B(_1617_));
 sg13g2_nor2_1 _3135_ (.A(_0210_),
    .B(net138),
    .Y(_0211_));
 sg13g2_a21oi_1 _3136_ (.A1(_0208_),
    .A2(_0210_),
    .Y(_0212_),
    .B1(_0211_));
 sg13g2_buf_1 _3137_ (.A(_1663_),
    .X(_0213_));
 sg13g2_nor2_1 _3138_ (.A(_1662_),
    .B(_0192_),
    .Y(_0214_));
 sg13g2_buf_2 _3139_ (.A(_0214_),
    .X(_0215_));
 sg13g2_buf_1 _3140_ (.A(_0215_),
    .X(_0216_));
 sg13g2_a22oi_1 _3141_ (.Y(_0217_),
    .B1(_1750_),
    .B2(net38),
    .A2(net178),
    .A1(net41));
 sg13g2_o21ai_1 _3142_ (.B1(_0217_),
    .Y(_0218_),
    .A1(_1627_),
    .A2(_0212_));
 sg13g2_nor3_1 _3143_ (.A(_0189_),
    .B(_1325_),
    .C(_0192_),
    .Y(_0219_));
 sg13g2_buf_1 _3144_ (.A(_0219_),
    .X(_0220_));
 sg13g2_buf_1 _3145_ (.A(net62),
    .X(_0221_));
 sg13g2_and3_1 _3146_ (.X(_0222_),
    .A(_0133_),
    .B(net48),
    .C(_0134_));
 sg13g2_nor3_1 _3147_ (.A(_0207_),
    .B(_0218_),
    .C(_0222_),
    .Y(_0223_));
 sg13g2_a21oi_1 _3148_ (.A1(_0196_),
    .A2(_0223_),
    .Y(_0224_),
    .B1(_1620_));
 sg13g2_nand3_1 _3149_ (.B(_0129_),
    .C(net130),
    .A(_0128_),
    .Y(_0225_));
 sg13g2_nand3_1 _3150_ (.B(_0127_),
    .C(net129),
    .A(_2249_),
    .Y(_0226_));
 sg13g2_nand3_1 _3151_ (.B(_0126_),
    .C(net128),
    .A(_2250_),
    .Y(_0227_));
 sg13g2_nand3_1 _3152_ (.B(_0125_),
    .C(net126),
    .A(_2251_),
    .Y(_0228_));
 sg13g2_nand3_1 _3153_ (.B(_0124_),
    .C(net125),
    .A(_2252_),
    .Y(_0229_));
 sg13g2_nand3_1 _3154_ (.B(_2256_),
    .C(net169),
    .A(_2253_),
    .Y(_0230_));
 sg13g2_nand3_1 _3155_ (.B(net179),
    .C(_2255_),
    .A(_2254_),
    .Y(_0231_));
 sg13g2_nand2b_1 _3156_ (.Y(_0232_),
    .B(_1838_),
    .A_N(_0023_));
 sg13g2_nand3_1 _3157_ (.B(_1845_),
    .C(_0232_),
    .A(_0231_),
    .Y(_0233_));
 sg13g2_nand3_1 _3158_ (.B(_0233_),
    .C(net164),
    .A(_0230_),
    .Y(_0234_));
 sg13g2_nand3_1 _3159_ (.B(_0234_),
    .C(net163),
    .A(_0229_),
    .Y(_0235_));
 sg13g2_nand3_1 _3160_ (.B(_0235_),
    .C(net158),
    .A(_0228_),
    .Y(_0236_));
 sg13g2_nand3_1 _3161_ (.B(_0236_),
    .C(net157),
    .A(_0227_),
    .Y(_0237_));
 sg13g2_nand3_1 _3162_ (.B(_0237_),
    .C(net151),
    .A(_0226_),
    .Y(_0238_));
 sg13g2_nand3_1 _3163_ (.B(_0238_),
    .C(net148),
    .A(_0225_),
    .Y(_0239_));
 sg13g2_nand3_1 _3164_ (.B(_0131_),
    .C(net131),
    .A(_0130_),
    .Y(_0240_));
 sg13g2_nand3_1 _3165_ (.B(_0240_),
    .C(net132),
    .A(_0239_),
    .Y(_0241_));
 sg13g2_nand3_1 _3166_ (.B(_0238_),
    .C(net131),
    .A(_0225_),
    .Y(_0242_));
 sg13g2_nand3_1 _3167_ (.B(_0237_),
    .C(net130),
    .A(_0226_),
    .Y(_0243_));
 sg13g2_nand3_1 _3168_ (.B(_0236_),
    .C(net129),
    .A(_0227_),
    .Y(_0244_));
 sg13g2_nand3_1 _3169_ (.B(_0235_),
    .C(net128),
    .A(_0228_),
    .Y(_0245_));
 sg13g2_nand3_1 _3170_ (.B(_0234_),
    .C(net126),
    .A(_0229_),
    .Y(_0246_));
 sg13g2_nand3_1 _3171_ (.B(_0233_),
    .C(net125),
    .A(_0230_),
    .Y(_0247_));
 sg13g2_nand3_1 _3172_ (.B(net169),
    .C(_0232_),
    .A(_0231_),
    .Y(_0248_));
 sg13g2_nand2_1 _3173_ (.Y(_0249_),
    .A(_0022_),
    .B(_1845_));
 sg13g2_nand3_1 _3174_ (.B(_1927_),
    .C(_0249_),
    .A(_0248_),
    .Y(_0250_));
 sg13g2_nand3_1 _3175_ (.B(_0250_),
    .C(net163),
    .A(_0247_),
    .Y(_0251_));
 sg13g2_nand3_1 _3176_ (.B(_0251_),
    .C(net158),
    .A(_0246_),
    .Y(_0252_));
 sg13g2_nand3_1 _3177_ (.B(_0252_),
    .C(net157),
    .A(_0245_),
    .Y(_0253_));
 sg13g2_nand3_1 _3178_ (.B(_0253_),
    .C(net151),
    .A(_0244_),
    .Y(_0254_));
 sg13g2_nand3_1 _3179_ (.B(_0254_),
    .C(net148),
    .A(_0243_),
    .Y(_0255_));
 sg13g2_buf_1 _3180_ (.A(net181),
    .X(_0256_));
 sg13g2_nand3_1 _3181_ (.B(_0255_),
    .C(net144),
    .A(_0242_),
    .Y(_0257_));
 sg13g2_buf_1 _3182_ (.A(_1693_),
    .X(_0258_));
 sg13g2_nand3_1 _3183_ (.B(_0257_),
    .C(net143),
    .A(_0241_),
    .Y(_0259_));
 sg13g2_nand3_1 _3184_ (.B(_0240_),
    .C(net144),
    .A(_0239_),
    .Y(_0260_));
 sg13g2_nand3_1 _3185_ (.B(_0134_),
    .C(_1700_),
    .A(_0133_),
    .Y(_0261_));
 sg13g2_nand3_1 _3186_ (.B(_0261_),
    .C(_1696_),
    .A(_0260_),
    .Y(_0262_));
 sg13g2_nand3_1 _3187_ (.B(_0262_),
    .C(net88),
    .A(_0259_),
    .Y(_0263_));
 sg13g2_nand3_1 _3188_ (.B(_0257_),
    .C(net87),
    .A(_0241_),
    .Y(_0264_));
 sg13g2_nand3_1 _3189_ (.B(_0255_),
    .C(net132),
    .A(_0242_),
    .Y(_0265_));
 sg13g2_nand3_1 _3190_ (.B(_0254_),
    .C(net131),
    .A(_0243_),
    .Y(_0266_));
 sg13g2_nand3_1 _3191_ (.B(_0253_),
    .C(net130),
    .A(_0244_),
    .Y(_0267_));
 sg13g2_nand3_1 _3192_ (.B(_0252_),
    .C(net129),
    .A(_0245_),
    .Y(_0268_));
 sg13g2_nand3_1 _3193_ (.B(_0251_),
    .C(net128),
    .A(_0246_),
    .Y(_0269_));
 sg13g2_nand3_1 _3194_ (.B(_0250_),
    .C(net126),
    .A(_0247_),
    .Y(_0270_));
 sg13g2_nand3_1 _3195_ (.B(net125),
    .C(_0249_),
    .A(_0248_),
    .Y(_0271_));
 sg13g2_nand2b_1 _3196_ (.Y(_0272_),
    .B(_1927_),
    .A_N(_0021_));
 sg13g2_nand3_1 _3197_ (.B(net163),
    .C(_0272_),
    .A(_0271_),
    .Y(_0273_));
 sg13g2_nand3_1 _3198_ (.B(_0273_),
    .C(_2006_),
    .A(_0270_),
    .Y(_0274_));
 sg13g2_nand3_1 _3199_ (.B(_0274_),
    .C(net157),
    .A(_0269_),
    .Y(_0275_));
 sg13g2_nand3_1 _3200_ (.B(_0275_),
    .C(net151),
    .A(_0268_),
    .Y(_0276_));
 sg13g2_nand3_1 _3201_ (.B(_0276_),
    .C(net148),
    .A(_0267_),
    .Y(_0277_));
 sg13g2_nand3_1 _3202_ (.B(_0277_),
    .C(net144),
    .A(_0266_),
    .Y(_0278_));
 sg13g2_nand3_1 _3203_ (.B(_0278_),
    .C(net143),
    .A(_0265_),
    .Y(_0279_));
 sg13g2_buf_1 _3204_ (.A(net165),
    .X(_0280_));
 sg13g2_nand3_1 _3205_ (.B(_0279_),
    .C(net100),
    .A(_0264_),
    .Y(_0281_));
 sg13g2_nand3_1 _3206_ (.B(_0281_),
    .C(net101),
    .A(_0263_),
    .Y(_0282_));
 sg13g2_nand3_1 _3207_ (.B(_0262_),
    .C(net100),
    .A(_0259_),
    .Y(_0283_));
 sg13g2_nand3_1 _3208_ (.B(_0261_),
    .C(net143),
    .A(_0260_),
    .Y(_0284_));
 sg13g2_nand3_1 _3209_ (.B(_0136_),
    .C(_1696_),
    .A(_0135_),
    .Y(_0285_));
 sg13g2_nand3_1 _3210_ (.B(_0285_),
    .C(_1691_),
    .A(_0284_),
    .Y(_0286_));
 sg13g2_nand3_1 _3211_ (.B(_0286_),
    .C(_1686_),
    .A(_0283_),
    .Y(_0287_));
 sg13g2_nand3_1 _3212_ (.B(_0287_),
    .C(net90),
    .A(_0282_),
    .Y(_0288_));
 sg13g2_nand3_1 _3213_ (.B(_0281_),
    .C(net89),
    .A(_0263_),
    .Y(_0289_));
 sg13g2_nand3_1 _3214_ (.B(_0279_),
    .C(net88),
    .A(_0264_),
    .Y(_0290_));
 sg13g2_nand3_1 _3215_ (.B(_0278_),
    .C(net87),
    .A(_0265_),
    .Y(_0291_));
 sg13g2_nand3_1 _3216_ (.B(_0277_),
    .C(net132),
    .A(_0266_),
    .Y(_0292_));
 sg13g2_nand3_1 _3217_ (.B(_0276_),
    .C(net131),
    .A(_0267_),
    .Y(_0293_));
 sg13g2_nand3_1 _3218_ (.B(_0275_),
    .C(net130),
    .A(_0268_),
    .Y(_0294_));
 sg13g2_nand3_1 _3219_ (.B(_0274_),
    .C(net129),
    .A(_0269_),
    .Y(_0295_));
 sg13g2_nand3_1 _3220_ (.B(_0273_),
    .C(net128),
    .A(_0270_),
    .Y(_0296_));
 sg13g2_nand3_1 _3221_ (.B(_1727_),
    .C(_0272_),
    .A(_0271_),
    .Y(_0297_));
 sg13g2_nand2_1 _3222_ (.Y(_0298_),
    .A(_0020_),
    .B(net163));
 sg13g2_nand3_1 _3223_ (.B(_2006_),
    .C(_0298_),
    .A(_0297_),
    .Y(_0299_));
 sg13g2_nand3_1 _3224_ (.B(_0299_),
    .C(net157),
    .A(_0296_),
    .Y(_0300_));
 sg13g2_nand3_1 _3225_ (.B(_0300_),
    .C(net151),
    .A(_0295_),
    .Y(_0301_));
 sg13g2_nand3_1 _3226_ (.B(_0301_),
    .C(net148),
    .A(_0294_),
    .Y(_0302_));
 sg13g2_nand3_1 _3227_ (.B(_0302_),
    .C(net144),
    .A(_0293_),
    .Y(_0303_));
 sg13g2_nand3_1 _3228_ (.B(_0303_),
    .C(net143),
    .A(_0292_),
    .Y(_0304_));
 sg13g2_nand3_1 _3229_ (.B(_0304_),
    .C(net100),
    .A(_0291_),
    .Y(_0305_));
 sg13g2_nand3_1 _3230_ (.B(_0305_),
    .C(net101),
    .A(_0290_),
    .Y(_0306_));
 sg13g2_buf_1 _3231_ (.A(net159),
    .X(_0307_));
 sg13g2_nand3_1 _3232_ (.B(_0306_),
    .C(net99),
    .A(_0289_),
    .Y(_0308_));
 sg13g2_buf_1 _3233_ (.A(net160),
    .X(_0309_));
 sg13g2_nand3_1 _3234_ (.B(_0308_),
    .C(_0309_),
    .A(_0288_),
    .Y(_0310_));
 sg13g2_nand3_1 _3235_ (.B(_0287_),
    .C(net99),
    .A(_0282_),
    .Y(_0311_));
 sg13g2_nand3_1 _3236_ (.B(_0286_),
    .C(net101),
    .A(_0283_),
    .Y(_0312_));
 sg13g2_nand3_1 _3237_ (.B(_0285_),
    .C(net100),
    .A(_0284_),
    .Y(_0313_));
 sg13g2_nand3_1 _3238_ (.B(_0138_),
    .C(net88),
    .A(_0137_),
    .Y(_0314_));
 sg13g2_nand3_1 _3239_ (.B(_0314_),
    .C(net89),
    .A(_0313_),
    .Y(_0315_));
 sg13g2_nand3_1 _3240_ (.B(_0315_),
    .C(net90),
    .A(_0312_),
    .Y(_0316_));
 sg13g2_nand3_1 _3241_ (.B(_0316_),
    .C(net54),
    .A(_0311_),
    .Y(_0317_));
 sg13g2_nand3_1 _3242_ (.B(_0317_),
    .C(net51),
    .A(_0310_),
    .Y(_0318_));
 sg13g2_nand3_1 _3243_ (.B(_0308_),
    .C(net54),
    .A(_0288_),
    .Y(_0319_));
 sg13g2_nand3_1 _3244_ (.B(_0306_),
    .C(_1681_),
    .A(_0289_),
    .Y(_0320_));
 sg13g2_nand3_1 _3245_ (.B(_0305_),
    .C(net89),
    .A(_0290_),
    .Y(_0321_));
 sg13g2_nand3_1 _3246_ (.B(_0304_),
    .C(net88),
    .A(_0291_),
    .Y(_0322_));
 sg13g2_nand3_1 _3247_ (.B(_0303_),
    .C(net87),
    .A(_0292_),
    .Y(_0323_));
 sg13g2_nand3_1 _3248_ (.B(_0302_),
    .C(net132),
    .A(_0293_),
    .Y(_0324_));
 sg13g2_nand3_1 _3249_ (.B(_0301_),
    .C(net131),
    .A(_0294_),
    .Y(_0325_));
 sg13g2_nand3_1 _3250_ (.B(_0300_),
    .C(net130),
    .A(_0295_),
    .Y(_0326_));
 sg13g2_nand3_1 _3251_ (.B(_0299_),
    .C(net129),
    .A(_0296_),
    .Y(_0327_));
 sg13g2_nand3_1 _3252_ (.B(_1718_),
    .C(_0298_),
    .A(_0297_),
    .Y(_0328_));
 sg13g2_nand2b_1 _3253_ (.Y(_0329_),
    .B(_1717_),
    .A_N(_0019_));
 sg13g2_nand3_1 _3254_ (.B(net157),
    .C(_0329_),
    .A(_0328_),
    .Y(_0330_));
 sg13g2_nand3_1 _3255_ (.B(_0330_),
    .C(_2179_),
    .A(_0327_),
    .Y(_0331_));
 sg13g2_nand3_1 _3256_ (.B(_0331_),
    .C(net148),
    .A(_0326_),
    .Y(_0332_));
 sg13g2_nand3_1 _3257_ (.B(_0332_),
    .C(net144),
    .A(_0325_),
    .Y(_0333_));
 sg13g2_nand3_1 _3258_ (.B(_0333_),
    .C(net143),
    .A(_0324_),
    .Y(_0334_));
 sg13g2_nand3_1 _3259_ (.B(_0334_),
    .C(net100),
    .A(_0323_),
    .Y(_0335_));
 sg13g2_nand3_1 _3260_ (.B(_0335_),
    .C(net101),
    .A(_0322_),
    .Y(_0336_));
 sg13g2_nand3_1 _3261_ (.B(_0336_),
    .C(net99),
    .A(_0321_),
    .Y(_0337_));
 sg13g2_nand3_1 _3262_ (.B(_0337_),
    .C(net98),
    .A(_0320_),
    .Y(_0338_));
 sg13g2_buf_1 _3263_ (.A(net116),
    .X(_0339_));
 sg13g2_nand3_1 _3264_ (.B(_0338_),
    .C(net61),
    .A(_0319_),
    .Y(_0340_));
 sg13g2_nand3_1 _3265_ (.B(_0340_),
    .C(net75),
    .A(_0318_),
    .Y(_0341_));
 sg13g2_nand3_1 _3266_ (.B(_0317_),
    .C(net61),
    .A(_0310_),
    .Y(_0342_));
 sg13g2_nand3_1 _3267_ (.B(_0316_),
    .C(net98),
    .A(_0311_),
    .Y(_0343_));
 sg13g2_nand3_1 _3268_ (.B(_0315_),
    .C(net99),
    .A(_0312_),
    .Y(_0344_));
 sg13g2_nand3_1 _3269_ (.B(_0314_),
    .C(net101),
    .A(_0313_),
    .Y(_0345_));
 sg13g2_nand3_1 _3270_ (.B(_0140_),
    .C(net89),
    .A(_0139_),
    .Y(_0346_));
 sg13g2_nand3_1 _3271_ (.B(_0346_),
    .C(net90),
    .A(_0345_),
    .Y(_0347_));
 sg13g2_nand3_1 _3272_ (.B(_0347_),
    .C(net54),
    .A(_0344_),
    .Y(_0348_));
 sg13g2_nand3_1 _3273_ (.B(_0348_),
    .C(_1798_),
    .A(_0343_),
    .Y(_0349_));
 sg13g2_nand3_1 _3274_ (.B(_0349_),
    .C(net52),
    .A(_0342_),
    .Y(_0350_));
 sg13g2_nand3_1 _3275_ (.B(_0350_),
    .C(net80),
    .A(_0341_),
    .Y(_0351_));
 sg13g2_nand3_1 _3276_ (.B(_0340_),
    .C(net52),
    .A(_0318_),
    .Y(_0352_));
 sg13g2_nand3_1 _3277_ (.B(_0338_),
    .C(net51),
    .A(_0319_),
    .Y(_0353_));
 sg13g2_nand3_1 _3278_ (.B(_0337_),
    .C(net54),
    .A(_0320_),
    .Y(_0354_));
 sg13g2_nand3_1 _3279_ (.B(_0336_),
    .C(_1681_),
    .A(_0321_),
    .Y(_0355_));
 sg13g2_nand3_1 _3280_ (.B(_0335_),
    .C(net89),
    .A(_0322_),
    .Y(_0356_));
 sg13g2_nand3_1 _3281_ (.B(_0334_),
    .C(net88),
    .A(_0323_),
    .Y(_0357_));
 sg13g2_nand3_1 _3282_ (.B(_0333_),
    .C(net87),
    .A(_0324_),
    .Y(_0358_));
 sg13g2_nand3_1 _3283_ (.B(_0332_),
    .C(net132),
    .A(_0325_),
    .Y(_0359_));
 sg13g2_nand3_1 _3284_ (.B(_0331_),
    .C(net131),
    .A(_0326_),
    .Y(_0360_));
 sg13g2_nand3_1 _3285_ (.B(_0330_),
    .C(net130),
    .A(_0327_),
    .Y(_0361_));
 sg13g2_nand3_1 _3286_ (.B(_1714_),
    .C(_0329_),
    .A(_0328_),
    .Y(_0362_));
 sg13g2_nand2_1 _3287_ (.Y(_0363_),
    .A(_0018_),
    .B(_1713_));
 sg13g2_nand3_1 _3288_ (.B(net151),
    .C(_0363_),
    .A(_0362_),
    .Y(_0364_));
 sg13g2_nand3_1 _3289_ (.B(_0364_),
    .C(net148),
    .A(_0361_),
    .Y(_0365_));
 sg13g2_nand3_1 _3290_ (.B(_0365_),
    .C(net144),
    .A(_0360_),
    .Y(_0366_));
 sg13g2_nand3_1 _3291_ (.B(_0366_),
    .C(net143),
    .A(_0359_),
    .Y(_0367_));
 sg13g2_nand3_1 _3292_ (.B(_0367_),
    .C(net100),
    .A(_0358_),
    .Y(_0368_));
 sg13g2_nand3_1 _3293_ (.B(_0368_),
    .C(net101),
    .A(_0357_),
    .Y(_0369_));
 sg13g2_nand3_1 _3294_ (.B(_0369_),
    .C(net99),
    .A(_0356_),
    .Y(_0370_));
 sg13g2_nand3_1 _3295_ (.B(_0370_),
    .C(net98),
    .A(_0355_),
    .Y(_0371_));
 sg13g2_nand3_1 _3296_ (.B(_0371_),
    .C(net61),
    .A(_0354_),
    .Y(_0372_));
 sg13g2_nand3_1 _3297_ (.B(_0372_),
    .C(net75),
    .A(_0353_),
    .Y(_0373_));
 sg13g2_nand3_1 _3298_ (.B(_0373_),
    .C(net110),
    .A(_0352_),
    .Y(_0374_));
 sg13g2_buf_1 _3299_ (.A(net115),
    .X(_0375_));
 sg13g2_nand3_1 _3300_ (.B(_0374_),
    .C(net60),
    .A(_0351_),
    .Y(_0376_));
 sg13g2_nand3_1 _3301_ (.B(_0350_),
    .C(net110),
    .A(_0341_),
    .Y(_0377_));
 sg13g2_nand3_1 _3302_ (.B(_0349_),
    .C(net75),
    .A(_0342_),
    .Y(_0378_));
 sg13g2_nand3_1 _3303_ (.B(_0348_),
    .C(net61),
    .A(_0343_),
    .Y(_0379_));
 sg13g2_nand3_1 _3304_ (.B(_0347_),
    .C(net98),
    .A(_0344_),
    .Y(_0380_));
 sg13g2_nand3_1 _3305_ (.B(_0346_),
    .C(net99),
    .A(_0345_),
    .Y(_0381_));
 sg13g2_nand3_1 _3306_ (.B(_0142_),
    .C(net90),
    .A(_0141_),
    .Y(_0382_));
 sg13g2_nand3_1 _3307_ (.B(_0382_),
    .C(net54),
    .A(_0381_),
    .Y(_0383_));
 sg13g2_nand3_1 _3308_ (.B(_0383_),
    .C(net51),
    .A(_0380_),
    .Y(_0384_));
 sg13g2_nand3_1 _3309_ (.B(_0384_),
    .C(net52),
    .A(_0379_),
    .Y(_0385_));
 sg13g2_nand3_1 _3310_ (.B(_0385_),
    .C(net80),
    .A(_0378_),
    .Y(_0386_));
 sg13g2_nand3_1 _3311_ (.B(_0386_),
    .C(net81),
    .A(_0377_),
    .Y(_0387_));
 sg13g2_nand3_1 _3312_ (.B(_0387_),
    .C(net82),
    .A(_0376_),
    .Y(_0388_));
 sg13g2_nand3_1 _3313_ (.B(_0374_),
    .C(net81),
    .A(_0351_),
    .Y(_0389_));
 sg13g2_nand3_1 _3314_ (.B(_0373_),
    .C(net80),
    .A(_0352_),
    .Y(_0390_));
 sg13g2_nand3_1 _3315_ (.B(_0372_),
    .C(_1792_),
    .A(_0353_),
    .Y(_0391_));
 sg13g2_nand3_1 _3316_ (.B(_0371_),
    .C(net51),
    .A(_0354_),
    .Y(_0392_));
 sg13g2_nand3_1 _3317_ (.B(_0370_),
    .C(net54),
    .A(_0355_),
    .Y(_0393_));
 sg13g2_nand3_1 _3318_ (.B(_0369_),
    .C(net90),
    .A(_0356_),
    .Y(_0394_));
 sg13g2_nand3_1 _3319_ (.B(_0368_),
    .C(net89),
    .A(_0357_),
    .Y(_0395_));
 sg13g2_nand3_1 _3320_ (.B(_0367_),
    .C(net88),
    .A(_0358_),
    .Y(_0396_));
 sg13g2_nand3_1 _3321_ (.B(_0366_),
    .C(net87),
    .A(_0359_),
    .Y(_0397_));
 sg13g2_nand3_1 _3322_ (.B(_0365_),
    .C(net132),
    .A(_0360_),
    .Y(_0398_));
 sg13g2_nand3_1 _3323_ (.B(_0364_),
    .C(net131),
    .A(_0361_),
    .Y(_0399_));
 sg13g2_nand3_1 _3324_ (.B(_1710_),
    .C(_0363_),
    .A(_0362_),
    .Y(_0400_));
 sg13g2_nand2b_1 _3325_ (.Y(_0401_),
    .B(_1709_),
    .A_N(_0017_));
 sg13g2_nand3_1 _3326_ (.B(_0132_),
    .C(_0401_),
    .A(_0400_),
    .Y(_0402_));
 sg13g2_nand3_1 _3327_ (.B(_0402_),
    .C(_0256_),
    .A(_0399_),
    .Y(_0403_));
 sg13g2_nand3_1 _3328_ (.B(_0403_),
    .C(_0258_),
    .A(_0398_),
    .Y(_0404_));
 sg13g2_nand3_1 _3329_ (.B(_0404_),
    .C(_0280_),
    .A(_0397_),
    .Y(_0405_));
 sg13g2_nand3_1 _3330_ (.B(_0405_),
    .C(_0197_),
    .A(_0396_),
    .Y(_0406_));
 sg13g2_nand3_1 _3331_ (.B(_0406_),
    .C(net99),
    .A(_0395_),
    .Y(_0407_));
 sg13g2_nand3_1 _3332_ (.B(_0407_),
    .C(net98),
    .A(_0394_),
    .Y(_0408_));
 sg13g2_nand3_1 _3333_ (.B(_0408_),
    .C(net61),
    .A(_0393_),
    .Y(_0409_));
 sg13g2_nand3_1 _3334_ (.B(_0409_),
    .C(net111),
    .A(_0392_),
    .Y(_0410_));
 sg13g2_nand3_1 _3335_ (.B(_0410_),
    .C(_2205_),
    .A(_0391_),
    .Y(_0411_));
 sg13g2_nand3_1 _3336_ (.B(_0411_),
    .C(net60),
    .A(_0390_),
    .Y(_0412_));
 sg13g2_nand3_1 _3337_ (.B(_0412_),
    .C(net72),
    .A(_0389_),
    .Y(_0413_));
 sg13g2_nand3_1 _3338_ (.B(_0413_),
    .C(net76),
    .A(_0388_),
    .Y(_0414_));
 sg13g2_nand3_1 _3339_ (.B(_0387_),
    .C(net72),
    .A(_0376_),
    .Y(_0415_));
 sg13g2_nand3_1 _3340_ (.B(_0386_),
    .C(net60),
    .A(_0377_),
    .Y(_0416_));
 sg13g2_nand3_1 _3341_ (.B(_0385_),
    .C(net110),
    .A(_0378_),
    .Y(_0417_));
 sg13g2_nand3_1 _3342_ (.B(_0384_),
    .C(net75),
    .A(_0379_),
    .Y(_0418_));
 sg13g2_nand3_1 _3343_ (.B(_0383_),
    .C(net61),
    .A(_0380_),
    .Y(_0419_));
 sg13g2_nand3_1 _3344_ (.B(_0382_),
    .C(net98),
    .A(_0381_),
    .Y(_0420_));
 sg13g2_nand3_1 _3345_ (.B(_0144_),
    .C(_1673_),
    .A(_0143_),
    .Y(_0421_));
 sg13g2_nand3_1 _3346_ (.B(_0421_),
    .C(_1798_),
    .A(_0420_),
    .Y(_0422_));
 sg13g2_nand3_1 _3347_ (.B(_0422_),
    .C(net52),
    .A(_0419_),
    .Y(_0423_));
 sg13g2_nand3_1 _3348_ (.B(_0423_),
    .C(net80),
    .A(_0418_),
    .Y(_0424_));
 sg13g2_nand3_1 _3349_ (.B(_0424_),
    .C(net81),
    .A(_0417_),
    .Y(_0425_));
 sg13g2_nand3_1 _3350_ (.B(_0425_),
    .C(net82),
    .A(_0416_),
    .Y(_0426_));
 sg13g2_nand3_1 _3351_ (.B(_0426_),
    .C(_1771_),
    .A(_0415_),
    .Y(_0427_));
 sg13g2_nand3_1 _3352_ (.B(_0427_),
    .C(net84),
    .A(_0414_),
    .Y(_0428_));
 sg13g2_nand3_1 _3353_ (.B(_0413_),
    .C(net53),
    .A(_0388_),
    .Y(_0429_));
 sg13g2_nand3_1 _3354_ (.B(_0412_),
    .C(net82),
    .A(_0389_),
    .Y(_0430_));
 sg13g2_nand3_1 _3355_ (.B(_0411_),
    .C(net81),
    .A(_0390_),
    .Y(_0431_));
 sg13g2_nand3_1 _3356_ (.B(_0410_),
    .C(net80),
    .A(_0391_),
    .Y(_0432_));
 sg13g2_nand3_1 _3357_ (.B(_0409_),
    .C(net52),
    .A(_0392_),
    .Y(_0433_));
 sg13g2_nand3_1 _3358_ (.B(_0408_),
    .C(net51),
    .A(_0393_),
    .Y(_0434_));
 sg13g2_nand3_1 _3359_ (.B(_0407_),
    .C(_1673_),
    .A(_0394_),
    .Y(_0435_));
 sg13g2_nand3_1 _3360_ (.B(_0406_),
    .C(net90),
    .A(_0395_),
    .Y(_0436_));
 sg13g2_nand3_1 _3361_ (.B(_0405_),
    .C(net89),
    .A(_0396_),
    .Y(_0437_));
 sg13g2_nand3_1 _3362_ (.B(_0404_),
    .C(net88),
    .A(_0397_),
    .Y(_0438_));
 sg13g2_nand3_1 _3363_ (.B(_0403_),
    .C(net87),
    .A(_0398_),
    .Y(_0439_));
 sg13g2_nand3_1 _3364_ (.B(_0402_),
    .C(_1700_),
    .A(_0399_),
    .Y(_0440_));
 sg13g2_nand3_1 _3365_ (.B(_1703_),
    .C(_0401_),
    .A(_0400_),
    .Y(_0441_));
 sg13g2_nand2_1 _3366_ (.Y(_0442_),
    .A(_0016_),
    .B(net180));
 sg13g2_nand3_1 _3367_ (.B(_0256_),
    .C(_0442_),
    .A(_0441_),
    .Y(_0443_));
 sg13g2_nand3_1 _3368_ (.B(_0443_),
    .C(_0258_),
    .A(_0440_),
    .Y(_0444_));
 sg13g2_nand3_1 _3369_ (.B(_0444_),
    .C(_0280_),
    .A(_0439_),
    .Y(_0445_));
 sg13g2_nand3_1 _3370_ (.B(_0445_),
    .C(net162),
    .A(_0438_),
    .Y(_0446_));
 sg13g2_nand3_1 _3371_ (.B(_0446_),
    .C(net159),
    .A(_0437_),
    .Y(_0447_));
 sg13g2_nand3_1 _3372_ (.B(_0447_),
    .C(net160),
    .A(_0436_),
    .Y(_0448_));
 sg13g2_nand3_1 _3373_ (.B(_0448_),
    .C(net116),
    .A(_0435_),
    .Y(_0449_));
 sg13g2_nand3_1 _3374_ (.B(_0449_),
    .C(net111),
    .A(_0434_),
    .Y(_0450_));
 sg13g2_nand3_1 _3375_ (.B(_0450_),
    .C(net113),
    .A(_0433_),
    .Y(_0451_));
 sg13g2_nand3_1 _3376_ (.B(_0451_),
    .C(net73),
    .A(_0432_),
    .Y(_0452_));
 sg13g2_nand3_1 _3377_ (.B(_0452_),
    .C(net72),
    .A(_0431_),
    .Y(_0453_));
 sg13g2_nand3_1 _3378_ (.B(_0453_),
    .C(net76),
    .A(_0430_),
    .Y(_0454_));
 sg13g2_nand3_1 _3379_ (.B(_0454_),
    .C(net71),
    .A(_0429_),
    .Y(_0455_));
 sg13g2_nand3_1 _3380_ (.B(_0455_),
    .C(net70),
    .A(_0428_),
    .Y(_0456_));
 sg13g2_nand3_1 _3381_ (.B(_0427_),
    .C(net71),
    .A(_0414_),
    .Y(_0457_));
 sg13g2_nand3_1 _3382_ (.B(_0426_),
    .C(net76),
    .A(_0415_),
    .Y(_0458_));
 sg13g2_nand3_1 _3383_ (.B(_0425_),
    .C(net72),
    .A(_0416_),
    .Y(_0459_));
 sg13g2_nand3_1 _3384_ (.B(_0424_),
    .C(net60),
    .A(_0417_),
    .Y(_0460_));
 sg13g2_nand3_1 _3385_ (.B(_0423_),
    .C(net110),
    .A(_0418_),
    .Y(_0461_));
 sg13g2_nand3_1 _3386_ (.B(_0422_),
    .C(net75),
    .A(_0419_),
    .Y(_0462_));
 sg13g2_nand3_1 _3387_ (.B(_0421_),
    .C(net61),
    .A(_0420_),
    .Y(_0463_));
 sg13g2_nand3_1 _3388_ (.B(_0146_),
    .C(net78),
    .A(_0145_),
    .Y(_0464_));
 sg13g2_nand3_1 _3389_ (.B(_0464_),
    .C(net52),
    .A(_0463_),
    .Y(_0465_));
 sg13g2_nand3_1 _3390_ (.B(_0465_),
    .C(net74),
    .A(_0462_),
    .Y(_0466_));
 sg13g2_nand3_1 _3391_ (.B(_0466_),
    .C(_1781_),
    .A(_0461_),
    .Y(_0467_));
 sg13g2_nand3_1 _3392_ (.B(_0467_),
    .C(_2247_),
    .A(_0460_),
    .Y(_0468_));
 sg13g2_nand3_1 _3393_ (.B(_0468_),
    .C(_1771_),
    .A(_0459_),
    .Y(_0469_));
 sg13g2_nand3_1 _3394_ (.B(_0469_),
    .C(net84),
    .A(_0458_),
    .Y(_0470_));
 sg13g2_nand3_1 _3395_ (.B(_0470_),
    .C(net85),
    .A(_0457_),
    .Y(_0471_));
 sg13g2_nand3_1 _3396_ (.B(_0471_),
    .C(net104),
    .A(_0456_),
    .Y(_0472_));
 sg13g2_nand3_1 _3397_ (.B(_0470_),
    .C(net70),
    .A(_0457_),
    .Y(_0473_));
 sg13g2_nand3_1 _3398_ (.B(_0469_),
    .C(net71),
    .A(_0458_),
    .Y(_0474_));
 sg13g2_nand3_1 _3399_ (.B(_0468_),
    .C(net67),
    .A(_0459_),
    .Y(_0475_));
 sg13g2_nand3_1 _3400_ (.B(_0467_),
    .C(_2211_),
    .A(_0460_),
    .Y(_0476_));
 sg13g2_nand3_1 _3401_ (.B(_0466_),
    .C(_2209_),
    .A(_0461_),
    .Y(_0477_));
 sg13g2_nand3_1 _3402_ (.B(_0465_),
    .C(net110),
    .A(_0462_),
    .Y(_0478_));
 sg13g2_nand3_1 _3403_ (.B(_0464_),
    .C(net111),
    .A(_0463_),
    .Y(_0479_));
 sg13g2_nand3_1 _3404_ (.B(_0148_),
    .C(net79),
    .A(_0147_),
    .Y(_0480_));
 sg13g2_nand3_1 _3405_ (.B(_0480_),
    .C(net74),
    .A(_0479_),
    .Y(_0481_));
 sg13g2_nand3_1 _3406_ (.B(_0481_),
    .C(_0156_),
    .A(_0478_),
    .Y(_0482_));
 sg13g2_nand3_1 _3407_ (.B(_0482_),
    .C(net69),
    .A(_0477_),
    .Y(_0483_));
 sg13g2_buf_1 _3408_ (.A(net83),
    .X(_0484_));
 sg13g2_nand3_1 _3409_ (.B(_0483_),
    .C(net47),
    .A(_0476_),
    .Y(_0485_));
 sg13g2_buf_1 _3410_ (.A(_1764_),
    .X(_0486_));
 sg13g2_nand3_1 _3411_ (.B(_0485_),
    .C(_0486_),
    .A(_0475_),
    .Y(_0487_));
 sg13g2_buf_1 _3412_ (.A(_1755_),
    .X(_0488_));
 sg13g2_buf_1 _3413_ (.A(_0488_),
    .X(_0489_));
 sg13g2_nand3_1 _3414_ (.B(_0487_),
    .C(net58),
    .A(_0474_),
    .Y(_0490_));
 sg13g2_buf_1 _3415_ (.A(net127),
    .X(_0491_));
 sg13g2_nand3_1 _3416_ (.B(_0490_),
    .C(net57),
    .A(_0473_),
    .Y(_0492_));
 sg13g2_buf_1 _3417_ (.A(_0168_),
    .X(_0493_));
 sg13g2_nand3_1 _3418_ (.B(_0492_),
    .C(net96),
    .A(_0472_),
    .Y(_0494_));
 sg13g2_nand3_1 _3419_ (.B(_0487_),
    .C(net70),
    .A(_0474_),
    .Y(_0495_));
 sg13g2_nand3_1 _3420_ (.B(_0483_),
    .C(net76),
    .A(_0476_),
    .Y(_0496_));
 sg13g2_nand3_1 _3421_ (.B(_0481_),
    .C(net60),
    .A(_0478_),
    .Y(_0497_));
 sg13g2_nand2_1 _3422_ (.Y(_0498_),
    .A(_0152_),
    .B(net80));
 sg13g2_nand3_1 _3423_ (.B(_0480_),
    .C(net110),
    .A(_0479_),
    .Y(_0499_));
 sg13g2_nand3_1 _3424_ (.B(_0499_),
    .C(net81),
    .A(_0498_),
    .Y(_0500_));
 sg13g2_nand3_1 _3425_ (.B(_0500_),
    .C(net82),
    .A(_0497_),
    .Y(_0501_));
 sg13g2_nand3_1 _3426_ (.B(_0482_),
    .C(net72),
    .A(_0477_),
    .Y(_0502_));
 sg13g2_nand3_1 _3427_ (.B(_0502_),
    .C(net53),
    .A(_0501_),
    .Y(_0503_));
 sg13g2_nand3_1 _3428_ (.B(_0503_),
    .C(net84),
    .A(_0496_),
    .Y(_0504_));
 sg13g2_nand3_1 _3429_ (.B(_0485_),
    .C(_2216_),
    .A(_0475_),
    .Y(_0505_));
 sg13g2_nand3_1 _3430_ (.B(_0505_),
    .C(net85),
    .A(_0504_),
    .Y(_0506_));
 sg13g2_nand3_1 _3431_ (.B(_0506_),
    .C(net86),
    .A(_0495_),
    .Y(_0507_));
 sg13g2_nand3_1 _3432_ (.B(_0490_),
    .C(net106),
    .A(_0473_),
    .Y(_0508_));
 sg13g2_buf_1 _3433_ (.A(net171),
    .X(_0509_));
 sg13g2_nand3_1 _3434_ (.B(_0508_),
    .C(net95),
    .A(_0507_),
    .Y(_0510_));
 sg13g2_buf_1 _3435_ (.A(_0194_),
    .X(_0511_));
 sg13g2_nand3_1 _3436_ (.B(_0510_),
    .C(net46),
    .A(_0494_),
    .Y(_0512_));
 sg13g2_nand3_1 _3437_ (.B(_0442_),
    .C(_0221_),
    .A(_0441_),
    .Y(_0513_));
 sg13g2_buf_1 _3438_ (.A(_0215_),
    .X(_0514_));
 sg13g2_a22oi_1 _3439_ (.Y(_0515_),
    .B1(net178),
    .B2(net37),
    .A2(_2202_),
    .A1(_0200_));
 sg13g2_buf_1 _3440_ (.A(_0189_),
    .X(_0516_));
 sg13g2_nor3_1 _3441_ (.A(_0516_),
    .B(_1598_),
    .C(_1589_),
    .Y(_0517_));
 sg13g2_a22oi_1 _3442_ (.Y(_0518_),
    .B1(_1588_),
    .B2(net55),
    .A2(net188),
    .A1(_0517_));
 sg13g2_inv_1 _3443_ (.Y(_0519_),
    .A(_0517_));
 sg13g2_buf_1 _3444_ (.A(net145),
    .X(_0520_));
 sg13g2_a21oi_1 _3445_ (.A1(_1598_),
    .A2(_1589_),
    .Y(_0521_),
    .B1(net94));
 sg13g2_a22oi_1 _3446_ (.Y(_0522_),
    .B1(_0519_),
    .B2(_0521_),
    .A2(net148),
    .A1(net42));
 sg13g2_and4_1 _3447_ (.A(_0513_),
    .B(_0515_),
    .C(_0518_),
    .D(_0522_),
    .X(_0523_));
 sg13g2_a21oi_1 _3448_ (.A1(_0512_),
    .A2(_0523_),
    .Y(_0524_),
    .B1(_1591_));
 sg13g2_nor2_1 _3449_ (.A(_0224_),
    .B(_0524_),
    .Y(_0525_));
 sg13g2_nand3_1 _3450_ (.B(_1699_),
    .C(_0442_),
    .A(_0441_),
    .Y(_0526_));
 sg13g2_nand2b_1 _3451_ (.Y(_0527_),
    .B(net181),
    .A_N(_0015_));
 sg13g2_nand3_1 _3452_ (.B(net133),
    .C(_0527_),
    .A(_0526_),
    .Y(_0528_));
 sg13g2_nand2_1 _3453_ (.Y(_0529_),
    .A(_0014_),
    .B(\ayayayayayaya.b[14] ));
 sg13g2_nand2_1 _3454_ (.Y(_0530_),
    .A(_0528_),
    .B(_0529_));
 sg13g2_nand2_1 _3455_ (.Y(_0531_),
    .A(_0530_),
    .B(net134));
 sg13g2_nand2_1 _3456_ (.Y(_0532_),
    .A(_0013_),
    .B(_1688_));
 sg13g2_nand2_1 _3457_ (.Y(_0533_),
    .A(_0531_),
    .B(_0532_));
 sg13g2_nand2_1 _3458_ (.Y(_0534_),
    .A(_0533_),
    .B(net135));
 sg13g2_nand2_1 _3459_ (.Y(_0535_),
    .A(_0012_),
    .B(net183));
 sg13g2_nand2_1 _3460_ (.Y(_0536_),
    .A(_0534_),
    .B(_0535_));
 sg13g2_nand2_1 _3461_ (.Y(_0537_),
    .A(_0536_),
    .B(net136));
 sg13g2_nand2_1 _3462_ (.Y(_0538_),
    .A(_0011_),
    .B(net184));
 sg13g2_nand2_1 _3463_ (.Y(_0539_),
    .A(_0537_),
    .B(_0538_));
 sg13g2_nand2_1 _3464_ (.Y(_0540_),
    .A(_0539_),
    .B(net137));
 sg13g2_nand2_1 _3465_ (.Y(_0541_),
    .A(_0010_),
    .B(net185));
 sg13g2_nand2_1 _3466_ (.Y(_0542_),
    .A(_0540_),
    .B(_0541_));
 sg13g2_nand2_1 _3467_ (.Y(_0543_),
    .A(_0542_),
    .B(_1796_));
 sg13g2_nand2_1 _3468_ (.Y(_0544_),
    .A(_0009_),
    .B(_1794_));
 sg13g2_nand2_1 _3469_ (.Y(_0545_),
    .A(_0543_),
    .B(_0544_));
 sg13g2_nand2_1 _3470_ (.Y(_0546_),
    .A(_0545_),
    .B(net118));
 sg13g2_nand2_1 _3471_ (.Y(_0547_),
    .A(_0008_),
    .B(_1788_));
 sg13g2_nand2_1 _3472_ (.Y(_0548_),
    .A(_0546_),
    .B(_0547_));
 sg13g2_nand2_1 _3473_ (.Y(_0549_),
    .A(_0548_),
    .B(net119));
 sg13g2_nand2_1 _3474_ (.Y(_0550_),
    .A(_0007_),
    .B(net174));
 sg13g2_nand2_1 _3475_ (.Y(_0551_),
    .A(_0549_),
    .B(_0550_));
 sg13g2_nand2_1 _3476_ (.Y(_0552_),
    .A(_0006_),
    .B(_1778_));
 sg13g2_inv_1 _3477_ (.Y(_0553_),
    .A(_0552_));
 sg13g2_a21oi_1 _3478_ (.A1(_0551_),
    .A2(net120),
    .Y(_0554_),
    .B1(_0553_));
 sg13g2_nand2_1 _3479_ (.Y(_0555_),
    .A(_0005_),
    .B(net153));
 sg13g2_o21ai_1 _3480_ (.B1(_0555_),
    .Y(_0556_),
    .A1(net114),
    .A2(_0554_));
 sg13g2_nand2_1 _3481_ (.Y(_0557_),
    .A(_0556_),
    .B(_1769_));
 sg13g2_nand2_1 _3482_ (.Y(_0558_),
    .A(_0004_),
    .B(_1767_));
 sg13g2_nand2_1 _3483_ (.Y(_0559_),
    .A(_0557_),
    .B(_0558_));
 sg13g2_nand2_1 _3484_ (.Y(_0560_),
    .A(_0559_),
    .B(net168));
 sg13g2_nand2_1 _3485_ (.Y(_0561_),
    .A(_0003_),
    .B(net175));
 sg13g2_nand2_1 _3486_ (.Y(_0562_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_nand2_1 _3487_ (.Y(_0563_),
    .A(_0562_),
    .B(net124));
 sg13g2_nand2_1 _3488_ (.Y(_0564_),
    .A(_0002_),
    .B(_1754_));
 sg13g2_nand2_1 _3489_ (.Y(_0565_),
    .A(_0563_),
    .B(_0564_));
 sg13g2_nand2_1 _3490_ (.Y(_0566_),
    .A(_0565_),
    .B(net103));
 sg13g2_nand2_1 _3491_ (.Y(_0567_),
    .A(_0001_),
    .B(net147));
 sg13g2_nand2_1 _3492_ (.Y(_0568_),
    .A(_0566_),
    .B(_0567_));
 sg13g2_nand2_1 _3493_ (.Y(_0569_),
    .A(_0568_),
    .B(net139));
 sg13g2_nand2_1 _3494_ (.Y(_0570_),
    .A(_0000_),
    .B(_1655_));
 sg13g2_inv_1 _3495_ (.Y(_0571_),
    .A(_0570_));
 sg13g2_nor2b_1 _3496_ (.A(_0571_),
    .B_N(_0194_),
    .Y(_0572_));
 sg13g2_nand2_1 _3497_ (.Y(_0573_),
    .A(_0569_),
    .B(_0572_));
 sg13g2_buf_1 _3498_ (.A(_1721_),
    .X(_0574_));
 sg13g2_nand2_1 _3499_ (.Y(_0575_),
    .A(\ayayayayayaya.b[15] ),
    .B(_1586_));
 sg13g2_inv_1 _3500_ (.Y(_0576_),
    .A(_0529_));
 sg13g2_a21oi_1 _3501_ (.A1(_0575_),
    .A2(_1694_),
    .Y(_0577_),
    .B1(_0576_));
 sg13g2_o21ai_1 _3502_ (.B1(_0532_),
    .Y(_0578_),
    .A1(_1688_),
    .A2(_0577_));
 sg13g2_inv_1 _3503_ (.Y(_0579_),
    .A(_0535_));
 sg13g2_a21oi_1 _3504_ (.A1(_0578_),
    .A2(_1684_),
    .Y(_0580_),
    .B1(_0579_));
 sg13g2_o21ai_1 _3505_ (.B1(_0538_),
    .Y(_0581_),
    .A1(net184),
    .A2(_0580_));
 sg13g2_inv_1 _3506_ (.Y(_0582_),
    .A(_0541_));
 sg13g2_a21oi_1 _3507_ (.A1(_0581_),
    .A2(net137),
    .Y(_0583_),
    .B1(_0582_));
 sg13g2_o21ai_1 _3508_ (.B1(_0544_),
    .Y(_0584_),
    .A1(net161),
    .A2(_0583_));
 sg13g2_inv_1 _3509_ (.Y(_0585_),
    .A(_0547_));
 sg13g2_a21oi_1 _3510_ (.A1(_0584_),
    .A2(_1789_),
    .Y(_0586_),
    .B1(_0585_));
 sg13g2_o21ai_1 _3511_ (.B1(_0550_),
    .Y(_0587_),
    .A1(net174),
    .A2(_0586_));
 sg13g2_a21oi_1 _3512_ (.A1(_0587_),
    .A2(_1779_),
    .Y(_0588_),
    .B1(_0553_));
 sg13g2_o21ai_1 _3513_ (.B1(_0555_),
    .Y(_0589_),
    .A1(net153),
    .A2(_0588_));
 sg13g2_inv_1 _3514_ (.Y(_0590_),
    .A(_0558_));
 sg13g2_a21oi_1 _3515_ (.A1(_0589_),
    .A2(net122),
    .Y(_0591_),
    .B1(_0590_));
 sg13g2_o21ai_1 _3516_ (.B1(_0561_),
    .Y(_0592_),
    .A1(_2214_),
    .A2(_0591_));
 sg13g2_inv_1 _3517_ (.Y(_0593_),
    .A(_0564_));
 sg13g2_a21oi_1 _3518_ (.A1(_0592_),
    .A2(net97),
    .Y(_0594_),
    .B1(_0593_));
 sg13g2_o21ai_1 _3519_ (.B1(_0567_),
    .Y(_0595_),
    .A1(net141),
    .A2(_0594_));
 sg13g2_buf_1 _3520_ (.A(net171),
    .X(_0596_));
 sg13g2_a21oi_1 _3521_ (.A1(_0595_),
    .A2(net93),
    .Y(_0597_),
    .B1(_0571_));
 sg13g2_buf_1 _3522_ (.A(net62),
    .X(_0598_));
 sg13g2_and3_1 _3523_ (.X(_0599_),
    .A(net172),
    .B(_1606_),
    .C(net187));
 sg13g2_nor2_1 _3524_ (.A(_1606_),
    .B(net187),
    .Y(_0600_));
 sg13g2_nor3_1 _3525_ (.A(net145),
    .B(_0600_),
    .C(_0599_),
    .Y(_0601_));
 sg13g2_a221oi_1 _3526_ (.B2(_0599_),
    .C1(_0601_),
    .B1(net188),
    .A1(_0168_),
    .Y(_0602_),
    .A2(net65));
 sg13g2_nand2_1 _3527_ (.Y(_0603_),
    .A(net37),
    .B(_0132_));
 sg13g2_buf_1 _3528_ (.A(_1655_),
    .X(_0604_));
 sg13g2_a22oi_1 _3529_ (.Y(_0605_),
    .B1(net140),
    .B2(net42),
    .A2(net187),
    .A1(_1369_));
 sg13g2_nand3_1 _3530_ (.B(_0603_),
    .C(_0605_),
    .A(_0602_),
    .Y(_0606_));
 sg13g2_a21oi_1 _3531_ (.A1(_0597_),
    .A2(net45),
    .Y(_0607_),
    .B1(_0606_));
 sg13g2_nand2_1 _3532_ (.Y(_0608_),
    .A(_0573_),
    .B(_0607_));
 sg13g2_nand3_1 _3533_ (.B(_0450_),
    .C(_2207_),
    .A(_0433_),
    .Y(_0609_));
 sg13g2_nand3_1 _3534_ (.B(_0449_),
    .C(net79),
    .A(_0434_),
    .Y(_0610_));
 sg13g2_nand3_1 _3535_ (.B(_0448_),
    .C(net78),
    .A(_0435_),
    .Y(_0611_));
 sg13g2_nand3_1 _3536_ (.B(_0447_),
    .C(net91),
    .A(_0436_),
    .Y(_0612_));
 sg13g2_nand3_1 _3537_ (.B(_0446_),
    .C(net136),
    .A(_0437_),
    .Y(_0613_));
 sg13g2_nand3_1 _3538_ (.B(_0445_),
    .C(_1685_),
    .A(_0438_),
    .Y(_0614_));
 sg13g2_nand3_1 _3539_ (.B(_0444_),
    .C(net88),
    .A(_0439_),
    .Y(_0615_));
 sg13g2_nand3_1 _3540_ (.B(_0443_),
    .C(net87),
    .A(_0440_),
    .Y(_0616_));
 sg13g2_nand3_1 _3541_ (.B(net182),
    .C(_0527_),
    .A(_0526_),
    .Y(_0617_));
 sg13g2_nand3_1 _3542_ (.B(_0617_),
    .C(_1905_),
    .A(_0616_),
    .Y(_0618_));
 sg13g2_nand3_1 _3543_ (.B(_0618_),
    .C(_1954_),
    .A(_0615_),
    .Y(_0619_));
 sg13g2_nand3_1 _3544_ (.B(_0619_),
    .C(_1985_),
    .A(_0614_),
    .Y(_0620_));
 sg13g2_nand3_1 _3545_ (.B(_0620_),
    .C(net160),
    .A(_0613_),
    .Y(_0621_));
 sg13g2_nand3_1 _3546_ (.B(_0621_),
    .C(net116),
    .A(_0612_),
    .Y(_0622_));
 sg13g2_nand3_1 _3547_ (.B(_0622_),
    .C(net111),
    .A(_0611_),
    .Y(_0623_));
 sg13g2_nand3_1 _3548_ (.B(_0623_),
    .C(net113),
    .A(_0610_),
    .Y(_0624_));
 sg13g2_nand3_1 _3549_ (.B(_0624_),
    .C(net68),
    .A(_0609_),
    .Y(_0625_));
 sg13g2_nand3_1 _3550_ (.B(_0623_),
    .C(net74),
    .A(_0610_),
    .Y(_0626_));
 sg13g2_nand3_1 _3551_ (.B(_0622_),
    .C(net79),
    .A(_0611_),
    .Y(_0627_));
 sg13g2_nand3_1 _3552_ (.B(_0621_),
    .C(_1797_),
    .A(_0612_),
    .Y(_0628_));
 sg13g2_nand3_1 _3553_ (.B(_0620_),
    .C(net91),
    .A(_0613_),
    .Y(_0629_));
 sg13g2_nand3_1 _3554_ (.B(_0619_),
    .C(_1680_),
    .A(_0614_),
    .Y(_0630_));
 sg13g2_nand3_1 _3555_ (.B(_0618_),
    .C(_1685_),
    .A(_0615_),
    .Y(_0631_));
 sg13g2_nand3_1 _3556_ (.B(_0617_),
    .C(net134),
    .A(_0616_),
    .Y(_0632_));
 sg13g2_nand3_1 _3557_ (.B(_1905_),
    .C(_0529_),
    .A(_0528_),
    .Y(_0633_));
 sg13g2_nand3_1 _3558_ (.B(_0633_),
    .C(net162),
    .A(_0632_),
    .Y(_0634_));
 sg13g2_nand3_1 _3559_ (.B(_0634_),
    .C(net159),
    .A(_0631_),
    .Y(_0635_));
 sg13g2_nand3_1 _3560_ (.B(_0635_),
    .C(_1974_),
    .A(_0630_),
    .Y(_0636_));
 sg13g2_nand3_1 _3561_ (.B(_0636_),
    .C(net116),
    .A(_0629_),
    .Y(_0637_));
 sg13g2_nand3_1 _3562_ (.B(_0637_),
    .C(net111),
    .A(_0628_),
    .Y(_0638_));
 sg13g2_nand3_1 _3563_ (.B(_0638_),
    .C(net113),
    .A(_0627_),
    .Y(_0639_));
 sg13g2_nand3_1 _3564_ (.B(_0639_),
    .C(net115),
    .A(_0626_),
    .Y(_0640_));
 sg13g2_nand3_1 _3565_ (.B(_0640_),
    .C(net82),
    .A(_0625_),
    .Y(_0641_));
 sg13g2_nand3_1 _3566_ (.B(_0638_),
    .C(_1786_),
    .A(_0627_),
    .Y(_0642_));
 sg13g2_nand3_1 _3567_ (.B(_0636_),
    .C(net51),
    .A(_0629_),
    .Y(_0643_));
 sg13g2_nand3_1 _3568_ (.B(_0634_),
    .C(net90),
    .A(_0631_),
    .Y(_0644_));
 sg13g2_nand2_1 _3569_ (.Y(_0645_),
    .A(_0533_),
    .B(_0197_));
 sg13g2_nand3_1 _3570_ (.B(_0633_),
    .C(_1686_),
    .A(_0632_),
    .Y(_0646_));
 sg13g2_nand3_1 _3571_ (.B(_0646_),
    .C(net99),
    .A(_0645_),
    .Y(_0647_));
 sg13g2_nand3_1 _3572_ (.B(_0647_),
    .C(net98),
    .A(_0644_),
    .Y(_0648_));
 sg13g2_nand3_1 _3573_ (.B(_0635_),
    .C(_1672_),
    .A(_0630_),
    .Y(_0649_));
 sg13g2_nand3_1 _3574_ (.B(_0649_),
    .C(net61),
    .A(_0648_),
    .Y(_0650_));
 sg13g2_nand3_1 _3575_ (.B(_0650_),
    .C(net75),
    .A(_0643_),
    .Y(_0651_));
 sg13g2_nand3_1 _3576_ (.B(_0637_),
    .C(net52),
    .A(_0628_),
    .Y(_0652_));
 sg13g2_nand3_1 _3577_ (.B(_0652_),
    .C(net113),
    .A(_0651_),
    .Y(_0653_));
 sg13g2_nand3_1 _3578_ (.B(_0653_),
    .C(_0375_),
    .A(_0642_),
    .Y(_0654_));
 sg13g2_nand3_1 _3579_ (.B(_0639_),
    .C(net68),
    .A(_0626_),
    .Y(_0655_));
 sg13g2_nand3_1 _3580_ (.B(_0655_),
    .C(net77),
    .A(_0654_),
    .Y(_0656_));
 sg13g2_nand3_1 _3581_ (.B(_0656_),
    .C(net53),
    .A(_0641_),
    .Y(_0657_));
 sg13g2_nand3_1 _3582_ (.B(_0655_),
    .C(net69),
    .A(_0654_),
    .Y(_0658_));
 sg13g2_nand3_1 _3583_ (.B(_0653_),
    .C(net81),
    .A(_0642_),
    .Y(_0659_));
 sg13g2_nand3_1 _3584_ (.B(_0652_),
    .C(net74),
    .A(_0651_),
    .Y(_0660_));
 sg13g2_nand3_1 _3585_ (.B(_0650_),
    .C(net52),
    .A(_0643_),
    .Y(_0661_));
 sg13g2_nand3_1 _3586_ (.B(_0649_),
    .C(_1797_),
    .A(_0648_),
    .Y(_0662_));
 sg13g2_nand3_1 _3587_ (.B(_0647_),
    .C(_1672_),
    .A(_0644_),
    .Y(_0663_));
 sg13g2_nand3_1 _3588_ (.B(_0646_),
    .C(_1680_),
    .A(_0645_),
    .Y(_0664_));
 sg13g2_nand3_1 _3589_ (.B(net159),
    .C(_0535_),
    .A(_0534_),
    .Y(_0665_));
 sg13g2_nand3_1 _3590_ (.B(_0665_),
    .C(net160),
    .A(_0664_),
    .Y(_0666_));
 sg13g2_nand3_1 _3591_ (.B(_0666_),
    .C(net116),
    .A(_0663_),
    .Y(_0667_));
 sg13g2_nand3_1 _3592_ (.B(_0667_),
    .C(_2201_),
    .A(_0662_),
    .Y(_0668_));
 sg13g2_nand3_1 _3593_ (.B(_0668_),
    .C(net113),
    .A(_0661_),
    .Y(_0669_));
 sg13g2_nand3_1 _3594_ (.B(_0669_),
    .C(net73),
    .A(_0660_),
    .Y(_0670_));
 sg13g2_nand3_1 _3595_ (.B(_0670_),
    .C(_2098_),
    .A(_0659_),
    .Y(_0671_));
 sg13g2_nand3_1 _3596_ (.B(_0671_),
    .C(net67),
    .A(_0658_),
    .Y(_0672_));
 sg13g2_nand3_1 _3597_ (.B(_0672_),
    .C(_1765_),
    .A(_0657_),
    .Y(_0673_));
 sg13g2_nand3_1 _3598_ (.B(_0670_),
    .C(_1776_),
    .A(_0659_),
    .Y(_0674_));
 sg13g2_nand3_1 _3599_ (.B(_0668_),
    .C(_1786_),
    .A(_0661_),
    .Y(_0675_));
 sg13g2_nand3_1 _3600_ (.B(_0666_),
    .C(net51),
    .A(_0663_),
    .Y(_0676_));
 sg13g2_nand2_1 _3601_ (.Y(_0677_),
    .A(_0539_),
    .B(net98));
 sg13g2_nand3_1 _3602_ (.B(_0665_),
    .C(net91),
    .A(_0664_),
    .Y(_0678_));
 sg13g2_nand3_1 _3603_ (.B(_0678_),
    .C(net116),
    .A(_0677_),
    .Y(_0679_));
 sg13g2_nand3_1 _3604_ (.B(_0679_),
    .C(net111),
    .A(_0676_),
    .Y(_0680_));
 sg13g2_nand3_1 _3605_ (.B(_0667_),
    .C(_1791_),
    .A(_0662_),
    .Y(_0681_));
 sg13g2_nand3_1 _3606_ (.B(_0681_),
    .C(_2112_),
    .A(_0680_),
    .Y(_0682_));
 sg13g2_nand3_1 _3607_ (.B(_0682_),
    .C(_0375_),
    .A(_0675_),
    .Y(_0683_));
 sg13g2_nand3_1 _3608_ (.B(_0669_),
    .C(net68),
    .A(_0660_),
    .Y(_0684_));
 sg13g2_nand3_1 _3609_ (.B(_0684_),
    .C(_2098_),
    .A(_0683_),
    .Y(_0685_));
 sg13g2_nand3_1 _3610_ (.B(_0685_),
    .C(_2127_),
    .A(_0674_),
    .Y(_0686_));
 sg13g2_nand3_1 _3611_ (.B(_0671_),
    .C(net47),
    .A(_0658_),
    .Y(_0687_));
 sg13g2_nand3_1 _3612_ (.B(_0687_),
    .C(net71),
    .A(_0686_),
    .Y(_0688_));
 sg13g2_nand3_1 _3613_ (.B(_0688_),
    .C(net58),
    .A(_0673_),
    .Y(_0689_));
 sg13g2_nand3_1 _3614_ (.B(_0687_),
    .C(net59),
    .A(_0686_),
    .Y(_0690_));
 sg13g2_nand3_1 _3615_ (.B(_0685_),
    .C(net47),
    .A(_0674_),
    .Y(_0691_));
 sg13g2_nand3_1 _3616_ (.B(_0684_),
    .C(_2247_),
    .A(_0683_),
    .Y(_0692_));
 sg13g2_nand3_1 _3617_ (.B(_0682_),
    .C(net68),
    .A(_0675_),
    .Y(_0693_));
 sg13g2_nand3_1 _3618_ (.B(_0681_),
    .C(net74),
    .A(_0680_),
    .Y(_0694_));
 sg13g2_nand3_1 _3619_ (.B(_0679_),
    .C(net79),
    .A(_0676_),
    .Y(_0695_));
 sg13g2_nand3_1 _3620_ (.B(_0678_),
    .C(net78),
    .A(_0677_),
    .Y(_0696_));
 sg13g2_nand3_1 _3621_ (.B(net116),
    .C(_0541_),
    .A(_0540_),
    .Y(_0697_));
 sg13g2_nand3_1 _3622_ (.B(_0697_),
    .C(net111),
    .A(_0696_),
    .Y(_0698_));
 sg13g2_nand3_1 _3623_ (.B(_0698_),
    .C(_2112_),
    .A(_0695_),
    .Y(_0699_));
 sg13g2_nand3_1 _3624_ (.B(_0699_),
    .C(net73),
    .A(_0694_),
    .Y(_0700_));
 sg13g2_nand3_1 _3625_ (.B(_0700_),
    .C(net77),
    .A(_0693_),
    .Y(_0701_));
 sg13g2_nand3_1 _3626_ (.B(_0701_),
    .C(net112),
    .A(_0692_),
    .Y(_0702_));
 sg13g2_nand3_1 _3627_ (.B(_0702_),
    .C(net66),
    .A(_0691_),
    .Y(_0703_));
 sg13g2_nand3_1 _3628_ (.B(_0703_),
    .C(net108),
    .A(_0690_),
    .Y(_0704_));
 sg13g2_nand3_1 _3629_ (.B(_0704_),
    .C(net57),
    .A(_0689_),
    .Y(_0705_));
 sg13g2_nand3_1 _3630_ (.B(_0703_),
    .C(net58),
    .A(_0690_),
    .Y(_0706_));
 sg13g2_nand3_1 _3631_ (.B(_0702_),
    .C(net59),
    .A(_0691_),
    .Y(_0707_));
 sg13g2_nand3_1 _3632_ (.B(_0701_),
    .C(net47),
    .A(_0692_),
    .Y(_0708_));
 sg13g2_nand3_1 _3633_ (.B(_0700_),
    .C(net69),
    .A(_0693_),
    .Y(_0709_));
 sg13g2_nand3_1 _3634_ (.B(_0699_),
    .C(net68),
    .A(_0694_),
    .Y(_0710_));
 sg13g2_nand3_1 _3635_ (.B(_0698_),
    .C(_2207_),
    .A(_0695_),
    .Y(_0711_));
 sg13g2_nand2_1 _3636_ (.Y(_0712_),
    .A(_0545_),
    .B(net75));
 sg13g2_nand3_1 _3637_ (.B(_0697_),
    .C(_1791_),
    .A(_0696_),
    .Y(_0713_));
 sg13g2_nand3_1 _3638_ (.B(_0713_),
    .C(net113),
    .A(_0712_),
    .Y(_0714_));
 sg13g2_nand3_1 _3639_ (.B(_0714_),
    .C(net73),
    .A(_0711_),
    .Y(_0715_));
 sg13g2_nand3_1 _3640_ (.B(_0715_),
    .C(net77),
    .A(_0710_),
    .Y(_0716_));
 sg13g2_nand3_1 _3641_ (.B(_0716_),
    .C(_2126_),
    .A(_0709_),
    .Y(_0717_));
 sg13g2_nand3_1 _3642_ (.B(_0717_),
    .C(net66),
    .A(_0708_),
    .Y(_0718_));
 sg13g2_nand3_1 _3643_ (.B(_0718_),
    .C(net108),
    .A(_0707_),
    .Y(_0719_));
 sg13g2_nand3_1 _3644_ (.B(_0719_),
    .C(net141),
    .A(_0706_),
    .Y(_0720_));
 sg13g2_nand3_1 _3645_ (.B(_0720_),
    .C(net139),
    .A(_0705_),
    .Y(_0721_));
 sg13g2_nand3_1 _3646_ (.B(_0719_),
    .C(net86),
    .A(_0706_),
    .Y(_0722_));
 sg13g2_nand3_1 _3647_ (.B(_0718_),
    .C(net85),
    .A(_0707_),
    .Y(_0723_));
 sg13g2_nand3_1 _3648_ (.B(_0717_),
    .C(net59),
    .A(_0708_),
    .Y(_0724_));
 sg13g2_nand3_1 _3649_ (.B(_0716_),
    .C(net53),
    .A(_0709_),
    .Y(_0725_));
 sg13g2_nand3_1 _3650_ (.B(_0715_),
    .C(net69),
    .A(_0710_),
    .Y(_0726_));
 sg13g2_nand3_1 _3651_ (.B(_0714_),
    .C(_1781_),
    .A(_0711_),
    .Y(_0727_));
 sg13g2_nand3_1 _3652_ (.B(_0713_),
    .C(net74),
    .A(_0712_),
    .Y(_0728_));
 sg13g2_nand3_1 _3653_ (.B(net113),
    .C(_0547_),
    .A(_0546_),
    .Y(_0729_));
 sg13g2_nand3_1 _3654_ (.B(_0729_),
    .C(net73),
    .A(_0728_),
    .Y(_0730_));
 sg13g2_nand3_1 _3655_ (.B(_0730_),
    .C(net77),
    .A(_0727_),
    .Y(_0731_));
 sg13g2_nand3_1 _3656_ (.B(_0731_),
    .C(net67),
    .A(_0726_),
    .Y(_0732_));
 sg13g2_nand3_1 _3657_ (.B(_0732_),
    .C(net66),
    .A(_0725_),
    .Y(_0733_));
 sg13g2_nand3_1 _3658_ (.B(_0733_),
    .C(net107),
    .A(_0724_),
    .Y(_0734_));
 sg13g2_nand3_1 _3659_ (.B(_0734_),
    .C(_0171_),
    .A(_0723_),
    .Y(_0735_));
 sg13g2_nand3_1 _3660_ (.B(_0735_),
    .C(_0493_),
    .A(_0722_),
    .Y(_0736_));
 sg13g2_nand3_1 _3661_ (.B(_0736_),
    .C(net46),
    .A(_0721_),
    .Y(_0737_));
 sg13g2_inv_2 _3662_ (.Y(_0738_),
    .A(_0215_));
 sg13g2_a22oi_1 _3663_ (.Y(_0739_),
    .B1(_2127_),
    .B2(net65),
    .A2(_2202_),
    .A1(_0213_));
 sg13g2_o21ai_1 _3664_ (.B1(_0739_),
    .Y(_0740_),
    .A1(_1728_),
    .A2(_0738_));
 sg13g2_nand2_1 _3665_ (.Y(_0741_),
    .A(net172),
    .B(_1652_));
 sg13g2_o21ai_1 _3666_ (.B1(\a[9] ),
    .Y(_0742_),
    .A1(_0741_),
    .A2(_1293_));
 sg13g2_a21oi_1 _3667_ (.A1(net94),
    .A2(_0741_),
    .Y(_0743_),
    .B1(_0742_));
 sg13g2_buf_1 _3668_ (.A(net56),
    .X(_0744_));
 sg13g2_inv_1 _3669_ (.Y(_0745_),
    .A(\a[9] ));
 sg13g2_nand2_1 _3670_ (.Y(_0746_),
    .A(net63),
    .B(_0745_));
 sg13g2_inv_1 _3671_ (.Y(_0747_),
    .A(_1652_));
 sg13g2_a21oi_1 _3672_ (.A1(_0744_),
    .A2(_0746_),
    .Y(_0748_),
    .B1(_0747_));
 sg13g2_inv_1 _3673_ (.Y(_0749_),
    .A(net62));
 sg13g2_nor2_1 _3674_ (.A(net133),
    .B(_0575_),
    .Y(_0750_));
 sg13g2_mux2_1 _3675_ (.A0(_0750_),
    .A1(_0577_),
    .S(_1688_),
    .X(_0751_));
 sg13g2_nand2b_1 _3676_ (.Y(_0752_),
    .B(_0750_),
    .A_N(_0044_));
 sg13g2_nor2_1 _3677_ (.A(net183),
    .B(_0752_),
    .Y(_0753_));
 sg13g2_a21oi_1 _3678_ (.A1(_0751_),
    .A2(net183),
    .Y(_0754_),
    .B1(_0753_));
 sg13g2_nor2_1 _3679_ (.A(net183),
    .B(_0751_),
    .Y(_0755_));
 sg13g2_a21oi_1 _3680_ (.A1(net183),
    .A2(_0578_),
    .Y(_0756_),
    .B1(_0755_));
 sg13g2_nor2_1 _3681_ (.A(_1679_),
    .B(_0756_),
    .Y(_0757_));
 sg13g2_a21oi_1 _3682_ (.A1(_1679_),
    .A2(_0754_),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_inv_1 _3683_ (.Y(_0759_),
    .A(_0758_));
 sg13g2_mux2_1 _3684_ (.A0(_0580_),
    .A1(_0756_),
    .S(_1679_),
    .X(_0760_));
 sg13g2_nor2_1 _3685_ (.A(_1671_),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_a21oi_1 _3686_ (.A1(net137),
    .A2(_0759_),
    .Y(_0762_),
    .B1(_0761_));
 sg13g2_nor2_1 _3687_ (.A(_1670_),
    .B(_0581_),
    .Y(_0763_));
 sg13g2_a21oi_1 _3688_ (.A1(_0760_),
    .A2(_1670_),
    .Y(_0764_),
    .B1(_0763_));
 sg13g2_nor2_1 _3689_ (.A(_1795_),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_a21o_1 _3690_ (.A2(net117),
    .A1(_0762_),
    .B1(_0765_),
    .X(_0766_));
 sg13g2_nor2_1 _3691_ (.A(_0043_),
    .B(_0752_),
    .Y(_0767_));
 sg13g2_nor2_1 _3692_ (.A(net184),
    .B(_0767_),
    .Y(_0768_));
 sg13g2_a21oi_1 _3693_ (.A1(_0754_),
    .A2(net184),
    .Y(_0769_),
    .B1(_0768_));
 sg13g2_nand2_1 _3694_ (.Y(_0770_),
    .A(_0769_),
    .B(_1670_));
 sg13g2_o21ai_1 _3695_ (.B1(_0770_),
    .Y(_0771_),
    .A1(_1670_),
    .A2(_0759_));
 sg13g2_nor2b_1 _3696_ (.A(net161),
    .B_N(_0771_),
    .Y(_0772_));
 sg13g2_a21o_1 _3697_ (.A2(net161),
    .A1(_0762_),
    .B1(_0772_),
    .X(_0773_));
 sg13g2_mux2_1 _3698_ (.A0(_0766_),
    .A1(_0773_),
    .S(net118),
    .X(_0774_));
 sg13g2_nand2b_1 _3699_ (.Y(_0775_),
    .B(_0767_),
    .A_N(_0042_));
 sg13g2_nor2_1 _3700_ (.A(net185),
    .B(_0775_),
    .Y(_0776_));
 sg13g2_a21oi_1 _3701_ (.A1(_0769_),
    .A2(net185),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_nor2_1 _3702_ (.A(_1795_),
    .B(_0771_),
    .Y(_0778_));
 sg13g2_a21oi_1 _3703_ (.A1(_1795_),
    .A2(_0777_),
    .Y(_0779_),
    .B1(_0778_));
 sg13g2_inv_1 _3704_ (.Y(_0780_),
    .A(_0779_));
 sg13g2_nor2_1 _3705_ (.A(net156),
    .B(_0780_),
    .Y(_0781_));
 sg13g2_a21o_1 _3706_ (.A2(net156),
    .A1(_0773_),
    .B1(_0781_),
    .X(_0782_));
 sg13g2_mux2_1 _3707_ (.A0(_0774_),
    .A1(_0782_),
    .S(_1784_),
    .X(_0783_));
 sg13g2_nor2_1 _3708_ (.A(_0041_),
    .B(_0775_),
    .Y(_0784_));
 sg13g2_nor2_1 _3709_ (.A(_1794_),
    .B(_0784_),
    .Y(_0785_));
 sg13g2_a21oi_1 _3710_ (.A1(_0777_),
    .A2(_1794_),
    .Y(_0786_),
    .B1(_0785_));
 sg13g2_nand2_1 _3711_ (.Y(_0787_),
    .A(_0786_),
    .B(_1789_));
 sg13g2_o21ai_1 _3712_ (.B1(_0787_),
    .Y(_0788_),
    .A1(_1789_),
    .A2(_0780_));
 sg13g2_nor2b_1 _3713_ (.A(net174),
    .B_N(_0788_),
    .Y(_0789_));
 sg13g2_a21o_1 _3714_ (.A2(net155),
    .A1(_0782_),
    .B1(_0789_),
    .X(_0790_));
 sg13g2_nor2b_1 _3715_ (.A(net154),
    .B_N(_0790_),
    .Y(_0791_));
 sg13g2_a21o_1 _3716_ (.A2(net154),
    .A1(_0783_),
    .B1(_0791_),
    .X(_0792_));
 sg13g2_nand2b_1 _3717_ (.Y(_0793_),
    .B(_0784_),
    .A_N(_0040_));
 sg13g2_nor2_1 _3718_ (.A(_1788_),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_a21oi_1 _3719_ (.A1(_0786_),
    .A2(_1788_),
    .Y(_0795_),
    .B1(_0794_));
 sg13g2_nor2_1 _3720_ (.A(_1784_),
    .B(_0788_),
    .Y(_0796_));
 sg13g2_a21oi_1 _3721_ (.A1(_1784_),
    .A2(_0795_),
    .Y(_0797_),
    .B1(_0796_));
 sg13g2_inv_1 _3722_ (.Y(_0798_),
    .A(_0797_));
 sg13g2_nor2_1 _3723_ (.A(_1778_),
    .B(_0798_),
    .Y(_0799_));
 sg13g2_a21o_1 _3724_ (.A2(net154),
    .A1(_0790_),
    .B1(_0799_),
    .X(_0800_));
 sg13g2_nor2b_1 _3725_ (.A(_1773_),
    .B_N(_0800_),
    .Y(_0801_));
 sg13g2_a21o_1 _3726_ (.A2(net153),
    .A1(_0792_),
    .B1(_0801_),
    .X(_0802_));
 sg13g2_nor2_1 _3727_ (.A(_0039_),
    .B(_0793_),
    .Y(_0803_));
 sg13g2_nor2_1 _3728_ (.A(_1783_),
    .B(_0803_),
    .Y(_0804_));
 sg13g2_a21oi_1 _3729_ (.A1(_0795_),
    .A2(net155),
    .Y(_0805_),
    .B1(_0804_));
 sg13g2_nand2_1 _3730_ (.Y(_0806_),
    .A(_0805_),
    .B(_1779_));
 sg13g2_o21ai_1 _3731_ (.B1(_0806_),
    .Y(_0807_),
    .A1(_1779_),
    .A2(_0798_));
 sg13g2_nor2b_1 _3732_ (.A(net153),
    .B_N(_0807_),
    .Y(_0808_));
 sg13g2_a21o_1 _3733_ (.A2(net153),
    .A1(_0800_),
    .B1(_0808_),
    .X(_0809_));
 sg13g2_nor2b_1 _3734_ (.A(_1767_),
    .B_N(_0809_),
    .Y(_0810_));
 sg13g2_a21o_1 _3735_ (.A2(net152),
    .A1(_0802_),
    .B1(_0810_),
    .X(_0811_));
 sg13g2_nand2_1 _3736_ (.Y(_0812_),
    .A(_0803_),
    .B(_0179_));
 sg13g2_nor2_1 _3737_ (.A(net154),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_a21oi_1 _3738_ (.A1(_0805_),
    .A2(_2092_),
    .Y(_0814_),
    .B1(_0813_));
 sg13g2_nor2_1 _3739_ (.A(net167),
    .B(_0807_),
    .Y(_0815_));
 sg13g2_a21oi_1 _3740_ (.A1(net167),
    .A2(_0814_),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_inv_1 _3741_ (.Y(_0817_),
    .A(_0816_));
 sg13g2_nor2_1 _3742_ (.A(_1767_),
    .B(_0817_),
    .Y(_0818_));
 sg13g2_a21o_1 _3743_ (.A2(net152),
    .A1(_0809_),
    .B1(_0818_),
    .X(_0819_));
 sg13g2_nor2b_1 _3744_ (.A(net175),
    .B_N(_0819_),
    .Y(_0820_));
 sg13g2_a21o_1 _3745_ (.A2(net150),
    .A1(_0811_),
    .B1(_0820_),
    .X(_0821_));
 sg13g2_nor2_1 _3746_ (.A(net117),
    .B(_0583_),
    .Y(_0822_));
 sg13g2_a21oi_1 _3747_ (.A1(_0764_),
    .A2(net117),
    .Y(_0823_),
    .B1(_0822_));
 sg13g2_nor2b_1 _3748_ (.A(_1788_),
    .B_N(_0766_),
    .Y(_0824_));
 sg13g2_a21o_1 _3749_ (.A2(_0823_),
    .A1(_1788_),
    .B1(_0824_),
    .X(_0825_));
 sg13g2_mux2_1 _3750_ (.A0(_0774_),
    .A1(_0825_),
    .S(net174),
    .X(_0826_));
 sg13g2_inv_1 _3751_ (.Y(_0827_),
    .A(_0826_));
 sg13g2_nor2_1 _3752_ (.A(net154),
    .B(_0783_),
    .Y(_0828_));
 sg13g2_a21oi_1 _3753_ (.A1(_0827_),
    .A2(net154),
    .Y(_0829_),
    .B1(_0828_));
 sg13g2_mux2_1 _3754_ (.A0(_0829_),
    .A1(_0792_),
    .S(net167),
    .X(_0830_));
 sg13g2_nor2b_1 _3755_ (.A(_1767_),
    .B_N(_0802_),
    .Y(_0831_));
 sg13g2_a21o_1 _3756_ (.A2(net152),
    .A1(_0830_),
    .B1(_0831_),
    .X(_0832_));
 sg13g2_nor2b_1 _3757_ (.A(net150),
    .B_N(_0811_),
    .Y(_0833_));
 sg13g2_a21o_1 _3758_ (.A2(net150),
    .A1(_0832_),
    .B1(_0833_),
    .X(_0834_));
 sg13g2_mux2_1 _3759_ (.A0(_0821_),
    .A1(_0834_),
    .S(net149),
    .X(_0835_));
 sg13g2_nor2_1 _3760_ (.A(_1789_),
    .B(_0584_),
    .Y(_0836_));
 sg13g2_a21oi_1 _3761_ (.A1(_0823_),
    .A2(net118),
    .Y(_0837_),
    .B1(_0836_));
 sg13g2_nor2_1 _3762_ (.A(net174),
    .B(_0825_),
    .Y(_0838_));
 sg13g2_a21oi_1 _3763_ (.A1(net174),
    .A2(_0837_),
    .Y(_0839_),
    .B1(_0838_));
 sg13g2_nor2_1 _3764_ (.A(net154),
    .B(_0827_),
    .Y(_0840_));
 sg13g2_a21o_1 _3765_ (.A2(_0839_),
    .A1(net154),
    .B1(_0840_),
    .X(_0841_));
 sg13g2_inv_1 _3766_ (.Y(_0842_),
    .A(_0841_));
 sg13g2_nor2_1 _3767_ (.A(net153),
    .B(_0829_),
    .Y(_0843_));
 sg13g2_a21oi_1 _3768_ (.A1(_0842_),
    .A2(net153),
    .Y(_0844_),
    .B1(_0843_));
 sg13g2_inv_1 _3769_ (.Y(_0845_),
    .A(_0844_));
 sg13g2_nor2_1 _3770_ (.A(net152),
    .B(_0830_),
    .Y(_0846_));
 sg13g2_a21oi_1 _3771_ (.A1(net152),
    .A2(_0845_),
    .Y(_0847_),
    .B1(_0846_));
 sg13g2_nor2b_1 _3772_ (.A(net175),
    .B_N(_0832_),
    .Y(_0848_));
 sg13g2_a21o_1 _3773_ (.A2(_0847_),
    .A1(net150),
    .B1(_0848_),
    .X(_0849_));
 sg13g2_mux2_1 _3774_ (.A0(_0834_),
    .A1(_0849_),
    .S(net149),
    .X(_0850_));
 sg13g2_mux2_1 _3775_ (.A0(_0835_),
    .A1(_0850_),
    .S(net147),
    .X(_0851_));
 sg13g2_nor2_1 _3776_ (.A(net140),
    .B(_0851_),
    .Y(_0852_));
 sg13g2_nor2_1 _3777_ (.A(_1784_),
    .B(_0586_),
    .Y(_0853_));
 sg13g2_a21oi_1 _3778_ (.A1(_0837_),
    .A2(_1784_),
    .Y(_0854_),
    .B1(_0853_));
 sg13g2_nor2b_1 _3779_ (.A(_1779_),
    .B_N(_0854_),
    .Y(_0855_));
 sg13g2_a21o_1 _3780_ (.A2(_1779_),
    .A1(_0839_),
    .B1(_0855_),
    .X(_0856_));
 sg13g2_nor2_1 _3781_ (.A(net167),
    .B(_0856_),
    .Y(_0857_));
 sg13g2_a21oi_1 _3782_ (.A1(_0842_),
    .A2(net167),
    .Y(_0858_),
    .B1(_0857_));
 sg13g2_nor2_1 _3783_ (.A(_1767_),
    .B(_0845_),
    .Y(_0859_));
 sg13g2_a21o_1 _3784_ (.A2(_0858_),
    .A1(net152),
    .B1(_0859_),
    .X(_0860_));
 sg13g2_mux2_1 _3785_ (.A0(_0847_),
    .A1(_0860_),
    .S(net175),
    .X(_0861_));
 sg13g2_mux2_1 _3786_ (.A0(_0861_),
    .A1(_0849_),
    .S(net97),
    .X(_0862_));
 sg13g2_mux2_1 _3787_ (.A0(_0862_),
    .A1(_0850_),
    .S(net170),
    .X(_0863_));
 sg13g2_nor2_1 _3788_ (.A(net93),
    .B(_0863_),
    .Y(_0864_));
 sg13g2_nor3_1 _3789_ (.A(_0749_),
    .B(_0852_),
    .C(_0864_),
    .Y(_0865_));
 sg13g2_nor4_1 _3790_ (.A(_0740_),
    .B(_0743_),
    .C(_0748_),
    .D(_0865_),
    .Y(_0866_));
 sg13g2_nand2_1 _3791_ (.Y(_0867_),
    .A(_0737_),
    .B(_0866_));
 sg13g2_a22oi_1 _3792_ (.Y(_0868_),
    .B1(_1542_),
    .B2(_0867_),
    .A2(_0608_),
    .A1(_1412_));
 sg13g2_nand2_1 _3793_ (.Y(net13),
    .A(_0525_),
    .B(_0868_));
 sg13g2_nand2_1 _3794_ (.Y(_0869_),
    .A(_0568_),
    .B(net96));
 sg13g2_nand2_1 _3795_ (.Y(_0870_),
    .A(_0562_),
    .B(net70));
 sg13g2_nand2_1 _3796_ (.Y(_0871_),
    .A(_0556_),
    .B(net76));
 sg13g2_nand2_1 _3797_ (.Y(_0872_),
    .A(_0554_),
    .B(_2211_));
 sg13g2_nand2_1 _3798_ (.Y(_0873_),
    .A(_0551_),
    .B(net60));
 sg13g2_nand3_1 _3799_ (.B(_0729_),
    .C(net68),
    .A(_0728_),
    .Y(_0874_));
 sg13g2_nand3_1 _3800_ (.B(_0874_),
    .C(net121),
    .A(_0873_),
    .Y(_0875_));
 sg13g2_nand3_1 _3801_ (.B(_0875_),
    .C(net83),
    .A(_0872_),
    .Y(_0876_));
 sg13g2_nand3_1 _3802_ (.B(net84),
    .C(_0876_),
    .A(_0871_),
    .Y(_0877_));
 sg13g2_nand3_1 _3803_ (.B(net66),
    .C(_0558_),
    .A(_0557_),
    .Y(_0878_));
 sg13g2_nand3_1 _3804_ (.B(_0878_),
    .C(net85),
    .A(_0877_),
    .Y(_0879_));
 sg13g2_nand3_1 _3805_ (.B(_0879_),
    .C(net57),
    .A(_0870_),
    .Y(_0880_));
 sg13g2_nand3_1 _3806_ (.B(net141),
    .C(_0564_),
    .A(_0563_),
    .Y(_0881_));
 sg13g2_nand3_1 _3807_ (.B(_0881_),
    .C(net102),
    .A(_0880_),
    .Y(_0882_));
 sg13g2_nand3_1 _3808_ (.B(_0882_),
    .C(net50),
    .A(_0869_),
    .Y(_0883_));
 sg13g2_inv_1 _3809_ (.Y(_0884_),
    .A(_1637_));
 sg13g2_nand2_1 _3810_ (.Y(_0885_),
    .A(net188),
    .B(net189));
 sg13g2_o21ai_1 _3811_ (.B1(net40),
    .Y(_0886_),
    .A1(_0884_),
    .A2(_0885_));
 sg13g2_nor2_1 _3812_ (.A(_1779_),
    .B(_0587_),
    .Y(_0887_));
 sg13g2_a21oi_1 _3813_ (.A1(_0854_),
    .A2(_1779_),
    .Y(_0888_),
    .B1(_0887_));
 sg13g2_nor2_1 _3814_ (.A(net167),
    .B(_0588_),
    .Y(_0889_));
 sg13g2_a21oi_1 _3815_ (.A1(_0888_),
    .A2(net167),
    .Y(_0890_),
    .B1(_0889_));
 sg13g2_nor2_1 _3816_ (.A(net122),
    .B(_0589_),
    .Y(_0891_));
 sg13g2_a21oi_1 _3817_ (.A1(_0890_),
    .A2(net122),
    .Y(_0892_),
    .B1(_0891_));
 sg13g2_nor2_1 _3818_ (.A(net168),
    .B(_0591_),
    .Y(_0893_));
 sg13g2_a21oi_1 _3819_ (.A1(_0892_),
    .A2(net168),
    .Y(_0894_),
    .B1(_0893_));
 sg13g2_nor2_1 _3820_ (.A(net97),
    .B(_0592_),
    .Y(_0895_));
 sg13g2_a21oi_1 _3821_ (.A1(_0894_),
    .A2(_0488_),
    .Y(_0896_),
    .B1(_0895_));
 sg13g2_nor2_1 _3822_ (.A(net170),
    .B(_0594_),
    .Y(_0897_));
 sg13g2_a21oi_1 _3823_ (.A1(_0896_),
    .A2(net127),
    .Y(_0898_),
    .B1(_0897_));
 sg13g2_nor2_1 _3824_ (.A(net146),
    .B(_0898_),
    .Y(_0899_));
 sg13g2_a21oi_1 _3825_ (.A1(net140),
    .A2(_0595_),
    .Y(_0900_),
    .B1(_0899_));
 sg13g2_inv_1 _3826_ (.Y(_0901_),
    .A(_1606_));
 sg13g2_a21oi_1 _3827_ (.A1(_0901_),
    .A2(_0884_),
    .Y(_0902_),
    .B1(net145));
 sg13g2_nand3_1 _3828_ (.B(_1606_),
    .C(_1637_),
    .A(net172),
    .Y(_0903_));
 sg13g2_a22oi_1 _3829_ (.Y(_0904_),
    .B1(_1588_),
    .B2(net37),
    .A2(_0903_),
    .A1(_0902_));
 sg13g2_a22oi_1 _3830_ (.Y(_0905_),
    .B1(_1478_),
    .B2(net49),
    .A2(net104),
    .A1(net42));
 sg13g2_nand2_1 _3831_ (.Y(_0906_),
    .A(_0904_),
    .B(_0905_));
 sg13g2_a221oi_1 _3832_ (.B2(net45),
    .C1(_0906_),
    .B1(_0900_),
    .A1(_1606_),
    .Y(_0907_),
    .A2(_0886_));
 sg13g2_a21oi_1 _3833_ (.A1(_0883_),
    .A2(_0907_),
    .Y(_0908_),
    .B1(_1423_));
 sg13g2_nand3_1 _3834_ (.B(_0508_),
    .C(net96),
    .A(_0507_),
    .Y(_0909_));
 sg13g2_nand3_1 _3835_ (.B(_0506_),
    .C(net104),
    .A(_0495_),
    .Y(_0910_));
 sg13g2_nand3_1 _3836_ (.B(_0505_),
    .C(net70),
    .A(_0504_),
    .Y(_0911_));
 sg13g2_nand3_1 _3837_ (.B(_0503_),
    .C(_2216_),
    .A(_0496_),
    .Y(_0912_));
 sg13g2_nand3_1 _3838_ (.B(_0502_),
    .C(net67),
    .A(_0501_),
    .Y(_0913_));
 sg13g2_nand3_1 _3839_ (.B(_0500_),
    .C(net72),
    .A(_0497_),
    .Y(_0914_));
 sg13g2_nand3_1 _3840_ (.B(_0499_),
    .C(_2209_),
    .A(_0498_),
    .Y(_0915_));
 sg13g2_nand3_1 _3841_ (.B(_0154_),
    .C(net68),
    .A(_0153_),
    .Y(_0916_));
 sg13g2_nand3_1 _3842_ (.B(_0916_),
    .C(net69),
    .A(_0915_),
    .Y(_0917_));
 sg13g2_nand3_1 _3843_ (.B(_0917_),
    .C(net47),
    .A(_0914_),
    .Y(_0918_));
 sg13g2_nand3_1 _3844_ (.B(_0918_),
    .C(net59),
    .A(_0913_),
    .Y(_0919_));
 sg13g2_nand3_1 _3845_ (.B(_0919_),
    .C(_0489_),
    .A(_0912_),
    .Y(_0920_));
 sg13g2_nand3_1 _3846_ (.B(_0920_),
    .C(_0174_),
    .A(_0911_),
    .Y(_0921_));
 sg13g2_nand3_1 _3847_ (.B(_0921_),
    .C(net95),
    .A(_0910_),
    .Y(_0922_));
 sg13g2_nand3_1 _3848_ (.B(_0922_),
    .C(net46),
    .A(_0909_),
    .Y(_0923_));
 sg13g2_nand2_1 _3849_ (.Y(_0924_),
    .A(_0209_),
    .B(\a[18] ));
 sg13g2_inv_1 _3850_ (.Y(_0925_),
    .A(_0924_));
 sg13g2_nand2_1 _3851_ (.Y(_0926_),
    .A(_0925_),
    .B(_1597_));
 sg13g2_nand2_1 _3852_ (.Y(_0927_),
    .A(_1661_),
    .B(net151));
 sg13g2_a21oi_1 _3853_ (.A1(_0926_),
    .A2(_0927_),
    .Y(_0928_),
    .B1(net138));
 sg13g2_a22oi_1 _3854_ (.Y(_0929_),
    .B1(_1617_),
    .B2(net37),
    .A2(_1652_),
    .A1(net49));
 sg13g2_a21oi_1 _3855_ (.A1(_1598_),
    .A2(_1601_),
    .Y(_0930_),
    .B1(net94));
 sg13g2_a22oi_1 _3856_ (.Y(_0931_),
    .B1(_0926_),
    .B2(_0930_),
    .A2(_1597_),
    .A1(_1564_));
 sg13g2_nand2_1 _3857_ (.Y(_0932_),
    .A(_0929_),
    .B(_0931_));
 sg13g2_and3_1 _3858_ (.X(_0933_),
    .A(_0399_),
    .B(net45),
    .C(_0402_));
 sg13g2_nor3_1 _3859_ (.A(_0928_),
    .B(_0932_),
    .C(_0933_),
    .Y(_0934_));
 sg13g2_a21oi_1 _3860_ (.A1(_0923_),
    .A2(_0934_),
    .Y(_0935_),
    .B1(_1591_));
 sg13g2_nor2_1 _3861_ (.A(_0908_),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_buf_1 _3862_ (.A(net146),
    .X(_0937_));
 sg13g2_nand3_1 _3863_ (.B(_0186_),
    .C(net92),
    .A(_0172_),
    .Y(_0938_));
 sg13g2_nand3_1 _3864_ (.B(net141),
    .C(_0185_),
    .A(_0173_),
    .Y(_0939_));
 sg13g2_nand3_1 _3865_ (.B(net108),
    .C(_0184_),
    .A(_0175_),
    .Y(_0940_));
 sg13g2_nand3_1 _3866_ (.B(net109),
    .C(_0183_),
    .A(_0176_),
    .Y(_0941_));
 sg13g2_nand3_1 _3867_ (.B(net112),
    .C(_0182_),
    .A(_0177_),
    .Y(_0942_));
 sg13g2_nand3_1 _3868_ (.B(net114),
    .C(_0181_),
    .A(_0178_),
    .Y(_0943_));
 sg13g2_nor2_1 _3869_ (.A(_0037_),
    .B(_0180_),
    .Y(_0944_));
 sg13g2_nand2_1 _3870_ (.Y(_0945_),
    .A(_0944_),
    .B(net121));
 sg13g2_nand3_1 _3871_ (.B(net83),
    .C(_0945_),
    .A(_0943_),
    .Y(_0946_));
 sg13g2_nand3_1 _3872_ (.B(net123),
    .C(_0946_),
    .A(_0942_),
    .Y(_0947_));
 sg13g2_nand3_1 _3873_ (.B(net124),
    .C(_0947_),
    .A(_0941_),
    .Y(_0948_));
 sg13g2_nand3_1 _3874_ (.B(_1723_),
    .C(_0948_),
    .A(_0940_),
    .Y(_0949_));
 sg13g2_nand3_1 _3875_ (.B(_0187_),
    .C(_0949_),
    .A(_0939_),
    .Y(_0950_));
 sg13g2_buf_1 _3876_ (.A(_0194_),
    .X(_0951_));
 sg13g2_nand3_1 _3877_ (.B(_0950_),
    .C(net44),
    .A(_0938_),
    .Y(_0952_));
 sg13g2_nand2_1 _3878_ (.Y(_0953_),
    .A(net189),
    .B(\a[26] ));
 sg13g2_inv_1 _3879_ (.Y(_0954_),
    .A(_0953_));
 sg13g2_nand2_1 _3880_ (.Y(_0955_),
    .A(_0954_),
    .B(_1626_));
 sg13g2_nand2_1 _3881_ (.Y(_0956_),
    .A(_1661_),
    .B(net177));
 sg13g2_a21oi_1 _3882_ (.A1(_0955_),
    .A2(_0956_),
    .Y(_0957_),
    .B1(net138));
 sg13g2_a21oi_1 _3883_ (.A1(_1627_),
    .A2(_1629_),
    .Y(_0958_),
    .B1(net145));
 sg13g2_a22oi_1 _3884_ (.Y(_0959_),
    .B1(\a[28] ),
    .B2(net37),
    .A2(_0955_),
    .A1(_0958_));
 sg13g2_a22oi_1 _3885_ (.Y(_0960_),
    .B1(\a[12] ),
    .B2(net49),
    .A2(_1626_),
    .A1(_1369_));
 sg13g2_nand2_1 _3886_ (.Y(_0961_),
    .A(_0959_),
    .B(_0960_));
 sg13g2_and3_1 _3887_ (.X(_0962_),
    .A(_2182_),
    .B(_0221_),
    .C(_2183_));
 sg13g2_nor3_1 _3888_ (.A(_0957_),
    .B(_0961_),
    .C(_0962_),
    .Y(_0963_));
 sg13g2_a21oi_1 _3889_ (.A1(_0952_),
    .A2(_0963_),
    .Y(_0964_),
    .B1(_1620_));
 sg13g2_nand3_1 _3890_ (.B(_0688_),
    .C(net107),
    .A(_0673_),
    .Y(_0965_));
 sg13g2_nand3_1 _3891_ (.B(_0656_),
    .C(net67),
    .A(_0641_),
    .Y(_0966_));
 sg13g2_nand3_1 _3892_ (.B(_0451_),
    .C(net68),
    .A(_0432_),
    .Y(_0967_));
 sg13g2_nand3_1 _3893_ (.B(_0624_),
    .C(net73),
    .A(_0609_),
    .Y(_0968_));
 sg13g2_nand3_1 _3894_ (.B(_0968_),
    .C(net121),
    .A(_0967_),
    .Y(_0969_));
 sg13g2_nand3_1 _3895_ (.B(_0640_),
    .C(net114),
    .A(_0625_),
    .Y(_0970_));
 sg13g2_nand3_1 _3896_ (.B(_0970_),
    .C(net47),
    .A(_0969_),
    .Y(_0971_));
 sg13g2_nand3_1 _3897_ (.B(_0971_),
    .C(net59),
    .A(_0966_),
    .Y(_0972_));
 sg13g2_nand3_1 _3898_ (.B(_0672_),
    .C(net66),
    .A(_0657_),
    .Y(_0973_));
 sg13g2_nand3_1 _3899_ (.B(_0973_),
    .C(net58),
    .A(_0972_),
    .Y(_0974_));
 sg13g2_nand3_1 _3900_ (.B(_0974_),
    .C(_0491_),
    .A(_0965_),
    .Y(_0975_));
 sg13g2_nand3_1 _3901_ (.B(_0704_),
    .C(net141),
    .A(_0689_),
    .Y(_0976_));
 sg13g2_nand3_1 _3902_ (.B(_0976_),
    .C(net95),
    .A(_0975_),
    .Y(_0977_));
 sg13g2_nand3_1 _3903_ (.B(_0720_),
    .C(net92),
    .A(_0705_),
    .Y(_0978_));
 sg13g2_nand3_1 _3904_ (.B(_0978_),
    .C(net50),
    .A(_0977_),
    .Y(_0979_));
 sg13g2_inv_2 _3905_ (.Y(_0980_),
    .A(_0885_));
 sg13g2_nand2_1 _3906_ (.Y(_0981_),
    .A(_0980_),
    .B(_1568_));
 sg13g2_a21oi_1 _3907_ (.A1(_0981_),
    .A2(net56),
    .Y(_0982_),
    .B1(_0745_));
 sg13g2_inv_1 _3908_ (.Y(_0983_),
    .A(_1568_));
 sg13g2_nand2_1 _3909_ (.Y(_0984_),
    .A(net172),
    .B(_1568_));
 sg13g2_nand2_1 _3910_ (.Y(_0985_),
    .A(net63),
    .B(_0984_));
 sg13g2_a22oi_1 _3911_ (.Y(_0986_),
    .B1(_0746_),
    .B2(_0985_),
    .A2(_0983_),
    .A1(_0745_));
 sg13g2_inv_1 _3912_ (.Y(_0987_),
    .A(\a[4] ));
 sg13g2_inv_1 _3913_ (.Y(_0988_),
    .A(_0198_));
 sg13g2_buf_1 _3914_ (.A(_0988_),
    .X(_0989_));
 sg13g2_a22oi_1 _3915_ (.Y(_0990_),
    .B1(\a[20] ),
    .B2(net38),
    .A2(_0339_),
    .A1(net41));
 sg13g2_o21ai_1 _3916_ (.B1(_0990_),
    .Y(_0991_),
    .A1(_0987_),
    .A2(net43));
 sg13g2_nor2_1 _3917_ (.A(_0037_),
    .B(_0812_),
    .Y(_0992_));
 sg13g2_nor2_1 _3918_ (.A(_2096_),
    .B(_0992_),
    .Y(_0993_));
 sg13g2_a21oi_1 _3919_ (.A1(_0814_),
    .A2(_2096_),
    .Y(_0994_),
    .B1(_0993_));
 sg13g2_nand2_1 _3920_ (.Y(_0995_),
    .A(_0994_),
    .B(net122));
 sg13g2_o21ai_1 _3921_ (.B1(_0995_),
    .Y(_0996_),
    .A1(net122),
    .A2(_0817_));
 sg13g2_nor2b_1 _3922_ (.A(net175),
    .B_N(_0996_),
    .Y(_0997_));
 sg13g2_a21o_1 _3923_ (.A2(net150),
    .A1(_0819_),
    .B1(_0997_),
    .X(_0998_));
 sg13g2_mux2_1 _3924_ (.A0(_0998_),
    .A1(_0821_),
    .S(net149),
    .X(_0999_));
 sg13g2_mux2_1 _3925_ (.A0(_0999_),
    .A1(_0835_),
    .S(net147),
    .X(_1000_));
 sg13g2_o21ai_1 _3926_ (.B1(net62),
    .Y(_1001_),
    .A1(net146),
    .A2(_1000_));
 sg13g2_nor2_1 _3927_ (.A(net93),
    .B(_0851_),
    .Y(_1002_));
 sg13g2_nor2_1 _3928_ (.A(_1001_),
    .B(_1002_),
    .Y(_1003_));
 sg13g2_nor4_1 _3929_ (.A(_0982_),
    .B(_0986_),
    .C(_0991_),
    .D(_1003_),
    .Y(_1004_));
 sg13g2_a21oi_1 _3930_ (.A1(_0979_),
    .A2(_1004_),
    .Y(_1005_),
    .B1(_1553_));
 sg13g2_nor2_1 _3931_ (.A(_0964_),
    .B(_1005_),
    .Y(_1006_));
 sg13g2_nand2_1 _3932_ (.Y(net14),
    .A(_0936_),
    .B(_1006_));
 sg13g2_nand3_1 _3933_ (.B(_0881_),
    .C(net105),
    .A(_0880_),
    .Y(_1007_));
 sg13g2_nand3_1 _3934_ (.B(_0879_),
    .C(net104),
    .A(_0870_),
    .Y(_1008_));
 sg13g2_nand3_1 _3935_ (.B(_0878_),
    .C(net107),
    .A(_0877_),
    .Y(_1009_));
 sg13g2_nand3_1 _3936_ (.B(net66),
    .C(_0876_),
    .A(_0871_),
    .Y(_1010_));
 sg13g2_nand3_1 _3937_ (.B(_0875_),
    .C(net67),
    .A(_0872_),
    .Y(_1011_));
 sg13g2_nand3_1 _3938_ (.B(_0730_),
    .C(_1775_),
    .A(_0727_),
    .Y(_1012_));
 sg13g2_nand3_1 _3939_ (.B(_0874_),
    .C(net114),
    .A(_0873_),
    .Y(_1013_));
 sg13g2_nand3_1 _3940_ (.B(_1013_),
    .C(_1770_),
    .A(_1012_),
    .Y(_1014_));
 sg13g2_nand3_1 _3941_ (.B(_1014_),
    .C(net123),
    .A(_1011_),
    .Y(_1015_));
 sg13g2_nand3_1 _3942_ (.B(_1015_),
    .C(net124),
    .A(_1010_),
    .Y(_1016_));
 sg13g2_nand3_1 _3943_ (.B(_1016_),
    .C(net103),
    .A(_1009_),
    .Y(_1017_));
 sg13g2_nand3_1 _3944_ (.B(_1017_),
    .C(net102),
    .A(_1008_),
    .Y(_1018_));
 sg13g2_nand3_1 _3945_ (.B(_1018_),
    .C(net50),
    .A(_1007_),
    .Y(_1019_));
 sg13g2_o21ai_1 _3946_ (.B1(net64),
    .Y(_1020_),
    .A1(net142),
    .A2(_0884_));
 sg13g2_o21ai_1 _3947_ (.B1(_1020_),
    .Y(_1021_),
    .A1(_0884_),
    .A2(_0885_));
 sg13g2_nor2_1 _3948_ (.A(_1773_),
    .B(_0856_),
    .Y(_1022_));
 sg13g2_a21oi_1 _3949_ (.A1(_1773_),
    .A2(_0888_),
    .Y(_1023_),
    .B1(_1022_));
 sg13g2_nor2b_1 _3950_ (.A(net122),
    .B_N(_0890_),
    .Y(_1024_));
 sg13g2_a21o_1 _3951_ (.A2(net122),
    .A1(_1023_),
    .B1(_1024_),
    .X(_1025_));
 sg13g2_nor2_1 _3952_ (.A(_1762_),
    .B(_1025_),
    .Y(_1026_));
 sg13g2_a21oi_1 _3953_ (.A1(_2214_),
    .A2(_0892_),
    .Y(_1027_),
    .B1(_1026_));
 sg13g2_mux2_1 _3954_ (.A0(_0894_),
    .A1(_1027_),
    .S(_1755_),
    .X(_1028_));
 sg13g2_nor2_1 _3955_ (.A(_1721_),
    .B(_1028_),
    .Y(_1029_));
 sg13g2_a21oi_1 _3956_ (.A1(net147),
    .A2(_0896_),
    .Y(_1030_),
    .B1(_1029_));
 sg13g2_mux2_1 _3957_ (.A0(_0898_),
    .A1(_1030_),
    .S(net93),
    .X(_1031_));
 sg13g2_inv_1 _3958_ (.Y(_1032_),
    .A(_1645_));
 sg13g2_a21oi_1 _3959_ (.A1(_1032_),
    .A2(net64),
    .Y(_1033_),
    .B1(_1369_));
 sg13g2_buf_1 _3960_ (.A(_1663_),
    .X(_1034_));
 sg13g2_nor2_1 _3961_ (.A(net103),
    .B(_0988_),
    .Y(_1035_));
 sg13g2_a221oi_1 _3962_ (.B2(_0215_),
    .C1(_1035_),
    .B1(_2179_),
    .A1(net39),
    .Y(_1036_),
    .A2(net70));
 sg13g2_o21ai_1 _3963_ (.B1(_1036_),
    .Y(_1037_),
    .A1(_0884_),
    .A2(_1033_));
 sg13g2_a221oi_1 _3964_ (.B2(net45),
    .C1(_1037_),
    .B1(_1031_),
    .A1(_1645_),
    .Y(_1038_),
    .A2(_1021_));
 sg13g2_a21oi_1 _3965_ (.A1(_1019_),
    .A2(_1038_),
    .Y(_1039_),
    .B1(_1423_));
 sg13g2_nand3_1 _3966_ (.B(_0921_),
    .C(net96),
    .A(_0910_),
    .Y(_1040_));
 sg13g2_nand3_1 _3967_ (.B(_0920_),
    .C(_0171_),
    .A(_0911_),
    .Y(_1041_));
 sg13g2_nand3_1 _3968_ (.B(_0919_),
    .C(_2220_),
    .A(_0912_),
    .Y(_1042_));
 sg13g2_nand3_1 _3969_ (.B(_0918_),
    .C(net71),
    .A(_0913_),
    .Y(_1043_));
 sg13g2_nand3_1 _3970_ (.B(_0917_),
    .C(_0159_),
    .A(_0914_),
    .Y(_1044_));
 sg13g2_nand3_1 _3971_ (.B(_0916_),
    .C(net72),
    .A(_0915_),
    .Y(_1045_));
 sg13g2_nand3_1 _3972_ (.B(_0157_),
    .C(net69),
    .A(_0155_),
    .Y(_1046_));
 sg13g2_nand3_1 _3973_ (.B(_1046_),
    .C(_0484_),
    .A(_1045_),
    .Y(_1047_));
 sg13g2_nand3_1 _3974_ (.B(_1047_),
    .C(_0486_),
    .A(_1044_),
    .Y(_1048_));
 sg13g2_nand3_1 _3975_ (.B(_1048_),
    .C(net58),
    .A(_1043_),
    .Y(_1049_));
 sg13g2_nand3_1 _3976_ (.B(_1049_),
    .C(_0174_),
    .A(_1042_),
    .Y(_1050_));
 sg13g2_nand3_1 _3977_ (.B(_1050_),
    .C(net95),
    .A(_1041_),
    .Y(_1051_));
 sg13g2_nand3_1 _3978_ (.B(_1051_),
    .C(_0511_),
    .A(_1040_),
    .Y(_1052_));
 sg13g2_a22oi_1 _3979_ (.Y(_1053_),
    .B1(_0339_),
    .B2(net65),
    .A2(_2009_),
    .A1(_1034_));
 sg13g2_o21ai_1 _3980_ (.B1(_1053_),
    .Y(_1054_),
    .A1(_1827_),
    .A2(_0738_));
 sg13g2_o21ai_1 _3981_ (.B1(\a[19] ),
    .Y(_1055_),
    .A1(_0924_),
    .A2(_1293_));
 sg13g2_a21oi_1 _3982_ (.A1(_0520_),
    .A2(_0924_),
    .Y(_1056_),
    .B1(_1055_));
 sg13g2_nand2_1 _3983_ (.Y(_1057_),
    .A(net63),
    .B(_1603_));
 sg13g2_a21oi_1 _3984_ (.A1(net40),
    .A2(_1057_),
    .Y(_1058_),
    .B1(_1601_));
 sg13g2_and3_1 _3985_ (.X(_1059_),
    .A(_0360_),
    .B(net48),
    .C(_0365_));
 sg13g2_nor4_1 _3986_ (.A(_1054_),
    .B(_1056_),
    .C(_1058_),
    .D(_1059_),
    .Y(_1060_));
 sg13g2_a21oi_1 _3987_ (.A1(_1052_),
    .A2(_1060_),
    .Y(_1061_),
    .B1(_1591_));
 sg13g2_nor2_1 _3988_ (.A(_1039_),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_nand3_1 _3989_ (.B(net147),
    .C(_0948_),
    .A(_0940_),
    .Y(_1063_));
 sg13g2_nand3_1 _3990_ (.B(net149),
    .C(_0947_),
    .A(_0941_),
    .Y(_1064_));
 sg13g2_nand3_1 _3991_ (.B(net109),
    .C(_0946_),
    .A(_0942_),
    .Y(_1065_));
 sg13g2_nand3_1 _3992_ (.B(net112),
    .C(_0945_),
    .A(_0943_),
    .Y(_1066_));
 sg13g2_inv_1 _3993_ (.Y(_1067_),
    .A(_0036_));
 sg13g2_nand2_1 _3994_ (.Y(_1068_),
    .A(_0944_),
    .B(_1067_));
 sg13g2_nand2_1 _3995_ (.Y(_1069_),
    .A(_1068_),
    .B(net83));
 sg13g2_nand3_1 _3996_ (.B(_1763_),
    .C(_1069_),
    .A(_1066_),
    .Y(_1070_));
 sg13g2_nand3_1 _3997_ (.B(net97),
    .C(_1070_),
    .A(_1065_),
    .Y(_1071_));
 sg13g2_nand3_1 _3998_ (.B(_1723_),
    .C(_1071_),
    .A(_1064_),
    .Y(_1072_));
 sg13g2_nand3_1 _3999_ (.B(net171),
    .C(_1072_),
    .A(_1063_),
    .Y(_1073_));
 sg13g2_nand2_1 _4000_ (.Y(_1074_),
    .A(_1073_),
    .B(_0194_));
 sg13g2_nand3_1 _4001_ (.B(_0604_),
    .C(_0949_),
    .A(_0939_),
    .Y(_1075_));
 sg13g2_nor2b_1 _4002_ (.A(_1074_),
    .B_N(_1075_),
    .Y(_1076_));
 sg13g2_a22oi_1 _4003_ (.Y(_1077_),
    .B1(net100),
    .B2(net65),
    .A2(net176),
    .A1(net39));
 sg13g2_o21ai_1 _4004_ (.B1(_1077_),
    .Y(_1078_),
    .A1(_1803_),
    .A2(_0738_));
 sg13g2_a21oi_1 _4005_ (.A1(net138),
    .A2(_0954_),
    .Y(_1079_),
    .B1(_1631_));
 sg13g2_o21ai_1 _4006_ (.B1(_1079_),
    .Y(_1080_),
    .A1(_0204_),
    .A2(_0954_));
 sg13g2_nor2_1 _4007_ (.A(\a[27] ),
    .B(net145),
    .Y(_1081_));
 sg13g2_o21ai_1 _4008_ (.B1(\a[26] ),
    .Y(_1082_),
    .A1(_1081_),
    .A2(_1369_));
 sg13g2_nand2_1 _4009_ (.Y(_1083_),
    .A(_1080_),
    .B(_1082_));
 sg13g2_and3_1 _4010_ (.X(_1084_),
    .A(_2072_),
    .B(net62),
    .C(_2073_));
 sg13g2_nor3_1 _4011_ (.A(_1078_),
    .B(_1083_),
    .C(_1084_),
    .Y(_1085_));
 sg13g2_nor2b_1 _4012_ (.A(_1076_),
    .B_N(_1085_),
    .Y(_1086_));
 sg13g2_nor2_1 _4013_ (.A(_1620_),
    .B(_1086_),
    .Y(_1087_));
 sg13g2_nand3_1 _4014_ (.B(_0452_),
    .C(net69),
    .A(_0431_),
    .Y(_1088_));
 sg13g2_nand3_1 _4015_ (.B(_0968_),
    .C(net77),
    .A(_0967_),
    .Y(_1089_));
 sg13g2_nand3_1 _4016_ (.B(_1089_),
    .C(_1770_),
    .A(_1088_),
    .Y(_1090_));
 sg13g2_nand3_1 _4017_ (.B(_0970_),
    .C(_2126_),
    .A(_0969_),
    .Y(_1091_));
 sg13g2_nand3_1 _4018_ (.B(_1091_),
    .C(net59),
    .A(_1090_),
    .Y(_1092_));
 sg13g2_nand3_1 _4019_ (.B(_0971_),
    .C(net66),
    .A(_0966_),
    .Y(_1093_));
 sg13g2_nand3_1 _4020_ (.B(_1093_),
    .C(net85),
    .A(_1092_),
    .Y(_1094_));
 sg13g2_nand3_1 _4021_ (.B(_0973_),
    .C(net107),
    .A(_0972_),
    .Y(_1095_));
 sg13g2_nand3_1 _4022_ (.B(_1095_),
    .C(net57),
    .A(_1094_),
    .Y(_1096_));
 sg13g2_nand3_1 _4023_ (.B(_0974_),
    .C(net106),
    .A(_0965_),
    .Y(_1097_));
 sg13g2_nand3_1 _4024_ (.B(_1097_),
    .C(net95),
    .A(_1096_),
    .Y(_1098_));
 sg13g2_nand3_1 _4025_ (.B(_0976_),
    .C(net92),
    .A(_0975_),
    .Y(_1099_));
 sg13g2_nand3_1 _4026_ (.B(_1099_),
    .C(net50),
    .A(_1098_),
    .Y(_1100_));
 sg13g2_inv_1 _4027_ (.Y(_1101_),
    .A(\a[11] ));
 sg13g2_a21oi_1 _4028_ (.A1(_0981_),
    .A2(_0985_),
    .Y(_1102_),
    .B1(_1101_));
 sg13g2_nand2_1 _4029_ (.Y(_1103_),
    .A(net63),
    .B(_1101_));
 sg13g2_a21oi_1 _4030_ (.A1(net40),
    .A2(_1103_),
    .Y(_1104_),
    .B1(_0983_));
 sg13g2_a22oi_1 _4031_ (.Y(_1105_),
    .B1(net164),
    .B2(_0216_),
    .A2(_0309_),
    .A1(_1034_));
 sg13g2_o21ai_1 _4032_ (.B1(_1105_),
    .Y(_1106_),
    .A1(_1776_),
    .A2(net43));
 sg13g2_nand2_1 _4033_ (.Y(_1107_),
    .A(_0992_),
    .B(_1067_));
 sg13g2_nor2_1 _4034_ (.A(net152),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_a21oi_1 _4035_ (.A1(_0994_),
    .A2(net152),
    .Y(_1109_),
    .B1(_1108_));
 sg13g2_nor2_1 _4036_ (.A(net168),
    .B(_0996_),
    .Y(_1110_));
 sg13g2_a21oi_1 _4037_ (.A1(net168),
    .A2(_1109_),
    .Y(_1111_),
    .B1(_1110_));
 sg13g2_inv_1 _4038_ (.Y(_1112_),
    .A(_1111_));
 sg13g2_nor2_1 _4039_ (.A(net149),
    .B(_1112_),
    .Y(_1113_));
 sg13g2_a21oi_1 _4040_ (.A1(_0998_),
    .A2(net149),
    .Y(_1114_),
    .B1(_1113_));
 sg13g2_nor2_1 _4041_ (.A(net170),
    .B(_0999_),
    .Y(_1115_));
 sg13g2_a21oi_1 _4042_ (.A1(net127),
    .A2(_1114_),
    .Y(_1116_),
    .B1(_1115_));
 sg13g2_nor2_1 _4043_ (.A(net146),
    .B(_1116_),
    .Y(_1117_));
 sg13g2_nor2_1 _4044_ (.A(net93),
    .B(_1000_),
    .Y(_1118_));
 sg13g2_nor3_1 _4045_ (.A(_0749_),
    .B(_1117_),
    .C(_1118_),
    .Y(_1119_));
 sg13g2_nor4_1 _4046_ (.A(_1102_),
    .B(_1104_),
    .C(_1106_),
    .D(_1119_),
    .Y(_1120_));
 sg13g2_a21oi_1 _4047_ (.A1(_1100_),
    .A2(_1120_),
    .Y(_1121_),
    .B1(_1553_));
 sg13g2_nor2_1 _4048_ (.A(_1087_),
    .B(_1121_),
    .Y(_1122_));
 sg13g2_nand2_1 _4049_ (.Y(net15),
    .A(_1062_),
    .B(_1122_));
 sg13g2_nand3_1 _4050_ (.B(_1017_),
    .C(net105),
    .A(_1008_),
    .Y(_1123_));
 sg13g2_nand3_1 _4051_ (.B(_1016_),
    .C(net104),
    .A(_1009_),
    .Y(_1124_));
 sg13g2_nand3_1 _4052_ (.B(_1015_),
    .C(net108),
    .A(_1010_),
    .Y(_1125_));
 sg13g2_nand3_1 _4053_ (.B(_0731_),
    .C(net47),
    .A(_0726_),
    .Y(_1126_));
 sg13g2_nand3_1 _4054_ (.B(_1013_),
    .C(net112),
    .A(_1012_),
    .Y(_1127_));
 sg13g2_nand3_1 _4055_ (.B(_1127_),
    .C(net123),
    .A(_1126_),
    .Y(_1128_));
 sg13g2_nand3_1 _4056_ (.B(_1014_),
    .C(_2215_),
    .A(_1011_),
    .Y(_1129_));
 sg13g2_nand3_1 _4057_ (.B(_1129_),
    .C(_1756_),
    .A(_1128_),
    .Y(_1130_));
 sg13g2_nand3_1 _4058_ (.B(_1130_),
    .C(net103),
    .A(_1125_),
    .Y(_1131_));
 sg13g2_nand3_1 _4059_ (.B(_1131_),
    .C(net102),
    .A(_1124_),
    .Y(_1132_));
 sg13g2_nand3_1 _4060_ (.B(_1132_),
    .C(net50),
    .A(_1123_),
    .Y(_1133_));
 sg13g2_nand2_1 _4061_ (.Y(_1134_),
    .A(_0980_),
    .B(\a[4] ));
 sg13g2_a21oi_1 _4062_ (.A1(_1134_),
    .A2(net56),
    .Y(_1135_),
    .B1(_1032_));
 sg13g2_nand2_1 _4063_ (.Y(_1136_),
    .A(net64),
    .B(_1032_));
 sg13g2_o21ai_1 _4064_ (.B1(net63),
    .Y(_1137_),
    .A1(net142),
    .A2(_0987_));
 sg13g2_a22oi_1 _4065_ (.Y(_1138_),
    .B1(_1136_),
    .B2(_1137_),
    .A2(_1032_),
    .A1(_0987_));
 sg13g2_a22oi_1 _4066_ (.Y(_1139_),
    .B1(_1597_),
    .B2(net38),
    .A2(net71),
    .A1(net39));
 sg13g2_o21ai_1 _4067_ (.B1(_1139_),
    .Y(_1140_),
    .A1(_0901_),
    .A2(net43));
 sg13g2_o21ai_1 _4068_ (.B1(net62),
    .Y(_1141_),
    .A1(net171),
    .A2(_1030_));
 sg13g2_nor2b_1 _4069_ (.A(_1768_),
    .B_N(_1023_),
    .Y(_1142_));
 sg13g2_a21o_1 _4070_ (.A2(_0858_),
    .A1(net122),
    .B1(_1142_),
    .X(_1143_));
 sg13g2_inv_1 _4071_ (.Y(_1144_),
    .A(_1143_));
 sg13g2_nor2_1 _4072_ (.A(net168),
    .B(_1025_),
    .Y(_1145_));
 sg13g2_a21oi_1 _4073_ (.A1(_1144_),
    .A2(net168),
    .Y(_1146_),
    .B1(_1145_));
 sg13g2_nor2b_1 _4074_ (.A(net97),
    .B_N(_1027_),
    .Y(_1147_));
 sg13g2_a21o_1 _4075_ (.A2(net97),
    .A1(_1146_),
    .B1(_1147_),
    .X(_1148_));
 sg13g2_mux2_1 _4076_ (.A0(_1028_),
    .A1(_1148_),
    .S(net170),
    .X(_1149_));
 sg13g2_nor2_1 _4077_ (.A(net140),
    .B(_1149_),
    .Y(_1150_));
 sg13g2_nor2_1 _4078_ (.A(_1141_),
    .B(_1150_),
    .Y(_1151_));
 sg13g2_nor4_1 _4079_ (.A(_1135_),
    .B(_1138_),
    .C(_1140_),
    .D(_1151_),
    .Y(_1152_));
 sg13g2_a21oi_1 _4080_ (.A1(_1133_),
    .A2(_1152_),
    .Y(_1153_),
    .B1(_1423_));
 sg13g2_nand3_1 _4081_ (.B(_1050_),
    .C(net96),
    .A(_1041_),
    .Y(_1154_));
 sg13g2_nand3_1 _4082_ (.B(_1048_),
    .C(net107),
    .A(_1043_),
    .Y(_1155_));
 sg13g2_nand3_1 _4083_ (.B(_1046_),
    .C(_0159_),
    .A(_1045_),
    .Y(_1156_));
 sg13g2_nand3_1 _4084_ (.B(_0158_),
    .C(net47),
    .A(_2248_),
    .Y(_1157_));
 sg13g2_nand3_1 _4085_ (.B(_1157_),
    .C(net59),
    .A(_1156_),
    .Y(_1158_));
 sg13g2_nand3_1 _4086_ (.B(_1047_),
    .C(_0161_),
    .A(_1044_),
    .Y(_1159_));
 sg13g2_nand3_1 _4087_ (.B(_1159_),
    .C(net58),
    .A(_1158_),
    .Y(_1160_));
 sg13g2_nand3_1 _4088_ (.B(_1160_),
    .C(net86),
    .A(_1155_),
    .Y(_1161_));
 sg13g2_nand3_1 _4089_ (.B(_1049_),
    .C(net106),
    .A(_1042_),
    .Y(_1162_));
 sg13g2_nand3_1 _4090_ (.B(_1162_),
    .C(_0509_),
    .A(_1161_),
    .Y(_1163_));
 sg13g2_nand3_1 _4091_ (.B(_1163_),
    .C(_0511_),
    .A(_1154_),
    .Y(_1164_));
 sg13g2_nand2_1 _4092_ (.Y(_1165_),
    .A(_0980_),
    .B(\a[20] ));
 sg13g2_a21oi_1 _4093_ (.A1(_1165_),
    .A2(_1380_),
    .Y(_1166_),
    .B1(_1603_));
 sg13g2_o21ai_1 _4094_ (.B1(_0208_),
    .Y(_1167_),
    .A1(_0516_),
    .A2(_1608_));
 sg13g2_a22oi_1 _4095_ (.Y(_1168_),
    .B1(_1057_),
    .B2(_1167_),
    .A2(_1603_),
    .A1(_1608_));
 sg13g2_a22oi_1 _4096_ (.Y(_1169_),
    .B1(_1626_),
    .B2(net38),
    .A2(net158),
    .A1(net41));
 sg13g2_o21ai_1 _4097_ (.B1(_1169_),
    .Y(_1170_),
    .A1(_0745_),
    .A2(net43));
 sg13g2_and3_1 _4098_ (.X(_1171_),
    .A(_0325_),
    .B(net48),
    .C(_0332_));
 sg13g2_nor4_1 _4099_ (.A(_1166_),
    .B(_1168_),
    .C(_1170_),
    .D(_1171_),
    .Y(_1172_));
 sg13g2_a21oi_1 _4100_ (.A1(_1164_),
    .A2(_1172_),
    .Y(_1173_),
    .B1(_1591_));
 sg13g2_nor2_1 _4101_ (.A(_1153_),
    .B(_1173_),
    .Y(_1174_));
 sg13g2_nand3_1 _4102_ (.B(_1093_),
    .C(_2219_),
    .A(_1092_),
    .Y(_1175_));
 sg13g2_nand3_1 _4103_ (.B(_0453_),
    .C(_0484_),
    .A(_0430_),
    .Y(_1176_));
 sg13g2_nand3_1 _4104_ (.B(_1089_),
    .C(net67),
    .A(_1088_),
    .Y(_1177_));
 sg13g2_nand3_1 _4105_ (.B(_1177_),
    .C(_1764_),
    .A(_1176_),
    .Y(_1178_));
 sg13g2_nand3_1 _4106_ (.B(_1091_),
    .C(_2215_),
    .A(_1090_),
    .Y(_1179_));
 sg13g2_nand3_1 _4107_ (.B(_1179_),
    .C(_1756_),
    .A(_1178_),
    .Y(_1180_));
 sg13g2_nand3_1 _4108_ (.B(_1180_),
    .C(net57),
    .A(_1175_),
    .Y(_1181_));
 sg13g2_nand3_1 _4109_ (.B(_1095_),
    .C(net106),
    .A(_1094_),
    .Y(_1182_));
 sg13g2_nand3_1 _4110_ (.B(_1182_),
    .C(net139),
    .A(_1181_),
    .Y(_1183_));
 sg13g2_nand3_1 _4111_ (.B(_1097_),
    .C(net105),
    .A(_1096_),
    .Y(_1184_));
 sg13g2_nand3_1 _4112_ (.B(_1184_),
    .C(net50),
    .A(_1183_),
    .Y(_1185_));
 sg13g2_nand2_1 _4113_ (.Y(_1186_),
    .A(_0980_),
    .B(\a[11] ));
 sg13g2_inv_1 _4114_ (.Y(_1187_),
    .A(\a[12] ));
 sg13g2_a21oi_1 _4115_ (.A1(_1186_),
    .A2(_1103_),
    .Y(_1188_),
    .B1(_1187_));
 sg13g2_o21ai_1 _4116_ (.B1(net64),
    .Y(_1189_),
    .A1(net142),
    .A2(_1187_));
 sg13g2_a21oi_1 _4117_ (.A1(_1189_),
    .A2(net40),
    .Y(_1190_),
    .B1(_1101_));
 sg13g2_inv_1 _4118_ (.Y(_1191_),
    .A(\a[5] ));
 sg13g2_a22oi_1 _4119_ (.Y(_1192_),
    .B1(_1610_),
    .B2(net38),
    .A2(_0307_),
    .A1(net41));
 sg13g2_o21ai_1 _4120_ (.B1(_1192_),
    .Y(_1193_),
    .A1(_1191_),
    .A2(net43));
 sg13g2_nor2_1 _4121_ (.A(_0035_),
    .B(_1107_),
    .Y(_1194_));
 sg13g2_nor2_1 _4122_ (.A(net175),
    .B(_1194_),
    .Y(_1195_));
 sg13g2_a21oi_1 _4123_ (.A1(_1109_),
    .A2(net150),
    .Y(_1196_),
    .B1(_1195_));
 sg13g2_nand2_1 _4124_ (.Y(_1197_),
    .A(_1196_),
    .B(_1755_));
 sg13g2_o21ai_1 _4125_ (.B1(_1197_),
    .Y(_1198_),
    .A1(net97),
    .A2(_1112_));
 sg13g2_nand2_1 _4126_ (.Y(_1199_),
    .A(_1198_),
    .B(_1722_));
 sg13g2_o21ai_1 _4127_ (.B1(_1199_),
    .Y(_1200_),
    .A1(net127),
    .A2(_1114_));
 sg13g2_nor2_1 _4128_ (.A(net146),
    .B(_1200_),
    .Y(_1201_));
 sg13g2_nor2_1 _4129_ (.A(net93),
    .B(_1116_),
    .Y(_1202_));
 sg13g2_nor3_1 _4130_ (.A(_0749_),
    .B(_1201_),
    .C(_1202_),
    .Y(_1203_));
 sg13g2_nor4_1 _4131_ (.A(_1188_),
    .B(_1190_),
    .C(_1193_),
    .D(_1203_),
    .Y(_1204_));
 sg13g2_nand2_1 _4132_ (.Y(_1205_),
    .A(_1185_),
    .B(_1204_));
 sg13g2_nand3_1 _4133_ (.B(net105),
    .C(_1072_),
    .A(_1063_),
    .Y(_1206_));
 sg13g2_nand3_1 _4134_ (.B(net141),
    .C(_1071_),
    .A(_1064_),
    .Y(_1207_));
 sg13g2_nand3_1 _4135_ (.B(net108),
    .C(_1070_),
    .A(_1065_),
    .Y(_1208_));
 sg13g2_nand3_1 _4136_ (.B(net109),
    .C(_1069_),
    .A(_1066_),
    .Y(_1209_));
 sg13g2_nor2_1 _4137_ (.A(_0035_),
    .B(_1068_),
    .Y(_1210_));
 sg13g2_nand2_1 _4138_ (.Y(_1211_),
    .A(_1210_),
    .B(net123));
 sg13g2_nand3_1 _4139_ (.B(net124),
    .C(_1211_),
    .A(_1209_),
    .Y(_1212_));
 sg13g2_nand3_1 _4140_ (.B(net103),
    .C(_1212_),
    .A(_1208_),
    .Y(_1213_));
 sg13g2_nand3_1 _4141_ (.B(_0596_),
    .C(_1213_),
    .A(_1207_),
    .Y(_1214_));
 sg13g2_nand3_1 _4142_ (.B(net44),
    .C(_1214_),
    .A(_1206_),
    .Y(_1215_));
 sg13g2_a21oi_1 _4143_ (.A1(_0980_),
    .A2(\a[27] ),
    .Y(_1216_),
    .B1(_1081_));
 sg13g2_nor2_1 _4144_ (.A(_1633_),
    .B(_1216_),
    .Y(_1217_));
 sg13g2_o21ai_1 _4145_ (.B1(net64),
    .Y(_1218_),
    .A1(net142),
    .A2(_1633_));
 sg13g2_a21oi_1 _4146_ (.A1(_1218_),
    .A2(_1380_),
    .Y(_1219_),
    .B1(_1631_));
 sg13g2_inv_1 _4147_ (.Y(_1220_),
    .A(_1578_));
 sg13g2_a22oi_1 _4148_ (.Y(_1221_),
    .B1(\a[29] ),
    .B2(_0215_),
    .A2(_1748_),
    .A1(net39));
 sg13g2_o21ai_1 _4149_ (.B1(_1221_),
    .Y(_1222_),
    .A1(_1220_),
    .A2(net43));
 sg13g2_and3_1 _4150_ (.X(_1223_),
    .A(_2014_),
    .B(net48),
    .C(_2015_));
 sg13g2_nor4_1 _4151_ (.A(_1217_),
    .B(_1219_),
    .C(_1222_),
    .D(_1223_),
    .Y(_1224_));
 sg13g2_a21oi_1 _4152_ (.A1(_1215_),
    .A2(_1224_),
    .Y(_1225_),
    .B1(_1620_));
 sg13g2_a21oi_1 _4153_ (.A1(_1205_),
    .A2(_1542_),
    .Y(_1226_),
    .B1(_1225_));
 sg13g2_nand2_1 _4154_ (.Y(net16),
    .A(_1174_),
    .B(_1226_));
 sg13g2_nand3_1 _4155_ (.B(_1129_),
    .C(net108),
    .A(_1128_),
    .Y(_1227_));
 sg13g2_nand3_1 _4156_ (.B(_0732_),
    .C(net123),
    .A(_0725_),
    .Y(_1228_));
 sg13g2_nand3_1 _4157_ (.B(_1127_),
    .C(net109),
    .A(_1126_),
    .Y(_1229_));
 sg13g2_nand3_1 _4158_ (.B(_1229_),
    .C(net124),
    .A(_1228_),
    .Y(_1230_));
 sg13g2_nand3_1 _4159_ (.B(_1230_),
    .C(net86),
    .A(_1227_),
    .Y(_1231_));
 sg13g2_nand3_1 _4160_ (.B(_1130_),
    .C(net106),
    .A(_1125_),
    .Y(_1232_));
 sg13g2_nand3_1 _4161_ (.B(_1232_),
    .C(net95),
    .A(_1231_),
    .Y(_1233_));
 sg13g2_nand3_1 _4162_ (.B(_1131_),
    .C(net92),
    .A(_1124_),
    .Y(_1234_));
 sg13g2_nand3_1 _4163_ (.B(_1234_),
    .C(_0951_),
    .A(_1233_),
    .Y(_1235_));
 sg13g2_a21oi_1 _4164_ (.A1(_1134_),
    .A2(_1137_),
    .Y(_1236_),
    .B1(_1191_));
 sg13g2_nand2_1 _4165_ (.Y(_1237_),
    .A(net63),
    .B(_1191_));
 sg13g2_a21oi_1 _4166_ (.A1(net40),
    .A2(_1237_),
    .Y(_1238_),
    .B1(_0987_));
 sg13g2_a22oi_1 _4167_ (.Y(_1239_),
    .B1(net70),
    .B2(net65),
    .A2(net76),
    .A1(net39));
 sg13g2_o21ai_1 _4168_ (.B1(_1239_),
    .Y(_1240_),
    .A1(_1715_),
    .A2(_0738_));
 sg13g2_nor2_1 _4169_ (.A(net175),
    .B(_0860_),
    .Y(_1241_));
 sg13g2_a21oi_1 _4170_ (.A1(net150),
    .A2(_1144_),
    .Y(_1242_),
    .B1(_1241_));
 sg13g2_nor2b_1 _4171_ (.A(_1755_),
    .B_N(_1146_),
    .Y(_1243_));
 sg13g2_a21o_1 _4172_ (.A2(_1242_),
    .A1(net97),
    .B1(_1243_),
    .X(_1244_));
 sg13g2_mux2_1 _4173_ (.A0(_1148_),
    .A1(_1244_),
    .S(net170),
    .X(_1245_));
 sg13g2_nor2_1 _4174_ (.A(net140),
    .B(_1245_),
    .Y(_1246_));
 sg13g2_o21ai_1 _4175_ (.B1(net62),
    .Y(_1247_),
    .A1(net171),
    .A2(_1149_));
 sg13g2_nor2_1 _4176_ (.A(_1246_),
    .B(_1247_),
    .Y(_1248_));
 sg13g2_nor4_1 _4177_ (.A(_1236_),
    .B(_1238_),
    .C(_1240_),
    .D(_1248_),
    .Y(_1249_));
 sg13g2_a21oi_1 _4178_ (.A1(_1235_),
    .A2(_1249_),
    .Y(_1250_),
    .B1(_1423_));
 sg13g2_nand3_1 _4179_ (.B(_1162_),
    .C(net96),
    .A(_1161_),
    .Y(_1251_));
 sg13g2_nand3_1 _4180_ (.B(_1159_),
    .C(net107),
    .A(_1158_),
    .Y(_1252_));
 sg13g2_nand3_1 _4181_ (.B(_0160_),
    .C(net59),
    .A(_2246_),
    .Y(_1253_));
 sg13g2_nand3_1 _4182_ (.B(_1157_),
    .C(_0161_),
    .A(_1156_),
    .Y(_1254_));
 sg13g2_nand3_1 _4183_ (.B(_1254_),
    .C(_0489_),
    .A(_1253_),
    .Y(_1255_));
 sg13g2_nand3_1 _4184_ (.B(_1255_),
    .C(_1724_),
    .A(_1252_),
    .Y(_1256_));
 sg13g2_nand3_1 _4185_ (.B(_1160_),
    .C(_0166_),
    .A(_1155_),
    .Y(_1257_));
 sg13g2_nand3_1 _4186_ (.B(_1257_),
    .C(_0509_),
    .A(_1256_),
    .Y(_1258_));
 sg13g2_nand3_1 _4187_ (.B(_1258_),
    .C(net46),
    .A(_1251_),
    .Y(_1259_));
 sg13g2_a21oi_1 _4188_ (.A1(_1165_),
    .A2(_1167_),
    .Y(_1261_),
    .B1(_1611_));
 sg13g2_nand2_1 _4189_ (.Y(_1262_),
    .A(net64),
    .B(_1611_));
 sg13g2_a21oi_1 _4190_ (.A1(_0744_),
    .A2(_1262_),
    .Y(_1263_),
    .B1(_1608_));
 sg13g2_a22oi_1 _4191_ (.Y(_1264_),
    .B1(net176),
    .B2(_0216_),
    .A2(net163),
    .A1(net41));
 sg13g2_o21ai_1 _4192_ (.B1(_1264_),
    .Y(_1265_),
    .A1(net54),
    .A2(_0989_));
 sg13g2_and3_1 _4193_ (.X(_1266_),
    .A(_0293_),
    .B(net48),
    .C(_0302_));
 sg13g2_nor4_1 _4194_ (.A(_1261_),
    .B(_1263_),
    .C(_1265_),
    .D(_1266_),
    .Y(_1267_));
 sg13g2_a21oi_1 _4195_ (.A1(_1259_),
    .A2(_1267_),
    .Y(_1268_),
    .B1(_1591_));
 sg13g2_nor2_1 _4196_ (.A(_1250_),
    .B(_1268_),
    .Y(_1269_));
 sg13g2_nand3_1 _4197_ (.B(_0454_),
    .C(_1765_),
    .A(_0429_),
    .Y(_1270_));
 sg13g2_nand3_1 _4198_ (.B(_1177_),
    .C(net71),
    .A(_1176_),
    .Y(_1272_));
 sg13g2_nand3_1 _4199_ (.B(_1272_),
    .C(_1757_),
    .A(_1270_),
    .Y(_1273_));
 sg13g2_nand3_1 _4200_ (.B(_1179_),
    .C(_0163_),
    .A(_1178_),
    .Y(_1274_));
 sg13g2_nand3_1 _4201_ (.B(_1274_),
    .C(net103),
    .A(_1273_),
    .Y(_1275_));
 sg13g2_nand3_1 _4202_ (.B(_1180_),
    .C(net141),
    .A(_1175_),
    .Y(_1276_));
 sg13g2_nand3_1 _4203_ (.B(_1276_),
    .C(net139),
    .A(_1275_),
    .Y(_1277_));
 sg13g2_nand3_1 _4204_ (.B(_1182_),
    .C(net92),
    .A(_1181_),
    .Y(_1278_));
 sg13g2_nand3_1 _4205_ (.B(_1278_),
    .C(_0195_),
    .A(_1277_),
    .Y(_1279_));
 sg13g2_nand2_1 _4206_ (.Y(_1280_),
    .A(_0980_),
    .B(_1578_));
 sg13g2_a21oi_1 _4207_ (.A1(_1280_),
    .A2(net40),
    .Y(_1281_),
    .B1(_1187_));
 sg13g2_a22oi_1 _4208_ (.Y(_1283_),
    .B1(net60),
    .B2(net49),
    .A2(net101),
    .A1(net41));
 sg13g2_nand2_1 _4209_ (.Y(_1284_),
    .A(_0209_),
    .B(_1578_));
 sg13g2_a21oi_1 _4210_ (.A1(_1187_),
    .A2(_1220_),
    .Y(_1285_),
    .B1(net145));
 sg13g2_o21ai_1 _4211_ (.B1(_1285_),
    .Y(_1286_),
    .A1(_1187_),
    .A2(_1284_));
 sg13g2_nand2_1 _4212_ (.Y(_1287_),
    .A(net37),
    .B(net166));
 sg13g2_nand3_1 _4213_ (.B(_1286_),
    .C(_1287_),
    .A(_1283_),
    .Y(_1288_));
 sg13g2_inv_1 _4214_ (.Y(_1289_),
    .A(_0034_));
 sg13g2_nand2_1 _4215_ (.Y(_1290_),
    .A(_1194_),
    .B(_1289_));
 sg13g2_nor2_1 _4216_ (.A(_2218_),
    .B(_1290_),
    .Y(_1291_));
 sg13g2_a21oi_1 _4217_ (.A1(_1196_),
    .A2(net149),
    .Y(_1292_),
    .B1(_1291_));
 sg13g2_nand2_1 _4218_ (.Y(_1294_),
    .A(_1198_),
    .B(net147));
 sg13g2_o21ai_1 _4219_ (.B1(_1294_),
    .Y(_1295_),
    .A1(net147),
    .A2(_1292_));
 sg13g2_nor2_1 _4220_ (.A(net140),
    .B(_1295_),
    .Y(_1296_));
 sg13g2_nor2_1 _4221_ (.A(net93),
    .B(_1200_),
    .Y(_1297_));
 sg13g2_nor3_1 _4222_ (.A(_0749_),
    .B(_1296_),
    .C(_1297_),
    .Y(_1298_));
 sg13g2_nor3_1 _4223_ (.A(_1281_),
    .B(_1288_),
    .C(_1298_),
    .Y(_1299_));
 sg13g2_nand2_1 _4224_ (.Y(_1300_),
    .A(_1279_),
    .B(_1299_));
 sg13g2_nand2_1 _4225_ (.Y(_1301_),
    .A(_1210_),
    .B(_1289_));
 sg13g2_a21o_1 _4226_ (.A2(_1211_),
    .A1(_1209_),
    .B1(net124),
    .X(_1302_));
 sg13g2_o21ai_1 _4227_ (.B1(_1302_),
    .Y(_1303_),
    .A1(net107),
    .A2(_1301_));
 sg13g2_nand2_1 _4228_ (.Y(_1305_),
    .A(_1303_),
    .B(net86));
 sg13g2_nand3_1 _4229_ (.B(net141),
    .C(_1212_),
    .A(_1208_),
    .Y(_1306_));
 sg13g2_nand3_1 _4230_ (.B(net95),
    .C(_1306_),
    .A(_1305_),
    .Y(_1307_));
 sg13g2_nand3_1 _4231_ (.B(net92),
    .C(_1213_),
    .A(_1207_),
    .Y(_1308_));
 sg13g2_nand3_1 _4232_ (.B(net44),
    .C(_1308_),
    .A(_1307_),
    .Y(_1309_));
 sg13g2_nand3_1 _4233_ (.B(_1940_),
    .C(_0220_),
    .A(_1939_),
    .Y(_1310_));
 sg13g2_nor3_1 _4234_ (.A(net142),
    .B(_1633_),
    .C(_1635_),
    .Y(_1311_));
 sg13g2_inv_1 _4235_ (.Y(_1312_),
    .A(_1311_));
 sg13g2_a21oi_1 _4236_ (.A1(_1633_),
    .A2(_1635_),
    .Y(_1313_),
    .B1(net94));
 sg13g2_a22oi_1 _4237_ (.Y(_1314_),
    .B1(_1312_),
    .B2(_1313_),
    .A2(net143),
    .A1(_0200_));
 sg13g2_a22oi_1 _4238_ (.Y(_1316_),
    .B1(_1759_),
    .B2(_0514_),
    .A2(_1750_),
    .A1(_1664_));
 sg13g2_a22oi_1 _4239_ (.Y(_1317_),
    .B1(\a[28] ),
    .B2(net55),
    .A2(net188),
    .A1(_1311_));
 sg13g2_and4_1 _4240_ (.A(_1310_),
    .B(_1314_),
    .C(_1316_),
    .D(_1317_),
    .X(_1318_));
 sg13g2_a21oi_1 _4241_ (.A1(_1309_),
    .A2(_1318_),
    .Y(_1319_),
    .B1(_1620_));
 sg13g2_a21oi_1 _4242_ (.A1(_1300_),
    .A2(_1542_),
    .Y(_1320_),
    .B1(_1319_));
 sg13g2_nand2_1 _4243_ (.Y(net17),
    .A(_1269_),
    .B(_1320_));
 sg13g2_nand3_1 _4244_ (.B(_1232_),
    .C(net105),
    .A(_1231_),
    .Y(_1321_));
 sg13g2_nand3_1 _4245_ (.B(_0733_),
    .C(net58),
    .A(_0724_),
    .Y(_1322_));
 sg13g2_nand3_1 _4246_ (.B(_1229_),
    .C(_2219_),
    .A(_1228_),
    .Y(_1323_));
 sg13g2_nand3_1 _4247_ (.B(_1323_),
    .C(net57),
    .A(_1322_),
    .Y(_1324_));
 sg13g2_nand3_1 _4248_ (.B(_1230_),
    .C(_0574_),
    .A(_1227_),
    .Y(_1326_));
 sg13g2_nand3_1 _4249_ (.B(_1326_),
    .C(net102),
    .A(_1324_),
    .Y(_1327_));
 sg13g2_nand3_1 _4250_ (.B(_1327_),
    .C(net44),
    .A(_1321_),
    .Y(_1328_));
 sg13g2_nand2_1 _4251_ (.Y(_1329_),
    .A(_0980_),
    .B(\a[6] ));
 sg13g2_a21oi_1 _4252_ (.A1(_1329_),
    .A2(net56),
    .Y(_1330_),
    .B1(_1191_));
 sg13g2_inv_1 _4253_ (.Y(_1331_),
    .A(\a[6] ));
 sg13g2_o21ai_1 _4254_ (.B1(net63),
    .Y(_1332_),
    .A1(net142),
    .A2(_1331_));
 sg13g2_a22oi_1 _4255_ (.Y(_1333_),
    .B1(_1237_),
    .B2(_1332_),
    .A2(_1331_),
    .A1(_1191_));
 sg13g2_inv_1 _4256_ (.Y(_1334_),
    .A(net41));
 sg13g2_a22oi_1 _4257_ (.Y(_1335_),
    .B1(\a[18] ),
    .B2(net38),
    .A2(_1637_),
    .A1(net65));
 sg13g2_o21ai_1 _4258_ (.B1(_1335_),
    .Y(_1337_),
    .A1(net82),
    .A2(_1334_));
 sg13g2_mux2_1 _4259_ (.A0(_1242_),
    .A1(_0861_),
    .S(_1755_),
    .X(_1338_));
 sg13g2_inv_1 _4260_ (.Y(_1339_),
    .A(_1338_));
 sg13g2_nor2_1 _4261_ (.A(net170),
    .B(_1244_),
    .Y(_1340_));
 sg13g2_a21oi_1 _4262_ (.A1(_1339_),
    .A2(net127),
    .Y(_1341_),
    .B1(_1340_));
 sg13g2_nor2_1 _4263_ (.A(net146),
    .B(_1341_),
    .Y(_1342_));
 sg13g2_nor2_1 _4264_ (.A(net93),
    .B(_1245_),
    .Y(_1343_));
 sg13g2_nor3_1 _4265_ (.A(_0749_),
    .B(_1342_),
    .C(_1343_),
    .Y(_1344_));
 sg13g2_nor4_1 _4266_ (.A(_1330_),
    .B(_1333_),
    .C(_1337_),
    .D(_1344_),
    .Y(_1345_));
 sg13g2_a21oi_1 _4267_ (.A1(_1328_),
    .A2(_1345_),
    .Y(_1346_),
    .B1(_1423_));
 sg13g2_nand3_1 _4268_ (.B(_1257_),
    .C(_0493_),
    .A(_1256_),
    .Y(_1348_));
 sg13g2_nand3_1 _4269_ (.B(_1254_),
    .C(_0163_),
    .A(_1253_),
    .Y(_1349_));
 sg13g2_nand3_1 _4270_ (.B(_0162_),
    .C(net58),
    .A(_2245_),
    .Y(_1350_));
 sg13g2_nand3_1 _4271_ (.B(_1350_),
    .C(net57),
    .A(_1349_),
    .Y(_1351_));
 sg13g2_nand3_1 _4272_ (.B(_1255_),
    .C(_0166_),
    .A(_1252_),
    .Y(_1352_));
 sg13g2_nand3_1 _4273_ (.B(_1352_),
    .C(_0187_),
    .A(_1351_),
    .Y(_1353_));
 sg13g2_nand3_1 _4274_ (.B(_1353_),
    .C(net46),
    .A(_1348_),
    .Y(_1354_));
 sg13g2_nand2_1 _4275_ (.Y(_1355_),
    .A(_1315_),
    .B(\a[22] ));
 sg13g2_inv_1 _4276_ (.Y(_1356_),
    .A(_1355_));
 sg13g2_nand2_1 _4277_ (.Y(_1357_),
    .A(_1356_),
    .B(_1610_));
 sg13g2_nand2_1 _4278_ (.Y(_1359_),
    .A(_1661_),
    .B(net164));
 sg13g2_a21oi_1 _4279_ (.A1(_1357_),
    .A2(_1359_),
    .Y(_1360_),
    .B1(_1658_));
 sg13g2_a21oi_1 _4280_ (.A1(_1611_),
    .A2(_1613_),
    .Y(_1361_),
    .B1(_0203_));
 sg13g2_a22oi_1 _4281_ (.Y(_1362_),
    .B1(\a[26] ),
    .B2(_0514_),
    .A2(_1357_),
    .A1(_1361_));
 sg13g2_a22oi_1 _4282_ (.Y(_1363_),
    .B1(_1568_),
    .B2(net49),
    .A2(_1610_),
    .A1(_1564_));
 sg13g2_nand2_1 _4283_ (.Y(_1364_),
    .A(_1362_),
    .B(_1363_));
 sg13g2_and3_1 _4284_ (.X(_1365_),
    .A(_0266_),
    .B(net45),
    .C(_0277_));
 sg13g2_nor3_1 _4285_ (.A(_1360_),
    .B(_1364_),
    .C(_1365_),
    .Y(_1366_));
 sg13g2_a21oi_1 _4286_ (.A1(_1354_),
    .A2(_1366_),
    .Y(_1367_),
    .B1(_1591_));
 sg13g2_nor2_1 _4287_ (.A(_1346_),
    .B(_1367_),
    .Y(_1368_));
 sg13g2_nor2_1 _4288_ (.A(_0033_),
    .B(_1290_),
    .Y(_1370_));
 sg13g2_nand2_1 _4289_ (.Y(_1371_),
    .A(_1370_),
    .B(net127));
 sg13g2_o21ai_1 _4290_ (.B1(_1371_),
    .Y(_1372_),
    .A1(net127),
    .A2(_1292_));
 sg13g2_o21ai_1 _4291_ (.B1(net45),
    .Y(_1373_),
    .A1(_0604_),
    .A2(_1372_));
 sg13g2_nor2_1 _4292_ (.A(_0596_),
    .B(_1295_),
    .Y(_1374_));
 sg13g2_o21ai_1 _4293_ (.B1(net56),
    .Y(_1375_),
    .A1(_1582_),
    .A2(net94));
 sg13g2_inv_1 _4294_ (.Y(_1376_),
    .A(_1284_));
 sg13g2_o21ai_1 _4295_ (.B1(_1280_),
    .Y(_1377_),
    .A1(net94),
    .A2(_1376_));
 sg13g2_a22oi_1 _4296_ (.Y(_1378_),
    .B1(\a[22] ),
    .B2(_0215_),
    .A2(net100),
    .A1(net39));
 sg13g2_o21ai_1 _4297_ (.B1(_1378_),
    .Y(_1379_),
    .A1(_1331_),
    .A2(net43));
 sg13g2_a221oi_1 _4298_ (.B2(_1377_),
    .C1(_1379_),
    .B1(_1582_),
    .A1(_1578_),
    .Y(_1381_),
    .A2(_1375_));
 sg13g2_o21ai_1 _4299_ (.B1(_1381_),
    .Y(_1382_),
    .A1(_1373_),
    .A2(_1374_));
 sg13g2_nand3_1 _4300_ (.B(_0455_),
    .C(_1757_),
    .A(_0428_),
    .Y(_1383_));
 sg13g2_nand3_1 _4301_ (.B(_1272_),
    .C(_2220_),
    .A(_1270_),
    .Y(_1384_));
 sg13g2_nand3_1 _4302_ (.B(_1384_),
    .C(_0491_),
    .A(_1383_),
    .Y(_1385_));
 sg13g2_nand3_1 _4303_ (.B(_1274_),
    .C(net106),
    .A(_1273_),
    .Y(_1386_));
 sg13g2_nand3_1 _4304_ (.B(_1386_),
    .C(net95),
    .A(_1385_),
    .Y(_1387_));
 sg13g2_nand3_1 _4305_ (.B(_1276_),
    .C(_0937_),
    .A(_1275_),
    .Y(_1388_));
 sg13g2_nand3_1 _4306_ (.B(_1388_),
    .C(net44),
    .A(_1387_),
    .Y(_1389_));
 sg13g2_nand2b_1 _4307_ (.Y(_1390_),
    .B(_1389_),
    .A_N(_1382_));
 sg13g2_nand3_1 _4308_ (.B(net105),
    .C(_1306_),
    .A(_1305_),
    .Y(_1392_));
 sg13g2_nand2_1 _4309_ (.Y(_1393_),
    .A(_1303_),
    .B(net104));
 sg13g2_nor2_1 _4310_ (.A(_0033_),
    .B(_1301_),
    .Y(_1394_));
 sg13g2_nand2_1 _4311_ (.Y(_1395_),
    .A(_1394_),
    .B(net86));
 sg13g2_nand3_1 _4312_ (.B(net102),
    .C(_1395_),
    .A(_1393_),
    .Y(_1396_));
 sg13g2_nand3_1 _4313_ (.B(_1396_),
    .C(net44),
    .A(_1392_),
    .Y(_1397_));
 sg13g2_nor3_1 _4314_ (.A(net142),
    .B(_1635_),
    .C(_1640_),
    .Y(_1398_));
 sg13g2_inv_1 _4315_ (.Y(_1399_),
    .A(_1398_));
 sg13g2_nand2_1 _4316_ (.Y(_1400_),
    .A(_1661_),
    .B(_1752_));
 sg13g2_a21oi_1 _4317_ (.A1(_1399_),
    .A2(_1400_),
    .Y(_1401_),
    .B1(net138));
 sg13g2_a22oi_1 _4318_ (.Y(_1403_),
    .B1(_1639_),
    .B2(_0215_),
    .A2(_1582_),
    .A1(_0199_));
 sg13g2_o21ai_1 _4319_ (.B1(_1403_),
    .Y(_1404_),
    .A1(_1635_),
    .A2(net56));
 sg13g2_nor2_1 _4320_ (.A(\a[29] ),
    .B(_1639_),
    .Y(_1405_));
 sg13g2_nor3_1 _4321_ (.A(net94),
    .B(_1405_),
    .C(_1398_),
    .Y(_1406_));
 sg13g2_and3_1 _4322_ (.X(_1407_),
    .A(_1879_),
    .B(net48),
    .C(_1883_));
 sg13g2_nor4_1 _4323_ (.A(_1401_),
    .B(_1404_),
    .C(_1406_),
    .D(_1407_),
    .Y(_1408_));
 sg13g2_a21oi_1 _4324_ (.A1(_1397_),
    .A2(_1408_),
    .Y(_1409_),
    .B1(_1620_));
 sg13g2_a21oi_1 _4325_ (.A1(_1390_),
    .A2(_1542_),
    .Y(_1410_),
    .B1(_1409_));
 sg13g2_nand2_1 _4326_ (.Y(net18),
    .A(_1368_),
    .B(_1410_));
 sg13g2_nand3_1 _4327_ (.B(_1326_),
    .C(_0169_),
    .A(_1324_),
    .Y(_1411_));
 sg13g2_nand3_1 _4328_ (.B(_0734_),
    .C(net103),
    .A(_0723_),
    .Y(_1413_));
 sg13g2_nand3_1 _4329_ (.B(_1323_),
    .C(_0574_),
    .A(_1322_),
    .Y(_1414_));
 sg13g2_nand3_1 _4330_ (.B(_1414_),
    .C(net102),
    .A(_1413_),
    .Y(_1415_));
 sg13g2_nand3_1 _4331_ (.B(_1415_),
    .C(_0951_),
    .A(_1411_),
    .Y(_1416_));
 sg13g2_inv_1 _4332_ (.Y(_1417_),
    .A(_1650_));
 sg13g2_a21oi_1 _4333_ (.A1(_1329_),
    .A2(_1332_),
    .Y(_1418_),
    .B1(_1417_));
 sg13g2_nand2_1 _4334_ (.Y(_1419_),
    .A(net64),
    .B(_1417_));
 sg13g2_a21oi_1 _4335_ (.A1(net40),
    .A2(_1419_),
    .Y(_1420_),
    .B1(_1331_));
 sg13g2_a22oi_1 _4336_ (.Y(_1421_),
    .B1(net158),
    .B2(net38),
    .A2(net60),
    .A1(net39));
 sg13g2_o21ai_1 _4337_ (.B1(_1421_),
    .Y(_1422_),
    .A1(net84),
    .A2(net43));
 sg13g2_o21ai_1 _4338_ (.B1(net62),
    .Y(_1424_),
    .A1(net171),
    .A2(_1341_));
 sg13g2_nor2_1 _4339_ (.A(_1721_),
    .B(_0862_),
    .Y(_1425_));
 sg13g2_a21oi_1 _4340_ (.A1(_1339_),
    .A2(net147),
    .Y(_1426_),
    .B1(_1425_));
 sg13g2_nor2_1 _4341_ (.A(net140),
    .B(_1426_),
    .Y(_1427_));
 sg13g2_nor2_1 _4342_ (.A(_1424_),
    .B(_1427_),
    .Y(_1428_));
 sg13g2_nor4_1 _4343_ (.A(_1418_),
    .B(_1420_),
    .C(_1422_),
    .D(_1428_),
    .Y(_1429_));
 sg13g2_a21oi_1 _4344_ (.A1(_1416_),
    .A2(_1429_),
    .Y(_1430_),
    .B1(_1423_));
 sg13g2_nand3_1 _4345_ (.B(_1352_),
    .C(_0169_),
    .A(_1351_),
    .Y(_1431_));
 sg13g2_nand3_1 _4346_ (.B(_0164_),
    .C(net57),
    .A(_2244_),
    .Y(_1432_));
 sg13g2_nand3_1 _4347_ (.B(_1350_),
    .C(net106),
    .A(_1349_),
    .Y(_1433_));
 sg13g2_nand3_1 _4348_ (.B(_1433_),
    .C(net102),
    .A(_1432_),
    .Y(_1435_));
 sg13g2_nand3_1 _4349_ (.B(_1435_),
    .C(net46),
    .A(_1431_),
    .Y(_1436_));
 sg13g2_a22oi_1 _4350_ (.Y(_1437_),
    .B1(_0307_),
    .B2(net49),
    .A2(net166),
    .A1(net41));
 sg13g2_o21ai_1 _4351_ (.B1(_1437_),
    .Y(_1438_),
    .A1(_1815_),
    .A2(_0738_));
 sg13g2_a21oi_1 _4352_ (.A1(_1615_),
    .A2(_0205_),
    .Y(_1439_),
    .B1(_1369_));
 sg13g2_a21oi_1 _4353_ (.A1(_1658_),
    .A2(_1356_),
    .Y(_1440_),
    .B1(_1615_));
 sg13g2_o21ai_1 _4354_ (.B1(_1440_),
    .Y(_1441_),
    .A1(_0205_),
    .A2(_1356_));
 sg13g2_o21ai_1 _4355_ (.B1(_1441_),
    .Y(_1442_),
    .A1(_1613_),
    .A2(_1439_));
 sg13g2_and3_1 _4356_ (.X(_1443_),
    .A(_0242_),
    .B(net48),
    .C(_0255_));
 sg13g2_nor3_1 _4357_ (.A(_1438_),
    .B(_1442_),
    .C(_1443_),
    .Y(_1444_));
 sg13g2_a21oi_1 _4358_ (.A1(_1436_),
    .A2(_1444_),
    .Y(_1446_),
    .B1(_1591_));
 sg13g2_nor2_1 _4359_ (.A(_1430_),
    .B(_1446_),
    .Y(_1447_));
 sg13g2_nand3_1 _4360_ (.B(_0471_),
    .C(_1724_),
    .A(_0456_),
    .Y(_1448_));
 sg13g2_nand3_1 _4361_ (.B(_1384_),
    .C(net104),
    .A(_1383_),
    .Y(_1449_));
 sg13g2_nand3_1 _4362_ (.B(_1449_),
    .C(net139),
    .A(_1448_),
    .Y(_1450_));
 sg13g2_nand3_1 _4363_ (.B(_1386_),
    .C(net92),
    .A(_1385_),
    .Y(_1451_));
 sg13g2_nand3_1 _4364_ (.B(_1451_),
    .C(_0195_),
    .A(_1450_),
    .Y(_1452_));
 sg13g2_inv_1 _4365_ (.Y(_1453_),
    .A(net186));
 sg13g2_inv_1 _4366_ (.Y(_1454_),
    .A(_1582_));
 sg13g2_nor3_1 _4367_ (.A(net142),
    .B(_1453_),
    .C(_1454_),
    .Y(_1455_));
 sg13g2_inv_1 _4368_ (.Y(_1457_),
    .A(_1455_));
 sg13g2_a21oi_1 _4369_ (.A1(_1453_),
    .A2(_1454_),
    .Y(_1458_),
    .B1(net94));
 sg13g2_nand2b_1 _4370_ (.Y(_1459_),
    .B(_0937_),
    .A_N(_1372_));
 sg13g2_nor3_1 _4371_ (.A(_0033_),
    .B(_0032_),
    .C(_1290_),
    .Y(_1460_));
 sg13g2_nor2_1 _4372_ (.A(net146),
    .B(_1460_),
    .Y(_1461_));
 sg13g2_nor2_1 _4373_ (.A(_0749_),
    .B(_1461_),
    .Y(_1462_));
 sg13g2_a21oi_1 _4374_ (.A1(net143),
    .A2(_1661_),
    .Y(_1463_),
    .B1(_1455_));
 sg13g2_nor2_1 _4375_ (.A(net80),
    .B(_0988_),
    .Y(_1464_));
 sg13g2_a221oi_1 _4376_ (.B2(net173),
    .C1(_1464_),
    .B1(_0215_),
    .A1(_1369_),
    .Y(_1465_),
    .A2(_1582_));
 sg13g2_o21ai_1 _4377_ (.B1(_1465_),
    .Y(_1466_),
    .A1(net138),
    .A2(_1463_));
 sg13g2_a221oi_1 _4378_ (.B2(_1462_),
    .C1(_1466_),
    .B1(_1459_),
    .A1(_1457_),
    .Y(_1468_),
    .A2(_1458_));
 sg13g2_nand2_1 _4379_ (.Y(_1469_),
    .A(_1452_),
    .B(_1468_));
 sg13g2_nand3_1 _4380_ (.B(net105),
    .C(_1395_),
    .A(_1393_),
    .Y(_1470_));
 sg13g2_nor3_1 _4381_ (.A(_0033_),
    .B(_0032_),
    .C(_1301_),
    .Y(_1471_));
 sg13g2_nand2b_1 _4382_ (.Y(_1472_),
    .B(net139),
    .A_N(_1471_));
 sg13g2_nand3_1 _4383_ (.B(net44),
    .C(_1472_),
    .A(_1470_),
    .Y(_1473_));
 sg13g2_nand3_1 _4384_ (.B(net48),
    .C(_1888_),
    .A(_1885_),
    .Y(_1474_));
 sg13g2_a22oi_1 _4385_ (.Y(_1475_),
    .B1(net144),
    .B2(net49),
    .A2(_1759_),
    .A1(net42));
 sg13g2_a22oi_1 _4386_ (.Y(_1476_),
    .B1(\ayayayayayaya.b[31] ),
    .B2(net37),
    .A2(_1639_),
    .A1(net55));
 sg13g2_nand3_1 _4387_ (.B(_1642_),
    .C(_1639_),
    .A(net172),
    .Y(_1477_));
 sg13g2_nor2_1 _4388_ (.A(net138),
    .B(_1477_),
    .Y(_1479_));
 sg13g2_nand2_1 _4389_ (.Y(_1480_),
    .A(_1643_),
    .B(_1640_));
 sg13g2_nand3_1 _4390_ (.B(net63),
    .C(_1480_),
    .A(_1477_),
    .Y(_1481_));
 sg13g2_nor2b_1 _4391_ (.A(_1479_),
    .B_N(_1481_),
    .Y(_1482_));
 sg13g2_and4_1 _4392_ (.A(_1474_),
    .B(_1475_),
    .C(_1476_),
    .D(_1482_),
    .X(_1483_));
 sg13g2_a21oi_1 _4393_ (.A1(_1473_),
    .A2(_1483_),
    .Y(_1484_),
    .B1(_1620_));
 sg13g2_a21oi_1 _4394_ (.A1(_1469_),
    .A2(_1542_),
    .Y(_1485_),
    .B1(_1484_));
 sg13g2_nand2_1 _4395_ (.Y(net19),
    .A(_1447_),
    .B(_1485_));
 sg13g2_nand3_1 _4396_ (.B(_0492_),
    .C(_1657_),
    .A(_0472_),
    .Y(_1486_));
 sg13g2_nand3_1 _4397_ (.B(_1449_),
    .C(net96),
    .A(_1448_),
    .Y(_1487_));
 sg13g2_nand3_1 _4398_ (.B(_1487_),
    .C(net46),
    .A(_1486_),
    .Y(_1489_));
 sg13g2_inv_1 _4399_ (.Y(_1490_),
    .A(_0031_));
 sg13g2_nand3_1 _4400_ (.B(_1490_),
    .C(net45),
    .A(_1460_),
    .Y(_1491_));
 sg13g2_nand2_1 _4401_ (.Y(_1492_),
    .A(net186),
    .B(net187));
 sg13g2_nand3_1 _4402_ (.B(net172),
    .C(_1659_),
    .A(net188),
    .Y(_1493_));
 sg13g2_nor2_1 _4403_ (.A(_1492_),
    .B(_1493_),
    .Y(_1494_));
 sg13g2_nand2_1 _4404_ (.Y(_1495_),
    .A(net186),
    .B(_1588_));
 sg13g2_nand3_1 _4405_ (.B(net172),
    .C(_1325_),
    .A(net188),
    .Y(_1496_));
 sg13g2_nor2_1 _4406_ (.A(_1495_),
    .B(_1496_),
    .Y(_1497_));
 sg13g2_o21ai_1 _4407_ (.B1(_1402_),
    .Y(_1498_),
    .A1(_1615_),
    .A2(_0738_));
 sg13g2_inv_1 _4408_ (.Y(_1499_),
    .A(_1495_));
 sg13g2_nand3_1 _4409_ (.B(net189),
    .C(_1325_),
    .A(_0204_),
    .Y(_1500_));
 sg13g2_nand2_1 _4410_ (.Y(_1501_),
    .A(_0204_),
    .B(_1661_));
 sg13g2_o21ai_1 _4411_ (.B1(_1501_),
    .Y(_1502_),
    .A1(_1499_),
    .A2(_1500_));
 sg13g2_o21ai_1 _4412_ (.B1(_1502_),
    .Y(_1503_),
    .A1(net186),
    .A2(_1588_));
 sg13g2_inv_1 _4413_ (.Y(_1504_),
    .A(_1492_));
 sg13g2_nand3_1 _4414_ (.B(net189),
    .C(_1659_),
    .A(_0204_),
    .Y(_1505_));
 sg13g2_nand2_1 _4415_ (.Y(_1506_),
    .A(_0204_),
    .B(_1336_));
 sg13g2_o21ai_1 _4416_ (.B1(_1506_),
    .Y(_1507_),
    .A1(_1504_),
    .A2(_1505_));
 sg13g2_o21ai_1 _4417_ (.B1(_1507_),
    .Y(_1508_),
    .A1(net186),
    .A2(net187));
 sg13g2_nand2_1 _4418_ (.Y(_1510_),
    .A(net55),
    .B(net186));
 sg13g2_a22oi_1 _4419_ (.Y(_1511_),
    .B1(_1650_),
    .B2(net65),
    .A2(net144),
    .A1(net39));
 sg13g2_nand4_1 _4420_ (.B(_1508_),
    .C(_1510_),
    .A(_1503_),
    .Y(_1512_),
    .D(_1511_));
 sg13g2_nor4_1 _4421_ (.A(_1494_),
    .B(_1497_),
    .C(_1498_),
    .D(_1512_),
    .Y(_1513_));
 sg13g2_nand3_1 _4422_ (.B(_1491_),
    .C(_1513_),
    .A(_1489_),
    .Y(_1514_));
 sg13g2_nand3_1 _4423_ (.B(_0735_),
    .C(net139),
    .A(_0722_),
    .Y(_1515_));
 sg13g2_nand3_1 _4424_ (.B(_1414_),
    .C(net92),
    .A(_1413_),
    .Y(_1516_));
 sg13g2_nand3_1 _4425_ (.B(_1516_),
    .C(net50),
    .A(_1515_),
    .Y(_1517_));
 sg13g2_nor2_1 _4426_ (.A(net171),
    .B(_1426_),
    .Y(_1518_));
 sg13g2_nor2_1 _4427_ (.A(net140),
    .B(_0863_),
    .Y(_1519_));
 sg13g2_nor2_1 _4428_ (.A(_1518_),
    .B(_1519_),
    .Y(_1521_));
 sg13g2_a22oi_1 _4429_ (.Y(_1522_),
    .B1(\a[19] ),
    .B2(net38),
    .A2(_1645_),
    .A1(net65));
 sg13g2_nand2_1 _4430_ (.Y(_1523_),
    .A(_1347_),
    .B(_0741_));
 sg13g2_nand3_1 _4431_ (.B(_1650_),
    .C(net188),
    .A(_1523_),
    .Y(_1524_));
 sg13g2_a21oi_1 _4432_ (.A1(_0747_),
    .A2(_1417_),
    .Y(_1525_),
    .B1(net145));
 sg13g2_o21ai_1 _4433_ (.B1(_1525_),
    .Y(_1526_),
    .A1(_1417_),
    .A2(_0741_));
 sg13g2_nand4_1 _4434_ (.B(_1524_),
    .C(_1531_),
    .A(_1522_),
    .Y(_1527_),
    .D(_1526_));
 sg13g2_a221oi_1 _4435_ (.B2(net45),
    .C1(_1527_),
    .B1(_1521_),
    .A1(_2205_),
    .Y(_1528_),
    .A2(net42));
 sg13g2_a21oi_1 _4436_ (.A1(_1517_),
    .A2(_1528_),
    .Y(_1529_),
    .B1(_1391_));
 sg13g2_nand2_1 _4437_ (.Y(_1530_),
    .A(_1514_),
    .B(_1529_));
 sg13g2_nand3_1 _4438_ (.B(_1490_),
    .C(net44),
    .A(_1471_),
    .Y(_1532_));
 sg13g2_nand2_1 _4439_ (.Y(_1533_),
    .A(_1892_),
    .B(_0598_));
 sg13g2_nand2_1 _4440_ (.Y(_1534_),
    .A(_1642_),
    .B(_1588_));
 sg13g2_nor2_1 _4441_ (.A(_1534_),
    .B(_1493_),
    .Y(_1535_));
 sg13g2_nand2_1 _4442_ (.Y(_1536_),
    .A(_1642_),
    .B(net187));
 sg13g2_nor2_1 _4443_ (.A(_1536_),
    .B(_1496_),
    .Y(_1537_));
 sg13g2_a21oi_1 _4444_ (.A1(_0738_),
    .A2(net56),
    .Y(_1538_),
    .B1(_1643_));
 sg13g2_a221oi_1 _4445_ (.B2(_0198_),
    .C1(_1531_),
    .B1(net186),
    .A1(_1663_),
    .Y(_1539_),
    .A2(\ayayayayayaya.b[31] ));
 sg13g2_inv_1 _4446_ (.Y(_1540_),
    .A(_1534_));
 sg13g2_o21ai_1 _4447_ (.B1(_1506_),
    .Y(_1541_),
    .A1(_1540_),
    .A2(_1505_));
 sg13g2_o21ai_1 _4448_ (.B1(_1541_),
    .Y(_1543_),
    .A1(_1642_),
    .A2(_1588_));
 sg13g2_inv_1 _4449_ (.Y(_1544_),
    .A(_1536_));
 sg13g2_o21ai_1 _4450_ (.B1(_1501_),
    .Y(_1545_),
    .A1(_1544_),
    .A2(_1500_));
 sg13g2_o21ai_1 _4451_ (.B1(_1545_),
    .Y(_1546_),
    .A1(_1642_),
    .A2(net187));
 sg13g2_nand3_1 _4452_ (.B(_1543_),
    .C(_1546_),
    .A(_1539_),
    .Y(_1547_));
 sg13g2_nor4_1 _4453_ (.A(_1535_),
    .B(_1537_),
    .C(_1538_),
    .D(_1547_),
    .Y(_1548_));
 sg13g2_nand3_1 _4454_ (.B(_1533_),
    .C(_1548_),
    .A(_1532_),
    .Y(_1549_));
 sg13g2_nand2_1 _4455_ (.Y(_1550_),
    .A(_1549_),
    .B(_1391_));
 sg13g2_nand3_1 _4456_ (.B(_1433_),
    .C(net96),
    .A(_1432_),
    .Y(_1551_));
 sg13g2_nand3_1 _4457_ (.B(_0167_),
    .C(_1657_),
    .A(_2243_),
    .Y(_1552_));
 sg13g2_nand3_1 _4458_ (.B(_1552_),
    .C(net46),
    .A(_1551_),
    .Y(_1554_));
 sg13g2_nand3_1 _4459_ (.B(_0240_),
    .C(_0598_),
    .A(_0239_),
    .Y(_1555_));
 sg13g2_a21oi_1 _4460_ (.A1(_0212_),
    .A2(net40),
    .Y(_1556_),
    .B1(_1615_));
 sg13g2_nor3_1 _4461_ (.A(_1618_),
    .B(\a[23] ),
    .C(_0520_),
    .Y(_1557_));
 sg13g2_a22oi_1 _4462_ (.Y(_1558_),
    .B1(\a[27] ),
    .B2(net37),
    .A2(net173),
    .A1(_0213_));
 sg13g2_o21ai_1 _4463_ (.B1(_1558_),
    .Y(_1559_),
    .A1(_1101_),
    .A2(_0989_));
 sg13g2_nor4_1 _4464_ (.A(_1402_),
    .B(_1556_),
    .C(_1557_),
    .D(_1559_),
    .Y(_1560_));
 sg13g2_nand3_1 _4465_ (.B(_1555_),
    .C(_1560_),
    .A(_1554_),
    .Y(_1561_));
 sg13g2_nand2b_1 _4466_ (.Y(_1562_),
    .B(_1561_),
    .A_N(_1550_));
 sg13g2_nand2_1 _4467_ (.Y(net20),
    .A(_1530_),
    .B(_1562_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _4469_ (.A(net12),
    .X(net5));
 sg13g2_buf_1 _4470_ (.A(net12),
    .X(net6));
 sg13g2_buf_1 _4471_ (.A(net12),
    .X(net7));
 sg13g2_buf_1 _4472_ (.A(net12),
    .X(net8));
 sg13g2_buf_1 _4473_ (.A(net12),
    .X(net9));
 sg13g2_buf_1 _4474_ (.A(net12),
    .X(net10));
 sg13g2_buf_1 _4475_ (.A(net12),
    .X(net11));
 sg13g2_buf_1 _4476_ (.A(net13),
    .X(net21));
 sg13g2_buf_1 _4477_ (.A(net14),
    .X(net22));
 sg13g2_buf_1 _4478_ (.A(net15),
    .X(net23));
 sg13g2_buf_1 _4479_ (.A(net16),
    .X(net24));
 sg13g2_buf_1 _4480_ (.A(net17),
    .X(net25));
 sg13g2_buf_1 _4481_ (.A(net18),
    .X(net26));
 sg13g2_buf_1 _4482_ (.A(net19),
    .X(net27));
 sg13g2_buf_1 _4483_ (.A(net20),
    .X(net28));
 sg13g2_dfrbp_1 \a[0]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net190),
    .D(_0060_),
    .Q_N(_0000_),
    .Q(\a[0] ));
 sg13g2_dfrbp_1 \a[10]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net191),
    .D(_0061_),
    .Q_N(_0010_),
    .Q(\a[10] ));
 sg13g2_dfrbp_1 \a[11]$_DFFE_PP_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net192),
    .D(_0062_),
    .Q_N(_0011_),
    .Q(\a[11] ));
 sg13g2_dfrbp_1 \a[12]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net193),
    .D(_0063_),
    .Q_N(_0012_),
    .Q(\a[12] ));
 sg13g2_dfrbp_1 \a[13]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net194),
    .D(_0064_),
    .Q_N(_0013_),
    .Q(\a[13] ));
 sg13g2_dfrbp_1 \a[14]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net195),
    .D(_0065_),
    .Q_N(_0014_),
    .Q(\a[14] ));
 sg13g2_dfrbp_1 \a[15]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net196),
    .D(_0066_),
    .Q_N(_0015_),
    .Q(\a[15] ));
 sg13g2_dfrbp_1 \a[16]$_DFFE_PP_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net197),
    .D(_0067_),
    .Q_N(_0016_),
    .Q(\a[16] ));
 sg13g2_dfrbp_1 \a[17]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net198),
    .D(_0068_),
    .Q_N(_0017_),
    .Q(\a[17] ));
 sg13g2_dfrbp_1 \a[18]$_DFFE_PP_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net199),
    .D(_0069_),
    .Q_N(_0018_),
    .Q(\a[18] ));
 sg13g2_dfrbp_1 \a[19]$_DFFE_PP_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net200),
    .D(_0070_),
    .Q_N(_0019_),
    .Q(\a[19] ));
 sg13g2_dfrbp_1 \a[1]$_DFFE_PP_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net201),
    .D(_0071_),
    .Q_N(_0001_),
    .Q(\a[1] ));
 sg13g2_dfrbp_1 \a[20]$_DFFE_PP_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net202),
    .D(_0072_),
    .Q_N(_0020_),
    .Q(\a[20] ));
 sg13g2_dfrbp_1 \a[21]$_DFFE_PP_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net203),
    .D(_0073_),
    .Q_N(_0021_),
    .Q(\a[21] ));
 sg13g2_dfrbp_1 \a[22]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net204),
    .D(_0074_),
    .Q_N(_0022_),
    .Q(\a[22] ));
 sg13g2_dfrbp_1 \a[23]$_DFFE_PP_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net205),
    .D(_0075_),
    .Q_N(_0023_),
    .Q(\a[23] ));
 sg13g2_dfrbp_1 \a[24]$_DFFE_PP_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net206),
    .D(_0076_),
    .Q_N(_0024_),
    .Q(\a[24] ));
 sg13g2_dfrbp_1 \a[25]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net207),
    .D(_0077_),
    .Q_N(_0025_),
    .Q(\a[25] ));
 sg13g2_dfrbp_1 \a[26]$_DFFE_PP_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net208),
    .D(_0078_),
    .Q_N(_0026_),
    .Q(\a[26] ));
 sg13g2_dfrbp_1 \a[27]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net209),
    .D(_0079_),
    .Q_N(_0027_),
    .Q(\a[27] ));
 sg13g2_dfrbp_1 \a[28]$_DFFE_PP_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net210),
    .D(_0080_),
    .Q_N(_0028_),
    .Q(\a[28] ));
 sg13g2_dfrbp_1 \a[29]$_DFFE_PP_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net211),
    .D(_0081_),
    .Q_N(_0029_),
    .Q(\a[29] ));
 sg13g2_dfrbp_1 \a[2]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net212),
    .D(_0082_),
    .Q_N(_0002_),
    .Q(\a[2] ));
 sg13g2_dfrbp_1 \a[30]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net213),
    .D(_0083_),
    .Q_N(_0030_),
    .Q(\a[30] ));
 sg13g2_dfrbp_1 \a[31]$_DFFE_PP_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net214),
    .D(_0084_),
    .Q_N(_2260_),
    .Q(\a[31] ));
 sg13g2_dfrbp_1 \a[3]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net215),
    .D(_0085_),
    .Q_N(_0003_),
    .Q(\a[3] ));
 sg13g2_dfrbp_1 \a[4]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net216),
    .D(_0086_),
    .Q_N(_0004_),
    .Q(\a[4] ));
 sg13g2_dfrbp_1 \a[5]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net217),
    .D(_0087_),
    .Q_N(_0005_),
    .Q(\a[5] ));
 sg13g2_dfrbp_1 \a[6]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net218),
    .D(_0088_),
    .Q_N(_0006_),
    .Q(\a[6] ));
 sg13g2_dfrbp_1 \a[7]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net219),
    .D(_0089_),
    .Q_N(_0007_),
    .Q(\a[7] ));
 sg13g2_dfrbp_1 \a[8]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net220),
    .D(_0090_),
    .Q_N(_0008_),
    .Q(\a[8] ));
 sg13g2_dfrbp_1 \a[9]$_DFFE_PP_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net221),
    .D(_0091_),
    .Q_N(_0009_),
    .Q(\a[9] ));
 sg13g2_dfrbp_1 \b[0]$_DFFE_PP_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net222),
    .D(_0092_),
    .Q_N(_0031_),
    .Q(\ayayayayayaya.b[0] ));
 sg13g2_dfrbp_1 \b[10]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net223),
    .D(_0093_),
    .Q_N(_0041_),
    .Q(\ayayayayayaya.b[10] ));
 sg13g2_dfrbp_1 \b[11]$_DFFE_PP_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net224),
    .D(_0094_),
    .Q_N(_0042_),
    .Q(\ayayayayayaya.b[11] ));
 sg13g2_dfrbp_1 \b[12]$_DFFE_PP_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net225),
    .D(_0095_),
    .Q_N(_0043_),
    .Q(\ayayayayayaya.b[12] ));
 sg13g2_dfrbp_1 \b[13]$_DFFE_PP_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net226),
    .D(_0096_),
    .Q_N(_0044_),
    .Q(\ayayayayayaya.b[13] ));
 sg13g2_dfrbp_1 \b[14]$_DFFE_PP_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net227),
    .D(_0097_),
    .Q_N(_0045_),
    .Q(\ayayayayayaya.b[14] ));
 sg13g2_dfrbp_1 \b[15]$_DFFE_PP_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net228),
    .D(_0098_),
    .Q_N(_0046_),
    .Q(\ayayayayayaya.b[15] ));
 sg13g2_dfrbp_1 \b[16]$_DFFE_PP_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net229),
    .D(_0099_),
    .Q_N(_0047_),
    .Q(\ayayayayayaya.b[16] ));
 sg13g2_dfrbp_1 \b[17]$_DFFE_PP_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net230),
    .D(_0100_),
    .Q_N(_0048_),
    .Q(\ayayayayayaya.b[17] ));
 sg13g2_dfrbp_1 \b[18]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net231),
    .D(_0101_),
    .Q_N(_0049_),
    .Q(\ayayayayayaya.b[18] ));
 sg13g2_dfrbp_1 \b[19]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net232),
    .D(_0102_),
    .Q_N(_0050_),
    .Q(\ayayayayayaya.b[19] ));
 sg13g2_dfrbp_1 \b[1]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net233),
    .D(_0103_),
    .Q_N(_0032_),
    .Q(\ayayayayayaya.b[1] ));
 sg13g2_dfrbp_1 \b[20]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net234),
    .D(_0104_),
    .Q_N(_0051_),
    .Q(\ayayayayayaya.b[20] ));
 sg13g2_dfrbp_1 \b[21]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net235),
    .D(_0105_),
    .Q_N(_0052_),
    .Q(\ayayayayayaya.b[21] ));
 sg13g2_dfrbp_1 \b[22]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net236),
    .D(_0106_),
    .Q_N(_0053_),
    .Q(\ayayayayayaya.b[22] ));
 sg13g2_dfrbp_1 \b[23]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net237),
    .D(_0107_),
    .Q_N(_0054_),
    .Q(\ayayayayayaya.b[23] ));
 sg13g2_dfrbp_1 \b[24]$_DFFE_PP_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net238),
    .D(_0108_),
    .Q_N(_0055_),
    .Q(\ayayayayayaya.b[24] ));
 sg13g2_dfrbp_1 \b[25]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net239),
    .D(_0109_),
    .Q_N(_0056_),
    .Q(\ayayayayayaya.b[25] ));
 sg13g2_dfrbp_1 \b[26]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net240),
    .D(_0110_),
    .Q_N(_0057_),
    .Q(\ayayayayayaya.b[26] ));
 sg13g2_dfrbp_1 \b[27]$_DFFE_PP_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net241),
    .D(_0111_),
    .Q_N(_0058_),
    .Q(\ayayayayayaya.b[27] ));
 sg13g2_dfrbp_1 \b[28]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net242),
    .D(_0112_),
    .Q_N(_0059_),
    .Q(\ayayayayayaya.b[28] ));
 sg13g2_dfrbp_1 \b[29]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net243),
    .D(_0113_),
    .Q_N(_2259_),
    .Q(\ayayayayayaya.b[29] ));
 sg13g2_dfrbp_1 \b[2]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net244),
    .D(_0114_),
    .Q_N(_0033_),
    .Q(\ayayayayayaya.b[2] ));
 sg13g2_dfrbp_1 \b[30]$_DFFE_PP_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net245),
    .D(_0115_),
    .Q_N(_2258_),
    .Q(\ayayayayayaya.b[30] ));
 sg13g2_dfrbp_1 \b[31]$_DFFE_PP_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net246),
    .D(_0116_),
    .Q_N(_2257_),
    .Q(\ayayayayayaya.b[31] ));
 sg13g2_dfrbp_1 \b[3]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net247),
    .D(_0117_),
    .Q_N(_0034_),
    .Q(\ayayayayayaya.b[3] ));
 sg13g2_dfrbp_1 \b[4]$_DFFE_PP_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net248),
    .D(_0118_),
    .Q_N(_0035_),
    .Q(\ayayayayayaya.b[4] ));
 sg13g2_dfrbp_1 \b[5]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net249),
    .D(_0119_),
    .Q_N(_0036_),
    .Q(\ayayayayayaya.b[5] ));
 sg13g2_dfrbp_1 \b[6]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net250),
    .D(_0120_),
    .Q_N(_0037_),
    .Q(\ayayayayayaya.b[6] ));
 sg13g2_dfrbp_1 \b[7]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net251),
    .D(_0121_),
    .Q_N(_0038_),
    .Q(\ayayayayayaya.b[7] ));
 sg13g2_dfrbp_1 \b[8]$_DFFE_PP_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net252),
    .D(_0122_),
    .Q_N(_0039_),
    .Q(\ayayayayayaya.b[8] ));
 sg13g2_dfrbp_1 \b[9]$_DFFE_PP_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net253),
    .D(_0123_),
    .Q_N(_0040_),
    .Q(\ayayayayayaya.b[9] ));
 sg13g2_buf_1 input1 (.A(ui_in[4]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[5]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[6]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[7]),
    .X(net4));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[0]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[1]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[2]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[3]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[4]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[5]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[6]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_oe[7]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[0]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[1]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[2]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[3]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[4]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[5]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[6]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[7]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[0]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[1]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[2]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[3]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[4]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[5]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[6]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout29 (.A(_1741_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1707_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1676_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1667_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1624_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1595_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1567_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1467_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0514_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0216_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1034_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0744_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0213_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1664_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0989_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0951_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0598_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0511_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0484_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0221_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0200_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0195_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1798_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1792_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1771_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1673_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1564_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1380_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0491_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0489_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0486_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0375_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0339_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0220_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0208_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0205_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0199_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0161_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0159_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0156_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_2247_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_2220_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_2216_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_2211_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2209_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2207_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_2202_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_2127_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_2098_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1797_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1791_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1786_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1781_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1776_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1770_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1765_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1757_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1724_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1696_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1691_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1686_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1681_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1672_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0937_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0596_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0520_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0509_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0493_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0488_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0309_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0307_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0280_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0197_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0187_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0174_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_0171_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0169_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0166_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0163_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_2219_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_2215_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_2205_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_2201_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_2126_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_2112_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_2097_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_2093_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_2086_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_1796_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_1790_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_1785_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_1780_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_1775_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_1769_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_1764_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_1756_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_1732_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_1728_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_1723_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_1719_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_1715_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_1711_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_1704_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_1700_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_1695_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_1690_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_1685_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_1680_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_1671_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_1658_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_1657_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_0604_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_0574_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_0516_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_0258_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_0256_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_0203_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_0168_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_0165_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_0132_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_2218_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_2214_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_2179_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_2125_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_2096_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_2092_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_2032_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_2029_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_2009_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_2006_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_1985_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_1974_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_1964_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_1954_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_1930_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_1927_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_1905_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_1845_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_1774_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_1763_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_1735_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_1722_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_1656_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_0209_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_1838_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_1783_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_1762_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_1746_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_1744_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_1742_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_1737_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_1702_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_1698_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_1693_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_1683_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_1678_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_1669_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_1586_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_1478_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_1293_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_1315_),
    .X(net189));
 sg13g2_tiehi \a[0]$_DFFE_PP__190  (.L_HI(net190));
 sg13g2_tiehi \a[10]$_DFFE_PP__191  (.L_HI(net191));
 sg13g2_tiehi \a[11]$_DFFE_PP__192  (.L_HI(net192));
 sg13g2_tiehi \a[12]$_DFFE_PP__193  (.L_HI(net193));
 sg13g2_tiehi \a[13]$_DFFE_PP__194  (.L_HI(net194));
 sg13g2_tiehi \a[14]$_DFFE_PP__195  (.L_HI(net195));
 sg13g2_tiehi \a[15]$_DFFE_PP__196  (.L_HI(net196));
 sg13g2_tiehi \a[16]$_DFFE_PP__197  (.L_HI(net197));
 sg13g2_tiehi \a[17]$_DFFE_PP__198  (.L_HI(net198));
 sg13g2_tiehi \a[18]$_DFFE_PP__199  (.L_HI(net199));
 sg13g2_tiehi \a[19]$_DFFE_PP__200  (.L_HI(net200));
 sg13g2_tiehi \a[1]$_DFFE_PP__201  (.L_HI(net201));
 sg13g2_tiehi \a[20]$_DFFE_PP__202  (.L_HI(net202));
 sg13g2_tiehi \a[21]$_DFFE_PP__203  (.L_HI(net203));
 sg13g2_tiehi \a[22]$_DFFE_PP__204  (.L_HI(net204));
 sg13g2_tiehi \a[23]$_DFFE_PP__205  (.L_HI(net205));
 sg13g2_tiehi \a[24]$_DFFE_PP__206  (.L_HI(net206));
 sg13g2_tiehi \a[25]$_DFFE_PP__207  (.L_HI(net207));
 sg13g2_tiehi \a[26]$_DFFE_PP__208  (.L_HI(net208));
 sg13g2_tiehi \a[27]$_DFFE_PP__209  (.L_HI(net209));
 sg13g2_tiehi \a[28]$_DFFE_PP__210  (.L_HI(net210));
 sg13g2_tiehi \a[29]$_DFFE_PP__211  (.L_HI(net211));
 sg13g2_tiehi \a[2]$_DFFE_PP__212  (.L_HI(net212));
 sg13g2_tiehi \a[30]$_DFFE_PP__213  (.L_HI(net213));
 sg13g2_tiehi \a[31]$_DFFE_PP__214  (.L_HI(net214));
 sg13g2_tiehi \a[3]$_DFFE_PP__215  (.L_HI(net215));
 sg13g2_tiehi \a[4]$_DFFE_PP__216  (.L_HI(net216));
 sg13g2_tiehi \a[5]$_DFFE_PP__217  (.L_HI(net217));
 sg13g2_tiehi \a[6]$_DFFE_PP__218  (.L_HI(net218));
 sg13g2_tiehi \a[7]$_DFFE_PP__219  (.L_HI(net219));
 sg13g2_tiehi \a[8]$_DFFE_PP__220  (.L_HI(net220));
 sg13g2_tiehi \a[9]$_DFFE_PP__221  (.L_HI(net221));
 sg13g2_tiehi \b[0]$_DFFE_PP__222  (.L_HI(net222));
 sg13g2_tiehi \b[10]$_DFFE_PP__223  (.L_HI(net223));
 sg13g2_tiehi \b[11]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \b[12]$_DFFE_PP__225  (.L_HI(net225));
 sg13g2_tiehi \b[13]$_DFFE_PP__226  (.L_HI(net226));
 sg13g2_tiehi \b[14]$_DFFE_PP__227  (.L_HI(net227));
 sg13g2_tiehi \b[15]$_DFFE_PP__228  (.L_HI(net228));
 sg13g2_tiehi \b[16]$_DFFE_PP__229  (.L_HI(net229));
 sg13g2_tiehi \b[17]$_DFFE_PP__230  (.L_HI(net230));
 sg13g2_tiehi \b[18]$_DFFE_PP__231  (.L_HI(net231));
 sg13g2_tiehi \b[19]$_DFFE_PP__232  (.L_HI(net232));
 sg13g2_tiehi \b[1]$_DFFE_PP__233  (.L_HI(net233));
 sg13g2_tiehi \b[20]$_DFFE_PP__234  (.L_HI(net234));
 sg13g2_tiehi \b[21]$_DFFE_PP__235  (.L_HI(net235));
 sg13g2_tiehi \b[22]$_DFFE_PP__236  (.L_HI(net236));
 sg13g2_tiehi \b[23]$_DFFE_PP__237  (.L_HI(net237));
 sg13g2_tiehi \b[24]$_DFFE_PP__238  (.L_HI(net238));
 sg13g2_tiehi \b[25]$_DFFE_PP__239  (.L_HI(net239));
 sg13g2_tiehi \b[26]$_DFFE_PP__240  (.L_HI(net240));
 sg13g2_tiehi \b[27]$_DFFE_PP__241  (.L_HI(net241));
 sg13g2_tiehi \b[28]$_DFFE_PP__242  (.L_HI(net242));
 sg13g2_tiehi \b[29]$_DFFE_PP__243  (.L_HI(net243));
 sg13g2_tiehi \b[2]$_DFFE_PP__244  (.L_HI(net244));
 sg13g2_tiehi \b[30]$_DFFE_PP__245  (.L_HI(net245));
 sg13g2_tiehi \b[31]$_DFFE_PP__246  (.L_HI(net246));
 sg13g2_tiehi \b[3]$_DFFE_PP__247  (.L_HI(net247));
 sg13g2_tiehi \b[4]$_DFFE_PP__248  (.L_HI(net248));
 sg13g2_tiehi \b[5]$_DFFE_PP__249  (.L_HI(net249));
 sg13g2_tiehi \b[6]$_DFFE_PP__250  (.L_HI(net250));
 sg13g2_tiehi \b[7]$_DFFE_PP__251  (.L_HI(net251));
 sg13g2_tiehi \b[8]$_DFFE_PP__252  (.L_HI(net252));
 sg13g2_tiehi \b[9]$_DFFE_PP__253  (.L_HI(net253));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_4 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_4 FILLER_4_252 ();
 sg13g2_fill_2 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_262 ();
 sg13g2_decap_8 FILLER_4_269 ();
 sg13g2_decap_8 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_283 ();
 sg13g2_decap_8 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_304 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_318 ();
 sg13g2_decap_8 FILLER_4_325 ();
 sg13g2_decap_8 FILLER_4_332 ();
 sg13g2_decap_8 FILLER_4_339 ();
 sg13g2_decap_4 FILLER_4_346 ();
 sg13g2_fill_2 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_370 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_8 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_4_412 ();
 sg13g2_decap_8 FILLER_4_419 ();
 sg13g2_decap_4 FILLER_4_426 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_fill_2 FILLER_5_63 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_decap_4 FILLER_5_77 ();
 sg13g2_fill_1 FILLER_5_81 ();
 sg13g2_fill_2 FILLER_5_90 ();
 sg13g2_fill_1 FILLER_5_92 ();
 sg13g2_decap_4 FILLER_5_101 ();
 sg13g2_decap_8 FILLER_5_113 ();
 sg13g2_fill_2 FILLER_5_120 ();
 sg13g2_decap_4 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_135 ();
 sg13g2_decap_8 FILLER_5_142 ();
 sg13g2_decap_8 FILLER_5_149 ();
 sg13g2_decap_8 FILLER_5_156 ();
 sg13g2_decap_4 FILLER_5_163 ();
 sg13g2_fill_2 FILLER_5_171 ();
 sg13g2_fill_1 FILLER_5_173 ();
 sg13g2_decap_8 FILLER_5_178 ();
 sg13g2_decap_8 FILLER_5_185 ();
 sg13g2_decap_8 FILLER_5_192 ();
 sg13g2_decap_8 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_5_206 ();
 sg13g2_decap_8 FILLER_5_213 ();
 sg13g2_decap_4 FILLER_5_220 ();
 sg13g2_fill_1 FILLER_5_224 ();
 sg13g2_fill_1 FILLER_5_240 ();
 sg13g2_fill_1 FILLER_5_246 ();
 sg13g2_fill_1 FILLER_5_252 ();
 sg13g2_fill_1 FILLER_5_257 ();
 sg13g2_fill_2 FILLER_5_263 ();
 sg13g2_fill_1 FILLER_5_265 ();
 sg13g2_decap_4 FILLER_5_279 ();
 sg13g2_fill_1 FILLER_5_283 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_4 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_fill_2 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_33 ();
 sg13g2_decap_4 FILLER_6_40 ();
 sg13g2_fill_1 FILLER_6_50 ();
 sg13g2_fill_1 FILLER_6_63 ();
 sg13g2_fill_1 FILLER_6_68 ();
 sg13g2_fill_1 FILLER_6_77 ();
 sg13g2_fill_1 FILLER_6_139 ();
 sg13g2_fill_2 FILLER_6_161 ();
 sg13g2_fill_1 FILLER_6_171 ();
 sg13g2_fill_1 FILLER_6_195 ();
 sg13g2_fill_2 FILLER_6_200 ();
 sg13g2_fill_2 FILLER_6_215 ();
 sg13g2_fill_1 FILLER_6_249 ();
 sg13g2_fill_1 FILLER_6_320 ();
 sg13g2_fill_2 FILLER_6_364 ();
 sg13g2_fill_1 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_6_409 ();
 sg13g2_decap_8 FILLER_6_416 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_15 ();
 sg13g2_fill_2 FILLER_7_22 ();
 sg13g2_fill_1 FILLER_7_63 ();
 sg13g2_fill_1 FILLER_7_69 ();
 sg13g2_fill_2 FILLER_7_87 ();
 sg13g2_fill_1 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_149 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_fill_2 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_222 ();
 sg13g2_fill_1 FILLER_7_228 ();
 sg13g2_fill_1 FILLER_7_255 ();
 sg13g2_fill_2 FILLER_7_261 ();
 sg13g2_fill_2 FILLER_7_281 ();
 sg13g2_fill_1 FILLER_7_302 ();
 sg13g2_fill_1 FILLER_7_307 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_fill_2 FILLER_7_326 ();
 sg13g2_fill_1 FILLER_7_332 ();
 sg13g2_fill_1 FILLER_7_346 ();
 sg13g2_fill_1 FILLER_7_352 ();
 sg13g2_fill_1 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_decap_8 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_7_414 ();
 sg13g2_decap_8 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_fill_2 FILLER_8_28 ();
 sg13g2_fill_2 FILLER_8_66 ();
 sg13g2_fill_2 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_165 ();
 sg13g2_fill_1 FILLER_8_183 ();
 sg13g2_fill_2 FILLER_8_206 ();
 sg13g2_fill_2 FILLER_8_228 ();
 sg13g2_fill_1 FILLER_8_230 ();
 sg13g2_fill_1 FILLER_8_236 ();
 sg13g2_fill_2 FILLER_8_254 ();
 sg13g2_fill_1 FILLER_8_273 ();
 sg13g2_fill_2 FILLER_8_310 ();
 sg13g2_fill_1 FILLER_8_312 ();
 sg13g2_fill_1 FILLER_8_325 ();
 sg13g2_fill_1 FILLER_8_336 ();
 sg13g2_fill_2 FILLER_8_361 ();
 sg13g2_fill_1 FILLER_8_384 ();
 sg13g2_fill_2 FILLER_8_403 ();
 sg13g2_fill_1 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_84 ();
 sg13g2_fill_2 FILLER_9_110 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_fill_2 FILLER_9_132 ();
 sg13g2_fill_1 FILLER_9_139 ();
 sg13g2_fill_1 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_155 ();
 sg13g2_fill_2 FILLER_9_215 ();
 sg13g2_fill_2 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_265 ();
 sg13g2_fill_1 FILLER_9_284 ();
 sg13g2_fill_2 FILLER_9_313 ();
 sg13g2_fill_2 FILLER_9_340 ();
 sg13g2_fill_1 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_415 ();
 sg13g2_decap_8 FILLER_9_422 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_fill_2 FILLER_10_97 ();
 sg13g2_fill_2 FILLER_10_108 ();
 sg13g2_fill_1 FILLER_10_110 ();
 sg13g2_fill_1 FILLER_10_128 ();
 sg13g2_fill_1 FILLER_10_133 ();
 sg13g2_decap_4 FILLER_10_150 ();
 sg13g2_fill_1 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_220 ();
 sg13g2_fill_2 FILLER_10_249 ();
 sg13g2_fill_2 FILLER_10_261 ();
 sg13g2_fill_2 FILLER_10_293 ();
 sg13g2_fill_1 FILLER_10_326 ();
 sg13g2_fill_2 FILLER_10_345 ();
 sg13g2_fill_1 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_415 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_fill_2 FILLER_11_88 ();
 sg13g2_fill_1 FILLER_11_94 ();
 sg13g2_fill_1 FILLER_11_165 ();
 sg13g2_fill_2 FILLER_11_206 ();
 sg13g2_fill_2 FILLER_11_232 ();
 sg13g2_fill_1 FILLER_11_234 ();
 sg13g2_fill_1 FILLER_11_240 ();
 sg13g2_fill_2 FILLER_11_261 ();
 sg13g2_fill_2 FILLER_11_292 ();
 sg13g2_fill_1 FILLER_11_294 ();
 sg13g2_fill_1 FILLER_11_313 ();
 sg13g2_fill_1 FILLER_11_318 ();
 sg13g2_fill_1 FILLER_11_329 ();
 sg13g2_fill_1 FILLER_11_362 ();
 sg13g2_fill_2 FILLER_11_368 ();
 sg13g2_fill_1 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_421 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_37 ();
 sg13g2_fill_1 FILLER_12_62 ();
 sg13g2_fill_1 FILLER_12_104 ();
 sg13g2_fill_2 FILLER_12_114 ();
 sg13g2_fill_1 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_137 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_154 ();
 sg13g2_fill_2 FILLER_12_159 ();
 sg13g2_fill_1 FILLER_12_181 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_fill_2 FILLER_12_198 ();
 sg13g2_fill_1 FILLER_12_200 ();
 sg13g2_fill_2 FILLER_12_211 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_224 ();
 sg13g2_fill_1 FILLER_12_226 ();
 sg13g2_fill_1 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_fill_1 FILLER_12_354 ();
 sg13g2_fill_1 FILLER_12_359 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_1 FILLER_13_30 ();
 sg13g2_fill_1 FILLER_13_58 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_fill_2 FILLER_13_82 ();
 sg13g2_fill_2 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_decap_4 FILLER_13_184 ();
 sg13g2_fill_2 FILLER_13_198 ();
 sg13g2_fill_1 FILLER_13_200 ();
 sg13g2_fill_1 FILLER_13_236 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_decap_4 FILLER_13_282 ();
 sg13g2_fill_1 FILLER_13_296 ();
 sg13g2_fill_2 FILLER_13_322 ();
 sg13g2_fill_1 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_374 ();
 sg13g2_fill_1 FILLER_13_419 ();
 sg13g2_fill_2 FILLER_13_424 ();
 sg13g2_fill_1 FILLER_13_426 ();
 sg13g2_fill_1 FILLER_14_27 ();
 sg13g2_fill_1 FILLER_14_104 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_fill_1 FILLER_14_115 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_fill_1 FILLER_14_130 ();
 sg13g2_fill_2 FILLER_14_156 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_fill_2 FILLER_14_164 ();
 sg13g2_fill_1 FILLER_14_171 ();
 sg13g2_fill_1 FILLER_14_177 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_fill_1 FILLER_14_209 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_233 ();
 sg13g2_fill_1 FILLER_14_239 ();
 sg13g2_fill_2 FILLER_14_245 ();
 sg13g2_fill_2 FILLER_14_267 ();
 sg13g2_fill_2 FILLER_14_328 ();
 sg13g2_fill_1 FILLER_14_340 ();
 sg13g2_fill_1 FILLER_14_346 ();
 sg13g2_fill_1 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_363 ();
 sg13g2_fill_1 FILLER_14_395 ();
 sg13g2_fill_1 FILLER_14_401 ();
 sg13g2_fill_2 FILLER_14_421 ();
 sg13g2_fill_1 FILLER_15_22 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_102 ();
 sg13g2_fill_1 FILLER_15_113 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_166 ();
 sg13g2_fill_2 FILLER_15_177 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_192 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_fill_1 FILLER_15_251 ();
 sg13g2_fill_1 FILLER_15_257 ();
 sg13g2_fill_1 FILLER_15_263 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_1 FILLER_15_275 ();
 sg13g2_fill_1 FILLER_15_281 ();
 sg13g2_fill_1 FILLER_15_287 ();
 sg13g2_fill_2 FILLER_15_293 ();
 sg13g2_fill_2 FILLER_15_305 ();
 sg13g2_fill_1 FILLER_15_317 ();
 sg13g2_fill_2 FILLER_15_328 ();
 sg13g2_fill_1 FILLER_15_335 ();
 sg13g2_fill_2 FILLER_15_341 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_fill_1 FILLER_16_26 ();
 sg13g2_fill_2 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_62 ();
 sg13g2_fill_2 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_fill_2 FILLER_16_140 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_fill_2 FILLER_16_208 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_fill_2 FILLER_16_227 ();
 sg13g2_fill_1 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_240 ();
 sg13g2_decap_4 FILLER_16_256 ();
 sg13g2_decap_4 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_274 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_fill_2 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_343 ();
 sg13g2_fill_2 FILLER_16_350 ();
 sg13g2_fill_1 FILLER_16_352 ();
 sg13g2_fill_2 FILLER_16_362 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_fill_2 FILLER_17_24 ();
 sg13g2_fill_1 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_61 ();
 sg13g2_fill_1 FILLER_17_74 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_2 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_166 ();
 sg13g2_fill_1 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_178 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_1 FILLER_17_209 ();
 sg13g2_decap_4 FILLER_17_230 ();
 sg13g2_fill_1 FILLER_17_234 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_4 FILLER_17_271 ();
 sg13g2_fill_2 FILLER_17_335 ();
 sg13g2_fill_2 FILLER_17_367 ();
 sg13g2_fill_1 FILLER_17_384 ();
 sg13g2_fill_1 FILLER_17_390 ();
 sg13g2_fill_1 FILLER_18_37 ();
 sg13g2_fill_1 FILLER_18_49 ();
 sg13g2_fill_1 FILLER_18_104 ();
 sg13g2_fill_2 FILLER_18_167 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_fill_2 FILLER_18_251 ();
 sg13g2_fill_1 FILLER_18_258 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_325 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_376 ();
 sg13g2_fill_2 FILLER_19_32 ();
 sg13g2_fill_1 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_76 ();
 sg13g2_fill_1 FILLER_19_82 ();
 sg13g2_fill_1 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_decap_4 FILLER_19_220 ();
 sg13g2_fill_1 FILLER_19_229 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_fill_2 FILLER_19_267 ();
 sg13g2_fill_2 FILLER_19_348 ();
 sg13g2_fill_2 FILLER_19_365 ();
 sg13g2_fill_2 FILLER_20_52 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_decap_4 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_244 ();
 sg13g2_decap_4 FILLER_20_251 ();
 sg13g2_fill_1 FILLER_20_255 ();
 sg13g2_decap_4 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_1 FILLER_20_395 ();
 sg13g2_fill_1 FILLER_21_50 ();
 sg13g2_fill_1 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_158 ();
 sg13g2_fill_2 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_237 ();
 sg13g2_decap_4 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_321 ();
 sg13g2_fill_1 FILLER_21_367 ();
 sg13g2_fill_2 FILLER_22_44 ();
 sg13g2_fill_2 FILLER_22_60 ();
 sg13g2_fill_1 FILLER_22_92 ();
 sg13g2_fill_1 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_117 ();
 sg13g2_fill_1 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_fill_1 FILLER_23_48 ();
 sg13g2_fill_1 FILLER_23_111 ();
 sg13g2_fill_1 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_fill_1 FILLER_23_229 ();
 sg13g2_fill_1 FILLER_23_234 ();
 sg13g2_fill_1 FILLER_23_239 ();
 sg13g2_fill_1 FILLER_23_244 ();
 sg13g2_decap_4 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_301 ();
 sg13g2_fill_1 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_391 ();
 sg13g2_fill_1 FILLER_23_402 ();
 sg13g2_fill_1 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_24_40 ();
 sg13g2_fill_1 FILLER_24_59 ();
 sg13g2_fill_1 FILLER_24_69 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_fill_1 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_189 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_258 ();
 sg13g2_fill_1 FILLER_24_280 ();
 sg13g2_fill_2 FILLER_24_389 ();
 sg13g2_fill_2 FILLER_24_395 ();
 sg13g2_fill_2 FILLER_25_121 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_fill_1 FILLER_25_276 ();
 sg13g2_fill_2 FILLER_25_332 ();
 sg13g2_fill_1 FILLER_25_391 ();
 sg13g2_fill_1 FILLER_25_397 ();
 sg13g2_fill_1 FILLER_25_403 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_fill_1 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_58 ();
 sg13g2_fill_2 FILLER_26_78 ();
 sg13g2_fill_2 FILLER_26_125 ();
 sg13g2_fill_1 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_1 FILLER_27_29 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_60 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_121 ();
 sg13g2_fill_1 FILLER_27_134 ();
 sg13g2_fill_1 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_191 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_241 ();
 sg13g2_fill_1 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_256 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_275 ();
 sg13g2_fill_1 FILLER_27_307 ();
 sg13g2_fill_1 FILLER_27_419 ();
 sg13g2_fill_2 FILLER_27_424 ();
 sg13g2_fill_1 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_83 ();
 sg13g2_fill_1 FILLER_28_115 ();
 sg13g2_fill_1 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_fill_1 FILLER_28_238 ();
 sg13g2_fill_2 FILLER_28_386 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_fill_1 FILLER_29_59 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_173 ();
 sg13g2_fill_1 FILLER_30_26 ();
 sg13g2_fill_1 FILLER_30_42 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_138 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_fill_1 FILLER_30_424 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_fill_1 FILLER_31_181 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_252 ();
 sg13g2_fill_2 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_fill_2 FILLER_31_286 ();
 sg13g2_fill_2 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_52 ();
 sg13g2_fill_1 FILLER_32_87 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_248 ();
 sg13g2_fill_1 FILLER_32_263 ();
 sg13g2_fill_1 FILLER_32_299 ();
 sg13g2_fill_1 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_fill_2 FILLER_32_393 ();
 sg13g2_fill_2 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_fill_2 FILLER_33_274 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_fill_1 FILLER_34_113 ();
 sg13g2_fill_1 FILLER_34_195 ();
 sg13g2_fill_2 FILLER_34_233 ();
 sg13g2_fill_2 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_289 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_1 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_386 ();
 sg13g2_fill_1 FILLER_34_392 ();
 sg13g2_fill_1 FILLER_34_398 ();
 sg13g2_fill_2 FILLER_35_30 ();
 sg13g2_fill_2 FILLER_35_46 ();
 sg13g2_fill_1 FILLER_35_52 ();
 sg13g2_fill_1 FILLER_35_63 ();
 sg13g2_fill_2 FILLER_35_74 ();
 sg13g2_fill_1 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_fill_1 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_134 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_fill_2 FILLER_35_193 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_209 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_fill_2 FILLER_36_295 ();
 sg13g2_fill_1 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_397 ();
 sg13g2_fill_2 FILLER_36_402 ();
 sg13g2_fill_2 FILLER_37_60 ();
 sg13g2_fill_1 FILLER_37_161 ();
 sg13g2_fill_1 FILLER_37_192 ();
 sg13g2_fill_2 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_2 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_41 ();
 sg13g2_fill_1 FILLER_38_157 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_fill_1 FILLER_38_403 ();
endmodule
