module tt_um_oled_frequency_counter (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire clknet_0_clk;
 wire net99;
 wire \counter.cnt_ref_enable ;
 wire \counter.cnt_x_digits[0] ;
 wire \counter.cnt_x_digits[10] ;
 wire \counter.cnt_x_digits[11] ;
 wire \counter.cnt_x_digits[12] ;
 wire \counter.cnt_x_digits[13] ;
 wire \counter.cnt_x_digits[14] ;
 wire \counter.cnt_x_digits[15] ;
 wire \counter.cnt_x_digits[16] ;
 wire \counter.cnt_x_digits[17] ;
 wire \counter.cnt_x_digits[18] ;
 wire \counter.cnt_x_digits[19] ;
 wire \counter.cnt_x_digits[1] ;
 wire \counter.cnt_x_digits[20] ;
 wire \counter.cnt_x_digits[21] ;
 wire \counter.cnt_x_digits[22] ;
 wire \counter.cnt_x_digits[23] ;
 wire \counter.cnt_x_digits[2] ;
 wire \counter.cnt_x_digits[3] ;
 wire \counter.cnt_x_digits[4] ;
 wire \counter.cnt_x_digits[5] ;
 wire \counter.cnt_x_digits[6] ;
 wire \counter.cnt_x_digits[7] ;
 wire \counter.cnt_x_digits[8] ;
 wire \counter.cnt_x_digits[9] ;
 wire \counter.counter_ref.digit_0.digit_out[0] ;
 wire \counter.counter_ref.digit_0.digit_out[1] ;
 wire \counter.counter_ref.digit_0.digit_out[2] ;
 wire \counter.counter_ref.digit_0.digit_out[3] ;
 wire \counter.counter_ref.digits_out[10] ;
 wire \counter.counter_ref.digits_out[11] ;
 wire \counter.counter_ref.digits_out[12] ;
 wire \counter.counter_ref.digits_out[13] ;
 wire \counter.counter_ref.digits_out[14] ;
 wire \counter.counter_ref.digits_out[15] ;
 wire \counter.counter_ref.digits_out[16] ;
 wire \counter.counter_ref.digits_out[17] ;
 wire \counter.counter_ref.digits_out[18] ;
 wire \counter.counter_ref.digits_out[19] ;
 wire \counter.counter_ref.digits_out[20] ;
 wire \counter.counter_ref.digits_out[21] ;
 wire \counter.counter_ref.digits_out[22] ;
 wire \counter.counter_ref.digits_out[23] ;
 wire \counter.counter_ref.digits_out[4] ;
 wire \counter.counter_ref.digits_out[5] ;
 wire \counter.counter_ref.digits_out[6] ;
 wire \counter.counter_ref.digits_out[7] ;
 wire \counter.counter_ref.digits_out[8] ;
 wire \counter.counter_ref.digits_out[9] ;
 wire \counter.oled_clk_out ;
 wire \counter.oled_csn_out ;
 wire \counter.oled_dc_out ;
 wire \counter.oled_driver.mc_exec.delay_cnt[0] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[10] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[11] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[12] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[13] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[14] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[15] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[16] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[1] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[2] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[3] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[4] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[5] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[6] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[7] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[8] ;
 wire \counter.oled_driver.mc_exec.delay_cnt[9] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[0] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[1] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[2] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[3] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[4] ;
 wire \counter.oled_driver.mc_exec.microcode_rom.address[5] ;
 wire \counter.oled_driver.mc_exec.oled_dc_out ;
 wire \counter.oled_driver.mc_exec.oled_rstn_out ;
 wire \counter.oled_driver.mc_exec.oled_vbatn_out ;
 wire \counter.oled_driver.mc_exec.oled_vcdn_out ;
 wire \counter.oled_driver.mc_exec.procedure_done_out ;
 wire \counter.oled_driver.mc_exec.procedure_offset_in[0] ;
 wire \counter.oled_driver.mc_exec.procedure_start_in ;
 wire \counter.oled_driver.mc_exec.reset_in ;
 wire \counter.oled_driver.mc_exec.spi_tx_trigger_out ;
 wire \counter.oled_driver.mc_exec.state_r[0] ;
 wire \counter.oled_driver.mc_exec.state_r[2] ;
 wire \counter.oled_driver.mc_exec.state_r[3] ;
 wire \counter.oled_driver.mc_exec.state_r[5] ;
 wire \counter.oled_driver.mc_exec.state_r[6] ;
 wire \counter.oled_driver.oled_mosi_out ;
 wire \counter.oled_driver.ready_out ;
 wire \counter.oled_driver.spi_data[0] ;
 wire \counter.oled_driver.spi_data[1] ;
 wire \counter.oled_driver.spi_data[2] ;
 wire \counter.oled_driver.spi_data[3] ;
 wire \counter.oled_driver.spi_data[4] ;
 wire \counter.oled_driver.spi_data[5] ;
 wire \counter.oled_driver.spi_data[6] ;
 wire \counter.oled_driver.spi_data[7] ;
 wire \counter.oled_driver.spi_deactivate_cs ;
 wire \counter.oled_driver.spi_driver.deactivate_cs_r ;
 wire \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ;
 wire \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ;
 wire \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ;
 wire \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[0] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[5] ;
 wire \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6] ;
 wire \counter.oled_driver.spi_driver.shift_reg.start_in ;
 wire \counter.oled_driver.spi_driver.state_r[0] ;
 wire \counter.oled_driver.spi_driver.state_r[1] ;
 wire \counter.oled_driver.state_r[0] ;
 wire \counter.oled_driver.state_r[2] ;
 wire \counter.oled_driver.state_r[4] ;
 wire \counter.oled_driver.sync_stb_in ;
 wire \counter.oled_driver.write_stb_in ;
 wire \counter.refresh_display ;
 wire \counter.state[0] ;
 wire \counter.state[1] ;
 wire \counter.streamer.digit_cnt_r[0] ;
 wire \counter.streamer.digit_cnt_r[1] ;
 wire \counter.streamer.digit_cnt_r[2] ;
 wire \counter.streamer.digits_r[0] ;
 wire \counter.streamer.digits_r[10] ;
 wire \counter.streamer.digits_r[11] ;
 wire \counter.streamer.digits_r[12] ;
 wire \counter.streamer.digits_r[13] ;
 wire \counter.streamer.digits_r[14] ;
 wire \counter.streamer.digits_r[15] ;
 wire \counter.streamer.digits_r[16] ;
 wire \counter.streamer.digits_r[17] ;
 wire \counter.streamer.digits_r[18] ;
 wire \counter.streamer.digits_r[19] ;
 wire \counter.streamer.digits_r[1] ;
 wire \counter.streamer.digits_r[20] ;
 wire \counter.streamer.digits_r[21] ;
 wire \counter.streamer.digits_r[22] ;
 wire \counter.streamer.digits_r[23] ;
 wire \counter.streamer.digits_r[2] ;
 wire \counter.streamer.digits_r[3] ;
 wire \counter.streamer.digits_r[4] ;
 wire \counter.streamer.digits_r[5] ;
 wire \counter.streamer.digits_r[6] ;
 wire \counter.streamer.digits_r[7] ;
 wire \counter.streamer.digits_r[8] ;
 wire \counter.streamer.digits_r[9] ;
 wire \counter.streamer.graphical_decoder.index_x_in[0] ;
 wire \counter.streamer.graphical_decoder.index_x_in[1] ;
 wire \counter.streamer.graphical_decoder.index_x_in[2] ;
 wire \counter.streamer.graphical_decoder.index_x_in[3] ;
 wire \counter.streamer.graphical_decoder.index_x_in[4] ;
 wire \counter.streamer.graphical_decoder.index_y_in[0] ;
 wire \counter.streamer.graphical_decoder.index_y_in[1] ;
 wire \counter.streamer.graphical_decoder.pattern_adg[1] ;
 wire \counter.streamer.graphical_decoder.pattern_adg[2] ;
 wire \counter.streamer.graphical_decoder.pattern_adg[3] ;
 wire \counter.streamer.graphical_decoder.pattern_adg[4] ;
 wire \counter.streamer.ready_out ;
 wire \counter.streamer.state_r[4] ;
 wire \counter.streamer.state_r[5] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _1310_ (.A(net1),
    .X(_0634_));
 sg13g2_inv_1 _1311_ (.Y(_0635_),
    .A(net78));
 sg13g2_buf_1 _1312_ (.A(_0635_),
    .X(_0636_));
 sg13g2_buf_1 _1313_ (.A(net63),
    .X(\counter.oled_driver.mc_exec.reset_in ));
 sg13g2_buf_2 _1314_ (.A(\counter.oled_driver.mc_exec.state_r[3] ),
    .X(_0637_));
 sg13g2_inv_1 _1315_ (.Y(_0638_),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[5] ));
 sg13g2_buf_2 _1316_ (.A(\counter.oled_driver.mc_exec.microcode_rom.address[2] ),
    .X(_0639_));
 sg13g2_buf_2 _1317_ (.A(\counter.oled_driver.mc_exec.microcode_rom.address[4] ),
    .X(_0640_));
 sg13g2_a21oi_2 _1318_ (.B1(_0640_),
    .Y(_0641_),
    .A2(_0639_),
    .A1(\counter.oled_driver.mc_exec.microcode_rom.address[3] ));
 sg13g2_nor2_2 _1319_ (.A(_0638_),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_buf_1 _1320_ (.A(\counter.oled_driver.spi_driver.state_r[0] ),
    .X(_0643_));
 sg13g2_nand2_1 _1321_ (.Y(_0644_),
    .A(net77),
    .B(\counter.oled_driver.mc_exec.procedure_start_in ));
 sg13g2_buf_2 _1322_ (.A(\counter.oled_driver.mc_exec.procedure_done_out ),
    .X(_0645_));
 sg13g2_buf_1 _1323_ (.A(_0645_),
    .X(_0646_));
 sg13g2_buf_1 _1324_ (.A(net62),
    .X(_0647_));
 sg13g2_a221oi_1 _1325_ (.B2(net47),
    .C1(\counter.oled_driver.mc_exec.state_r[0] ),
    .B1(_0644_),
    .A1(_0637_),
    .Y(_0648_),
    .A2(_0642_));
 sg13g2_buf_1 _1326_ (.A(\counter.oled_driver.mc_exec.state_r[2] ),
    .X(_0649_));
 sg13g2_inv_1 _1327_ (.Y(_0650_),
    .A(net76));
 sg13g2_o21ai_1 _1328_ (.B1(_0042_),
    .Y(_0651_),
    .A1(_0638_),
    .A2(_0641_));
 sg13g2_buf_2 _1329_ (.A(_0651_),
    .X(_0652_));
 sg13g2_buf_2 _1330_ (.A(_0037_),
    .X(_0653_));
 sg13g2_inv_1 _1331_ (.Y(_0654_),
    .A(_0653_));
 sg13g2_buf_1 _1332_ (.A(_0038_),
    .X(_0655_));
 sg13g2_buf_2 _1333_ (.A(_0039_),
    .X(_0656_));
 sg13g2_a21oi_1 _1334_ (.A1(_0654_),
    .A2(net75),
    .Y(_0657_),
    .B1(_0656_));
 sg13g2_o21ai_1 _1335_ (.B1(net78),
    .Y(_0658_),
    .A1(_0642_),
    .A2(_0657_));
 sg13g2_nor4_1 _1336_ (.A(_0040_),
    .B(_0650_),
    .C(_0652_),
    .D(_0658_),
    .Y(_0659_));
 sg13g2_buf_2 _1337_ (.A(_0033_),
    .X(_0660_));
 sg13g2_a21o_1 _1338_ (.A2(_0639_),
    .A1(\counter.oled_driver.mc_exec.microcode_rom.address[3] ),
    .B1(_0640_),
    .X(_0661_));
 sg13g2_nand2_1 _1339_ (.Y(_0662_),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[5] ),
    .B(_0661_));
 sg13g2_buf_1 _1340_ (.A(_0662_),
    .X(_0663_));
 sg13g2_and2_1 _1341_ (.A(_0660_),
    .B(net37),
    .X(_0664_));
 sg13g2_nor3_2 _1342_ (.A(_0040_),
    .B(_0653_),
    .C(_0656_),
    .Y(_0665_));
 sg13g2_buf_2 _1343_ (.A(_0034_),
    .X(_0666_));
 sg13g2_buf_1 _1344_ (.A(_0035_),
    .X(_0667_));
 sg13g2_buf_1 _1345_ (.A(_0036_),
    .X(_0668_));
 sg13g2_nor4_1 _1346_ (.A(_0666_),
    .B(net74),
    .C(net73),
    .D(net75),
    .Y(_0669_));
 sg13g2_nand4_1 _1347_ (.B(_0664_),
    .C(_0665_),
    .A(_0659_),
    .Y(_0670_),
    .D(_0669_));
 sg13g2_o21ai_1 _1348_ (.B1(_0670_),
    .Y(_0019_),
    .A1(net63),
    .A2(_0648_));
 sg13g2_a22oi_1 _1349_ (.Y(_0671_),
    .B1(\counter.oled_driver.state_r[2] ),
    .B2(net47),
    .A2(\counter.oled_driver.state_r[4] ),
    .A1(_0643_));
 sg13g2_buf_1 _1350_ (.A(\counter.oled_driver.ready_out ),
    .X(_0672_));
 sg13g2_buf_1 _1351_ (.A(_0672_),
    .X(_0673_));
 sg13g2_nor2_1 _1352_ (.A(\counter.oled_driver.sync_stb_in ),
    .B(\counter.oled_driver.write_stb_in ),
    .Y(_0674_));
 sg13g2_nand2_1 _1353_ (.Y(_0675_),
    .A(_0673_),
    .B(_0674_));
 sg13g2_buf_1 _1354_ (.A(_0635_),
    .X(_0676_));
 sg13g2_a21oi_1 _1355_ (.A1(_0671_),
    .A2(_0675_),
    .Y(_0026_),
    .B1(_0676_));
 sg13g2_inv_1 _1356_ (.Y(_0677_),
    .A(net77));
 sg13g2_nor2_1 _1357_ (.A(_0677_),
    .B(_0051_),
    .Y(_0678_));
 sg13g2_and2_1 _1358_ (.A(net61),
    .B(\counter.oled_driver.sync_stb_in ),
    .X(_0679_));
 sg13g2_a221oi_1 _1359_ (.B2(_0678_),
    .C1(_0679_),
    .B1(\counter.oled_driver.state_r[0] ),
    .A1(\counter.oled_driver.mc_exec.procedure_start_in ),
    .Y(_0680_),
    .A2(net47));
 sg13g2_nor2_1 _1360_ (.A(net48),
    .B(_0680_),
    .Y(_0025_));
 sg13g2_inv_1 _1361_ (.Y(_0681_),
    .A(\counter.oled_driver.mc_exec.delay_cnt[4] ));
 sg13g2_nor4_1 _1362_ (.A(\counter.oled_driver.mc_exec.delay_cnt[1] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[0] ),
    .C(\counter.oled_driver.mc_exec.delay_cnt[3] ),
    .D(\counter.oled_driver.mc_exec.delay_cnt[2] ),
    .Y(_0682_));
 sg13g2_nor3_1 _1363_ (.A(\counter.oled_driver.mc_exec.delay_cnt[5] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[6] ),
    .C(\counter.oled_driver.mc_exec.delay_cnt[10] ),
    .Y(_0683_));
 sg13g2_nor3_1 _1364_ (.A(\counter.oled_driver.mc_exec.delay_cnt[7] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[9] ),
    .C(\counter.oled_driver.mc_exec.delay_cnt[8] ),
    .Y(_0684_));
 sg13g2_nand4_1 _1365_ (.B(_0682_),
    .C(_0683_),
    .A(_0681_),
    .Y(_0685_),
    .D(_0684_));
 sg13g2_nor3_1 _1366_ (.A(\counter.oled_driver.mc_exec.delay_cnt[11] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[12] ),
    .C(_0685_),
    .Y(_0686_));
 sg13g2_nor2b_1 _1367_ (.A(\counter.oled_driver.mc_exec.delay_cnt[13] ),
    .B_N(_0686_),
    .Y(_0687_));
 sg13g2_nand2b_1 _1368_ (.Y(_0688_),
    .B(_0687_),
    .A_N(\counter.oled_driver.mc_exec.delay_cnt[14] ));
 sg13g2_nor2_1 _1369_ (.A(\counter.oled_driver.mc_exec.delay_cnt[15] ),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_nand3_1 _1370_ (.B(\counter.oled_driver.mc_exec.state_r[6] ),
    .C(_0689_),
    .A(_0052_),
    .Y(_0690_));
 sg13g2_inv_1 _1371_ (.Y(_0691_),
    .A(_0040_));
 sg13g2_nor4_2 _1372_ (.A(_0666_),
    .B(_0035_),
    .C(net73),
    .Y(_0692_),
    .D(_0660_));
 sg13g2_o21ai_1 _1373_ (.B1(_0665_),
    .Y(_0693_),
    .A1(net75),
    .A2(_0692_));
 sg13g2_nor2_1 _1374_ (.A(_0650_),
    .B(_0642_),
    .Y(_0694_));
 sg13g2_nand2_1 _1375_ (.Y(_0695_),
    .A(_0042_),
    .B(_0694_));
 sg13g2_a21oi_1 _1376_ (.A1(_0691_),
    .A2(_0693_),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_a21oi_1 _1377_ (.A1(net77),
    .A2(\counter.oled_driver.mc_exec.state_r[5] ),
    .Y(_0697_),
    .B1(_0696_));
 sg13g2_a21oi_1 _1378_ (.A1(_0690_),
    .A2(_0697_),
    .Y(_0018_),
    .B1(net60));
 sg13g2_nand2_1 _1379_ (.Y(_0698_),
    .A(net77),
    .B(\counter.oled_driver.mc_exec.spi_tx_trigger_out ));
 sg13g2_nand2_1 _1380_ (.Y(_0699_),
    .A(net76),
    .B(_0652_));
 sg13g2_a21oi_1 _1381_ (.A1(_0698_),
    .A2(_0699_),
    .Y(_0016_),
    .B1(net60));
 sg13g2_and4_1 _1382_ (.A(net1),
    .B(\counter.oled_driver.spi_driver.state_r[0] ),
    .C(\counter.oled_driver.mc_exec.procedure_start_in ),
    .D(_0645_),
    .X(_0700_));
 sg13g2_buf_1 _1383_ (.A(_0634_),
    .X(_0701_));
 sg13g2_nand2_1 _1384_ (.Y(_0702_),
    .A(_0665_),
    .B(_0669_));
 sg13g2_a22oi_1 _1385_ (.Y(_0703_),
    .B1(_0659_),
    .B2(_0702_),
    .A2(_0637_),
    .A1(net72));
 sg13g2_nor2_1 _1386_ (.A(_0642_),
    .B(_0703_),
    .Y(_0704_));
 sg13g2_or2_1 _1387_ (.X(_0017_),
    .B(_0704_),
    .A(_0700_));
 sg13g2_a22oi_1 _1388_ (.Y(_0705_),
    .B1(\counter.oled_driver.spi_deactivate_cs ),
    .B2(net77),
    .A2(\counter.oled_driver.write_stb_in ),
    .A1(net61));
 sg13g2_nor2_1 _1389_ (.A(\counter.oled_driver.mc_exec.reset_in ),
    .B(_0705_),
    .Y(_0024_));
 sg13g2_buf_2 _1390_ (.A(\counter.streamer.ready_out ),
    .X(_0706_));
 sg13g2_nand2b_2 _1391_ (.Y(_0707_),
    .B(_0706_),
    .A_N(\counter.refresh_display ));
 sg13g2_buf_1 _1392_ (.A(\counter.counter_ref.digits_out[21] ),
    .X(_0708_));
 sg13g2_nor2b_1 _1393_ (.A(\counter.counter_ref.digits_out[22] ),
    .B_N(\counter.counter_ref.digits_out[23] ),
    .Y(_0709_));
 sg13g2_nand3b_1 _1394_ (.B(_0709_),
    .C(\counter.counter_ref.digits_out[20] ),
    .Y(_0710_),
    .A_N(_0708_));
 sg13g2_inv_1 _1395_ (.Y(_0711_),
    .A(_0710_));
 sg13g2_buf_1 _1396_ (.A(\counter.counter_ref.digits_out[17] ),
    .X(_0712_));
 sg13g2_inv_1 _1397_ (.Y(_0713_),
    .A(\counter.counter_ref.digits_out[13] ));
 sg13g2_nor2b_1 _1398_ (.A(\counter.counter_ref.digits_out[14] ),
    .B_N(\counter.counter_ref.digits_out[15] ),
    .Y(_0714_));
 sg13g2_nand4_1 _1399_ (.B(_0713_),
    .C(\counter.counter_ref.digits_out[16] ),
    .A(\counter.counter_ref.digits_out[12] ),
    .Y(_0715_),
    .D(_0714_));
 sg13g2_nand2b_1 _1400_ (.Y(_0716_),
    .B(net1),
    .A_N(\counter.state[0] ));
 sg13g2_buf_1 _1401_ (.A(_0716_),
    .X(_0717_));
 sg13g2_inv_1 _1402_ (.Y(_0718_),
    .A(\counter.counter_ref.digits_out[18] ));
 sg13g2_nand2_1 _1403_ (.Y(_0719_),
    .A(_0718_),
    .B(\counter.counter_ref.digits_out[19] ));
 sg13g2_or4_1 _1404_ (.A(_0712_),
    .B(_0715_),
    .C(net59),
    .D(_0719_),
    .X(_0720_));
 sg13g2_buf_1 _1405_ (.A(\counter.cnt_ref_enable ),
    .X(_0721_));
 sg13g2_nand2b_1 _1406_ (.Y(_0722_),
    .B(\counter.counter_ref.digits_out[11] ),
    .A_N(\counter.counter_ref.digits_out[10] ));
 sg13g2_inv_1 _1407_ (.Y(_0723_),
    .A(\counter.counter_ref.digits_out[5] ));
 sg13g2_nor2b_1 _1408_ (.A(\counter.counter_ref.digits_out[6] ),
    .B_N(\counter.counter_ref.digits_out[7] ),
    .Y(_0724_));
 sg13g2_nand4_1 _1409_ (.B(_0723_),
    .C(\counter.counter_ref.digits_out[8] ),
    .A(\counter.counter_ref.digits_out[4] ),
    .Y(_0725_),
    .D(_0724_));
 sg13g2_inv_1 _1410_ (.Y(_0726_),
    .A(\counter.counter_ref.digit_0.digit_out[0] ));
 sg13g2_buf_1 _1411_ (.A(\counter.counter_ref.digit_0.digit_out[1] ),
    .X(_0727_));
 sg13g2_nand2b_1 _1412_ (.Y(_0728_),
    .B(\counter.counter_ref.digit_0.digit_out[3] ),
    .A_N(\counter.counter_ref.digit_0.digit_out[2] ));
 sg13g2_nor4_2 _1413_ (.A(_0726_),
    .B(_0727_),
    .C(net59),
    .Y(_0729_),
    .D(_0728_));
 sg13g2_inv_1 _1414_ (.Y(_0730_),
    .A(_0729_));
 sg13g2_nor4_2 _1415_ (.A(\counter.counter_ref.digits_out[9] ),
    .B(_0722_),
    .C(_0725_),
    .Y(_0731_),
    .D(_0730_));
 sg13g2_nand2_1 _1416_ (.Y(_0732_),
    .A(_0721_),
    .B(_0731_));
 sg13g2_nor2_2 _1417_ (.A(_0720_),
    .B(_0732_),
    .Y(_0733_));
 sg13g2_a22oi_1 _1418_ (.Y(_0734_),
    .B1(_0711_),
    .B2(_0733_),
    .A2(_0707_),
    .A1(\counter.state[1] ));
 sg13g2_nor2_1 _1419_ (.A(net48),
    .B(_0734_),
    .Y(_0028_));
 sg13g2_buf_1 _1420_ (.A(net72),
    .X(_0735_));
 sg13g2_buf_1 _1421_ (.A(\counter.refresh_display ),
    .X(_0736_));
 sg13g2_buf_1 _1422_ (.A(_0706_),
    .X(_0737_));
 sg13g2_nand3b_1 _1423_ (.B(\counter.state[1] ),
    .C(net57),
    .Y(_0738_),
    .A_N(net70));
 sg13g2_nand2b_1 _1424_ (.Y(_0739_),
    .B(\counter.state[0] ),
    .A_N(net57));
 sg13g2_nand3_1 _1425_ (.B(_0738_),
    .C(_0739_),
    .A(net58),
    .Y(_0027_));
 sg13g2_inv_1 _1426_ (.Y(_0740_),
    .A(\counter.oled_driver.state_r[0] ));
 sg13g2_o21ai_1 _1427_ (.B1(net58),
    .Y(_0023_),
    .A1(_0740_),
    .A2(_0678_));
 sg13g2_buf_1 _1428_ (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ),
    .X(_0741_));
 sg13g2_nor3_1 _1429_ (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ),
    .B(_0741_),
    .C(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ),
    .Y(_0742_));
 sg13g2_nor2b_1 _1430_ (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ),
    .B_N(_0742_),
    .Y(_0743_));
 sg13g2_buf_1 _1431_ (.A(_0743_),
    .X(_0744_));
 sg13g2_buf_1 _1432_ (.A(net36),
    .X(_0745_));
 sg13g2_nand2_1 _1433_ (.Y(_0746_),
    .A(net72),
    .B(net30));
 sg13g2_mux2_1 _1434_ (.A0(\counter.oled_driver.mc_exec.spi_tx_trigger_out ),
    .A1(\counter.oled_driver.spi_deactivate_cs ),
    .S(net62),
    .X(_0747_));
 sg13g2_buf_1 _1435_ (.A(\counter.oled_driver.spi_driver.shift_reg.start_in ),
    .X(_0748_));
 sg13g2_buf_1 _1436_ (.A(net69),
    .X(_0749_));
 sg13g2_a21oi_1 _1437_ (.A1(net77),
    .A2(_0747_),
    .Y(_0750_),
    .B1(net56));
 sg13g2_nor2_1 _1438_ (.A(_0746_),
    .B(_0750_),
    .Y(_0022_));
 sg13g2_inv_1 _1439_ (.Y(_0751_),
    .A(\counter.streamer.graphical_decoder.index_x_in[3] ));
 sg13g2_buf_2 _1440_ (.A(\counter.streamer.graphical_decoder.index_x_in[2] ),
    .X(_0752_));
 sg13g2_buf_1 _1441_ (.A(\counter.streamer.graphical_decoder.index_x_in[1] ),
    .X(_0753_));
 sg13g2_buf_2 _1442_ (.A(\counter.streamer.graphical_decoder.index_x_in[0] ),
    .X(_0754_));
 sg13g2_nor2_1 _1443_ (.A(net68),
    .B(_0754_),
    .Y(_0755_));
 sg13g2_nand4_1 _1444_ (.B(_0752_),
    .C(\counter.streamer.graphical_decoder.index_x_in[4] ),
    .A(_0751_),
    .Y(_0756_),
    .D(_0755_));
 sg13g2_buf_1 _1445_ (.A(\counter.streamer.graphical_decoder.index_y_in[0] ),
    .X(_0757_));
 sg13g2_buf_1 _1446_ (.A(\counter.streamer.graphical_decoder.index_y_in[1] ),
    .X(_0758_));
 sg13g2_buf_1 _1447_ (.A(_0758_),
    .X(_0759_));
 sg13g2_buf_8 _1448_ (.A(\counter.streamer.digit_cnt_r[0] ),
    .X(_0760_));
 sg13g2_buf_8 _1449_ (.A(\counter.streamer.digit_cnt_r[1] ),
    .X(_0761_));
 sg13g2_buf_8 _1450_ (.A(_0761_),
    .X(_0762_));
 sg13g2_buf_1 _1451_ (.A(\counter.streamer.digit_cnt_r[2] ),
    .X(_0763_));
 sg13g2_nor3_1 _1452_ (.A(net66),
    .B(_0762_),
    .C(net65),
    .Y(_0764_));
 sg13g2_nand3_1 _1453_ (.B(net55),
    .C(_0764_),
    .A(net67),
    .Y(_0765_));
 sg13g2_nor2_1 _1454_ (.A(_0756_),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_buf_1 _1455_ (.A(\counter.streamer.state_r[5] ),
    .X(_0767_));
 sg13g2_nor2b_1 _1456_ (.A(_0050_),
    .B_N(net64),
    .Y(_0768_));
 sg13g2_a21oi_1 _1457_ (.A1(_0766_),
    .A2(_0768_),
    .Y(_0769_),
    .B1(_0679_));
 sg13g2_nor2_1 _1458_ (.A(\counter.oled_driver.mc_exec.reset_in ),
    .B(_0769_),
    .Y(_0030_));
 sg13g2_and2_1 _1459_ (.A(_0743_),
    .B(_0747_),
    .X(_0770_));
 sg13g2_a21oi_1 _1460_ (.A1(\counter.oled_driver.spi_driver.state_r[1] ),
    .A2(net30),
    .Y(_0771_),
    .B1(_0636_));
 sg13g2_o21ai_1 _1461_ (.B1(_0771_),
    .Y(_0021_),
    .A1(_0677_),
    .A2(_0770_));
 sg13g2_nor2_1 _1462_ (.A(_0710_),
    .B(_0720_),
    .Y(_0772_));
 sg13g2_nand2_1 _1463_ (.Y(_0773_),
    .A(_0731_),
    .B(_0772_));
 sg13g2_nand2_1 _1464_ (.Y(_0774_),
    .A(net71),
    .B(_0773_));
 sg13g2_buf_1 _1465_ (.A(_0706_),
    .X(_0775_));
 sg13g2_nand2_1 _1466_ (.Y(_0776_),
    .A(net53),
    .B(\counter.state[0] ));
 sg13g2_a21oi_1 _1467_ (.A1(_0774_),
    .A2(_0776_),
    .Y(_0029_),
    .B1(net60));
 sg13g2_a22oi_1 _1468_ (.Y(_0777_),
    .B1(\counter.oled_driver.write_stb_in ),
    .B2(net61),
    .A2(net70),
    .A1(net57));
 sg13g2_o21ai_1 _1469_ (.B1(_0768_),
    .Y(_0778_),
    .A1(_0756_),
    .A2(_0765_));
 sg13g2_buf_1 _1470_ (.A(net63),
    .X(_0779_));
 sg13g2_a21oi_1 _1471_ (.A1(_0777_),
    .A2(_0778_),
    .Y(_0031_),
    .B1(net46));
 sg13g2_nor3_1 _1472_ (.A(_0040_),
    .B(_0650_),
    .C(_0652_),
    .Y(_0780_));
 sg13g2_nand2_1 _1473_ (.Y(_0781_),
    .A(_0052_),
    .B(_0689_));
 sg13g2_a22oi_1 _1474_ (.Y(_0782_),
    .B1(_0781_),
    .B2(\counter.oled_driver.mc_exec.state_r[6] ),
    .A2(_0780_),
    .A1(_0656_));
 sg13g2_nor2_1 _1475_ (.A(net48),
    .B(_0782_),
    .Y(_0020_));
 sg13g2_a21oi_1 _1476_ (.A1(net61),
    .A2(\counter.streamer.state_r[4] ),
    .Y(_0783_),
    .B1(\counter.oled_driver.mc_exec.state_r[0] ));
 sg13g2_a21oi_1 _1477_ (.A1(_0707_),
    .A2(_0783_),
    .Y(_0032_),
    .B1(net46));
 sg13g2_or4_1 _1478_ (.A(_0666_),
    .B(_0035_),
    .C(_0036_),
    .D(_0660_),
    .X(_0784_));
 sg13g2_nor3_1 _1479_ (.A(_0653_),
    .B(net75),
    .C(_0784_),
    .Y(_0785_));
 sg13g2_o21ai_1 _1480_ (.B1(net75),
    .Y(_0786_),
    .A1(_0653_),
    .A2(_0784_));
 sg13g2_nand2b_1 _1481_ (.Y(_0787_),
    .B(_0786_),
    .A_N(_0785_));
 sg13g2_o21ai_1 _1482_ (.B1(net76),
    .Y(_0788_),
    .A1(_0642_),
    .A2(_0787_));
 sg13g2_buf_2 _1483_ (.A(\counter.oled_driver.mc_exec.microcode_rom.address[1] ),
    .X(_0789_));
 sg13g2_nor2b_1 _1484_ (.A(_0058_),
    .B_N(_0640_),
    .Y(_0790_));
 sg13g2_nand4_1 _1485_ (.B(_0639_),
    .C(_0789_),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[3] ),
    .Y(_0791_),
    .D(_0790_));
 sg13g2_xnor2_1 _1486_ (.Y(_0792_),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[5] ),
    .B(_0791_));
 sg13g2_a22oi_1 _1487_ (.Y(_0793_),
    .B1(_0792_),
    .B2(_0637_),
    .A2(\counter.oled_driver.mc_exec.procedure_offset_in[0] ),
    .A1(_0645_));
 sg13g2_inv_1 _1488_ (.Y(_0794_),
    .A(_0051_));
 sg13g2_nor3_2 _1489_ (.A(\counter.oled_driver.mc_exec.state_r[2] ),
    .B(_0637_),
    .C(_0794_),
    .Y(_0795_));
 sg13g2_a21oi_1 _1490_ (.A1(_0788_),
    .A2(_0793_),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_inv_1 _1491_ (.Y(_0797_),
    .A(_0042_));
 sg13g2_a21oi_1 _1492_ (.A1(\counter.oled_driver.mc_exec.microcode_rom.address[5] ),
    .A2(_0661_),
    .Y(_0798_),
    .B1(_0797_));
 sg13g2_inv_1 _1493_ (.Y(_0799_),
    .A(_0645_));
 sg13g2_or3_1 _1494_ (.A(\counter.oled_driver.mc_exec.state_r[0] ),
    .B(\counter.oled_driver.mc_exec.state_r[2] ),
    .C(_0637_),
    .X(_0800_));
 sg13g2_a21oi_1 _1495_ (.A1(_0799_),
    .A2(_0800_),
    .Y(_0801_),
    .B1(_0700_));
 sg13g2_nor3_1 _1496_ (.A(_0638_),
    .B(_0054_),
    .C(_0641_),
    .Y(_0802_));
 sg13g2_nor4_1 _1497_ (.A(\counter.oled_driver.mc_exec.state_r[2] ),
    .B(_0798_),
    .C(_0801_),
    .D(_0802_),
    .Y(_0803_));
 sg13g2_buf_1 _1498_ (.A(_0053_),
    .X(_0804_));
 sg13g2_nor2_1 _1499_ (.A(_0652_),
    .B(_0801_),
    .Y(_0805_));
 sg13g2_and2_1 _1500_ (.A(_0804_),
    .B(_0805_),
    .X(_0806_));
 sg13g2_nor4_1 _1501_ (.A(_0691_),
    .B(_0656_),
    .C(_0652_),
    .D(_0785_),
    .Y(_0807_));
 sg13g2_nor2_1 _1502_ (.A(_0666_),
    .B(_0660_),
    .Y(_0808_));
 sg13g2_nand2_1 _1503_ (.Y(_0809_),
    .A(_0035_),
    .B(net73));
 sg13g2_o21ai_1 _1504_ (.B1(_0654_),
    .Y(_0810_),
    .A1(_0808_),
    .A2(_0809_));
 sg13g2_a21oi_1 _1505_ (.A1(net75),
    .A2(_0810_),
    .Y(_0811_),
    .B1(_0801_));
 sg13g2_and2_1 _1506_ (.A(_0807_),
    .B(_0811_),
    .X(_0812_));
 sg13g2_or3_1 _1507_ (.A(_0803_),
    .B(_0806_),
    .C(_0812_),
    .X(_0813_));
 sg13g2_buf_2 _1508_ (.A(_0813_),
    .X(_0814_));
 sg13g2_mux2_1 _1509_ (.A0(\counter.oled_driver.mc_exec.microcode_rom.address[5] ),
    .A1(_0796_),
    .S(_0814_),
    .X(_0815_));
 sg13g2_nand2_2 _1510_ (.Y(_0816_),
    .A(net78),
    .B(_0815_));
 sg13g2_inv_1 _1511_ (.Y(_0148_),
    .A(_0816_));
 sg13g2_buf_1 _1512_ (.A(\counter.oled_driver.mc_exec.microcode_rom.address[0] ),
    .X(_0817_));
 sg13g2_nand2_1 _1513_ (.Y(_0818_),
    .A(_0789_),
    .B(_0817_));
 sg13g2_xor2_1 _1514_ (.B(_0818_),
    .A(_0056_),
    .X(_0819_));
 sg13g2_nor2_1 _1515_ (.A(_0054_),
    .B(_0795_),
    .Y(_0820_));
 sg13g2_nor3_1 _1516_ (.A(_0666_),
    .B(net74),
    .C(_0660_),
    .Y(_0821_));
 sg13g2_nor2b_1 _1517_ (.A(_0808_),
    .B_N(net74),
    .Y(_0822_));
 sg13g2_or3_1 _1518_ (.A(_0642_),
    .B(_0821_),
    .C(_0822_),
    .X(_0823_));
 sg13g2_a22oi_1 _1519_ (.Y(_0824_),
    .B1(_0823_),
    .B2(net76),
    .A2(_0820_),
    .A1(_0819_));
 sg13g2_a221oi_1 _1520_ (.B2(_0811_),
    .C1(_0803_),
    .B1(_0807_),
    .A1(_0804_),
    .Y(_0825_),
    .A2(_0805_));
 sg13g2_buf_2 _1521_ (.A(_0825_),
    .X(_0826_));
 sg13g2_mux2_1 _1522_ (.A0(_0824_),
    .A1(_0056_),
    .S(_0826_),
    .X(_0827_));
 sg13g2_buf_2 _1523_ (.A(_0827_),
    .X(_0828_));
 sg13g2_xor2_1 _1524_ (.B(_0660_),
    .A(_0666_),
    .X(_0829_));
 sg13g2_a21o_1 _1525_ (.A2(_0829_),
    .A1(_0662_),
    .B1(_0804_),
    .X(_0830_));
 sg13g2_xor2_1 _1526_ (.B(_0817_),
    .A(_0789_),
    .X(_0831_));
 sg13g2_nand2b_1 _1527_ (.Y(_0832_),
    .B(_0831_),
    .A_N(_0054_));
 sg13g2_a21oi_1 _1528_ (.A1(_0830_),
    .A2(_0832_),
    .Y(_0833_),
    .B1(_0795_));
 sg13g2_inv_1 _1529_ (.Y(_0834_),
    .A(_0059_));
 sg13g2_mux2_1 _1530_ (.A0(_0833_),
    .A1(_0834_),
    .S(_0826_),
    .X(_0835_));
 sg13g2_buf_2 _1531_ (.A(_0835_),
    .X(_0836_));
 sg13g2_nor2b_1 _1532_ (.A(_0828_),
    .B_N(_0836_),
    .Y(_0837_));
 sg13g2_nand2_1 _1533_ (.Y(_0838_),
    .A(_0645_),
    .B(\counter.oled_driver.mc_exec.procedure_offset_in[0] ));
 sg13g2_nand2_1 _1534_ (.Y(_0839_),
    .A(_0817_),
    .B(_0838_));
 sg13g2_nand3_1 _1535_ (.B(_0662_),
    .C(_0838_),
    .A(_0660_),
    .Y(_0840_));
 sg13g2_nor2_1 _1536_ (.A(_0051_),
    .B(_0838_),
    .Y(_0841_));
 sg13g2_a221oi_1 _1537_ (.B2(net76),
    .C1(_0841_),
    .B1(_0840_),
    .A1(_0637_),
    .Y(_0842_),
    .A2(_0839_));
 sg13g2_mux2_1 _1538_ (.A0(_0842_),
    .A1(_0058_),
    .S(_0826_),
    .X(_0843_));
 sg13g2_buf_8 _1539_ (.A(_0843_),
    .X(_0844_));
 sg13g2_inv_2 _1540_ (.Y(_0845_),
    .A(_0844_));
 sg13g2_xor2_1 _1541_ (.B(_0821_),
    .A(net73),
    .X(_0846_));
 sg13g2_o21ai_1 _1542_ (.B1(_0649_),
    .Y(_0847_),
    .A1(_0642_),
    .A2(_0846_));
 sg13g2_nand3_1 _1543_ (.B(_0789_),
    .C(_0817_),
    .A(_0639_),
    .Y(_0848_));
 sg13g2_xor2_1 _1544_ (.B(_0848_),
    .A(_0057_),
    .X(_0849_));
 sg13g2_nand2b_1 _1545_ (.Y(_0850_),
    .B(_0849_),
    .A_N(_0054_));
 sg13g2_a21o_1 _1546_ (.A2(_0850_),
    .A1(_0847_),
    .B1(_0795_),
    .X(_0851_));
 sg13g2_mux2_1 _1547_ (.A0(_0851_),
    .A1(_0057_),
    .S(_0826_),
    .X(_0852_));
 sg13g2_buf_1 _1548_ (.A(_0852_),
    .X(_0853_));
 sg13g2_o21ai_1 _1549_ (.B1(net21),
    .Y(_0854_),
    .A1(_0837_),
    .A2(net19));
 sg13g2_buf_1 _1550_ (.A(_0815_),
    .X(_0855_));
 sg13g2_nor2_1 _1551_ (.A(_0635_),
    .B(net18),
    .Y(_0856_));
 sg13g2_buf_1 _1552_ (.A(_0856_),
    .X(_0857_));
 sg13g2_buf_8 _1553_ (.A(_0826_),
    .X(_0858_));
 sg13g2_nand2b_1 _1554_ (.Y(_0859_),
    .B(net24),
    .A_N(_0057_));
 sg13g2_o21ai_1 _1555_ (.B1(_0859_),
    .Y(_0860_),
    .A1(net24),
    .A2(_0851_));
 sg13g2_buf_1 _1556_ (.A(_0860_),
    .X(_0861_));
 sg13g2_buf_1 _1557_ (.A(_0828_),
    .X(_0862_));
 sg13g2_nor2_1 _1558_ (.A(_0640_),
    .B(_0058_),
    .Y(_0863_));
 sg13g2_nand4_1 _1559_ (.B(_0639_),
    .C(_0789_),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[3] ),
    .Y(_0864_),
    .D(_0817_));
 sg13g2_xor2_1 _1560_ (.B(_0864_),
    .A(_0640_),
    .X(_0865_));
 sg13g2_or2_1 _1561_ (.X(_0866_),
    .B(_0865_),
    .A(_0054_));
 sg13g2_xnor2_1 _1562_ (.Y(_0867_),
    .A(_0653_),
    .B(_0692_));
 sg13g2_a21o_1 _1563_ (.A2(_0867_),
    .A1(_0662_),
    .B1(_0804_),
    .X(_0868_));
 sg13g2_a21oi_2 _1564_ (.B1(_0795_),
    .Y(_0869_),
    .A2(_0868_),
    .A1(_0866_));
 sg13g2_nor3_1 _1565_ (.A(net24),
    .B(_0842_),
    .C(_0869_),
    .Y(_0870_));
 sg13g2_a21o_1 _1566_ (.A2(_0863_),
    .A1(net24),
    .B1(_0870_),
    .X(_0871_));
 sg13g2_or2_1 _1567_ (.X(_0872_),
    .B(_0871_),
    .A(_0862_));
 sg13g2_nor2_1 _1568_ (.A(net13),
    .B(_0872_),
    .Y(_0873_));
 sg13g2_a22oi_1 _1569_ (.Y(_0874_),
    .B1(net12),
    .B2(_0873_),
    .A2(_0854_),
    .A1(_0148_));
 sg13g2_buf_1 _1570_ (.A(net72),
    .X(_0875_));
 sg13g2_buf_1 _1571_ (.A(_0836_),
    .X(_0876_));
 sg13g2_and2_1 _1572_ (.A(_0853_),
    .B(_0828_),
    .X(_0877_));
 sg13g2_buf_1 _1573_ (.A(_0877_),
    .X(_0878_));
 sg13g2_mux2_1 _1574_ (.A0(_0869_),
    .A1(_0640_),
    .S(net24),
    .X(_0879_));
 sg13g2_buf_8 _1575_ (.A(_0879_),
    .X(_0880_));
 sg13g2_nor2_1 _1576_ (.A(net22),
    .B(net15),
    .Y(_0881_));
 sg13g2_a22oi_1 _1577_ (.Y(_0882_),
    .B1(_0881_),
    .B2(net13),
    .A2(_0878_),
    .A1(net16));
 sg13g2_o21ai_1 _1578_ (.B1(_0837_),
    .Y(_0883_),
    .A1(net18),
    .A2(net13));
 sg13g2_o21ai_1 _1579_ (.B1(_0883_),
    .Y(_0884_),
    .A1(_0855_),
    .A2(_0882_));
 sg13g2_nand3_1 _1580_ (.B(net19),
    .C(_0884_),
    .A(net52),
    .Y(_0885_));
 sg13g2_buf_1 _1581_ (.A(_0844_),
    .X(_0886_));
 sg13g2_inv_1 _1582_ (.Y(_0887_),
    .A(_0828_));
 sg13g2_and2_1 _1583_ (.A(_0640_),
    .B(_0858_),
    .X(_0888_));
 sg13g2_a21oi_2 _1584_ (.B1(_0888_),
    .Y(_0889_),
    .A2(_0869_),
    .A1(_0814_));
 sg13g2_nor2_1 _1585_ (.A(net22),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_nand2_1 _1586_ (.Y(_0891_),
    .A(net22),
    .B(_0828_));
 sg13g2_nor2_1 _1587_ (.A(_0891_),
    .B(net15),
    .Y(_0892_));
 sg13g2_a21o_1 _1588_ (.A2(_0890_),
    .A1(_0887_),
    .B1(_0892_),
    .X(_0893_));
 sg13g2_nand3_1 _1589_ (.B(net12),
    .C(_0893_),
    .A(net14),
    .Y(_0894_));
 sg13g2_nand3_1 _1590_ (.B(_0885_),
    .C(_0894_),
    .A(_0874_),
    .Y(_0000_));
 sg13g2_nor2b_1 _1591_ (.A(net21),
    .B_N(net16),
    .Y(_0895_));
 sg13g2_nor2_1 _1592_ (.A(_0887_),
    .B(net19),
    .Y(_0896_));
 sg13g2_nor2_1 _1593_ (.A(net21),
    .B(_0828_),
    .Y(_0897_));
 sg13g2_nor2_1 _1594_ (.A(_0878_),
    .B(_0897_),
    .Y(_0898_));
 sg13g2_nor2_1 _1595_ (.A(net16),
    .B(net14),
    .Y(_0899_));
 sg13g2_a221oi_1 _1596_ (.B2(_0899_),
    .C1(net15),
    .B1(_0898_),
    .A1(_0895_),
    .Y(_0900_),
    .A2(_0896_));
 sg13g2_nand2_2 _1597_ (.Y(_0901_),
    .A(net78),
    .B(net15));
 sg13g2_nor2_1 _1598_ (.A(_0860_),
    .B(net22),
    .Y(_0902_));
 sg13g2_xnor2_1 _1599_ (.Y(_0903_),
    .A(_0824_),
    .B(_0842_));
 sg13g2_xor2_1 _1600_ (.B(_0058_),
    .A(_0056_),
    .X(_0904_));
 sg13g2_nand2_1 _1601_ (.Y(_0905_),
    .A(_0858_),
    .B(_0904_));
 sg13g2_o21ai_1 _1602_ (.B1(_0905_),
    .Y(_0906_),
    .A1(net24),
    .A2(_0903_));
 sg13g2_mux2_1 _1603_ (.A0(net16),
    .A1(_0902_),
    .S(_0906_),
    .X(_0907_));
 sg13g2_o21ai_1 _1604_ (.B1(net12),
    .Y(_0908_),
    .A1(_0901_),
    .A2(_0907_));
 sg13g2_nor2_1 _1605_ (.A(_0828_),
    .B(_0844_),
    .Y(_0909_));
 sg13g2_nand2b_1 _1606_ (.Y(_0910_),
    .B(_0844_),
    .A_N(net22));
 sg13g2_nand2_1 _1607_ (.Y(_0911_),
    .A(net72),
    .B(_0910_));
 sg13g2_nor2_2 _1608_ (.A(_0816_),
    .B(net13),
    .Y(_0912_));
 sg13g2_o21ai_1 _1609_ (.B1(_0912_),
    .Y(_0913_),
    .A1(_0909_),
    .A2(_0911_));
 sg13g2_o21ai_1 _1610_ (.B1(_0913_),
    .Y(_0001_),
    .A1(_0900_),
    .A2(_0908_));
 sg13g2_nand3_1 _1611_ (.B(net18),
    .C(net17),
    .A(net78),
    .Y(_0914_));
 sg13g2_nand3_1 _1612_ (.B(_0887_),
    .C(_0886_),
    .A(net21),
    .Y(_0915_));
 sg13g2_a21o_1 _1613_ (.A2(_0915_),
    .A1(_0914_),
    .B1(_0876_),
    .X(_0916_));
 sg13g2_nand3_1 _1614_ (.B(net14),
    .C(_0891_),
    .A(_0816_),
    .Y(_0917_));
 sg13g2_o21ai_1 _1615_ (.B1(net13),
    .Y(_0918_),
    .A1(_0886_),
    .A2(_0891_));
 sg13g2_inv_1 _1616_ (.Y(_0919_),
    .A(_0918_));
 sg13g2_a21oi_1 _1617_ (.A1(_0917_),
    .A2(_0919_),
    .Y(_0920_),
    .B1(_0901_));
 sg13g2_a21oi_1 _1618_ (.A1(net21),
    .A2(_0876_),
    .Y(_0921_),
    .B1(_0816_));
 sg13g2_o21ai_1 _1619_ (.B1(_0921_),
    .Y(_0922_),
    .A1(net14),
    .A2(_0878_));
 sg13g2_nand2b_1 _1620_ (.Y(_0923_),
    .B(_0835_),
    .A_N(_0828_));
 sg13g2_nor2_1 _1621_ (.A(_0923_),
    .B(net19),
    .Y(_0924_));
 sg13g2_or2_1 _1622_ (.X(_0925_),
    .B(_0844_),
    .A(_0835_));
 sg13g2_buf_1 _1623_ (.A(_0925_),
    .X(_0926_));
 sg13g2_nand2_1 _1624_ (.Y(_0927_),
    .A(_0889_),
    .B(_0926_));
 sg13g2_o21ai_1 _1625_ (.B1(_0857_),
    .Y(_0928_),
    .A1(_0924_),
    .A2(_0927_));
 sg13g2_a22oi_1 _1626_ (.Y(_0002_),
    .B1(_0922_),
    .B2(_0928_),
    .A2(_0920_),
    .A1(_0916_));
 sg13g2_nor2_1 _1627_ (.A(_0923_),
    .B(_0844_),
    .Y(_0929_));
 sg13g2_nor3_1 _1628_ (.A(_0901_),
    .B(_0902_),
    .C(_0929_),
    .Y(_0930_));
 sg13g2_nand2b_1 _1629_ (.Y(_0931_),
    .B(net12),
    .A_N(_0930_));
 sg13g2_nand2_1 _1630_ (.Y(_0932_),
    .A(_0860_),
    .B(net17));
 sg13g2_a21oi_1 _1631_ (.A1(net14),
    .A2(_0932_),
    .Y(_0933_),
    .B1(net16));
 sg13g2_nor2_1 _1632_ (.A(_0880_),
    .B(_0933_),
    .Y(_0934_));
 sg13g2_o21ai_1 _1633_ (.B1(_0922_),
    .Y(_0003_),
    .A1(_0931_),
    .A2(_0934_));
 sg13g2_nand2_1 _1634_ (.Y(_0935_),
    .A(net16),
    .B(net14));
 sg13g2_nor2_1 _1635_ (.A(_0878_),
    .B(_0935_),
    .Y(_0936_));
 sg13g2_nor2_1 _1636_ (.A(_0926_),
    .B(_0932_),
    .Y(_0937_));
 sg13g2_nor3_1 _1637_ (.A(_0880_),
    .B(_0936_),
    .C(_0937_),
    .Y(_0938_));
 sg13g2_inv_2 _1638_ (.Y(_0147_),
    .A(_0901_));
 sg13g2_nand2_1 _1639_ (.Y(_0939_),
    .A(_0923_),
    .B(_0147_));
 sg13g2_nor2_1 _1640_ (.A(_0861_),
    .B(_0926_),
    .Y(_0940_));
 sg13g2_o21ai_1 _1641_ (.B1(net12),
    .Y(_0941_),
    .A1(_0939_),
    .A2(_0940_));
 sg13g2_nor2_1 _1642_ (.A(net17),
    .B(_0910_),
    .Y(_0942_));
 sg13g2_nand2_1 _1643_ (.Y(_0943_),
    .A(_0912_),
    .B(_0942_));
 sg13g2_o21ai_1 _1644_ (.B1(_0943_),
    .Y(_0004_),
    .A1(_0938_),
    .A2(_0941_));
 sg13g2_nand2_1 _1645_ (.Y(_0944_),
    .A(net18),
    .B(net14));
 sg13g2_nand3b_1 _1646_ (.B(_0889_),
    .C(_0929_),
    .Y(_0945_),
    .A_N(net18));
 sg13g2_a21oi_1 _1647_ (.A1(_0944_),
    .A2(_0945_),
    .Y(_0946_),
    .B1(_0853_));
 sg13g2_o21ai_1 _1648_ (.B1(_0902_),
    .Y(_0947_),
    .A1(net18),
    .A2(_0871_));
 sg13g2_a21oi_1 _1649_ (.A1(_0891_),
    .A2(_0926_),
    .Y(_0948_),
    .B1(net21));
 sg13g2_nor2_1 _1650_ (.A(_0855_),
    .B(_0889_),
    .Y(_0949_));
 sg13g2_o21ai_1 _1651_ (.B1(_0949_),
    .Y(_0950_),
    .A1(_0924_),
    .A2(_0948_));
 sg13g2_nand3_1 _1652_ (.B(_0947_),
    .C(_0950_),
    .A(net72),
    .Y(_0951_));
 sg13g2_nor2_1 _1653_ (.A(net22),
    .B(net19),
    .Y(_0952_));
 sg13g2_nor3_1 _1654_ (.A(net18),
    .B(_0860_),
    .C(_0844_),
    .Y(_0953_));
 sg13g2_o21ai_1 _1655_ (.B1(_0889_),
    .Y(_0954_),
    .A1(_0952_),
    .A2(_0953_));
 sg13g2_a21oi_1 _1656_ (.A1(_0944_),
    .A2(_0954_),
    .Y(_0955_),
    .B1(_0887_));
 sg13g2_or3_1 _1657_ (.A(_0946_),
    .B(_0951_),
    .C(_0955_),
    .X(_0005_));
 sg13g2_a21oi_1 _1658_ (.A1(_0837_),
    .A2(_0901_),
    .Y(_0956_),
    .B1(net19));
 sg13g2_nor2_1 _1659_ (.A(net21),
    .B(_0956_),
    .Y(_0957_));
 sg13g2_and2_1 _1660_ (.A(net22),
    .B(net15),
    .X(_0958_));
 sg13g2_or2_1 _1661_ (.X(_0959_),
    .B(_0958_),
    .A(_0881_));
 sg13g2_nand2b_1 _1662_ (.Y(_0960_),
    .B(net78),
    .A_N(net18));
 sg13g2_a221oi_1 _1663_ (.B2(net17),
    .C1(_0960_),
    .B1(_0959_),
    .A1(net15),
    .Y(_0961_),
    .A2(_0942_));
 sg13g2_nand2b_1 _1664_ (.Y(_0962_),
    .B(_0961_),
    .A_N(_0871_));
 sg13g2_o21ai_1 _1665_ (.B1(_0943_),
    .Y(_0006_),
    .A1(_0957_),
    .A2(_0962_));
 sg13g2_nand2_1 _1666_ (.Y(_0963_),
    .A(_0862_),
    .B(_0845_));
 sg13g2_mux2_1 _1667_ (.A0(_0963_),
    .A1(net19),
    .S(_0890_),
    .X(_0964_));
 sg13g2_nand4_1 _1668_ (.B(_0857_),
    .C(_0872_),
    .A(_0861_),
    .Y(_0965_),
    .D(_0964_));
 sg13g2_o21ai_1 _1669_ (.B1(_0889_),
    .Y(_0966_),
    .A1(net17),
    .A2(_0952_));
 sg13g2_a21oi_1 _1670_ (.A1(net16),
    .A2(_0896_),
    .Y(_0967_),
    .B1(net13));
 sg13g2_nand3_1 _1671_ (.B(_0966_),
    .C(_0967_),
    .A(net12),
    .Y(_0968_));
 sg13g2_nand3_1 _1672_ (.B(_0912_),
    .C(_0952_),
    .A(net17),
    .Y(_0969_));
 sg13g2_nand3_1 _1673_ (.B(_0968_),
    .C(_0969_),
    .A(_0965_),
    .Y(_0007_));
 sg13g2_o21ai_1 _1674_ (.B1(_0897_),
    .Y(_0970_),
    .A1(_0899_),
    .A2(_0958_));
 sg13g2_nand2_1 _1675_ (.Y(_0971_),
    .A(net17),
    .B(_0844_));
 sg13g2_o21ai_1 _1676_ (.B1(_0971_),
    .Y(_0972_),
    .A1(net13),
    .A2(_0909_));
 sg13g2_nor2_1 _1677_ (.A(net21),
    .B(net22),
    .Y(_0973_));
 sg13g2_o21ai_1 _1678_ (.B1(net15),
    .Y(_0974_),
    .A1(net14),
    .A2(_0973_));
 sg13g2_o21ai_1 _1679_ (.B1(_0974_),
    .Y(_0975_),
    .A1(net15),
    .A2(_0972_));
 sg13g2_nand3_1 _1680_ (.B(_0970_),
    .C(_0975_),
    .A(net12),
    .Y(_0976_));
 sg13g2_o21ai_1 _1681_ (.B1(_0912_),
    .Y(_0977_),
    .A1(_0911_),
    .A2(_0929_));
 sg13g2_nand2_1 _1682_ (.Y(_0008_),
    .A(_0976_),
    .B(_0977_));
 sg13g2_or2_1 _1683_ (.X(_0978_),
    .B(_0966_),
    .A(net13));
 sg13g2_nand2_1 _1684_ (.Y(_0979_),
    .A(net16),
    .B(net19));
 sg13g2_nand4_1 _1685_ (.B(_0147_),
    .C(_0910_),
    .A(_0897_),
    .Y(_0980_),
    .D(_0979_));
 sg13g2_and2_1 _1686_ (.A(net12),
    .B(_0980_),
    .X(_0981_));
 sg13g2_nand3_1 _1687_ (.B(net17),
    .C(_0899_),
    .A(net52),
    .Y(_0982_));
 sg13g2_a22oi_1 _1688_ (.Y(_0009_),
    .B1(_0982_),
    .B2(_0912_),
    .A2(_0981_),
    .A1(_0978_));
 sg13g2_nand2_1 _1689_ (.Y(_0983_),
    .A(net72),
    .B(_0677_));
 sg13g2_nor2_1 _1690_ (.A(\counter.oled_driver.mc_exec.state_r[5] ),
    .B(\counter.oled_driver.mc_exec.spi_tx_trigger_out ),
    .Y(_0984_));
 sg13g2_nor2_1 _1691_ (.A(_0983_),
    .B(_0984_),
    .Y(_0010_));
 sg13g2_nor2_1 _1692_ (.A(\counter.oled_driver.state_r[4] ),
    .B(\counter.oled_driver.spi_deactivate_cs ),
    .Y(_0985_));
 sg13g2_nor2_1 _1693_ (.A(_0983_),
    .B(_0985_),
    .Y(_0013_));
 sg13g2_nand2b_1 _1694_ (.Y(_0986_),
    .B(net72),
    .A_N(net61));
 sg13g2_nor2_1 _1695_ (.A(net64),
    .B(\counter.oled_driver.write_stb_in ),
    .Y(_0987_));
 sg13g2_nor2_1 _1696_ (.A(_0986_),
    .B(_0987_),
    .Y(_0015_));
 sg13g2_nor2_1 _1697_ (.A(\counter.oled_driver.sync_stb_in ),
    .B(\counter.streamer.state_r[4] ),
    .Y(_0988_));
 sg13g2_nor2_1 _1698_ (.A(_0986_),
    .B(_0988_),
    .Y(_0014_));
 sg13g2_buf_1 _1699_ (.A(_0635_),
    .X(_0989_));
 sg13g2_nor2_1 _1700_ (.A(\counter.oled_driver.mc_exec.procedure_start_in ),
    .B(\counter.oled_driver.state_r[2] ),
    .Y(_0990_));
 sg13g2_nor3_1 _1701_ (.A(net51),
    .B(net47),
    .C(_0990_),
    .Y(_0012_));
 sg13g2_nand2b_1 _1702_ (.Y(_0991_),
    .B(_0701_),
    .A_N(net30));
 sg13g2_nor2_1 _1703_ (.A(\counter.oled_driver.spi_driver.state_r[1] ),
    .B(net56),
    .Y(_0992_));
 sg13g2_nor2_1 _1704_ (.A(_0991_),
    .B(_0992_),
    .Y(_0011_));
 sg13g2_buf_1 _1705_ (.A(net59),
    .X(_0993_));
 sg13g2_inv_1 _1706_ (.Y(_0073_),
    .A(_0993_));
 sg13g2_xor2_1 _1707_ (.B(\counter.cnt_x_digits[0] ),
    .A(_0721_),
    .X(_0098_));
 sg13g2_inv_2 _1708_ (.Y(_0994_),
    .A(\counter.cnt_x_digits[1] ));
 sg13g2_and2_1 _1709_ (.A(\counter.cnt_ref_enable ),
    .B(\counter.cnt_x_digits[0] ),
    .X(_0995_));
 sg13g2_buf_8 _1710_ (.A(_0995_),
    .X(_0996_));
 sg13g2_nand2_1 _1711_ (.Y(_0997_),
    .A(net71),
    .B(\counter.cnt_x_digits[0] ));
 sg13g2_nor2b_1 _1712_ (.A(\counter.cnt_x_digits[2] ),
    .B_N(\counter.cnt_x_digits[3] ),
    .Y(_0998_));
 sg13g2_or3_1 _1713_ (.A(\counter.cnt_x_digits[1] ),
    .B(_0997_),
    .C(_0998_),
    .X(_0999_));
 sg13g2_o21ai_1 _1714_ (.B1(_0999_),
    .Y(_0099_),
    .A1(_0994_),
    .A2(_0996_));
 sg13g2_nand2_1 _1715_ (.Y(_1000_),
    .A(\counter.cnt_x_digits[1] ),
    .B(_0996_));
 sg13g2_xnor2_1 _1716_ (.Y(_0100_),
    .A(\counter.cnt_x_digits[2] ),
    .B(_1000_));
 sg13g2_nor2b_1 _1717_ (.A(\counter.cnt_x_digits[3] ),
    .B_N(\counter.cnt_x_digits[2] ),
    .Y(_1001_));
 sg13g2_a21oi_1 _1718_ (.A1(_0996_),
    .A2(_1001_),
    .Y(_1002_),
    .B1(_0998_));
 sg13g2_nor2b_1 _1719_ (.A(\counter.cnt_x_digits[1] ),
    .B_N(\counter.cnt_x_digits[2] ),
    .Y(_1003_));
 sg13g2_o21ai_1 _1720_ (.B1(\counter.cnt_x_digits[3] ),
    .Y(_1004_),
    .A1(_0997_),
    .A2(_1003_));
 sg13g2_o21ai_1 _1721_ (.B1(_1004_),
    .Y(_0101_),
    .A1(_0994_),
    .A2(_1002_));
 sg13g2_and3_1 _1722_ (.X(_1005_),
    .A(_0994_),
    .B(_0996_),
    .C(_0998_));
 sg13g2_xor2_1 _1723_ (.B(_1005_),
    .A(\counter.cnt_x_digits[4] ),
    .X(_0102_));
 sg13g2_buf_2 _1724_ (.A(\counter.cnt_x_digits[5] ),
    .X(_1006_));
 sg13g2_nand4_1 _1725_ (.B(\counter.cnt_x_digits[4] ),
    .C(_0996_),
    .A(_0994_),
    .Y(_1007_),
    .D(_0998_));
 sg13g2_buf_2 _1726_ (.A(_1007_),
    .X(_1008_));
 sg13g2_nor2b_1 _1727_ (.A(\counter.cnt_x_digits[6] ),
    .B_N(\counter.cnt_x_digits[7] ),
    .Y(_1009_));
 sg13g2_nor3_1 _1728_ (.A(_1006_),
    .B(_1008_),
    .C(_1009_),
    .Y(_1010_));
 sg13g2_a21o_1 _1729_ (.A2(_1008_),
    .A1(_1006_),
    .B1(_1010_),
    .X(_0103_));
 sg13g2_nand3_1 _1730_ (.B(_1006_),
    .C(_1005_),
    .A(\counter.cnt_x_digits[4] ),
    .Y(_1011_));
 sg13g2_xnor2_1 _1731_ (.Y(_0104_),
    .A(\counter.cnt_x_digits[6] ),
    .B(_1011_));
 sg13g2_inv_1 _1732_ (.Y(_1012_),
    .A(\counter.cnt_x_digits[6] ));
 sg13g2_nor2_1 _1733_ (.A(_1006_),
    .B(_1012_),
    .Y(_1013_));
 sg13g2_o21ai_1 _1734_ (.B1(\counter.cnt_x_digits[7] ),
    .Y(_1014_),
    .A1(_1008_),
    .A2(_1013_));
 sg13g2_nor3_1 _1735_ (.A(_1012_),
    .B(\counter.cnt_x_digits[7] ),
    .C(_1008_),
    .Y(_1015_));
 sg13g2_o21ai_1 _1736_ (.B1(_1006_),
    .Y(_1016_),
    .A1(_1009_),
    .A2(_1015_));
 sg13g2_nand2_1 _1737_ (.Y(_0105_),
    .A(_1014_),
    .B(_1016_));
 sg13g2_buf_2 _1738_ (.A(\counter.cnt_x_digits[8] ),
    .X(_1017_));
 sg13g2_nand2_1 _1739_ (.Y(_1018_),
    .A(_1012_),
    .B(\counter.cnt_x_digits[7] ));
 sg13g2_nor3_2 _1740_ (.A(_1006_),
    .B(_1008_),
    .C(_1018_),
    .Y(_1019_));
 sg13g2_xor2_1 _1741_ (.B(_1019_),
    .A(_1017_),
    .X(_0106_));
 sg13g2_buf_2 _1742_ (.A(\counter.cnt_x_digits[9] ),
    .X(_1020_));
 sg13g2_nand2b_1 _1743_ (.Y(_1021_),
    .B(\counter.cnt_x_digits[11] ),
    .A_N(\counter.cnt_x_digits[10] ));
 sg13g2_nand3_1 _1744_ (.B(_1019_),
    .C(_1021_),
    .A(_1017_),
    .Y(_1022_));
 sg13g2_nand2_1 _1745_ (.Y(_1023_),
    .A(_1017_),
    .B(_1019_));
 sg13g2_nand2_1 _1746_ (.Y(_1024_),
    .A(_1020_),
    .B(_1023_));
 sg13g2_o21ai_1 _1747_ (.B1(_1024_),
    .Y(_0107_),
    .A1(_1020_),
    .A2(_1022_));
 sg13g2_nand3_1 _1748_ (.B(_1020_),
    .C(_1019_),
    .A(_1017_),
    .Y(_1025_));
 sg13g2_xnor2_1 _1749_ (.Y(_0108_),
    .A(\counter.cnt_x_digits[10] ),
    .B(_1025_));
 sg13g2_nor2b_1 _1750_ (.A(_1020_),
    .B_N(\counter.cnt_x_digits[10] ),
    .Y(_1026_));
 sg13g2_o21ai_1 _1751_ (.B1(\counter.cnt_x_digits[11] ),
    .Y(_1027_),
    .A1(_1023_),
    .A2(_1026_));
 sg13g2_nand2b_1 _1752_ (.Y(_1028_),
    .B(\counter.cnt_x_digits[10] ),
    .A_N(\counter.cnt_x_digits[11] ));
 sg13g2_o21ai_1 _1753_ (.B1(_1021_),
    .Y(_1029_),
    .A1(_1023_),
    .A2(_1028_));
 sg13g2_nand2_1 _1754_ (.Y(_1030_),
    .A(_1020_),
    .B(_1029_));
 sg13g2_nand2_1 _1755_ (.Y(_0109_),
    .A(_1027_),
    .B(_1030_));
 sg13g2_nor3_1 _1756_ (.A(_1020_),
    .B(_1023_),
    .C(_1021_),
    .Y(_1031_));
 sg13g2_xor2_1 _1757_ (.B(_1031_),
    .A(\counter.cnt_x_digits[12] ),
    .X(_0110_));
 sg13g2_nor3_1 _1758_ (.A(_1006_),
    .B(_1008_),
    .C(_1018_),
    .Y(_1032_));
 sg13g2_nor2_1 _1759_ (.A(_1020_),
    .B(_1021_),
    .Y(_1033_));
 sg13g2_nand4_1 _1760_ (.B(\counter.cnt_x_digits[12] ),
    .C(_1032_),
    .A(_1017_),
    .Y(_1034_),
    .D(_1033_));
 sg13g2_buf_2 _1761_ (.A(_1034_),
    .X(_1035_));
 sg13g2_buf_2 _1762_ (.A(\counter.cnt_x_digits[13] ),
    .X(_1036_));
 sg13g2_nand2b_1 _1763_ (.Y(_1037_),
    .B(\counter.cnt_x_digits[15] ),
    .A_N(\counter.cnt_x_digits[14] ));
 sg13g2_nand2b_1 _1764_ (.Y(_1038_),
    .B(_1037_),
    .A_N(_1036_));
 sg13g2_nand2_1 _1765_ (.Y(_1039_),
    .A(_1036_),
    .B(_1035_));
 sg13g2_o21ai_1 _1766_ (.B1(_1039_),
    .Y(_0111_),
    .A1(_1035_),
    .A2(_1038_));
 sg13g2_nand3_1 _1767_ (.B(_1036_),
    .C(_1031_),
    .A(\counter.cnt_x_digits[12] ),
    .Y(_1040_));
 sg13g2_xnor2_1 _1768_ (.Y(_0112_),
    .A(\counter.cnt_x_digits[14] ),
    .B(_1040_));
 sg13g2_nor2b_1 _1769_ (.A(_1036_),
    .B_N(\counter.cnt_x_digits[14] ),
    .Y(_1041_));
 sg13g2_o21ai_1 _1770_ (.B1(\counter.cnt_x_digits[15] ),
    .Y(_1042_),
    .A1(_1035_),
    .A2(_1041_));
 sg13g2_nand2b_1 _1771_ (.Y(_1043_),
    .B(\counter.cnt_x_digits[14] ),
    .A_N(\counter.cnt_x_digits[15] ));
 sg13g2_o21ai_1 _1772_ (.B1(_1037_),
    .Y(_1044_),
    .A1(_1035_),
    .A2(_1043_));
 sg13g2_nand2_1 _1773_ (.Y(_1045_),
    .A(_1036_),
    .B(_1044_));
 sg13g2_nand2_1 _1774_ (.Y(_0113_),
    .A(_1042_),
    .B(_1045_));
 sg13g2_inv_1 _1775_ (.Y(_1046_),
    .A(\counter.cnt_x_digits[16] ));
 sg13g2_nor3_1 _1776_ (.A(_1036_),
    .B(_1035_),
    .C(_1037_),
    .Y(_1047_));
 sg13g2_xnor2_1 _1777_ (.Y(_0114_),
    .A(_1046_),
    .B(_1047_));
 sg13g2_inv_1 _1778_ (.Y(_1048_),
    .A(\counter.cnt_x_digits[19] ));
 sg13g2_nor2_1 _1779_ (.A(\counter.cnt_x_digits[18] ),
    .B(_1048_),
    .Y(_1049_));
 sg13g2_nor2_1 _1780_ (.A(\counter.cnt_x_digits[17] ),
    .B(_1049_),
    .Y(_1050_));
 sg13g2_nor4_2 _1781_ (.A(_1036_),
    .B(_1046_),
    .C(_1035_),
    .Y(_1051_),
    .D(_1037_));
 sg13g2_mux2_1 _1782_ (.A0(\counter.cnt_x_digits[17] ),
    .A1(_1050_),
    .S(_1051_),
    .X(_0115_));
 sg13g2_nand2_1 _1783_ (.Y(_1052_),
    .A(\counter.cnt_x_digits[17] ),
    .B(_1051_));
 sg13g2_xnor2_1 _1784_ (.Y(_0116_),
    .A(\counter.cnt_x_digits[18] ),
    .B(_1052_));
 sg13g2_inv_1 _1785_ (.Y(_1053_),
    .A(\counter.cnt_x_digits[17] ));
 sg13g2_nor2b_1 _1786_ (.A(\counter.cnt_x_digits[19] ),
    .B_N(\counter.cnt_x_digits[18] ),
    .Y(_1054_));
 sg13g2_a21oi_1 _1787_ (.A1(_1051_),
    .A2(_1054_),
    .Y(_1055_),
    .B1(_1049_));
 sg13g2_nand2_1 _1788_ (.Y(_1056_),
    .A(_1053_),
    .B(\counter.cnt_x_digits[18] ));
 sg13g2_a21o_1 _1789_ (.A2(_1056_),
    .A1(_1051_),
    .B1(_1048_),
    .X(_1057_));
 sg13g2_o21ai_1 _1790_ (.B1(_1057_),
    .Y(_0117_),
    .A1(_1053_),
    .A2(_1055_));
 sg13g2_and3_1 _1791_ (.X(_1058_),
    .A(_1053_),
    .B(_1051_),
    .C(_1049_));
 sg13g2_xor2_1 _1792_ (.B(_1058_),
    .A(\counter.cnt_x_digits[20] ),
    .X(_0118_));
 sg13g2_inv_1 _1793_ (.Y(_1059_),
    .A(\counter.cnt_x_digits[21] ));
 sg13g2_and2_1 _1794_ (.A(\counter.cnt_x_digits[20] ),
    .B(_1058_),
    .X(_1060_));
 sg13g2_buf_8 _1795_ (.A(_1060_),
    .X(_1061_));
 sg13g2_inv_1 _1796_ (.Y(_1062_),
    .A(\counter.cnt_x_digits[22] ));
 sg13g2_nand2_1 _1797_ (.Y(_1063_),
    .A(_1062_),
    .B(\counter.cnt_x_digits[23] ));
 sg13g2_nand3_1 _1798_ (.B(_1061_),
    .C(_1063_),
    .A(_1059_),
    .Y(_1064_));
 sg13g2_o21ai_1 _1799_ (.B1(_1064_),
    .Y(_0119_),
    .A1(_1059_),
    .A2(_1061_));
 sg13g2_nand2_1 _1800_ (.Y(_1065_),
    .A(\counter.cnt_x_digits[21] ),
    .B(_1061_));
 sg13g2_xnor2_1 _1801_ (.Y(_0120_),
    .A(\counter.cnt_x_digits[22] ),
    .B(_1065_));
 sg13g2_o21ai_1 _1802_ (.B1(_1061_),
    .Y(_1066_),
    .A1(\counter.cnt_x_digits[21] ),
    .A2(_1062_));
 sg13g2_nand3b_1 _1803_ (.B(_1061_),
    .C(\counter.cnt_x_digits[22] ),
    .Y(_1067_),
    .A_N(\counter.cnt_x_digits[23] ));
 sg13g2_a21oi_1 _1804_ (.A1(_1063_),
    .A2(_1067_),
    .Y(_1068_),
    .B1(_1059_));
 sg13g2_a21o_1 _1805_ (.A2(_1066_),
    .A1(\counter.cnt_x_digits[23] ),
    .B1(_1068_),
    .X(_0121_));
 sg13g2_xnor2_1 _1806_ (.Y(_1069_),
    .A(\counter.counter_ref.digit_0.digit_out[0] ),
    .B(net71));
 sg13g2_nor2_1 _1807_ (.A(_0993_),
    .B(_1069_),
    .Y(_0074_));
 sg13g2_nand2_1 _1808_ (.Y(_1070_),
    .A(\counter.counter_ref.digit_0.digit_out[0] ),
    .B(net71));
 sg13g2_nor2b_1 _1809_ (.A(\counter.counter_ref.digit_0.digit_out[2] ),
    .B_N(\counter.counter_ref.digit_0.digit_out[3] ),
    .Y(_1071_));
 sg13g2_nor3_1 _1810_ (.A(_0727_),
    .B(_1071_),
    .C(_1070_),
    .Y(_1072_));
 sg13g2_a21oi_1 _1811_ (.A1(_0727_),
    .A2(_1070_),
    .Y(_1073_),
    .B1(_1072_));
 sg13g2_nor2_1 _1812_ (.A(net45),
    .B(_1073_),
    .Y(_0075_));
 sg13g2_inv_1 _1813_ (.Y(_1074_),
    .A(\counter.counter_ref.digit_0.digit_out[2] ));
 sg13g2_nand3_1 _1814_ (.B(_0727_),
    .C(net71),
    .A(\counter.counter_ref.digit_0.digit_out[0] ),
    .Y(_1075_));
 sg13g2_xnor2_1 _1815_ (.Y(_1076_),
    .A(_1074_),
    .B(_1075_));
 sg13g2_nor2_1 _1816_ (.A(net45),
    .B(_1076_),
    .Y(_0076_));
 sg13g2_nor2_1 _1817_ (.A(_0727_),
    .B(_1074_),
    .Y(_1077_));
 sg13g2_o21ai_1 _1818_ (.B1(\counter.counter_ref.digit_0.digit_out[3] ),
    .Y(_1078_),
    .A1(_1070_),
    .A2(_1077_));
 sg13g2_nor3_1 _1819_ (.A(_1074_),
    .B(\counter.counter_ref.digit_0.digit_out[3] ),
    .C(_1070_),
    .Y(_1079_));
 sg13g2_o21ai_1 _1820_ (.B1(_0727_),
    .Y(_1080_),
    .A1(_1071_),
    .A2(_1079_));
 sg13g2_buf_1 _1821_ (.A(net59),
    .X(_1081_));
 sg13g2_a21oi_1 _1822_ (.A1(_1078_),
    .A2(_1080_),
    .Y(_0077_),
    .B1(net44));
 sg13g2_nand2_1 _1823_ (.Y(_1082_),
    .A(net71),
    .B(_0729_));
 sg13g2_xor2_1 _1824_ (.B(_1082_),
    .A(\counter.counter_ref.digits_out[4] ),
    .X(_1083_));
 sg13g2_nor2_1 _1825_ (.A(net45),
    .B(_1083_),
    .Y(_0078_));
 sg13g2_nand3_1 _1826_ (.B(net71),
    .C(_0729_),
    .A(\counter.counter_ref.digits_out[4] ),
    .Y(_1084_));
 sg13g2_buf_1 _1827_ (.A(_1084_),
    .X(_1085_));
 sg13g2_nor3_1 _1828_ (.A(\counter.counter_ref.digits_out[5] ),
    .B(_0724_),
    .C(_1085_),
    .Y(_1086_));
 sg13g2_a21oi_1 _1829_ (.A1(\counter.counter_ref.digits_out[5] ),
    .A2(_1085_),
    .Y(_1087_),
    .B1(_1086_));
 sg13g2_nor2_1 _1830_ (.A(net45),
    .B(_1087_),
    .Y(_0079_));
 sg13g2_nor2_1 _1831_ (.A(_0723_),
    .B(_1085_),
    .Y(_1088_));
 sg13g2_xnor2_1 _1832_ (.Y(_1089_),
    .A(\counter.counter_ref.digits_out[6] ),
    .B(_1088_));
 sg13g2_nor2_1 _1833_ (.A(net45),
    .B(_1089_),
    .Y(_0080_));
 sg13g2_inv_1 _1834_ (.Y(_1090_),
    .A(\counter.counter_ref.digits_out[6] ));
 sg13g2_nor2_1 _1835_ (.A(\counter.counter_ref.digits_out[5] ),
    .B(_1090_),
    .Y(_1091_));
 sg13g2_o21ai_1 _1836_ (.B1(\counter.counter_ref.digits_out[7] ),
    .Y(_1092_),
    .A1(_1085_),
    .A2(_1091_));
 sg13g2_nor3_1 _1837_ (.A(_1090_),
    .B(\counter.counter_ref.digits_out[7] ),
    .C(_1085_),
    .Y(_1093_));
 sg13g2_o21ai_1 _1838_ (.B1(\counter.counter_ref.digits_out[5] ),
    .Y(_1094_),
    .A1(_0724_),
    .A2(_1093_));
 sg13g2_a21oi_1 _1839_ (.A1(_1092_),
    .A2(_1094_),
    .Y(_0081_),
    .B1(net44));
 sg13g2_nand2_1 _1840_ (.Y(_1095_),
    .A(_0723_),
    .B(_0724_));
 sg13g2_nor2_1 _1841_ (.A(_1085_),
    .B(_1095_),
    .Y(_1096_));
 sg13g2_xnor2_1 _1842_ (.Y(_1097_),
    .A(\counter.counter_ref.digits_out[8] ),
    .B(_1096_));
 sg13g2_nor2_1 _1843_ (.A(net45),
    .B(_1097_),
    .Y(_0082_));
 sg13g2_o21ai_1 _1844_ (.B1(\counter.counter_ref.digits_out[9] ),
    .Y(_1098_),
    .A1(_0725_),
    .A2(_1082_));
 sg13g2_nor2_1 _1845_ (.A(_0725_),
    .B(_1082_),
    .Y(_1099_));
 sg13g2_nand3b_1 _1846_ (.B(_0722_),
    .C(_1099_),
    .Y(_1100_),
    .A_N(\counter.counter_ref.digits_out[9] ));
 sg13g2_a21oi_1 _1847_ (.A1(_1098_),
    .A2(_1100_),
    .Y(_0083_),
    .B1(net59));
 sg13g2_nand2_1 _1848_ (.Y(_1101_),
    .A(\counter.counter_ref.digits_out[9] ),
    .B(_1099_));
 sg13g2_xor2_1 _1849_ (.B(_1101_),
    .A(\counter.counter_ref.digits_out[10] ),
    .X(_1102_));
 sg13g2_nor2_1 _1850_ (.A(net45),
    .B(_1102_),
    .Y(_0084_));
 sg13g2_and2_1 _1851_ (.A(net71),
    .B(_0731_),
    .X(_1103_));
 sg13g2_buf_1 _1852_ (.A(_1103_),
    .X(_1104_));
 sg13g2_nand3_1 _1853_ (.B(\counter.counter_ref.digits_out[10] ),
    .C(_1099_),
    .A(\counter.counter_ref.digits_out[9] ),
    .Y(_1105_));
 sg13g2_xor2_1 _1854_ (.B(_1105_),
    .A(\counter.counter_ref.digits_out[11] ),
    .X(_1106_));
 sg13g2_nor3_1 _1855_ (.A(net59),
    .B(_1104_),
    .C(_1106_),
    .Y(_0085_));
 sg13g2_xnor2_1 _1856_ (.Y(_1107_),
    .A(\counter.counter_ref.digits_out[12] ),
    .B(_1104_));
 sg13g2_nor2_1 _1857_ (.A(net45),
    .B(_1107_),
    .Y(_0086_));
 sg13g2_nand2_2 _1858_ (.Y(_1108_),
    .A(\counter.counter_ref.digits_out[12] ),
    .B(_1104_));
 sg13g2_nor3_1 _1859_ (.A(\counter.counter_ref.digits_out[13] ),
    .B(_0714_),
    .C(_1108_),
    .Y(_1109_));
 sg13g2_a21oi_1 _1860_ (.A1(\counter.counter_ref.digits_out[13] ),
    .A2(_1108_),
    .Y(_1110_),
    .B1(_1109_));
 sg13g2_nor2_1 _1861_ (.A(_1081_),
    .B(_1110_),
    .Y(_0087_));
 sg13g2_nor2_1 _1862_ (.A(_0713_),
    .B(_1108_),
    .Y(_1111_));
 sg13g2_xnor2_1 _1863_ (.Y(_1112_),
    .A(\counter.counter_ref.digits_out[14] ),
    .B(_1111_));
 sg13g2_nor2_1 _1864_ (.A(net44),
    .B(_1112_),
    .Y(_0088_));
 sg13g2_inv_1 _1865_ (.Y(_1113_),
    .A(\counter.counter_ref.digits_out[14] ));
 sg13g2_nor2_1 _1866_ (.A(\counter.counter_ref.digits_out[13] ),
    .B(_1113_),
    .Y(_1114_));
 sg13g2_o21ai_1 _1867_ (.B1(\counter.counter_ref.digits_out[15] ),
    .Y(_1115_),
    .A1(_1108_),
    .A2(_1114_));
 sg13g2_nor3_1 _1868_ (.A(_1113_),
    .B(\counter.counter_ref.digits_out[15] ),
    .C(_1108_),
    .Y(_1116_));
 sg13g2_o21ai_1 _1869_ (.B1(\counter.counter_ref.digits_out[13] ),
    .Y(_1117_),
    .A1(_0714_),
    .A2(_1116_));
 sg13g2_a21oi_1 _1870_ (.A1(_1115_),
    .A2(_1117_),
    .Y(_0089_),
    .B1(net59));
 sg13g2_and4_1 _1871_ (.A(\counter.counter_ref.digits_out[12] ),
    .B(_0713_),
    .C(_0714_),
    .D(_1104_),
    .X(_1118_));
 sg13g2_xnor2_1 _1872_ (.Y(_1119_),
    .A(\counter.counter_ref.digits_out[16] ),
    .B(_1118_));
 sg13g2_nor2_1 _1873_ (.A(_1081_),
    .B(_1119_),
    .Y(_0090_));
 sg13g2_nand2b_1 _1874_ (.Y(_1120_),
    .B(_1104_),
    .A_N(_0715_));
 sg13g2_nand2_1 _1875_ (.Y(_1121_),
    .A(_0712_),
    .B(_1120_));
 sg13g2_nor2_1 _1876_ (.A(_0715_),
    .B(_0732_),
    .Y(_1122_));
 sg13g2_nand3b_1 _1877_ (.B(_0719_),
    .C(_1122_),
    .Y(_1123_),
    .A_N(_0712_));
 sg13g2_a21oi_1 _1878_ (.A1(_1121_),
    .A2(_1123_),
    .Y(_0091_),
    .B1(net59));
 sg13g2_nand2_1 _1879_ (.Y(_1124_),
    .A(_0712_),
    .B(_1122_));
 sg13g2_xnor2_1 _1880_ (.Y(_1125_),
    .A(_0718_),
    .B(_1124_));
 sg13g2_nor2_1 _1881_ (.A(net44),
    .B(_1125_),
    .Y(_0092_));
 sg13g2_o21ai_1 _1882_ (.B1(_1122_),
    .Y(_1126_),
    .A1(_0712_),
    .A2(_0718_));
 sg13g2_nand2b_1 _1883_ (.Y(_1127_),
    .B(\counter.counter_ref.digits_out[18] ),
    .A_N(\counter.counter_ref.digits_out[19] ));
 sg13g2_o21ai_1 _1884_ (.B1(_0719_),
    .Y(_1128_),
    .A1(_1120_),
    .A2(_1127_));
 sg13g2_a22oi_1 _1885_ (.Y(_1129_),
    .B1(_1128_),
    .B2(_0712_),
    .A2(_1126_),
    .A1(\counter.counter_ref.digits_out[19] ));
 sg13g2_nor2_1 _1886_ (.A(net44),
    .B(_1129_),
    .Y(_0093_));
 sg13g2_xnor2_1 _1887_ (.Y(_1130_),
    .A(\counter.counter_ref.digits_out[20] ),
    .B(_0733_));
 sg13g2_nor2_1 _1888_ (.A(net44),
    .B(_1130_),
    .Y(_0094_));
 sg13g2_nand2_1 _1889_ (.Y(_1131_),
    .A(\counter.counter_ref.digits_out[20] ),
    .B(_0733_));
 sg13g2_nor3_1 _1890_ (.A(_0708_),
    .B(_0709_),
    .C(_1131_),
    .Y(_1132_));
 sg13g2_a21oi_1 _1891_ (.A1(_0708_),
    .A2(_1131_),
    .Y(_1133_),
    .B1(_1132_));
 sg13g2_nor2_1 _1892_ (.A(net44),
    .B(_1133_),
    .Y(_0095_));
 sg13g2_inv_1 _1893_ (.Y(_1134_),
    .A(\counter.counter_ref.digits_out[22] ));
 sg13g2_nand3_1 _1894_ (.B(_0708_),
    .C(_0733_),
    .A(\counter.counter_ref.digits_out[20] ),
    .Y(_1135_));
 sg13g2_xnor2_1 _1895_ (.Y(_1136_),
    .A(_1134_),
    .B(_1135_));
 sg13g2_nor2_1 _1896_ (.A(net44),
    .B(_1136_),
    .Y(_0096_));
 sg13g2_nor2_1 _1897_ (.A(_0708_),
    .B(_1134_),
    .Y(_1137_));
 sg13g2_o21ai_1 _1898_ (.B1(\counter.counter_ref.digits_out[23] ),
    .Y(_1138_),
    .A1(_1131_),
    .A2(_1137_));
 sg13g2_nor3_1 _1899_ (.A(_1134_),
    .B(\counter.counter_ref.digits_out[23] ),
    .C(_1131_),
    .Y(_1139_));
 sg13g2_o21ai_1 _1900_ (.B1(_0708_),
    .Y(_1140_),
    .A1(_0709_),
    .A2(_1139_));
 sg13g2_a21oi_1 _1901_ (.A1(_1138_),
    .A2(_1140_),
    .Y(_0097_),
    .B1(_0717_));
 sg13g2_nand2b_1 _1902_ (.Y(_1141_),
    .B(_0749_),
    .A_N(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ));
 sg13g2_nand2_1 _1903_ (.Y(_1142_),
    .A(net58),
    .B(_0072_));
 sg13g2_a21oi_1 _1904_ (.A1(_0742_),
    .A2(_1141_),
    .Y(_0160_),
    .B1(_1142_));
 sg13g2_xnor2_1 _1905_ (.Y(_1143_),
    .A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ),
    .B(_0741_));
 sg13g2_nor2_1 _1906_ (.A(net48),
    .B(_1143_),
    .Y(_0161_));
 sg13g2_nand2_1 _1907_ (.Y(_1144_),
    .A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ),
    .B(_0741_));
 sg13g2_xor2_1 _1908_ (.B(_1144_),
    .A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ),
    .X(_1145_));
 sg13g2_nor2_1 _1909_ (.A(net48),
    .B(_1145_),
    .Y(_0162_));
 sg13g2_o21ai_1 _1910_ (.B1(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ),
    .Y(_1146_),
    .A1(_0741_),
    .A2(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ));
 sg13g2_nor2b_1 _1911_ (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ),
    .B_N(_1146_),
    .Y(_1147_));
 sg13g2_and4_1 _1912_ (.A(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ),
    .B(_0741_),
    .C(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ),
    .D(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ),
    .X(_1148_));
 sg13g2_a21oi_1 _1913_ (.A1(_0741_),
    .A2(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ),
    .Y(_1149_),
    .B1(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ));
 sg13g2_nor4_1 _1914_ (.A(net63),
    .B(_1147_),
    .C(_1148_),
    .D(_1149_),
    .Y(_0163_));
 sg13g2_nand3_1 _1915_ (.B(_0758_),
    .C(_0672_),
    .A(\counter.streamer.graphical_decoder.index_y_in[0] ),
    .Y(_1150_));
 sg13g2_o21ai_1 _1916_ (.B1(_0707_),
    .Y(_1151_),
    .A1(net64),
    .A2(_0706_));
 sg13g2_a21o_1 _1917_ (.A2(_1150_),
    .A1(net64),
    .B1(_1151_),
    .X(_1152_));
 sg13g2_buf_1 _1918_ (.A(_1152_),
    .X(_1153_));
 sg13g2_a21oi_2 _1919_ (.B1(net29),
    .Y(_1154_),
    .A2(_0756_),
    .A1(net64));
 sg13g2_nand2b_1 _1920_ (.Y(_1155_),
    .B(net78),
    .A_N(_1154_));
 sg13g2_nand2_1 _1921_ (.Y(_1156_),
    .A(net68),
    .B(_0754_));
 sg13g2_xnor2_1 _1922_ (.Y(_1157_),
    .A(_0061_),
    .B(_1156_));
 sg13g2_nand2_1 _1923_ (.Y(_1158_),
    .A(_0752_),
    .B(net29));
 sg13g2_o21ai_1 _1924_ (.B1(_1158_),
    .Y(_1159_),
    .A1(net29),
    .A2(_1157_));
 sg13g2_nand2b_1 _1925_ (.Y(_1160_),
    .B(_1159_),
    .A_N(_1155_));
 sg13g2_nand2_1 _1926_ (.Y(_1161_),
    .A(_0753_),
    .B(_0752_));
 sg13g2_nor3_1 _1927_ (.A(_0062_),
    .B(net29),
    .C(_1161_),
    .Y(_1162_));
 sg13g2_xnor2_1 _1928_ (.Y(_1163_),
    .A(\counter.streamer.graphical_decoder.index_x_in[3] ),
    .B(_1162_));
 sg13g2_or2_1 _1929_ (.X(_1164_),
    .B(_1163_),
    .A(_1155_));
 sg13g2_nand4_1 _1930_ (.B(_0754_),
    .C(\counter.streamer.graphical_decoder.index_x_in[3] ),
    .A(net68),
    .Y(_1165_),
    .D(_0752_));
 sg13g2_xnor2_1 _1931_ (.Y(_1166_),
    .A(_0060_),
    .B(_1165_));
 sg13g2_nor2_1 _1932_ (.A(net29),
    .B(_1166_),
    .Y(_0211_));
 sg13g2_a21oi_1 _1933_ (.A1(\counter.streamer.graphical_decoder.index_x_in[4] ),
    .A2(net29),
    .Y(_0212_),
    .B1(_0211_));
 sg13g2_nor2_1 _1934_ (.A(_1155_),
    .B(_0212_),
    .Y(_0208_));
 sg13g2_a21oi_1 _1935_ (.A1(_1160_),
    .A2(_1164_),
    .Y(_0200_),
    .B1(_0208_));
 sg13g2_xnor2_1 _1936_ (.Y(_0213_),
    .A(_0754_),
    .B(net29));
 sg13g2_inv_1 _1937_ (.Y(_0214_),
    .A(net68));
 sg13g2_nand2_1 _1938_ (.Y(_0215_),
    .A(_0214_),
    .B(_0754_));
 sg13g2_inv_1 _1939_ (.Y(_0216_),
    .A(_0754_));
 sg13g2_nand2_1 _1940_ (.Y(_0217_),
    .A(net68),
    .B(_0216_));
 sg13g2_o21ai_1 _1941_ (.B1(_0217_),
    .Y(_0218_),
    .A1(net29),
    .A2(_0215_));
 sg13g2_a22oi_1 _1942_ (.Y(_0219_),
    .B1(_0218_),
    .B2(_0767_),
    .A2(_1153_),
    .A1(net68));
 sg13g2_nor2_1 _1943_ (.A(_0635_),
    .B(_0219_),
    .Y(_0205_));
 sg13g2_inv_1 _1944_ (.Y(_0206_),
    .A(_1160_));
 sg13g2_o21ai_1 _1945_ (.B1(_0206_),
    .Y(_0220_),
    .A1(_0213_),
    .A2(_0205_));
 sg13g2_and2_1 _1946_ (.A(_0206_),
    .B(_0205_),
    .X(_0221_));
 sg13g2_nor2b_1 _1947_ (.A(_1163_),
    .B_N(_0213_),
    .Y(_0222_));
 sg13g2_a221oi_1 _1948_ (.B2(_0222_),
    .C1(_0208_),
    .B1(_0221_),
    .A1(_1164_),
    .Y(_0201_),
    .A2(_0220_));
 sg13g2_nand2_1 _1949_ (.Y(_0223_),
    .A(_1163_),
    .B(_0221_));
 sg13g2_inv_1 _1950_ (.Y(_0207_),
    .A(_1164_));
 sg13g2_nand2b_1 _1951_ (.Y(_0224_),
    .B(_0207_),
    .A_N(_0221_));
 sg13g2_a21oi_1 _1952_ (.A1(_0223_),
    .A2(_0224_),
    .Y(_0203_),
    .B1(_0208_));
 sg13g2_nor2b_1 _1953_ (.A(_1155_),
    .B_N(_0213_),
    .Y(_0204_));
 sg13g2_a21o_1 _1954_ (.A2(_0204_),
    .A1(_0205_),
    .B1(_0220_),
    .X(_0225_));
 sg13g2_and2_1 _1955_ (.A(_0203_),
    .B(_0225_),
    .X(_0202_));
 sg13g2_nor2b_1 _1956_ (.A(_0040_),
    .B_N(_0656_),
    .Y(_0226_));
 sg13g2_or3_1 _1957_ (.A(_0804_),
    .B(_0652_),
    .C(_0226_),
    .X(_0227_));
 sg13g2_buf_1 _1958_ (.A(_0055_),
    .X(_0228_));
 sg13g2_nor2_1 _1959_ (.A(\counter.oled_driver.mc_exec.state_r[0] ),
    .B(net76),
    .Y(_0229_));
 sg13g2_nand2_1 _1960_ (.Y(_0230_),
    .A(_0228_),
    .B(_0229_));
 sg13g2_nand3_1 _1961_ (.B(_0227_),
    .C(_0230_),
    .A(_0699_),
    .Y(_0231_));
 sg13g2_buf_2 _1962_ (.A(_0231_),
    .X(_0232_));
 sg13g2_buf_1 _1963_ (.A(_0232_),
    .X(_0233_));
 sg13g2_inv_1 _1964_ (.Y(_0234_),
    .A(\counter.oled_driver.mc_exec.state_r[6] ));
 sg13g2_nor3_1 _1965_ (.A(\counter.oled_driver.mc_exec.delay_cnt[0] ),
    .B(_0234_),
    .C(net23),
    .Y(_0235_));
 sg13g2_a21oi_1 _1966_ (.A1(\counter.oled_driver.mc_exec.delay_cnt[0] ),
    .A2(net23),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_nor2_1 _1967_ (.A(net48),
    .B(_0236_),
    .Y(_0122_));
 sg13g2_nor2_1 _1968_ (.A(net76),
    .B(\counter.oled_driver.mc_exec.state_r[6] ),
    .Y(_0237_));
 sg13g2_nor2_1 _1969_ (.A(_0228_),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_o21ai_1 _1970_ (.B1(net78),
    .Y(_0239_),
    .A1(_0232_),
    .A2(_0238_));
 sg13g2_buf_1 _1971_ (.A(_0239_),
    .X(_0240_));
 sg13g2_nand2_1 _1972_ (.Y(_0241_),
    .A(_0681_),
    .B(_0682_));
 sg13g2_or3_1 _1973_ (.A(\counter.oled_driver.mc_exec.delay_cnt[5] ),
    .B(_0241_),
    .C(_0232_),
    .X(_0242_));
 sg13g2_or2_1 _1974_ (.X(_0243_),
    .B(_0242_),
    .A(\counter.oled_driver.mc_exec.delay_cnt[6] ));
 sg13g2_buf_2 _1975_ (.A(_0243_),
    .X(_0244_));
 sg13g2_nor3_1 _1976_ (.A(\counter.oled_driver.mc_exec.delay_cnt[7] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[8] ),
    .C(_0244_),
    .Y(_0245_));
 sg13g2_nand2b_1 _1977_ (.Y(_0246_),
    .B(_0245_),
    .A_N(\counter.oled_driver.mc_exec.delay_cnt[9] ));
 sg13g2_xor2_1 _1978_ (.B(_0246_),
    .A(\counter.oled_driver.mc_exec.delay_cnt[10] ),
    .X(_0247_));
 sg13g2_nor2_1 _1979_ (.A(_0240_),
    .B(_0247_),
    .Y(_0123_));
 sg13g2_xor2_1 _1980_ (.B(_0685_),
    .A(\counter.oled_driver.mc_exec.delay_cnt[11] ),
    .X(_0248_));
 sg13g2_nand2b_1 _1981_ (.Y(_0249_),
    .B(_0664_),
    .A_N(_0804_));
 sg13g2_o21ai_1 _1982_ (.B1(_0249_),
    .Y(_0250_),
    .A1(_0228_),
    .A2(_0248_));
 sg13g2_nor2_1 _1983_ (.A(_0232_),
    .B(_0237_),
    .Y(_0251_));
 sg13g2_a22oi_1 _1984_ (.Y(_0252_),
    .B1(_0250_),
    .B2(_0251_),
    .A2(net23),
    .A1(\counter.oled_driver.mc_exec.delay_cnt[11] ));
 sg13g2_nor2_1 _1985_ (.A(net48),
    .B(_0252_),
    .Y(_0124_));
 sg13g2_buf_1 _1986_ (.A(net63),
    .X(_0253_));
 sg13g2_o21ai_1 _1987_ (.B1(\counter.oled_driver.mc_exec.delay_cnt[12] ),
    .Y(_0254_),
    .A1(\counter.oled_driver.mc_exec.delay_cnt[11] ),
    .A2(_0685_));
 sg13g2_nor2b_1 _1988_ (.A(_0686_),
    .B_N(_0254_),
    .Y(_0255_));
 sg13g2_nor2_1 _1989_ (.A(_0804_),
    .B(_0642_),
    .Y(_0256_));
 sg13g2_nand2_1 _1990_ (.Y(_0257_),
    .A(_0666_),
    .B(_0256_));
 sg13g2_o21ai_1 _1991_ (.B1(_0257_),
    .Y(_0258_),
    .A1(_0228_),
    .A2(_0255_));
 sg13g2_a22oi_1 _1992_ (.Y(_0259_),
    .B1(_0251_),
    .B2(_0258_),
    .A2(net23),
    .A1(\counter.oled_driver.mc_exec.delay_cnt[12] ));
 sg13g2_nor2_1 _1993_ (.A(net43),
    .B(_0259_),
    .Y(_0125_));
 sg13g2_a22oi_1 _1994_ (.Y(_0260_),
    .B1(_0238_),
    .B2(_0687_),
    .A2(_0694_),
    .A1(net74));
 sg13g2_nor2b_1 _1995_ (.A(_0686_),
    .B_N(_0238_),
    .Y(_0261_));
 sg13g2_o21ai_1 _1996_ (.B1(\counter.oled_driver.mc_exec.delay_cnt[13] ),
    .Y(_0262_),
    .A1(_0232_),
    .A2(_0261_));
 sg13g2_o21ai_1 _1997_ (.B1(_0262_),
    .Y(_0263_),
    .A1(net23),
    .A2(_0260_));
 sg13g2_and2_1 _1998_ (.A(net58),
    .B(_0263_),
    .X(_0126_));
 sg13g2_nand2b_1 _1999_ (.Y(_0264_),
    .B(\counter.oled_driver.mc_exec.delay_cnt[14] ),
    .A_N(_0687_));
 sg13g2_a21oi_1 _2000_ (.A1(_0688_),
    .A2(_0264_),
    .Y(_0265_),
    .B1(_0228_));
 sg13g2_nand2_1 _2001_ (.Y(_0266_),
    .A(net73),
    .B(net37));
 sg13g2_nor2b_1 _2002_ (.A(_0265_),
    .B_N(_0266_),
    .Y(_0267_));
 sg13g2_a21oi_1 _2003_ (.A1(\counter.oled_driver.mc_exec.state_r[6] ),
    .A2(_0265_),
    .Y(_0268_),
    .B1(net76));
 sg13g2_nor3_1 _2004_ (.A(_0232_),
    .B(_0267_),
    .C(_0268_),
    .Y(_0269_));
 sg13g2_a21oi_1 _2005_ (.A1(\counter.oled_driver.mc_exec.delay_cnt[14] ),
    .A2(net23),
    .Y(_0270_),
    .B1(_0269_));
 sg13g2_nor2_1 _2006_ (.A(net43),
    .B(_0270_),
    .Y(_0127_));
 sg13g2_xor2_1 _2007_ (.B(_0688_),
    .A(\counter.oled_driver.mc_exec.delay_cnt[15] ),
    .X(_0271_));
 sg13g2_nand2_1 _2008_ (.Y(_0272_),
    .A(_0653_),
    .B(_0256_));
 sg13g2_o21ai_1 _2009_ (.B1(_0272_),
    .Y(_0273_),
    .A1(_0228_),
    .A2(_0271_));
 sg13g2_a22oi_1 _2010_ (.Y(_0274_),
    .B1(_0251_),
    .B2(_0273_),
    .A2(net23),
    .A1(\counter.oled_driver.mc_exec.delay_cnt[15] ));
 sg13g2_nor2_1 _2011_ (.A(net43),
    .B(_0274_),
    .Y(_0128_));
 sg13g2_nor2b_1 _2012_ (.A(\counter.oled_driver.mc_exec.delay_cnt[16] ),
    .B_N(_0233_),
    .Y(_0275_));
 sg13g2_xnor2_1 _2013_ (.Y(_0276_),
    .A(_0052_),
    .B(_0689_));
 sg13g2_a221oi_1 _2014_ (.B2(_0276_),
    .C1(_0233_),
    .B1(_0238_),
    .A1(net75),
    .Y(_0277_),
    .A2(_0694_));
 sg13g2_nor3_1 _2015_ (.A(net63),
    .B(_0275_),
    .C(_0277_),
    .Y(_0129_));
 sg13g2_nor2_1 _2016_ (.A(\counter.oled_driver.mc_exec.delay_cnt[0] ),
    .B(_0232_),
    .Y(_0278_));
 sg13g2_xnor2_1 _2017_ (.Y(_0279_),
    .A(\counter.oled_driver.mc_exec.delay_cnt[1] ),
    .B(_0278_));
 sg13g2_nor2_1 _2018_ (.A(net20),
    .B(_0279_),
    .Y(_0130_));
 sg13g2_nand2b_1 _2019_ (.Y(_0280_),
    .B(_0278_),
    .A_N(\counter.oled_driver.mc_exec.delay_cnt[1] ));
 sg13g2_xor2_1 _2020_ (.B(_0280_),
    .A(\counter.oled_driver.mc_exec.delay_cnt[2] ),
    .X(_0281_));
 sg13g2_nor2_1 _2021_ (.A(net20),
    .B(_0281_),
    .Y(_0131_));
 sg13g2_or3_1 _2022_ (.A(\counter.oled_driver.mc_exec.delay_cnt[3] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[2] ),
    .C(_0280_),
    .X(_0282_));
 sg13g2_o21ai_1 _2023_ (.B1(\counter.oled_driver.mc_exec.delay_cnt[3] ),
    .Y(_0283_),
    .A1(\counter.oled_driver.mc_exec.delay_cnt[2] ),
    .A2(_0280_));
 sg13g2_a21oi_1 _2024_ (.A1(_0282_),
    .A2(_0283_),
    .Y(_0132_),
    .B1(net20));
 sg13g2_xnor2_1 _2025_ (.Y(_0284_),
    .A(_0681_),
    .B(_0282_));
 sg13g2_nor2_1 _2026_ (.A(net20),
    .B(_0284_),
    .Y(_0133_));
 sg13g2_o21ai_1 _2027_ (.B1(\counter.oled_driver.mc_exec.delay_cnt[5] ),
    .Y(_0285_),
    .A1(_0241_),
    .A2(net23));
 sg13g2_a21oi_1 _2028_ (.A1(_0242_),
    .A2(_0285_),
    .Y(_0134_),
    .B1(net20));
 sg13g2_nand2_1 _2029_ (.Y(_0286_),
    .A(\counter.oled_driver.mc_exec.delay_cnt[6] ),
    .B(_0242_));
 sg13g2_a21oi_1 _2030_ (.A1(_0244_),
    .A2(_0286_),
    .Y(_0135_),
    .B1(net20));
 sg13g2_xor2_1 _2031_ (.B(_0244_),
    .A(\counter.oled_driver.mc_exec.delay_cnt[7] ),
    .X(_0287_));
 sg13g2_nor2_1 _2032_ (.A(net20),
    .B(_0287_),
    .Y(_0136_));
 sg13g2_or3_1 _2033_ (.A(\counter.oled_driver.mc_exec.delay_cnt[7] ),
    .B(\counter.oled_driver.mc_exec.delay_cnt[8] ),
    .C(_0244_),
    .X(_0288_));
 sg13g2_o21ai_1 _2034_ (.B1(\counter.oled_driver.mc_exec.delay_cnt[8] ),
    .Y(_0289_),
    .A1(\counter.oled_driver.mc_exec.delay_cnt[7] ),
    .A2(_0244_));
 sg13g2_a21oi_1 _2035_ (.A1(_0288_),
    .A2(_0289_),
    .Y(_0137_),
    .B1(net20));
 sg13g2_nand2b_1 _2036_ (.Y(_0290_),
    .B(\counter.oled_driver.mc_exec.delay_cnt[9] ),
    .A_N(_0245_));
 sg13g2_a21oi_1 _2037_ (.A1(_0246_),
    .A2(_0290_),
    .Y(_0138_),
    .B1(_0240_));
 sg13g2_nand2_1 _2038_ (.Y(_0291_),
    .A(_0660_),
    .B(net37));
 sg13g2_nand2_1 _2039_ (.Y(_0292_),
    .A(net75),
    .B(_0665_));
 sg13g2_nor2_1 _2040_ (.A(_0695_),
    .B(_0292_),
    .Y(_0293_));
 sg13g2_nand3_1 _2041_ (.B(net73),
    .C(_0293_),
    .A(net74),
    .Y(_0294_));
 sg13g2_nand2_1 _2042_ (.Y(_0295_),
    .A(\counter.oled_driver.mc_exec.oled_dc_out ),
    .B(_0294_));
 sg13g2_o21ai_1 _2043_ (.B1(_0295_),
    .Y(_0296_),
    .A1(_0291_),
    .A2(_0294_));
 sg13g2_and2_1 _2044_ (.A(net58),
    .B(_0296_),
    .X(_0139_));
 sg13g2_nor3_1 _2045_ (.A(_0667_),
    .B(net73),
    .C(_0292_),
    .Y(_0297_));
 sg13g2_o21ai_1 _2046_ (.B1(_0691_),
    .Y(_0298_),
    .A1(_0656_),
    .A2(_0297_));
 sg13g2_nand3_1 _2047_ (.B(_0256_),
    .C(_0298_),
    .A(_0042_),
    .Y(_0299_));
 sg13g2_o21ai_1 _2048_ (.B1(_0649_),
    .Y(_0300_),
    .A1(_0652_),
    .A2(_0226_));
 sg13g2_nand3b_1 _2049_ (.B(_0299_),
    .C(_0300_),
    .Y(_0301_),
    .A_N(_0229_));
 sg13g2_nor2_1 _2050_ (.A(_0249_),
    .B(_0301_),
    .Y(_0302_));
 sg13g2_a21oi_1 _2051_ (.A1(\counter.oled_driver.mc_exec.oled_rstn_out ),
    .A2(_0301_),
    .Y(_0303_),
    .B1(_0302_));
 sg13g2_nor2_1 _2052_ (.A(net43),
    .B(_0303_),
    .Y(_0140_));
 sg13g2_nand2_1 _2053_ (.Y(_0304_),
    .A(net74),
    .B(_0293_));
 sg13g2_nor3_1 _2054_ (.A(net73),
    .B(_0291_),
    .C(_0304_),
    .Y(_0305_));
 sg13g2_o21ai_1 _2055_ (.B1(\counter.oled_driver.mc_exec.oled_vbatn_out ),
    .Y(_0306_),
    .A1(_0668_),
    .A2(_0304_));
 sg13g2_nand3b_1 _2056_ (.B(net58),
    .C(_0306_),
    .Y(_0141_),
    .A_N(_0305_));
 sg13g2_nand2_1 _2057_ (.Y(_0307_),
    .A(_0668_),
    .B(_0293_));
 sg13g2_nor3_1 _2058_ (.A(_0667_),
    .B(_0291_),
    .C(_0307_),
    .Y(_0308_));
 sg13g2_o21ai_1 _2059_ (.B1(\counter.oled_driver.mc_exec.oled_vcdn_out ),
    .Y(_0309_),
    .A1(net74),
    .A2(_0307_));
 sg13g2_nand3b_1 _2060_ (.B(_0735_),
    .C(_0309_),
    .Y(_0142_),
    .A_N(_0308_));
 sg13g2_o21ai_1 _2061_ (.B1(net52),
    .Y(_0310_),
    .A1(_0817_),
    .A2(_0814_));
 sg13g2_a21oi_1 _2062_ (.A1(_0814_),
    .A2(_0842_),
    .Y(_0143_),
    .B1(_0310_));
 sg13g2_nand2_1 _2063_ (.Y(_0311_),
    .A(_0814_),
    .B(_0833_));
 sg13g2_nand2_1 _2064_ (.Y(_0312_),
    .A(_0789_),
    .B(net24));
 sg13g2_a21oi_1 _2065_ (.A1(_0311_),
    .A2(_0312_),
    .Y(_0144_),
    .B1(net46));
 sg13g2_o21ai_1 _2066_ (.B1(net52),
    .Y(_0313_),
    .A1(_0639_),
    .A2(_0814_));
 sg13g2_a21oi_1 _2067_ (.A1(_0814_),
    .A2(_0824_),
    .Y(_0145_),
    .B1(_0313_));
 sg13g2_inv_1 _2068_ (.Y(_0314_),
    .A(\counter.oled_driver.mc_exec.microcode_rom.address[3] ));
 sg13g2_mux2_1 _2069_ (.A0(_0851_),
    .A1(_0314_),
    .S(net24),
    .X(_0315_));
 sg13g2_nor2_1 _2070_ (.A(net43),
    .B(_0315_),
    .Y(_0146_));
 sg13g2_o21ai_1 _2071_ (.B1(net61),
    .Y(_0316_),
    .A1(\counter.oled_driver.sync_stb_in ),
    .A2(\counter.oled_driver.mc_exec.procedure_offset_in[0] ));
 sg13g2_nand2_1 _2072_ (.Y(_0317_),
    .A(_0740_),
    .B(\counter.oled_driver.mc_exec.procedure_offset_in[0] ));
 sg13g2_a21oi_1 _2073_ (.A1(_0316_),
    .A2(_0317_),
    .Y(_0149_),
    .B1(_0779_));
 sg13g2_nand2_1 _2074_ (.Y(_0318_),
    .A(net1),
    .B(net77));
 sg13g2_nand2b_1 _2075_ (.Y(_0319_),
    .B(\counter.oled_driver.write_stb_in ),
    .A_N(\counter.oled_driver.sync_stb_in ));
 sg13g2_nor3_1 _2076_ (.A(_0672_),
    .B(\counter.oled_driver.state_r[4] ),
    .C(\counter.oled_driver.state_r[0] ),
    .Y(_0320_));
 sg13g2_a221oi_1 _2077_ (.B2(_0672_),
    .C1(_0320_),
    .B1(_0319_),
    .A1(\counter.oled_driver.state_r[4] ),
    .Y(_0321_),
    .A2(_0318_));
 sg13g2_buf_1 _2078_ (.A(_0321_),
    .X(_0322_));
 sg13g2_inv_1 _2079_ (.Y(_0323_),
    .A(_0322_));
 sg13g2_nor2_1 _2080_ (.A(_0760_),
    .B(net65),
    .Y(_0324_));
 sg13g2_mux2_1 _2081_ (.A0(\counter.streamer.digits_r[1] ),
    .A1(\counter.streamer.digits_r[9] ),
    .S(net54),
    .X(_0325_));
 sg13g2_nand2_1 _2082_ (.Y(_0326_),
    .A(_0324_),
    .B(_0325_));
 sg13g2_nor2b_1 _2083_ (.A(net54),
    .B_N(\counter.streamer.digit_cnt_r[2] ),
    .Y(_0327_));
 sg13g2_mux2_1 _2084_ (.A0(\counter.streamer.digits_r[17] ),
    .A1(\counter.streamer.digits_r[21] ),
    .S(net66),
    .X(_0328_));
 sg13g2_mux2_1 _2085_ (.A0(\counter.streamer.digits_r[5] ),
    .A1(\counter.streamer.digits_r[13] ),
    .S(net54),
    .X(_0329_));
 sg13g2_nor2b_1 _2086_ (.A(net65),
    .B_N(net66),
    .Y(_0330_));
 sg13g2_a22oi_1 _2087_ (.Y(_0331_),
    .B1(_0329_),
    .B2(_0330_),
    .A2(_0328_),
    .A1(_0327_));
 sg13g2_and2_1 _2088_ (.A(_0326_),
    .B(_0331_),
    .X(_0332_));
 sg13g2_buf_8 _2089_ (.A(_0332_),
    .X(_0333_));
 sg13g2_mux2_1 _2090_ (.A0(\counter.streamer.digits_r[2] ),
    .A1(\counter.streamer.digits_r[18] ),
    .S(\counter.streamer.digit_cnt_r[2] ),
    .X(_0334_));
 sg13g2_nor2b_1 _2091_ (.A(net65),
    .B_N(\counter.streamer.digits_r[10] ),
    .Y(_0335_));
 sg13g2_mux2_1 _2092_ (.A0(\counter.streamer.digits_r[6] ),
    .A1(\counter.streamer.digits_r[22] ),
    .S(\counter.streamer.digit_cnt_r[2] ),
    .X(_0336_));
 sg13g2_nor2b_1 _2093_ (.A(net65),
    .B_N(\counter.streamer.digits_r[14] ),
    .Y(_0337_));
 sg13g2_mux4_1 _2094_ (.S0(net54),
    .A0(_0334_),
    .A1(_0335_),
    .A2(_0336_),
    .A3(_0337_),
    .S1(net66),
    .X(_0338_));
 sg13g2_buf_1 _2095_ (.A(_0338_),
    .X(_0339_));
 sg13g2_nand2b_1 _2096_ (.Y(_0340_),
    .B(_0760_),
    .A_N(net65));
 sg13g2_mux2_1 _2097_ (.A0(_0069_),
    .A1(_0071_),
    .S(_0761_),
    .X(_0341_));
 sg13g2_nor2_1 _2098_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sg13g2_mux2_1 _2099_ (.A0(_0068_),
    .A1(_0070_),
    .S(_0761_),
    .X(_0343_));
 sg13g2_nor2b_1 _2100_ (.A(_0343_),
    .B_N(_0324_),
    .Y(_0344_));
 sg13g2_mux2_1 _2101_ (.A0(\counter.streamer.digits_r[19] ),
    .A1(\counter.streamer.digits_r[23] ),
    .S(\counter.streamer.digit_cnt_r[0] ),
    .X(_0345_));
 sg13g2_and3_1 _2102_ (.X(_0346_),
    .A(net65),
    .B(_0067_),
    .C(_0345_));
 sg13g2_or3_1 _2103_ (.A(_0342_),
    .B(_0344_),
    .C(_0346_),
    .X(_0347_));
 sg13g2_buf_1 _2104_ (.A(_0347_),
    .X(_0348_));
 sg13g2_buf_8 _2105_ (.A(net28),
    .X(_0349_));
 sg13g2_mux2_1 _2106_ (.A0(\counter.streamer.digits_r[0] ),
    .A1(\counter.streamer.digits_r[8] ),
    .S(_0761_),
    .X(_0350_));
 sg13g2_nand2_1 _2107_ (.Y(_0351_),
    .A(_0324_),
    .B(_0350_));
 sg13g2_mux2_1 _2108_ (.A0(\counter.streamer.digits_r[16] ),
    .A1(\counter.streamer.digits_r[20] ),
    .S(\counter.streamer.digit_cnt_r[0] ),
    .X(_0352_));
 sg13g2_mux2_1 _2109_ (.A0(\counter.streamer.digits_r[4] ),
    .A1(\counter.streamer.digits_r[12] ),
    .S(_0761_),
    .X(_0353_));
 sg13g2_a22oi_1 _2110_ (.Y(_0354_),
    .B1(_0353_),
    .B2(_0330_),
    .A2(_0352_),
    .A1(_0327_));
 sg13g2_and2_1 _2111_ (.A(_0351_),
    .B(_0354_),
    .X(_0355_));
 sg13g2_buf_2 _2112_ (.A(_0355_),
    .X(_0356_));
 sg13g2_nand3_1 _2113_ (.B(net26),
    .C(_0356_),
    .A(net31),
    .Y(_0357_));
 sg13g2_o21ai_1 _2114_ (.B1(_0357_),
    .Y(_0358_),
    .A1(net31),
    .A2(net26));
 sg13g2_nor2_1 _2115_ (.A(net26),
    .B(net27),
    .Y(_0359_));
 sg13g2_inv_1 _2116_ (.Y(_0360_),
    .A(_0338_));
 sg13g2_nor2_1 _2117_ (.A(_0360_),
    .B(_0356_),
    .Y(_0361_));
 sg13g2_o21ai_1 _2118_ (.B1(_0752_),
    .Y(_0362_),
    .A1(net68),
    .A2(_0754_));
 sg13g2_inv_1 _2119_ (.Y(_0363_),
    .A(\counter.streamer.graphical_decoder.index_x_in[4] ));
 sg13g2_a21oi_1 _2120_ (.A1(_0751_),
    .A2(_0362_),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_a221oi_1 _2121_ (.B2(_0361_),
    .C1(_0364_),
    .B1(_0359_),
    .A1(net27),
    .Y(_0365_),
    .A2(_0358_));
 sg13g2_inv_1 _2122_ (.Y(_0366_),
    .A(_0758_));
 sg13g2_buf_1 _2123_ (.A(_0366_),
    .X(_0367_));
 sg13g2_nor2_1 _2124_ (.A(net67),
    .B(net42),
    .Y(_0368_));
 sg13g2_and2_1 _2125_ (.A(_0365_),
    .B(_0368_),
    .X(_0369_));
 sg13g2_inv_1 _2126_ (.Y(_0370_),
    .A(_0066_));
 sg13g2_and2_1 _2127_ (.A(_0672_),
    .B(_0322_),
    .X(_0371_));
 sg13g2_buf_1 _2128_ (.A(_0371_),
    .X(_0372_));
 sg13g2_and2_1 _2129_ (.A(_0370_),
    .B(net25),
    .X(_0373_));
 sg13g2_a22oi_1 _2130_ (.Y(_0374_),
    .B1(_0369_),
    .B2(_0373_),
    .A2(_0323_),
    .A1(\counter.oled_driver.spi_data[0] ));
 sg13g2_buf_1 _2131_ (.A(_0043_),
    .X(_0375_));
 sg13g2_nand2_2 _2132_ (.Y(_0376_),
    .A(_0326_),
    .B(_0331_));
 sg13g2_nor3_1 _2133_ (.A(_0360_),
    .B(net28),
    .C(_0376_),
    .Y(_0377_));
 sg13g2_o21ai_1 _2134_ (.B1(_0758_),
    .Y(_0378_),
    .A1(_0375_),
    .A2(_0377_));
 sg13g2_nand3_1 _2135_ (.B(_0326_),
    .C(_0331_),
    .A(_0758_),
    .Y(_0379_));
 sg13g2_a221oi_1 _2136_ (.B2(net28),
    .C1(_0356_),
    .B1(_0379_),
    .A1(net31),
    .Y(_0380_),
    .A2(net27));
 sg13g2_nand2b_1 _2137_ (.Y(_0381_),
    .B(_0060_),
    .A_N(_0754_));
 sg13g2_a21oi_1 _2138_ (.A1(_0062_),
    .A2(_0381_),
    .Y(_0382_),
    .B1(_0214_));
 sg13g2_o21ai_1 _2139_ (.B1(\counter.streamer.graphical_decoder.index_x_in[3] ),
    .Y(_0383_),
    .A1(_0752_),
    .A2(_0382_));
 sg13g2_and2_1 _2140_ (.A(_0363_),
    .B(_0383_),
    .X(_0384_));
 sg13g2_nor2b_1 _2141_ (.A(_0380_),
    .B_N(_0384_),
    .Y(_0385_));
 sg13g2_nand2_2 _2142_ (.Y(_0386_),
    .A(_0351_),
    .B(_0354_));
 sg13g2_and4_1 _2143_ (.A(net31),
    .B(net28),
    .C(net27),
    .D(_0386_),
    .X(_0387_));
 sg13g2_nor3_1 _2144_ (.A(net31),
    .B(_0348_),
    .C(net27),
    .Y(_0388_));
 sg13g2_o21ai_1 _2145_ (.B1(_0375_),
    .Y(_0389_),
    .A1(_0387_),
    .A2(_0388_));
 sg13g2_nand3_1 _2146_ (.B(_0385_),
    .C(_0389_),
    .A(_0378_),
    .Y(_0390_));
 sg13g2_nand4_1 _2147_ (.B(_0338_),
    .C(_0333_),
    .A(_0375_),
    .Y(_0391_),
    .D(_0386_));
 sg13g2_nor2_1 _2148_ (.A(_0375_),
    .B(_0338_),
    .Y(_0392_));
 sg13g2_nand3_1 _2149_ (.B(_0356_),
    .C(_0392_),
    .A(_0376_),
    .Y(_0393_));
 sg13g2_a21o_1 _2150_ (.A2(_0393_),
    .A1(_0391_),
    .B1(net28),
    .X(_0394_));
 sg13g2_buf_2 _2151_ (.A(_0394_),
    .X(_0395_));
 sg13g2_and2_1 _2152_ (.A(net28),
    .B(_0356_),
    .X(_0396_));
 sg13g2_and3_1 _2153_ (.X(_0397_),
    .A(_0338_),
    .B(_0351_),
    .C(_0354_));
 sg13g2_a21o_1 _2154_ (.A2(_0386_),
    .A1(net28),
    .B1(_0397_),
    .X(_0398_));
 sg13g2_nor4_1 _2155_ (.A(_0375_),
    .B(_0342_),
    .C(_0344_),
    .D(_0346_),
    .Y(_0399_));
 sg13g2_nor3_1 _2156_ (.A(net27),
    .B(_0392_),
    .C(_0399_),
    .Y(_0400_));
 sg13g2_a221oi_1 _2157_ (.B2(_0400_),
    .C1(_0384_),
    .B1(_0398_),
    .A1(_0339_),
    .Y(_0401_),
    .A2(_0396_));
 sg13g2_buf_2 _2158_ (.A(_0401_),
    .X(_0402_));
 sg13g2_nand2_1 _2159_ (.Y(_0403_),
    .A(_0395_),
    .B(_0402_));
 sg13g2_a221oi_1 _2160_ (.B2(_0354_),
    .C1(net26),
    .B1(_0351_),
    .A1(net31),
    .Y(_0404_),
    .A2(net27));
 sg13g2_nand3_1 _2161_ (.B(_0363_),
    .C(_0383_),
    .A(_0366_),
    .Y(_0405_));
 sg13g2_nor4_1 _2162_ (.A(_0387_),
    .B(_0388_),
    .C(_0404_),
    .D(_0405_),
    .Y(_0406_));
 sg13g2_or4_1 _2163_ (.A(_0360_),
    .B(net28),
    .C(_0376_),
    .D(_0356_),
    .X(_0407_));
 sg13g2_o21ai_1 _2164_ (.B1(_0397_),
    .Y(_0408_),
    .A1(_0349_),
    .A2(_0376_));
 sg13g2_inv_1 _2165_ (.Y(_0409_),
    .A(_0375_));
 sg13g2_a21oi_1 _2166_ (.A1(_0363_),
    .A2(_0383_),
    .Y(_0410_),
    .B1(_0409_));
 sg13g2_nand3_1 _2167_ (.B(_0376_),
    .C(_0386_),
    .A(_0349_),
    .Y(_0411_));
 sg13g2_and4_1 _2168_ (.A(_0407_),
    .B(_0408_),
    .C(_0410_),
    .D(_0411_),
    .X(_0412_));
 sg13g2_o21ai_1 _2169_ (.B1(_0757_),
    .Y(_0413_),
    .A1(_0406_),
    .A2(_0412_));
 sg13g2_inv_1 _2170_ (.Y(_0414_),
    .A(_0044_));
 sg13g2_or3_1 _2171_ (.A(_0414_),
    .B(_0406_),
    .C(_0412_),
    .X(_0415_));
 sg13g2_a22oi_1 _2172_ (.Y(_0416_),
    .B1(_0413_),
    .B2(_0415_),
    .A2(_0403_),
    .A1(_0390_));
 sg13g2_buf_1 _2173_ (.A(_0416_),
    .X(_0417_));
 sg13g2_xnor2_1 _2174_ (.Y(_0418_),
    .A(net42),
    .B(net11));
 sg13g2_inv_1 _2175_ (.Y(_0419_),
    .A(_0061_));
 sg13g2_inv_1 _2176_ (.Y(_0420_),
    .A(_0045_));
 sg13g2_and4_1 _2177_ (.A(_0419_),
    .B(_0420_),
    .C(_0395_),
    .D(_0402_),
    .X(_0421_));
 sg13g2_and4_1 _2178_ (.A(_0061_),
    .B(_0045_),
    .C(_0395_),
    .D(_0402_),
    .X(_0422_));
 sg13g2_nor2_1 _2179_ (.A(_0753_),
    .B(_0061_),
    .Y(_0423_));
 sg13g2_and4_1 _2180_ (.A(_0378_),
    .B(_0385_),
    .C(_0389_),
    .D(_0423_),
    .X(_0424_));
 sg13g2_nor2_1 _2181_ (.A(_0214_),
    .B(_0419_),
    .Y(_0425_));
 sg13g2_and4_1 _2182_ (.A(_0378_),
    .B(_0385_),
    .C(_0389_),
    .D(_0425_),
    .X(_0426_));
 sg13g2_or4_1 _2183_ (.A(_0421_),
    .B(_0422_),
    .C(_0424_),
    .D(_0426_),
    .X(_0427_));
 sg13g2_buf_8 _2184_ (.A(_0427_),
    .X(_0428_));
 sg13g2_nand3_1 _2185_ (.B(_0418_),
    .C(_0428_),
    .A(net25),
    .Y(_0429_));
 sg13g2_a21oi_1 _2186_ (.A1(_0374_),
    .A2(_0429_),
    .Y(_0150_),
    .B1(_0779_));
 sg13g2_nand3_1 _2187_ (.B(_0395_),
    .C(_0402_),
    .A(_0062_),
    .Y(_0430_));
 sg13g2_nand4_1 _2188_ (.B(_0378_),
    .C(_0385_),
    .A(net68),
    .Y(_0431_),
    .D(_0389_));
 sg13g2_a21o_1 _2189_ (.A2(_0430_),
    .A1(_0216_),
    .B1(_0431_),
    .X(_0432_));
 sg13g2_or2_1 _2190_ (.X(_0433_),
    .B(_0430_),
    .A(_0420_));
 sg13g2_a21oi_1 _2191_ (.A1(_0432_),
    .A2(_0433_),
    .Y(_0434_),
    .B1(_0419_));
 sg13g2_nor2b_1 _2192_ (.A(net11),
    .B_N(_0428_),
    .Y(_0435_));
 sg13g2_o21ai_1 _2193_ (.B1(net55),
    .Y(_0436_),
    .A1(_0434_),
    .A2(_0435_));
 sg13g2_inv_1 _2194_ (.Y(_0437_),
    .A(_0046_));
 sg13g2_xnor2_1 _2195_ (.Y(_0438_),
    .A(net26),
    .B(_0356_));
 sg13g2_nand3b_1 _2196_ (.B(_0386_),
    .C(_0360_),
    .Y(_0439_),
    .A_N(net26));
 sg13g2_o21ai_1 _2197_ (.B1(_0439_),
    .Y(_0440_),
    .A1(_0360_),
    .A2(_0438_));
 sg13g2_nor3_1 _2198_ (.A(_0757_),
    .B(_0759_),
    .C(_0364_),
    .Y(_0441_));
 sg13g2_o21ai_1 _2199_ (.B1(_0441_),
    .Y(_0442_),
    .A1(_0339_),
    .A2(_0411_));
 sg13g2_a21oi_2 _2200_ (.B1(_0442_),
    .Y(_0443_),
    .A2(_0440_),
    .A1(_0333_));
 sg13g2_nor2b_1 _2201_ (.A(_0322_),
    .B_N(\counter.oled_driver.spi_data[1] ),
    .Y(_0444_));
 sg13g2_a221oi_1 _2202_ (.B2(\counter.streamer.graphical_decoder.pattern_adg[1] ),
    .C1(_0444_),
    .B1(_0443_),
    .A1(_0437_),
    .Y(_0445_),
    .A2(_0369_));
 sg13g2_nand3_1 _2203_ (.B(net11),
    .C(_0428_),
    .A(net42),
    .Y(_0446_));
 sg13g2_and2_1 _2204_ (.A(_0445_),
    .B(_0446_),
    .X(_0447_));
 sg13g2_o21ai_1 _2205_ (.B1(net52),
    .Y(_0448_),
    .A1(net25),
    .A2(_0444_));
 sg13g2_a21oi_1 _2206_ (.A1(_0436_),
    .A2(_0447_),
    .Y(_0151_),
    .B1(_0448_));
 sg13g2_nor2b_1 _2207_ (.A(_0322_),
    .B_N(\counter.oled_driver.spi_data[2] ),
    .Y(_0449_));
 sg13g2_a21oi_1 _2208_ (.A1(_0370_),
    .A2(_0443_),
    .Y(_0450_),
    .B1(_0449_));
 sg13g2_o21ai_1 _2209_ (.B1(_0428_),
    .Y(_0451_),
    .A1(net55),
    .A2(net11));
 sg13g2_nand4_1 _2210_ (.B(_0420_),
    .C(_0395_),
    .A(_0062_),
    .Y(_0452_),
    .D(_0402_));
 sg13g2_o21ai_1 _2211_ (.B1(_0452_),
    .Y(_0453_),
    .A1(_0215_),
    .A2(_0390_));
 sg13g2_nand3_1 _2212_ (.B(net11),
    .C(_0453_),
    .A(net55),
    .Y(_0454_));
 sg13g2_nand2b_1 _2213_ (.Y(_0455_),
    .B(_0454_),
    .A_N(_0451_));
 sg13g2_o21ai_1 _2214_ (.B1(net52),
    .Y(_0456_),
    .A1(net25),
    .A2(_0449_));
 sg13g2_a21oi_1 _2215_ (.A1(_0450_),
    .A2(_0455_),
    .Y(_0152_),
    .B1(_0456_));
 sg13g2_nand2_1 _2216_ (.Y(_0457_),
    .A(net11),
    .B(_0428_));
 sg13g2_nand3b_1 _2217_ (.B(net55),
    .C(\counter.streamer.graphical_decoder.index_y_in[0] ),
    .Y(_0458_),
    .A_N(_0364_));
 sg13g2_nand2_1 _2218_ (.Y(_0459_),
    .A(net31),
    .B(_0386_));
 sg13g2_nand3_1 _2219_ (.B(net26),
    .C(_0356_),
    .A(_0360_),
    .Y(_0460_));
 sg13g2_a21oi_1 _2220_ (.A1(_0459_),
    .A2(_0460_),
    .Y(_0461_),
    .B1(net27));
 sg13g2_nor2_1 _2221_ (.A(net31),
    .B(_0386_),
    .Y(_0462_));
 sg13g2_nor4_1 _2222_ (.A(net26),
    .B(_0376_),
    .C(_0361_),
    .D(_0462_),
    .Y(_0463_));
 sg13g2_nor3_2 _2223_ (.A(_0458_),
    .B(_0461_),
    .C(_0463_),
    .Y(_0464_));
 sg13g2_nor2b_1 _2224_ (.A(_0322_),
    .B_N(\counter.oled_driver.spi_data[3] ),
    .Y(_0465_));
 sg13g2_a221oi_1 _2225_ (.B2(\counter.streamer.graphical_decoder.pattern_adg[4] ),
    .C1(_0465_),
    .B1(_0464_),
    .A1(_0437_),
    .Y(_0466_),
    .A2(_0443_));
 sg13g2_and2_1 _2226_ (.A(_0457_),
    .B(_0466_),
    .X(_0467_));
 sg13g2_a21o_1 _2227_ (.A2(_0433_),
    .A1(_0432_),
    .B1(_0419_),
    .X(_0468_));
 sg13g2_nand2b_1 _2228_ (.Y(_0469_),
    .B(_0428_),
    .A_N(_0453_));
 sg13g2_mux2_1 _2229_ (.A0(_0468_),
    .A1(_0469_),
    .S(_0759_),
    .X(_0470_));
 sg13g2_o21ai_1 _2230_ (.B1(net52),
    .Y(_0471_),
    .A1(net25),
    .A2(_0465_));
 sg13g2_a21oi_1 _2231_ (.A1(_0467_),
    .A2(_0470_),
    .Y(_0153_),
    .B1(_0471_));
 sg13g2_nor2b_1 _2232_ (.A(_0322_),
    .B_N(\counter.oled_driver.spi_data[4] ),
    .Y(_0472_));
 sg13g2_a221oi_1 _2233_ (.B2(\counter.streamer.graphical_decoder.pattern_adg[3] ),
    .C1(_0472_),
    .B1(_0464_),
    .A1(\counter.streamer.graphical_decoder.pattern_adg[4] ),
    .Y(_0473_),
    .A2(_0443_));
 sg13g2_and2_1 _2234_ (.A(_0457_),
    .B(_0473_),
    .X(_0474_));
 sg13g2_mux2_1 _2235_ (.A0(_0468_),
    .A1(_0469_),
    .S(net42),
    .X(_0475_));
 sg13g2_o21ai_1 _2236_ (.B1(net52),
    .Y(_0476_),
    .A1(_0372_),
    .A2(_0472_));
 sg13g2_a21oi_1 _2237_ (.A1(_0474_),
    .A2(_0475_),
    .Y(_0154_),
    .B1(_0476_));
 sg13g2_nor2_1 _2238_ (.A(_0214_),
    .B(_0062_),
    .Y(_0477_));
 sg13g2_nor4_1 _2239_ (.A(\counter.streamer.graphical_decoder.index_x_in[3] ),
    .B(_0752_),
    .C(_0363_),
    .D(_0477_),
    .Y(_0478_));
 sg13g2_nand2b_1 _2240_ (.Y(_0479_),
    .B(net54),
    .A_N(_0060_));
 sg13g2_nor4_2 _2241_ (.A(_0340_),
    .B(_0458_),
    .C(_0478_),
    .Y(_0480_),
    .D(_0479_));
 sg13g2_a221oi_1 _2242_ (.B2(_0370_),
    .C1(_0480_),
    .B1(_0464_),
    .A1(\counter.oled_driver.spi_data[5] ),
    .Y(_0481_),
    .A2(_0323_));
 sg13g2_o21ai_1 _2243_ (.B1(_0428_),
    .Y(_0482_),
    .A1(_0367_),
    .A2(net11));
 sg13g2_nand3_1 _2244_ (.B(_0417_),
    .C(_0453_),
    .A(_0367_),
    .Y(_0483_));
 sg13g2_nand2b_1 _2245_ (.Y(_0484_),
    .B(_0483_),
    .A_N(_0482_));
 sg13g2_nor2b_1 _2246_ (.A(_0322_),
    .B_N(\counter.oled_driver.spi_data[5] ),
    .Y(_0485_));
 sg13g2_o21ai_1 _2247_ (.B1(_0875_),
    .Y(_0486_),
    .A1(net25),
    .A2(_0485_));
 sg13g2_a21oi_1 _2248_ (.A1(_0481_),
    .A2(_0484_),
    .Y(_0155_),
    .B1(_0486_));
 sg13g2_a21oi_1 _2249_ (.A1(\counter.oled_driver.spi_data[6] ),
    .A2(_0323_),
    .Y(_0487_),
    .B1(net25));
 sg13g2_a221oi_1 _2250_ (.B2(\counter.streamer.graphical_decoder.pattern_adg[1] ),
    .C1(_0480_),
    .B1(_0464_),
    .A1(\counter.oled_driver.spi_data[6] ),
    .Y(_0488_),
    .A2(_0323_));
 sg13g2_nand3_1 _2251_ (.B(\counter.streamer.graphical_decoder.pattern_adg[3] ),
    .C(_0365_),
    .A(net67),
    .Y(_0489_));
 sg13g2_nand3_1 _2252_ (.B(_0488_),
    .C(_0489_),
    .A(net42),
    .Y(_0490_));
 sg13g2_nor3_1 _2253_ (.A(_0434_),
    .B(_0435_),
    .C(_0490_),
    .Y(_0491_));
 sg13g2_and3_1 _2254_ (.X(_0492_),
    .A(net55),
    .B(_0457_),
    .C(_0488_));
 sg13g2_nor4_1 _2255_ (.A(_0636_),
    .B(_0487_),
    .C(_0491_),
    .D(_0492_),
    .Y(_0156_));
 sg13g2_nand2b_1 _2256_ (.Y(_0493_),
    .B(_0428_),
    .A_N(net11));
 sg13g2_and2_1 _2257_ (.A(net67),
    .B(\counter.streamer.graphical_decoder.pattern_adg[2] ),
    .X(_0494_));
 sg13g2_a21oi_1 _2258_ (.A1(_0365_),
    .A2(_0494_),
    .Y(_0495_),
    .B1(net55));
 sg13g2_nor2_1 _2259_ (.A(net42),
    .B(_0480_),
    .Y(_0496_));
 sg13g2_nand2_1 _2260_ (.Y(_0497_),
    .A(_0701_),
    .B(net25));
 sg13g2_a221oi_1 _2261_ (.B2(_0457_),
    .C1(_0497_),
    .B1(_0496_),
    .A1(_0493_),
    .Y(_0498_),
    .A2(_0495_));
 sg13g2_nand3_1 _2262_ (.B(\counter.oled_driver.spi_data[7] ),
    .C(_0323_),
    .A(_0875_),
    .Y(_0499_));
 sg13g2_nand2b_1 _2263_ (.Y(_0157_),
    .B(_0499_),
    .A_N(_0498_));
 sg13g2_o21ai_1 _2264_ (.B1(net36),
    .Y(_0500_),
    .A1(_0677_),
    .A2(_0747_));
 sg13g2_nand2_1 _2265_ (.Y(_0501_),
    .A(\counter.oled_csn_out ),
    .B(_0500_));
 sg13g2_nand3_1 _2266_ (.B(\counter.oled_driver.spi_driver.deactivate_cs_r ),
    .C(_0770_),
    .A(\counter.oled_driver.spi_driver.state_r[1] ),
    .Y(_0502_));
 sg13g2_nor2b_1 _2267_ (.A(\counter.oled_driver.spi_driver.state_r[1] ),
    .B_N(\counter.oled_csn_out ),
    .Y(_0503_));
 sg13g2_and4_1 _2268_ (.A(_0634_),
    .B(\counter.oled_driver.spi_driver.state_r[1] ),
    .C(\counter.oled_driver.spi_driver.deactivate_cs_r ),
    .D(_0743_),
    .X(_0504_));
 sg13g2_o21ai_1 _2269_ (.B1(_0677_),
    .Y(_0505_),
    .A1(_0503_),
    .A2(_0504_));
 sg13g2_nand4_1 _2270_ (.B(_0501_),
    .C(_0502_),
    .A(_0735_),
    .Y(_0158_),
    .D(_0505_));
 sg13g2_nand4_1 _2271_ (.B(_0799_),
    .C(\counter.oled_driver.mc_exec.spi_tx_trigger_out ),
    .A(_0643_),
    .Y(_0506_),
    .D(net36));
 sg13g2_a21oi_1 _2272_ (.A1(_0041_),
    .A2(net37),
    .Y(_0507_),
    .B1(_0506_));
 sg13g2_a21oi_1 _2273_ (.A1(net77),
    .A2(_0770_),
    .Y(_0508_),
    .B1(\counter.oled_driver.spi_driver.deactivate_cs_r ));
 sg13g2_nor3_1 _2274_ (.A(net63),
    .B(_0507_),
    .C(_0508_),
    .Y(_0159_));
 sg13g2_nor2_1 _2275_ (.A(net62),
    .B(_0291_),
    .Y(_0509_));
 sg13g2_a21oi_1 _2276_ (.A1(_0647_),
    .A2(\counter.oled_driver.spi_data[0] ),
    .Y(_0510_),
    .B1(_0509_));
 sg13g2_nand2_1 _2277_ (.Y(_0511_),
    .A(_0749_),
    .B(_0510_));
 sg13g2_o21ai_1 _2278_ (.B1(_0511_),
    .Y(_0512_),
    .A1(net56),
    .A2(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[0] ));
 sg13g2_nor2_1 _2279_ (.A(_0746_),
    .B(_0512_),
    .Y(_0164_));
 sg13g2_nor2b_1 _2280_ (.A(net62),
    .B_N(_0666_),
    .Y(_0513_));
 sg13g2_a22oi_1 _2281_ (.Y(_0514_),
    .B1(net37),
    .B2(_0513_),
    .A2(\counter.oled_driver.spi_data[1] ),
    .A1(net47));
 sg13g2_nor2_1 _2282_ (.A(net69),
    .B(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1] ),
    .Y(_0515_));
 sg13g2_a21oi_1 _2283_ (.A1(net56),
    .A2(_0514_),
    .Y(_0516_),
    .B1(_0515_));
 sg13g2_nor2b_1 _2284_ (.A(net36),
    .B_N(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[0] ),
    .Y(_0517_));
 sg13g2_a21oi_1 _2285_ (.A1(net30),
    .A2(_0516_),
    .Y(_0518_),
    .B1(_0517_));
 sg13g2_nor2_1 _2286_ (.A(net43),
    .B(_0518_),
    .Y(_0165_));
 sg13g2_inv_1 _2287_ (.Y(_0519_),
    .A(_0047_));
 sg13g2_nor2b_1 _2288_ (.A(net62),
    .B_N(net74),
    .Y(_0520_));
 sg13g2_a22oi_1 _2289_ (.Y(_0521_),
    .B1(net37),
    .B2(_0520_),
    .A2(_0519_),
    .A1(net47));
 sg13g2_nor2_1 _2290_ (.A(net69),
    .B(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2] ),
    .Y(_0522_));
 sg13g2_a21oi_1 _2291_ (.A1(net56),
    .A2(_0521_),
    .Y(_0523_),
    .B1(_0522_));
 sg13g2_nor2b_1 _2292_ (.A(net36),
    .B_N(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1] ),
    .Y(_0524_));
 sg13g2_a21oi_1 _2293_ (.A1(net30),
    .A2(_0523_),
    .Y(_0525_),
    .B1(_0524_));
 sg13g2_nor2_1 _2294_ (.A(net43),
    .B(_0525_),
    .Y(_0166_));
 sg13g2_mux2_1 _2295_ (.A0(_0048_),
    .A1(_0266_),
    .S(_0799_),
    .X(_0526_));
 sg13g2_nor2_1 _2296_ (.A(_0748_),
    .B(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3] ),
    .Y(_0527_));
 sg13g2_a21oi_1 _2297_ (.A1(net56),
    .A2(_0526_),
    .Y(_0528_),
    .B1(_0527_));
 sg13g2_nor2b_1 _2298_ (.A(_0744_),
    .B_N(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2] ),
    .Y(_0529_));
 sg13g2_a21oi_1 _2299_ (.A1(net30),
    .A2(_0528_),
    .Y(_0530_),
    .B1(_0529_));
 sg13g2_nor2_1 _2300_ (.A(net43),
    .B(_0530_),
    .Y(_0167_));
 sg13g2_nor2_1 _2301_ (.A(_0646_),
    .B(_0654_),
    .Y(_0531_));
 sg13g2_a22oi_1 _2302_ (.Y(_0532_),
    .B1(net37),
    .B2(_0531_),
    .A2(\counter.oled_driver.spi_data[4] ),
    .A1(net47));
 sg13g2_nor2_1 _2303_ (.A(_0748_),
    .B(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4] ),
    .Y(_0533_));
 sg13g2_a21oi_1 _2304_ (.A1(net56),
    .A2(_0532_),
    .Y(_0534_),
    .B1(_0533_));
 sg13g2_nor2b_1 _2305_ (.A(_0744_),
    .B_N(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3] ),
    .Y(_0535_));
 sg13g2_a21oi_1 _2306_ (.A1(net30),
    .A2(_0534_),
    .Y(_0536_),
    .B1(_0535_));
 sg13g2_nor2_1 _2307_ (.A(_0253_),
    .B(_0536_),
    .Y(_0168_));
 sg13g2_and3_1 _2308_ (.X(_0537_),
    .A(_0799_),
    .B(_0655_),
    .C(net37));
 sg13g2_a21oi_1 _2309_ (.A1(_0647_),
    .A2(\counter.oled_driver.spi_data[5] ),
    .Y(_0538_),
    .B1(_0537_));
 sg13g2_nor2_1 _2310_ (.A(net69),
    .B(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[5] ),
    .Y(_0539_));
 sg13g2_a21oi_1 _2311_ (.A1(net56),
    .A2(_0538_),
    .Y(_0540_),
    .B1(_0539_));
 sg13g2_nor2b_1 _2312_ (.A(net36),
    .B_N(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4] ),
    .Y(_0541_));
 sg13g2_a21oi_1 _2313_ (.A1(_0745_),
    .A2(_0540_),
    .Y(_0542_),
    .B1(_0541_));
 sg13g2_nor2_1 _2314_ (.A(_0253_),
    .B(_0542_),
    .Y(_0169_));
 sg13g2_nor2b_1 _2315_ (.A(net62),
    .B_N(_0656_),
    .Y(_0543_));
 sg13g2_a22oi_1 _2316_ (.Y(_0544_),
    .B1(_0663_),
    .B2(_0543_),
    .A2(\counter.oled_driver.spi_data[6] ),
    .A1(net62));
 sg13g2_nor2_1 _2317_ (.A(net69),
    .B(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6] ),
    .Y(_0545_));
 sg13g2_a21oi_1 _2318_ (.A1(net69),
    .A2(_0544_),
    .Y(_0546_),
    .B1(_0545_));
 sg13g2_nor2b_1 _2319_ (.A(net36),
    .B_N(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[5] ),
    .Y(_0547_));
 sg13g2_a21oi_1 _2320_ (.A1(_0745_),
    .A2(_0546_),
    .Y(_0548_),
    .B1(_0547_));
 sg13g2_nor2_1 _2321_ (.A(net60),
    .B(_0548_),
    .Y(_0170_));
 sg13g2_inv_1 _2322_ (.Y(_0549_),
    .A(_0049_));
 sg13g2_nor2_1 _2323_ (.A(net62),
    .B(_0691_),
    .Y(_0550_));
 sg13g2_a22oi_1 _2324_ (.Y(_0551_),
    .B1(_0663_),
    .B2(_0550_),
    .A2(_0549_),
    .A1(_0646_));
 sg13g2_nor2_1 _2325_ (.A(net69),
    .B(\counter.oled_driver.oled_mosi_out ),
    .Y(_0552_));
 sg13g2_a21oi_1 _2326_ (.A1(net69),
    .A2(_0551_),
    .Y(_0553_),
    .B1(_0552_));
 sg13g2_nor2b_1 _2327_ (.A(net36),
    .B_N(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6] ),
    .Y(_0554_));
 sg13g2_a21oi_1 _2328_ (.A1(net30),
    .A2(_0553_),
    .Y(_0555_),
    .B1(_0554_));
 sg13g2_nor2_1 _2329_ (.A(_0676_),
    .B(_0555_),
    .Y(_0171_));
 sg13g2_buf_1 _2330_ (.A(net70),
    .X(_0556_));
 sg13g2_nand3b_1 _2331_ (.B(\counter.state[1] ),
    .C(_0774_),
    .Y(_0557_),
    .A_N(net57));
 sg13g2_nor4_1 _2332_ (.A(\counter.state[1] ),
    .B(_0710_),
    .C(_0720_),
    .D(_0732_),
    .Y(_0558_));
 sg13g2_a21oi_1 _2333_ (.A1(net50),
    .A2(_0557_),
    .Y(_0559_),
    .B1(_0558_));
 sg13g2_nor2_1 _2334_ (.A(net60),
    .B(_0559_),
    .Y(_0172_));
 sg13g2_nor2_1 _2335_ (.A(net66),
    .B(_1154_),
    .Y(_0560_));
 sg13g2_inv_1 _2336_ (.Y(_0561_),
    .A(_1154_));
 sg13g2_nor4_1 _2337_ (.A(_0064_),
    .B(_0063_),
    .C(_0764_),
    .D(_0561_),
    .Y(_0562_));
 sg13g2_o21ai_1 _2338_ (.B1(net58),
    .Y(_0173_),
    .A1(_0560_),
    .A2(_0562_));
 sg13g2_nor3_1 _2339_ (.A(net66),
    .B(net54),
    .C(_0065_),
    .Y(_0563_));
 sg13g2_a22oi_1 _2340_ (.Y(_0564_),
    .B1(_1154_),
    .B2(_0563_),
    .A2(net54),
    .A1(net66));
 sg13g2_inv_1 _2341_ (.Y(_0565_),
    .A(_0564_));
 sg13g2_a22oi_1 _2342_ (.Y(_0566_),
    .B1(_0565_),
    .B2(net64),
    .A2(_0561_),
    .A1(_0762_));
 sg13g2_nor2_1 _2343_ (.A(net60),
    .B(_0566_),
    .Y(_0174_));
 sg13g2_nor2_1 _2344_ (.A(net66),
    .B(net54),
    .Y(_0567_));
 sg13g2_nand3_1 _2345_ (.B(_0567_),
    .C(_1154_),
    .A(net65),
    .Y(_0568_));
 sg13g2_or2_1 _2346_ (.X(_0569_),
    .B(_0567_),
    .A(_0763_));
 sg13g2_a21oi_1 _2347_ (.A1(_0568_),
    .A2(_0569_),
    .Y(_0570_),
    .B1(_0063_));
 sg13g2_nor2_1 _2348_ (.A(_0763_),
    .B(_1154_),
    .Y(_0571_));
 sg13g2_o21ai_1 _2349_ (.B1(net58),
    .Y(_0175_),
    .A1(_0570_),
    .A2(_0571_));
 sg13g2_nand3_1 _2350_ (.B(net50),
    .C(\counter.cnt_x_digits[0] ),
    .A(net53),
    .Y(_0572_));
 sg13g2_nand2_2 _2351_ (.Y(_0573_),
    .A(_0706_),
    .B(net70));
 sg13g2_buf_1 _2352_ (.A(_0573_),
    .X(_0574_));
 sg13g2_nand2_1 _2353_ (.Y(_0575_),
    .A(\counter.streamer.digits_r[0] ),
    .B(net41));
 sg13g2_a21oi_1 _2354_ (.A1(_0572_),
    .A2(_0575_),
    .Y(_0176_),
    .B1(net46));
 sg13g2_nand3_1 _2355_ (.B(net50),
    .C(\counter.cnt_x_digits[10] ),
    .A(net53),
    .Y(_0576_));
 sg13g2_nand2_1 _2356_ (.Y(_0577_),
    .A(\counter.streamer.digits_r[10] ),
    .B(net41));
 sg13g2_a21oi_1 _2357_ (.A1(_0576_),
    .A2(_0577_),
    .Y(_0177_),
    .B1(net46));
 sg13g2_nand3_1 _2358_ (.B(net50),
    .C(\counter.cnt_x_digits[11] ),
    .A(net53),
    .Y(_0578_));
 sg13g2_nand2_1 _2359_ (.Y(_0579_),
    .A(\counter.streamer.digits_r[11] ),
    .B(net41));
 sg13g2_a21oi_1 _2360_ (.A1(_0578_),
    .A2(_0579_),
    .Y(_0178_),
    .B1(net46));
 sg13g2_nand3_1 _2361_ (.B(net50),
    .C(\counter.cnt_x_digits[12] ),
    .A(net53),
    .Y(_0580_));
 sg13g2_nand2_1 _2362_ (.Y(_0581_),
    .A(\counter.streamer.digits_r[12] ),
    .B(net41));
 sg13g2_a21oi_1 _2363_ (.A1(_0580_),
    .A2(_0581_),
    .Y(_0179_),
    .B1(net46));
 sg13g2_nand3_1 _2364_ (.B(net50),
    .C(_1036_),
    .A(net53),
    .Y(_0582_));
 sg13g2_nand2_1 _2365_ (.Y(_0583_),
    .A(\counter.streamer.digits_r[13] ),
    .B(net41));
 sg13g2_a21oi_1 _2366_ (.A1(_0582_),
    .A2(_0583_),
    .Y(_0180_),
    .B1(net46));
 sg13g2_nand3_1 _2367_ (.B(net50),
    .C(\counter.cnt_x_digits[14] ),
    .A(net53),
    .Y(_0584_));
 sg13g2_nand2_1 _2368_ (.Y(_0585_),
    .A(\counter.streamer.digits_r[14] ),
    .B(net41));
 sg13g2_buf_1 _2369_ (.A(net63),
    .X(_0586_));
 sg13g2_a21oi_1 _2370_ (.A1(_0584_),
    .A2(_0585_),
    .Y(_0181_),
    .B1(net40));
 sg13g2_nand3_1 _2371_ (.B(net50),
    .C(\counter.cnt_x_digits[15] ),
    .A(net53),
    .Y(_0587_));
 sg13g2_nand2_1 _2372_ (.Y(_0588_),
    .A(\counter.streamer.digits_r[15] ),
    .B(net41));
 sg13g2_a21oi_1 _2373_ (.A1(_0587_),
    .A2(_0588_),
    .Y(_0182_),
    .B1(net40));
 sg13g2_nand3_1 _2374_ (.B(_0556_),
    .C(\counter.cnt_x_digits[16] ),
    .A(_0775_),
    .Y(_0589_));
 sg13g2_nand2_1 _2375_ (.Y(_0590_),
    .A(\counter.streamer.digits_r[16] ),
    .B(net41));
 sg13g2_a21oi_1 _2376_ (.A1(_0589_),
    .A2(_0590_),
    .Y(_0183_),
    .B1(net40));
 sg13g2_nand3_1 _2377_ (.B(_0556_),
    .C(\counter.cnt_x_digits[17] ),
    .A(_0775_),
    .Y(_0591_));
 sg13g2_nand2_1 _2378_ (.Y(_0592_),
    .A(\counter.streamer.digits_r[17] ),
    .B(_0574_));
 sg13g2_a21oi_1 _2379_ (.A1(_0591_),
    .A2(_0592_),
    .Y(_0184_),
    .B1(net40));
 sg13g2_buf_1 _2380_ (.A(net57),
    .X(_0593_));
 sg13g2_buf_1 _2381_ (.A(_0736_),
    .X(_0594_));
 sg13g2_nand3_1 _2382_ (.B(net49),
    .C(\counter.cnt_x_digits[18] ),
    .A(net39),
    .Y(_0595_));
 sg13g2_nand2_1 _2383_ (.Y(_0596_),
    .A(\counter.streamer.digits_r[18] ),
    .B(_0574_));
 sg13g2_a21oi_1 _2384_ (.A1(_0595_),
    .A2(_0596_),
    .Y(_0185_),
    .B1(_0586_));
 sg13g2_nand3_1 _2385_ (.B(net49),
    .C(\counter.cnt_x_digits[19] ),
    .A(net39),
    .Y(_0597_));
 sg13g2_buf_1 _2386_ (.A(_0573_),
    .X(_0598_));
 sg13g2_nand2_1 _2387_ (.Y(_0599_),
    .A(\counter.streamer.digits_r[19] ),
    .B(net38));
 sg13g2_a21oi_1 _2388_ (.A1(_0597_),
    .A2(_0599_),
    .Y(_0186_),
    .B1(net40));
 sg13g2_nand3_1 _2389_ (.B(net49),
    .C(\counter.cnt_x_digits[1] ),
    .A(net39),
    .Y(_0600_));
 sg13g2_nand2_1 _2390_ (.Y(_0601_),
    .A(\counter.streamer.digits_r[1] ),
    .B(_0598_));
 sg13g2_a21oi_1 _2391_ (.A1(_0600_),
    .A2(_0601_),
    .Y(_0187_),
    .B1(_0586_));
 sg13g2_nand3_1 _2392_ (.B(net49),
    .C(\counter.cnt_x_digits[20] ),
    .A(net39),
    .Y(_0602_));
 sg13g2_nand2_1 _2393_ (.Y(_0603_),
    .A(\counter.streamer.digits_r[20] ),
    .B(net38));
 sg13g2_a21oi_1 _2394_ (.A1(_0602_),
    .A2(_0603_),
    .Y(_0188_),
    .B1(net40));
 sg13g2_nand3_1 _2395_ (.B(net49),
    .C(\counter.cnt_x_digits[21] ),
    .A(net39),
    .Y(_0604_));
 sg13g2_nand2_1 _2396_ (.Y(_0605_),
    .A(\counter.streamer.digits_r[21] ),
    .B(net38));
 sg13g2_a21oi_1 _2397_ (.A1(_0604_),
    .A2(_0605_),
    .Y(_0189_),
    .B1(net40));
 sg13g2_nand3_1 _2398_ (.B(_0594_),
    .C(\counter.cnt_x_digits[22] ),
    .A(_0593_),
    .Y(_0606_));
 sg13g2_nand2_1 _2399_ (.Y(_0607_),
    .A(\counter.streamer.digits_r[22] ),
    .B(_0598_));
 sg13g2_a21oi_1 _2400_ (.A1(_0606_),
    .A2(_0607_),
    .Y(_0190_),
    .B1(net40));
 sg13g2_nand3_1 _2401_ (.B(_0594_),
    .C(\counter.cnt_x_digits[23] ),
    .A(_0593_),
    .Y(_0608_));
 sg13g2_nand2_1 _2402_ (.Y(_0609_),
    .A(\counter.streamer.digits_r[23] ),
    .B(net38));
 sg13g2_a21oi_1 _2403_ (.A1(_0608_),
    .A2(_0609_),
    .Y(_0191_),
    .B1(_0989_));
 sg13g2_nand3_1 _2404_ (.B(net49),
    .C(\counter.cnt_x_digits[2] ),
    .A(net39),
    .Y(_0610_));
 sg13g2_nand2_1 _2405_ (.Y(_0611_),
    .A(\counter.streamer.digits_r[2] ),
    .B(net38));
 sg13g2_a21oi_1 _2406_ (.A1(_0610_),
    .A2(_0611_),
    .Y(_0192_),
    .B1(net51));
 sg13g2_nand3_1 _2407_ (.B(net49),
    .C(\counter.cnt_x_digits[3] ),
    .A(net39),
    .Y(_0612_));
 sg13g2_nand2_1 _2408_ (.Y(_0613_),
    .A(\counter.streamer.digits_r[3] ),
    .B(net38));
 sg13g2_a21oi_1 _2409_ (.A1(_0612_),
    .A2(_0613_),
    .Y(_0193_),
    .B1(net51));
 sg13g2_nand3_1 _2410_ (.B(net49),
    .C(\counter.cnt_x_digits[4] ),
    .A(net39),
    .Y(_0614_));
 sg13g2_nand2_1 _2411_ (.Y(_0615_),
    .A(\counter.streamer.digits_r[4] ),
    .B(net38));
 sg13g2_a21oi_1 _2412_ (.A1(_0614_),
    .A2(_0615_),
    .Y(_0194_),
    .B1(net51));
 sg13g2_nand3_1 _2413_ (.B(_0736_),
    .C(_1006_),
    .A(_0737_),
    .Y(_0616_));
 sg13g2_nand2_1 _2414_ (.Y(_0617_),
    .A(\counter.streamer.digits_r[5] ),
    .B(net38));
 sg13g2_a21oi_1 _2415_ (.A1(_0616_),
    .A2(_0617_),
    .Y(_0195_),
    .B1(net51));
 sg13g2_nand3_1 _2416_ (.B(net70),
    .C(\counter.cnt_x_digits[6] ),
    .A(net57),
    .Y(_0618_));
 sg13g2_nand2_1 _2417_ (.Y(_0619_),
    .A(\counter.streamer.digits_r[6] ),
    .B(_0573_));
 sg13g2_a21oi_1 _2418_ (.A1(_0618_),
    .A2(_0619_),
    .Y(_0196_),
    .B1(net51));
 sg13g2_nand3_1 _2419_ (.B(net70),
    .C(\counter.cnt_x_digits[7] ),
    .A(net57),
    .Y(_0620_));
 sg13g2_nand2_1 _2420_ (.Y(_0621_),
    .A(\counter.streamer.digits_r[7] ),
    .B(_0573_));
 sg13g2_a21oi_1 _2421_ (.A1(_0620_),
    .A2(_0621_),
    .Y(_0197_),
    .B1(net51));
 sg13g2_nand3_1 _2422_ (.B(net70),
    .C(_1017_),
    .A(net57),
    .Y(_0622_));
 sg13g2_nand2_1 _2423_ (.Y(_0623_),
    .A(\counter.streamer.digits_r[8] ),
    .B(_0573_));
 sg13g2_a21oi_1 _2424_ (.A1(_0622_),
    .A2(_0623_),
    .Y(_0198_),
    .B1(net51));
 sg13g2_nand3_1 _2425_ (.B(net70),
    .C(_1020_),
    .A(_0737_),
    .Y(_0624_));
 sg13g2_nand2_1 _2426_ (.Y(_0625_),
    .A(\counter.streamer.digits_r[9] ),
    .B(_0573_));
 sg13g2_a21oi_1 _2427_ (.A1(_0624_),
    .A2(_0625_),
    .Y(_0199_),
    .B1(_0989_));
 sg13g2_nand2_1 _2428_ (.Y(_0626_),
    .A(net61),
    .B(_0707_));
 sg13g2_nand2b_1 _2429_ (.Y(_0627_),
    .B(net67),
    .A_N(_0673_));
 sg13g2_o21ai_1 _2430_ (.B1(_0627_),
    .Y(_0628_),
    .A1(net67),
    .A2(_0626_));
 sg13g2_a22oi_1 _2431_ (.Y(_0629_),
    .B1(_0628_),
    .B2(net64),
    .A2(_1151_),
    .A1(net67));
 sg13g2_nor2_1 _2432_ (.A(net60),
    .B(_0629_),
    .Y(_0209_));
 sg13g2_and2_1 _2433_ (.A(net67),
    .B(net61),
    .X(_0630_));
 sg13g2_nand3_1 _2434_ (.B(_0707_),
    .C(_0630_),
    .A(net42),
    .Y(_0631_));
 sg13g2_o21ai_1 _2435_ (.B1(_0631_),
    .Y(_0632_),
    .A1(net42),
    .A2(_0630_));
 sg13g2_a22oi_1 _2436_ (.Y(_0633_),
    .B1(_0632_),
    .B2(net64),
    .A2(_1151_),
    .A1(net55));
 sg13g2_nor2_1 _2437_ (.A(net60),
    .B(_0633_),
    .Y(_0210_));
 sg13g2_nor2_1 _2438_ (.A(clknet_5_19__leaf_clk),
    .B(_0991_),
    .Y(\counter.oled_clk_out ));
 sg13g2_or2_1 _2439_ (.X(\counter.oled_dc_out ),
    .B(\counter.oled_driver.mc_exec.oled_dc_out ),
    .A(net47));
 sg13g2_dfrbp_1 _2440_ (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net99),
    .D(_0000_),
    .Q_N(_1279_),
    .Q(_0033_));
 sg13g2_dfrbp_1 _2441_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net100),
    .D(_0001_),
    .Q_N(_1280_),
    .Q(_0034_));
 sg13g2_dfrbp_1 _2442_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net101),
    .D(_0002_),
    .Q_N(_1281_),
    .Q(_0035_));
 sg13g2_dfrbp_1 _2443_ (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net102),
    .D(_0003_),
    .Q_N(_1282_),
    .Q(_0036_));
 sg13g2_dfrbp_1 _2444_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net103),
    .D(_0004_),
    .Q_N(_1283_),
    .Q(_0037_));
 sg13g2_dfrbp_1 _2445_ (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net104),
    .D(_0005_),
    .Q_N(_1284_),
    .Q(_0038_));
 sg13g2_dfrbp_1 _2446_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net105),
    .D(_0006_),
    .Q_N(_1285_),
    .Q(_0039_));
 sg13g2_dfrbp_1 _2447_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net106),
    .D(_0007_),
    .Q_N(_1286_),
    .Q(_0040_));
 sg13g2_dfrbp_1 _2448_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net107),
    .D(_0008_),
    .Q_N(_1287_),
    .Q(_0041_));
 sg13g2_dfrbp_1 _2449_ (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net108),
    .D(_0009_),
    .Q_N(_1278_),
    .Q(_0042_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _2440__99 (.L_HI(net99));
 sg13g2_buf_1 _2452_ (.A(net83),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2453_ (.A(net84),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2454_ (.A(net85),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2455_ (.A(net86),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2456_ (.A(net87),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2457_ (.A(net88),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2458_ (.A(net89),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2459_ (.A(net90),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2460_ (.A(net91),
    .X(uio_out[0]));
 sg13g2_buf_1 _2461_ (.A(net92),
    .X(uio_out[1]));
 sg13g2_buf_1 _2462_ (.A(net93),
    .X(uio_out[2]));
 sg13g2_buf_1 _2463_ (.A(net94),
    .X(uio_out[3]));
 sg13g2_buf_1 _2464_ (.A(net95),
    .X(uio_out[4]));
 sg13g2_buf_1 _2465_ (.A(net96),
    .X(uio_out[5]));
 sg13g2_buf_1 _2466_ (.A(net97),
    .X(uio_out[6]));
 sg13g2_buf_1 _2467_ (.A(net98),
    .X(uio_out[7]));
 sg13g2_buf_1 _2468_ (.A(\counter.oled_driver.mc_exec.oled_rstn_out ),
    .X(net3));
 sg13g2_buf_1 _2469_ (.A(\counter.oled_driver.mc_exec.oled_vbatn_out ),
    .X(net4));
 sg13g2_buf_1 _2470_ (.A(\counter.oled_driver.mc_exec.oled_vcdn_out ),
    .X(net5));
 sg13g2_buf_1 _2471_ (.A(\counter.oled_csn_out ),
    .X(net6));
 sg13g2_buf_1 _2472_ (.A(\counter.oled_dc_out ),
    .X(net7));
 sg13g2_buf_1 _2473_ (.A(\counter.oled_clk_out ),
    .X(net8));
 sg13g2_buf_1 _2474_ (.A(\counter.oled_driver.oled_mosi_out ),
    .X(net9));
 sg13g2_buf_1 _2475_ (.A(ui_in[7]),
    .X(net10));
 sg13g2_dfrbp_1 \counter.counter_ref.digit_0.digit_out[0]$_SDFFE_PP0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net109),
    .D(_0074_),
    .Q_N(_1277_),
    .Q(\counter.counter_ref.digit_0.digit_out[0] ));
 sg13g2_dfrbp_1 \counter.counter_ref.digit_0.digit_out[1]$_SDFFE_PP0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net110),
    .D(_0075_),
    .Q_N(_1276_),
    .Q(\counter.counter_ref.digit_0.digit_out[1] ));
 sg13g2_dfrbp_1 \counter.counter_ref.digit_0.digit_out[2]$_SDFFE_PP0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net111),
    .D(_0076_),
    .Q_N(_1275_),
    .Q(\counter.counter_ref.digit_0.digit_out[2] ));
 sg13g2_dfrbp_1 \counter.counter_ref.digit_0.digit_out[3]$_SDFFE_PP0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net112),
    .D(_0077_),
    .Q_N(_1274_),
    .Q(\counter.counter_ref.digit_0.digit_out[3] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[1].digit_x.digit_out[0]$_SDFFE_PP0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net113),
    .D(_0078_),
    .Q_N(_1273_),
    .Q(\counter.counter_ref.digits_out[4] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[1].digit_x.digit_out[1]$_SDFFE_PP0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net114),
    .D(_0079_),
    .Q_N(_1272_),
    .Q(\counter.counter_ref.digits_out[5] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[1].digit_x.digit_out[2]$_SDFFE_PP0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net115),
    .D(_0080_),
    .Q_N(_1271_),
    .Q(\counter.counter_ref.digits_out[6] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[1].digit_x.digit_out[3]$_SDFFE_PP0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net116),
    .D(_0081_),
    .Q_N(_1270_),
    .Q(\counter.counter_ref.digits_out[7] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[2].digit_x.digit_out[0]$_SDFFE_PP0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net117),
    .D(_0082_),
    .Q_N(_1269_),
    .Q(\counter.counter_ref.digits_out[8] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[2].digit_x.digit_out[1]$_SDFFE_PP0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net118),
    .D(_0083_),
    .Q_N(_1268_),
    .Q(\counter.counter_ref.digits_out[9] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[2].digit_x.digit_out[2]$_SDFFE_PP0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net119),
    .D(_0084_),
    .Q_N(_1267_),
    .Q(\counter.counter_ref.digits_out[10] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[2].digit_x.digit_out[3]$_SDFFE_PP0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net120),
    .D(_0085_),
    .Q_N(_1266_),
    .Q(\counter.counter_ref.digits_out[11] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[3].digit_x.digit_out[0]$_SDFFE_PP0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net121),
    .D(_0086_),
    .Q_N(_1265_),
    .Q(\counter.counter_ref.digits_out[12] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[3].digit_x.digit_out[1]$_SDFFE_PP0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net122),
    .D(_0087_),
    .Q_N(_1264_),
    .Q(\counter.counter_ref.digits_out[13] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[3].digit_x.digit_out[2]$_SDFFE_PP0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net123),
    .D(_0088_),
    .Q_N(_1263_),
    .Q(\counter.counter_ref.digits_out[14] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[3].digit_x.digit_out[3]$_SDFFE_PP0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net124),
    .D(_0089_),
    .Q_N(_1262_),
    .Q(\counter.counter_ref.digits_out[15] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[4].digit_x.digit_out[0]$_SDFFE_PP0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net125),
    .D(_0090_),
    .Q_N(_1261_),
    .Q(\counter.counter_ref.digits_out[16] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[4].digit_x.digit_out[1]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net126),
    .D(_0091_),
    .Q_N(_1260_),
    .Q(\counter.counter_ref.digits_out[17] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[4].digit_x.digit_out[2]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net127),
    .D(_0092_),
    .Q_N(_1259_),
    .Q(\counter.counter_ref.digits_out[18] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[4].digit_x.digit_out[3]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net128),
    .D(_0093_),
    .Q_N(_1258_),
    .Q(\counter.counter_ref.digits_out[19] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[5].digit_x.digit_out[0]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net129),
    .D(_0094_),
    .Q_N(_1257_),
    .Q(\counter.counter_ref.digits_out[20] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[5].digit_x.digit_out[1]$_SDFFE_PP0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net130),
    .D(_0095_),
    .Q_N(_1256_),
    .Q(\counter.counter_ref.digits_out[21] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[5].digit_x.digit_out[2]$_SDFFE_PP0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net131),
    .D(_0096_),
    .Q_N(_1255_),
    .Q(\counter.counter_ref.digits_out[22] ));
 sg13g2_dfrbp_1 \counter.counter_ref.genblk1[5].digit_x.digit_out[3]$_SDFFE_PP0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net132),
    .D(_0097_),
    .Q_N(_1254_),
    .Q(\counter.counter_ref.digits_out[23] ));
 sg13g2_dfrbp_1 \counter.counter_x.digit_0.digit_out[0]$_DFFE_PP0P_  (.CLK(net80),
    .RESET_B(net33),
    .D(_0098_),
    .Q_N(_1253_),
    .Q(\counter.cnt_x_digits[0] ));
 sg13g2_dfrbp_1 \counter.counter_x.digit_0.digit_out[1]$_DFFE_PP0P_  (.CLK(net80),
    .RESET_B(net33),
    .D(_0099_),
    .Q_N(_1252_),
    .Q(\counter.cnt_x_digits[1] ));
 sg13g2_dfrbp_1 \counter.counter_x.digit_0.digit_out[2]$_DFFE_PP0P_  (.CLK(net80),
    .RESET_B(net34),
    .D(_0100_),
    .Q_N(_1251_),
    .Q(\counter.cnt_x_digits[2] ));
 sg13g2_dfrbp_1 \counter.counter_x.digit_0.digit_out[3]$_DFFE_PP0P_  (.CLK(net80),
    .RESET_B(net34),
    .D(_0101_),
    .Q_N(_1250_),
    .Q(\counter.cnt_x_digits[3] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[1].digit_x.digit_out[0]$_DFFE_PP0P_  (.CLK(net82),
    .RESET_B(net35),
    .D(_0102_),
    .Q_N(_1249_),
    .Q(\counter.cnt_x_digits[4] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[1].digit_x.digit_out[1]$_DFFE_PP0P_  (.CLK(net79),
    .RESET_B(net32),
    .D(_0103_),
    .Q_N(_1248_),
    .Q(\counter.cnt_x_digits[5] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[1].digit_x.digit_out[2]$_DFFE_PP0P_  (.CLK(net81),
    .RESET_B(net34),
    .D(_0104_),
    .Q_N(_1247_),
    .Q(\counter.cnt_x_digits[6] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[1].digit_x.digit_out[3]$_DFFE_PP0P_  (.CLK(net79),
    .RESET_B(net32),
    .D(_0105_),
    .Q_N(_1246_),
    .Q(\counter.cnt_x_digits[7] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[2].digit_x.digit_out[0]$_DFFE_PP0P_  (.CLK(net79),
    .RESET_B(net32),
    .D(_0106_),
    .Q_N(_1245_),
    .Q(\counter.cnt_x_digits[8] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[2].digit_x.digit_out[1]$_DFFE_PP0P_  (.CLK(net79),
    .RESET_B(net32),
    .D(_0107_),
    .Q_N(_1244_),
    .Q(\counter.cnt_x_digits[9] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[2].digit_x.digit_out[2]$_DFFE_PP0P_  (.CLK(net79),
    .RESET_B(net32),
    .D(_0108_),
    .Q_N(_1243_),
    .Q(\counter.cnt_x_digits[10] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[2].digit_x.digit_out[3]$_DFFE_PP0P_  (.CLK(net79),
    .RESET_B(net32),
    .D(_0109_),
    .Q_N(_1242_),
    .Q(\counter.cnt_x_digits[11] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[3].digit_x.digit_out[0]$_DFFE_PP0P_  (.CLK(net79),
    .RESET_B(net32),
    .D(_0110_),
    .Q_N(_1241_),
    .Q(\counter.cnt_x_digits[12] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[3].digit_x.digit_out[1]$_DFFE_PP0P_  (.CLK(net79),
    .RESET_B(net32),
    .D(_0111_),
    .Q_N(_1240_),
    .Q(\counter.cnt_x_digits[13] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[3].digit_x.digit_out[2]$_DFFE_PP0P_  (.CLK(net80),
    .RESET_B(net33),
    .D(_0112_),
    .Q_N(_1239_),
    .Q(\counter.cnt_x_digits[14] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[3].digit_x.digit_out[3]$_DFFE_PP0P_  (.CLK(net80),
    .RESET_B(net33),
    .D(_0113_),
    .Q_N(_1238_),
    .Q(\counter.cnt_x_digits[15] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[4].digit_x.digit_out[0]$_DFFE_PP0P_  (.CLK(net80),
    .RESET_B(net33),
    .D(_0114_),
    .Q_N(_1237_),
    .Q(\counter.cnt_x_digits[16] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[4].digit_x.digit_out[1]$_DFFE_PP0P_  (.CLK(net81),
    .RESET_B(net33),
    .D(_0115_),
    .Q_N(_1236_),
    .Q(\counter.cnt_x_digits[17] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[4].digit_x.digit_out[2]$_DFFE_PP0P_  (.CLK(net81),
    .RESET_B(net34),
    .D(_0116_),
    .Q_N(_1235_),
    .Q(\counter.cnt_x_digits[18] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[4].digit_x.digit_out[3]$_DFFE_PP0P_  (.CLK(net81),
    .RESET_B(net33),
    .D(_0117_),
    .Q_N(_1234_),
    .Q(\counter.cnt_x_digits[19] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[5].digit_x.digit_out[0]$_DFFE_PP0P_  (.CLK(net82),
    .RESET_B(net35),
    .D(_0118_),
    .Q_N(_1233_),
    .Q(\counter.cnt_x_digits[20] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[5].digit_x.digit_out[1]$_DFFE_PP0P_  (.CLK(net82),
    .RESET_B(net35),
    .D(_0119_),
    .Q_N(_1232_),
    .Q(\counter.cnt_x_digits[21] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[5].digit_x.digit_out[2]$_DFFE_PP0P_  (.CLK(net82),
    .RESET_B(net35),
    .D(_0120_),
    .Q_N(_1231_),
    .Q(\counter.cnt_x_digits[22] ));
 sg13g2_dfrbp_1 \counter.counter_x.genblk1[5].digit_x.digit_out[3]$_DFFE_PP0P_  (.CLK(net82),
    .RESET_B(net35),
    .D(_0121_),
    .Q_N(_1230_),
    .Q(\counter.cnt_x_digits[23] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[0]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net133),
    .D(_0122_),
    .Q_N(_1229_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[0] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[10]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net134),
    .D(_0123_),
    .Q_N(_1228_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[10] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[11]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net135),
    .D(_0124_),
    .Q_N(_1227_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[11] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[12]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net136),
    .D(_0125_),
    .Q_N(_1226_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[12] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[13]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net137),
    .D(_0126_),
    .Q_N(_1225_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[13] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[14]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net138),
    .D(_0127_),
    .Q_N(_1224_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[14] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[15]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net139),
    .D(_0128_),
    .Q_N(_1223_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[15] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[16]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net140),
    .D(_0129_),
    .Q_N(_0052_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[16] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[1]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net141),
    .D(_0130_),
    .Q_N(_1222_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[1] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[2]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net142),
    .D(_0131_),
    .Q_N(_1221_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[2] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[3]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net143),
    .D(_0132_),
    .Q_N(_1220_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[3] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[4]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net144),
    .D(_0133_),
    .Q_N(_1219_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[4] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[5]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net145),
    .D(_0134_),
    .Q_N(_1218_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[5] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[6]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net146),
    .D(_0135_),
    .Q_N(_1217_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[6] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[7]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net147),
    .D(_0136_),
    .Q_N(_1216_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[7] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[8]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net148),
    .D(_0137_),
    .Q_N(_1215_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[8] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.delay_cnt[9]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net149),
    .D(_0138_),
    .Q_N(_1214_),
    .Q(\counter.oled_driver.mc_exec.delay_cnt[9] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.oled_dc_out$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net150),
    .D(_0139_),
    .Q_N(_1213_),
    .Q(\counter.oled_driver.mc_exec.oled_dc_out ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.oled_rstn_out$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net151),
    .D(_0140_),
    .Q_N(_1212_),
    .Q(\counter.oled_driver.mc_exec.oled_rstn_out ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.oled_vbatn_out$_SDFFE_PN1P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net152),
    .D(_0141_),
    .Q_N(_1211_),
    .Q(\counter.oled_driver.mc_exec.oled_vbatn_out ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.oled_vcdn_out$_SDFFE_PN1P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net153),
    .D(_0142_),
    .Q_N(_1210_),
    .Q(\counter.oled_driver.mc_exec.oled_vcdn_out ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.rom_index_r[0]$_SDFFE_PN0N_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net154),
    .D(_0143_),
    .Q_N(_0058_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[0] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.rom_index_r[1]$_SDFFE_PN0N_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net155),
    .D(_0144_),
    .Q_N(_0059_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[1] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.rom_index_r[2]$_SDFFE_PN0N_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net156),
    .D(_0145_),
    .Q_N(_0056_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[2] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.rom_index_r[3]$_SDFFE_PN0N_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net157),
    .D(_0146_),
    .Q_N(_0057_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[3] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.rom_index_r[4]$_SDFFE_PN0N_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net158),
    .D(_0147_),
    .Q_N(_1209_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[4] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.rom_index_r[5]$_SDFFE_PN0N_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net159),
    .D(_0148_),
    .Q_N(_1288_),
    .Q(\counter.oled_driver.mc_exec.microcode_rom.address[5] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.state_r[1]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net160),
    .D(_0016_),
    .Q_N(_1289_),
    .Q(\counter.oled_driver.mc_exec.spi_tx_trigger_out ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.state_r[2]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net161),
    .D(_0017_),
    .Q_N(_0053_),
    .Q(\counter.oled_driver.mc_exec.state_r[2] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.state_r[3]$_DFF_P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net162),
    .D(_0018_),
    .Q_N(_0054_),
    .Q(\counter.oled_driver.mc_exec.state_r[3] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.state_r[4]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net163),
    .D(_0019_),
    .Q_N(_0051_),
    .Q(\counter.oled_driver.mc_exec.procedure_done_out ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.state_r[5]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net164),
    .D(_0010_),
    .Q_N(_1290_),
    .Q(\counter.oled_driver.mc_exec.state_r[5] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_exec.state_r[6]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net165),
    .D(_0020_),
    .Q_N(_0055_),
    .Q(\counter.oled_driver.mc_exec.state_r[6] ));
 sg13g2_dfrbp_1 \counter.oled_driver.mc_procedure_offset[0]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net166),
    .D(_0149_),
    .Q_N(_1208_),
    .Q(\counter.oled_driver.mc_exec.procedure_offset_in[0] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_data[0]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net167),
    .D(_0150_),
    .Q_N(_1207_),
    .Q(\counter.oled_driver.spi_data[0] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_data[1]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net168),
    .D(_0151_),
    .Q_N(_1206_),
    .Q(\counter.oled_driver.spi_data[1] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_data[2]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net169),
    .D(_0152_),
    .Q_N(_0047_),
    .Q(\counter.oled_driver.spi_data[2] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_data[3]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net170),
    .D(_0153_),
    .Q_N(_0048_),
    .Q(\counter.oled_driver.spi_data[3] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_data[4]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net171),
    .D(_0154_),
    .Q_N(_1205_),
    .Q(\counter.oled_driver.spi_data[4] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_data[5]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net172),
    .D(_0155_),
    .Q_N(_1204_),
    .Q(\counter.oled_driver.spi_data[5] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_data[6]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net173),
    .D(_0156_),
    .Q_N(_1203_),
    .Q(\counter.oled_driver.spi_data[6] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_data[7]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net174),
    .D(_0157_),
    .Q_N(_0049_),
    .Q(\counter.oled_driver.spi_data[7] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.chip_select_r$_SDFFE_PN1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net175),
    .D(_0158_),
    .Q_N(_1202_),
    .Q(\counter.oled_csn_out ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.deactivate_cs_r$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net176),
    .D(_0159_),
    .Q_N(_1201_),
    .Q(\counter.oled_driver.spi_driver.deactivate_cs_r ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0]$_SDFFE_PP0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net177),
    .D(_0160_),
    .Q_N(_0072_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1]$_SDFFE_PP0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net178),
    .D(_0161_),
    .Q_N(_1200_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2]$_SDFFE_PP0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net179),
    .D(_0162_),
    .Q_N(_1199_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3]$_SDFFE_PP0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net180),
    .D(_0163_),
    .Q_N(_1198_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[0]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net181),
    .D(_0164_),
    .Q_N(_1197_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[0] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net182),
    .D(_0165_),
    .Q_N(_1196_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net183),
    .D(_0166_),
    .Q_N(_1195_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net184),
    .D(_0167_),
    .Q_N(_1194_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net185),
    .D(_0168_),
    .Q_N(_1193_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[5]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net186),
    .D(_0169_),
    .Q_N(_1192_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[5] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net187),
    .D(_0170_),
    .Q_N(_1191_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[7]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net188),
    .D(_0171_),
    .Q_N(_1291_),
    .Q(\counter.oled_driver.oled_mosi_out ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.state_r[0]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net189),
    .D(_0021_),
    .Q_N(_1292_),
    .Q(\counter.oled_driver.spi_driver.state_r[0] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.state_r[1]$_DFF_P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net190),
    .D(_0011_),
    .Q_N(_1293_),
    .Q(\counter.oled_driver.spi_driver.state_r[1] ));
 sg13g2_dfrbp_1 \counter.oled_driver.spi_driver.state_r[2]$_DFF_P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net191),
    .D(_0022_),
    .Q_N(_1294_),
    .Q(\counter.oled_driver.spi_driver.shift_reg.start_in ));
 sg13g2_dfrbp_1 \counter.oled_driver.state_r[0]$_DFF_P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net192),
    .D(_0023_),
    .Q_N(_1295_),
    .Q(\counter.oled_driver.state_r[0] ));
 sg13g2_dfrbp_1 \counter.oled_driver.state_r[1]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net193),
    .D(_0024_),
    .Q_N(_1296_),
    .Q(\counter.oled_driver.spi_deactivate_cs ));
 sg13g2_dfrbp_1 \counter.oled_driver.state_r[2]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net194),
    .D(_0012_),
    .Q_N(_1297_),
    .Q(\counter.oled_driver.state_r[2] ));
 sg13g2_dfrbp_1 \counter.oled_driver.state_r[3]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net195),
    .D(_0025_),
    .Q_N(_1298_),
    .Q(\counter.oled_driver.mc_exec.procedure_start_in ));
 sg13g2_dfrbp_1 \counter.oled_driver.state_r[4]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net196),
    .D(_0013_),
    .Q_N(_1299_),
    .Q(\counter.oled_driver.state_r[4] ));
 sg13g2_dfrbp_1 \counter.oled_driver.state_r[5]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net197),
    .D(_0026_),
    .Q_N(_0050_),
    .Q(\counter.oled_driver.ready_out ));
 sg13g2_dfrbp_1 \counter.refresh_display$_SDFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net198),
    .D(_0172_),
    .Q_N(_1300_),
    .Q(\counter.refresh_display ));
 sg13g2_dfrbp_1 \counter.state[0]$_DFF_P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net199),
    .D(_0027_),
    .Q_N(_1301_),
    .Q(\counter.state[0] ));
 sg13g2_dfrbp_1 \counter.state[1]$_DFF_P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net200),
    .D(_0028_),
    .Q_N(_1302_),
    .Q(\counter.state[1] ));
 sg13g2_dfrbp_1 \counter.state[2]$_DFF_P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net201),
    .D(_0029_),
    .Q_N(_1190_),
    .Q(\counter.cnt_ref_enable ));
 sg13g2_dfrbp_1 \counter.streamer.digit_cnt_r[0]$_SDFFE_PN1P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net202),
    .D(_0173_),
    .Q_N(_0064_),
    .Q(\counter.streamer.digit_cnt_r[0] ));
 sg13g2_dfrbp_1 \counter.streamer.digit_cnt_r[1]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net203),
    .D(_0174_),
    .Q_N(_0067_),
    .Q(\counter.streamer.digit_cnt_r[1] ));
 sg13g2_dfrbp_1 \counter.streamer.digit_cnt_r[2]$_SDFFE_PN1P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net204),
    .D(_0175_),
    .Q_N(_0065_),
    .Q(\counter.streamer.digit_cnt_r[2] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[0]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net205),
    .D(_0176_),
    .Q_N(_1189_),
    .Q(\counter.streamer.digits_r[0] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[10]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net206),
    .D(_0177_),
    .Q_N(_1188_),
    .Q(\counter.streamer.digits_r[10] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[11]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net207),
    .D(_0178_),
    .Q_N(_0070_),
    .Q(\counter.streamer.digits_r[11] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[12]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net208),
    .D(_0179_),
    .Q_N(_1187_),
    .Q(\counter.streamer.digits_r[12] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[13]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net209),
    .D(_0180_),
    .Q_N(_1186_),
    .Q(\counter.streamer.digits_r[13] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[14]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net210),
    .D(_0181_),
    .Q_N(_1185_),
    .Q(\counter.streamer.digits_r[14] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[15]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net211),
    .D(_0182_),
    .Q_N(_0071_),
    .Q(\counter.streamer.digits_r[15] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[16]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net212),
    .D(_0183_),
    .Q_N(_1184_),
    .Q(\counter.streamer.digits_r[16] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[17]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net213),
    .D(_0184_),
    .Q_N(_1183_),
    .Q(\counter.streamer.digits_r[17] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[18]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net214),
    .D(_0185_),
    .Q_N(_1182_),
    .Q(\counter.streamer.digits_r[18] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[19]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net215),
    .D(_0186_),
    .Q_N(_1181_),
    .Q(\counter.streamer.digits_r[19] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[1]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net216),
    .D(_0187_),
    .Q_N(_1180_),
    .Q(\counter.streamer.digits_r[1] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[20]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net217),
    .D(_0188_),
    .Q_N(_1179_),
    .Q(\counter.streamer.digits_r[20] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[21]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net218),
    .D(_0189_),
    .Q_N(_1178_),
    .Q(\counter.streamer.digits_r[21] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[22]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net219),
    .D(_0190_),
    .Q_N(_1177_),
    .Q(\counter.streamer.digits_r[22] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[23]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net220),
    .D(_0191_),
    .Q_N(_1176_),
    .Q(\counter.streamer.digits_r[23] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[2]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net221),
    .D(_0192_),
    .Q_N(_1175_),
    .Q(\counter.streamer.digits_r[2] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[3]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net222),
    .D(_0193_),
    .Q_N(_0068_),
    .Q(\counter.streamer.digits_r[3] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[4]$_SDFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net223),
    .D(_0194_),
    .Q_N(_1174_),
    .Q(\counter.streamer.digits_r[4] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[5]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net224),
    .D(_0195_),
    .Q_N(_1173_),
    .Q(\counter.streamer.digits_r[5] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[6]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net225),
    .D(_0196_),
    .Q_N(_1172_),
    .Q(\counter.streamer.digits_r[6] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[7]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net226),
    .D(_0197_),
    .Q_N(_0069_),
    .Q(\counter.streamer.digits_r[7] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[8]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net227),
    .D(_0198_),
    .Q_N(_1171_),
    .Q(\counter.streamer.digits_r[8] ));
 sg13g2_dfrbp_1 \counter.streamer.digits_r[9]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net228),
    .D(_0199_),
    .Q_N(_1170_),
    .Q(\counter.streamer.digits_r[9] ));
 sg13g2_dfrbp_1 \counter.streamer.graphical_decoder.pattern_adg[1]$_SDFF_PP0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net229),
    .D(_0200_),
    .Q_N(_1169_),
    .Q(\counter.streamer.graphical_decoder.pattern_adg[1] ));
 sg13g2_dfrbp_1 \counter.streamer.graphical_decoder.pattern_adg[2]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net230),
    .D(_0201_),
    .Q_N(_0066_),
    .Q(\counter.streamer.graphical_decoder.pattern_adg[2] ));
 sg13g2_dfrbp_1 \counter.streamer.graphical_decoder.pattern_adg[4]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net231),
    .D(_0202_),
    .Q_N(_1168_),
    .Q(\counter.streamer.graphical_decoder.pattern_adg[4] ));
 sg13g2_dfrbp_1 \counter.streamer.graphical_decoder.pattern_adg[6]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net232),
    .D(_0203_),
    .Q_N(_0046_),
    .Q(\counter.streamer.graphical_decoder.pattern_adg[3] ));
 sg13g2_dfrbp_1 \counter.streamer.state_r[0]$_DFF_P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net233),
    .D(net48),
    .Q_N(_1303_),
    .Q(\counter.oled_driver.mc_exec.state_r[0] ));
 sg13g2_dfrbp_1 \counter.streamer.state_r[1]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net234),
    .D(_0030_),
    .Q_N(_1304_),
    .Q(\counter.oled_driver.sync_stb_in ));
 sg13g2_dfrbp_1 \counter.streamer.state_r[2]$_DFF_P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net235),
    .D(_0031_),
    .Q_N(_1305_),
    .Q(\counter.oled_driver.write_stb_in ));
 sg13g2_dfrbp_1 \counter.streamer.state_r[3]$_DFF_P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net236),
    .D(_0032_),
    .Q_N(_1306_),
    .Q(\counter.streamer.ready_out ));
 sg13g2_dfrbp_1 \counter.streamer.state_r[4]$_DFF_P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net237),
    .D(_0014_),
    .Q_N(_1307_),
    .Q(\counter.streamer.state_r[4] ));
 sg13g2_dfrbp_1 \counter.streamer.state_r[5]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net238),
    .D(_0015_),
    .Q_N(_0063_),
    .Q(\counter.streamer.state_r[5] ));
 sg13g2_dfrbp_1 \counter.streamer.x_index_r[0]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net239),
    .D(_0204_),
    .Q_N(_0062_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[0] ));
 sg13g2_dfrbp_1 \counter.streamer.x_index_r[1]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net240),
    .D(_0205_),
    .Q_N(_0045_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[1] ));
 sg13g2_dfrbp_1 \counter.streamer.x_index_r[2]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net241),
    .D(_0206_),
    .Q_N(_0061_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[2] ));
 sg13g2_dfrbp_1 \counter.streamer.x_index_r[3]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net242),
    .D(_0207_),
    .Q_N(_1167_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[3] ));
 sg13g2_dfrbp_1 \counter.streamer.x_index_r[4]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net243),
    .D(_0208_),
    .Q_N(_0060_),
    .Q(\counter.streamer.graphical_decoder.index_x_in[4] ));
 sg13g2_dfrbp_1 \counter.streamer.y_index_r[0]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net244),
    .D(_0209_),
    .Q_N(_0044_),
    .Q(\counter.streamer.graphical_decoder.index_y_in[0] ));
 sg13g2_dfrbp_1 \counter.streamer.y_index_r[1]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net245),
    .D(_0210_),
    .Q_N(_0043_),
    .Q(\counter.streamer.graphical_decoder.index_y_in[1] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout11 (.A(_0417_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_0857_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0861_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_0886_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_0880_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0876_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0862_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0855_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0845_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0240_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0853_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0836_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0233_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0858_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0372_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0349_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0333_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0348_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1153_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0745_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0339_),
    .X(net31));
 sg13g2_buf_4 fanout32 (.X(net32),
    .A(net33));
 sg13g2_buf_4 fanout33 (.X(net33),
    .A(net35));
 sg13g2_buf_2 fanout34 (.A(net35),
    .X(net34));
 sg13g2_buf_4 fanout35 (.X(net35),
    .A(_0073_));
 sg13g2_buf_2 fanout36 (.A(_0744_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0663_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0598_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0593_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0586_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0574_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0367_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0253_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1081_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0993_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0779_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0647_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(\counter.oled_driver.mc_exec.reset_in ),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0594_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0556_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0989_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0875_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0775_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0762_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0759_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0749_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0737_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0735_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0717_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0676_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0673_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0646_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0636_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0767_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0763_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0760_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0757_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0753_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0748_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0736_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0721_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0701_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0668_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0667_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0655_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0649_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0643_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0634_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(net80),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(net82),
    .X(net80));
 sg13g2_buf_1 fanout81 (.A(net82),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(net2),
    .X(net82));
 sg13g2_tielo _2452__83 (.L_LO(net83));
 sg13g2_tielo _2453__84 (.L_LO(net84));
 sg13g2_tielo _2454__85 (.L_LO(net85));
 sg13g2_tielo _2455__86 (.L_LO(net86));
 sg13g2_tielo _2456__87 (.L_LO(net87));
 sg13g2_tielo _2457__88 (.L_LO(net88));
 sg13g2_tielo _2458__89 (.L_LO(net89));
 sg13g2_tielo _2459__90 (.L_LO(net90));
 sg13g2_tielo _2460__91 (.L_LO(net91));
 sg13g2_tielo _2461__92 (.L_LO(net92));
 sg13g2_tielo _2462__93 (.L_LO(net93));
 sg13g2_tielo _2463__94 (.L_LO(net94));
 sg13g2_tielo _2464__95 (.L_LO(net95));
 sg13g2_tielo _2465__96 (.L_LO(net96));
 sg13g2_tielo _2466__97 (.L_LO(net97));
 sg13g2_tielo _2467__98 (.L_LO(net98));
 sg13g2_tiehi _2441__100 (.L_HI(net100));
 sg13g2_tiehi _2442__101 (.L_HI(net101));
 sg13g2_tiehi _2443__102 (.L_HI(net102));
 sg13g2_tiehi _2444__103 (.L_HI(net103));
 sg13g2_tiehi _2445__104 (.L_HI(net104));
 sg13g2_tiehi _2446__105 (.L_HI(net105));
 sg13g2_tiehi _2447__106 (.L_HI(net106));
 sg13g2_tiehi _2448__107 (.L_HI(net107));
 sg13g2_tiehi _2449__108 (.L_HI(net108));
 sg13g2_tiehi \counter.counter_ref.digit_0.digit_out[0]$_SDFFE_PP0P__109  (.L_HI(net109));
 sg13g2_tiehi \counter.counter_ref.digit_0.digit_out[1]$_SDFFE_PP0P__110  (.L_HI(net110));
 sg13g2_tiehi \counter.counter_ref.digit_0.digit_out[2]$_SDFFE_PP0P__111  (.L_HI(net111));
 sg13g2_tiehi \counter.counter_ref.digit_0.digit_out[3]$_SDFFE_PP0P__112  (.L_HI(net112));
 sg13g2_tiehi \counter.counter_ref.genblk1[1].digit_x.digit_out[0]$_SDFFE_PP0P__113  (.L_HI(net113));
 sg13g2_tiehi \counter.counter_ref.genblk1[1].digit_x.digit_out[1]$_SDFFE_PP0P__114  (.L_HI(net114));
 sg13g2_tiehi \counter.counter_ref.genblk1[1].digit_x.digit_out[2]$_SDFFE_PP0P__115  (.L_HI(net115));
 sg13g2_tiehi \counter.counter_ref.genblk1[1].digit_x.digit_out[3]$_SDFFE_PP0P__116  (.L_HI(net116));
 sg13g2_tiehi \counter.counter_ref.genblk1[2].digit_x.digit_out[0]$_SDFFE_PP0P__117  (.L_HI(net117));
 sg13g2_tiehi \counter.counter_ref.genblk1[2].digit_x.digit_out[1]$_SDFFE_PP0P__118  (.L_HI(net118));
 sg13g2_tiehi \counter.counter_ref.genblk1[2].digit_x.digit_out[2]$_SDFFE_PP0P__119  (.L_HI(net119));
 sg13g2_tiehi \counter.counter_ref.genblk1[2].digit_x.digit_out[3]$_SDFFE_PP0P__120  (.L_HI(net120));
 sg13g2_tiehi \counter.counter_ref.genblk1[3].digit_x.digit_out[0]$_SDFFE_PP0P__121  (.L_HI(net121));
 sg13g2_tiehi \counter.counter_ref.genblk1[3].digit_x.digit_out[1]$_SDFFE_PP0P__122  (.L_HI(net122));
 sg13g2_tiehi \counter.counter_ref.genblk1[3].digit_x.digit_out[2]$_SDFFE_PP0P__123  (.L_HI(net123));
 sg13g2_tiehi \counter.counter_ref.genblk1[3].digit_x.digit_out[3]$_SDFFE_PP0P__124  (.L_HI(net124));
 sg13g2_tiehi \counter.counter_ref.genblk1[4].digit_x.digit_out[0]$_SDFFE_PP0P__125  (.L_HI(net125));
 sg13g2_tiehi \counter.counter_ref.genblk1[4].digit_x.digit_out[1]$_SDFFE_PP0P__126  (.L_HI(net126));
 sg13g2_tiehi \counter.counter_ref.genblk1[4].digit_x.digit_out[2]$_SDFFE_PP0P__127  (.L_HI(net127));
 sg13g2_tiehi \counter.counter_ref.genblk1[4].digit_x.digit_out[3]$_SDFFE_PP0P__128  (.L_HI(net128));
 sg13g2_tiehi \counter.counter_ref.genblk1[5].digit_x.digit_out[0]$_SDFFE_PP0P__129  (.L_HI(net129));
 sg13g2_tiehi \counter.counter_ref.genblk1[5].digit_x.digit_out[1]$_SDFFE_PP0P__130  (.L_HI(net130));
 sg13g2_tiehi \counter.counter_ref.genblk1[5].digit_x.digit_out[2]$_SDFFE_PP0P__131  (.L_HI(net131));
 sg13g2_tiehi \counter.counter_ref.genblk1[5].digit_x.digit_out[3]$_SDFFE_PP0P__132  (.L_HI(net132));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[0]$_SDFFE_PN0P__133  (.L_HI(net133));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[10]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[11]$_SDFFE_PN0P__135  (.L_HI(net135));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[12]$_SDFFE_PN0P__136  (.L_HI(net136));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[13]$_SDFFE_PN0P__137  (.L_HI(net137));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[14]$_SDFFE_PN0P__138  (.L_HI(net138));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[15]$_SDFFE_PN0P__139  (.L_HI(net139));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[16]$_SDFFE_PN0P__140  (.L_HI(net140));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[1]$_SDFFE_PN0P__141  (.L_HI(net141));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[2]$_SDFFE_PN0P__142  (.L_HI(net142));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[3]$_SDFFE_PN0P__143  (.L_HI(net143));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[4]$_SDFFE_PN0P__144  (.L_HI(net144));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[5]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[6]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[7]$_SDFFE_PN0P__147  (.L_HI(net147));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[8]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \counter.oled_driver.mc_exec.delay_cnt[9]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \counter.oled_driver.mc_exec.oled_dc_out$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \counter.oled_driver.mc_exec.oled_rstn_out$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \counter.oled_driver.mc_exec.oled_vbatn_out$_SDFFE_PN1P__152  (.L_HI(net152));
 sg13g2_tiehi \counter.oled_driver.mc_exec.oled_vcdn_out$_SDFFE_PN1P__153  (.L_HI(net153));
 sg13g2_tiehi \counter.oled_driver.mc_exec.rom_index_r[0]$_SDFFE_PN0N__154  (.L_HI(net154));
 sg13g2_tiehi \counter.oled_driver.mc_exec.rom_index_r[1]$_SDFFE_PN0N__155  (.L_HI(net155));
 sg13g2_tiehi \counter.oled_driver.mc_exec.rom_index_r[2]$_SDFFE_PN0N__156  (.L_HI(net156));
 sg13g2_tiehi \counter.oled_driver.mc_exec.rom_index_r[3]$_SDFFE_PN0N__157  (.L_HI(net157));
 sg13g2_tiehi \counter.oled_driver.mc_exec.rom_index_r[4]$_SDFFE_PN0N__158  (.L_HI(net158));
 sg13g2_tiehi \counter.oled_driver.mc_exec.rom_index_r[5]$_SDFFE_PN0N__159  (.L_HI(net159));
 sg13g2_tiehi \counter.oled_driver.mc_exec.state_r[1]$_DFF_P__160  (.L_HI(net160));
 sg13g2_tiehi \counter.oled_driver.mc_exec.state_r[2]$_DFF_P__161  (.L_HI(net161));
 sg13g2_tiehi \counter.oled_driver.mc_exec.state_r[3]$_DFF_P__162  (.L_HI(net162));
 sg13g2_tiehi \counter.oled_driver.mc_exec.state_r[4]$_DFF_P__163  (.L_HI(net163));
 sg13g2_tiehi \counter.oled_driver.mc_exec.state_r[5]$_DFF_P__164  (.L_HI(net164));
 sg13g2_tiehi \counter.oled_driver.mc_exec.state_r[6]$_DFF_P__165  (.L_HI(net165));
 sg13g2_tiehi \counter.oled_driver.mc_procedure_offset[0]$_SDFFE_PN0P__166  (.L_HI(net166));
 sg13g2_tiehi \counter.oled_driver.spi_data[0]$_SDFFE_PN0P__167  (.L_HI(net167));
 sg13g2_tiehi \counter.oled_driver.spi_data[1]$_SDFFE_PN0P__168  (.L_HI(net168));
 sg13g2_tiehi \counter.oled_driver.spi_data[2]$_SDFFE_PN0P__169  (.L_HI(net169));
 sg13g2_tiehi \counter.oled_driver.spi_data[3]$_SDFFE_PN0P__170  (.L_HI(net170));
 sg13g2_tiehi \counter.oled_driver.spi_data[4]$_SDFFE_PN0P__171  (.L_HI(net171));
 sg13g2_tiehi \counter.oled_driver.spi_data[5]$_SDFFE_PN0P__172  (.L_HI(net172));
 sg13g2_tiehi \counter.oled_driver.spi_data[6]$_SDFFE_PN0P__173  (.L_HI(net173));
 sg13g2_tiehi \counter.oled_driver.spi_data[7]$_SDFFE_PN0P__174  (.L_HI(net174));
 sg13g2_tiehi \counter.oled_driver.spi_driver.chip_select_r$_SDFFE_PN1P__175  (.L_HI(net175));
 sg13g2_tiehi \counter.oled_driver.spi_driver.deactivate_cs_r$_SDFFE_PN0P__176  (.L_HI(net176));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[0]$_SDFFE_PP0P__177  (.L_HI(net177));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[1]$_SDFFE_PP0P__178  (.L_HI(net178));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[2]$_SDFFE_PP0P__179  (.L_HI(net179));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.bit_counter_r[3]$_SDFFE_PP0P__180  (.L_HI(net180));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[0]$_SDFFE_PN0P__181  (.L_HI(net181));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[1]$_SDFFE_PN0P__182  (.L_HI(net182));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[2]$_SDFFE_PN0P__183  (.L_HI(net183));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[3]$_SDFFE_PN0P__184  (.L_HI(net184));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[4]$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[5]$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[6]$_SDFFE_PN0P__187  (.L_HI(net187));
 sg13g2_tiehi \counter.oled_driver.spi_driver.shift_reg.shadow_reg_r[7]$_SDFFE_PN0P__188  (.L_HI(net188));
 sg13g2_tiehi \counter.oled_driver.spi_driver.state_r[0]$_DFF_P__189  (.L_HI(net189));
 sg13g2_tiehi \counter.oled_driver.spi_driver.state_r[1]$_DFF_P__190  (.L_HI(net190));
 sg13g2_tiehi \counter.oled_driver.spi_driver.state_r[2]$_DFF_P__191  (.L_HI(net191));
 sg13g2_tiehi \counter.oled_driver.state_r[0]$_DFF_P__192  (.L_HI(net192));
 sg13g2_tiehi \counter.oled_driver.state_r[1]$_DFF_P__193  (.L_HI(net193));
 sg13g2_tiehi \counter.oled_driver.state_r[2]$_DFF_P__194  (.L_HI(net194));
 sg13g2_tiehi \counter.oled_driver.state_r[3]$_DFF_P__195  (.L_HI(net195));
 sg13g2_tiehi \counter.oled_driver.state_r[4]$_DFF_P__196  (.L_HI(net196));
 sg13g2_tiehi \counter.oled_driver.state_r[5]$_DFF_P__197  (.L_HI(net197));
 sg13g2_tiehi \counter.refresh_display$_SDFFE_PN0P__198  (.L_HI(net198));
 sg13g2_tiehi \counter.state[0]$_DFF_P__199  (.L_HI(net199));
 sg13g2_tiehi \counter.state[1]$_DFF_P__200  (.L_HI(net200));
 sg13g2_tiehi \counter.state[2]$_DFF_P__201  (.L_HI(net201));
 sg13g2_tiehi \counter.streamer.digit_cnt_r[0]$_SDFFE_PN1P__202  (.L_HI(net202));
 sg13g2_tiehi \counter.streamer.digit_cnt_r[1]$_SDFFE_PN0P__203  (.L_HI(net203));
 sg13g2_tiehi \counter.streamer.digit_cnt_r[2]$_SDFFE_PN1P__204  (.L_HI(net204));
 sg13g2_tiehi \counter.streamer.digits_r[0]$_SDFFE_PN0P__205  (.L_HI(net205));
 sg13g2_tiehi \counter.streamer.digits_r[10]$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \counter.streamer.digits_r[11]$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_tiehi \counter.streamer.digits_r[12]$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \counter.streamer.digits_r[13]$_SDFFE_PN0P__209  (.L_HI(net209));
 sg13g2_tiehi \counter.streamer.digits_r[14]$_SDFFE_PN0P__210  (.L_HI(net210));
 sg13g2_tiehi \counter.streamer.digits_r[15]$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \counter.streamer.digits_r[16]$_SDFFE_PN0P__212  (.L_HI(net212));
 sg13g2_tiehi \counter.streamer.digits_r[17]$_SDFFE_PN0P__213  (.L_HI(net213));
 sg13g2_tiehi \counter.streamer.digits_r[18]$_SDFFE_PN0P__214  (.L_HI(net214));
 sg13g2_tiehi \counter.streamer.digits_r[19]$_SDFFE_PN0P__215  (.L_HI(net215));
 sg13g2_tiehi \counter.streamer.digits_r[1]$_SDFFE_PN0P__216  (.L_HI(net216));
 sg13g2_tiehi \counter.streamer.digits_r[20]$_SDFFE_PN0P__217  (.L_HI(net217));
 sg13g2_tiehi \counter.streamer.digits_r[21]$_SDFFE_PN0P__218  (.L_HI(net218));
 sg13g2_tiehi \counter.streamer.digits_r[22]$_SDFFE_PN0P__219  (.L_HI(net219));
 sg13g2_tiehi \counter.streamer.digits_r[23]$_SDFFE_PN0P__220  (.L_HI(net220));
 sg13g2_tiehi \counter.streamer.digits_r[2]$_SDFFE_PN0P__221  (.L_HI(net221));
 sg13g2_tiehi \counter.streamer.digits_r[3]$_SDFFE_PN0P__222  (.L_HI(net222));
 sg13g2_tiehi \counter.streamer.digits_r[4]$_SDFFE_PN0P__223  (.L_HI(net223));
 sg13g2_tiehi \counter.streamer.digits_r[5]$_SDFFE_PN0P__224  (.L_HI(net224));
 sg13g2_tiehi \counter.streamer.digits_r[6]$_SDFFE_PN0P__225  (.L_HI(net225));
 sg13g2_tiehi \counter.streamer.digits_r[7]$_SDFFE_PN0P__226  (.L_HI(net226));
 sg13g2_tiehi \counter.streamer.digits_r[8]$_SDFFE_PN0P__227  (.L_HI(net227));
 sg13g2_tiehi \counter.streamer.digits_r[9]$_SDFFE_PN0P__228  (.L_HI(net228));
 sg13g2_tiehi \counter.streamer.graphical_decoder.pattern_adg[1]$_SDFF_PP0__229  (.L_HI(net229));
 sg13g2_tiehi \counter.streamer.graphical_decoder.pattern_adg[2]$_SDFF_PP0__230  (.L_HI(net230));
 sg13g2_tiehi \counter.streamer.graphical_decoder.pattern_adg[4]$_SDFF_PP0__231  (.L_HI(net231));
 sg13g2_tiehi \counter.streamer.graphical_decoder.pattern_adg[6]$_SDFF_PP0__232  (.L_HI(net232));
 sg13g2_tiehi \counter.streamer.state_r[0]$_DFF_P__233  (.L_HI(net233));
 sg13g2_tiehi \counter.streamer.state_r[1]$_DFF_P__234  (.L_HI(net234));
 sg13g2_tiehi \counter.streamer.state_r[2]$_DFF_P__235  (.L_HI(net235));
 sg13g2_tiehi \counter.streamer.state_r[3]$_DFF_P__236  (.L_HI(net236));
 sg13g2_tiehi \counter.streamer.state_r[4]$_DFF_P__237  (.L_HI(net237));
 sg13g2_tiehi \counter.streamer.state_r[5]$_DFF_P__238  (.L_HI(net238));
 sg13g2_tiehi \counter.streamer.x_index_r[0]$_SDFFE_PN0P__239  (.L_HI(net239));
 sg13g2_tiehi \counter.streamer.x_index_r[1]$_SDFFE_PN0P__240  (.L_HI(net240));
 sg13g2_tiehi \counter.streamer.x_index_r[2]$_SDFFE_PN0P__241  (.L_HI(net241));
 sg13g2_tiehi \counter.streamer.x_index_r[3]$_SDFFE_PN0P__242  (.L_HI(net242));
 sg13g2_tiehi \counter.streamer.x_index_r[4]$_SDFFE_PN0P__243  (.L_HI(net243));
 sg13g2_tiehi \counter.streamer.y_index_r[0]$_SDFFE_PN0P__244  (.L_HI(net244));
 sg13g2_tiehi \counter.streamer.y_index_r[1]$_SDFFE_PN0P__245  (.L_HI(net245));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_31__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_fill_2 FILLER_11_427 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_fill_2 FILLER_15_427 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_4 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_decap_8 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_16_415 ();
 sg13g2_decap_8 FILLER_16_422 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_fill_2 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_237 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_fill_2 FILLER_18_224 ();
 sg13g2_fill_2 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_fill_1 FILLER_18_284 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_295 ();
 sg13g2_decap_4 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_8 FILLER_18_356 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_8 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_18_412 ();
 sg13g2_decap_8 FILLER_18_419 ();
 sg13g2_decap_4 FILLER_18_426 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_4 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_257 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_fill_2 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_224 ();
 sg13g2_decap_4 FILLER_20_229 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_fill_1 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_fill_1 FILLER_20_282 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_decap_8 FILLER_20_309 ();
 sg13g2_decap_8 FILLER_20_316 ();
 sg13g2_decap_8 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_330 ();
 sg13g2_decap_8 FILLER_20_337 ();
 sg13g2_decap_8 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_decap_8 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_20_414 ();
 sg13g2_decap_8 FILLER_20_421 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_fill_1 FILLER_21_254 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_1 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_4 FILLER_22_217 ();
 sg13g2_decap_4 FILLER_22_262 ();
 sg13g2_fill_1 FILLER_22_270 ();
 sg13g2_fill_2 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_decap_4 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_314 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_8 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_22_412 ();
 sg13g2_decap_8 FILLER_22_419 ();
 sg13g2_decap_4 FILLER_22_426 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_4 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_255 ();
 sg13g2_decap_8 FILLER_23_260 ();
 sg13g2_decap_8 FILLER_23_267 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_282 ();
 sg13g2_fill_1 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_314 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_fill_2 FILLER_23_342 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_decap_8 FILLER_23_391 ();
 sg13g2_decap_8 FILLER_23_398 ();
 sg13g2_decap_8 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_23_412 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_decap_4 FILLER_23_426 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_fill_2 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_237 ();
 sg13g2_decap_4 FILLER_24_244 ();
 sg13g2_fill_2 FILLER_24_248 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_268 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_fill_2 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_8 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_24_412 ();
 sg13g2_decap_8 FILLER_24_419 ();
 sg13g2_decap_4 FILLER_24_426 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_fill_2 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_fill_2 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_fill_1 FILLER_25_285 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_fill_1 FILLER_25_299 ();
 sg13g2_fill_2 FILLER_25_304 ();
 sg13g2_decap_8 FILLER_25_310 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_324 ();
 sg13g2_decap_4 FILLER_25_331 ();
 sg13g2_fill_2 FILLER_25_348 ();
 sg13g2_decap_8 FILLER_25_381 ();
 sg13g2_decap_8 FILLER_25_388 ();
 sg13g2_decap_8 FILLER_25_395 ();
 sg13g2_decap_8 FILLER_25_402 ();
 sg13g2_decap_8 FILLER_25_409 ();
 sg13g2_decap_8 FILLER_25_416 ();
 sg13g2_decap_8 FILLER_25_423 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_4 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_decap_4 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_238 ();
 sg13g2_decap_4 FILLER_26_247 ();
 sg13g2_fill_2 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_261 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_4 FILLER_26_280 ();
 sg13g2_fill_2 FILLER_26_293 ();
 sg13g2_decap_4 FILLER_26_306 ();
 sg13g2_decap_4 FILLER_26_336 ();
 sg13g2_fill_1 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_8 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_decap_8 FILLER_26_417 ();
 sg13g2_decap_4 FILLER_26_424 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_fill_2 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_decap_8 FILLER_27_334 ();
 sg13g2_fill_2 FILLER_27_341 ();
 sg13g2_fill_1 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_decap_4 FILLER_27_359 ();
 sg13g2_fill_1 FILLER_27_363 ();
 sg13g2_decap_4 FILLER_27_372 ();
 sg13g2_fill_2 FILLER_27_376 ();
 sg13g2_decap_8 FILLER_27_404 ();
 sg13g2_decap_8 FILLER_27_411 ();
 sg13g2_decap_8 FILLER_27_418 ();
 sg13g2_decap_4 FILLER_27_425 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_173 ();
 sg13g2_decap_4 FILLER_28_180 ();
 sg13g2_decap_8 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_237 ();
 sg13g2_fill_2 FILLER_28_251 ();
 sg13g2_decap_8 FILLER_28_275 ();
 sg13g2_decap_4 FILLER_28_282 ();
 sg13g2_fill_2 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_293 ();
 sg13g2_decap_8 FILLER_28_303 ();
 sg13g2_decap_4 FILLER_28_310 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_fill_1 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_352 ();
 sg13g2_fill_1 FILLER_28_354 ();
 sg13g2_fill_2 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_407 ();
 sg13g2_decap_4 FILLER_28_414 ();
 sg13g2_fill_1 FILLER_28_418 ();
 sg13g2_decap_4 FILLER_28_424 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_4 FILLER_29_133 ();
 sg13g2_fill_2 FILLER_29_168 ();
 sg13g2_fill_1 FILLER_29_170 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_decap_4 FILLER_29_191 ();
 sg13g2_decap_4 FILLER_29_220 ();
 sg13g2_decap_4 FILLER_29_229 ();
 sg13g2_decap_4 FILLER_29_237 ();
 sg13g2_fill_2 FILLER_29_241 ();
 sg13g2_fill_1 FILLER_29_262 ();
 sg13g2_decap_8 FILLER_29_269 ();
 sg13g2_decap_8 FILLER_29_276 ();
 sg13g2_decap_4 FILLER_29_283 ();
 sg13g2_fill_2 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_4 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_decap_4 FILLER_29_330 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_369 ();
 sg13g2_decap_4 FILLER_29_379 ();
 sg13g2_fill_1 FILLER_29_383 ();
 sg13g2_fill_1 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_4 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_208 ();
 sg13g2_decap_4 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_264 ();
 sg13g2_decap_8 FILLER_30_271 ();
 sg13g2_decap_4 FILLER_30_278 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_fill_1 FILLER_30_298 ();
 sg13g2_decap_4 FILLER_30_304 ();
 sg13g2_fill_2 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_349 ();
 sg13g2_decap_8 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_30_363 ();
 sg13g2_decap_8 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_377 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_fill_1 FILLER_30_409 ();
 sg13g2_fill_1 FILLER_30_415 ();
 sg13g2_decap_8 FILLER_30_421 ();
 sg13g2_fill_2 FILLER_30_428 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_4 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_decap_4 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_decap_4 FILLER_31_215 ();
 sg13g2_fill_1 FILLER_31_219 ();
 sg13g2_decap_4 FILLER_31_250 ();
 sg13g2_fill_1 FILLER_31_254 ();
 sg13g2_decap_4 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_321 ();
 sg13g2_fill_1 FILLER_31_323 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_fill_2 FILLER_31_395 ();
 sg13g2_fill_1 FILLER_31_397 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_4 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_158 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_fill_2 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_fill_2 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_4 FILLER_32_256 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_295 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_decap_8 FILLER_32_311 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_4 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_4 FILLER_32_357 ();
 sg13g2_fill_1 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_414 ();
 sg13g2_decap_8 FILLER_32_421 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_fill_2 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_160 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_decap_8 FILLER_33_218 ();
 sg13g2_decap_4 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_decap_8 FILLER_33_237 ();
 sg13g2_decap_8 FILLER_33_244 ();
 sg13g2_decap_8 FILLER_33_251 ();
 sg13g2_decap_4 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_262 ();
 sg13g2_decap_4 FILLER_33_275 ();
 sg13g2_fill_2 FILLER_33_299 ();
 sg13g2_decap_8 FILLER_33_309 ();
 sg13g2_decap_8 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_323 ();
 sg13g2_decap_8 FILLER_33_330 ();
 sg13g2_decap_8 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_357 ();
 sg13g2_decap_4 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_371 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_1 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_4 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_176 ();
 sg13g2_fill_2 FILLER_34_183 ();
 sg13g2_decap_8 FILLER_34_198 ();
 sg13g2_fill_2 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_decap_8 FILLER_34_219 ();
 sg13g2_decap_8 FILLER_34_226 ();
 sg13g2_decap_4 FILLER_34_241 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_264 ();
 sg13g2_decap_4 FILLER_34_271 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_285 ();
 sg13g2_fill_2 FILLER_34_290 ();
 sg13g2_fill_1 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_296 ();
 sg13g2_decap_8 FILLER_34_303 ();
 sg13g2_decap_8 FILLER_34_310 ();
 sg13g2_fill_2 FILLER_34_317 ();
 sg13g2_decap_4 FILLER_34_397 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_4 FILLER_35_203 ();
 sg13g2_decap_4 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_271 ();
 sg13g2_decap_4 FILLER_35_278 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_291 ();
 sg13g2_decap_4 FILLER_35_298 ();
 sg13g2_fill_1 FILLER_35_302 ();
 sg13g2_decap_8 FILLER_35_337 ();
 sg13g2_fill_2 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_346 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_2 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_414 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_decap_4 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_decap_8 FILLER_36_181 ();
 sg13g2_decap_4 FILLER_36_188 ();
 sg13g2_fill_2 FILLER_36_192 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_decap_4 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_decap_4 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_349 ();
 sg13g2_decap_4 FILLER_36_356 ();
 sg13g2_fill_1 FILLER_36_360 ();
 sg13g2_decap_4 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_370 ();
 sg13g2_decap_8 FILLER_36_379 ();
 sg13g2_fill_2 FILLER_36_386 ();
 sg13g2_fill_1 FILLER_36_388 ();
 sg13g2_decap_4 FILLER_36_394 ();
 sg13g2_fill_1 FILLER_36_402 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_decap_4 FILLER_37_221 ();
 sg13g2_fill_2 FILLER_37_225 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_fill_1 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_282 ();
 sg13g2_fill_2 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_295 ();
 sg13g2_fill_1 FILLER_37_297 ();
 sg13g2_fill_2 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_4 FILLER_37_333 ();
 sg13g2_fill_1 FILLER_37_337 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_4 FILLER_37_386 ();
 sg13g2_fill_1 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_decap_8 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_4 FILLER_38_161 ();
 sg13g2_fill_2 FILLER_38_165 ();
 sg13g2_fill_1 FILLER_38_209 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_fill_2 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_246 ();
 sg13g2_fill_1 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_280 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_decap_4 FILLER_38_293 ();
 sg13g2_decap_4 FILLER_38_301 ();
 sg13g2_fill_1 FILLER_38_305 ();
 sg13g2_decap_4 FILLER_38_311 ();
 sg13g2_fill_1 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_fill_2 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_4 FILLER_38_364 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_fill_2 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_403 ();
 sg13g2_decap_8 FILLER_38_412 ();
 sg13g2_decap_8 FILLER_38_419 ();
 sg13g2_decap_4 FILLER_38_426 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_fill_2 FILLER_39_140 ();
 sg13g2_fill_1 FILLER_39_142 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_fill_2 FILLER_39_168 ();
 sg13g2_fill_1 FILLER_39_170 ();
 sg13g2_fill_1 FILLER_39_176 ();
 sg13g2_decap_4 FILLER_39_185 ();
 sg13g2_fill_1 FILLER_39_195 ();
 sg13g2_fill_1 FILLER_39_201 ();
 sg13g2_decap_4 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_225 ();
 sg13g2_decap_8 FILLER_39_232 ();
 sg13g2_decap_8 FILLER_39_239 ();
 sg13g2_decap_8 FILLER_39_246 ();
 sg13g2_decap_8 FILLER_39_253 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_decap_8 FILLER_39_271 ();
 sg13g2_decap_4 FILLER_39_278 ();
 sg13g2_fill_2 FILLER_39_288 ();
 sg13g2_fill_1 FILLER_39_290 ();
 sg13g2_decap_8 FILLER_39_298 ();
 sg13g2_fill_1 FILLER_39_305 ();
 sg13g2_fill_2 FILLER_39_354 ();
 sg13g2_fill_1 FILLER_39_356 ();
 sg13g2_decap_8 FILLER_39_361 ();
 sg13g2_decap_8 FILLER_39_368 ();
 sg13g2_decap_8 FILLER_39_375 ();
 sg13g2_decap_8 FILLER_39_382 ();
 sg13g2_fill_1 FILLER_39_389 ();
 sg13g2_fill_1 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_237 ();
 sg13g2_decap_8 FILLER_40_244 ();
 sg13g2_fill_2 FILLER_40_251 ();
 sg13g2_decap_8 FILLER_40_257 ();
 sg13g2_fill_1 FILLER_40_264 ();
 sg13g2_decap_8 FILLER_40_300 ();
 sg13g2_fill_1 FILLER_40_312 ();
 sg13g2_fill_1 FILLER_40_317 ();
 sg13g2_fill_1 FILLER_40_344 ();
 sg13g2_fill_1 FILLER_40_371 ();
 sg13g2_fill_2 FILLER_40_402 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_fill_1 FILLER_41_154 ();
 sg13g2_fill_1 FILLER_41_185 ();
 sg13g2_fill_1 FILLER_41_192 ();
 sg13g2_fill_2 FILLER_41_201 ();
 sg13g2_fill_2 FILLER_41_207 ();
 sg13g2_fill_1 FILLER_41_209 ();
 sg13g2_decap_8 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_222 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_4 FILLER_41_287 ();
 sg13g2_fill_1 FILLER_41_291 ();
 sg13g2_decap_8 FILLER_41_304 ();
 sg13g2_fill_2 FILLER_41_311 ();
 sg13g2_fill_1 FILLER_41_313 ();
 sg13g2_decap_8 FILLER_41_326 ();
 sg13g2_decap_8 FILLER_41_333 ();
 sg13g2_decap_4 FILLER_41_387 ();
 sg13g2_fill_2 FILLER_41_391 ();
 sg13g2_fill_2 FILLER_41_398 ();
 sg13g2_decap_4 FILLER_41_417 ();
 sg13g2_decap_4 FILLER_41_425 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_4 FILLER_42_154 ();
 sg13g2_fill_1 FILLER_42_188 ();
 sg13g2_fill_1 FILLER_42_194 ();
 sg13g2_fill_1 FILLER_42_205 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_fill_1 FILLER_42_231 ();
 sg13g2_fill_1 FILLER_42_236 ();
 sg13g2_fill_2 FILLER_42_257 ();
 sg13g2_fill_1 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_264 ();
 sg13g2_decap_8 FILLER_42_271 ();
 sg13g2_decap_8 FILLER_42_278 ();
 sg13g2_fill_1 FILLER_42_285 ();
 sg13g2_fill_2 FILLER_42_293 ();
 sg13g2_fill_1 FILLER_42_295 ();
 sg13g2_fill_2 FILLER_42_301 ();
 sg13g2_decap_4 FILLER_42_307 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_decap_8 FILLER_42_327 ();
 sg13g2_decap_4 FILLER_42_339 ();
 sg13g2_fill_1 FILLER_42_343 ();
 sg13g2_fill_2 FILLER_42_349 ();
 sg13g2_fill_2 FILLER_42_360 ();
 sg13g2_fill_1 FILLER_42_362 ();
 sg13g2_fill_1 FILLER_42_367 ();
 sg13g2_fill_1 FILLER_42_378 ();
 sg13g2_fill_1 FILLER_42_393 ();
 sg13g2_decap_4 FILLER_42_399 ();
 sg13g2_fill_1 FILLER_42_403 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_fill_2 FILLER_43_119 ();
 sg13g2_decap_4 FILLER_43_147 ();
 sg13g2_fill_2 FILLER_43_151 ();
 sg13g2_decap_4 FILLER_43_160 ();
 sg13g2_fill_2 FILLER_43_164 ();
 sg13g2_fill_2 FILLER_43_170 ();
 sg13g2_decap_4 FILLER_43_176 ();
 sg13g2_fill_2 FILLER_43_180 ();
 sg13g2_fill_1 FILLER_43_194 ();
 sg13g2_fill_1 FILLER_43_218 ();
 sg13g2_fill_2 FILLER_43_223 ();
 sg13g2_fill_1 FILLER_43_225 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_fill_1 FILLER_43_252 ();
 sg13g2_decap_4 FILLER_43_268 ();
 sg13g2_fill_2 FILLER_43_272 ();
 sg13g2_decap_8 FILLER_43_304 ();
 sg13g2_fill_2 FILLER_43_311 ();
 sg13g2_fill_1 FILLER_43_313 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_fill_1 FILLER_43_343 ();
 sg13g2_decap_4 FILLER_43_353 ();
 sg13g2_fill_1 FILLER_43_361 ();
 sg13g2_decap_4 FILLER_43_369 ();
 sg13g2_decap_4 FILLER_43_377 ();
 sg13g2_decap_8 FILLER_43_407 ();
 sg13g2_fill_1 FILLER_43_426 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_fill_2 FILLER_44_126 ();
 sg13g2_fill_1 FILLER_44_128 ();
 sg13g2_decap_4 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_167 ();
 sg13g2_decap_8 FILLER_44_174 ();
 sg13g2_decap_8 FILLER_44_181 ();
 sg13g2_decap_4 FILLER_44_193 ();
 sg13g2_fill_1 FILLER_44_210 ();
 sg13g2_fill_2 FILLER_44_237 ();
 sg13g2_fill_1 FILLER_44_244 ();
 sg13g2_fill_1 FILLER_44_250 ();
 sg13g2_fill_1 FILLER_44_265 ();
 sg13g2_decap_8 FILLER_44_271 ();
 sg13g2_decap_8 FILLER_44_278 ();
 sg13g2_fill_1 FILLER_44_285 ();
 sg13g2_fill_2 FILLER_44_290 ();
 sg13g2_fill_1 FILLER_44_292 ();
 sg13g2_decap_8 FILLER_44_298 ();
 sg13g2_decap_8 FILLER_44_305 ();
 sg13g2_fill_1 FILLER_44_312 ();
 sg13g2_decap_4 FILLER_44_328 ();
 sg13g2_fill_2 FILLER_44_332 ();
 sg13g2_fill_2 FILLER_44_339 ();
 sg13g2_fill_1 FILLER_44_341 ();
 sg13g2_fill_1 FILLER_44_368 ();
 sg13g2_decap_8 FILLER_44_373 ();
 sg13g2_decap_8 FILLER_44_380 ();
 sg13g2_decap_8 FILLER_44_387 ();
 sg13g2_fill_2 FILLER_44_394 ();
 sg13g2_fill_1 FILLER_44_396 ();
 sg13g2_decap_4 FILLER_44_401 ();
 sg13g2_fill_2 FILLER_44_405 ();
 sg13g2_fill_2 FILLER_44_428 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_4 FILLER_45_98 ();
 sg13g2_fill_1 FILLER_45_102 ();
 sg13g2_decap_4 FILLER_45_138 ();
 sg13g2_fill_1 FILLER_45_142 ();
 sg13g2_decap_4 FILLER_45_160 ();
 sg13g2_decap_4 FILLER_45_168 ();
 sg13g2_fill_2 FILLER_45_172 ();
 sg13g2_decap_8 FILLER_45_179 ();
 sg13g2_decap_8 FILLER_45_186 ();
 sg13g2_fill_2 FILLER_45_193 ();
 sg13g2_fill_1 FILLER_45_195 ();
 sg13g2_decap_4 FILLER_45_204 ();
 sg13g2_fill_2 FILLER_45_208 ();
 sg13g2_fill_1 FILLER_45_215 ();
 sg13g2_fill_2 FILLER_45_255 ();
 sg13g2_fill_1 FILLER_45_257 ();
 sg13g2_decap_8 FILLER_45_284 ();
 sg13g2_decap_4 FILLER_45_291 ();
 sg13g2_decap_8 FILLER_45_304 ();
 sg13g2_decap_4 FILLER_45_311 ();
 sg13g2_fill_2 FILLER_45_315 ();
 sg13g2_fill_2 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_fill_2 FILLER_45_357 ();
 sg13g2_fill_2 FILLER_45_363 ();
 sg13g2_fill_2 FILLER_45_370 ();
 sg13g2_fill_2 FILLER_45_382 ();
 sg13g2_fill_1 FILLER_45_384 ();
 sg13g2_decap_4 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_fill_2 FILLER_45_427 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_4 FILLER_46_105 ();
 sg13g2_fill_2 FILLER_46_109 ();
 sg13g2_decap_8 FILLER_46_115 ();
 sg13g2_decap_4 FILLER_46_125 ();
 sg13g2_fill_1 FILLER_46_129 ();
 sg13g2_decap_4 FILLER_46_135 ();
 sg13g2_fill_2 FILLER_46_139 ();
 sg13g2_decap_8 FILLER_46_146 ();
 sg13g2_fill_2 FILLER_46_153 ();
 sg13g2_fill_2 FILLER_46_211 ();
 sg13g2_decap_4 FILLER_46_225 ();
 sg13g2_fill_1 FILLER_46_229 ();
 sg13g2_fill_2 FILLER_46_234 ();
 sg13g2_decap_8 FILLER_46_251 ();
 sg13g2_decap_8 FILLER_46_258 ();
 sg13g2_fill_1 FILLER_46_265 ();
 sg13g2_decap_8 FILLER_46_278 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_fill_1 FILLER_46_287 ();
 sg13g2_fill_1 FILLER_46_318 ();
 sg13g2_fill_1 FILLER_46_345 ();
 sg13g2_fill_1 FILLER_46_351 ();
 sg13g2_decap_8 FILLER_46_409 ();
 sg13g2_decap_8 FILLER_46_416 ();
 sg13g2_decap_8 FILLER_46_423 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_167 ();
 sg13g2_decap_8 FILLER_47_174 ();
 sg13g2_decap_8 FILLER_47_181 ();
 sg13g2_decap_8 FILLER_47_192 ();
 sg13g2_fill_1 FILLER_47_199 ();
 sg13g2_decap_8 FILLER_47_211 ();
 sg13g2_fill_1 FILLER_47_218 ();
 sg13g2_decap_8 FILLER_47_223 ();
 sg13g2_decap_8 FILLER_47_230 ();
 sg13g2_decap_8 FILLER_47_237 ();
 sg13g2_decap_8 FILLER_47_244 ();
 sg13g2_decap_8 FILLER_47_251 ();
 sg13g2_decap_4 FILLER_47_258 ();
 sg13g2_decap_8 FILLER_47_296 ();
 sg13g2_decap_4 FILLER_47_303 ();
 sg13g2_fill_1 FILLER_47_307 ();
 sg13g2_decap_8 FILLER_47_324 ();
 sg13g2_decap_8 FILLER_47_331 ();
 sg13g2_decap_4 FILLER_47_342 ();
 sg13g2_decap_8 FILLER_47_355 ();
 sg13g2_decap_4 FILLER_47_362 ();
 sg13g2_fill_1 FILLER_47_366 ();
 sg13g2_decap_4 FILLER_47_389 ();
 sg13g2_decap_4 FILLER_47_398 ();
 sg13g2_fill_2 FILLER_47_402 ();
 sg13g2_decap_4 FILLER_47_408 ();
 sg13g2_fill_1 FILLER_47_412 ();
 sg13g2_decap_8 FILLER_47_417 ();
 sg13g2_decap_4 FILLER_47_424 ();
 sg13g2_fill_2 FILLER_47_428 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_fill_1 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_143 ();
 sg13g2_fill_1 FILLER_48_150 ();
 sg13g2_decap_8 FILLER_48_165 ();
 sg13g2_decap_8 FILLER_48_172 ();
 sg13g2_fill_1 FILLER_48_179 ();
 sg13g2_decap_8 FILLER_48_183 ();
 sg13g2_decap_8 FILLER_48_190 ();
 sg13g2_decap_4 FILLER_48_197 ();
 sg13g2_fill_1 FILLER_48_201 ();
 sg13g2_fill_1 FILLER_48_206 ();
 sg13g2_decap_4 FILLER_48_216 ();
 sg13g2_fill_1 FILLER_48_220 ();
 sg13g2_decap_8 FILLER_48_225 ();
 sg13g2_decap_8 FILLER_48_232 ();
 sg13g2_decap_8 FILLER_48_239 ();
 sg13g2_decap_8 FILLER_48_246 ();
 sg13g2_decap_8 FILLER_48_253 ();
 sg13g2_decap_4 FILLER_48_286 ();
 sg13g2_decap_4 FILLER_48_298 ();
 sg13g2_fill_2 FILLER_48_302 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_fill_2 FILLER_48_361 ();
 sg13g2_fill_1 FILLER_48_367 ();
 sg13g2_fill_1 FILLER_48_377 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_fill_2 FILLER_49_112 ();
 sg13g2_fill_1 FILLER_49_145 ();
 sg13g2_fill_2 FILLER_49_172 ();
 sg13g2_fill_2 FILLER_49_213 ();
 sg13g2_fill_1 FILLER_49_215 ();
 sg13g2_fill_2 FILLER_49_220 ();
 sg13g2_fill_1 FILLER_49_222 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_fill_2 FILLER_49_288 ();
 sg13g2_fill_1 FILLER_49_290 ();
 sg13g2_fill_1 FILLER_49_327 ();
 sg13g2_fill_1 FILLER_49_342 ();
 sg13g2_fill_2 FILLER_49_347 ();
 sg13g2_fill_1 FILLER_49_349 ();
 sg13g2_decap_8 FILLER_49_376 ();
 sg13g2_fill_2 FILLER_49_383 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_fill_1 FILLER_50_130 ();
 sg13g2_fill_1 FILLER_50_166 ();
 sg13g2_fill_2 FILLER_50_171 ();
 sg13g2_decap_4 FILLER_50_179 ();
 sg13g2_decap_4 FILLER_50_187 ();
 sg13g2_fill_1 FILLER_50_195 ();
 sg13g2_fill_2 FILLER_50_210 ();
 sg13g2_decap_8 FILLER_50_248 ();
 sg13g2_fill_1 FILLER_50_255 ();
 sg13g2_fill_1 FILLER_50_261 ();
 sg13g2_fill_1 FILLER_50_265 ();
 sg13g2_fill_1 FILLER_50_275 ();
 sg13g2_decap_4 FILLER_50_307 ();
 sg13g2_fill_1 FILLER_50_388 ();
 sg13g2_fill_2 FILLER_50_394 ();
 sg13g2_decap_4 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_50_411 ();
 sg13g2_decap_8 FILLER_50_418 ();
 sg13g2_decap_4 FILLER_50_425 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_fill_1 FILLER_51_119 ();
 sg13g2_decap_4 FILLER_51_125 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_148 ();
 sg13g2_decap_8 FILLER_51_155 ();
 sg13g2_fill_1 FILLER_51_167 ();
 sg13g2_fill_1 FILLER_51_176 ();
 sg13g2_fill_1 FILLER_51_193 ();
 sg13g2_decap_8 FILLER_51_208 ();
 sg13g2_decap_8 FILLER_51_215 ();
 sg13g2_decap_4 FILLER_51_226 ();
 sg13g2_decap_4 FILLER_51_234 ();
 sg13g2_decap_8 FILLER_51_242 ();
 sg13g2_decap_8 FILLER_51_249 ();
 sg13g2_decap_8 FILLER_51_256 ();
 sg13g2_fill_1 FILLER_51_263 ();
 sg13g2_fill_2 FILLER_51_268 ();
 sg13g2_fill_1 FILLER_51_270 ();
 sg13g2_decap_8 FILLER_51_275 ();
 sg13g2_fill_2 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_284 ();
 sg13g2_fill_2 FILLER_51_294 ();
 sg13g2_fill_1 FILLER_51_296 ();
 sg13g2_fill_1 FILLER_51_302 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_decap_8 FILLER_51_314 ();
 sg13g2_decap_8 FILLER_51_321 ();
 sg13g2_fill_1 FILLER_51_328 ();
 sg13g2_decap_8 FILLER_51_333 ();
 sg13g2_fill_1 FILLER_51_345 ();
 sg13g2_fill_2 FILLER_51_351 ();
 sg13g2_fill_2 FILLER_51_357 ();
 sg13g2_fill_2 FILLER_51_363 ();
 sg13g2_fill_1 FILLER_51_395 ();
 sg13g2_fill_2 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_403 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_fill_1 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_130 ();
 sg13g2_decap_8 FILLER_52_137 ();
 sg13g2_decap_8 FILLER_52_144 ();
 sg13g2_decap_8 FILLER_52_151 ();
 sg13g2_fill_2 FILLER_52_158 ();
 sg13g2_fill_2 FILLER_52_171 ();
 sg13g2_fill_1 FILLER_52_177 ();
 sg13g2_fill_1 FILLER_52_182 ();
 sg13g2_fill_2 FILLER_52_186 ();
 sg13g2_decap_8 FILLER_52_196 ();
 sg13g2_fill_1 FILLER_52_203 ();
 sg13g2_fill_1 FILLER_52_211 ();
 sg13g2_fill_1 FILLER_52_217 ();
 sg13g2_fill_2 FILLER_52_223 ();
 sg13g2_fill_1 FILLER_52_255 ();
 sg13g2_decap_8 FILLER_52_272 ();
 sg13g2_fill_2 FILLER_52_283 ();
 sg13g2_fill_2 FILLER_52_293 ();
 sg13g2_fill_1 FILLER_52_295 ();
 sg13g2_decap_4 FILLER_52_327 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_fill_2 FILLER_52_364 ();
 sg13g2_fill_1 FILLER_52_366 ();
 sg13g2_fill_2 FILLER_52_397 ();
 sg13g2_fill_1 FILLER_52_399 ();
 sg13g2_decap_4 FILLER_52_414 ();
 sg13g2_fill_1 FILLER_52_418 ();
 sg13g2_decap_8 FILLER_52_423 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_4 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_fill_2 FILLER_53_143 ();
 sg13g2_fill_1 FILLER_53_145 ();
 sg13g2_decap_4 FILLER_53_151 ();
 sg13g2_fill_2 FILLER_53_155 ();
 sg13g2_decap_8 FILLER_53_164 ();
 sg13g2_fill_2 FILLER_53_171 ();
 sg13g2_decap_4 FILLER_53_182 ();
 sg13g2_fill_2 FILLER_53_191 ();
 sg13g2_fill_1 FILLER_53_198 ();
 sg13g2_fill_2 FILLER_53_203 ();
 sg13g2_fill_1 FILLER_53_216 ();
 sg13g2_decap_4 FILLER_53_225 ();
 sg13g2_fill_1 FILLER_53_229 ();
 sg13g2_decap_4 FILLER_53_238 ();
 sg13g2_fill_2 FILLER_53_242 ();
 sg13g2_fill_2 FILLER_53_252 ();
 sg13g2_fill_1 FILLER_53_254 ();
 sg13g2_decap_8 FILLER_53_311 ();
 sg13g2_decap_8 FILLER_53_318 ();
 sg13g2_decap_8 FILLER_53_325 ();
 sg13g2_decap_4 FILLER_53_332 ();
 sg13g2_fill_1 FILLER_53_336 ();
 sg13g2_decap_8 FILLER_53_360 ();
 sg13g2_decap_8 FILLER_53_367 ();
 sg13g2_fill_2 FILLER_53_374 ();
 sg13g2_fill_2 FILLER_53_381 ();
 sg13g2_fill_2 FILLER_53_395 ();
 sg13g2_decap_8 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_53_414 ();
 sg13g2_decap_8 FILLER_53_421 ();
 sg13g2_fill_2 FILLER_53_428 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_fill_2 FILLER_54_112 ();
 sg13g2_fill_1 FILLER_54_114 ();
 sg13g2_decap_8 FILLER_54_155 ();
 sg13g2_fill_1 FILLER_54_162 ();
 sg13g2_fill_1 FILLER_54_171 ();
 sg13g2_fill_2 FILLER_54_177 ();
 sg13g2_fill_1 FILLER_54_186 ();
 sg13g2_decap_8 FILLER_54_226 ();
 sg13g2_decap_8 FILLER_54_246 ();
 sg13g2_decap_4 FILLER_54_253 ();
 sg13g2_fill_2 FILLER_54_283 ();
 sg13g2_fill_1 FILLER_54_285 ();
 sg13g2_decap_4 FILLER_54_296 ();
 sg13g2_fill_1 FILLER_54_300 ();
 sg13g2_decap_4 FILLER_54_310 ();
 sg13g2_fill_2 FILLER_54_314 ();
 sg13g2_decap_8 FILLER_54_321 ();
 sg13g2_fill_2 FILLER_54_328 ();
 sg13g2_decap_4 FILLER_54_334 ();
 sg13g2_fill_2 FILLER_54_338 ();
 sg13g2_fill_2 FILLER_54_344 ();
 sg13g2_decap_4 FILLER_54_350 ();
 sg13g2_fill_2 FILLER_54_354 ();
 sg13g2_decap_8 FILLER_54_360 ();
 sg13g2_decap_8 FILLER_54_367 ();
 sg13g2_decap_8 FILLER_54_374 ();
 sg13g2_decap_8 FILLER_54_381 ();
 sg13g2_decap_8 FILLER_54_388 ();
 sg13g2_decap_4 FILLER_54_395 ();
 sg13g2_fill_1 FILLER_54_399 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_4 FILLER_55_112 ();
 sg13g2_fill_2 FILLER_55_126 ();
 sg13g2_fill_1 FILLER_55_128 ();
 sg13g2_fill_1 FILLER_55_146 ();
 sg13g2_decap_4 FILLER_55_157 ();
 sg13g2_fill_2 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_176 ();
 sg13g2_fill_2 FILLER_55_183 ();
 sg13g2_fill_2 FILLER_55_227 ();
 sg13g2_fill_1 FILLER_55_229 ();
 sg13g2_decap_4 FILLER_55_256 ();
 sg13g2_fill_2 FILLER_55_260 ();
 sg13g2_decap_4 FILLER_55_290 ();
 sg13g2_fill_1 FILLER_55_294 ();
 sg13g2_fill_2 FILLER_55_299 ();
 sg13g2_fill_1 FILLER_55_301 ();
 sg13g2_fill_2 FILLER_55_332 ();
 sg13g2_fill_1 FILLER_55_334 ();
 sg13g2_fill_2 FILLER_55_379 ();
 sg13g2_fill_2 FILLER_55_385 ();
 sg13g2_fill_1 FILLER_55_387 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_fill_1 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_406 ();
 sg13g2_fill_2 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_419 ();
 sg13g2_decap_4 FILLER_55_426 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_4 FILLER_56_105 ();
 sg13g2_fill_2 FILLER_56_109 ();
 sg13g2_decap_4 FILLER_56_124 ();
 sg13g2_fill_1 FILLER_56_128 ();
 sg13g2_fill_1 FILLER_56_134 ();
 sg13g2_decap_4 FILLER_56_143 ();
 sg13g2_decap_8 FILLER_56_151 ();
 sg13g2_decap_8 FILLER_56_158 ();
 sg13g2_fill_2 FILLER_56_170 ();
 sg13g2_fill_1 FILLER_56_172 ();
 sg13g2_decap_4 FILLER_56_184 ();
 sg13g2_fill_1 FILLER_56_188 ();
 sg13g2_fill_2 FILLER_56_199 ();
 sg13g2_fill_1 FILLER_56_201 ();
 sg13g2_decap_4 FILLER_56_232 ();
 sg13g2_fill_2 FILLER_56_236 ();
 sg13g2_fill_2 FILLER_56_242 ();
 sg13g2_fill_1 FILLER_56_248 ();
 sg13g2_decap_8 FILLER_56_253 ();
 sg13g2_decap_8 FILLER_56_260 ();
 sg13g2_decap_4 FILLER_56_267 ();
 sg13g2_fill_1 FILLER_56_271 ();
 sg13g2_fill_1 FILLER_56_281 ();
 sg13g2_fill_2 FILLER_56_288 ();
 sg13g2_fill_2 FILLER_56_295 ();
 sg13g2_decap_4 FILLER_56_305 ();
 sg13g2_fill_1 FILLER_56_309 ();
 sg13g2_fill_2 FILLER_56_319 ();
 sg13g2_fill_1 FILLER_56_321 ();
 sg13g2_fill_2 FILLER_56_326 ();
 sg13g2_fill_1 FILLER_56_343 ();
 sg13g2_fill_1 FILLER_56_348 ();
 sg13g2_fill_2 FILLER_56_353 ();
 sg13g2_fill_2 FILLER_56_360 ();
 sg13g2_fill_2 FILLER_56_400 ();
 sg13g2_decap_8 FILLER_56_406 ();
 sg13g2_decap_8 FILLER_56_413 ();
 sg13g2_decap_8 FILLER_56_420 ();
 sg13g2_fill_2 FILLER_56_427 ();
 sg13g2_fill_1 FILLER_56_429 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_124 ();
 sg13g2_decap_8 FILLER_57_131 ();
 sg13g2_fill_2 FILLER_57_138 ();
 sg13g2_fill_1 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_159 ();
 sg13g2_decap_4 FILLER_57_166 ();
 sg13g2_fill_2 FILLER_57_170 ();
 sg13g2_fill_2 FILLER_57_192 ();
 sg13g2_fill_1 FILLER_57_194 ();
 sg13g2_decap_8 FILLER_57_204 ();
 sg13g2_fill_1 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_229 ();
 sg13g2_decap_8 FILLER_57_236 ();
 sg13g2_fill_2 FILLER_57_277 ();
 sg13g2_fill_2 FILLER_57_291 ();
 sg13g2_fill_1 FILLER_57_328 ();
 sg13g2_fill_1 FILLER_57_334 ();
 sg13g2_fill_1 FILLER_57_339 ();
 sg13g2_fill_2 FILLER_57_343 ();
 sg13g2_decap_4 FILLER_57_351 ();
 sg13g2_decap_4 FILLER_57_368 ();
 sg13g2_fill_1 FILLER_57_372 ();
 sg13g2_decap_8 FILLER_57_377 ();
 sg13g2_fill_1 FILLER_57_388 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_4 FILLER_58_112 ();
 sg13g2_fill_1 FILLER_58_116 ();
 sg13g2_decap_8 FILLER_58_121 ();
 sg13g2_decap_8 FILLER_58_128 ();
 sg13g2_decap_8 FILLER_58_135 ();
 sg13g2_decap_8 FILLER_58_142 ();
 sg13g2_decap_8 FILLER_58_149 ();
 sg13g2_decap_8 FILLER_58_156 ();
 sg13g2_decap_8 FILLER_58_163 ();
 sg13g2_decap_8 FILLER_58_170 ();
 sg13g2_decap_4 FILLER_58_177 ();
 sg13g2_decap_4 FILLER_58_186 ();
 sg13g2_fill_2 FILLER_58_194 ();
 sg13g2_fill_1 FILLER_58_196 ();
 sg13g2_decap_4 FILLER_58_202 ();
 sg13g2_fill_2 FILLER_58_206 ();
 sg13g2_decap_8 FILLER_58_212 ();
 sg13g2_decap_4 FILLER_58_219 ();
 sg13g2_fill_1 FILLER_58_223 ();
 sg13g2_decap_8 FILLER_58_233 ();
 sg13g2_fill_2 FILLER_58_240 ();
 sg13g2_decap_8 FILLER_58_252 ();
 sg13g2_decap_4 FILLER_58_263 ();
 sg13g2_decap_4 FILLER_58_276 ();
 sg13g2_fill_1 FILLER_58_280 ();
 sg13g2_fill_2 FILLER_58_315 ();
 sg13g2_fill_1 FILLER_58_317 ();
 sg13g2_decap_4 FILLER_58_323 ();
 sg13g2_fill_2 FILLER_58_359 ();
 sg13g2_decap_4 FILLER_58_366 ();
 sg13g2_fill_2 FILLER_58_378 ();
 sg13g2_decap_8 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_392 ();
 sg13g2_decap_4 FILLER_58_399 ();
 sg13g2_fill_1 FILLER_58_413 ();
 sg13g2_decap_8 FILLER_58_418 ();
 sg13g2_decap_4 FILLER_58_425 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_4 FILLER_59_105 ();
 sg13g2_fill_1 FILLER_59_109 ();
 sg13g2_fill_2 FILLER_59_124 ();
 sg13g2_fill_1 FILLER_59_126 ();
 sg13g2_decap_4 FILLER_59_151 ();
 sg13g2_fill_1 FILLER_59_155 ();
 sg13g2_decap_8 FILLER_59_160 ();
 sg13g2_decap_4 FILLER_59_171 ();
 sg13g2_fill_1 FILLER_59_175 ();
 sg13g2_fill_2 FILLER_59_194 ();
 sg13g2_fill_1 FILLER_59_214 ();
 sg13g2_decap_4 FILLER_59_226 ();
 sg13g2_fill_2 FILLER_59_230 ();
 sg13g2_fill_2 FILLER_59_236 ();
 sg13g2_fill_1 FILLER_59_238 ();
 sg13g2_fill_2 FILLER_59_248 ();
 sg13g2_decap_8 FILLER_59_276 ();
 sg13g2_fill_2 FILLER_59_283 ();
 sg13g2_fill_1 FILLER_59_285 ();
 sg13g2_fill_2 FILLER_59_291 ();
 sg13g2_fill_1 FILLER_59_293 ();
 sg13g2_decap_8 FILLER_59_307 ();
 sg13g2_decap_4 FILLER_59_314 ();
 sg13g2_fill_2 FILLER_59_318 ();
 sg13g2_fill_2 FILLER_59_329 ();
 sg13g2_fill_1 FILLER_59_345 ();
 sg13g2_fill_2 FILLER_59_350 ();
 sg13g2_fill_1 FILLER_59_391 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_decap_8 FILLER_59_420 ();
 sg13g2_fill_2 FILLER_59_427 ();
 sg13g2_fill_1 FILLER_59_429 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_4 FILLER_60_98 ();
 sg13g2_fill_2 FILLER_60_102 ();
 sg13g2_fill_2 FILLER_60_123 ();
 sg13g2_fill_1 FILLER_60_140 ();
 sg13g2_fill_2 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_223 ();
 sg13g2_fill_1 FILLER_60_235 ();
 sg13g2_fill_2 FILLER_60_241 ();
 sg13g2_fill_1 FILLER_60_258 ();
 sg13g2_decap_8 FILLER_60_271 ();
 sg13g2_decap_8 FILLER_60_278 ();
 sg13g2_decap_8 FILLER_60_285 ();
 sg13g2_fill_2 FILLER_60_292 ();
 sg13g2_fill_2 FILLER_60_303 ();
 sg13g2_decap_8 FILLER_60_315 ();
 sg13g2_fill_2 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_60_324 ();
 sg13g2_fill_2 FILLER_60_330 ();
 sg13g2_fill_1 FILLER_60_332 ();
 sg13g2_decap_4 FILLER_60_338 ();
 sg13g2_decap_8 FILLER_60_346 ();
 sg13g2_decap_4 FILLER_60_353 ();
 sg13g2_decap_8 FILLER_60_361 ();
 sg13g2_fill_1 FILLER_60_368 ();
 sg13g2_decap_8 FILLER_60_374 ();
 sg13g2_fill_1 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_60_386 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_60_422 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_fill_1 FILLER_61_98 ();
 sg13g2_fill_1 FILLER_61_103 ();
 sg13g2_fill_1 FILLER_61_109 ();
 sg13g2_fill_2 FILLER_61_123 ();
 sg13g2_fill_1 FILLER_61_125 ();
 sg13g2_fill_1 FILLER_61_146 ();
 sg13g2_fill_1 FILLER_61_152 ();
 sg13g2_fill_1 FILLER_61_158 ();
 sg13g2_fill_2 FILLER_61_185 ();
 sg13g2_decap_8 FILLER_61_192 ();
 sg13g2_decap_4 FILLER_61_199 ();
 sg13g2_fill_1 FILLER_61_203 ();
 sg13g2_decap_4 FILLER_61_213 ();
 sg13g2_fill_2 FILLER_61_267 ();
 sg13g2_fill_1 FILLER_61_269 ();
 sg13g2_decap_8 FILLER_61_274 ();
 sg13g2_decap_8 FILLER_61_281 ();
 sg13g2_decap_4 FILLER_61_288 ();
 sg13g2_fill_1 FILLER_61_292 ();
 sg13g2_fill_2 FILLER_61_297 ();
 sg13g2_fill_1 FILLER_61_299 ();
 sg13g2_decap_4 FILLER_61_306 ();
 sg13g2_fill_1 FILLER_61_310 ();
 sg13g2_fill_1 FILLER_61_330 ();
 sg13g2_fill_2 FILLER_61_337 ();
 sg13g2_fill_1 FILLER_61_339 ();
 sg13g2_fill_1 FILLER_61_344 ();
 sg13g2_decap_8 FILLER_61_349 ();
 sg13g2_decap_8 FILLER_61_356 ();
 sg13g2_decap_8 FILLER_61_363 ();
 sg13g2_decap_8 FILLER_61_370 ();
 sg13g2_decap_8 FILLER_61_377 ();
 sg13g2_fill_2 FILLER_61_384 ();
 sg13g2_fill_1 FILLER_61_386 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_decap_4 FILLER_61_398 ();
 sg13g2_fill_2 FILLER_61_402 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_fill_2 FILLER_62_98 ();
 sg13g2_fill_1 FILLER_62_100 ();
 sg13g2_fill_1 FILLER_62_105 ();
 sg13g2_fill_1 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_125 ();
 sg13g2_fill_1 FILLER_62_132 ();
 sg13g2_fill_1 FILLER_62_138 ();
 sg13g2_fill_1 FILLER_62_144 ();
 sg13g2_fill_2 FILLER_62_154 ();
 sg13g2_fill_2 FILLER_62_160 ();
 sg13g2_fill_1 FILLER_62_193 ();
 sg13g2_decap_8 FILLER_62_199 ();
 sg13g2_decap_8 FILLER_62_206 ();
 sg13g2_decap_8 FILLER_62_213 ();
 sg13g2_decap_4 FILLER_62_220 ();
 sg13g2_decap_8 FILLER_62_228 ();
 sg13g2_fill_2 FILLER_62_235 ();
 sg13g2_fill_1 FILLER_62_237 ();
 sg13g2_fill_2 FILLER_62_248 ();
 sg13g2_decap_4 FILLER_62_276 ();
 sg13g2_fill_2 FILLER_62_280 ();
 sg13g2_decap_4 FILLER_62_312 ();
 sg13g2_decap_4 FILLER_62_321 ();
 sg13g2_fill_2 FILLER_62_330 ();
 sg13g2_fill_1 FILLER_62_332 ();
 sg13g2_decap_4 FILLER_62_368 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_decap_4 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_415 ();
 sg13g2_fill_1 FILLER_62_426 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_4 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_109 ();
 sg13g2_decap_4 FILLER_63_115 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_fill_2 FILLER_63_140 ();
 sg13g2_fill_1 FILLER_63_142 ();
 sg13g2_fill_2 FILLER_63_153 ();
 sg13g2_decap_4 FILLER_63_159 ();
 sg13g2_fill_1 FILLER_63_163 ();
 sg13g2_decap_8 FILLER_63_173 ();
 sg13g2_decap_8 FILLER_63_180 ();
 sg13g2_decap_8 FILLER_63_187 ();
 sg13g2_decap_8 FILLER_63_194 ();
 sg13g2_decap_8 FILLER_63_204 ();
 sg13g2_fill_2 FILLER_63_211 ();
 sg13g2_decap_4 FILLER_63_217 ();
 sg13g2_fill_2 FILLER_63_221 ();
 sg13g2_fill_2 FILLER_63_227 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_fill_2 FILLER_63_252 ();
 sg13g2_fill_1 FILLER_63_254 ();
 sg13g2_decap_8 FILLER_63_264 ();
 sg13g2_decap_8 FILLER_63_271 ();
 sg13g2_decap_4 FILLER_63_278 ();
 sg13g2_fill_2 FILLER_63_287 ();
 sg13g2_fill_1 FILLER_63_289 ();
 sg13g2_decap_8 FILLER_63_298 ();
 sg13g2_decap_8 FILLER_63_305 ();
 sg13g2_decap_4 FILLER_63_312 ();
 sg13g2_fill_2 FILLER_63_316 ();
 sg13g2_decap_8 FILLER_63_324 ();
 sg13g2_decap_4 FILLER_63_342 ();
 sg13g2_decap_8 FILLER_63_355 ();
 sg13g2_fill_1 FILLER_63_362 ();
 sg13g2_fill_2 FILLER_63_401 ();
 sg13g2_fill_1 FILLER_63_417 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_fill_2 FILLER_64_105 ();
 sg13g2_fill_1 FILLER_64_126 ();
 sg13g2_fill_1 FILLER_64_135 ();
 sg13g2_decap_4 FILLER_64_154 ();
 sg13g2_fill_1 FILLER_64_158 ();
 sg13g2_fill_2 FILLER_64_193 ();
 sg13g2_fill_1 FILLER_64_195 ();
 sg13g2_decap_8 FILLER_64_206 ();
 sg13g2_decap_4 FILLER_64_213 ();
 sg13g2_fill_1 FILLER_64_221 ();
 sg13g2_fill_1 FILLER_64_254 ();
 sg13g2_fill_2 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_308 ();
 sg13g2_decap_8 FILLER_64_315 ();
 sg13g2_fill_1 FILLER_64_326 ();
 sg13g2_fill_1 FILLER_64_331 ();
 sg13g2_fill_2 FILLER_64_381 ();
 sg13g2_decap_8 FILLER_64_398 ();
 sg13g2_decap_8 FILLER_64_405 ();
 sg13g2_decap_8 FILLER_64_412 ();
 sg13g2_decap_8 FILLER_64_419 ();
 sg13g2_decap_4 FILLER_64_426 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_4 FILLER_65_105 ();
 sg13g2_fill_1 FILLER_65_114 ();
 sg13g2_decap_4 FILLER_65_128 ();
 sg13g2_fill_2 FILLER_65_132 ();
 sg13g2_fill_2 FILLER_65_158 ();
 sg13g2_fill_2 FILLER_65_225 ();
 sg13g2_fill_1 FILLER_65_232 ();
 sg13g2_decap_8 FILLER_65_268 ();
 sg13g2_decap_4 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_279 ();
 sg13g2_decap_4 FILLER_65_285 ();
 sg13g2_fill_2 FILLER_65_289 ();
 sg13g2_fill_1 FILLER_65_310 ();
 sg13g2_decap_4 FILLER_65_319 ();
 sg13g2_fill_1 FILLER_65_323 ();
 sg13g2_fill_1 FILLER_65_329 ();
 sg13g2_fill_1 FILLER_65_346 ();
 sg13g2_fill_2 FILLER_65_352 ();
 sg13g2_fill_1 FILLER_65_354 ();
 sg13g2_fill_1 FILLER_65_362 ();
 sg13g2_fill_1 FILLER_65_371 ();
 sg13g2_fill_2 FILLER_65_382 ();
 sg13g2_decap_4 FILLER_65_425 ();
 sg13g2_fill_1 FILLER_65_429 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_fill_1 FILLER_66_105 ();
 sg13g2_fill_2 FILLER_66_111 ();
 sg13g2_fill_1 FILLER_66_122 ();
 sg13g2_fill_1 FILLER_66_128 ();
 sg13g2_fill_1 FILLER_66_133 ();
 sg13g2_fill_2 FILLER_66_151 ();
 sg13g2_decap_8 FILLER_66_158 ();
 sg13g2_fill_2 FILLER_66_165 ();
 sg13g2_fill_1 FILLER_66_167 ();
 sg13g2_decap_8 FILLER_66_172 ();
 sg13g2_decap_8 FILLER_66_179 ();
 sg13g2_fill_1 FILLER_66_186 ();
 sg13g2_decap_8 FILLER_66_192 ();
 sg13g2_fill_1 FILLER_66_199 ();
 sg13g2_fill_2 FILLER_66_204 ();
 sg13g2_fill_1 FILLER_66_220 ();
 sg13g2_fill_1 FILLER_66_225 ();
 sg13g2_decap_8 FILLER_66_257 ();
 sg13g2_decap_4 FILLER_66_264 ();
 sg13g2_fill_1 FILLER_66_268 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_4 FILLER_66_280 ();
 sg13g2_fill_2 FILLER_66_284 ();
 sg13g2_fill_2 FILLER_66_291 ();
 sg13g2_fill_1 FILLER_66_331 ();
 sg13g2_fill_2 FILLER_66_342 ();
 sg13g2_decap_8 FILLER_66_359 ();
 sg13g2_decap_8 FILLER_66_366 ();
 sg13g2_fill_1 FILLER_66_386 ();
 sg13g2_fill_2 FILLER_66_392 ();
 sg13g2_fill_1 FILLER_66_394 ();
 sg13g2_decap_4 FILLER_66_400 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_fill_1 FILLER_67_116 ();
 sg13g2_fill_1 FILLER_67_125 ();
 sg13g2_fill_1 FILLER_67_140 ();
 sg13g2_fill_2 FILLER_67_151 ();
 sg13g2_fill_1 FILLER_67_153 ();
 sg13g2_decap_8 FILLER_67_159 ();
 sg13g2_fill_2 FILLER_67_166 ();
 sg13g2_decap_8 FILLER_67_172 ();
 sg13g2_fill_1 FILLER_67_179 ();
 sg13g2_decap_4 FILLER_67_215 ();
 sg13g2_fill_2 FILLER_67_236 ();
 sg13g2_fill_1 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_247 ();
 sg13g2_decap_4 FILLER_67_254 ();
 sg13g2_fill_2 FILLER_67_258 ();
 sg13g2_decap_4 FILLER_67_320 ();
 sg13g2_fill_2 FILLER_67_324 ();
 sg13g2_decap_8 FILLER_67_335 ();
 sg13g2_decap_4 FILLER_67_342 ();
 sg13g2_fill_2 FILLER_67_346 ();
 sg13g2_fill_2 FILLER_67_351 ();
 sg13g2_fill_1 FILLER_67_353 ();
 sg13g2_decap_4 FILLER_67_359 ();
 sg13g2_fill_1 FILLER_67_363 ();
 sg13g2_fill_2 FILLER_67_377 ();
 sg13g2_fill_1 FILLER_67_379 ();
 sg13g2_fill_1 FILLER_67_390 ();
 sg13g2_decap_4 FILLER_67_396 ();
 sg13g2_decap_8 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_67_415 ();
 sg13g2_decap_8 FILLER_67_422 ();
 sg13g2_fill_1 FILLER_67_429 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_fill_2 FILLER_68_105 ();
 sg13g2_fill_1 FILLER_68_115 ();
 sg13g2_fill_2 FILLER_68_125 ();
 sg13g2_fill_1 FILLER_68_131 ();
 sg13g2_fill_2 FILLER_68_136 ();
 sg13g2_decap_8 FILLER_68_155 ();
 sg13g2_decap_8 FILLER_68_162 ();
 sg13g2_decap_8 FILLER_68_169 ();
 sg13g2_decap_8 FILLER_68_176 ();
 sg13g2_fill_2 FILLER_68_183 ();
 sg13g2_fill_1 FILLER_68_185 ();
 sg13g2_decap_4 FILLER_68_194 ();
 sg13g2_decap_8 FILLER_68_202 ();
 sg13g2_decap_4 FILLER_68_223 ();
 sg13g2_decap_8 FILLER_68_233 ();
 sg13g2_decap_4 FILLER_68_240 ();
 sg13g2_fill_2 FILLER_68_244 ();
 sg13g2_fill_2 FILLER_68_285 ();
 sg13g2_fill_1 FILLER_68_287 ();
 sg13g2_fill_2 FILLER_68_306 ();
 sg13g2_decap_8 FILLER_68_318 ();
 sg13g2_fill_2 FILLER_68_325 ();
 sg13g2_fill_1 FILLER_68_327 ();
 sg13g2_decap_8 FILLER_68_332 ();
 sg13g2_fill_1 FILLER_68_339 ();
 sg13g2_fill_2 FILLER_68_352 ();
 sg13g2_fill_1 FILLER_68_366 ();
 sg13g2_fill_1 FILLER_68_388 ();
 sg13g2_decap_8 FILLER_68_409 ();
 sg13g2_decap_8 FILLER_68_416 ();
 sg13g2_decap_8 FILLER_68_423 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_fill_2 FILLER_69_119 ();
 sg13g2_decap_4 FILLER_69_139 ();
 sg13g2_decap_4 FILLER_69_148 ();
 sg13g2_fill_2 FILLER_69_152 ();
 sg13g2_decap_8 FILLER_69_184 ();
 sg13g2_decap_8 FILLER_69_195 ();
 sg13g2_decap_4 FILLER_69_202 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_decap_4 FILLER_69_216 ();
 sg13g2_decap_8 FILLER_69_225 ();
 sg13g2_decap_4 FILLER_69_232 ();
 sg13g2_fill_1 FILLER_69_236 ();
 sg13g2_fill_1 FILLER_69_242 ();
 sg13g2_decap_8 FILLER_69_248 ();
 sg13g2_decap_8 FILLER_69_255 ();
 sg13g2_decap_8 FILLER_69_262 ();
 sg13g2_decap_8 FILLER_69_269 ();
 sg13g2_decap_8 FILLER_69_276 ();
 sg13g2_decap_8 FILLER_69_283 ();
 sg13g2_decap_4 FILLER_69_298 ();
 sg13g2_fill_1 FILLER_69_302 ();
 sg13g2_fill_1 FILLER_69_313 ();
 sg13g2_fill_1 FILLER_69_356 ();
 sg13g2_fill_1 FILLER_69_362 ();
 sg13g2_fill_2 FILLER_69_368 ();
 sg13g2_fill_1 FILLER_69_376 ();
 sg13g2_fill_2 FILLER_69_382 ();
 sg13g2_fill_2 FILLER_69_399 ();
 sg13g2_decap_8 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_69_412 ();
 sg13g2_decap_8 FILLER_69_419 ();
 sg13g2_decap_4 FILLER_69_426 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_4 FILLER_70_105 ();
 sg13g2_fill_2 FILLER_70_122 ();
 sg13g2_fill_1 FILLER_70_128 ();
 sg13g2_fill_1 FILLER_70_144 ();
 sg13g2_decap_4 FILLER_70_150 ();
 sg13g2_fill_1 FILLER_70_154 ();
 sg13g2_decap_4 FILLER_70_185 ();
 sg13g2_fill_2 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_195 ();
 sg13g2_fill_2 FILLER_70_212 ();
 sg13g2_decap_8 FILLER_70_225 ();
 sg13g2_fill_1 FILLER_70_232 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_decap_8 FILLER_70_252 ();
 sg13g2_decap_4 FILLER_70_259 ();
 sg13g2_fill_2 FILLER_70_263 ();
 sg13g2_decap_8 FILLER_70_268 ();
 sg13g2_decap_8 FILLER_70_279 ();
 sg13g2_fill_1 FILLER_70_286 ();
 sg13g2_decap_8 FILLER_70_297 ();
 sg13g2_decap_8 FILLER_70_304 ();
 sg13g2_decap_4 FILLER_70_311 ();
 sg13g2_fill_2 FILLER_70_315 ();
 sg13g2_decap_4 FILLER_70_330 ();
 sg13g2_fill_1 FILLER_70_346 ();
 sg13g2_fill_2 FILLER_70_350 ();
 sg13g2_fill_1 FILLER_70_399 ();
 sg13g2_fill_1 FILLER_70_406 ();
 sg13g2_decap_8 FILLER_70_411 ();
 sg13g2_decap_8 FILLER_70_418 ();
 sg13g2_decap_4 FILLER_70_425 ();
 sg13g2_fill_1 FILLER_70_429 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_4 FILLER_71_105 ();
 sg13g2_decap_4 FILLER_71_153 ();
 sg13g2_fill_1 FILLER_71_157 ();
 sg13g2_decap_8 FILLER_71_184 ();
 sg13g2_decap_8 FILLER_71_191 ();
 sg13g2_fill_1 FILLER_71_198 ();
 sg13g2_decap_4 FILLER_71_263 ();
 sg13g2_fill_2 FILLER_71_267 ();
 sg13g2_decap_8 FILLER_71_304 ();
 sg13g2_decap_4 FILLER_71_311 ();
 sg13g2_decap_8 FILLER_71_325 ();
 sg13g2_decap_8 FILLER_71_332 ();
 sg13g2_fill_2 FILLER_71_339 ();
 sg13g2_decap_8 FILLER_71_357 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_decap_4 FILLER_71_378 ();
 sg13g2_fill_1 FILLER_71_392 ();
 sg13g2_fill_1 FILLER_71_401 ();
 sg13g2_decap_8 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_71_414 ();
 sg13g2_decap_8 FILLER_71_421 ();
 sg13g2_fill_2 FILLER_71_428 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_4 FILLER_72_112 ();
 sg13g2_fill_2 FILLER_72_125 ();
 sg13g2_fill_1 FILLER_72_132 ();
 sg13g2_fill_1 FILLER_72_146 ();
 sg13g2_decap_8 FILLER_72_152 ();
 sg13g2_decap_4 FILLER_72_159 ();
 sg13g2_fill_1 FILLER_72_163 ();
 sg13g2_decap_4 FILLER_72_172 ();
 sg13g2_fill_2 FILLER_72_176 ();
 sg13g2_fill_1 FILLER_72_209 ();
 sg13g2_fill_1 FILLER_72_249 ();
 sg13g2_fill_1 FILLER_72_255 ();
 sg13g2_fill_1 FILLER_72_287 ();
 sg13g2_decap_4 FILLER_72_312 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_decap_4 FILLER_72_328 ();
 sg13g2_decap_4 FILLER_72_338 ();
 sg13g2_fill_1 FILLER_72_342 ();
 sg13g2_fill_2 FILLER_72_347 ();
 sg13g2_fill_1 FILLER_72_349 ();
 sg13g2_fill_2 FILLER_72_368 ();
 sg13g2_fill_1 FILLER_72_370 ();
 sg13g2_decap_8 FILLER_72_376 ();
 sg13g2_decap_4 FILLER_72_383 ();
 sg13g2_fill_2 FILLER_72_387 ();
 sg13g2_decap_8 FILLER_72_394 ();
 sg13g2_decap_8 FILLER_72_401 ();
 sg13g2_decap_8 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_72_415 ();
 sg13g2_decap_8 FILLER_72_422 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_4 FILLER_73_105 ();
 sg13g2_fill_2 FILLER_73_109 ();
 sg13g2_fill_2 FILLER_73_115 ();
 sg13g2_decap_8 FILLER_73_144 ();
 sg13g2_decap_8 FILLER_73_159 ();
 sg13g2_decap_8 FILLER_73_166 ();
 sg13g2_decap_8 FILLER_73_173 ();
 sg13g2_decap_4 FILLER_73_184 ();
 sg13g2_fill_1 FILLER_73_197 ();
 sg13g2_fill_1 FILLER_73_227 ();
 sg13g2_fill_1 FILLER_73_238 ();
 sg13g2_fill_2 FILLER_73_252 ();
 sg13g2_fill_1 FILLER_73_254 ();
 sg13g2_fill_1 FILLER_73_281 ();
 sg13g2_fill_1 FILLER_73_287 ();
 sg13g2_fill_1 FILLER_73_293 ();
 sg13g2_decap_4 FILLER_73_304 ();
 sg13g2_decap_4 FILLER_73_328 ();
 sg13g2_fill_2 FILLER_73_336 ();
 sg13g2_fill_1 FILLER_73_338 ();
 sg13g2_fill_2 FILLER_73_346 ();
 sg13g2_fill_1 FILLER_73_348 ();
 sg13g2_fill_1 FILLER_73_353 ();
 sg13g2_fill_2 FILLER_73_359 ();
 sg13g2_decap_4 FILLER_73_366 ();
 sg13g2_decap_8 FILLER_73_374 ();
 sg13g2_decap_8 FILLER_73_381 ();
 sg13g2_fill_1 FILLER_73_388 ();
 sg13g2_decap_8 FILLER_73_394 ();
 sg13g2_decap_8 FILLER_73_401 ();
 sg13g2_decap_8 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_73_415 ();
 sg13g2_decap_8 FILLER_73_422 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_fill_1 FILLER_74_134 ();
 sg13g2_fill_1 FILLER_74_141 ();
 sg13g2_fill_2 FILLER_74_146 ();
 sg13g2_fill_2 FILLER_74_153 ();
 sg13g2_fill_2 FILLER_74_207 ();
 sg13g2_decap_8 FILLER_74_213 ();
 sg13g2_fill_1 FILLER_74_220 ();
 sg13g2_decap_4 FILLER_74_229 ();
 sg13g2_decap_8 FILLER_74_237 ();
 sg13g2_decap_8 FILLER_74_244 ();
 sg13g2_decap_8 FILLER_74_251 ();
 sg13g2_fill_2 FILLER_74_258 ();
 sg13g2_fill_1 FILLER_74_260 ();
 sg13g2_fill_1 FILLER_74_265 ();
 sg13g2_decap_4 FILLER_74_274 ();
 sg13g2_fill_2 FILLER_74_278 ();
 sg13g2_decap_4 FILLER_74_320 ();
 sg13g2_fill_1 FILLER_74_324 ();
 sg13g2_fill_1 FILLER_74_369 ();
 sg13g2_fill_2 FILLER_74_376 ();
 sg13g2_fill_1 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_decap_8 FILLER_74_406 ();
 sg13g2_decap_8 FILLER_74_413 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_fill_2 FILLER_74_427 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_4 FILLER_75_119 ();
 sg13g2_decap_4 FILLER_75_128 ();
 sg13g2_fill_2 FILLER_75_137 ();
 sg13g2_decap_8 FILLER_75_178 ();
 sg13g2_fill_2 FILLER_75_185 ();
 sg13g2_fill_2 FILLER_75_191 ();
 sg13g2_fill_1 FILLER_75_193 ();
 sg13g2_decap_4 FILLER_75_220 ();
 sg13g2_fill_2 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_fill_2 FILLER_75_287 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_decap_8 FILLER_75_295 ();
 sg13g2_decap_8 FILLER_75_302 ();
 sg13g2_decap_8 FILLER_75_309 ();
 sg13g2_decap_8 FILLER_75_316 ();
 sg13g2_fill_2 FILLER_75_323 ();
 sg13g2_fill_1 FILLER_75_325 ();
 sg13g2_fill_2 FILLER_75_331 ();
 sg13g2_decap_8 FILLER_75_337 ();
 sg13g2_fill_2 FILLER_75_344 ();
 sg13g2_fill_2 FILLER_75_351 ();
 sg13g2_fill_1 FILLER_75_360 ();
 sg13g2_fill_1 FILLER_75_373 ();
 sg13g2_decap_8 FILLER_75_404 ();
 sg13g2_decap_8 FILLER_75_411 ();
 sg13g2_decap_8 FILLER_75_418 ();
 sg13g2_decap_4 FILLER_75_425 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_fill_1 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_159 ();
 sg13g2_decap_8 FILLER_76_166 ();
 sg13g2_decap_8 FILLER_76_173 ();
 sg13g2_decap_8 FILLER_76_180 ();
 sg13g2_decap_8 FILLER_76_187 ();
 sg13g2_decap_4 FILLER_76_194 ();
 sg13g2_fill_2 FILLER_76_198 ();
 sg13g2_decap_4 FILLER_76_204 ();
 sg13g2_fill_1 FILLER_76_208 ();
 sg13g2_decap_8 FILLER_76_218 ();
 sg13g2_decap_8 FILLER_76_225 ();
 sg13g2_fill_2 FILLER_76_232 ();
 sg13g2_fill_1 FILLER_76_234 ();
 sg13g2_decap_8 FILLER_76_291 ();
 sg13g2_decap_8 FILLER_76_298 ();
 sg13g2_decap_4 FILLER_76_305 ();
 sg13g2_fill_2 FILLER_76_312 ();
 sg13g2_fill_1 FILLER_76_340 ();
 sg13g2_decap_4 FILLER_76_361 ();
 sg13g2_fill_1 FILLER_76_377 ();
 sg13g2_decap_8 FILLER_76_394 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_decap_8 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_76_415 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_178 ();
 sg13g2_decap_8 FILLER_77_185 ();
 sg13g2_decap_8 FILLER_77_192 ();
 sg13g2_fill_2 FILLER_77_199 ();
 sg13g2_fill_2 FILLER_77_220 ();
 sg13g2_fill_1 FILLER_77_222 ();
 sg13g2_decap_8 FILLER_77_230 ();
 sg13g2_decap_8 FILLER_77_237 ();
 sg13g2_decap_8 FILLER_77_247 ();
 sg13g2_decap_8 FILLER_77_254 ();
 sg13g2_decap_8 FILLER_77_261 ();
 sg13g2_decap_4 FILLER_77_268 ();
 sg13g2_decap_8 FILLER_77_276 ();
 sg13g2_decap_8 FILLER_77_283 ();
 sg13g2_fill_2 FILLER_77_336 ();
 sg13g2_fill_1 FILLER_77_338 ();
 sg13g2_fill_2 FILLER_77_370 ();
 sg13g2_fill_2 FILLER_77_375 ();
 sg13g2_fill_1 FILLER_77_377 ();
 sg13g2_fill_2 FILLER_77_382 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_fill_2 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_fill_2 FILLER_78_154 ();
 sg13g2_decap_4 FILLER_78_160 ();
 sg13g2_fill_2 FILLER_78_171 ();
 sg13g2_decap_4 FILLER_78_263 ();
 sg13g2_fill_1 FILLER_78_267 ();
 sg13g2_fill_1 FILLER_78_325 ();
 sg13g2_fill_2 FILLER_78_356 ();
 sg13g2_decap_4 FILLER_78_363 ();
 sg13g2_fill_2 FILLER_78_367 ();
 sg13g2_decap_8 FILLER_78_373 ();
 sg13g2_decap_4 FILLER_78_380 ();
 sg13g2_fill_1 FILLER_78_384 ();
 sg13g2_decap_8 FILLER_78_389 ();
 sg13g2_decap_8 FILLER_78_396 ();
 sg13g2_decap_8 FILLER_78_403 ();
 sg13g2_decap_8 FILLER_78_410 ();
 sg13g2_decap_8 FILLER_78_417 ();
 sg13g2_decap_4 FILLER_78_424 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_4 FILLER_79_70 ();
 sg13g2_fill_2 FILLER_79_74 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_116 ();
 sg13g2_decap_8 FILLER_79_123 ();
 sg13g2_decap_8 FILLER_79_130 ();
 sg13g2_decap_8 FILLER_79_137 ();
 sg13g2_decap_8 FILLER_79_144 ();
 sg13g2_decap_8 FILLER_79_151 ();
 sg13g2_decap_8 FILLER_79_158 ();
 sg13g2_decap_8 FILLER_79_165 ();
 sg13g2_fill_1 FILLER_79_172 ();
 sg13g2_decap_4 FILLER_79_181 ();
 sg13g2_decap_4 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_197 ();
 sg13g2_decap_8 FILLER_79_204 ();
 sg13g2_fill_1 FILLER_79_211 ();
 sg13g2_decap_4 FILLER_79_221 ();
 sg13g2_fill_1 FILLER_79_225 ();
 sg13g2_decap_4 FILLER_79_264 ();
 sg13g2_fill_1 FILLER_79_268 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_4 FILLER_79_280 ();
 sg13g2_fill_2 FILLER_79_284 ();
 sg13g2_decap_4 FILLER_79_290 ();
 sg13g2_fill_2 FILLER_79_294 ();
 sg13g2_fill_1 FILLER_79_300 ();
 sg13g2_fill_1 FILLER_79_305 ();
 sg13g2_fill_1 FILLER_79_311 ();
 sg13g2_fill_2 FILLER_79_334 ();
 sg13g2_decap_4 FILLER_79_340 ();
 sg13g2_fill_2 FILLER_79_344 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_4 FILLER_79_357 ();
 sg13g2_fill_1 FILLER_79_361 ();
 sg13g2_decap_8 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_79_409 ();
 sg13g2_decap_8 FILLER_79_416 ();
 sg13g2_decap_8 FILLER_79_423 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_fill_2 FILLER_80_77 ();
 sg13g2_fill_1 FILLER_80_87 ();
 sg13g2_fill_2 FILLER_80_112 ();
 sg13g2_fill_1 FILLER_80_114 ();
 sg13g2_decap_8 FILLER_80_179 ();
 sg13g2_fill_1 FILLER_80_186 ();
 sg13g2_decap_8 FILLER_80_195 ();
 sg13g2_decap_4 FILLER_80_202 ();
 sg13g2_fill_2 FILLER_80_206 ();
 sg13g2_decap_4 FILLER_80_212 ();
 sg13g2_decap_4 FILLER_80_232 ();
 sg13g2_fill_2 FILLER_80_236 ();
 sg13g2_decap_8 FILLER_80_266 ();
 sg13g2_decap_4 FILLER_80_273 ();
 sg13g2_fill_2 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_305 ();
 sg13g2_decap_8 FILLER_80_312 ();
 sg13g2_decap_4 FILLER_80_319 ();
 sg13g2_fill_1 FILLER_80_323 ();
 sg13g2_decap_8 FILLER_80_327 ();
 sg13g2_decap_8 FILLER_80_334 ();
 sg13g2_decap_8 FILLER_80_341 ();
 sg13g2_decap_8 FILLER_80_348 ();
 sg13g2_decap_8 FILLER_80_355 ();
 sg13g2_fill_1 FILLER_80_362 ();
 sg13g2_decap_8 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_374 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_fill_2 FILLER_80_388 ();
 sg13g2_fill_1 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 sg13g2_decap_8 FILLER_80_409 ();
 sg13g2_decap_8 FILLER_80_416 ();
 sg13g2_decap_8 FILLER_80_423 ();
endmodule
