module tt_um_urish_simon (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire clknet_0_clk;
 wire net91;
 wire \simon1.button_released ;
 wire \simon1.lfsr_capture[0] ;
 wire \simon1.lfsr_capture[10] ;
 wire \simon1.lfsr_capture[11] ;
 wire \simon1.lfsr_capture[12] ;
 wire \simon1.lfsr_capture[13] ;
 wire \simon1.lfsr_capture[14] ;
 wire \simon1.lfsr_capture[15] ;
 wire \simon1.lfsr_capture[16] ;
 wire \simon1.lfsr_capture[17] ;
 wire \simon1.lfsr_capture[18] ;
 wire \simon1.lfsr_capture[19] ;
 wire \simon1.lfsr_capture[1] ;
 wire \simon1.lfsr_capture[20] ;
 wire \simon1.lfsr_capture[21] ;
 wire \simon1.lfsr_capture[22] ;
 wire \simon1.lfsr_capture[23] ;
 wire \simon1.lfsr_capture[24] ;
 wire \simon1.lfsr_capture[25] ;
 wire \simon1.lfsr_capture[26] ;
 wire \simon1.lfsr_capture[27] ;
 wire \simon1.lfsr_capture[28] ;
 wire \simon1.lfsr_capture[29] ;
 wire \simon1.lfsr_capture[2] ;
 wire \simon1.lfsr_capture[30] ;
 wire \simon1.lfsr_capture[31] ;
 wire \simon1.lfsr_capture[3] ;
 wire \simon1.lfsr_capture[4] ;
 wire \simon1.lfsr_capture[5] ;
 wire \simon1.lfsr_capture[6] ;
 wire \simon1.lfsr_capture[7] ;
 wire \simon1.lfsr_capture[8] ;
 wire \simon1.lfsr_capture[9] ;
 wire \simon1.lfsr_cycles[0] ;
 wire \simon1.lfsr_cycles[1] ;
 wire \simon1.lfsr_inst.lfsr_out[0] ;
 wire \simon1.lfsr_inst.lfsr_out[10] ;
 wire \simon1.lfsr_inst.lfsr_out[11] ;
 wire \simon1.lfsr_inst.lfsr_out[12] ;
 wire \simon1.lfsr_inst.lfsr_out[13] ;
 wire \simon1.lfsr_inst.lfsr_out[14] ;
 wire \simon1.lfsr_inst.lfsr_out[15] ;
 wire \simon1.lfsr_inst.lfsr_out[16] ;
 wire \simon1.lfsr_inst.lfsr_out[17] ;
 wire \simon1.lfsr_inst.lfsr_out[18] ;
 wire \simon1.lfsr_inst.lfsr_out[19] ;
 wire \simon1.lfsr_inst.lfsr_out[1] ;
 wire \simon1.lfsr_inst.lfsr_out[20] ;
 wire \simon1.lfsr_inst.lfsr_out[21] ;
 wire \simon1.lfsr_inst.lfsr_out[22] ;
 wire \simon1.lfsr_inst.lfsr_out[23] ;
 wire \simon1.lfsr_inst.lfsr_out[24] ;
 wire \simon1.lfsr_inst.lfsr_out[25] ;
 wire \simon1.lfsr_inst.lfsr_out[26] ;
 wire \simon1.lfsr_inst.lfsr_out[27] ;
 wire \simon1.lfsr_inst.lfsr_out[28] ;
 wire \simon1.lfsr_inst.lfsr_out[29] ;
 wire \simon1.lfsr_inst.lfsr_out[2] ;
 wire \simon1.lfsr_inst.lfsr_out[30] ;
 wire \simon1.lfsr_inst.lfsr_out[31] ;
 wire \simon1.lfsr_inst.lfsr_out[3] ;
 wire \simon1.lfsr_inst.lfsr_out[4] ;
 wire \simon1.lfsr_inst.lfsr_out[5] ;
 wire \simon1.lfsr_inst.lfsr_out[6] ;
 wire \simon1.lfsr_inst.lfsr_out[7] ;
 wire \simon1.lfsr_inst.lfsr_out[8] ;
 wire \simon1.lfsr_inst.lfsr_out[9] ;
 wire \simon1.lfsr_inst.load_enable ;
 wire \simon1.lfsr_stopped ;
 wire \simon1.millis_counter[0] ;
 wire \simon1.millis_counter[1] ;
 wire \simon1.millis_counter[2] ;
 wire \simon1.millis_counter[3] ;
 wire \simon1.millis_counter[4] ;
 wire \simon1.millis_counter[5] ;
 wire \simon1.millis_counter[6] ;
 wire \simon1.millis_counter[7] ;
 wire \simon1.millis_counter[8] ;
 wire \simon1.millis_counter[9] ;
 wire \simon1.prev_btn[0] ;
 wire \simon1.prev_btn[1] ;
 wire \simon1.prev_btn[2] ;
 wire \simon1.prev_btn[3] ;
 wire \simon1.score_ena ;
 wire \simon1.score_inc ;
 wire \simon1.score_inst.active_digit ;
 wire \simon1.score_inst.ones[0] ;
 wire \simon1.score_inst.ones[1] ;
 wire \simon1.score_inst.ones[2] ;
 wire \simon1.score_inst.ones[3] ;
 wire \simon1.score_inst.tens[0] ;
 wire \simon1.score_inst.tens[1] ;
 wire \simon1.score_inst.tens[2] ;
 wire \simon1.score_inst.tens[3] ;
 wire \simon1.score_rst ;
 wire \simon1.seq_counter[0] ;
 wire \simon1.seq_counter[1] ;
 wire \simon1.seq_counter[2] ;
 wire \simon1.seq_counter[3] ;
 wire \simon1.seq_counter[4] ;
 wire \simon1.seq_counter[5] ;
 wire \simon1.seq_counter[6] ;
 wire \simon1.seq_length[0] ;
 wire \simon1.seq_length[1] ;
 wire \simon1.seq_length[2] ;
 wire \simon1.seq_length[3] ;
 wire \simon1.seq_length[4] ;
 wire \simon1.seq_length[5] ;
 wire \simon1.seq_length[6] ;
 wire \simon1.sound ;
 wire \simon1.sound_freq[0] ;
 wire \simon1.sound_freq[1] ;
 wire \simon1.sound_freq[2] ;
 wire \simon1.sound_freq[3] ;
 wire \simon1.sound_freq[4] ;
 wire \simon1.sound_freq[5] ;
 wire \simon1.sound_freq[6] ;
 wire \simon1.sound_freq[7] ;
 wire \simon1.sound_freq[8] ;
 wire \simon1.sound_freq[9] ;
 wire \simon1.sound_gen_inst.tick_counter[0] ;
 wire \simon1.sound_gen_inst.tick_counter[10] ;
 wire \simon1.sound_gen_inst.tick_counter[11] ;
 wire \simon1.sound_gen_inst.tick_counter[12] ;
 wire \simon1.sound_gen_inst.tick_counter[13] ;
 wire \simon1.sound_gen_inst.tick_counter[14] ;
 wire \simon1.sound_gen_inst.tick_counter[15] ;
 wire \simon1.sound_gen_inst.tick_counter[16] ;
 wire \simon1.sound_gen_inst.tick_counter[17] ;
 wire \simon1.sound_gen_inst.tick_counter[18] ;
 wire \simon1.sound_gen_inst.tick_counter[19] ;
 wire \simon1.sound_gen_inst.tick_counter[1] ;
 wire \simon1.sound_gen_inst.tick_counter[20] ;
 wire \simon1.sound_gen_inst.tick_counter[21] ;
 wire \simon1.sound_gen_inst.tick_counter[22] ;
 wire \simon1.sound_gen_inst.tick_counter[23] ;
 wire \simon1.sound_gen_inst.tick_counter[24] ;
 wire \simon1.sound_gen_inst.tick_counter[25] ;
 wire \simon1.sound_gen_inst.tick_counter[26] ;
 wire \simon1.sound_gen_inst.tick_counter[27] ;
 wire \simon1.sound_gen_inst.tick_counter[28] ;
 wire \simon1.sound_gen_inst.tick_counter[29] ;
 wire \simon1.sound_gen_inst.tick_counter[2] ;
 wire \simon1.sound_gen_inst.tick_counter[30] ;
 wire \simon1.sound_gen_inst.tick_counter[31] ;
 wire \simon1.sound_gen_inst.tick_counter[3] ;
 wire \simon1.sound_gen_inst.tick_counter[4] ;
 wire \simon1.sound_gen_inst.tick_counter[5] ;
 wire \simon1.sound_gen_inst.tick_counter[6] ;
 wire \simon1.sound_gen_inst.tick_counter[7] ;
 wire \simon1.sound_gen_inst.tick_counter[8] ;
 wire \simon1.sound_gen_inst.tick_counter[9] ;
 wire \simon1.state[0] ;
 wire \simon1.state[1] ;
 wire \simon1.state[2] ;
 wire \simon1.state[3] ;
 wire \simon1.state[4] ;
 wire \simon1.state[5] ;
 wire \simon1.state[6] ;
 wire \simon1.state[7] ;
 wire \simon1.state[8] ;
 wire \simon1.tick_counter[0] ;
 wire \simon1.tick_counter[10] ;
 wire \simon1.tick_counter[11] ;
 wire \simon1.tick_counter[12] ;
 wire \simon1.tick_counter[13] ;
 wire \simon1.tick_counter[14] ;
 wire \simon1.tick_counter[15] ;
 wire \simon1.tick_counter[1] ;
 wire \simon1.tick_counter[2] ;
 wire \simon1.tick_counter[3] ;
 wire \simon1.tick_counter[4] ;
 wire \simon1.tick_counter[5] ;
 wire \simon1.tick_counter[6] ;
 wire \simon1.tick_counter[7] ;
 wire \simon1.tick_counter[8] ;
 wire \simon1.tick_counter[9] ;
 wire \simon1.tone_sequence_counter[0] ;
 wire \simon1.tone_sequence_counter[1] ;
 wire \simon1.tone_sequence_counter[2] ;
 wire \simon1.user_input[0] ;
 wire \simon1.user_input[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_2 _1612_ (.A(\simon1.tone_sequence_counter[0] ),
    .X(_0933_));
 sg13g2_buf_1 _1613_ (.A(\simon1.tone_sequence_counter[1] ),
    .X(_0934_));
 sg13g2_nand2_1 _1614_ (.Y(_0935_),
    .A(_0933_),
    .B(_0934_));
 sg13g2_or2_1 _1615_ (.X(_0936_),
    .B(_0935_),
    .A(_0026_));
 sg13g2_buf_2 _1616_ (.A(_0936_),
    .X(_0937_));
 sg13g2_buf_1 _1617_ (.A(ui_in[0]),
    .X(_0938_));
 sg13g2_buf_1 _1618_ (.A(ui_in[1]),
    .X(_0939_));
 sg13g2_buf_2 _1619_ (.A(ui_in[2]),
    .X(_0940_));
 sg13g2_buf_2 _1620_ (.A(ui_in[3]),
    .X(_0941_));
 sg13g2_nor3_2 _1621_ (.A(net86),
    .B(_0940_),
    .C(_0941_),
    .Y(_0942_));
 sg13g2_nor2b_2 _1622_ (.A(net87),
    .B_N(_0942_),
    .Y(_0943_));
 sg13g2_buf_1 _1623_ (.A(\simon1.state[1] ),
    .X(_0944_));
 sg13g2_o21ai_1 _1624_ (.B1(_0944_),
    .Y(_0945_),
    .A1(_0937_),
    .A2(_0943_));
 sg13g2_buf_2 _1625_ (.A(\simon1.state[4] ),
    .X(_0946_));
 sg13g2_buf_2 _1626_ (.A(\simon1.lfsr_inst.lfsr_out[1] ),
    .X(_0947_));
 sg13g2_buf_1 _1627_ (.A(\simon1.user_input[1] ),
    .X(_0948_));
 sg13g2_xnor2_1 _1628_ (.Y(_0949_),
    .A(_0947_),
    .B(net83));
 sg13g2_buf_1 _1629_ (.A(\simon1.lfsr_inst.lfsr_out[0] ),
    .X(_0950_));
 sg13g2_buf_1 _1630_ (.A(\simon1.user_input[0] ),
    .X(_0951_));
 sg13g2_xnor2_1 _1631_ (.Y(_0952_),
    .A(net82),
    .B(net81));
 sg13g2_nand2_1 _1632_ (.Y(_0953_),
    .A(_0949_),
    .B(_0952_));
 sg13g2_buf_2 _1633_ (.A(\simon1.millis_counter[2] ),
    .X(_0954_));
 sg13g2_and2_1 _1634_ (.A(_0954_),
    .B(\simon1.millis_counter[5] ),
    .X(_0955_));
 sg13g2_buf_1 _1635_ (.A(\simon1.millis_counter[0] ),
    .X(_0956_));
 sg13g2_buf_2 _1636_ (.A(\simon1.millis_counter[1] ),
    .X(_0957_));
 sg13g2_buf_1 _1637_ (.A(\simon1.millis_counter[8] ),
    .X(_0958_));
 sg13g2_nand2b_1 _1638_ (.Y(_0959_),
    .B(_0958_),
    .A_N(\simon1.millis_counter[9] ));
 sg13g2_nor3_1 _1639_ (.A(net80),
    .B(_0957_),
    .C(_0959_),
    .Y(_0960_));
 sg13g2_buf_1 _1640_ (.A(\simon1.millis_counter[3] ),
    .X(_0961_));
 sg13g2_nor2b_1 _1641_ (.A(\simon1.millis_counter[4] ),
    .B_N(_0961_),
    .Y(_0962_));
 sg13g2_buf_1 _1642_ (.A(\simon1.millis_counter[6] ),
    .X(_0963_));
 sg13g2_nor2_1 _1643_ (.A(\simon1.millis_counter[7] ),
    .B(_0963_),
    .Y(_0964_));
 sg13g2_and4_1 _1644_ (.A(_0955_),
    .B(_0960_),
    .C(_0962_),
    .D(_0964_),
    .X(_0965_));
 sg13g2_buf_1 _1645_ (.A(_0965_),
    .X(_0966_));
 sg13g2_nand3_1 _1646_ (.B(_0953_),
    .C(_0966_),
    .A(_0946_),
    .Y(_0967_));
 sg13g2_buf_1 _1647_ (.A(net1),
    .X(_0968_));
 sg13g2_inv_2 _1648_ (.Y(_0969_),
    .A(net85));
 sg13g2_buf_1 _1649_ (.A(_0969_),
    .X(_0970_));
 sg13g2_buf_1 _1650_ (.A(net61),
    .X(_0971_));
 sg13g2_a21oi_1 _1651_ (.A1(_0945_),
    .A2(_0967_),
    .Y(_0001_),
    .B1(net48));
 sg13g2_buf_1 _1652_ (.A(net85),
    .X(_0972_));
 sg13g2_buf_1 _1653_ (.A(net79),
    .X(_0973_));
 sg13g2_buf_1 _1654_ (.A(\simon1.state[0] ),
    .X(_0974_));
 sg13g2_nand2_1 _1655_ (.Y(_0975_),
    .A(_0974_),
    .B(_0943_));
 sg13g2_nand2_1 _1656_ (.Y(_0000_),
    .A(net60),
    .B(_0975_));
 sg13g2_buf_1 _1657_ (.A(\simon1.seq_counter[0] ),
    .X(_0976_));
 sg13g2_inv_1 _1658_ (.Y(_0977_),
    .A(_0976_));
 sg13g2_buf_2 _1659_ (.A(\simon1.seq_length[0] ),
    .X(_0978_));
 sg13g2_xor2_1 _1660_ (.B(_0027_),
    .A(\simon1.seq_counter[2] ),
    .X(_0979_));
 sg13g2_buf_2 _1661_ (.A(\simon1.seq_counter[1] ),
    .X(_0980_));
 sg13g2_buf_2 _1662_ (.A(\simon1.seq_length[1] ),
    .X(_0981_));
 sg13g2_xnor2_1 _1663_ (.Y(_0982_),
    .A(_0980_),
    .B(_0981_));
 sg13g2_nand4_1 _1664_ (.B(_0978_),
    .C(_0979_),
    .A(_0977_),
    .Y(_0983_),
    .D(_0982_));
 sg13g2_nor2b_1 _1665_ (.A(_0980_),
    .B_N(_0981_),
    .Y(_0984_));
 sg13g2_nor2_1 _1666_ (.A(_0981_),
    .B(_0979_),
    .Y(_0985_));
 sg13g2_a22oi_1 _1667_ (.Y(_0986_),
    .B1(_0985_),
    .B2(_0980_),
    .A2(_0984_),
    .A1(_0979_));
 sg13g2_or3_1 _1668_ (.A(_0977_),
    .B(_0978_),
    .C(_0986_),
    .X(_0987_));
 sg13g2_and3_1 _1669_ (.X(_0988_),
    .A(_0976_),
    .B(_0980_),
    .C(\simon1.seq_counter[2] ));
 sg13g2_buf_2 _1670_ (.A(_0988_),
    .X(_0989_));
 sg13g2_buf_1 _1671_ (.A(\simon1.seq_counter[4] ),
    .X(_0990_));
 sg13g2_xnor2_1 _1672_ (.Y(_0991_),
    .A(_0990_),
    .B(_0029_));
 sg13g2_and3_1 _1673_ (.X(_0992_),
    .A(_0028_),
    .B(_0989_),
    .C(_0991_));
 sg13g2_nor3_1 _1674_ (.A(_0028_),
    .B(_0989_),
    .C(_0991_),
    .Y(_0993_));
 sg13g2_buf_2 _1675_ (.A(\simon1.seq_counter[3] ),
    .X(_0994_));
 sg13g2_o21ai_1 _1676_ (.B1(_0994_),
    .Y(_0995_),
    .A1(_0992_),
    .A2(_0993_));
 sg13g2_xnor2_1 _1677_ (.Y(_0996_),
    .A(_0028_),
    .B(_0989_));
 sg13g2_or3_1 _1678_ (.A(_0994_),
    .B(_0991_),
    .C(_0996_),
    .X(_0997_));
 sg13g2_xor2_1 _1679_ (.B(_0031_),
    .A(\simon1.seq_counter[6] ),
    .X(_0998_));
 sg13g2_inv_1 _1680_ (.Y(_0999_),
    .A(_0030_));
 sg13g2_nand3_1 _1681_ (.B(_0990_),
    .C(_0989_),
    .A(_0994_),
    .Y(_1000_));
 sg13g2_xnor2_1 _1682_ (.Y(_1001_),
    .A(_0999_),
    .B(_1000_));
 sg13g2_nand3_1 _1683_ (.B(_0999_),
    .C(_1000_),
    .A(\simon1.seq_counter[5] ),
    .Y(_1002_));
 sg13g2_o21ai_1 _1684_ (.B1(_1002_),
    .Y(_1003_),
    .A1(\simon1.seq_counter[5] ),
    .A2(_1001_));
 sg13g2_nand4_1 _1685_ (.B(_0990_),
    .C(\simon1.seq_counter[5] ),
    .A(_0994_),
    .Y(_1004_),
    .D(_0989_));
 sg13g2_nor4_1 _1686_ (.A(_0999_),
    .B(\simon1.seq_counter[6] ),
    .C(_0031_),
    .D(_1004_),
    .Y(_1005_));
 sg13g2_a21oi_1 _1687_ (.A1(_0998_),
    .A2(_1003_),
    .Y(_1006_),
    .B1(_1005_));
 sg13g2_a221oi_1 _1688_ (.B2(_0997_),
    .C1(_1006_),
    .B1(_0995_),
    .A1(_0983_),
    .Y(_1007_),
    .A2(_0987_));
 sg13g2_buf_1 _1689_ (.A(_1007_),
    .X(_1008_));
 sg13g2_nand2_1 _1690_ (.Y(_1009_),
    .A(net79),
    .B(net20));
 sg13g2_buf_1 _1691_ (.A(_0946_),
    .X(_1010_));
 sg13g2_nand4_1 _1692_ (.B(_0960_),
    .C(_0962_),
    .A(_0955_),
    .Y(_1011_),
    .D(_0964_));
 sg13g2_nor2_2 _1693_ (.A(_0953_),
    .B(_1011_),
    .Y(_1012_));
 sg13g2_nand2_2 _1694_ (.Y(_1013_),
    .A(net59),
    .B(_1012_));
 sg13g2_inv_1 _1695_ (.Y(_1014_),
    .A(\simon1.millis_counter[4] ));
 sg13g2_inv_1 _1696_ (.Y(_1015_),
    .A(\simon1.millis_counter[7] ));
 sg13g2_nor4_1 _1697_ (.A(_1014_),
    .B(\simon1.millis_counter[5] ),
    .C(_1015_),
    .D(_0963_),
    .Y(_1016_));
 sg13g2_or2_1 _1698_ (.X(_1017_),
    .B(_0958_),
    .A(\simon1.millis_counter[9] ));
 sg13g2_nand2b_1 _1699_ (.Y(_1018_),
    .B(_0957_),
    .A_N(net80));
 sg13g2_nand2b_1 _1700_ (.Y(_1019_),
    .B(_0954_),
    .A_N(_0961_));
 sg13g2_nor3_1 _1701_ (.A(_1017_),
    .B(_1018_),
    .C(_1019_),
    .Y(_1020_));
 sg13g2_nand2_1 _1702_ (.Y(_1021_),
    .A(_1016_),
    .B(_1020_));
 sg13g2_nor2_1 _1703_ (.A(_0937_),
    .B(_1021_),
    .Y(_1022_));
 sg13g2_buf_1 _1704_ (.A(\simon1.state[8] ),
    .X(_1023_));
 sg13g2_buf_1 _1705_ (.A(_1023_),
    .X(_1024_));
 sg13g2_nand3b_1 _1706_ (.B(net79),
    .C(net58),
    .Y(_1025_),
    .A_N(_1022_));
 sg13g2_o21ai_1 _1707_ (.B1(_1025_),
    .Y(_0008_),
    .A1(_1009_),
    .A2(_1013_));
 sg13g2_buf_1 _1708_ (.A(\simon1.state[3] ),
    .X(_1026_));
 sg13g2_inv_1 _1709_ (.Y(_1027_),
    .A(_1026_));
 sg13g2_buf_2 _1710_ (.A(\simon1.state[7] ),
    .X(_1028_));
 sg13g2_nor2_1 _1711_ (.A(_0954_),
    .B(_0961_),
    .Y(_1029_));
 sg13g2_nand3_1 _1712_ (.B(_1016_),
    .C(_1029_),
    .A(_0960_),
    .Y(_1030_));
 sg13g2_nand2_1 _1713_ (.Y(_1031_),
    .A(_1028_),
    .B(_1030_));
 sg13g2_a21oi_1 _1714_ (.A1(_1027_),
    .A2(_1031_),
    .Y(_0007_),
    .B1(net48));
 sg13g2_buf_1 _1715_ (.A(net61),
    .X(_1032_));
 sg13g2_nor2_1 _1716_ (.A(\simon1.millis_counter[5] ),
    .B(_1018_),
    .Y(_1033_));
 sg13g2_xnor2_1 _1717_ (.Y(_1034_),
    .A(net86),
    .B(\simon1.prev_btn[1] ));
 sg13g2_xnor2_1 _1718_ (.Y(_1035_),
    .A(net87),
    .B(\simon1.prev_btn[0] ));
 sg13g2_xnor2_1 _1719_ (.Y(_1036_),
    .A(_0941_),
    .B(\simon1.prev_btn[3] ));
 sg13g2_xnor2_1 _1720_ (.Y(_1037_),
    .A(_0940_),
    .B(\simon1.prev_btn[2] ));
 sg13g2_nand4_1 _1721_ (.B(_1035_),
    .C(_1036_),
    .A(_1034_),
    .Y(_1038_),
    .D(_1037_));
 sg13g2_nand2_1 _1722_ (.Y(_1039_),
    .A(_1014_),
    .B(_0961_));
 sg13g2_nor2_1 _1723_ (.A(_0954_),
    .B(_1039_),
    .Y(_1040_));
 sg13g2_nor3_1 _1724_ (.A(\simon1.millis_counter[7] ),
    .B(_0963_),
    .C(_1017_),
    .Y(_1041_));
 sg13g2_nand4_1 _1725_ (.B(_1038_),
    .C(_1040_),
    .A(_1033_),
    .Y(_1042_),
    .D(_1041_));
 sg13g2_nand2_1 _1726_ (.Y(_1043_),
    .A(\simon1.button_released ),
    .B(_0943_));
 sg13g2_nor2_1 _1727_ (.A(net20),
    .B(_1013_),
    .Y(_1044_));
 sg13g2_a22oi_1 _1728_ (.Y(_1045_),
    .B1(_1043_),
    .B2(_1044_),
    .A2(_1042_),
    .A1(\simon1.state[6] ));
 sg13g2_nor2_1 _1729_ (.A(net47),
    .B(_1045_),
    .Y(_0006_));
 sg13g2_nor2_1 _1730_ (.A(net80),
    .B(_0957_),
    .Y(_1046_));
 sg13g2_nand3b_1 _1731_ (.B(_0958_),
    .C(_1046_),
    .Y(_1047_),
    .A_N(\simon1.millis_counter[9] ));
 sg13g2_nand2_1 _1732_ (.Y(_1048_),
    .A(\simon1.millis_counter[4] ),
    .B(\simon1.millis_counter[5] ));
 sg13g2_nand2_1 _1733_ (.Y(_1049_),
    .A(\simon1.millis_counter[7] ),
    .B(_0963_));
 sg13g2_nor4_1 _1734_ (.A(_1047_),
    .B(_1019_),
    .C(_1048_),
    .D(_1049_),
    .Y(_1050_));
 sg13g2_buf_1 _1735_ (.A(\simon1.state[5] ),
    .X(_1051_));
 sg13g2_nand2b_1 _1736_ (.Y(_1052_),
    .B(_1051_),
    .A_N(_1050_));
 sg13g2_inv_1 _1737_ (.Y(_1053_),
    .A(_0944_));
 sg13g2_nor2_1 _1738_ (.A(_1053_),
    .B(_0937_),
    .Y(_1054_));
 sg13g2_nand2b_2 _1739_ (.Y(_1055_),
    .B(_0942_),
    .A_N(net87));
 sg13g2_o21ai_1 _1740_ (.B1(_1055_),
    .Y(_1056_),
    .A1(_0974_),
    .A2(_1054_));
 sg13g2_a21oi_1 _1741_ (.A1(_1052_),
    .A2(_1056_),
    .Y(_0005_),
    .B1(net48));
 sg13g2_xor2_1 _1742_ (.B(_0941_),
    .A(_0940_),
    .X(_1057_));
 sg13g2_o21ai_1 _1743_ (.B1(net86),
    .Y(_1058_),
    .A1(_0940_),
    .A2(_0941_));
 sg13g2_o21ai_1 _1744_ (.B1(_1058_),
    .Y(_1059_),
    .A1(net86),
    .A2(_1057_));
 sg13g2_nor2_1 _1745_ (.A(net87),
    .B(_1059_),
    .Y(_1060_));
 sg13g2_a21oi_1 _1746_ (.A1(net87),
    .A2(_0942_),
    .Y(_1061_),
    .B1(_1060_));
 sg13g2_buf_1 _1747_ (.A(\simon1.state[2] ),
    .X(_1062_));
 sg13g2_nand2_2 _1748_ (.Y(_1063_),
    .A(_1062_),
    .B(_1055_));
 sg13g2_nand2_2 _1749_ (.Y(_1064_),
    .A(_0946_),
    .B(_1011_));
 sg13g2_o21ai_1 _1750_ (.B1(_1064_),
    .Y(_1065_),
    .A1(_1061_),
    .A2(_1063_));
 sg13g2_and2_1 _1751_ (.A(net60),
    .B(_1065_),
    .X(_0004_));
 sg13g2_nor4_1 _1752_ (.A(_1047_),
    .B(_1019_),
    .C(_1048_),
    .D(_1049_),
    .Y(_1066_));
 sg13g2_inv_1 _1753_ (.Y(_1067_),
    .A(_1028_));
 sg13g2_nor2_1 _1754_ (.A(_1067_),
    .B(_1030_),
    .Y(_1068_));
 sg13g2_inv_1 _1755_ (.Y(_1069_),
    .A(_1068_));
 sg13g2_nor2_1 _1756_ (.A(_1008_),
    .B(_1069_),
    .Y(_1070_));
 sg13g2_a221oi_1 _1757_ (.B2(_1051_),
    .C1(_1070_),
    .B1(_1066_),
    .A1(net58),
    .Y(_1071_),
    .A2(_1022_));
 sg13g2_nor2_1 _1758_ (.A(net47),
    .B(_1071_),
    .Y(_0003_));
 sg13g2_or2_1 _1759_ (.X(_1072_),
    .B(_1013_),
    .A(net20));
 sg13g2_inv_1 _1760_ (.Y(_1073_),
    .A(\simon1.state[6] ));
 sg13g2_nor2_1 _1761_ (.A(_1073_),
    .B(_1042_),
    .Y(_1074_));
 sg13g2_a221oi_1 _1762_ (.B2(net20),
    .C1(_1074_),
    .B1(_1068_),
    .A1(net78),
    .Y(_1075_),
    .A2(_1061_));
 sg13g2_o21ai_1 _1763_ (.B1(_1075_),
    .Y(_1076_),
    .A1(_1043_),
    .A2(_1072_));
 sg13g2_and2_1 _1764_ (.A(net60),
    .B(_1076_),
    .X(_0002_));
 sg13g2_buf_4 _1765_ (.X(_1077_),
    .A(ui_in[4]));
 sg13g2_buf_1 _1766_ (.A(\simon1.score_inst.active_digit ),
    .X(_1078_));
 sg13g2_xor2_1 _1767_ (.B(_1078_),
    .A(_1077_),
    .X(_0011_));
 sg13g2_inv_1 _1768_ (.Y(_0010_),
    .A(_0011_));
 sg13g2_buf_2 _1769_ (.A(\simon1.score_inst.ones[1] ),
    .X(_1079_));
 sg13g2_nand2b_1 _1770_ (.Y(_1080_),
    .B(_1079_),
    .A_N(net77));
 sg13g2_buf_1 _1771_ (.A(\simon1.score_inst.tens[1] ),
    .X(_1081_));
 sg13g2_nand2_1 _1772_ (.Y(_1082_),
    .A(net77),
    .B(_1081_));
 sg13g2_nand3_1 _1773_ (.B(_1080_),
    .C(_1082_),
    .A(\simon1.score_ena ),
    .Y(_1083_));
 sg13g2_buf_2 _1774_ (.A(_1083_),
    .X(_1084_));
 sg13g2_inv_1 _1775_ (.Y(_1085_),
    .A(_1084_));
 sg13g2_inv_1 _1776_ (.Y(_1086_),
    .A(\simon1.score_inst.tens[2] ));
 sg13g2_nor2_1 _1777_ (.A(\simon1.score_inst.ones[2] ),
    .B(net77),
    .Y(_1087_));
 sg13g2_a21oi_1 _1778_ (.A1(net77),
    .A2(_1086_),
    .Y(_1088_),
    .B1(_1087_));
 sg13g2_or2_1 _1779_ (.X(_1089_),
    .B(_1088_),
    .A(_0014_));
 sg13g2_buf_2 _1780_ (.A(_1089_),
    .X(_1090_));
 sg13g2_inv_1 _1781_ (.Y(_1091_),
    .A(\simon1.score_inst.ones[3] ));
 sg13g2_nand2_1 _1782_ (.Y(_1092_),
    .A(net77),
    .B(\simon1.score_inst.tens[3] ));
 sg13g2_o21ai_1 _1783_ (.B1(_1092_),
    .Y(_1093_),
    .A1(_1091_),
    .A2(net77));
 sg13g2_nor3_1 _1784_ (.A(_0014_),
    .B(_1093_),
    .C(_1088_),
    .Y(_1094_));
 sg13g2_nand2b_1 _1785_ (.Y(_1095_),
    .B(\simon1.score_inst.ones[0] ),
    .A_N(net77));
 sg13g2_nand2_1 _1786_ (.Y(_1096_),
    .A(net77),
    .B(\simon1.score_inst.tens[0] ));
 sg13g2_nand3_1 _1787_ (.B(_1095_),
    .C(_1096_),
    .A(\simon1.score_ena ),
    .Y(_1097_));
 sg13g2_buf_2 _1788_ (.A(_1097_),
    .X(_1098_));
 sg13g2_mux2_1 _1789_ (.A0(_1090_),
    .A1(_1094_),
    .S(_1098_),
    .X(_1099_));
 sg13g2_nor2_2 _1790_ (.A(_0014_),
    .B(_1093_),
    .Y(_1100_));
 sg13g2_nor2_2 _1791_ (.A(_1090_),
    .B(_1084_),
    .Y(_1101_));
 sg13g2_nor2_1 _1792_ (.A(_1100_),
    .B(_1101_),
    .Y(_1102_));
 sg13g2_a21oi_1 _1793_ (.A1(_1085_),
    .A2(_1099_),
    .Y(_1103_),
    .B1(_1102_));
 sg13g2_xor2_1 _1794_ (.B(_1103_),
    .A(_1077_),
    .X(_0213_));
 sg13g2_xor2_1 _1795_ (.B(_1098_),
    .A(_1084_),
    .X(_1104_));
 sg13g2_a21oi_1 _1796_ (.A1(_1090_),
    .A2(_1104_),
    .Y(_1105_),
    .B1(_1102_));
 sg13g2_xor2_1 _1797_ (.B(_1105_),
    .A(_1077_),
    .X(_0214_));
 sg13g2_o21ai_1 _1798_ (.B1(_1100_),
    .Y(_1106_),
    .A1(_1090_),
    .A2(_1098_));
 sg13g2_nor2b_1 _1799_ (.A(_1101_),
    .B_N(_1106_),
    .Y(_1107_));
 sg13g2_xnor2_1 _1800_ (.Y(_0215_),
    .A(_1077_),
    .B(_1107_));
 sg13g2_nand2_1 _1801_ (.Y(_1108_),
    .A(_1090_),
    .B(_1084_));
 sg13g2_nand2_1 _1802_ (.Y(_1109_),
    .A(_1100_),
    .B(_1101_));
 sg13g2_nand2_1 _1803_ (.Y(_1110_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_nor2_1 _1804_ (.A(_1084_),
    .B(_1098_),
    .Y(_1111_));
 sg13g2_a221oi_1 _1805_ (.B2(_1090_),
    .C1(_1102_),
    .B1(_1111_),
    .A1(_1098_),
    .Y(_1112_),
    .A2(_1110_));
 sg13g2_xor2_1 _1806_ (.B(_1112_),
    .A(_1077_),
    .X(_0216_));
 sg13g2_a21oi_1 _1807_ (.A1(_1100_),
    .A2(_1084_),
    .Y(_1113_),
    .B1(_1101_));
 sg13g2_nor2_1 _1808_ (.A(_1098_),
    .B(_1113_),
    .Y(_1114_));
 sg13g2_xor2_1 _1809_ (.B(_1114_),
    .A(_1077_),
    .X(_0217_));
 sg13g2_and2_1 _1810_ (.A(_1100_),
    .B(_1090_),
    .X(_1115_));
 sg13g2_o21ai_1 _1811_ (.B1(_1098_),
    .Y(_1116_),
    .A1(_1084_),
    .A2(_1094_));
 sg13g2_o21ai_1 _1812_ (.B1(_1116_),
    .Y(_1117_),
    .A1(_1101_),
    .A2(_1115_));
 sg13g2_xnor2_1 _1813_ (.Y(_0218_),
    .A(_1077_),
    .B(_1117_));
 sg13g2_nand3_1 _1814_ (.B(_1084_),
    .C(_1098_),
    .A(_1090_),
    .Y(_1118_));
 sg13g2_nand3b_1 _1815_ (.B(_1109_),
    .C(_1118_),
    .Y(_1119_),
    .A_N(_1102_));
 sg13g2_xnor2_1 _1816_ (.Y(_0219_),
    .A(_1077_),
    .B(_1119_));
 sg13g2_inv_1 _1817_ (.Y(_1120_),
    .A(_0933_));
 sg13g2_buf_1 _1818_ (.A(\simon1.tone_sequence_counter[2] ),
    .X(_1121_));
 sg13g2_inv_1 _1819_ (.Y(_1122_),
    .A(net76));
 sg13g2_nor2_2 _1820_ (.A(_0933_),
    .B(_0934_),
    .Y(_1123_));
 sg13g2_nand2_2 _1821_ (.Y(_1124_),
    .A(\simon1.tone_sequence_counter[2] ),
    .B(_1123_));
 sg13g2_nand2_1 _1822_ (.Y(_1125_),
    .A(_0944_),
    .B(_1124_));
 sg13g2_a21oi_1 _1823_ (.A1(_1122_),
    .A2(_0966_),
    .Y(_1126_),
    .B1(_1125_));
 sg13g2_nand3_1 _1824_ (.B(_0958_),
    .C(\simon1.millis_counter[5] ),
    .A(\simon1.millis_counter[9] ),
    .Y(_1127_));
 sg13g2_nand3_1 _1825_ (.B(_0963_),
    .C(_1046_),
    .A(\simon1.millis_counter[7] ),
    .Y(_1128_));
 sg13g2_nor4_2 _1826_ (.A(_0954_),
    .B(_1039_),
    .C(_1127_),
    .Y(_1129_),
    .D(_1128_));
 sg13g2_inv_1 _1827_ (.Y(_1130_),
    .A(_1124_));
 sg13g2_nand2b_1 _1828_ (.Y(_1131_),
    .B(_1130_),
    .A_N(_1129_));
 sg13g2_nor2_1 _1829_ (.A(_0033_),
    .B(_1131_),
    .Y(_1132_));
 sg13g2_and2_1 _1830_ (.A(_1023_),
    .B(_1021_),
    .X(_1133_));
 sg13g2_nand2_1 _1831_ (.Y(_1134_),
    .A(_1053_),
    .B(_0032_));
 sg13g2_o21ai_1 _1832_ (.B1(net1),
    .Y(_1135_),
    .A1(_1051_),
    .A2(_1134_));
 sg13g2_nor4_2 _1833_ (.A(_1126_),
    .B(_1132_),
    .C(_1133_),
    .Y(_1136_),
    .D(_1135_));
 sg13g2_nor2_1 _1834_ (.A(_0944_),
    .B(_1023_),
    .Y(_1137_));
 sg13g2_nor2_1 _1835_ (.A(_0933_),
    .B(_1137_),
    .Y(_1138_));
 sg13g2_nand2_1 _1836_ (.Y(_1139_),
    .A(_1136_),
    .B(_1138_));
 sg13g2_o21ai_1 _1837_ (.B1(_1139_),
    .Y(_0208_),
    .A1(_1120_),
    .A2(_1136_));
 sg13g2_inv_1 _1838_ (.Y(_1140_),
    .A(net84));
 sg13g2_nor2_1 _1839_ (.A(_1122_),
    .B(_0033_),
    .Y(_1141_));
 sg13g2_o21ai_1 _1840_ (.B1(_1136_),
    .Y(_1142_),
    .A1(_0933_),
    .A2(_1141_));
 sg13g2_inv_1 _1841_ (.Y(_1143_),
    .A(_0033_));
 sg13g2_a21oi_1 _1842_ (.A1(_0944_),
    .A2(_1143_),
    .Y(_1144_),
    .B1(net58));
 sg13g2_a21o_1 _1843_ (.A2(net84),
    .A1(_0933_),
    .B1(_1144_),
    .X(_1145_));
 sg13g2_a22oi_1 _1844_ (.Y(_0209_),
    .B1(_1145_),
    .B2(_1136_),
    .A2(_1142_),
    .A1(_1140_));
 sg13g2_nand2_1 _1845_ (.Y(_1146_),
    .A(_0026_),
    .B(_0935_));
 sg13g2_a22oi_1 _1846_ (.Y(_1147_),
    .B1(_1146_),
    .B2(_0937_),
    .A2(_1141_),
    .A1(_1123_));
 sg13g2_nor2_1 _1847_ (.A(_1144_),
    .B(_1147_),
    .Y(_1148_));
 sg13g2_nand2_1 _1848_ (.Y(_1149_),
    .A(_1136_),
    .B(_1148_));
 sg13g2_o21ai_1 _1849_ (.B1(_1149_),
    .Y(_0210_),
    .A1(_1122_),
    .A2(_1136_));
 sg13g2_nor4_1 _1850_ (.A(\simon1.lfsr_inst.lfsr_out[19] ),
    .B(\simon1.lfsr_inst.lfsr_out[22] ),
    .C(\simon1.lfsr_inst.lfsr_out[25] ),
    .D(\simon1.lfsr_inst.lfsr_out[27] ),
    .Y(_1150_));
 sg13g2_nor4_1 _1851_ (.A(\simon1.lfsr_inst.lfsr_out[18] ),
    .B(\simon1.lfsr_inst.lfsr_out[21] ),
    .C(\simon1.lfsr_inst.lfsr_out[20] ),
    .D(\simon1.lfsr_inst.lfsr_out[23] ),
    .Y(_1151_));
 sg13g2_nor4_1 _1852_ (.A(\simon1.lfsr_inst.lfsr_out[3] ),
    .B(\simon1.lfsr_inst.lfsr_out[2] ),
    .C(\simon1.lfsr_inst.lfsr_out[24] ),
    .D(\simon1.lfsr_inst.lfsr_out[30] ),
    .Y(_1152_));
 sg13g2_nor4_1 _1853_ (.A(\simon1.lfsr_inst.lfsr_out[26] ),
    .B(\simon1.lfsr_inst.lfsr_out[29] ),
    .C(\simon1.lfsr_inst.lfsr_out[28] ),
    .D(\simon1.lfsr_inst.lfsr_out[31] ),
    .Y(_1153_));
 sg13g2_nand4_1 _1854_ (.B(_1151_),
    .C(_1152_),
    .A(_1150_),
    .Y(_1154_),
    .D(_1153_));
 sg13g2_nor4_1 _1855_ (.A(\simon1.lfsr_inst.lfsr_out[9] ),
    .B(\simon1.lfsr_inst.lfsr_out[8] ),
    .C(\simon1.lfsr_inst.lfsr_out[10] ),
    .D(\simon1.lfsr_inst.lfsr_out[16] ),
    .Y(_1155_));
 sg13g2_nor4_1 _1856_ (.A(\simon1.lfsr_inst.lfsr_out[5] ),
    .B(\simon1.lfsr_inst.lfsr_out[4] ),
    .C(\simon1.lfsr_inst.lfsr_out[7] ),
    .D(\simon1.lfsr_inst.lfsr_out[6] ),
    .Y(_1156_));
 sg13g2_nor4_1 _1857_ (.A(\simon1.lfsr_inst.lfsr_out[13] ),
    .B(\simon1.lfsr_inst.lfsr_out[12] ),
    .C(\simon1.lfsr_inst.lfsr_out[15] ),
    .D(\simon1.lfsr_inst.lfsr_out[14] ),
    .Y(_1157_));
 sg13g2_nor4_1 _1858_ (.A(net82),
    .B(_0947_),
    .C(\simon1.lfsr_inst.lfsr_out[11] ),
    .D(\simon1.lfsr_inst.lfsr_out[17] ),
    .Y(_1158_));
 sg13g2_nand4_1 _1859_ (.B(_1156_),
    .C(_1157_),
    .A(_1155_),
    .Y(_1159_),
    .D(_1158_));
 sg13g2_o21ai_1 _1860_ (.B1(net1),
    .Y(_1160_),
    .A1(_1154_),
    .A2(_1159_));
 sg13g2_buf_1 _1861_ (.A(_1160_),
    .X(_1161_));
 sg13g2_buf_1 _1862_ (.A(_1161_),
    .X(_1162_));
 sg13g2_buf_1 _1863_ (.A(\simon1.lfsr_inst.load_enable ),
    .X(_1163_));
 sg13g2_buf_1 _1864_ (.A(_1163_),
    .X(_1164_));
 sg13g2_buf_1 _1865_ (.A(net57),
    .X(_1165_));
 sg13g2_inv_1 _1866_ (.Y(_1166_),
    .A(\simon1.lfsr_stopped ));
 sg13g2_nor3_1 _1867_ (.A(\simon1.lfsr_cycles[0] ),
    .B(\simon1.lfsr_cycles[1] ),
    .C(_1166_),
    .Y(_1167_));
 sg13g2_inv_2 _1868_ (.Y(_1168_),
    .A(_0947_));
 sg13g2_xnor2_1 _1869_ (.Y(_1169_),
    .A(\simon1.lfsr_inst.lfsr_out[21] ),
    .B(\simon1.lfsr_inst.lfsr_out[31] ));
 sg13g2_xnor2_1 _1870_ (.Y(_1170_),
    .A(_1168_),
    .B(_1169_));
 sg13g2_nor2_1 _1871_ (.A(_1167_),
    .B(_1170_),
    .Y(_1171_));
 sg13g2_xnor2_1 _1872_ (.Y(_1172_),
    .A(net82),
    .B(_1171_));
 sg13g2_nor2_1 _1873_ (.A(net46),
    .B(_1172_),
    .Y(_1173_));
 sg13g2_a21oi_1 _1874_ (.A1(net46),
    .A2(\simon1.lfsr_capture[0] ),
    .Y(_1174_),
    .B1(_1173_));
 sg13g2_nor2_1 _1875_ (.A(net30),
    .B(_1174_),
    .Y(_0075_));
 sg13g2_buf_1 _1876_ (.A(_1161_),
    .X(_1175_));
 sg13g2_nand2b_1 _1877_ (.Y(_1176_),
    .B(_1167_),
    .A_N(_1163_));
 sg13g2_buf_1 _1878_ (.A(_1176_),
    .X(_1177_));
 sg13g2_buf_1 _1879_ (.A(net41),
    .X(_1178_));
 sg13g2_nor2_1 _1880_ (.A(\simon1.lfsr_inst.lfsr_out[10] ),
    .B(net39),
    .Y(_1179_));
 sg13g2_nor2b_1 _1881_ (.A(_1163_),
    .B_N(_1167_),
    .Y(_1180_));
 sg13g2_buf_2 _1882_ (.A(_1180_),
    .X(_1181_));
 sg13g2_buf_1 _1883_ (.A(_1181_),
    .X(_1182_));
 sg13g2_mux2_1 _1884_ (.A0(\simon1.lfsr_inst.lfsr_out[9] ),
    .A1(\simon1.lfsr_capture[10] ),
    .S(net46),
    .X(_1183_));
 sg13g2_nor2_1 _1885_ (.A(net38),
    .B(_1183_),
    .Y(_1184_));
 sg13g2_nor3_1 _1886_ (.A(_1175_),
    .B(_1179_),
    .C(_1184_),
    .Y(_0076_));
 sg13g2_buf_1 _1887_ (.A(net41),
    .X(_1185_));
 sg13g2_buf_1 _1888_ (.A(net41),
    .X(_1186_));
 sg13g2_buf_1 _1889_ (.A(_1163_),
    .X(_1187_));
 sg13g2_buf_1 _1890_ (.A(_1163_),
    .X(_1188_));
 sg13g2_nand2b_1 _1891_ (.Y(_1189_),
    .B(net55),
    .A_N(\simon1.lfsr_capture[11] ));
 sg13g2_o21ai_1 _1892_ (.B1(_1189_),
    .Y(_1190_),
    .A1(net56),
    .A2(\simon1.lfsr_inst.lfsr_out[10] ));
 sg13g2_nand2_1 _1893_ (.Y(_1191_),
    .A(net36),
    .B(_1190_));
 sg13g2_o21ai_1 _1894_ (.B1(_1191_),
    .Y(_1192_),
    .A1(\simon1.lfsr_inst.lfsr_out[11] ),
    .A2(net37));
 sg13g2_nand2b_1 _1895_ (.Y(_0077_),
    .B(_1192_),
    .A_N(_1162_));
 sg13g2_buf_1 _1896_ (.A(_1163_),
    .X(_1193_));
 sg13g2_nand2b_1 _1897_ (.Y(_1194_),
    .B(net55),
    .A_N(\simon1.lfsr_capture[12] ));
 sg13g2_o21ai_1 _1898_ (.B1(_1194_),
    .Y(_1195_),
    .A1(net54),
    .A2(\simon1.lfsr_inst.lfsr_out[11] ));
 sg13g2_nand2_1 _1899_ (.Y(_1196_),
    .A(net36),
    .B(_1195_));
 sg13g2_o21ai_1 _1900_ (.B1(_1196_),
    .Y(_1197_),
    .A1(\simon1.lfsr_inst.lfsr_out[12] ),
    .A2(net37));
 sg13g2_nand2b_1 _1901_ (.Y(_0078_),
    .B(_1197_),
    .A_N(_1162_));
 sg13g2_nand2b_1 _1902_ (.Y(_1198_),
    .B(net55),
    .A_N(\simon1.lfsr_capture[13] ));
 sg13g2_o21ai_1 _1903_ (.B1(_1198_),
    .Y(_1199_),
    .A1(net54),
    .A2(\simon1.lfsr_inst.lfsr_out[12] ));
 sg13g2_nand2_1 _1904_ (.Y(_1200_),
    .A(net36),
    .B(_1199_));
 sg13g2_o21ai_1 _1905_ (.B1(_1200_),
    .Y(_1201_),
    .A1(\simon1.lfsr_inst.lfsr_out[13] ),
    .A2(net37));
 sg13g2_nand2b_1 _1906_ (.Y(_0079_),
    .B(_1201_),
    .A_N(net30));
 sg13g2_nand2b_1 _1907_ (.Y(_1202_),
    .B(net55),
    .A_N(\simon1.lfsr_capture[14] ));
 sg13g2_o21ai_1 _1908_ (.B1(_1202_),
    .Y(_1203_),
    .A1(net54),
    .A2(\simon1.lfsr_inst.lfsr_out[13] ));
 sg13g2_nand2_1 _1909_ (.Y(_1204_),
    .A(_1186_),
    .B(_1203_));
 sg13g2_o21ai_1 _1910_ (.B1(_1204_),
    .Y(_1205_),
    .A1(\simon1.lfsr_inst.lfsr_out[14] ),
    .A2(_1185_));
 sg13g2_nand2b_1 _1911_ (.Y(_0080_),
    .B(_1205_),
    .A_N(net30));
 sg13g2_nand2b_1 _1912_ (.Y(_1206_),
    .B(_1188_),
    .A_N(\simon1.lfsr_capture[15] ));
 sg13g2_o21ai_1 _1913_ (.B1(_1206_),
    .Y(_1207_),
    .A1(net54),
    .A2(\simon1.lfsr_inst.lfsr_out[14] ));
 sg13g2_nand2_1 _1914_ (.Y(_1208_),
    .A(_1186_),
    .B(_1207_));
 sg13g2_o21ai_1 _1915_ (.B1(_1208_),
    .Y(_1209_),
    .A1(\simon1.lfsr_inst.lfsr_out[15] ),
    .A2(_1185_));
 sg13g2_nand2b_1 _1916_ (.Y(_0081_),
    .B(_1209_),
    .A_N(net30));
 sg13g2_nor2_1 _1917_ (.A(\simon1.lfsr_inst.lfsr_out[16] ),
    .B(net39),
    .Y(_1210_));
 sg13g2_mux2_1 _1918_ (.A0(\simon1.lfsr_inst.lfsr_out[15] ),
    .A1(\simon1.lfsr_capture[16] ),
    .S(net46),
    .X(_1211_));
 sg13g2_nor2_1 _1919_ (.A(net38),
    .B(_1211_),
    .Y(_1212_));
 sg13g2_nor3_1 _1920_ (.A(_1175_),
    .B(_1210_),
    .C(_1212_),
    .Y(_0082_));
 sg13g2_nor2_1 _1921_ (.A(\simon1.lfsr_inst.lfsr_out[17] ),
    .B(net39),
    .Y(_1213_));
 sg13g2_mux2_1 _1922_ (.A0(\simon1.lfsr_inst.lfsr_out[16] ),
    .A1(\simon1.lfsr_capture[17] ),
    .S(net46),
    .X(_1214_));
 sg13g2_nor2_1 _1923_ (.A(net38),
    .B(_1214_),
    .Y(_1215_));
 sg13g2_nor3_1 _1924_ (.A(net29),
    .B(_1213_),
    .C(_1215_),
    .Y(_0083_));
 sg13g2_buf_1 _1925_ (.A(_1161_),
    .X(_1216_));
 sg13g2_nor2_1 _1926_ (.A(\simon1.lfsr_inst.lfsr_out[18] ),
    .B(_1178_),
    .Y(_1217_));
 sg13g2_mux2_1 _1927_ (.A0(\simon1.lfsr_inst.lfsr_out[17] ),
    .A1(\simon1.lfsr_capture[18] ),
    .S(net46),
    .X(_1218_));
 sg13g2_nor2_1 _1928_ (.A(net38),
    .B(_1218_),
    .Y(_1219_));
 sg13g2_nor3_1 _1929_ (.A(net28),
    .B(_1217_),
    .C(_1219_),
    .Y(_0084_));
 sg13g2_nand2b_1 _1930_ (.Y(_1220_),
    .B(_1188_),
    .A_N(\simon1.lfsr_capture[19] ));
 sg13g2_o21ai_1 _1931_ (.B1(_1220_),
    .Y(_1221_),
    .A1(_1193_),
    .A2(\simon1.lfsr_inst.lfsr_out[18] ));
 sg13g2_nand2_1 _1932_ (.Y(_1222_),
    .A(net36),
    .B(_1221_));
 sg13g2_o21ai_1 _1933_ (.B1(_1222_),
    .Y(_1223_),
    .A1(\simon1.lfsr_inst.lfsr_out[19] ),
    .A2(net37));
 sg13g2_nand2b_1 _1934_ (.Y(_0085_),
    .B(_1223_),
    .A_N(net30));
 sg13g2_nand2b_1 _1935_ (.Y(_1224_),
    .B(_1164_),
    .A_N(\simon1.lfsr_capture[1] ));
 sg13g2_o21ai_1 _1936_ (.B1(_1224_),
    .Y(_1225_),
    .A1(net82),
    .A2(net56));
 sg13g2_nand2_1 _1937_ (.Y(_1226_),
    .A(net36),
    .B(_1225_));
 sg13g2_o21ai_1 _1938_ (.B1(_1226_),
    .Y(_1227_),
    .A1(_0947_),
    .A2(net37));
 sg13g2_nand2b_1 _1939_ (.Y(_0086_),
    .B(_1227_),
    .A_N(net30));
 sg13g2_nor2_1 _1940_ (.A(\simon1.lfsr_inst.lfsr_out[20] ),
    .B(_1178_),
    .Y(_1228_));
 sg13g2_mux2_1 _1941_ (.A0(\simon1.lfsr_inst.lfsr_out[19] ),
    .A1(\simon1.lfsr_capture[20] ),
    .S(net46),
    .X(_1229_));
 sg13g2_nor2_1 _1942_ (.A(net38),
    .B(_1229_),
    .Y(_1230_));
 sg13g2_nor3_1 _1943_ (.A(_1216_),
    .B(_1228_),
    .C(_1230_),
    .Y(_0087_));
 sg13g2_buf_1 _1944_ (.A(_1177_),
    .X(_1231_));
 sg13g2_nor2_1 _1945_ (.A(\simon1.lfsr_inst.lfsr_out[21] ),
    .B(net35),
    .Y(_1232_));
 sg13g2_mux2_1 _1946_ (.A0(\simon1.lfsr_inst.lfsr_out[20] ),
    .A1(\simon1.lfsr_capture[21] ),
    .S(_1165_),
    .X(_1233_));
 sg13g2_nor2_1 _1947_ (.A(_1182_),
    .B(_1233_),
    .Y(_1234_));
 sg13g2_nor3_1 _1948_ (.A(_1216_),
    .B(_1232_),
    .C(_1234_),
    .Y(_0088_));
 sg13g2_nand2b_1 _1949_ (.Y(_1235_),
    .B(_1164_),
    .A_N(\simon1.lfsr_capture[22] ));
 sg13g2_o21ai_1 _1950_ (.B1(_1235_),
    .Y(_1236_),
    .A1(_1193_),
    .A2(\simon1.lfsr_inst.lfsr_out[21] ));
 sg13g2_nand2_1 _1951_ (.Y(_1237_),
    .A(net36),
    .B(_1236_));
 sg13g2_o21ai_1 _1952_ (.B1(_1237_),
    .Y(_1238_),
    .A1(\simon1.lfsr_inst.lfsr_out[22] ),
    .A2(net37));
 sg13g2_nand2b_1 _1953_ (.Y(_0089_),
    .B(_1238_),
    .A_N(net30));
 sg13g2_nor2_1 _1954_ (.A(\simon1.lfsr_inst.lfsr_out[23] ),
    .B(net35),
    .Y(_1239_));
 sg13g2_mux2_1 _1955_ (.A0(\simon1.lfsr_inst.lfsr_out[22] ),
    .A1(\simon1.lfsr_capture[23] ),
    .S(_1165_),
    .X(_1240_));
 sg13g2_nor2_1 _1956_ (.A(_1182_),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_nor3_1 _1957_ (.A(net28),
    .B(_1239_),
    .C(_1241_),
    .Y(_0090_));
 sg13g2_nor2_1 _1958_ (.A(\simon1.lfsr_inst.lfsr_out[24] ),
    .B(_1231_),
    .Y(_1242_));
 sg13g2_mux2_1 _1959_ (.A0(\simon1.lfsr_inst.lfsr_out[23] ),
    .A1(\simon1.lfsr_capture[24] ),
    .S(_1187_),
    .X(_1243_));
 sg13g2_nor2_1 _1960_ (.A(net38),
    .B(_1243_),
    .Y(_1244_));
 sg13g2_nor3_1 _1961_ (.A(net28),
    .B(_1242_),
    .C(_1244_),
    .Y(_0091_));
 sg13g2_nor2_1 _1962_ (.A(\simon1.lfsr_inst.lfsr_out[25] ),
    .B(_1231_),
    .Y(_1245_));
 sg13g2_mux2_1 _1963_ (.A0(\simon1.lfsr_inst.lfsr_out[24] ),
    .A1(\simon1.lfsr_capture[25] ),
    .S(net56),
    .X(_1246_));
 sg13g2_nor2_1 _1964_ (.A(net38),
    .B(_1246_),
    .Y(_1247_));
 sg13g2_nor3_1 _1965_ (.A(net28),
    .B(_1245_),
    .C(_1247_),
    .Y(_0092_));
 sg13g2_nor2_1 _1966_ (.A(\simon1.lfsr_inst.lfsr_out[26] ),
    .B(net35),
    .Y(_1248_));
 sg13g2_mux2_1 _1967_ (.A0(\simon1.lfsr_inst.lfsr_out[25] ),
    .A1(\simon1.lfsr_capture[26] ),
    .S(_1187_),
    .X(_1249_));
 sg13g2_nor2_1 _1968_ (.A(net38),
    .B(_1249_),
    .Y(_1250_));
 sg13g2_nor3_1 _1969_ (.A(net28),
    .B(_1248_),
    .C(_1250_),
    .Y(_0093_));
 sg13g2_nor2_1 _1970_ (.A(\simon1.lfsr_inst.lfsr_out[27] ),
    .B(net35),
    .Y(_1251_));
 sg13g2_mux2_1 _1971_ (.A0(\simon1.lfsr_inst.lfsr_out[26] ),
    .A1(\simon1.lfsr_capture[27] ),
    .S(net56),
    .X(_1252_));
 sg13g2_nor2_1 _1972_ (.A(_1181_),
    .B(_1252_),
    .Y(_1253_));
 sg13g2_nor3_1 _1973_ (.A(net28),
    .B(_1251_),
    .C(_1253_),
    .Y(_0094_));
 sg13g2_nor2_1 _1974_ (.A(\simon1.lfsr_inst.lfsr_out[28] ),
    .B(net35),
    .Y(_1254_));
 sg13g2_mux2_1 _1975_ (.A0(\simon1.lfsr_inst.lfsr_out[27] ),
    .A1(\simon1.lfsr_capture[28] ),
    .S(net56),
    .X(_1255_));
 sg13g2_nor2_1 _1976_ (.A(_1181_),
    .B(_1255_),
    .Y(_1256_));
 sg13g2_nor3_1 _1977_ (.A(net28),
    .B(_1254_),
    .C(_1256_),
    .Y(_0095_));
 sg13g2_nand2b_1 _1978_ (.Y(_1257_),
    .B(net57),
    .A_N(\simon1.lfsr_capture[29] ));
 sg13g2_o21ai_1 _1979_ (.B1(_1257_),
    .Y(_1258_),
    .A1(net54),
    .A2(\simon1.lfsr_inst.lfsr_out[28] ));
 sg13g2_nand2_1 _1980_ (.Y(_1259_),
    .A(net36),
    .B(_1258_));
 sg13g2_o21ai_1 _1981_ (.B1(_1259_),
    .Y(_1260_),
    .A1(\simon1.lfsr_inst.lfsr_out[29] ),
    .A2(net37));
 sg13g2_nand2b_1 _1982_ (.Y(_0096_),
    .B(_1260_),
    .A_N(net29));
 sg13g2_nor2_1 _1983_ (.A(_1168_),
    .B(net55),
    .Y(_1261_));
 sg13g2_a21oi_1 _1984_ (.A1(net46),
    .A2(\simon1.lfsr_capture[2] ),
    .Y(_1262_),
    .B1(_1261_));
 sg13g2_nor2_1 _1985_ (.A(_1181_),
    .B(_1262_),
    .Y(_1263_));
 sg13g2_a21oi_1 _1986_ (.A1(\simon1.lfsr_inst.lfsr_out[2] ),
    .A2(_1181_),
    .Y(_1264_),
    .B1(_1263_));
 sg13g2_nor2_1 _1987_ (.A(net30),
    .B(_1264_),
    .Y(_0097_));
 sg13g2_nor2_1 _1988_ (.A(\simon1.lfsr_inst.lfsr_out[30] ),
    .B(net35),
    .Y(_1265_));
 sg13g2_mux2_1 _1989_ (.A0(\simon1.lfsr_inst.lfsr_out[29] ),
    .A1(\simon1.lfsr_capture[30] ),
    .S(net56),
    .X(_1266_));
 sg13g2_nor2_1 _1990_ (.A(_1181_),
    .B(_1266_),
    .Y(_1267_));
 sg13g2_nor3_1 _1991_ (.A(net28),
    .B(_1265_),
    .C(_1267_),
    .Y(_0098_));
 sg13g2_nor2_1 _1992_ (.A(\simon1.lfsr_inst.lfsr_out[31] ),
    .B(net35),
    .Y(_1268_));
 sg13g2_mux2_1 _1993_ (.A0(\simon1.lfsr_inst.lfsr_out[30] ),
    .A1(\simon1.lfsr_capture[31] ),
    .S(net56),
    .X(_1269_));
 sg13g2_nor2_1 _1994_ (.A(_1181_),
    .B(_1269_),
    .Y(_1270_));
 sg13g2_nor3_1 _1995_ (.A(_1161_),
    .B(_1268_),
    .C(_1270_),
    .Y(_0099_));
 sg13g2_nand2b_1 _1996_ (.Y(_1271_),
    .B(net57),
    .A_N(\simon1.lfsr_capture[3] ));
 sg13g2_o21ai_1 _1997_ (.B1(_1271_),
    .Y(_1272_),
    .A1(net54),
    .A2(\simon1.lfsr_inst.lfsr_out[2] ));
 sg13g2_nand2_1 _1998_ (.Y(_1273_),
    .A(net36),
    .B(_1272_));
 sg13g2_o21ai_1 _1999_ (.B1(_1273_),
    .Y(_1274_),
    .A1(\simon1.lfsr_inst.lfsr_out[3] ),
    .A2(net37));
 sg13g2_nand2b_1 _2000_ (.Y(_0100_),
    .B(_1274_),
    .A_N(net29));
 sg13g2_nand2b_1 _2001_ (.Y(_1275_),
    .B(net57),
    .A_N(\simon1.lfsr_capture[4] ));
 sg13g2_o21ai_1 _2002_ (.B1(_1275_),
    .Y(_1276_),
    .A1(net54),
    .A2(\simon1.lfsr_inst.lfsr_out[3] ));
 sg13g2_nand2_1 _2003_ (.Y(_1277_),
    .A(net41),
    .B(_1276_));
 sg13g2_o21ai_1 _2004_ (.B1(_1277_),
    .Y(_1278_),
    .A1(\simon1.lfsr_inst.lfsr_out[4] ),
    .A2(net39));
 sg13g2_nand2b_1 _2005_ (.Y(_0101_),
    .B(_1278_),
    .A_N(net29));
 sg13g2_nand2b_1 _2006_ (.Y(_1279_),
    .B(net57),
    .A_N(\simon1.lfsr_capture[5] ));
 sg13g2_o21ai_1 _2007_ (.B1(_1279_),
    .Y(_1280_),
    .A1(net54),
    .A2(\simon1.lfsr_inst.lfsr_out[4] ));
 sg13g2_nand2_1 _2008_ (.Y(_1281_),
    .A(net41),
    .B(_1280_));
 sg13g2_o21ai_1 _2009_ (.B1(_1281_),
    .Y(_1282_),
    .A1(\simon1.lfsr_inst.lfsr_out[5] ),
    .A2(net39));
 sg13g2_nand2b_1 _2010_ (.Y(_0102_),
    .B(_1282_),
    .A_N(net29));
 sg13g2_nand2b_1 _2011_ (.Y(_1283_),
    .B(net57),
    .A_N(\simon1.lfsr_capture[6] ));
 sg13g2_o21ai_1 _2012_ (.B1(_1283_),
    .Y(_1284_),
    .A1(net55),
    .A2(\simon1.lfsr_inst.lfsr_out[5] ));
 sg13g2_nand2_1 _2013_ (.Y(_1285_),
    .A(net41),
    .B(_1284_));
 sg13g2_o21ai_1 _2014_ (.B1(_1285_),
    .Y(_1286_),
    .A1(\simon1.lfsr_inst.lfsr_out[6] ),
    .A2(net39));
 sg13g2_nand2b_1 _2015_ (.Y(_0103_),
    .B(_1286_),
    .A_N(net29));
 sg13g2_nand2b_1 _2016_ (.Y(_1287_),
    .B(net57),
    .A_N(\simon1.lfsr_capture[7] ));
 sg13g2_o21ai_1 _2017_ (.B1(_1287_),
    .Y(_1288_),
    .A1(net55),
    .A2(\simon1.lfsr_inst.lfsr_out[6] ));
 sg13g2_nand2_1 _2018_ (.Y(_1289_),
    .A(net41),
    .B(_1288_));
 sg13g2_o21ai_1 _2019_ (.B1(_1289_),
    .Y(_1290_),
    .A1(\simon1.lfsr_inst.lfsr_out[7] ),
    .A2(net39));
 sg13g2_nand2b_1 _2020_ (.Y(_0104_),
    .B(_1290_),
    .A_N(net29));
 sg13g2_nor2_1 _2021_ (.A(\simon1.lfsr_inst.lfsr_out[8] ),
    .B(net35),
    .Y(_1291_));
 sg13g2_mux2_1 _2022_ (.A0(\simon1.lfsr_inst.lfsr_out[7] ),
    .A1(\simon1.lfsr_capture[8] ),
    .S(net56),
    .X(_1292_));
 sg13g2_nor2_1 _2023_ (.A(_1181_),
    .B(_1292_),
    .Y(_1293_));
 sg13g2_nor3_1 _2024_ (.A(_1161_),
    .B(_1291_),
    .C(_1293_),
    .Y(_0105_));
 sg13g2_nand2b_1 _2025_ (.Y(_1294_),
    .B(net57),
    .A_N(\simon1.lfsr_capture[9] ));
 sg13g2_o21ai_1 _2026_ (.B1(_1294_),
    .Y(_1295_),
    .A1(net55),
    .A2(\simon1.lfsr_inst.lfsr_out[8] ));
 sg13g2_nand2_1 _2027_ (.Y(_1296_),
    .A(net41),
    .B(_1295_));
 sg13g2_o21ai_1 _2028_ (.B1(_1296_),
    .Y(_1297_),
    .A1(\simon1.lfsr_inst.lfsr_out[9] ),
    .A2(net39));
 sg13g2_nand2b_1 _2029_ (.Y(_0106_),
    .B(_1297_),
    .A_N(net29));
 sg13g2_inv_1 _2030_ (.Y(_1298_),
    .A(_0012_));
 sg13g2_nand2b_1 _2031_ (.Y(_1299_),
    .B(net85),
    .A_N(\simon1.score_rst ));
 sg13g2_buf_1 _2032_ (.A(_1299_),
    .X(_1300_));
 sg13g2_nor2_1 _2033_ (.A(_1298_),
    .B(net53),
    .Y(_0125_));
 sg13g2_xnor2_1 _2034_ (.Y(_1301_),
    .A(\simon1.score_inst.ones[0] ),
    .B(\simon1.score_inc ));
 sg13g2_nor2_1 _2035_ (.A(net53),
    .B(_1301_),
    .Y(_0126_));
 sg13g2_nand2_2 _2036_ (.Y(_1302_),
    .A(\simon1.score_inst.ones[0] ),
    .B(\simon1.score_inc ));
 sg13g2_nor2_1 _2037_ (.A(\simon1.score_inst.ones[2] ),
    .B(_1091_),
    .Y(_1303_));
 sg13g2_nor3_1 _2038_ (.A(_1079_),
    .B(_1302_),
    .C(_1303_),
    .Y(_1304_));
 sg13g2_a21oi_1 _2039_ (.A1(_1079_),
    .A2(_1302_),
    .Y(_1305_),
    .B1(_1304_));
 sg13g2_nor2_1 _2040_ (.A(net53),
    .B(_1305_),
    .Y(_0127_));
 sg13g2_inv_1 _2041_ (.Y(_1306_),
    .A(\simon1.score_inst.ones[2] ));
 sg13g2_nand3_1 _2042_ (.B(_1079_),
    .C(\simon1.score_inc ),
    .A(\simon1.score_inst.ones[0] ),
    .Y(_1307_));
 sg13g2_xnor2_1 _2043_ (.Y(_1308_),
    .A(_1306_),
    .B(_1307_));
 sg13g2_nor2_1 _2044_ (.A(net53),
    .B(_1308_),
    .Y(_0128_));
 sg13g2_nor2_1 _2045_ (.A(_1079_),
    .B(_1306_),
    .Y(_1309_));
 sg13g2_o21ai_1 _2046_ (.B1(\simon1.score_inst.ones[3] ),
    .Y(_1310_),
    .A1(_1302_),
    .A2(_1309_));
 sg13g2_nor3_1 _2047_ (.A(_1306_),
    .B(\simon1.score_inst.ones[3] ),
    .C(_1302_),
    .Y(_1311_));
 sg13g2_o21ai_1 _2048_ (.B1(_1079_),
    .Y(_1312_),
    .A1(_1303_),
    .A2(_1311_));
 sg13g2_a21oi_1 _2049_ (.A1(_1310_),
    .A2(_1312_),
    .Y(_0129_),
    .B1(net53));
 sg13g2_nor4_2 _2050_ (.A(_1079_),
    .B(\simon1.score_inst.ones[2] ),
    .C(_1091_),
    .Y(_1313_),
    .D(_1302_));
 sg13g2_xnor2_1 _2051_ (.Y(_1314_),
    .A(\simon1.score_inst.tens[0] ),
    .B(_1313_));
 sg13g2_nor2_1 _2052_ (.A(_1300_),
    .B(_1314_),
    .Y(_0130_));
 sg13g2_nand2_1 _2053_ (.Y(_1315_),
    .A(\simon1.score_inst.tens[0] ),
    .B(_1313_));
 sg13g2_nor2b_1 _2054_ (.A(\simon1.score_inst.tens[2] ),
    .B_N(\simon1.score_inst.tens[3] ),
    .Y(_1316_));
 sg13g2_nor3_1 _2055_ (.A(_1081_),
    .B(_1315_),
    .C(_1316_),
    .Y(_1317_));
 sg13g2_a21oi_1 _2056_ (.A1(_1081_),
    .A2(_1315_),
    .Y(_1318_),
    .B1(_1317_));
 sg13g2_nor2_1 _2057_ (.A(net53),
    .B(_1318_),
    .Y(_0131_));
 sg13g2_nand3_1 _2058_ (.B(_1081_),
    .C(_1313_),
    .A(\simon1.score_inst.tens[0] ),
    .Y(_1319_));
 sg13g2_xnor2_1 _2059_ (.Y(_1320_),
    .A(_1086_),
    .B(_1319_));
 sg13g2_nor2_1 _2060_ (.A(net53),
    .B(_1320_),
    .Y(_0132_));
 sg13g2_nor2_1 _2061_ (.A(_1081_),
    .B(_1086_),
    .Y(_1321_));
 sg13g2_o21ai_1 _2062_ (.B1(\simon1.score_inst.tens[3] ),
    .Y(_1322_),
    .A1(_1315_),
    .A2(_1321_));
 sg13g2_nor3_1 _2063_ (.A(_1086_),
    .B(\simon1.score_inst.tens[3] ),
    .C(_1315_),
    .Y(_1323_));
 sg13g2_o21ai_1 _2064_ (.B1(_1081_),
    .Y(_1324_),
    .A1(_1316_),
    .A2(_1323_));
 sg13g2_a21oi_1 _2065_ (.A1(_1322_),
    .A2(_1324_),
    .Y(_0133_),
    .B1(net53));
 sg13g2_buf_1 _2066_ (.A(\simon1.sound_freq[5] ),
    .X(_1325_));
 sg13g2_buf_2 _2067_ (.A(\simon1.sound_freq[4] ),
    .X(_1326_));
 sg13g2_nor2_1 _2068_ (.A(net75),
    .B(_1326_),
    .Y(_1327_));
 sg13g2_buf_2 _2069_ (.A(\simon1.sound_freq[9] ),
    .X(_1328_));
 sg13g2_buf_1 _2070_ (.A(\simon1.sound_freq[8] ),
    .X(_1329_));
 sg13g2_nor2_1 _2071_ (.A(_1328_),
    .B(net74),
    .Y(_1330_));
 sg13g2_buf_2 _2072_ (.A(\simon1.sound_freq[7] ),
    .X(_1331_));
 sg13g2_buf_1 _2073_ (.A(\simon1.sound_freq[6] ),
    .X(_1332_));
 sg13g2_nor2_1 _2074_ (.A(_1331_),
    .B(net73),
    .Y(_1333_));
 sg13g2_buf_2 _2075_ (.A(\simon1.sound_freq[2] ),
    .X(_1334_));
 sg13g2_nor4_1 _2076_ (.A(\simon1.sound_freq[0] ),
    .B(\simon1.sound_freq[1] ),
    .C(\simon1.sound_freq[3] ),
    .D(_1334_),
    .Y(_1335_));
 sg13g2_nand4_1 _2077_ (.B(_1330_),
    .C(_1333_),
    .A(_1327_),
    .Y(_1336_),
    .D(_1335_));
 sg13g2_buf_2 _2078_ (.A(_1336_),
    .X(_1337_));
 sg13g2_buf_1 _2079_ (.A(_1337_),
    .X(_1338_));
 sg13g2_nand2_2 _2080_ (.Y(_1339_),
    .A(net85),
    .B(net34));
 sg13g2_buf_1 _2081_ (.A(\simon1.sound_gen_inst.tick_counter[13] ),
    .X(_1340_));
 sg13g2_nand2_1 _2082_ (.Y(_1341_),
    .A(\simon1.sound_gen_inst.tick_counter[14] ),
    .B(net72));
 sg13g2_buf_1 _2083_ (.A(\simon1.sound_gen_inst.tick_counter[7] ),
    .X(_1342_));
 sg13g2_buf_1 _2084_ (.A(\simon1.sound_gen_inst.tick_counter[8] ),
    .X(_1343_));
 sg13g2_nand2_1 _2085_ (.Y(_1344_),
    .A(net71),
    .B(net70));
 sg13g2_nor2_1 _2086_ (.A(_1341_),
    .B(_1344_),
    .Y(_1345_));
 sg13g2_buf_8 _2087_ (.A(\simon1.sound_gen_inst.tick_counter[3] ),
    .X(_1346_));
 sg13g2_inv_1 _2088_ (.Y(_1347_),
    .A(_1346_));
 sg13g2_buf_2 _2089_ (.A(\simon1.sound_gen_inst.tick_counter[2] ),
    .X(_1348_));
 sg13g2_buf_2 _2090_ (.A(\simon1.sound_gen_inst.tick_counter[15] ),
    .X(_1349_));
 sg13g2_nor4_1 _2091_ (.A(\simon1.sound_gen_inst.tick_counter[0] ),
    .B(_1347_),
    .C(_1348_),
    .D(_1349_),
    .Y(_1350_));
 sg13g2_buf_1 _2092_ (.A(\simon1.sound_gen_inst.tick_counter[12] ),
    .X(_1351_));
 sg13g2_buf_1 _2093_ (.A(\simon1.sound_gen_inst.tick_counter[11] ),
    .X(_1352_));
 sg13g2_buf_1 _2094_ (.A(\simon1.sound_gen_inst.tick_counter[10] ),
    .X(_1353_));
 sg13g2_buf_1 _2095_ (.A(\simon1.sound_gen_inst.tick_counter[9] ),
    .X(_1354_));
 sg13g2_nor4_1 _2096_ (.A(_1351_),
    .B(net69),
    .C(_1353_),
    .D(net68),
    .Y(_1355_));
 sg13g2_buf_1 _2097_ (.A(\simon1.sound_gen_inst.tick_counter[6] ),
    .X(_1356_));
 sg13g2_buf_1 _2098_ (.A(\simon1.sound_gen_inst.tick_counter[4] ),
    .X(_1357_));
 sg13g2_buf_1 _2099_ (.A(\simon1.sound_gen_inst.tick_counter[5] ),
    .X(_1358_));
 sg13g2_inv_1 _2100_ (.Y(_1359_),
    .A(net65));
 sg13g2_nor4_1 _2101_ (.A(\simon1.sound_gen_inst.tick_counter[1] ),
    .B(net67),
    .C(net66),
    .D(_1359_),
    .Y(_1360_));
 sg13g2_and4_1 _2102_ (.A(_1345_),
    .B(_1350_),
    .C(_1355_),
    .D(_1360_),
    .X(_1361_));
 sg13g2_buf_1 _2103_ (.A(\simon1.sound_gen_inst.tick_counter[23] ),
    .X(_1362_));
 sg13g2_inv_1 _2104_ (.Y(_1363_),
    .A(_1362_));
 sg13g2_buf_1 _2105_ (.A(\simon1.sound_gen_inst.tick_counter[27] ),
    .X(_1364_));
 sg13g2_nor4_1 _2106_ (.A(\simon1.sound_gen_inst.tick_counter[31] ),
    .B(\simon1.sound_gen_inst.tick_counter[29] ),
    .C(\simon1.sound_gen_inst.tick_counter[28] ),
    .D(_1364_),
    .Y(_1365_));
 sg13g2_nand3b_1 _2107_ (.B(_1363_),
    .C(_1365_),
    .Y(_1366_),
    .A_N(\simon1.sound_gen_inst.tick_counter[30] ));
 sg13g2_buf_1 _2108_ (.A(\simon1.sound_gen_inst.tick_counter[18] ),
    .X(_1367_));
 sg13g2_buf_1 _2109_ (.A(\simon1.sound_gen_inst.tick_counter[16] ),
    .X(_1368_));
 sg13g2_nor3_1 _2110_ (.A(net64),
    .B(\simon1.sound_gen_inst.tick_counter[17] ),
    .C(_1368_),
    .Y(_1369_));
 sg13g2_buf_2 _2111_ (.A(\simon1.sound_gen_inst.tick_counter[24] ),
    .X(_1370_));
 sg13g2_nor4_1 _2112_ (.A(_1349_),
    .B(\simon1.sound_gen_inst.tick_counter[26] ),
    .C(\simon1.sound_gen_inst.tick_counter[25] ),
    .D(_1370_),
    .Y(_1371_));
 sg13g2_buf_1 _2113_ (.A(\simon1.sound_gen_inst.tick_counter[22] ),
    .X(_1372_));
 sg13g2_buf_2 _2114_ (.A(\simon1.sound_gen_inst.tick_counter[21] ),
    .X(_1373_));
 sg13g2_buf_1 _2115_ (.A(\simon1.sound_gen_inst.tick_counter[20] ),
    .X(_1374_));
 sg13g2_buf_1 _2116_ (.A(\simon1.sound_gen_inst.tick_counter[19] ),
    .X(_1375_));
 sg13g2_nor4_1 _2117_ (.A(_1372_),
    .B(_1373_),
    .C(_1374_),
    .D(_1375_),
    .Y(_1376_));
 sg13g2_nand3_1 _2118_ (.B(_1371_),
    .C(_1376_),
    .A(_1369_),
    .Y(_1377_));
 sg13g2_inv_1 _2119_ (.Y(_1378_),
    .A(net67));
 sg13g2_o21ai_1 _2120_ (.B1(net65),
    .Y(_1379_),
    .A1(_1346_),
    .A2(net66));
 sg13g2_a21o_1 _2121_ (.A2(_1379_),
    .A1(_1378_),
    .B1(_1344_),
    .X(_1380_));
 sg13g2_a21oi_1 _2122_ (.A1(_1355_),
    .A2(_1380_),
    .Y(_1381_),
    .B1(_1341_));
 sg13g2_or4_1 _2123_ (.A(_1361_),
    .B(_1366_),
    .C(_1377_),
    .D(_1381_),
    .X(_1382_));
 sg13g2_buf_1 _2124_ (.A(_1382_),
    .X(_1383_));
 sg13g2_mux2_1 _2125_ (.A0(\simon1.sound ),
    .A1(_0013_),
    .S(net27),
    .X(_1384_));
 sg13g2_nor2b_1 _2126_ (.A(_1339_),
    .B_N(_1384_),
    .Y(_0159_));
 sg13g2_inv_1 _2127_ (.Y(_1385_),
    .A(_0035_));
 sg13g2_inv_1 _2128_ (.Y(_1386_),
    .A(\simon1.tick_counter[0] ));
 sg13g2_nor4_1 _2129_ (.A(_1386_),
    .B(\simon1.tick_counter[8] ),
    .C(\simon1.tick_counter[10] ),
    .D(\simon1.tick_counter[11] ),
    .Y(_1387_));
 sg13g2_nor4_1 _2130_ (.A(\simon1.tick_counter[12] ),
    .B(\simon1.tick_counter[13] ),
    .C(\simon1.tick_counter[14] ),
    .D(\simon1.tick_counter[15] ),
    .Y(_1388_));
 sg13g2_nor4_1 _2131_ (.A(\simon1.tick_counter[2] ),
    .B(\simon1.tick_counter[3] ),
    .C(\simon1.tick_counter[6] ),
    .D(\simon1.tick_counter[7] ),
    .Y(_1389_));
 sg13g2_nand2_1 _2132_ (.Y(_1390_),
    .A(\simon1.tick_counter[4] ),
    .B(\simon1.tick_counter[5] ));
 sg13g2_nor3_1 _2133_ (.A(\simon1.tick_counter[1] ),
    .B(\simon1.tick_counter[9] ),
    .C(_1390_),
    .Y(_1391_));
 sg13g2_and4_1 _2134_ (.A(_1387_),
    .B(_1388_),
    .C(_1389_),
    .D(_1391_),
    .X(_1392_));
 sg13g2_buf_1 _2135_ (.A(_1392_),
    .X(_1393_));
 sg13g2_nand2b_1 _2136_ (.Y(_1394_),
    .B(net85),
    .A_N(_1393_));
 sg13g2_buf_1 _2137_ (.A(_1394_),
    .X(_1395_));
 sg13g2_buf_1 _2138_ (.A(_1395_),
    .X(_1396_));
 sg13g2_nor2_1 _2139_ (.A(_1385_),
    .B(net25),
    .Y(_0192_));
 sg13g2_inv_1 _2140_ (.Y(_1397_),
    .A(\simon1.tick_counter[8] ));
 sg13g2_nand4_1 _2141_ (.B(\simon1.tick_counter[1] ),
    .C(\simon1.tick_counter[2] ),
    .A(\simon1.tick_counter[0] ),
    .Y(_1398_),
    .D(\simon1.tick_counter[3] ));
 sg13g2_nor2_1 _2142_ (.A(_1390_),
    .B(_1398_),
    .Y(_1399_));
 sg13g2_nand3_1 _2143_ (.B(\simon1.tick_counter[7] ),
    .C(_1399_),
    .A(\simon1.tick_counter[6] ),
    .Y(_1400_));
 sg13g2_nor2_1 _2144_ (.A(_1397_),
    .B(_1400_),
    .Y(_1401_));
 sg13g2_nand2_1 _2145_ (.Y(_1402_),
    .A(\simon1.tick_counter[9] ),
    .B(_1401_));
 sg13g2_xor2_1 _2146_ (.B(_1402_),
    .A(\simon1.tick_counter[10] ),
    .X(_1403_));
 sg13g2_nor2_1 _2147_ (.A(net25),
    .B(_1403_),
    .Y(_0193_));
 sg13g2_inv_1 _2148_ (.Y(_1404_),
    .A(\simon1.tick_counter[11] ));
 sg13g2_nand3_1 _2149_ (.B(\simon1.tick_counter[10] ),
    .C(_1401_),
    .A(\simon1.tick_counter[9] ),
    .Y(_1405_));
 sg13g2_xnor2_1 _2150_ (.Y(_1406_),
    .A(_1404_),
    .B(_1405_));
 sg13g2_nor2_1 _2151_ (.A(net25),
    .B(_1406_),
    .Y(_0194_));
 sg13g2_nor2_2 _2152_ (.A(_1404_),
    .B(_1405_),
    .Y(_1407_));
 sg13g2_xnor2_1 _2153_ (.Y(_1408_),
    .A(\simon1.tick_counter[12] ),
    .B(_1407_));
 sg13g2_nor2_1 _2154_ (.A(net25),
    .B(_1408_),
    .Y(_0195_));
 sg13g2_nand2_1 _2155_ (.Y(_1409_),
    .A(\simon1.tick_counter[12] ),
    .B(_1407_));
 sg13g2_xor2_1 _2156_ (.B(_1409_),
    .A(\simon1.tick_counter[13] ),
    .X(_1410_));
 sg13g2_nor2_1 _2157_ (.A(net25),
    .B(_1410_),
    .Y(_0196_));
 sg13g2_nand3_1 _2158_ (.B(\simon1.tick_counter[13] ),
    .C(_1407_),
    .A(\simon1.tick_counter[12] ),
    .Y(_1411_));
 sg13g2_xor2_1 _2159_ (.B(_1411_),
    .A(\simon1.tick_counter[14] ),
    .X(_1412_));
 sg13g2_nor2_1 _2160_ (.A(_1396_),
    .B(_1412_),
    .Y(_0197_));
 sg13g2_nand4_1 _2161_ (.B(\simon1.tick_counter[13] ),
    .C(\simon1.tick_counter[14] ),
    .A(\simon1.tick_counter[12] ),
    .Y(_1413_),
    .D(_1407_));
 sg13g2_xor2_1 _2162_ (.B(_1413_),
    .A(\simon1.tick_counter[15] ),
    .X(_1414_));
 sg13g2_nor2_1 _2163_ (.A(_1396_),
    .B(_1414_),
    .Y(_0198_));
 sg13g2_xnor2_1 _2164_ (.Y(_1415_),
    .A(\simon1.tick_counter[0] ),
    .B(\simon1.tick_counter[1] ));
 sg13g2_nor2_1 _2165_ (.A(net25),
    .B(_1415_),
    .Y(_0199_));
 sg13g2_nand2_1 _2166_ (.Y(_1416_),
    .A(\simon1.tick_counter[0] ),
    .B(\simon1.tick_counter[1] ));
 sg13g2_xor2_1 _2167_ (.B(_1416_),
    .A(\simon1.tick_counter[2] ),
    .X(_1417_));
 sg13g2_nor2_1 _2168_ (.A(net25),
    .B(_1417_),
    .Y(_0200_));
 sg13g2_nand3_1 _2169_ (.B(\simon1.tick_counter[1] ),
    .C(\simon1.tick_counter[2] ),
    .A(\simon1.tick_counter[0] ),
    .Y(_1418_));
 sg13g2_xor2_1 _2170_ (.B(_1418_),
    .A(\simon1.tick_counter[3] ),
    .X(_1419_));
 sg13g2_nor2_1 _2171_ (.A(net25),
    .B(_1419_),
    .Y(_0201_));
 sg13g2_inv_1 _2172_ (.Y(_1420_),
    .A(\simon1.tick_counter[4] ));
 sg13g2_xnor2_1 _2173_ (.Y(_1421_),
    .A(_1420_),
    .B(_1398_));
 sg13g2_nor2_1 _2174_ (.A(_1395_),
    .B(_1421_),
    .Y(_0202_));
 sg13g2_nor2_1 _2175_ (.A(_1420_),
    .B(_1398_),
    .Y(_1422_));
 sg13g2_xnor2_1 _2176_ (.Y(_1423_),
    .A(\simon1.tick_counter[5] ),
    .B(_1422_));
 sg13g2_nor2_1 _2177_ (.A(_1395_),
    .B(_1423_),
    .Y(_0203_));
 sg13g2_xnor2_1 _2178_ (.Y(_1424_),
    .A(\simon1.tick_counter[6] ),
    .B(_1399_));
 sg13g2_nor2_1 _2179_ (.A(_1395_),
    .B(_1424_),
    .Y(_0204_));
 sg13g2_nand2_1 _2180_ (.Y(_1425_),
    .A(\simon1.tick_counter[6] ),
    .B(_1399_));
 sg13g2_xor2_1 _2181_ (.B(_1425_),
    .A(\simon1.tick_counter[7] ),
    .X(_1426_));
 sg13g2_nor2_1 _2182_ (.A(_1395_),
    .B(_1426_),
    .Y(_0205_));
 sg13g2_xnor2_1 _2183_ (.Y(_1427_),
    .A(_1397_),
    .B(_1400_));
 sg13g2_nor2_1 _2184_ (.A(_1395_),
    .B(_1427_),
    .Y(_0206_));
 sg13g2_xnor2_1 _2185_ (.Y(_1428_),
    .A(\simon1.tick_counter[9] ),
    .B(_1401_));
 sg13g2_nor2_1 _2186_ (.A(_1395_),
    .B(_1428_),
    .Y(_0207_));
 sg13g2_inv_1 _2187_ (.Y(_1429_),
    .A(_0946_));
 sg13g2_nand2_1 _2188_ (.Y(_1430_),
    .A(net80),
    .B(_0957_));
 sg13g2_a21oi_1 _2189_ (.A1(_1029_),
    .A2(_1430_),
    .Y(_1431_),
    .B1(_1048_));
 sg13g2_nand2b_1 _2190_ (.Y(_1432_),
    .B(_1041_),
    .A_N(_1431_));
 sg13g2_buf_1 _2191_ (.A(_0009_),
    .X(_1433_));
 sg13g2_a21oi_1 _2192_ (.A1(_1038_),
    .A2(_1432_),
    .Y(_1434_),
    .B1(_1433_));
 sg13g2_o21ai_1 _2193_ (.B1(\simon1.button_released ),
    .Y(_1435_),
    .A1(_1063_),
    .A2(_1434_));
 sg13g2_a21oi_1 _2194_ (.A1(net78),
    .A2(_0943_),
    .Y(_1436_),
    .B1(_1434_));
 sg13g2_buf_1 _2195_ (.A(net85),
    .X(_1437_));
 sg13g2_o21ai_1 _2196_ (.B1(_1437_),
    .Y(_1438_),
    .A1(\simon1.button_released ),
    .A2(_1436_));
 sg13g2_a21oi_1 _2197_ (.A1(net52),
    .A2(_1435_),
    .Y(_0036_),
    .B1(_1438_));
 sg13g2_inv_1 _2198_ (.Y(_1439_),
    .A(\simon1.state[2] ));
 sg13g2_nor3_1 _2199_ (.A(_0946_),
    .B(_1028_),
    .C(_1026_),
    .Y(_0220_));
 sg13g2_nand3_1 _2200_ (.B(_1137_),
    .C(_0220_),
    .A(_1439_),
    .Y(_0221_));
 sg13g2_nor2_1 _2201_ (.A(_0974_),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_nor2_1 _2202_ (.A(_0025_),
    .B(_0966_),
    .Y(_0223_));
 sg13g2_nor2_2 _2203_ (.A(_0222_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_nor2_1 _2204_ (.A(_1055_),
    .B(_0221_),
    .Y(_0225_));
 sg13g2_o21ai_1 _2205_ (.B1(net59),
    .Y(_0226_),
    .A1(net81),
    .A2(net83));
 sg13g2_nor2_1 _2206_ (.A(net82),
    .B(_0947_),
    .Y(_0227_));
 sg13g2_a21o_1 _2207_ (.A2(_0227_),
    .A1(_1026_),
    .B1(net59),
    .X(_0228_));
 sg13g2_nor2_1 _2208_ (.A(_0021_),
    .B(_0945_),
    .Y(_0229_));
 sg13g2_a221oi_1 _2209_ (.B2(_0228_),
    .C1(_0229_),
    .B1(_0226_),
    .A1(_1017_),
    .Y(_0230_),
    .A2(_0225_));
 sg13g2_buf_1 _2210_ (.A(net85),
    .X(_0231_));
 sg13g2_o21ai_1 _2211_ (.B1(net62),
    .Y(_0232_),
    .A1(net9),
    .A2(_0224_));
 sg13g2_a21oi_1 _2212_ (.A1(_0224_),
    .A2(_0230_),
    .Y(_0037_),
    .B1(_0232_));
 sg13g2_nor2b_1 _2213_ (.A(net83),
    .B_N(net81),
    .Y(_0233_));
 sg13g2_nand2_1 _2214_ (.Y(_0234_),
    .A(_1026_),
    .B(net82));
 sg13g2_nor3_1 _2215_ (.A(net59),
    .B(_0947_),
    .C(_0234_),
    .Y(_0235_));
 sg13g2_a221oi_1 _2216_ (.B2(net59),
    .C1(_0235_),
    .B1(_0233_),
    .A1(_0959_),
    .Y(_0236_),
    .A2(_0225_));
 sg13g2_nor2b_1 _2217_ (.A(_0229_),
    .B_N(_0236_),
    .Y(_0237_));
 sg13g2_o21ai_1 _2218_ (.B1(net62),
    .Y(_0238_),
    .A1(net10),
    .A2(_0224_));
 sg13g2_a21oi_1 _2219_ (.A1(_0224_),
    .A2(_0237_),
    .Y(_0038_),
    .B1(_0238_));
 sg13g2_nor2b_1 _2220_ (.A(net81),
    .B_N(net83),
    .Y(_0239_));
 sg13g2_nand2b_1 _2221_ (.Y(_0240_),
    .B(\simon1.millis_counter[9] ),
    .A_N(_0958_));
 sg13g2_nand2_1 _2222_ (.Y(_0241_),
    .A(net52),
    .B(_1026_));
 sg13g2_nor2_1 _2223_ (.A(net82),
    .B(_1168_),
    .Y(_0242_));
 sg13g2_nor2b_1 _2224_ (.A(_0241_),
    .B_N(_0242_),
    .Y(_0243_));
 sg13g2_a221oi_1 _2225_ (.B2(_0225_),
    .C1(_0243_),
    .B1(_0240_),
    .A1(net59),
    .Y(_0244_),
    .A2(_0239_));
 sg13g2_nor2b_1 _2226_ (.A(_0229_),
    .B_N(_0244_),
    .Y(_0245_));
 sg13g2_o21ai_1 _2227_ (.B1(net62),
    .Y(_0246_),
    .A1(net11),
    .A2(_0224_));
 sg13g2_a21oi_1 _2228_ (.A1(_0224_),
    .A2(_0245_),
    .Y(_0039_),
    .B1(_0246_));
 sg13g2_nand2_1 _2229_ (.Y(_0247_),
    .A(\simon1.millis_counter[9] ),
    .B(_0958_));
 sg13g2_nand2_1 _2230_ (.Y(_0248_),
    .A(net81),
    .B(net83));
 sg13g2_nand2_1 _2231_ (.Y(_0249_),
    .A(_1010_),
    .B(_0248_));
 sg13g2_o21ai_1 _2232_ (.B1(net52),
    .Y(_0250_),
    .A1(_1168_),
    .A2(_0234_));
 sg13g2_a221oi_1 _2233_ (.B2(_0250_),
    .C1(_0229_),
    .B1(_0249_),
    .A1(_0247_),
    .Y(_0251_),
    .A2(_0225_));
 sg13g2_o21ai_1 _2234_ (.B1(net62),
    .Y(_0252_),
    .A1(net12),
    .A2(_0224_));
 sg13g2_a21oi_1 _2235_ (.A1(_0224_),
    .A2(_0251_),
    .Y(_0040_),
    .B1(_0252_));
 sg13g2_inv_1 _2236_ (.Y(_0253_),
    .A(net82));
 sg13g2_nand2_1 _2237_ (.Y(_0254_),
    .A(_1051_),
    .B(_1066_));
 sg13g2_buf_2 _2238_ (.A(_0254_),
    .X(_0255_));
 sg13g2_buf_1 _2239_ (.A(_0255_),
    .X(_0256_));
 sg13g2_nand2_1 _2240_ (.Y(_0257_),
    .A(\simon1.lfsr_capture[0] ),
    .B(net24));
 sg13g2_o21ai_1 _2241_ (.B1(_0257_),
    .Y(_0258_),
    .A1(_0253_),
    .A2(net24));
 sg13g2_and2_1 _2242_ (.A(net60),
    .B(_0258_),
    .X(_0041_));
 sg13g2_mux2_1 _2243_ (.A0(\simon1.lfsr_inst.lfsr_out[10] ),
    .A1(\simon1.lfsr_capture[10] ),
    .S(net24),
    .X(_0259_));
 sg13g2_and2_1 _2244_ (.A(net60),
    .B(_0259_),
    .X(_0042_));
 sg13g2_mux2_1 _2245_ (.A0(\simon1.lfsr_inst.lfsr_out[11] ),
    .A1(\simon1.lfsr_capture[11] ),
    .S(net24),
    .X(_0260_));
 sg13g2_and2_1 _2246_ (.A(net60),
    .B(_0260_),
    .X(_0043_));
 sg13g2_mux2_1 _2247_ (.A0(\simon1.lfsr_inst.lfsr_out[12] ),
    .A1(\simon1.lfsr_capture[12] ),
    .S(net24),
    .X(_0261_));
 sg13g2_and2_1 _2248_ (.A(net60),
    .B(_0261_),
    .X(_0044_));
 sg13g2_mux2_1 _2249_ (.A0(\simon1.lfsr_inst.lfsr_out[13] ),
    .A1(\simon1.lfsr_capture[13] ),
    .S(net24),
    .X(_0262_));
 sg13g2_and2_1 _2250_ (.A(net60),
    .B(_0262_),
    .X(_0045_));
 sg13g2_mux2_1 _2251_ (.A0(\simon1.lfsr_inst.lfsr_out[14] ),
    .A1(\simon1.lfsr_capture[14] ),
    .S(_0256_),
    .X(_0263_));
 sg13g2_and2_1 _2252_ (.A(_0973_),
    .B(_0263_),
    .X(_0046_));
 sg13g2_mux2_1 _2253_ (.A0(\simon1.lfsr_inst.lfsr_out[15] ),
    .A1(\simon1.lfsr_capture[15] ),
    .S(_0256_),
    .X(_0264_));
 sg13g2_and2_1 _2254_ (.A(_0973_),
    .B(_0264_),
    .X(_0047_));
 sg13g2_buf_1 _2255_ (.A(net79),
    .X(_0265_));
 sg13g2_buf_1 _2256_ (.A(_0255_),
    .X(_0266_));
 sg13g2_mux2_1 _2257_ (.A0(\simon1.lfsr_inst.lfsr_out[16] ),
    .A1(\simon1.lfsr_capture[16] ),
    .S(net23),
    .X(_0267_));
 sg13g2_and2_1 _2258_ (.A(_0265_),
    .B(_0267_),
    .X(_0048_));
 sg13g2_mux2_1 _2259_ (.A0(\simon1.lfsr_inst.lfsr_out[17] ),
    .A1(\simon1.lfsr_capture[17] ),
    .S(net23),
    .X(_0268_));
 sg13g2_and2_1 _2260_ (.A(net51),
    .B(_0268_),
    .X(_0049_));
 sg13g2_mux2_1 _2261_ (.A0(\simon1.lfsr_inst.lfsr_out[18] ),
    .A1(\simon1.lfsr_capture[18] ),
    .S(net23),
    .X(_0269_));
 sg13g2_and2_1 _2262_ (.A(net51),
    .B(_0269_),
    .X(_0050_));
 sg13g2_mux2_1 _2263_ (.A0(\simon1.lfsr_inst.lfsr_out[19] ),
    .A1(\simon1.lfsr_capture[19] ),
    .S(net23),
    .X(_0270_));
 sg13g2_and2_1 _2264_ (.A(_0265_),
    .B(_0270_),
    .X(_0051_));
 sg13g2_nand2_1 _2265_ (.Y(_0271_),
    .A(\simon1.lfsr_capture[1] ),
    .B(net24));
 sg13g2_o21ai_1 _2266_ (.B1(_0271_),
    .Y(_0272_),
    .A1(_1168_),
    .A2(net24));
 sg13g2_and2_1 _2267_ (.A(net51),
    .B(_0272_),
    .X(_0052_));
 sg13g2_mux2_1 _2268_ (.A0(\simon1.lfsr_inst.lfsr_out[20] ),
    .A1(\simon1.lfsr_capture[20] ),
    .S(_0266_),
    .X(_0273_));
 sg13g2_and2_1 _2269_ (.A(net51),
    .B(_0273_),
    .X(_0053_));
 sg13g2_mux2_1 _2270_ (.A0(\simon1.lfsr_inst.lfsr_out[21] ),
    .A1(\simon1.lfsr_capture[21] ),
    .S(_0266_),
    .X(_0274_));
 sg13g2_and2_1 _2271_ (.A(net51),
    .B(_0274_),
    .X(_0054_));
 sg13g2_mux2_1 _2272_ (.A0(\simon1.lfsr_inst.lfsr_out[22] ),
    .A1(\simon1.lfsr_capture[22] ),
    .S(net23),
    .X(_0275_));
 sg13g2_and2_1 _2273_ (.A(net51),
    .B(_0275_),
    .X(_0055_));
 sg13g2_mux2_1 _2274_ (.A0(\simon1.lfsr_inst.lfsr_out[23] ),
    .A1(\simon1.lfsr_capture[23] ),
    .S(net23),
    .X(_0276_));
 sg13g2_and2_1 _2275_ (.A(net51),
    .B(_0276_),
    .X(_0056_));
 sg13g2_mux2_1 _2276_ (.A0(\simon1.lfsr_inst.lfsr_out[24] ),
    .A1(\simon1.lfsr_capture[24] ),
    .S(net23),
    .X(_0277_));
 sg13g2_and2_1 _2277_ (.A(net51),
    .B(_0277_),
    .X(_0057_));
 sg13g2_buf_1 _2278_ (.A(_0972_),
    .X(_0278_));
 sg13g2_mux2_1 _2279_ (.A0(\simon1.lfsr_inst.lfsr_out[25] ),
    .A1(\simon1.lfsr_capture[25] ),
    .S(net23),
    .X(_0279_));
 sg13g2_and2_1 _2280_ (.A(_0278_),
    .B(_0279_),
    .X(_0058_));
 sg13g2_buf_1 _2281_ (.A(_0255_),
    .X(_0280_));
 sg13g2_mux2_1 _2282_ (.A0(\simon1.lfsr_inst.lfsr_out[26] ),
    .A1(\simon1.lfsr_capture[26] ),
    .S(_0280_),
    .X(_0281_));
 sg13g2_and2_1 _2283_ (.A(net50),
    .B(_0281_),
    .X(_0059_));
 sg13g2_mux2_1 _2284_ (.A0(\simon1.lfsr_inst.lfsr_out[27] ),
    .A1(\simon1.lfsr_capture[27] ),
    .S(net22),
    .X(_0282_));
 sg13g2_and2_1 _2285_ (.A(net50),
    .B(_0282_),
    .X(_0060_));
 sg13g2_mux2_1 _2286_ (.A0(\simon1.lfsr_inst.lfsr_out[28] ),
    .A1(\simon1.lfsr_capture[28] ),
    .S(net22),
    .X(_0283_));
 sg13g2_and2_1 _2287_ (.A(net50),
    .B(_0283_),
    .X(_0061_));
 sg13g2_mux2_1 _2288_ (.A0(\simon1.lfsr_inst.lfsr_out[29] ),
    .A1(\simon1.lfsr_capture[29] ),
    .S(net22),
    .X(_0284_));
 sg13g2_and2_1 _2289_ (.A(net50),
    .B(_0284_),
    .X(_0062_));
 sg13g2_mux2_1 _2290_ (.A0(\simon1.lfsr_inst.lfsr_out[2] ),
    .A1(\simon1.lfsr_capture[2] ),
    .S(_0280_),
    .X(_0285_));
 sg13g2_and2_1 _2291_ (.A(_0278_),
    .B(_0285_),
    .X(_0063_));
 sg13g2_mux2_1 _2292_ (.A0(\simon1.lfsr_inst.lfsr_out[30] ),
    .A1(\simon1.lfsr_capture[30] ),
    .S(net22),
    .X(_0286_));
 sg13g2_and2_1 _2293_ (.A(net50),
    .B(_0286_),
    .X(_0064_));
 sg13g2_mux2_1 _2294_ (.A0(\simon1.lfsr_inst.lfsr_out[31] ),
    .A1(\simon1.lfsr_capture[31] ),
    .S(net22),
    .X(_0287_));
 sg13g2_and2_1 _2295_ (.A(net50),
    .B(_0287_),
    .X(_0065_));
 sg13g2_mux2_1 _2296_ (.A0(\simon1.lfsr_inst.lfsr_out[3] ),
    .A1(\simon1.lfsr_capture[3] ),
    .S(net22),
    .X(_0288_));
 sg13g2_and2_1 _2297_ (.A(net50),
    .B(_0288_),
    .X(_0066_));
 sg13g2_mux2_1 _2298_ (.A0(\simon1.lfsr_inst.lfsr_out[4] ),
    .A1(\simon1.lfsr_capture[4] ),
    .S(net22),
    .X(_0289_));
 sg13g2_and2_1 _2299_ (.A(net50),
    .B(_0289_),
    .X(_0067_));
 sg13g2_mux2_1 _2300_ (.A0(\simon1.lfsr_inst.lfsr_out[5] ),
    .A1(\simon1.lfsr_capture[5] ),
    .S(net22),
    .X(_0290_));
 sg13g2_and2_1 _2301_ (.A(net63),
    .B(_0290_),
    .X(_0068_));
 sg13g2_mux2_1 _2302_ (.A0(\simon1.lfsr_inst.lfsr_out[6] ),
    .A1(\simon1.lfsr_capture[6] ),
    .S(_0255_),
    .X(_0291_));
 sg13g2_and2_1 _2303_ (.A(net63),
    .B(_0291_),
    .X(_0069_));
 sg13g2_mux2_1 _2304_ (.A0(\simon1.lfsr_inst.lfsr_out[7] ),
    .A1(\simon1.lfsr_capture[7] ),
    .S(_0255_),
    .X(_0292_));
 sg13g2_and2_1 _2305_ (.A(net63),
    .B(_0292_),
    .X(_0070_));
 sg13g2_mux2_1 _2306_ (.A0(\simon1.lfsr_inst.lfsr_out[8] ),
    .A1(\simon1.lfsr_capture[8] ),
    .S(_0255_),
    .X(_0293_));
 sg13g2_and2_1 _2307_ (.A(net63),
    .B(_0293_),
    .X(_0071_));
 sg13g2_mux2_1 _2308_ (.A0(\simon1.lfsr_inst.lfsr_out[9] ),
    .A1(\simon1.lfsr_capture[9] ),
    .S(_0255_),
    .X(_0294_));
 sg13g2_and2_1 _2309_ (.A(net63),
    .B(_0294_),
    .X(_0072_));
 sg13g2_nand3_1 _2310_ (.B(_0972_),
    .C(_0241_),
    .A(\simon1.lfsr_cycles[1] ),
    .Y(_0295_));
 sg13g2_nor3_1 _2311_ (.A(\simon1.lfsr_cycles[0] ),
    .B(_1044_),
    .C(_0295_),
    .Y(_0073_));
 sg13g2_a21oi_1 _2312_ (.A1(\simon1.lfsr_cycles[0] ),
    .A2(\simon1.lfsr_cycles[1] ),
    .Y(_0296_),
    .B1(_1026_));
 sg13g2_a21oi_1 _2313_ (.A1(_1072_),
    .A2(_0296_),
    .Y(_0074_),
    .B1(net48));
 sg13g2_a21oi_1 _2314_ (.A1(_1013_),
    .A2(_1069_),
    .Y(_0107_),
    .B1(_1009_));
 sg13g2_nor2_1 _2315_ (.A(_0944_),
    .B(_0974_),
    .Y(_0297_));
 sg13g2_nand2_1 _2316_ (.Y(_0298_),
    .A(_0945_),
    .B(_1064_));
 sg13g2_a221oi_1 _2317_ (.B2(_1429_),
    .C1(_0298_),
    .B1(_0297_),
    .A1(_0974_),
    .Y(_0299_),
    .A2(_0943_));
 sg13g2_nand2b_1 _2318_ (.Y(_0300_),
    .B(_0299_),
    .A_N(_1012_));
 sg13g2_a22oi_1 _2319_ (.Y(_0301_),
    .B1(_0300_),
    .B2(\simon1.lfsr_stopped ),
    .A2(_0299_),
    .A1(_1433_));
 sg13g2_nor2_1 _2320_ (.A(net47),
    .B(_0301_),
    .Y(_0108_));
 sg13g2_inv_1 _2321_ (.Y(_0302_),
    .A(_0953_));
 sg13g2_a21oi_1 _2322_ (.A1(_0946_),
    .A2(_0302_),
    .Y(_0303_),
    .B1(_1028_));
 sg13g2_nand2_1 _2323_ (.Y(_0304_),
    .A(_0966_),
    .B(_1124_));
 sg13g2_nand2_1 _2324_ (.Y(_0305_),
    .A(_1023_),
    .B(_1021_));
 sg13g2_nand2_1 _2325_ (.Y(_0306_),
    .A(_1073_),
    .B(_0222_));
 sg13g2_nand4_1 _2326_ (.B(_1031_),
    .C(_0305_),
    .A(_0975_),
    .Y(_0307_),
    .D(_0306_));
 sg13g2_a21oi_1 _2327_ (.A1(_0298_),
    .A2(_0304_),
    .Y(_0308_),
    .B1(_0307_));
 sg13g2_o21ai_1 _2328_ (.B1(_0308_),
    .Y(_0309_),
    .A1(_1008_),
    .A2(_0303_));
 sg13g2_buf_1 _2329_ (.A(_0309_),
    .X(_0310_));
 sg13g2_and2_1 _2330_ (.A(\simon1.state[6] ),
    .B(_1038_),
    .X(_0311_));
 sg13g2_a21o_1 _2331_ (.A2(_0310_),
    .A1(_1393_),
    .B1(_0311_),
    .X(_0312_));
 sg13g2_buf_1 _2332_ (.A(_0312_),
    .X(_0313_));
 sg13g2_nand2b_2 _2333_ (.Y(_0314_),
    .B(_0310_),
    .A_N(_1393_));
 sg13g2_nand2_1 _2334_ (.Y(_0315_),
    .A(net80),
    .B(_0314_));
 sg13g2_o21ai_1 _2335_ (.B1(_0315_),
    .Y(_0316_),
    .A1(net80),
    .A2(_0313_));
 sg13g2_nor2_1 _2336_ (.A(net47),
    .B(_0316_),
    .Y(_0109_));
 sg13g2_inv_1 _2337_ (.Y(_0317_),
    .A(_0015_));
 sg13g2_nor2b_2 _2338_ (.A(_1393_),
    .B_N(_0310_),
    .Y(_0318_));
 sg13g2_xor2_1 _2339_ (.B(_0957_),
    .A(net80),
    .X(_0319_));
 sg13g2_a22oi_1 _2340_ (.Y(_0320_),
    .B1(_0313_),
    .B2(_0319_),
    .A2(_0318_),
    .A1(_0317_));
 sg13g2_nor2_1 _2341_ (.A(net47),
    .B(_0320_),
    .Y(_0110_));
 sg13g2_buf_1 _2342_ (.A(_0969_),
    .X(_0321_));
 sg13g2_nand2b_1 _2343_ (.Y(_0322_),
    .B(_0016_),
    .A_N(_1393_));
 sg13g2_a21oi_1 _2344_ (.A1(_0310_),
    .A2(_0322_),
    .Y(_0323_),
    .B1(_0311_));
 sg13g2_nor3_1 _2345_ (.A(_0016_),
    .B(_1430_),
    .C(_0318_),
    .Y(_0324_));
 sg13g2_and2_1 _2346_ (.A(_0016_),
    .B(_1430_),
    .X(_0325_));
 sg13g2_nor4_1 _2347_ (.A(net49),
    .B(_0323_),
    .C(_0324_),
    .D(_0325_),
    .Y(_0111_));
 sg13g2_and3_1 _2348_ (.X(_0326_),
    .A(_0956_),
    .B(_0957_),
    .C(_0954_));
 sg13g2_buf_1 _2349_ (.A(_0326_),
    .X(_0327_));
 sg13g2_a21o_1 _2350_ (.A2(_0327_),
    .A1(_0314_),
    .B1(_0017_),
    .X(_0328_));
 sg13g2_or2_1 _2351_ (.X(_0329_),
    .B(_0311_),
    .A(_1393_));
 sg13g2_buf_1 _2352_ (.A(_0329_),
    .X(_0330_));
 sg13g2_nand3_1 _2353_ (.B(_0327_),
    .C(_0330_),
    .A(_0017_),
    .Y(_0331_));
 sg13g2_o21ai_1 _2354_ (.B1(net85),
    .Y(_0332_),
    .A1(_0310_),
    .A2(_0311_));
 sg13g2_a21oi_1 _2355_ (.A1(_0328_),
    .A2(_0331_),
    .Y(_0112_),
    .B1(_0332_));
 sg13g2_and2_1 _2356_ (.A(_0961_),
    .B(_0327_),
    .X(_0333_));
 sg13g2_nand2_1 _2357_ (.Y(_0334_),
    .A(_0330_),
    .B(_0333_));
 sg13g2_nand2_1 _2358_ (.Y(_0335_),
    .A(_0961_),
    .B(_0327_));
 sg13g2_nor2_1 _2359_ (.A(_0018_),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_a221oi_1 _2360_ (.B2(_0314_),
    .C1(_0332_),
    .B1(_0336_),
    .A1(_0018_),
    .Y(_0113_),
    .A2(_0334_));
 sg13g2_inv_1 _2361_ (.Y(_0337_),
    .A(_0019_));
 sg13g2_nor2_1 _2362_ (.A(_1014_),
    .B(_0335_),
    .Y(_0338_));
 sg13g2_xnor2_1 _2363_ (.Y(_0339_),
    .A(_0019_),
    .B(_0338_));
 sg13g2_a22oi_1 _2364_ (.Y(_0340_),
    .B1(_0313_),
    .B2(_0339_),
    .A2(_0318_),
    .A1(_0337_));
 sg13g2_nor2_1 _2365_ (.A(net47),
    .B(_0340_),
    .Y(_0114_));
 sg13g2_nor2_1 _2366_ (.A(_1048_),
    .B(_0335_),
    .Y(_0341_));
 sg13g2_nand2_1 _2367_ (.Y(_0342_),
    .A(_0330_),
    .B(_0341_));
 sg13g2_nand2b_1 _2368_ (.Y(_0343_),
    .B(_0333_),
    .A_N(_1048_));
 sg13g2_nor2_1 _2369_ (.A(_0020_),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_a221oi_1 _2370_ (.B2(_0314_),
    .C1(_0332_),
    .B1(_0344_),
    .A1(_0020_),
    .Y(_0115_),
    .A2(_0342_));
 sg13g2_inv_1 _2371_ (.Y(_0345_),
    .A(_0021_));
 sg13g2_nand2_1 _2372_ (.Y(_0346_),
    .A(_0963_),
    .B(_0341_));
 sg13g2_xnor2_1 _2373_ (.Y(_0347_),
    .A(_0345_),
    .B(_0346_));
 sg13g2_a22oi_1 _2374_ (.Y(_0348_),
    .B1(_0313_),
    .B2(_0347_),
    .A2(_0318_),
    .A1(_0345_));
 sg13g2_nor2_1 _2375_ (.A(net47),
    .B(_0348_),
    .Y(_0116_));
 sg13g2_nor2_1 _2376_ (.A(_1049_),
    .B(_0343_),
    .Y(_0349_));
 sg13g2_nand3_1 _2377_ (.B(_0330_),
    .C(_0349_),
    .A(_0022_),
    .Y(_0350_));
 sg13g2_a21o_1 _2378_ (.A2(_0349_),
    .A1(_0314_),
    .B1(_0022_),
    .X(_0351_));
 sg13g2_a21oi_1 _2379_ (.A1(_0350_),
    .A2(_0351_),
    .Y(_0117_),
    .B1(_0332_));
 sg13g2_inv_1 _2380_ (.Y(_0352_),
    .A(_0023_));
 sg13g2_nand2_1 _2381_ (.Y(_0353_),
    .A(_0958_),
    .B(_0349_));
 sg13g2_xnor2_1 _2382_ (.Y(_0354_),
    .A(_0352_),
    .B(_0353_));
 sg13g2_a22oi_1 _2383_ (.Y(_0355_),
    .B1(_0313_),
    .B2(_0354_),
    .A2(_0318_),
    .A1(_0352_));
 sg13g2_nor2_1 _2384_ (.A(net47),
    .B(_0355_),
    .Y(_0118_));
 sg13g2_a22oi_1 _2385_ (.Y(_0356_),
    .B1(\simon1.prev_btn[0] ),
    .B2(_1063_),
    .A2(net78),
    .A1(net87));
 sg13g2_nor2_1 _2386_ (.A(_1032_),
    .B(_0356_),
    .Y(_0119_));
 sg13g2_a22oi_1 _2387_ (.Y(_0357_),
    .B1(\simon1.prev_btn[1] ),
    .B2(_1063_),
    .A2(net78),
    .A1(net86));
 sg13g2_nor2_1 _2388_ (.A(_1032_),
    .B(_0357_),
    .Y(_0120_));
 sg13g2_buf_1 _2389_ (.A(net61),
    .X(_0358_));
 sg13g2_a22oi_1 _2390_ (.Y(_0359_),
    .B1(\simon1.prev_btn[2] ),
    .B2(_1063_),
    .A2(net78),
    .A1(_0940_));
 sg13g2_nor2_1 _2391_ (.A(_0358_),
    .B(_0359_),
    .Y(_0121_));
 sg13g2_a22oi_1 _2392_ (.Y(_0360_),
    .B1(\simon1.prev_btn[3] ),
    .B2(_1063_),
    .A2(net78),
    .A1(_0941_));
 sg13g2_nor2_1 _2393_ (.A(_0358_),
    .B(_0360_),
    .Y(_0122_));
 sg13g2_a21oi_1 _2394_ (.A1(_0974_),
    .A2(_1055_),
    .Y(_0361_),
    .B1(\simon1.score_ena ));
 sg13g2_nor2_1 _2395_ (.A(net45),
    .B(_0361_),
    .Y(_0123_));
 sg13g2_nor2_1 _2396_ (.A(_1009_),
    .B(_1013_),
    .Y(_0124_));
 sg13g2_and3_1 _2397_ (.X(_0134_),
    .A(_1437_),
    .B(_1051_),
    .C(_1050_));
 sg13g2_nand2b_1 _2398_ (.Y(_0362_),
    .B(_1030_),
    .A_N(_0025_));
 sg13g2_o21ai_1 _2399_ (.B1(_0362_),
    .Y(_0363_),
    .A1(_1433_),
    .A2(_0966_));
 sg13g2_nand2b_1 _2400_ (.Y(_0364_),
    .B(_0937_),
    .A_N(_0032_));
 sg13g2_o21ai_1 _2401_ (.B1(_0305_),
    .Y(_0365_),
    .A1(_1021_),
    .A2(_0364_));
 sg13g2_or3_1 _2402_ (.A(_1028_),
    .B(_1023_),
    .C(_1051_),
    .X(_0366_));
 sg13g2_o21ai_1 _2403_ (.B1(_0967_),
    .Y(_0367_),
    .A1(_1010_),
    .A2(_0366_));
 sg13g2_nor3_1 _2404_ (.A(_0363_),
    .B(_0365_),
    .C(_0367_),
    .Y(_0368_));
 sg13g2_inv_1 _2405_ (.Y(_0369_),
    .A(_1433_));
 sg13g2_nand3_1 _2406_ (.B(net20),
    .C(_1012_),
    .A(_0369_),
    .Y(_0370_));
 sg13g2_nand2_1 _2407_ (.Y(_0371_),
    .A(_0368_),
    .B(_0370_));
 sg13g2_buf_1 _2408_ (.A(_0371_),
    .X(_0372_));
 sg13g2_inv_1 _2409_ (.Y(_0373_),
    .A(net20));
 sg13g2_a21oi_1 _2410_ (.A1(_1028_),
    .A2(_0373_),
    .Y(_0374_),
    .B1(net59));
 sg13g2_nor3_1 _2411_ (.A(_0976_),
    .B(net17),
    .C(_0374_),
    .Y(_0375_));
 sg13g2_a21oi_1 _2412_ (.A1(_0976_),
    .A2(net17),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_nor2_1 _2413_ (.A(net45),
    .B(_0376_),
    .Y(_0135_));
 sg13g2_nand2_1 _2414_ (.Y(_0377_),
    .A(_1433_),
    .B(net20));
 sg13g2_a22oi_1 _2415_ (.Y(_0378_),
    .B1(_0377_),
    .B2(_1028_),
    .A2(_0369_),
    .A1(net59));
 sg13g2_nor2_2 _2416_ (.A(_0372_),
    .B(_0378_),
    .Y(_0379_));
 sg13g2_xor2_1 _2417_ (.B(_0980_),
    .A(_0976_),
    .X(_0380_));
 sg13g2_a22oi_1 _2418_ (.Y(_0381_),
    .B1(_0379_),
    .B2(_0380_),
    .A2(net17),
    .A1(_0980_));
 sg13g2_nor2_1 _2419_ (.A(net45),
    .B(_0381_),
    .Y(_0136_));
 sg13g2_nand2_1 _2420_ (.Y(_0382_),
    .A(_0976_),
    .B(_0980_));
 sg13g2_xnor2_1 _2421_ (.Y(_0383_),
    .A(\simon1.seq_counter[2] ),
    .B(_0382_));
 sg13g2_a22oi_1 _2422_ (.Y(_0384_),
    .B1(_0379_),
    .B2(_0383_),
    .A2(net17),
    .A1(\simon1.seq_counter[2] ));
 sg13g2_nor2_1 _2423_ (.A(net45),
    .B(_0384_),
    .Y(_0137_));
 sg13g2_xor2_1 _2424_ (.B(_0989_),
    .A(_0994_),
    .X(_0385_));
 sg13g2_a22oi_1 _2425_ (.Y(_0386_),
    .B1(_0379_),
    .B2(_0385_),
    .A2(net17),
    .A1(_0994_));
 sg13g2_nor2_1 _2426_ (.A(net45),
    .B(_0386_),
    .Y(_0138_));
 sg13g2_nand2_1 _2427_ (.Y(_0387_),
    .A(_0994_),
    .B(_0989_));
 sg13g2_xnor2_1 _2428_ (.Y(_0388_),
    .A(_0990_),
    .B(_0387_));
 sg13g2_a22oi_1 _2429_ (.Y(_0389_),
    .B1(_0379_),
    .B2(_0388_),
    .A2(net17),
    .A1(_0990_));
 sg13g2_nor2_1 _2430_ (.A(net45),
    .B(_0389_),
    .Y(_0139_));
 sg13g2_xnor2_1 _2431_ (.Y(_0390_),
    .A(\simon1.seq_counter[5] ),
    .B(_1000_));
 sg13g2_a22oi_1 _2432_ (.Y(_0391_),
    .B1(_0379_),
    .B2(_0390_),
    .A2(net17),
    .A1(\simon1.seq_counter[5] ));
 sg13g2_nor2_1 _2433_ (.A(net45),
    .B(_0391_),
    .Y(_0140_));
 sg13g2_xnor2_1 _2434_ (.Y(_0392_),
    .A(\simon1.seq_counter[6] ),
    .B(_1004_));
 sg13g2_a22oi_1 _2435_ (.Y(_0393_),
    .B1(_0379_),
    .B2(_0392_),
    .A2(net17),
    .A1(\simon1.seq_counter[6] ));
 sg13g2_nor2_1 _2436_ (.A(net45),
    .B(_0393_),
    .Y(_0141_));
 sg13g2_buf_1 _2437_ (.A(net61),
    .X(_0394_));
 sg13g2_nor2_1 _2438_ (.A(_1433_),
    .B(net20),
    .Y(_0395_));
 sg13g2_or2_1 _2439_ (.X(_0396_),
    .B(_1051_),
    .A(_0946_));
 sg13g2_o21ai_1 _2440_ (.B1(_0396_),
    .Y(_0397_),
    .A1(net52),
    .A2(_1012_));
 sg13g2_a21o_1 _2441_ (.A2(_0395_),
    .A1(_1012_),
    .B1(_0397_),
    .X(_0398_));
 sg13g2_buf_1 _2442_ (.A(_0398_),
    .X(_0399_));
 sg13g2_nor2_1 _2443_ (.A(_1013_),
    .B(_0395_),
    .Y(_0400_));
 sg13g2_mux2_1 _2444_ (.A0(net16),
    .A1(_0400_),
    .S(_0978_),
    .X(_0401_));
 sg13g2_nor2_1 _2445_ (.A(net44),
    .B(_0401_),
    .Y(_0142_));
 sg13g2_nor3_1 _2446_ (.A(_0978_),
    .B(_1013_),
    .C(_0395_),
    .Y(_0402_));
 sg13g2_o21ai_1 _2447_ (.B1(_0981_),
    .Y(_0403_),
    .A1(net16),
    .A2(_0402_));
 sg13g2_nand3b_1 _2448_ (.B(_0400_),
    .C(_0978_),
    .Y(_0404_),
    .A_N(_0981_));
 sg13g2_a21oi_1 _2449_ (.A1(_0403_),
    .A2(_0404_),
    .Y(_0143_),
    .B1(net48));
 sg13g2_nand2_1 _2450_ (.Y(_0405_),
    .A(_0978_),
    .B(_0981_));
 sg13g2_xor2_1 _2451_ (.B(_0405_),
    .A(_0027_),
    .X(_0406_));
 sg13g2_a22oi_1 _2452_ (.Y(_0407_),
    .B1(_0406_),
    .B2(_0400_),
    .A2(_0399_),
    .A1(\simon1.seq_length[2] ));
 sg13g2_nor2_1 _2453_ (.A(net44),
    .B(_0407_),
    .Y(_0144_));
 sg13g2_nand3_1 _2454_ (.B(_0981_),
    .C(\simon1.seq_length[2] ),
    .A(_0978_),
    .Y(_0408_));
 sg13g2_xnor2_1 _2455_ (.Y(_0409_),
    .A(_0028_),
    .B(_0408_));
 sg13g2_nor3_1 _2456_ (.A(net52),
    .B(net16),
    .C(_0409_),
    .Y(_0410_));
 sg13g2_a21oi_1 _2457_ (.A1(\simon1.seq_length[3] ),
    .A2(_0399_),
    .Y(_0411_),
    .B1(_0410_));
 sg13g2_nor2_1 _2458_ (.A(net44),
    .B(_0411_),
    .Y(_0145_));
 sg13g2_inv_1 _2459_ (.Y(_0412_),
    .A(\simon1.seq_length[3] ));
 sg13g2_nor2_1 _2460_ (.A(_0412_),
    .B(_0408_),
    .Y(_0413_));
 sg13g2_xor2_1 _2461_ (.B(_0413_),
    .A(_0029_),
    .X(_0414_));
 sg13g2_nor3_1 _2462_ (.A(net52),
    .B(net16),
    .C(_0414_),
    .Y(_0415_));
 sg13g2_a21o_1 _2463_ (.A2(net16),
    .A1(\simon1.seq_length[4] ),
    .B1(_0415_),
    .X(_0416_));
 sg13g2_and2_1 _2464_ (.A(net63),
    .B(_0416_),
    .X(_0146_));
 sg13g2_nand2_1 _2465_ (.Y(_0417_),
    .A(\simon1.seq_length[4] ),
    .B(_0413_));
 sg13g2_xnor2_1 _2466_ (.Y(_0418_),
    .A(_0030_),
    .B(_0417_));
 sg13g2_nor3_1 _2467_ (.A(net52),
    .B(net16),
    .C(_0418_),
    .Y(_0419_));
 sg13g2_a21o_1 _2468_ (.A2(net16),
    .A1(\simon1.seq_length[5] ),
    .B1(_0419_),
    .X(_0420_));
 sg13g2_and2_1 _2469_ (.A(net63),
    .B(_0420_),
    .X(_0147_));
 sg13g2_nand3_1 _2470_ (.B(\simon1.seq_length[5] ),
    .C(_0413_),
    .A(\simon1.seq_length[4] ),
    .Y(_0421_));
 sg13g2_xnor2_1 _2471_ (.Y(_0422_),
    .A(_0031_),
    .B(_0421_));
 sg13g2_nor3_1 _2472_ (.A(net52),
    .B(_0398_),
    .C(_0422_),
    .Y(_0423_));
 sg13g2_a21o_1 _2473_ (.A2(net16),
    .A1(\simon1.seq_length[6] ),
    .B1(_0423_),
    .X(_0424_));
 sg13g2_and2_1 _2474_ (.A(net63),
    .B(_0424_),
    .X(_0148_));
 sg13g2_nor2_1 _2475_ (.A(_0937_),
    .B(_0943_),
    .Y(_0425_));
 sg13g2_nor2b_1 _2476_ (.A(_0425_),
    .B_N(_1126_),
    .Y(_0426_));
 sg13g2_nor2b_1 _2477_ (.A(_1134_),
    .B_N(_0220_),
    .Y(_0427_));
 sg13g2_nor4_1 _2478_ (.A(_1133_),
    .B(_0223_),
    .C(_0426_),
    .D(_0427_),
    .Y(_0428_));
 sg13g2_buf_1 _2479_ (.A(_0428_),
    .X(_0429_));
 sg13g2_buf_1 _2480_ (.A(net19),
    .X(_0430_));
 sg13g2_nand2_1 _2481_ (.Y(_0431_),
    .A(_1122_),
    .B(net84));
 sg13g2_nor2_1 _2482_ (.A(_0026_),
    .B(_1120_),
    .Y(_0432_));
 sg13g2_o21ai_1 _2483_ (.B1(_1124_),
    .Y(_0433_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_o21ai_1 _2484_ (.B1(_1120_),
    .Y(_0434_),
    .A1(_0956_),
    .A2(_1131_));
 sg13g2_nor2_2 _2485_ (.A(_1053_),
    .B(_0425_),
    .Y(_0435_));
 sg13g2_a22oi_1 _2486_ (.Y(_0436_),
    .B1(_0434_),
    .B2(_0435_),
    .A2(_0433_),
    .A1(net58));
 sg13g2_o21ai_1 _2487_ (.B1(net62),
    .Y(_0437_),
    .A1(\simon1.sound_freq[0] ),
    .A2(net18));
 sg13g2_a21oi_1 _2488_ (.A1(_0430_),
    .A2(_0436_),
    .Y(_0149_),
    .B1(_0437_));
 sg13g2_nand2b_1 _2489_ (.Y(_0438_),
    .B(\simon1.sound_freq[1] ),
    .A_N(net19));
 sg13g2_nor2_1 _2490_ (.A(_1120_),
    .B(net84),
    .Y(_0439_));
 sg13g2_a21oi_1 _2491_ (.A1(_1121_),
    .A2(net84),
    .Y(_0440_),
    .B1(_0439_));
 sg13g2_or2_1 _2492_ (.X(_0441_),
    .B(_0239_),
    .A(_0233_));
 sg13g2_nor2_1 _2493_ (.A(_1429_),
    .B(_0966_),
    .Y(_0442_));
 sg13g2_nor4_1 _2494_ (.A(_0946_),
    .B(_1028_),
    .C(_0944_),
    .D(_1023_),
    .Y(_0443_));
 sg13g2_buf_1 _2495_ (.A(_0443_),
    .X(_0444_));
 sg13g2_a221oi_1 _2496_ (.B2(_0442_),
    .C1(net43),
    .B1(_0441_),
    .A1(net58),
    .Y(_0445_),
    .A2(_0440_));
 sg13g2_o21ai_1 _2497_ (.B1(_1130_),
    .Y(_0446_),
    .A1(_1129_),
    .A2(_0319_));
 sg13g2_nand2_1 _2498_ (.Y(_0447_),
    .A(_0435_),
    .B(_0446_));
 sg13g2_xnor2_1 _2499_ (.Y(_0448_),
    .A(_0950_),
    .B(_0947_));
 sg13g2_a22oi_1 _2500_ (.Y(_0449_),
    .B1(_0448_),
    .B2(net43),
    .A2(_0447_),
    .A1(_0445_));
 sg13g2_nand2_1 _2501_ (.Y(_0450_),
    .A(net18),
    .B(_0449_));
 sg13g2_buf_1 _2502_ (.A(net61),
    .X(_0451_));
 sg13g2_a21oi_1 _2503_ (.A1(_0438_),
    .A2(_0450_),
    .Y(_0150_),
    .B1(net42));
 sg13g2_nor2_1 _2504_ (.A(_1334_),
    .B(net18),
    .Y(_0452_));
 sg13g2_nor2b_1 _2505_ (.A(_1046_),
    .B_N(_0954_),
    .Y(_0453_));
 sg13g2_nor3_1 _2506_ (.A(net80),
    .B(_0957_),
    .C(_0954_),
    .Y(_0454_));
 sg13g2_o21ai_1 _2507_ (.B1(net76),
    .Y(_0455_),
    .A1(_0453_),
    .A2(_0454_));
 sg13g2_nand3_1 _2508_ (.B(_1123_),
    .C(_0455_),
    .A(_0435_),
    .Y(_0456_));
 sg13g2_o21ai_1 _2509_ (.B1(_0456_),
    .Y(_0457_),
    .A1(net83),
    .A2(_1064_));
 sg13g2_a21oi_1 _2510_ (.A1(_1168_),
    .A2(net43),
    .Y(_0458_),
    .B1(_0457_));
 sg13g2_and2_1 _2511_ (.A(net19),
    .B(_0458_),
    .X(_0459_));
 sg13g2_nor3_1 _2512_ (.A(net49),
    .B(_0452_),
    .C(_0459_),
    .Y(_0151_));
 sg13g2_xnor2_1 _2513_ (.Y(_0460_),
    .A(_0017_),
    .B(_0453_));
 sg13g2_o21ai_1 _2514_ (.B1(_1130_),
    .Y(_0461_),
    .A1(_1129_),
    .A2(_0460_));
 sg13g2_nand2_1 _2515_ (.Y(_0462_),
    .A(_0435_),
    .B(_0461_));
 sg13g2_nand2_1 _2516_ (.Y(_0463_),
    .A(_1120_),
    .B(net84));
 sg13g2_nand2_1 _2517_ (.Y(_0464_),
    .A(net58),
    .B(_0463_));
 sg13g2_a21oi_1 _2518_ (.A1(net76),
    .A2(_0933_),
    .Y(_0465_),
    .B1(_0464_));
 sg13g2_a221oi_1 _2519_ (.B2(net43),
    .C1(_0465_),
    .B1(_0242_),
    .A1(_0442_),
    .Y(_0466_),
    .A2(_0239_));
 sg13g2_nand3_1 _2520_ (.B(_0462_),
    .C(_0466_),
    .A(net19),
    .Y(_0467_));
 sg13g2_o21ai_1 _2521_ (.B1(_0467_),
    .Y(_0468_),
    .A1(\simon1.sound_freq[3] ),
    .A2(_0430_));
 sg13g2_nor2_1 _2522_ (.A(net44),
    .B(_0468_),
    .Y(_0152_));
 sg13g2_nand2_1 _2523_ (.Y(_0469_),
    .A(net76),
    .B(_0439_));
 sg13g2_o21ai_1 _2524_ (.B1(_0469_),
    .Y(_0470_),
    .A1(net76),
    .A2(_0463_));
 sg13g2_nor2_1 _2525_ (.A(_0945_),
    .B(_1131_),
    .Y(_0471_));
 sg13g2_o21ai_1 _2526_ (.B1(_0017_),
    .Y(_0472_),
    .A1(_1046_),
    .A2(_1019_));
 sg13g2_xor2_1 _2527_ (.B(_0472_),
    .A(_0018_),
    .X(_0473_));
 sg13g2_nand3_1 _2528_ (.B(_0947_),
    .C(net43),
    .A(_0950_),
    .Y(_0474_));
 sg13g2_o21ai_1 _2529_ (.B1(_0474_),
    .Y(_0475_),
    .A1(_1064_),
    .A2(_0248_));
 sg13g2_a221oi_1 _2530_ (.B2(_0473_),
    .C1(_0475_),
    .B1(_0471_),
    .A1(net58),
    .Y(_0476_),
    .A2(_0470_));
 sg13g2_o21ai_1 _2531_ (.B1(net62),
    .Y(_0477_),
    .A1(_1326_),
    .A2(net19));
 sg13g2_a21oi_1 _2532_ (.A1(net18),
    .A2(_0476_),
    .Y(_0153_),
    .B1(_0477_));
 sg13g2_nand2b_1 _2533_ (.Y(_0478_),
    .B(net75),
    .A_N(_0429_));
 sg13g2_nor3_1 _2534_ (.A(\simon1.millis_counter[4] ),
    .B(_0961_),
    .C(_0453_),
    .Y(_0479_));
 sg13g2_nor2_1 _2535_ (.A(_1124_),
    .B(_0479_),
    .Y(_0480_));
 sg13g2_nor4_1 _2536_ (.A(_0933_),
    .B(_0033_),
    .C(net43),
    .D(_0480_),
    .Y(_0481_));
 sg13g2_nand2_1 _2537_ (.Y(_0482_),
    .A(net18),
    .B(_0481_));
 sg13g2_a21oi_1 _2538_ (.A1(_0478_),
    .A2(_0482_),
    .Y(_0154_),
    .B1(net42));
 sg13g2_a21o_1 _2539_ (.A2(_0026_),
    .A1(net76),
    .B1(_1123_),
    .X(_0483_));
 sg13g2_nor3_1 _2540_ (.A(_1053_),
    .B(net84),
    .C(_0480_),
    .Y(_0484_));
 sg13g2_a221oi_1 _2541_ (.B2(net58),
    .C1(_0484_),
    .B1(_0483_),
    .A1(_0253_),
    .Y(_0485_),
    .A2(_0444_));
 sg13g2_o21ai_1 _2542_ (.B1(_0485_),
    .Y(_0486_),
    .A1(net81),
    .A2(_1064_));
 sg13g2_nand2_1 _2543_ (.Y(_0487_),
    .A(net18),
    .B(_0486_));
 sg13g2_nand2b_1 _2544_ (.Y(_0488_),
    .B(net73),
    .A_N(_0429_));
 sg13g2_a21oi_1 _2545_ (.A1(_0487_),
    .A2(_0488_),
    .Y(_0155_),
    .B1(net42));
 sg13g2_inv_1 _2546_ (.Y(_0489_),
    .A(_1331_));
 sg13g2_nor3_1 _2547_ (.A(net81),
    .B(net83),
    .C(_1064_),
    .Y(_0490_));
 sg13g2_nand2_1 _2548_ (.Y(_0491_),
    .A(_1130_),
    .B(_0479_));
 sg13g2_nor2b_1 _2549_ (.A(net76),
    .B_N(_1023_),
    .Y(_0492_));
 sg13g2_nand2b_1 _2550_ (.Y(_0493_),
    .B(_0463_),
    .A_N(_0439_));
 sg13g2_a21oi_1 _2551_ (.A1(_0492_),
    .A2(_0493_),
    .Y(_0494_),
    .B1(net43));
 sg13g2_o21ai_1 _2552_ (.B1(_0494_),
    .Y(_0495_),
    .A1(_0945_),
    .A2(_0491_));
 sg13g2_nand2b_1 _2553_ (.Y(_0496_),
    .B(net43),
    .A_N(_0227_));
 sg13g2_o21ai_1 _2554_ (.B1(_0496_),
    .Y(_0497_),
    .A1(_0490_),
    .A2(_0495_));
 sg13g2_mux2_1 _2555_ (.A0(_0489_),
    .A1(_0497_),
    .S(net19),
    .X(_0498_));
 sg13g2_nor2_1 _2556_ (.A(net44),
    .B(_0498_),
    .Y(_0156_));
 sg13g2_inv_1 _2557_ (.Y(_0499_),
    .A(_0472_));
 sg13g2_nand3_1 _2558_ (.B(_0471_),
    .C(_0499_),
    .A(_0018_),
    .Y(_0500_));
 sg13g2_nand2_1 _2559_ (.Y(_0501_),
    .A(net76),
    .B(_0024_));
 sg13g2_nand4_1 _2560_ (.B(_0937_),
    .C(_0431_),
    .A(_1024_),
    .Y(_0502_),
    .D(_0501_));
 sg13g2_o21ai_1 _2561_ (.B1(_0442_),
    .Y(_0503_),
    .A1(net81),
    .A2(net83));
 sg13g2_nand4_1 _2562_ (.B(_0500_),
    .C(_0502_),
    .A(_0496_),
    .Y(_0504_),
    .D(_0503_));
 sg13g2_nand2_1 _2563_ (.Y(_0505_),
    .A(net18),
    .B(_0504_));
 sg13g2_nand2b_1 _2564_ (.Y(_0506_),
    .B(net74),
    .A_N(net19));
 sg13g2_a21oi_1 _2565_ (.A1(_0505_),
    .A2(_0506_),
    .Y(_0157_),
    .B1(_0451_));
 sg13g2_xor2_1 _2566_ (.B(net84),
    .A(_1121_),
    .X(_0507_));
 sg13g2_o21ai_1 _2567_ (.B1(_1130_),
    .Y(_0508_),
    .A1(_1129_),
    .A2(_0479_));
 sg13g2_a221oi_1 _2568_ (.B2(_0435_),
    .C1(_0475_),
    .B1(_0508_),
    .A1(_1024_),
    .Y(_0509_),
    .A2(_0507_));
 sg13g2_o21ai_1 _2569_ (.B1(_0231_),
    .Y(_0510_),
    .A1(_1328_),
    .A2(net19));
 sg13g2_a21oi_1 _2570_ (.A1(net18),
    .A2(_0509_),
    .Y(_0158_),
    .B1(_0510_));
 sg13g2_xnor2_1 _2571_ (.Y(_0511_),
    .A(\simon1.sound_gen_inst.tick_counter[0] ),
    .B(\simon1.sound_freq[0] ));
 sg13g2_nor2_1 _2572_ (.A(_0394_),
    .B(_0511_),
    .Y(_0160_));
 sg13g2_nor2_1 _2573_ (.A(_1353_),
    .B(net34),
    .Y(_0512_));
 sg13g2_and4_1 _2574_ (.A(_1327_),
    .B(_1330_),
    .C(_1333_),
    .D(_1335_),
    .X(_0513_));
 sg13g2_buf_1 _2575_ (.A(_0513_),
    .X(_0514_));
 sg13g2_buf_1 _2576_ (.A(net40),
    .X(_0515_));
 sg13g2_nor3_1 _2577_ (.A(_1361_),
    .B(_1366_),
    .C(_1377_),
    .Y(_0516_));
 sg13g2_inv_1 _2578_ (.Y(_0517_),
    .A(_1381_));
 sg13g2_xnor2_1 _2579_ (.Y(_0518_),
    .A(net74),
    .B(net70));
 sg13g2_nand3_1 _2580_ (.B(net66),
    .C(\simon1.sound_gen_inst.tick_counter[5] ),
    .A(_1326_),
    .Y(_0519_));
 sg13g2_a21oi_1 _2581_ (.A1(_1331_),
    .A2(net71),
    .Y(_0520_),
    .B1(\simon1.sound_freq[5] ));
 sg13g2_a221oi_1 _2582_ (.B2(_1326_),
    .C1(net65),
    .B1(net66),
    .A1(_1331_),
    .Y(_0521_),
    .A2(net71));
 sg13g2_a21o_1 _2583_ (.A2(_0520_),
    .A1(_0519_),
    .B1(_0521_),
    .X(_0522_));
 sg13g2_o21ai_1 _2584_ (.B1(net71),
    .Y(_0523_),
    .A1(\simon1.sound_freq[6] ),
    .A2(\simon1.sound_gen_inst.tick_counter[6] ));
 sg13g2_and2_1 _2585_ (.A(_0489_),
    .B(_0523_),
    .X(_0524_));
 sg13g2_a21o_1 _2586_ (.A2(_0522_),
    .A1(_1378_),
    .B1(_0524_),
    .X(_0525_));
 sg13g2_a21oi_1 _2587_ (.A1(_0519_),
    .A2(_0520_),
    .Y(_0526_),
    .B1(_0521_));
 sg13g2_or2_1 _2588_ (.X(_0527_),
    .B(net71),
    .A(net67));
 sg13g2_a21oi_1 _2589_ (.A1(_0526_),
    .A2(_0527_),
    .Y(_0528_),
    .B1(_1332_));
 sg13g2_inv_1 _2590_ (.Y(_0529_),
    .A(\simon1.sound_freq[3] ));
 sg13g2_a21oi_1 _2591_ (.A1(_1334_),
    .A2(_1348_),
    .Y(_0530_),
    .B1(_1346_));
 sg13g2_nand3_1 _2592_ (.B(_1346_),
    .C(_1348_),
    .A(_1334_),
    .Y(_0531_));
 sg13g2_o21ai_1 _2593_ (.B1(_0531_),
    .Y(_0532_),
    .A1(_0529_),
    .A2(_0530_));
 sg13g2_nor2_1 _2594_ (.A(\simon1.sound_freq[1] ),
    .B(\simon1.sound_gen_inst.tick_counter[1] ),
    .Y(_0533_));
 sg13g2_a22oi_1 _2595_ (.Y(_0534_),
    .B1(\simon1.sound_freq[1] ),
    .B2(\simon1.sound_gen_inst.tick_counter[1] ),
    .A2(\simon1.sound_freq[0] ),
    .A1(\simon1.sound_gen_inst.tick_counter[0] ));
 sg13g2_xnor2_1 _2596_ (.Y(_0535_),
    .A(\simon1.sound_freq[3] ),
    .B(_1346_));
 sg13g2_xnor2_1 _2597_ (.Y(_0536_),
    .A(_1334_),
    .B(_1348_));
 sg13g2_nor4_1 _2598_ (.A(_0533_),
    .B(_0534_),
    .C(_0535_),
    .D(_0536_),
    .Y(_0537_));
 sg13g2_xnor2_1 _2599_ (.Y(_0538_),
    .A(_1326_),
    .B(net66));
 sg13g2_xnor2_1 _2600_ (.Y(_0539_),
    .A(net75),
    .B(net65));
 sg13g2_xnor2_1 _2601_ (.Y(_0540_),
    .A(_1331_),
    .B(net71));
 sg13g2_xnor2_1 _2602_ (.Y(_0541_),
    .A(\simon1.sound_freq[6] ),
    .B(\simon1.sound_gen_inst.tick_counter[6] ));
 sg13g2_nor4_2 _2603_ (.A(_0538_),
    .B(_0539_),
    .C(_0540_),
    .Y(_0542_),
    .D(_0541_));
 sg13g2_o21ai_1 _2604_ (.B1(_0542_),
    .Y(_0543_),
    .A1(_0532_),
    .A2(_0537_));
 sg13g2_o21ai_1 _2605_ (.B1(_0543_),
    .Y(_0544_),
    .A1(_0525_),
    .A2(_0528_));
 sg13g2_xnor2_1 _2606_ (.Y(_0545_),
    .A(_0518_),
    .B(_0544_));
 sg13g2_inv_1 _2607_ (.Y(_0546_),
    .A(net75));
 sg13g2_nand2_1 _2608_ (.Y(_0547_),
    .A(_1334_),
    .B(_1348_));
 sg13g2_o21ai_1 _2609_ (.B1(_0547_),
    .Y(_0548_),
    .A1(_0533_),
    .A2(_0534_));
 sg13g2_buf_2 _2610_ (.A(_0548_),
    .X(_0549_));
 sg13g2_nor2_1 _2611_ (.A(_1334_),
    .B(_1348_),
    .Y(_0550_));
 sg13g2_nor3_2 _2612_ (.A(_0538_),
    .B(_0550_),
    .C(_0535_),
    .Y(_0551_));
 sg13g2_nor2_2 _2613_ (.A(_1326_),
    .B(net66),
    .Y(_0552_));
 sg13g2_a22oi_1 _2614_ (.Y(_0553_),
    .B1(net66),
    .B2(_1326_),
    .A2(_1346_),
    .A1(\simon1.sound_freq[3] ));
 sg13g2_buf_1 _2615_ (.A(_0553_),
    .X(_0554_));
 sg13g2_nor2_1 _2616_ (.A(_0552_),
    .B(_0554_),
    .Y(_0555_));
 sg13g2_a21oi_2 _2617_ (.B1(_0555_),
    .Y(_0556_),
    .A2(_0551_),
    .A1(_0549_));
 sg13g2_or2_1 _2618_ (.X(_0557_),
    .B(_0537_),
    .A(_0532_));
 sg13g2_buf_8 _2619_ (.A(_0557_),
    .X(_0558_));
 sg13g2_and4_1 _2620_ (.A(net75),
    .B(_1326_),
    .C(net66),
    .D(net65),
    .X(_0559_));
 sg13g2_a221oi_1 _2621_ (.B2(_0559_),
    .C1(_0541_),
    .B1(_0558_),
    .A1(_0546_),
    .Y(_0560_),
    .A2(_0556_));
 sg13g2_nand2_2 _2622_ (.Y(_0561_),
    .A(_1359_),
    .B(_0556_));
 sg13g2_or2_1 _2623_ (.X(_0562_),
    .B(_1348_),
    .A(_1334_));
 sg13g2_buf_1 _2624_ (.A(_0562_),
    .X(_0563_));
 sg13g2_and2_1 _2625_ (.A(_0549_),
    .B(_0563_),
    .X(_0564_));
 sg13g2_and4_1 _2626_ (.A(net75),
    .B(net65),
    .C(_0555_),
    .D(_0535_),
    .X(_0565_));
 sg13g2_nand2_1 _2627_ (.Y(_0566_),
    .A(net75),
    .B(net65));
 sg13g2_or4_1 _2628_ (.A(_0552_),
    .B(_0554_),
    .C(_0535_),
    .D(_0566_),
    .X(_0567_));
 sg13g2_a21oi_1 _2629_ (.A1(_0549_),
    .A2(_0563_),
    .Y(_0568_),
    .B1(_0567_));
 sg13g2_a221oi_1 _2630_ (.B2(_0565_),
    .C1(_0568_),
    .B1(_0564_),
    .A1(_0546_),
    .Y(_0569_),
    .A2(_1359_));
 sg13g2_and3_1 _2631_ (.X(_0570_),
    .A(_0560_),
    .B(_0561_),
    .C(_0569_));
 sg13g2_xor2_1 _2632_ (.B(net67),
    .A(net73),
    .X(_0571_));
 sg13g2_xnor2_1 _2633_ (.Y(_0572_),
    .A(_0538_),
    .B(_0558_));
 sg13g2_nand3_1 _2634_ (.B(_0563_),
    .C(_0535_),
    .A(_0549_),
    .Y(_0573_));
 sg13g2_a21o_1 _2635_ (.A2(_0563_),
    .A1(_0549_),
    .B1(_0535_),
    .X(_0574_));
 sg13g2_nand2_2 _2636_ (.Y(_0575_),
    .A(_0573_),
    .B(_0574_));
 sg13g2_nor4_2 _2637_ (.A(_0571_),
    .B(_0572_),
    .C(_0575_),
    .Y(_0576_),
    .D(_0561_));
 sg13g2_nand3_1 _2638_ (.B(_0573_),
    .C(_0574_),
    .A(_1359_),
    .Y(_0577_));
 sg13g2_o21ai_1 _2639_ (.B1(_0535_),
    .Y(_0578_),
    .A1(_0552_),
    .A2(_0554_));
 sg13g2_a21oi_1 _2640_ (.A1(_0549_),
    .A2(_0563_),
    .Y(_0579_),
    .B1(_0578_));
 sg13g2_a21oi_1 _2641_ (.A1(_1359_),
    .A2(_0556_),
    .Y(_0580_),
    .B1(_0579_));
 sg13g2_nand2_1 _2642_ (.Y(_0581_),
    .A(_0546_),
    .B(_0541_));
 sg13g2_a221oi_1 _2643_ (.B2(_0580_),
    .C1(_0581_),
    .B1(_0577_),
    .A1(_0572_),
    .Y(_0582_),
    .A2(_0561_));
 sg13g2_nor2_1 _2644_ (.A(\simon1.sound_freq[6] ),
    .B(net67),
    .Y(_0583_));
 sg13g2_a21oi_1 _2645_ (.A1(net73),
    .A2(net67),
    .Y(_0584_),
    .B1(_1358_));
 sg13g2_o21ai_1 _2646_ (.B1(_0584_),
    .Y(_0585_),
    .A1(_0552_),
    .A2(_0554_));
 sg13g2_a21oi_1 _2647_ (.A1(net73),
    .A2(net67),
    .Y(_0586_),
    .B1(net75));
 sg13g2_o21ai_1 _2648_ (.B1(_0586_),
    .Y(_0587_),
    .A1(_0552_),
    .A2(_0554_));
 sg13g2_a22oi_1 _2649_ (.Y(_0588_),
    .B1(_0585_),
    .B2(_0587_),
    .A2(_0551_),
    .A1(_0549_));
 sg13g2_nand2_1 _2650_ (.Y(_0589_),
    .A(_0546_),
    .B(_1359_));
 sg13g2_a21oi_1 _2651_ (.A1(net73),
    .A2(net67),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_nor3_1 _2652_ (.A(_0583_),
    .B(_0588_),
    .C(_0590_),
    .Y(_0591_));
 sg13g2_xor2_1 _2653_ (.B(_0591_),
    .A(_0540_),
    .X(_0592_));
 sg13g2_nor4_2 _2654_ (.A(_0570_),
    .B(_0576_),
    .C(_0582_),
    .Y(_0593_),
    .D(_0592_));
 sg13g2_xnor2_1 _2655_ (.Y(_0594_),
    .A(_1328_),
    .B(net68));
 sg13g2_a21o_1 _2656_ (.A2(_0551_),
    .A1(_0549_),
    .B1(_0555_),
    .X(_0595_));
 sg13g2_nor4_2 _2657_ (.A(_0518_),
    .B(_0539_),
    .C(_0540_),
    .Y(_0596_),
    .D(_0541_));
 sg13g2_or2_1 _2658_ (.X(_0597_),
    .B(net70),
    .A(net74));
 sg13g2_a22oi_1 _2659_ (.Y(_0598_),
    .B1(net71),
    .B2(_1331_),
    .A2(_1356_),
    .A1(_1332_));
 sg13g2_o21ai_1 _2660_ (.B1(_0598_),
    .Y(_0599_),
    .A1(_0583_),
    .A2(_0566_));
 sg13g2_or2_1 _2661_ (.X(_0600_),
    .B(net71),
    .A(_1331_));
 sg13g2_and2_1 _2662_ (.A(net74),
    .B(net70),
    .X(_0601_));
 sg13g2_a21o_1 _2663_ (.A2(_0600_),
    .A1(_0599_),
    .B1(_0601_),
    .X(_0602_));
 sg13g2_a22oi_1 _2664_ (.Y(_0603_),
    .B1(_0597_),
    .B2(_0602_),
    .A2(_0596_),
    .A1(_0595_));
 sg13g2_xnor2_1 _2665_ (.Y(_0604_),
    .A(_0594_),
    .B(_0603_));
 sg13g2_inv_1 _2666_ (.Y(_0605_),
    .A(_0604_));
 sg13g2_a221oi_1 _2667_ (.B2(_0593_),
    .C1(_0605_),
    .B1(_0545_),
    .A1(_0516_),
    .Y(_0606_),
    .A2(_0517_));
 sg13g2_buf_1 _2668_ (.A(_0606_),
    .X(_0607_));
 sg13g2_inv_1 _2669_ (.Y(_0608_),
    .A(_1328_));
 sg13g2_o21ai_1 _2670_ (.B1(net68),
    .Y(_0609_),
    .A1(\simon1.sound_freq[8] ),
    .A2(\simon1.sound_gen_inst.tick_counter[8] ));
 sg13g2_nor3_1 _2671_ (.A(net74),
    .B(net68),
    .C(net70),
    .Y(_0610_));
 sg13g2_a21o_1 _2672_ (.A2(_0609_),
    .A1(_0608_),
    .B1(_0610_),
    .X(_0611_));
 sg13g2_buf_1 _2673_ (.A(_0611_),
    .X(_0612_));
 sg13g2_buf_1 _2674_ (.A(_0612_),
    .X(_0613_));
 sg13g2_a21oi_1 _2675_ (.A1(_1378_),
    .A2(_0522_),
    .Y(_0614_),
    .B1(_0524_));
 sg13g2_a21o_1 _2676_ (.A2(_0527_),
    .A1(_0526_),
    .B1(net73),
    .X(_0615_));
 sg13g2_a21o_1 _2677_ (.A2(net70),
    .A1(net74),
    .B1(net68),
    .X(_0616_));
 sg13g2_and3_1 _2678_ (.X(_0617_),
    .A(_1329_),
    .B(net68),
    .C(net70));
 sg13g2_a21o_1 _2679_ (.A2(_0616_),
    .A1(_1328_),
    .B1(_0617_),
    .X(_0618_));
 sg13g2_a221oi_1 _2680_ (.B2(_0542_),
    .C1(_0618_),
    .B1(_0558_),
    .A1(_0614_),
    .Y(_0619_),
    .A2(_0615_));
 sg13g2_buf_2 _2681_ (.A(_0619_),
    .X(_0620_));
 sg13g2_buf_8 _2682_ (.A(_0620_),
    .X(_0621_));
 sg13g2_buf_1 _2683_ (.A(_0034_),
    .X(_0622_));
 sg13g2_o21ai_1 _2684_ (.B1(_0622_),
    .Y(_0623_),
    .A1(net32),
    .A2(net21));
 sg13g2_nor2_1 _2685_ (.A(net32),
    .B(net21),
    .Y(_0624_));
 sg13g2_nand2b_1 _2686_ (.Y(_0625_),
    .B(_0624_),
    .A_N(_0622_));
 sg13g2_nand2_1 _2687_ (.Y(_0626_),
    .A(_0623_),
    .B(_0625_));
 sg13g2_xnor2_1 _2688_ (.Y(_0627_),
    .A(_0607_),
    .B(_0626_));
 sg13g2_nor2_1 _2689_ (.A(net33),
    .B(_0627_),
    .Y(_0628_));
 sg13g2_nor3_1 _2690_ (.A(net49),
    .B(_0512_),
    .C(_0628_),
    .Y(_0161_));
 sg13g2_buf_1 _2691_ (.A(_0514_),
    .X(_0629_));
 sg13g2_mux2_1 _2692_ (.A0(_0625_),
    .A1(_0623_),
    .S(_0607_),
    .X(_0630_));
 sg13g2_nor2_1 _2693_ (.A(net31),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_xnor2_1 _2694_ (.Y(_0632_),
    .A(net69),
    .B(_0631_));
 sg13g2_nor2_1 _2695_ (.A(_0394_),
    .B(_0632_),
    .Y(_0162_));
 sg13g2_nand3b_1 _2696_ (.B(_0624_),
    .C(net69),
    .Y(_0633_),
    .A_N(_1353_));
 sg13g2_nand3_1 _2697_ (.B(_1353_),
    .C(_0624_),
    .A(net69),
    .Y(_0634_));
 sg13g2_nand2b_1 _2698_ (.Y(_0635_),
    .B(_0607_),
    .A_N(_0622_));
 sg13g2_mux2_1 _2699_ (.A0(_0633_),
    .A1(_0634_),
    .S(_0635_),
    .X(_0636_));
 sg13g2_inv_2 _2700_ (.Y(_0637_),
    .A(net27));
 sg13g2_a21oi_1 _2701_ (.A1(_0545_),
    .A2(_0593_),
    .Y(_0638_),
    .B1(_0637_));
 sg13g2_nand2_1 _2702_ (.Y(_0639_),
    .A(_0604_),
    .B(_0638_));
 sg13g2_nor2b_1 _2703_ (.A(_1352_),
    .B_N(_0622_),
    .Y(_0640_));
 sg13g2_o21ai_1 _2704_ (.B1(_0640_),
    .Y(_0641_),
    .A1(net32),
    .A2(_0620_));
 sg13g2_or2_1 _2705_ (.X(_0642_),
    .B(_0641_),
    .A(_0639_));
 sg13g2_inv_1 _2706_ (.Y(_0643_),
    .A(_1351_));
 sg13g2_nor2_1 _2707_ (.A(_0969_),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_nand3_1 _2708_ (.B(_0642_),
    .C(_0644_),
    .A(_0636_),
    .Y(_0645_));
 sg13g2_nor3_1 _2709_ (.A(_0969_),
    .B(_1351_),
    .C(_0514_),
    .Y(_0646_));
 sg13g2_nand2b_1 _2710_ (.Y(_0647_),
    .B(_0646_),
    .A_N(_0636_));
 sg13g2_nor2_1 _2711_ (.A(_0639_),
    .B(_0641_),
    .Y(_0648_));
 sg13g2_a22oi_1 _2712_ (.Y(_0649_),
    .B1(_0646_),
    .B2(_0648_),
    .A2(_0644_),
    .A1(net33));
 sg13g2_nand3_1 _2713_ (.B(_0647_),
    .C(_0649_),
    .A(_0645_),
    .Y(_0163_));
 sg13g2_nand2b_1 _2714_ (.Y(_0650_),
    .B(_0596_),
    .A_N(_0594_));
 sg13g2_nor2_1 _2715_ (.A(_0556_),
    .B(_0650_),
    .Y(_0651_));
 sg13g2_a21oi_1 _2716_ (.A1(_0599_),
    .A2(_0600_),
    .Y(_0652_),
    .B1(_1343_));
 sg13g2_nand3b_1 _2717_ (.B(net68),
    .C(_1328_),
    .Y(_0653_),
    .A_N(_0622_));
 sg13g2_nor2b_1 _2718_ (.A(net74),
    .B_N(_0653_),
    .Y(_0654_));
 sg13g2_nand3_1 _2719_ (.B(_0599_),
    .C(_0600_),
    .A(_1343_),
    .Y(_0655_));
 sg13g2_nor2_1 _2720_ (.A(_1328_),
    .B(net68),
    .Y(_0656_));
 sg13g2_a221oi_1 _2721_ (.B2(_0655_),
    .C1(_0656_),
    .B1(_0654_),
    .A1(_0652_),
    .Y(_0657_),
    .A2(_0653_));
 sg13g2_inv_1 _2722_ (.Y(_0658_),
    .A(net69));
 sg13g2_nor3_1 _2723_ (.A(_0643_),
    .B(_0658_),
    .C(_0622_),
    .Y(_0659_));
 sg13g2_o21ai_1 _2724_ (.B1(_0659_),
    .Y(_0660_),
    .A1(_0651_),
    .A2(_0657_));
 sg13g2_nand3_1 _2725_ (.B(net69),
    .C(_1353_),
    .A(_1351_),
    .Y(_0661_));
 sg13g2_nor3_1 _2726_ (.A(net32),
    .B(_0621_),
    .C(_0661_),
    .Y(_0662_));
 sg13g2_nand2b_1 _2727_ (.Y(_0663_),
    .B(_0662_),
    .A_N(_0660_));
 sg13g2_or2_1 _2728_ (.X(_0664_),
    .B(_0622_),
    .A(_1353_));
 sg13g2_or4_1 _2729_ (.A(_0658_),
    .B(net32),
    .C(_0620_),
    .D(_0664_),
    .X(_0665_));
 sg13g2_a21o_1 _2730_ (.A2(_0665_),
    .A1(_0641_),
    .B1(_1351_),
    .X(_0666_));
 sg13g2_a221oi_1 _2731_ (.B2(_0666_),
    .C1(_0605_),
    .B1(_0663_),
    .A1(_0545_),
    .Y(_0667_),
    .A2(_0593_));
 sg13g2_nor2_2 _2732_ (.A(_0637_),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_xor2_1 _2733_ (.B(_0668_),
    .A(_0660_),
    .X(_0669_));
 sg13g2_o21ai_1 _2734_ (.B1(_1340_),
    .Y(_0670_),
    .A1(net33),
    .A2(_0669_));
 sg13g2_or3_1 _2735_ (.A(net72),
    .B(net31),
    .C(_0669_),
    .X(_0671_));
 sg13g2_a21oi_1 _2736_ (.A1(_0670_),
    .A2(_0671_),
    .Y(_0164_),
    .B1(_0451_));
 sg13g2_inv_1 _2737_ (.Y(_0672_),
    .A(\simon1.sound_gen_inst.tick_counter[14] ));
 sg13g2_nor2_1 _2738_ (.A(net49),
    .B(_0672_),
    .Y(_0673_));
 sg13g2_nor2_1 _2739_ (.A(_0970_),
    .B(\simon1.sound_gen_inst.tick_counter[14] ),
    .Y(_0674_));
 sg13g2_nand2_1 _2740_ (.Y(_0675_),
    .A(net72),
    .B(_0662_));
 sg13g2_nand3b_1 _2741_ (.B(_0596_),
    .C(_0659_),
    .Y(_0676_),
    .A_N(_0594_));
 sg13g2_o21ai_1 _2742_ (.B1(net72),
    .Y(_0677_),
    .A1(_0556_),
    .A2(_0676_));
 sg13g2_a21o_1 _2743_ (.A2(_0657_),
    .A1(_0659_),
    .B1(_0677_),
    .X(_0678_));
 sg13g2_or3_1 _2744_ (.A(_0613_),
    .B(_0621_),
    .C(_0661_),
    .X(_0679_));
 sg13g2_nand2b_1 _2745_ (.Y(_0680_),
    .B(_0679_),
    .A_N(_0678_));
 sg13g2_mux2_1 _2746_ (.A0(_0675_),
    .A1(_0680_),
    .S(_0668_),
    .X(_0681_));
 sg13g2_inv_1 _2747_ (.Y(_0682_),
    .A(_0663_));
 sg13g2_nor2_1 _2748_ (.A(net72),
    .B(_0660_),
    .Y(_0683_));
 sg13g2_a22oi_1 _2749_ (.Y(_0684_),
    .B1(_0668_),
    .B2(_0683_),
    .A2(_0682_),
    .A1(net72));
 sg13g2_a21oi_1 _2750_ (.A1(_0681_),
    .A2(_0684_),
    .Y(_0685_),
    .B1(net31));
 sg13g2_mux2_1 _2751_ (.A0(_0673_),
    .A1(_0674_),
    .S(_0685_),
    .X(_0165_));
 sg13g2_nand2_1 _2752_ (.Y(_0686_),
    .A(net27),
    .B(_0604_));
 sg13g2_a221oi_1 _2753_ (.B2(_0666_),
    .C1(_0686_),
    .B1(_0663_),
    .A1(_0545_),
    .Y(_0687_),
    .A2(_0593_));
 sg13g2_buf_1 _2754_ (.A(_0687_),
    .X(_0688_));
 sg13g2_nor3_1 _2755_ (.A(\simon1.sound_gen_inst.tick_counter[14] ),
    .B(_0679_),
    .C(_0678_),
    .Y(_0689_));
 sg13g2_nor3_1 _2756_ (.A(_0672_),
    .B(_0662_),
    .C(_0678_),
    .Y(_0690_));
 sg13g2_nor3_1 _2757_ (.A(_0672_),
    .B(net72),
    .C(_0660_),
    .Y(_0691_));
 sg13g2_nor4_2 _2758_ (.A(_0637_),
    .B(_0689_),
    .C(_0690_),
    .Y(_0692_),
    .D(_0691_));
 sg13g2_nor2_1 _2759_ (.A(_0688_),
    .B(_0692_),
    .Y(_0693_));
 sg13g2_nand3b_1 _2760_ (.B(net69),
    .C(_1351_),
    .Y(_0694_),
    .A_N(_0622_));
 sg13g2_nor4_2 _2761_ (.A(_1341_),
    .B(_0613_),
    .C(_0620_),
    .Y(_0695_),
    .D(_0694_));
 sg13g2_nor3_1 _2762_ (.A(net40),
    .B(_0693_),
    .C(_0695_),
    .Y(_0696_));
 sg13g2_xnor2_1 _2763_ (.Y(_0697_),
    .A(_1349_),
    .B(_0696_));
 sg13g2_nor2_1 _2764_ (.A(net44),
    .B(_0697_),
    .Y(_0166_));
 sg13g2_nor2_1 _2765_ (.A(net49),
    .B(_1368_),
    .Y(_0698_));
 sg13g2_inv_1 _2766_ (.Y(_0699_),
    .A(_1368_));
 sg13g2_nor2_1 _2767_ (.A(_0970_),
    .B(_0699_),
    .Y(_0700_));
 sg13g2_nand3_1 _2768_ (.B(\simon1.sound_gen_inst.tick_counter[14] ),
    .C(net72),
    .A(_1349_),
    .Y(_0701_));
 sg13g2_or3_1 _2769_ (.A(_0612_),
    .B(_0661_),
    .C(_0701_),
    .X(_0702_));
 sg13g2_buf_1 _2770_ (.A(_0702_),
    .X(_0703_));
 sg13g2_a21oi_1 _2771_ (.A1(_1328_),
    .A2(_0616_),
    .Y(_0704_),
    .B1(_0617_));
 sg13g2_nand2_1 _2772_ (.Y(_0705_),
    .A(net69),
    .B(_1353_));
 sg13g2_nor2_1 _2773_ (.A(_0704_),
    .B(_0705_),
    .Y(_0706_));
 sg13g2_a221oi_1 _2774_ (.B2(_0542_),
    .C1(_0706_),
    .B1(_0558_),
    .A1(_0614_),
    .Y(_0707_),
    .A2(_0615_));
 sg13g2_buf_2 _2775_ (.A(_0707_),
    .X(_0708_));
 sg13g2_nor2_1 _2776_ (.A(net26),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_xnor2_1 _2777_ (.Y(_0710_),
    .A(_1349_),
    .B(_0695_));
 sg13g2_o21ai_1 _2778_ (.B1(_0710_),
    .Y(_0711_),
    .A1(_0688_),
    .A2(_0692_));
 sg13g2_xnor2_1 _2779_ (.Y(_0712_),
    .A(_0709_),
    .B(_0711_));
 sg13g2_nand2_1 _2780_ (.Y(_0713_),
    .A(net34),
    .B(_0712_));
 sg13g2_mux2_1 _2781_ (.A0(_0698_),
    .A1(_0700_),
    .S(_0713_),
    .X(_0167_));
 sg13g2_or3_1 _2782_ (.A(_1368_),
    .B(net40),
    .C(_0709_),
    .X(_0714_));
 sg13g2_or2_1 _2783_ (.X(_0715_),
    .B(_0701_),
    .A(_0694_));
 sg13g2_buf_1 _2784_ (.A(_0715_),
    .X(_0716_));
 sg13g2_or3_1 _2785_ (.A(net32),
    .B(net21),
    .C(_0716_),
    .X(_0717_));
 sg13g2_or4_1 _2786_ (.A(_0699_),
    .B(_0513_),
    .C(_0709_),
    .D(_0717_),
    .X(_0718_));
 sg13g2_o21ai_1 _2787_ (.B1(_0718_),
    .Y(_0719_),
    .A1(_0711_),
    .A2(_0714_));
 sg13g2_xnor2_1 _2788_ (.Y(_0720_),
    .A(\simon1.sound_gen_inst.tick_counter[17] ),
    .B(_0719_));
 sg13g2_nor2_1 _2789_ (.A(net44),
    .B(_0720_),
    .Y(_0168_));
 sg13g2_nand2_1 _2790_ (.Y(_0721_),
    .A(\simon1.sound_gen_inst.tick_counter[17] ),
    .B(_1368_));
 sg13g2_or2_1 _2791_ (.X(_0722_),
    .B(_0721_),
    .A(net26));
 sg13g2_or2_1 _2792_ (.X(_0723_),
    .B(_0722_),
    .A(_0708_));
 sg13g2_xor2_1 _2793_ (.B(_0695_),
    .A(_1349_),
    .X(_0724_));
 sg13g2_a22oi_1 _2794_ (.Y(_0725_),
    .B1(_0558_),
    .B2(_0542_),
    .A2(_0615_),
    .A1(_0614_));
 sg13g2_or2_1 _2795_ (.X(_0726_),
    .B(_0705_),
    .A(_0704_));
 sg13g2_buf_1 _2796_ (.A(_0726_),
    .X(_0727_));
 sg13g2_nand2_1 _2797_ (.Y(_0728_),
    .A(_0725_),
    .B(_0727_));
 sg13g2_or2_1 _2798_ (.X(_0729_),
    .B(_0721_),
    .A(_0716_));
 sg13g2_nor2_1 _2799_ (.A(net26),
    .B(_0729_),
    .Y(_0730_));
 sg13g2_nor3_1 _2800_ (.A(_0699_),
    .B(net26),
    .C(_0708_),
    .Y(_0731_));
 sg13g2_nand2_1 _2801_ (.Y(_0732_),
    .A(_0699_),
    .B(_0727_));
 sg13g2_nand2_1 _2802_ (.Y(_0733_),
    .A(_0699_),
    .B(net26));
 sg13g2_o21ai_1 _2803_ (.B1(_0733_),
    .Y(_0734_),
    .A1(_0544_),
    .A2(_0732_));
 sg13g2_a221oi_1 _2804_ (.B2(_0717_),
    .C1(_0734_),
    .B1(_0731_),
    .A1(_0728_),
    .Y(_0735_),
    .A2(_0730_));
 sg13g2_nand2b_1 _2805_ (.Y(_0736_),
    .B(_0730_),
    .A_N(_0708_));
 sg13g2_and2_1 _2806_ (.A(\simon1.sound_gen_inst.tick_counter[17] ),
    .B(_0736_),
    .X(_0737_));
 sg13g2_nor3_2 _2807_ (.A(_0724_),
    .B(_0735_),
    .C(_0737_),
    .Y(_0738_));
 sg13g2_o21ai_1 _2808_ (.B1(_0738_),
    .Y(_0739_),
    .A1(_0688_),
    .A2(_0692_));
 sg13g2_xnor2_1 _2809_ (.Y(_0740_),
    .A(_0723_),
    .B(_0739_));
 sg13g2_o21ai_1 _2810_ (.B1(net64),
    .Y(_0741_),
    .A1(net31),
    .A2(_0740_));
 sg13g2_or3_1 _2811_ (.A(_1367_),
    .B(net31),
    .C(_0740_),
    .X(_0742_));
 sg13g2_a21oi_1 _2812_ (.A1(_0741_),
    .A2(_0742_),
    .Y(_0169_),
    .B1(net42));
 sg13g2_nand3b_1 _2813_ (.B(_1337_),
    .C(_0723_),
    .Y(_0743_),
    .A_N(net64));
 sg13g2_nor3_1 _2814_ (.A(net32),
    .B(net21),
    .C(_0729_),
    .Y(_0744_));
 sg13g2_nand4_1 _2815_ (.B(_1337_),
    .C(_0736_),
    .A(net64),
    .Y(_0745_),
    .D(_0744_));
 sg13g2_o21ai_1 _2816_ (.B1(_0745_),
    .Y(_0746_),
    .A1(_0739_),
    .A2(_0743_));
 sg13g2_xnor2_1 _2817_ (.Y(_0747_),
    .A(_1375_),
    .B(_0746_));
 sg13g2_nor2_1 _2818_ (.A(net44),
    .B(_0747_),
    .Y(_0170_));
 sg13g2_nand2_1 _2819_ (.Y(_0748_),
    .A(\simon1.sound_gen_inst.tick_counter[0] ),
    .B(\simon1.sound_freq[0] ));
 sg13g2_xnor2_1 _2820_ (.Y(_0749_),
    .A(\simon1.sound_freq[1] ),
    .B(\simon1.sound_gen_inst.tick_counter[1] ));
 sg13g2_xnor2_1 _2821_ (.Y(_0750_),
    .A(_0748_),
    .B(_0749_));
 sg13g2_nor2_1 _2822_ (.A(net48),
    .B(_0750_),
    .Y(_0171_));
 sg13g2_or2_1 _2823_ (.X(_0751_),
    .B(_0692_),
    .A(_0688_));
 sg13g2_buf_2 _2824_ (.A(_0751_),
    .X(_0752_));
 sg13g2_or2_1 _2825_ (.X(_0753_),
    .B(net64),
    .A(_1375_));
 sg13g2_nand2_1 _2826_ (.Y(_0754_),
    .A(_1375_),
    .B(net64));
 sg13g2_nor2b_1 _2827_ (.A(_1375_),
    .B_N(net64),
    .Y(_0755_));
 sg13g2_o21ai_1 _2828_ (.B1(_0755_),
    .Y(_0756_),
    .A1(_0694_),
    .A2(_0701_));
 sg13g2_o21ai_1 _2829_ (.B1(_0756_),
    .Y(_0757_),
    .A1(_0716_),
    .A2(_0754_));
 sg13g2_nor3_1 _2830_ (.A(_0703_),
    .B(_0721_),
    .C(_0757_),
    .Y(_0758_));
 sg13g2_nor4_1 _2831_ (.A(_0703_),
    .B(_0727_),
    .C(_0721_),
    .D(_0757_),
    .Y(_0759_));
 sg13g2_a221oi_1 _2832_ (.B2(_0544_),
    .C1(_0759_),
    .B1(_0758_),
    .A1(_0753_),
    .Y(_0760_),
    .A2(_0722_));
 sg13g2_nand3_1 _2833_ (.B(_0725_),
    .C(_0727_),
    .A(_0753_),
    .Y(_0761_));
 sg13g2_and4_1 _2834_ (.A(_0752_),
    .B(_0738_),
    .C(_0760_),
    .D(_0761_),
    .X(_0762_));
 sg13g2_inv_1 _2835_ (.Y(_0763_),
    .A(_1374_));
 sg13g2_nor2_1 _2836_ (.A(_0763_),
    .B(_0706_),
    .Y(_0764_));
 sg13g2_nor3_1 _2837_ (.A(_0612_),
    .B(_0661_),
    .C(_0701_),
    .Y(_0765_));
 sg13g2_and4_1 _2838_ (.A(_1375_),
    .B(net64),
    .C(\simon1.sound_gen_inst.tick_counter[17] ),
    .D(_1368_),
    .X(_0766_));
 sg13g2_buf_1 _2839_ (.A(_0766_),
    .X(_0767_));
 sg13g2_a21oi_1 _2840_ (.A1(_0765_),
    .A2(_0767_),
    .Y(_0768_),
    .B1(_0763_));
 sg13g2_a21oi_1 _2841_ (.A1(_0725_),
    .A2(_0764_),
    .Y(_0769_),
    .B1(_0768_));
 sg13g2_or4_1 _2842_ (.A(_1374_),
    .B(_0708_),
    .C(_0722_),
    .D(_0754_),
    .X(_0770_));
 sg13g2_nand2_1 _2843_ (.Y(_0771_),
    .A(_0769_),
    .B(_0770_));
 sg13g2_xnor2_1 _2844_ (.Y(_0772_),
    .A(_0762_),
    .B(_0771_));
 sg13g2_nand3_1 _2845_ (.B(_1374_),
    .C(net33),
    .A(net62),
    .Y(_0773_));
 sg13g2_o21ai_1 _2846_ (.B1(_0773_),
    .Y(_0172_),
    .A1(_1339_),
    .A2(_0772_));
 sg13g2_nor4_1 _2847_ (.A(_0763_),
    .B(_0716_),
    .C(_0721_),
    .D(_0754_),
    .Y(_0774_));
 sg13g2_o21ai_1 _2848_ (.B1(_0774_),
    .Y(_0775_),
    .A1(_0651_),
    .A2(_0657_));
 sg13g2_nand4_1 _2849_ (.B(_0761_),
    .C(_0769_),
    .A(_0760_),
    .Y(_0776_),
    .D(_0770_));
 sg13g2_nor4_1 _2850_ (.A(_0724_),
    .B(_0735_),
    .C(_0737_),
    .D(_0776_),
    .Y(_0777_));
 sg13g2_o21ai_1 _2851_ (.B1(_0777_),
    .Y(_0778_),
    .A1(_0688_),
    .A2(_0692_));
 sg13g2_xnor2_1 _2852_ (.Y(_0779_),
    .A(_0775_),
    .B(_0778_));
 sg13g2_o21ai_1 _2853_ (.B1(_1373_),
    .Y(_0780_),
    .A1(net31),
    .A2(_0779_));
 sg13g2_or3_1 _2854_ (.A(_1373_),
    .B(net31),
    .C(_0779_),
    .X(_0781_));
 sg13g2_a21oi_1 _2855_ (.A1(_0780_),
    .A2(_0781_),
    .Y(_0173_),
    .B1(net42));
 sg13g2_xnor2_1 _2856_ (.Y(_0782_),
    .A(_1373_),
    .B(_0775_));
 sg13g2_nand3_1 _2857_ (.B(_1374_),
    .C(_0767_),
    .A(_1373_),
    .Y(_0783_));
 sg13g2_nor3_2 _2858_ (.A(net21),
    .B(net26),
    .C(_0783_),
    .Y(_0784_));
 sg13g2_o21ai_1 _2859_ (.B1(_0784_),
    .Y(_0785_),
    .A1(_0778_),
    .A2(_0782_));
 sg13g2_or4_1 _2860_ (.A(net40),
    .B(_0778_),
    .C(_0784_),
    .D(_0782_),
    .X(_0786_));
 sg13g2_nand3_1 _2861_ (.B(_0785_),
    .C(_0786_),
    .A(_1372_),
    .Y(_0787_));
 sg13g2_a21o_1 _2862_ (.A2(_0786_),
    .A1(_0785_),
    .B1(_1372_),
    .X(_0788_));
 sg13g2_a21oi_1 _2863_ (.A1(_0787_),
    .A2(_0788_),
    .Y(_0174_),
    .B1(net42));
 sg13g2_or2_1 _2864_ (.X(_0789_),
    .B(_0737_),
    .A(_0735_));
 sg13g2_nand4_1 _2865_ (.B(_1373_),
    .C(_1374_),
    .A(_1372_),
    .Y(_0790_),
    .D(_0767_));
 sg13g2_nor2_1 _2866_ (.A(_0716_),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_nand2b_1 _2867_ (.Y(_0792_),
    .B(_0791_),
    .A_N(_0612_));
 sg13g2_or2_1 _2868_ (.X(_0793_),
    .B(_0792_),
    .A(_0620_));
 sg13g2_buf_2 _2869_ (.A(_0793_),
    .X(_0794_));
 sg13g2_xor2_1 _2870_ (.B(_0784_),
    .A(_1372_),
    .X(_0795_));
 sg13g2_nor3_1 _2871_ (.A(_0776_),
    .B(_0782_),
    .C(_0795_),
    .Y(_0796_));
 sg13g2_nand3b_1 _2872_ (.B(_0794_),
    .C(_0796_),
    .Y(_0797_),
    .A_N(_0789_));
 sg13g2_nor2_1 _2873_ (.A(net21),
    .B(_0792_),
    .Y(_0798_));
 sg13g2_and4_1 _2874_ (.A(_1372_),
    .B(_1373_),
    .C(_1374_),
    .D(_0767_),
    .X(_0799_));
 sg13g2_nand2_1 _2875_ (.Y(_0800_),
    .A(_0709_),
    .B(_0799_));
 sg13g2_nand2_1 _2876_ (.Y(_0801_),
    .A(_0798_),
    .B(_0800_));
 sg13g2_o21ai_1 _2877_ (.B1(_0801_),
    .Y(_0802_),
    .A1(_0711_),
    .A2(_0797_));
 sg13g2_a21o_1 _2878_ (.A2(_0802_),
    .A1(net34),
    .B1(_1363_),
    .X(_0803_));
 sg13g2_nand3_1 _2879_ (.B(net34),
    .C(_0802_),
    .A(_1363_),
    .Y(_0804_));
 sg13g2_a21oi_1 _2880_ (.A1(_0803_),
    .A2(_0804_),
    .Y(_0175_),
    .B1(net42));
 sg13g2_and2_1 _2881_ (.A(net79),
    .B(_1370_),
    .X(_0805_));
 sg13g2_nor2_1 _2882_ (.A(net61),
    .B(_1370_),
    .Y(_0806_));
 sg13g2_nand2b_1 _2883_ (.Y(_0807_),
    .B(_0796_),
    .A_N(_0739_));
 sg13g2_nand3_1 _2884_ (.B(_1337_),
    .C(_0794_),
    .A(_1363_),
    .Y(_0808_));
 sg13g2_nor3_2 _2885_ (.A(net26),
    .B(_0708_),
    .C(_0790_),
    .Y(_0809_));
 sg13g2_nand4_1 _2886_ (.B(_1337_),
    .C(_0794_),
    .A(_1362_),
    .Y(_0810_),
    .D(_0809_));
 sg13g2_o21ai_1 _2887_ (.B1(_0810_),
    .Y(_0811_),
    .A1(_0807_),
    .A2(_0808_));
 sg13g2_mux2_1 _2888_ (.A0(_0805_),
    .A1(_0806_),
    .S(_0811_),
    .X(_0176_));
 sg13g2_nand3_1 _2889_ (.B(_1362_),
    .C(_0791_),
    .A(_1370_),
    .Y(_0812_));
 sg13g2_nor3_1 _2890_ (.A(net32),
    .B(net21),
    .C(_0812_),
    .Y(_0813_));
 sg13g2_xnor2_1 _2891_ (.Y(_0814_),
    .A(\simon1.sound_gen_inst.tick_counter[25] ),
    .B(_0813_));
 sg13g2_nor4_1 _2892_ (.A(_1370_),
    .B(_1363_),
    .C(_0794_),
    .D(_0809_),
    .Y(_0815_));
 sg13g2_nand4_1 _2893_ (.B(_1362_),
    .C(_0765_),
    .A(_1370_),
    .Y(_0816_),
    .D(_0799_));
 sg13g2_nor3_1 _2894_ (.A(_0708_),
    .B(_0794_),
    .C(_0816_),
    .Y(_0817_));
 sg13g2_nor3_1 _2895_ (.A(_1370_),
    .B(_1362_),
    .C(_0798_),
    .Y(_0818_));
 sg13g2_or3_1 _2896_ (.A(_0815_),
    .B(_0817_),
    .C(_0818_),
    .X(_0819_));
 sg13g2_nand4_1 _2897_ (.B(_0738_),
    .C(_0796_),
    .A(_0752_),
    .Y(_0820_),
    .D(_0819_));
 sg13g2_xnor2_1 _2898_ (.Y(_0821_),
    .A(_0814_),
    .B(_0820_));
 sg13g2_nand3_1 _2899_ (.B(\simon1.sound_gen_inst.tick_counter[25] ),
    .C(net33),
    .A(net62),
    .Y(_0822_));
 sg13g2_o21ai_1 _2900_ (.B1(_0822_),
    .Y(_0177_),
    .A1(_1339_),
    .A2(_0821_));
 sg13g2_inv_1 _2901_ (.Y(_0823_),
    .A(\simon1.sound_gen_inst.tick_counter[26] ));
 sg13g2_nor2_1 _2902_ (.A(_0782_),
    .B(_0795_),
    .Y(_0824_));
 sg13g2_nor2b_1 _2903_ (.A(_0776_),
    .B_N(_0814_),
    .Y(_0825_));
 sg13g2_nand4_1 _2904_ (.B(_0824_),
    .C(_0819_),
    .A(_0738_),
    .Y(_0826_),
    .D(_0825_));
 sg13g2_nand3_1 _2905_ (.B(_1370_),
    .C(_1362_),
    .A(\simon1.sound_gen_inst.tick_counter[25] ),
    .Y(_0827_));
 sg13g2_buf_1 _2906_ (.A(_0827_),
    .X(_0828_));
 sg13g2_nor4_2 _2907_ (.A(net26),
    .B(_0708_),
    .C(_0790_),
    .Y(_0829_),
    .D(_0828_));
 sg13g2_nor4_1 _2908_ (.A(net40),
    .B(_0693_),
    .C(_0826_),
    .D(_0829_),
    .Y(_0830_));
 sg13g2_and4_1 _2909_ (.A(_0738_),
    .B(_0824_),
    .C(_0819_),
    .D(_0825_),
    .X(_0831_));
 sg13g2_buf_1 _2910_ (.A(_0831_),
    .X(_0832_));
 sg13g2_inv_1 _2911_ (.Y(_0833_),
    .A(_0829_));
 sg13g2_a21oi_1 _2912_ (.A1(_0752_),
    .A2(_0832_),
    .Y(_0834_),
    .B1(_0833_));
 sg13g2_or3_1 _2913_ (.A(_0823_),
    .B(_0830_),
    .C(_0834_),
    .X(_0835_));
 sg13g2_o21ai_1 _2914_ (.B1(_0823_),
    .Y(_0836_),
    .A1(_0830_),
    .A2(_0834_));
 sg13g2_a21oi_1 _2915_ (.A1(_0835_),
    .A2(_0836_),
    .Y(_0178_),
    .B1(net42));
 sg13g2_nor2_1 _2916_ (.A(net61),
    .B(_1364_),
    .Y(_0837_));
 sg13g2_and2_1 _2917_ (.A(net79),
    .B(_1364_),
    .X(_0838_));
 sg13g2_nor3_1 _2918_ (.A(_0823_),
    .B(_0794_),
    .C(_0828_),
    .Y(_0839_));
 sg13g2_nand3_1 _2919_ (.B(_0809_),
    .C(_0832_),
    .A(_0752_),
    .Y(_0840_));
 sg13g2_o21ai_1 _2920_ (.B1(\simon1.sound_gen_inst.tick_counter[26] ),
    .Y(_0841_),
    .A1(net21),
    .A2(_0792_));
 sg13g2_mux2_1 _2921_ (.A0(\simon1.sound_gen_inst.tick_counter[26] ),
    .A1(_0841_),
    .S(_0829_),
    .X(_0842_));
 sg13g2_nor2_1 _2922_ (.A(net40),
    .B(_0842_),
    .Y(_0843_));
 sg13g2_nor2_1 _2923_ (.A(_0693_),
    .B(_0826_),
    .Y(_0844_));
 sg13g2_a22oi_1 _2924_ (.Y(_0845_),
    .B1(_0843_),
    .B2(_0844_),
    .A2(_0840_),
    .A1(_0839_));
 sg13g2_mux2_1 _2925_ (.A0(_0837_),
    .A1(_0838_),
    .S(_0845_),
    .X(_0179_));
 sg13g2_nor2_1 _2926_ (.A(_1364_),
    .B(_0842_),
    .Y(_0846_));
 sg13g2_nand3_1 _2927_ (.B(_0728_),
    .C(_0799_),
    .A(_0765_),
    .Y(_0847_));
 sg13g2_and2_1 _2928_ (.A(_1364_),
    .B(\simon1.sound_gen_inst.tick_counter[26] ),
    .X(_0848_));
 sg13g2_nand2b_1 _2929_ (.Y(_0849_),
    .B(_0848_),
    .A_N(_0828_));
 sg13g2_nor2_1 _2930_ (.A(_0847_),
    .B(_0849_),
    .Y(_0850_));
 sg13g2_nand3_1 _2931_ (.B(_0829_),
    .C(_0848_),
    .A(_0798_),
    .Y(_0851_));
 sg13g2_o21ai_1 _2932_ (.B1(_0851_),
    .Y(_0852_),
    .A1(_1364_),
    .A2(_0842_));
 sg13g2_nand3_1 _2933_ (.B(_0832_),
    .C(_0852_),
    .A(_0752_),
    .Y(_0853_));
 sg13g2_nand2_1 _2934_ (.Y(_0854_),
    .A(_0968_),
    .B(\simon1.sound_gen_inst.tick_counter[28] ));
 sg13g2_a221oi_1 _2935_ (.B2(_0853_),
    .C1(_0854_),
    .B1(_0850_),
    .A1(_0844_),
    .Y(_0855_),
    .A2(_0846_));
 sg13g2_nor3_1 _2936_ (.A(_0969_),
    .B(\simon1.sound_gen_inst.tick_counter[28] ),
    .C(net40),
    .Y(_0856_));
 sg13g2_nand3_1 _2937_ (.B(_0853_),
    .C(_0856_),
    .A(_0850_),
    .Y(_0857_));
 sg13g2_inv_1 _2938_ (.Y(_0858_),
    .A(\simon1.sound_gen_inst.tick_counter[28] ));
 sg13g2_nor2_1 _2939_ (.A(_0969_),
    .B(_0858_),
    .Y(_0859_));
 sg13g2_nor4_1 _2940_ (.A(_1364_),
    .B(_0693_),
    .C(_0826_),
    .D(_0842_),
    .Y(_0860_));
 sg13g2_a22oi_1 _2941_ (.Y(_0861_),
    .B1(_0856_),
    .B2(_0860_),
    .A2(_0859_),
    .A1(net33));
 sg13g2_nand3b_1 _2942_ (.B(_0857_),
    .C(_0861_),
    .Y(_0180_),
    .A_N(_0855_));
 sg13g2_nand2_1 _2943_ (.Y(_0862_),
    .A(\simon1.sound_gen_inst.tick_counter[28] ),
    .B(_0848_));
 sg13g2_nor4_1 _2944_ (.A(_0717_),
    .B(_0790_),
    .C(_0828_),
    .D(_0862_),
    .Y(_0863_));
 sg13g2_xnor2_1 _2945_ (.Y(_0864_),
    .A(\simon1.sound_gen_inst.tick_counter[29] ),
    .B(_0863_));
 sg13g2_nor4_1 _2946_ (.A(_0794_),
    .B(_0800_),
    .C(_0828_),
    .D(_0862_),
    .Y(_0865_));
 sg13g2_a21o_1 _2947_ (.A2(_0846_),
    .A1(_0858_),
    .B1(_0865_),
    .X(_0866_));
 sg13g2_nand3_1 _2948_ (.B(_0832_),
    .C(_0866_),
    .A(_0752_),
    .Y(_0867_));
 sg13g2_xnor2_1 _2949_ (.Y(_0868_),
    .A(_0864_),
    .B(_0867_));
 sg13g2_nand3_1 _2950_ (.B(\simon1.sound_gen_inst.tick_counter[29] ),
    .C(net33),
    .A(net79),
    .Y(_0869_));
 sg13g2_o21ai_1 _2951_ (.B1(_0869_),
    .Y(_0181_),
    .A1(_1339_),
    .A2(_0868_));
 sg13g2_nor2_1 _2952_ (.A(_0533_),
    .B(_0534_),
    .Y(_0870_));
 sg13g2_xor2_1 _2953_ (.B(_0536_),
    .A(_0870_),
    .X(_0871_));
 sg13g2_nor2_1 _2954_ (.A(net48),
    .B(_0871_),
    .Y(_0182_));
 sg13g2_and2_1 _2955_ (.A(net79),
    .B(\simon1.sound_gen_inst.tick_counter[30] ),
    .X(_0872_));
 sg13g2_nor2_1 _2956_ (.A(_0969_),
    .B(\simon1.sound_gen_inst.tick_counter[30] ),
    .Y(_0873_));
 sg13g2_nor2_1 _2957_ (.A(_0828_),
    .B(_0862_),
    .Y(_0874_));
 sg13g2_nand2_1 _2958_ (.Y(_0875_),
    .A(\simon1.sound_gen_inst.tick_counter[29] ),
    .B(_0874_));
 sg13g2_nor2_1 _2959_ (.A(_0847_),
    .B(_0875_),
    .Y(_0876_));
 sg13g2_nor2_1 _2960_ (.A(net40),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_and4_1 _2961_ (.A(_0752_),
    .B(_0832_),
    .C(_0864_),
    .D(_0866_),
    .X(_0878_));
 sg13g2_mux2_1 _2962_ (.A0(_0876_),
    .A1(_0877_),
    .S(_0878_),
    .X(_0879_));
 sg13g2_mux2_1 _2963_ (.A0(_0872_),
    .A1(_0873_),
    .S(_0879_),
    .X(_0183_));
 sg13g2_nor2_1 _2964_ (.A(net61),
    .B(\simon1.sound_gen_inst.tick_counter[31] ),
    .Y(_0880_));
 sg13g2_and2_1 _2965_ (.A(_0968_),
    .B(\simon1.sound_gen_inst.tick_counter[31] ),
    .X(_0881_));
 sg13g2_inv_1 _2966_ (.Y(_0882_),
    .A(_0875_));
 sg13g2_nand4_1 _2967_ (.B(_1337_),
    .C(_0798_),
    .A(\simon1.sound_gen_inst.tick_counter[30] ),
    .Y(_0883_),
    .D(_0882_));
 sg13g2_nand4_1 _2968_ (.B(_0794_),
    .C(_0809_),
    .A(\simon1.sound_gen_inst.tick_counter[30] ),
    .Y(_0884_),
    .D(_0882_));
 sg13g2_o21ai_1 _2969_ (.B1(_0884_),
    .Y(_0885_),
    .A1(\simon1.sound_gen_inst.tick_counter[30] ),
    .A2(_0876_));
 sg13g2_nand4_1 _2970_ (.B(_0864_),
    .C(_0866_),
    .A(_1337_),
    .Y(_0886_),
    .D(_0885_));
 sg13g2_mux2_1 _2971_ (.A0(_0883_),
    .A1(_0886_),
    .S(_0844_),
    .X(_0887_));
 sg13g2_mux2_1 _2972_ (.A0(_0880_),
    .A1(_0881_),
    .S(_0887_),
    .X(_0184_));
 sg13g2_xnor2_1 _2973_ (.Y(_0888_),
    .A(net27),
    .B(_0575_));
 sg13g2_o21ai_1 _2974_ (.B1(_0231_),
    .Y(_0889_),
    .A1(_1346_),
    .A2(net34));
 sg13g2_a21oi_1 _2975_ (.A1(net34),
    .A2(_0888_),
    .Y(_0185_),
    .B1(_0889_));
 sg13g2_nand2_1 _2976_ (.Y(_0890_),
    .A(_1357_),
    .B(net33));
 sg13g2_nor2_1 _2977_ (.A(_0637_),
    .B(_0575_),
    .Y(_0891_));
 sg13g2_xor2_1 _2978_ (.B(_0891_),
    .A(_0572_),
    .X(_0892_));
 sg13g2_nand2_1 _2979_ (.Y(_0893_),
    .A(net34),
    .B(_0892_));
 sg13g2_a21oi_1 _2980_ (.A1(_0890_),
    .A2(_0893_),
    .Y(_0186_),
    .B1(net49));
 sg13g2_o21ai_1 _2981_ (.B1(net27),
    .Y(_0894_),
    .A1(_0572_),
    .A2(_0575_));
 sg13g2_xnor2_1 _2982_ (.Y(_0895_),
    .A(_0546_),
    .B(_0556_));
 sg13g2_xnor2_1 _2983_ (.Y(_0896_),
    .A(_0894_),
    .B(_0895_));
 sg13g2_nor2_1 _2984_ (.A(_0629_),
    .B(_0896_),
    .Y(_0897_));
 sg13g2_xnor2_1 _2985_ (.Y(_0898_),
    .A(_1358_),
    .B(_0897_));
 sg13g2_nor2_1 _2986_ (.A(net48),
    .B(_0898_),
    .Y(_0187_));
 sg13g2_nor3_1 _2987_ (.A(_0572_),
    .B(_0575_),
    .C(_0561_),
    .Y(_0899_));
 sg13g2_a221oi_1 _2988_ (.B2(_0580_),
    .C1(_1325_),
    .B1(_0577_),
    .A1(_0572_),
    .Y(_0900_),
    .A2(_0561_));
 sg13g2_o21ai_1 _2989_ (.B1(net27),
    .Y(_0901_),
    .A1(_0899_),
    .A2(_0900_));
 sg13g2_nor2_1 _2990_ (.A(net27),
    .B(_0556_),
    .Y(_0902_));
 sg13g2_o21ai_1 _2991_ (.B1(_0902_),
    .Y(_0903_),
    .A1(_1325_),
    .A2(net65));
 sg13g2_o21ai_1 _2992_ (.B1(_0595_),
    .Y(_0904_),
    .A1(_0572_),
    .A2(_0575_));
 sg13g2_a21o_1 _2993_ (.A2(_0904_),
    .A1(net27),
    .B1(_0566_),
    .X(_0905_));
 sg13g2_nand3_1 _2994_ (.B(_0903_),
    .C(_0905_),
    .A(_0901_),
    .Y(_0906_));
 sg13g2_xnor2_1 _2995_ (.Y(_0907_),
    .A(net73),
    .B(_0906_));
 sg13g2_nor2_1 _2996_ (.A(net31),
    .B(_0907_),
    .Y(_0908_));
 sg13g2_xnor2_1 _2997_ (.Y(_0909_),
    .A(_1356_),
    .B(_0908_));
 sg13g2_nor2_1 _2998_ (.A(_0971_),
    .B(_0909_),
    .Y(_0188_));
 sg13g2_nand2_1 _2999_ (.Y(_0910_),
    .A(_1342_),
    .B(_0515_));
 sg13g2_nand2_1 _3000_ (.Y(_0911_),
    .A(_1383_),
    .B(_0593_));
 sg13g2_or3_1 _3001_ (.A(_0570_),
    .B(_0576_),
    .C(_0582_),
    .X(_0912_));
 sg13g2_o21ai_1 _3002_ (.B1(_0592_),
    .Y(_0913_),
    .A1(_0637_),
    .A2(_0912_));
 sg13g2_nand3_1 _3003_ (.B(_0911_),
    .C(_0913_),
    .A(_1338_),
    .Y(_0914_));
 sg13g2_a21oi_1 _3004_ (.A1(_0910_),
    .A2(_0914_),
    .Y(_0189_),
    .B1(_0321_));
 sg13g2_xnor2_1 _3005_ (.Y(_0915_),
    .A(_1329_),
    .B(_0544_));
 sg13g2_xnor2_1 _3006_ (.Y(_0916_),
    .A(_0911_),
    .B(_0915_));
 sg13g2_nor2_1 _3007_ (.A(_0629_),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_xnor2_1 _3008_ (.Y(_0918_),
    .A(net70),
    .B(_0917_));
 sg13g2_nor2_1 _3009_ (.A(_0971_),
    .B(_0918_),
    .Y(_0190_));
 sg13g2_nand2_1 _3010_ (.Y(_0919_),
    .A(_1354_),
    .B(_0515_));
 sg13g2_nor2_1 _3011_ (.A(_0604_),
    .B(_0638_),
    .Y(_0920_));
 sg13g2_o21ai_1 _3012_ (.B1(_1338_),
    .Y(_0921_),
    .A1(_0607_),
    .A2(_0920_));
 sg13g2_a21oi_1 _3013_ (.A1(_0919_),
    .A2(_0921_),
    .Y(_0191_),
    .B1(_0321_));
 sg13g2_xnor2_1 _3014_ (.Y(_0922_),
    .A(net86),
    .B(_0941_));
 sg13g2_nor3_1 _3015_ (.A(net87),
    .B(_0940_),
    .C(_0922_),
    .Y(_0923_));
 sg13g2_a21oi_1 _3016_ (.A1(net78),
    .A2(_0923_),
    .Y(_0924_),
    .B1(_0951_));
 sg13g2_xnor2_1 _3017_ (.Y(_0925_),
    .A(net87),
    .B(_0940_));
 sg13g2_nor4_1 _3018_ (.A(_0939_),
    .B(_0941_),
    .C(_1439_),
    .D(_0925_),
    .Y(_0926_));
 sg13g2_nor3_1 _3019_ (.A(net49),
    .B(_0924_),
    .C(_0926_),
    .Y(_0211_));
 sg13g2_a21oi_1 _3020_ (.A1(_1062_),
    .A2(_1057_),
    .Y(_0927_),
    .B1(_0948_));
 sg13g2_nor2_1 _3021_ (.A(_0940_),
    .B(_0941_),
    .Y(_0928_));
 sg13g2_nand2_1 _3022_ (.Y(_0929_),
    .A(_0938_),
    .B(net86));
 sg13g2_nand3_1 _3023_ (.B(_0928_),
    .C(_0929_),
    .A(net78),
    .Y(_0930_));
 sg13g2_nor2_1 _3024_ (.A(_0938_),
    .B(net86),
    .Y(_0931_));
 sg13g2_a21oi_1 _3025_ (.A1(_0948_),
    .A2(_0930_),
    .Y(_0932_),
    .B1(_0931_));
 sg13g2_nor3_1 _3026_ (.A(net49),
    .B(_0927_),
    .C(_0932_),
    .Y(_0212_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _3029__91 (.L_HI(net91));
 sg13g2_buf_1 _3029_ (.A(net91),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3030_ (.A(net92),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3031_ (.A(net93),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3032_ (.A(net94),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3033_ (.A(net95),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3034_ (.A(net96),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3035_ (.A(net97),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3036_ (.A(net88),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3037_ (.A(net89),
    .X(uio_out[7]));
 sg13g2_buf_1 _3038_ (.A(\simon1.sound ),
    .X(net13));
 sg13g2_buf_1 _3039_ (.A(net90),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \simon1.button_released$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net98),
    .D(_0036_),
    .Q_N(_1595_),
    .Q(\simon1.button_released ));
 sg13g2_dfrbp_1 \simon1.led[0]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net99),
    .D(_0037_),
    .Q_N(_1594_),
    .Q(net9));
 sg13g2_dfrbp_1 \simon1.led[1]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net100),
    .D(_0038_),
    .Q_N(_1593_),
    .Q(net10));
 sg13g2_dfrbp_1 \simon1.led[2]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net101),
    .D(_0039_),
    .Q_N(_1592_),
    .Q(net11));
 sg13g2_dfrbp_1 \simon1.led[3]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net102),
    .D(_0040_),
    .Q_N(_1591_),
    .Q(net12));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[0]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net103),
    .D(_0041_),
    .Q_N(_1590_),
    .Q(\simon1.lfsr_capture[0] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[10]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net104),
    .D(_0042_),
    .Q_N(_1589_),
    .Q(\simon1.lfsr_capture[10] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[11]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net105),
    .D(_0043_),
    .Q_N(_1588_),
    .Q(\simon1.lfsr_capture[11] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[12]$_SDFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net106),
    .D(_0044_),
    .Q_N(_1587_),
    .Q(\simon1.lfsr_capture[12] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[13]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net107),
    .D(_0045_),
    .Q_N(_1586_),
    .Q(\simon1.lfsr_capture[13] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[14]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net108),
    .D(_0046_),
    .Q_N(_1585_),
    .Q(\simon1.lfsr_capture[14] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[15]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net109),
    .D(_0047_),
    .Q_N(_1584_),
    .Q(\simon1.lfsr_capture[15] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[16]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net110),
    .D(_0048_),
    .Q_N(_1583_),
    .Q(\simon1.lfsr_capture[16] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[17]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net111),
    .D(_0049_),
    .Q_N(_1582_),
    .Q(\simon1.lfsr_capture[17] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[18]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net112),
    .D(_0050_),
    .Q_N(_1581_),
    .Q(\simon1.lfsr_capture[18] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[19]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net113),
    .D(_0051_),
    .Q_N(_1580_),
    .Q(\simon1.lfsr_capture[19] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[1]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net114),
    .D(_0052_),
    .Q_N(_1579_),
    .Q(\simon1.lfsr_capture[1] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[20]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net115),
    .D(_0053_),
    .Q_N(_1578_),
    .Q(\simon1.lfsr_capture[20] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[21]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net116),
    .D(_0054_),
    .Q_N(_1577_),
    .Q(\simon1.lfsr_capture[21] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[22]$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net117),
    .D(_0055_),
    .Q_N(_1576_),
    .Q(\simon1.lfsr_capture[22] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[23]$_SDFFE_PN0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net118),
    .D(_0056_),
    .Q_N(_1575_),
    .Q(\simon1.lfsr_capture[23] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[24]$_SDFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net119),
    .D(_0057_),
    .Q_N(_1574_),
    .Q(\simon1.lfsr_capture[24] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[25]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net120),
    .D(_0058_),
    .Q_N(_1573_),
    .Q(\simon1.lfsr_capture[25] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[26]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net121),
    .D(_0059_),
    .Q_N(_1572_),
    .Q(\simon1.lfsr_capture[26] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[27]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net122),
    .D(_0060_),
    .Q_N(_1571_),
    .Q(\simon1.lfsr_capture[27] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[28]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net123),
    .D(_0061_),
    .Q_N(_1570_),
    .Q(\simon1.lfsr_capture[28] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[29]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net124),
    .D(_0062_),
    .Q_N(_1569_),
    .Q(\simon1.lfsr_capture[29] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[2]$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net125),
    .D(_0063_),
    .Q_N(_1568_),
    .Q(\simon1.lfsr_capture[2] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[30]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net126),
    .D(_0064_),
    .Q_N(_1567_),
    .Q(\simon1.lfsr_capture[30] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[31]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net127),
    .D(_0065_),
    .Q_N(_1566_),
    .Q(\simon1.lfsr_capture[31] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[3]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net128),
    .D(_0066_),
    .Q_N(_1565_),
    .Q(\simon1.lfsr_capture[3] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[4]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net129),
    .D(_0067_),
    .Q_N(_1564_),
    .Q(\simon1.lfsr_capture[4] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[5]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net130),
    .D(_0068_),
    .Q_N(_1563_),
    .Q(\simon1.lfsr_capture[5] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[6]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net131),
    .D(_0069_),
    .Q_N(_1562_),
    .Q(\simon1.lfsr_capture[6] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[7]$_SDFFE_PN0P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net132),
    .D(_0070_),
    .Q_N(_1561_),
    .Q(\simon1.lfsr_capture[7] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[8]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net133),
    .D(_0071_),
    .Q_N(_1560_),
    .Q(\simon1.lfsr_capture[8] ));
 sg13g2_dfrbp_1 \simon1.lfsr_capture[9]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net134),
    .D(_0072_),
    .Q_N(_1559_),
    .Q(\simon1.lfsr_capture[9] ));
 sg13g2_dfrbp_1 \simon1.lfsr_cycles[0]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net135),
    .D(_0073_),
    .Q_N(_1558_),
    .Q(\simon1.lfsr_cycles[0] ));
 sg13g2_dfrbp_1 \simon1.lfsr_cycles[1]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net136),
    .D(_0074_),
    .Q_N(_1557_),
    .Q(\simon1.lfsr_cycles[1] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[0]$_SDFFE_PP0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net137),
    .D(_0075_),
    .Q_N(_1556_),
    .Q(\simon1.lfsr_inst.lfsr_out[0] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[10]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net138),
    .D(_0076_),
    .Q_N(_1555_),
    .Q(\simon1.lfsr_inst.lfsr_out[10] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[11]$_SDFFE_PP1P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net139),
    .D(_0077_),
    .Q_N(_1554_),
    .Q(\simon1.lfsr_inst.lfsr_out[11] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[12]$_SDFFE_PP1P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net140),
    .D(_0078_),
    .Q_N(_1553_),
    .Q(\simon1.lfsr_inst.lfsr_out[12] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[13]$_SDFFE_PP1P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net141),
    .D(_0079_),
    .Q_N(_1552_),
    .Q(\simon1.lfsr_inst.lfsr_out[13] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[14]$_SDFFE_PP1P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net142),
    .D(_0080_),
    .Q_N(_1551_),
    .Q(\simon1.lfsr_inst.lfsr_out[14] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[15]$_SDFFE_PP1P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net143),
    .D(_0081_),
    .Q_N(_1550_),
    .Q(\simon1.lfsr_inst.lfsr_out[15] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[16]$_SDFFE_PP0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net144),
    .D(_0082_),
    .Q_N(_1549_),
    .Q(\simon1.lfsr_inst.lfsr_out[16] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[17]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net145),
    .D(_0083_),
    .Q_N(_1548_),
    .Q(\simon1.lfsr_inst.lfsr_out[17] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[18]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net146),
    .D(_0084_),
    .Q_N(_1547_),
    .Q(\simon1.lfsr_inst.lfsr_out[18] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[19]$_SDFFE_PP1P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net147),
    .D(_0085_),
    .Q_N(_1546_),
    .Q(\simon1.lfsr_inst.lfsr_out[19] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[1]$_SDFFE_PP1P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net148),
    .D(_0086_),
    .Q_N(_1545_),
    .Q(\simon1.lfsr_inst.lfsr_out[1] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[20]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net149),
    .D(_0087_),
    .Q_N(_1544_),
    .Q(\simon1.lfsr_inst.lfsr_out[20] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[21]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net150),
    .D(_0088_),
    .Q_N(_1543_),
    .Q(\simon1.lfsr_inst.lfsr_out[21] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[22]$_SDFFE_PP1P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net151),
    .D(_0089_),
    .Q_N(_1542_),
    .Q(\simon1.lfsr_inst.lfsr_out[22] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[23]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net152),
    .D(_0090_),
    .Q_N(_1541_),
    .Q(\simon1.lfsr_inst.lfsr_out[23] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[24]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net153),
    .D(_0091_),
    .Q_N(_1540_),
    .Q(\simon1.lfsr_inst.lfsr_out[24] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[25]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net154),
    .D(_0092_),
    .Q_N(_1539_),
    .Q(\simon1.lfsr_inst.lfsr_out[25] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[26]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net155),
    .D(_0093_),
    .Q_N(_1538_),
    .Q(\simon1.lfsr_inst.lfsr_out[26] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[27]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net156),
    .D(_0094_),
    .Q_N(_1537_),
    .Q(\simon1.lfsr_inst.lfsr_out[27] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[28]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net157),
    .D(_0095_),
    .Q_N(_1536_),
    .Q(\simon1.lfsr_inst.lfsr_out[28] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[29]$_SDFFE_PP1P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net158),
    .D(_0096_),
    .Q_N(_1535_),
    .Q(\simon1.lfsr_inst.lfsr_out[29] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[2]$_SDFFE_PP0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net159),
    .D(_0097_),
    .Q_N(_1534_),
    .Q(\simon1.lfsr_inst.lfsr_out[2] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[30]$_SDFFE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net160),
    .D(_0098_),
    .Q_N(_1533_),
    .Q(\simon1.lfsr_inst.lfsr_out[30] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[31]$_SDFFE_PP0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net161),
    .D(_0099_),
    .Q_N(_1532_),
    .Q(\simon1.lfsr_inst.lfsr_out[31] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[3]$_SDFFE_PP1P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net162),
    .D(_0100_),
    .Q_N(_1531_),
    .Q(\simon1.lfsr_inst.lfsr_out[3] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[4]$_SDFFE_PP1P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net163),
    .D(_0101_),
    .Q_N(_1530_),
    .Q(\simon1.lfsr_inst.lfsr_out[4] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[5]$_SDFFE_PP1P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net164),
    .D(_0102_),
    .Q_N(_1529_),
    .Q(\simon1.lfsr_inst.lfsr_out[5] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[6]$_SDFFE_PP1P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net165),
    .D(_0103_),
    .Q_N(_1528_),
    .Q(\simon1.lfsr_inst.lfsr_out[6] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[7]$_SDFFE_PP1P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net166),
    .D(_0104_),
    .Q_N(_1527_),
    .Q(\simon1.lfsr_inst.lfsr_out[7] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[8]$_SDFFE_PP0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net167),
    .D(_0105_),
    .Q_N(_1526_),
    .Q(\simon1.lfsr_inst.lfsr_out[8] ));
 sg13g2_dfrbp_1 \simon1.lfsr_inst.lfsr_out[9]$_SDFFE_PP1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net168),
    .D(_0106_),
    .Q_N(_1525_),
    .Q(\simon1.lfsr_inst.lfsr_out[9] ));
 sg13g2_dfrbp_1 \simon1.lfsr_rewind$_SDFF_PN0_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net169),
    .D(_0107_),
    .Q_N(_1524_),
    .Q(\simon1.lfsr_inst.load_enable ));
 sg13g2_dfrbp_1 \simon1.lfsr_stopped$_SDFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net170),
    .D(_0108_),
    .Q_N(_1523_),
    .Q(\simon1.lfsr_stopped ));
 sg13g2_dfrbp_1 \simon1.millis_counter[0]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net171),
    .D(_0109_),
    .Q_N(_1522_),
    .Q(\simon1.millis_counter[0] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[1]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net172),
    .D(_0110_),
    .Q_N(_0015_),
    .Q(\simon1.millis_counter[1] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[2]$_SDFF_PN0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net173),
    .D(_0111_),
    .Q_N(_0016_),
    .Q(\simon1.millis_counter[2] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[3]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net174),
    .D(_0112_),
    .Q_N(_0017_),
    .Q(\simon1.millis_counter[3] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[4]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net175),
    .D(_0113_),
    .Q_N(_0018_),
    .Q(\simon1.millis_counter[4] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[5]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net176),
    .D(_0114_),
    .Q_N(_0019_),
    .Q(\simon1.millis_counter[5] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[6]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net177),
    .D(_0115_),
    .Q_N(_0020_),
    .Q(\simon1.millis_counter[6] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[7]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net178),
    .D(_0116_),
    .Q_N(_0021_),
    .Q(\simon1.millis_counter[7] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[8]$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net179),
    .D(_0117_),
    .Q_N(_0022_),
    .Q(\simon1.millis_counter[8] ));
 sg13g2_dfrbp_1 \simon1.millis_counter[9]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net180),
    .D(_0118_),
    .Q_N(_0023_),
    .Q(\simon1.millis_counter[9] ));
 sg13g2_dfrbp_1 \simon1.prev_btn[0]$_SDFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net181),
    .D(_0119_),
    .Q_N(_1521_),
    .Q(\simon1.prev_btn[0] ));
 sg13g2_dfrbp_1 \simon1.prev_btn[1]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net182),
    .D(_0120_),
    .Q_N(_1520_),
    .Q(\simon1.prev_btn[1] ));
 sg13g2_dfrbp_1 \simon1.prev_btn[2]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net183),
    .D(_0121_),
    .Q_N(_1519_),
    .Q(\simon1.prev_btn[2] ));
 sg13g2_dfrbp_1 \simon1.prev_btn[3]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net184),
    .D(_0122_),
    .Q_N(_1518_),
    .Q(\simon1.prev_btn[3] ));
 sg13g2_dfrbp_1 \simon1.score_ena$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net185),
    .D(_0123_),
    .Q_N(_0014_),
    .Q(\simon1.score_ena ));
 sg13g2_dfrbp_1 \simon1.score_inc$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net186),
    .D(_0124_),
    .Q_N(_1517_),
    .Q(\simon1.score_inc ));
 sg13g2_dfrbp_1 \simon1.score_inst.active_digit$_SDFF_PP0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net187),
    .D(_0125_),
    .Q_N(_0012_),
    .Q(\simon1.score_inst.active_digit ));
 sg13g2_dfrbp_1 \simon1.score_inst.digits[0]$_DFF_P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net188),
    .D(_0010_),
    .Q_N(_1596_),
    .Q(net14));
 sg13g2_dfrbp_1 \simon1.score_inst.digits[1]$_DFF_P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net189),
    .D(_0011_),
    .Q_N(_1516_),
    .Q(net15));
 sg13g2_dfrbp_1 \simon1.score_inst.ones[0]$_SDFFE_PP0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net190),
    .D(_0126_),
    .Q_N(_1515_),
    .Q(\simon1.score_inst.ones[0] ));
 sg13g2_dfrbp_1 \simon1.score_inst.ones[1]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net191),
    .D(_0127_),
    .Q_N(_1514_),
    .Q(\simon1.score_inst.ones[1] ));
 sg13g2_dfrbp_1 \simon1.score_inst.ones[2]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net192),
    .D(_0128_),
    .Q_N(_1513_),
    .Q(\simon1.score_inst.ones[2] ));
 sg13g2_dfrbp_1 \simon1.score_inst.ones[3]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net193),
    .D(_0129_),
    .Q_N(_1597_),
    .Q(\simon1.score_inst.ones[3] ));
 sg13g2_dfrbp_1 \simon1.score_inst.segments[0]$_DFF_P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net194),
    .D(_0213_),
    .Q_N(_1598_),
    .Q(net2));
 sg13g2_dfrbp_1 \simon1.score_inst.segments[1]$_DFF_P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net195),
    .D(_0214_),
    .Q_N(_1599_),
    .Q(net3));
 sg13g2_dfrbp_1 \simon1.score_inst.segments[2]$_DFF_P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net196),
    .D(_0215_),
    .Q_N(_1600_),
    .Q(net4));
 sg13g2_dfrbp_1 \simon1.score_inst.segments[3]$_DFF_P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net197),
    .D(_0216_),
    .Q_N(_1601_),
    .Q(net5));
 sg13g2_dfrbp_1 \simon1.score_inst.segments[4]$_DFF_P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net198),
    .D(_0217_),
    .Q_N(_1602_),
    .Q(net6));
 sg13g2_dfrbp_1 \simon1.score_inst.segments[5]$_DFF_P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net199),
    .D(_0218_),
    .Q_N(_1603_),
    .Q(net7));
 sg13g2_dfrbp_1 \simon1.score_inst.segments[6]$_DFF_P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net200),
    .D(_0219_),
    .Q_N(_1512_),
    .Q(net8));
 sg13g2_dfrbp_1 \simon1.score_inst.tens[0]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net201),
    .D(_0130_),
    .Q_N(_1511_),
    .Q(\simon1.score_inst.tens[0] ));
 sg13g2_dfrbp_1 \simon1.score_inst.tens[1]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net202),
    .D(_0131_),
    .Q_N(_1510_),
    .Q(\simon1.score_inst.tens[1] ));
 sg13g2_dfrbp_1 \simon1.score_inst.tens[2]$_SDFFE_PP0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net203),
    .D(_0132_),
    .Q_N(_1509_),
    .Q(\simon1.score_inst.tens[2] ));
 sg13g2_dfrbp_1 \simon1.score_inst.tens[3]$_SDFFE_PP0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net204),
    .D(_0133_),
    .Q_N(_1508_),
    .Q(\simon1.score_inst.tens[3] ));
 sg13g2_dfrbp_1 \simon1.score_rst$_SDFF_PN0_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net205),
    .D(_0134_),
    .Q_N(_1507_),
    .Q(\simon1.score_rst ));
 sg13g2_dfrbp_1 \simon1.seq_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net206),
    .D(_0135_),
    .Q_N(_1506_),
    .Q(\simon1.seq_counter[0] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net207),
    .D(_0136_),
    .Q_N(_1505_),
    .Q(\simon1.seq_counter[1] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net208),
    .D(_0137_),
    .Q_N(_1504_),
    .Q(\simon1.seq_counter[2] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net209),
    .D(_0138_),
    .Q_N(_1503_),
    .Q(\simon1.seq_counter[3] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net210),
    .D(_0139_),
    .Q_N(_1502_),
    .Q(\simon1.seq_counter[4] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net211),
    .D(_0140_),
    .Q_N(_1501_),
    .Q(\simon1.seq_counter[5] ));
 sg13g2_dfrbp_1 \simon1.seq_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net212),
    .D(_0141_),
    .Q_N(_1500_),
    .Q(\simon1.seq_counter[6] ));
 sg13g2_dfrbp_1 \simon1.seq_length[0]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net213),
    .D(_0142_),
    .Q_N(_1499_),
    .Q(\simon1.seq_length[0] ));
 sg13g2_dfrbp_1 \simon1.seq_length[1]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net214),
    .D(_0143_),
    .Q_N(_1498_),
    .Q(\simon1.seq_length[1] ));
 sg13g2_dfrbp_1 \simon1.seq_length[2]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net215),
    .D(_0144_),
    .Q_N(_0027_),
    .Q(\simon1.seq_length[2] ));
 sg13g2_dfrbp_1 \simon1.seq_length[3]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net216),
    .D(_0145_),
    .Q_N(_0028_),
    .Q(\simon1.seq_length[3] ));
 sg13g2_dfrbp_1 \simon1.seq_length[4]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net217),
    .D(_0146_),
    .Q_N(_0029_),
    .Q(\simon1.seq_length[4] ));
 sg13g2_dfrbp_1 \simon1.seq_length[5]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net218),
    .D(_0147_),
    .Q_N(_0030_),
    .Q(\simon1.seq_length[5] ));
 sg13g2_dfrbp_1 \simon1.seq_length[6]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net219),
    .D(_0148_),
    .Q_N(_0031_),
    .Q(\simon1.seq_length[6] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[0]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net220),
    .D(_0149_),
    .Q_N(_1497_),
    .Q(\simon1.sound_freq[0] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[1]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net221),
    .D(_0150_),
    .Q_N(_1496_),
    .Q(\simon1.sound_freq[1] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[2]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net222),
    .D(_0151_),
    .Q_N(_1495_),
    .Q(\simon1.sound_freq[2] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[3]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net223),
    .D(_0152_),
    .Q_N(_1494_),
    .Q(\simon1.sound_freq[3] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[4]$_SDFFE_PN0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net224),
    .D(_0153_),
    .Q_N(_1493_),
    .Q(\simon1.sound_freq[4] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[5]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net225),
    .D(_0154_),
    .Q_N(_1492_),
    .Q(\simon1.sound_freq[5] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[6]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net226),
    .D(_0155_),
    .Q_N(_1491_),
    .Q(\simon1.sound_freq[6] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[7]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net227),
    .D(_0156_),
    .Q_N(_1490_),
    .Q(\simon1.sound_freq[7] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[8]$_SDFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net228),
    .D(_0157_),
    .Q_N(_1489_),
    .Q(\simon1.sound_freq[8] ));
 sg13g2_dfrbp_1 \simon1.sound_freq[9]$_SDFFE_PN0P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net229),
    .D(_0158_),
    .Q_N(_1488_),
    .Q(\simon1.sound_freq[9] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.sound$_SDFFE_PP0N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net230),
    .D(_0159_),
    .Q_N(_0013_),
    .Q(\simon1.sound ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[0]$_SDFFE_PN0N_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net231),
    .D(_0160_),
    .Q_N(_1487_),
    .Q(\simon1.sound_gen_inst.tick_counter[0] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[10]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net232),
    .D(_0161_),
    .Q_N(_0034_),
    .Q(\simon1.sound_gen_inst.tick_counter[10] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[11]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net233),
    .D(_0162_),
    .Q_N(_1486_),
    .Q(\simon1.sound_gen_inst.tick_counter[11] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[12]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net234),
    .D(_0163_),
    .Q_N(_1485_),
    .Q(\simon1.sound_gen_inst.tick_counter[12] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[13]$_SDFFE_PN0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net235),
    .D(_0164_),
    .Q_N(_1484_),
    .Q(\simon1.sound_gen_inst.tick_counter[13] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[14]$_SDFFE_PN0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net236),
    .D(_0165_),
    .Q_N(_1483_),
    .Q(\simon1.sound_gen_inst.tick_counter[14] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[15]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net237),
    .D(_0166_),
    .Q_N(_1482_),
    .Q(\simon1.sound_gen_inst.tick_counter[15] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[16]$_SDFFE_PN0N_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net238),
    .D(_0167_),
    .Q_N(_1481_),
    .Q(\simon1.sound_gen_inst.tick_counter[16] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[17]$_SDFFE_PN0N_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net239),
    .D(_0168_),
    .Q_N(_1480_),
    .Q(\simon1.sound_gen_inst.tick_counter[17] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[18]$_SDFFE_PN0N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net240),
    .D(_0169_),
    .Q_N(_1479_),
    .Q(\simon1.sound_gen_inst.tick_counter[18] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[19]$_SDFFE_PN0N_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net241),
    .D(_0170_),
    .Q_N(_1478_),
    .Q(\simon1.sound_gen_inst.tick_counter[19] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[1]$_SDFFE_PN0N_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net242),
    .D(_0171_),
    .Q_N(_1477_),
    .Q(\simon1.sound_gen_inst.tick_counter[1] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[20]$_SDFFE_PN0N_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net243),
    .D(_0172_),
    .Q_N(_1476_),
    .Q(\simon1.sound_gen_inst.tick_counter[20] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[21]$_SDFFE_PN0N_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net244),
    .D(_0173_),
    .Q_N(_1475_),
    .Q(\simon1.sound_gen_inst.tick_counter[21] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[22]$_SDFFE_PN0N_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net245),
    .D(_0174_),
    .Q_N(_1474_),
    .Q(\simon1.sound_gen_inst.tick_counter[22] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[23]$_SDFFE_PN0N_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net246),
    .D(_0175_),
    .Q_N(_1473_),
    .Q(\simon1.sound_gen_inst.tick_counter[23] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[24]$_SDFFE_PN0N_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net247),
    .D(_0176_),
    .Q_N(_1472_),
    .Q(\simon1.sound_gen_inst.tick_counter[24] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[25]$_SDFFE_PN0N_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net248),
    .D(_0177_),
    .Q_N(_1471_),
    .Q(\simon1.sound_gen_inst.tick_counter[25] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[26]$_SDFFE_PN0N_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net249),
    .D(_0178_),
    .Q_N(_1470_),
    .Q(\simon1.sound_gen_inst.tick_counter[26] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[27]$_SDFFE_PN0N_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net250),
    .D(_0179_),
    .Q_N(_1469_),
    .Q(\simon1.sound_gen_inst.tick_counter[27] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[28]$_SDFFE_PN0N_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net251),
    .D(_0180_),
    .Q_N(_1468_),
    .Q(\simon1.sound_gen_inst.tick_counter[28] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[29]$_SDFFE_PN0N_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net252),
    .D(_0181_),
    .Q_N(_1467_),
    .Q(\simon1.sound_gen_inst.tick_counter[29] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[2]$_SDFFE_PN0N_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net253),
    .D(_0182_),
    .Q_N(_1466_),
    .Q(\simon1.sound_gen_inst.tick_counter[2] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[30]$_SDFFE_PN0N_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net254),
    .D(_0183_),
    .Q_N(_1465_),
    .Q(\simon1.sound_gen_inst.tick_counter[30] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[31]$_SDFFE_PN0N_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net255),
    .D(_0184_),
    .Q_N(_1464_),
    .Q(\simon1.sound_gen_inst.tick_counter[31] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[3]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net256),
    .D(_0185_),
    .Q_N(_1463_),
    .Q(\simon1.sound_gen_inst.tick_counter[3] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[4]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net257),
    .D(_0186_),
    .Q_N(_1462_),
    .Q(\simon1.sound_gen_inst.tick_counter[4] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[5]$_SDFFE_PN0N_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net258),
    .D(_0187_),
    .Q_N(_1461_),
    .Q(\simon1.sound_gen_inst.tick_counter[5] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[6]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net259),
    .D(_0188_),
    .Q_N(_1460_),
    .Q(\simon1.sound_gen_inst.tick_counter[6] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[7]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net260),
    .D(_0189_),
    .Q_N(_1459_),
    .Q(\simon1.sound_gen_inst.tick_counter[7] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[8]$_SDFFE_PN0N_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net261),
    .D(_0190_),
    .Q_N(_1458_),
    .Q(\simon1.sound_gen_inst.tick_counter[8] ));
 sg13g2_dfrbp_1 \simon1.sound_gen_inst.tick_counter[9]$_SDFFE_PN0N_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net262),
    .D(_0191_),
    .Q_N(_1604_),
    .Q(\simon1.sound_gen_inst.tick_counter[9] ));
 sg13g2_dfrbp_1 \simon1.state[0]$_DFF_P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net263),
    .D(_0000_),
    .Q_N(_1605_),
    .Q(\simon1.state[0] ));
 sg13g2_dfrbp_1 \simon1.state[1]$_DFF_P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net264),
    .D(_0001_),
    .Q_N(_0033_),
    .Q(\simon1.state[1] ));
 sg13g2_dfrbp_1 \simon1.state[2]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net265),
    .D(_0002_),
    .Q_N(_1606_),
    .Q(\simon1.state[2] ));
 sg13g2_dfrbp_1 \simon1.state[3]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net266),
    .D(_0003_),
    .Q_N(_1607_),
    .Q(\simon1.state[3] ));
 sg13g2_dfrbp_1 \simon1.state[4]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net267),
    .D(_0004_),
    .Q_N(_0009_),
    .Q(\simon1.state[4] ));
 sg13g2_dfrbp_1 \simon1.state[5]$_DFF_P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net268),
    .D(_0005_),
    .Q_N(_1608_),
    .Q(\simon1.state[5] ));
 sg13g2_dfrbp_1 \simon1.state[6]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net269),
    .D(_0006_),
    .Q_N(_1609_),
    .Q(\simon1.state[6] ));
 sg13g2_dfrbp_1 \simon1.state[7]$_DFF_P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net270),
    .D(_0007_),
    .Q_N(_0025_),
    .Q(\simon1.state[7] ));
 sg13g2_dfrbp_1 \simon1.state[8]$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net271),
    .D(_0008_),
    .Q_N(_0032_),
    .Q(\simon1.state[8] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[0]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net272),
    .D(_0192_),
    .Q_N(_0035_),
    .Q(\simon1.tick_counter[0] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[10]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net273),
    .D(_0193_),
    .Q_N(_1457_),
    .Q(\simon1.tick_counter[10] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[11]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net274),
    .D(_0194_),
    .Q_N(_1456_),
    .Q(\simon1.tick_counter[11] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[12]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net275),
    .D(_0195_),
    .Q_N(_1455_),
    .Q(\simon1.tick_counter[12] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[13]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net276),
    .D(_0196_),
    .Q_N(_1454_),
    .Q(\simon1.tick_counter[13] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[14]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net277),
    .D(_0197_),
    .Q_N(_1453_),
    .Q(\simon1.tick_counter[14] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[15]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net278),
    .D(_0198_),
    .Q_N(_1452_),
    .Q(\simon1.tick_counter[15] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[1]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net279),
    .D(_0199_),
    .Q_N(_1451_),
    .Q(\simon1.tick_counter[1] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[2]$_SDFF_PP0_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net280),
    .D(_0200_),
    .Q_N(_1450_),
    .Q(\simon1.tick_counter[2] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[3]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net281),
    .D(_0201_),
    .Q_N(_1449_),
    .Q(\simon1.tick_counter[3] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[4]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net282),
    .D(_0202_),
    .Q_N(_1448_),
    .Q(\simon1.tick_counter[4] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[5]$_SDFF_PP0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net283),
    .D(_0203_),
    .Q_N(_1447_),
    .Q(\simon1.tick_counter[5] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[6]$_SDFF_PP0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net284),
    .D(_0204_),
    .Q_N(_1446_),
    .Q(\simon1.tick_counter[6] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[7]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net285),
    .D(_0205_),
    .Q_N(_1445_),
    .Q(\simon1.tick_counter[7] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[8]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net286),
    .D(_0206_),
    .Q_N(_1444_),
    .Q(\simon1.tick_counter[8] ));
 sg13g2_dfrbp_1 \simon1.tick_counter[9]$_SDFF_PP0_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net287),
    .D(_0207_),
    .Q_N(_1443_),
    .Q(\simon1.tick_counter[9] ));
 sg13g2_dfrbp_1 \simon1.tone_sequence_counter[0]$_DFFE_PP_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net288),
    .D(_0208_),
    .Q_N(_0024_),
    .Q(\simon1.tone_sequence_counter[0] ));
 sg13g2_dfrbp_1 \simon1.tone_sequence_counter[1]$_DFFE_PP_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net289),
    .D(_0209_),
    .Q_N(_1442_),
    .Q(\simon1.tone_sequence_counter[1] ));
 sg13g2_dfrbp_1 \simon1.tone_sequence_counter[2]$_DFFE_PP_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net290),
    .D(_0210_),
    .Q_N(_0026_),
    .Q(\simon1.tone_sequence_counter[2] ));
 sg13g2_dfrbp_1 \simon1.user_input[0]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net291),
    .D(_0211_),
    .Q_N(_1441_),
    .Q(\simon1.user_input[0] ));
 sg13g2_dfrbp_1 \simon1.user_input[1]$_SDFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net292),
    .D(_0212_),
    .Q_N(_1440_),
    .Q(\simon1.user_input[1] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uio_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[0]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[1]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[2]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[3]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[4]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[5]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[6]));
 sg13g2_buf_2 fanout16 (.A(_0399_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0372_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0430_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0429_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_1008_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0621_),
    .X(net21));
 sg13g2_buf_4 fanout22 (.X(net22),
    .A(_0280_));
 sg13g2_buf_4 fanout23 (.X(net23),
    .A(_0266_));
 sg13g2_buf_2 fanout24 (.A(_0256_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1396_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0703_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1383_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1216_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1175_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1162_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0629_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0613_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0515_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1338_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1231_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1186_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1185_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1182_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1178_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0514_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1177_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0451_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0444_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0394_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0358_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1165_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1032_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_0971_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_0321_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0278_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0265_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1429_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1300_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1193_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1188_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1187_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1164_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1024_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1010_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0973_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0970_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0231_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1437_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1367_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1358_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1357_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1356_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1354_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1352_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1343_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1342_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_1340_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1332_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1329_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1325_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1121_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1078_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1062_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0972_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0956_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0951_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0950_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0948_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0934_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0968_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0939_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0938_),
    .X(net87));
 sg13g2_tielo _3036__88 (.L_LO(net88));
 sg13g2_tielo _3037__89 (.L_LO(net89));
 sg13g2_tielo _3039__90 (.L_LO(net90));
 sg13g2_tiehi _3030__92 (.L_HI(net92));
 sg13g2_tiehi _3031__93 (.L_HI(net93));
 sg13g2_tiehi _3032__94 (.L_HI(net94));
 sg13g2_tiehi _3033__95 (.L_HI(net95));
 sg13g2_tiehi _3034__96 (.L_HI(net96));
 sg13g2_tiehi _3035__97 (.L_HI(net97));
 sg13g2_tiehi \simon1.button_released$_SDFFE_PN0P__98  (.L_HI(net98));
 sg13g2_tiehi \simon1.led[0]$_SDFFE_PN0P__99  (.L_HI(net99));
 sg13g2_tiehi \simon1.led[1]$_SDFFE_PN0P__100  (.L_HI(net100));
 sg13g2_tiehi \simon1.led[2]$_SDFFE_PN0P__101  (.L_HI(net101));
 sg13g2_tiehi \simon1.led[3]$_SDFFE_PN0P__102  (.L_HI(net102));
 sg13g2_tiehi \simon1.lfsr_capture[0]$_SDFFE_PN0P__103  (.L_HI(net103));
 sg13g2_tiehi \simon1.lfsr_capture[10]$_SDFFE_PN0P__104  (.L_HI(net104));
 sg13g2_tiehi \simon1.lfsr_capture[11]$_SDFFE_PN0P__105  (.L_HI(net105));
 sg13g2_tiehi \simon1.lfsr_capture[12]$_SDFFE_PN0P__106  (.L_HI(net106));
 sg13g2_tiehi \simon1.lfsr_capture[13]$_SDFFE_PN0P__107  (.L_HI(net107));
 sg13g2_tiehi \simon1.lfsr_capture[14]$_SDFFE_PN0P__108  (.L_HI(net108));
 sg13g2_tiehi \simon1.lfsr_capture[15]$_SDFFE_PN0P__109  (.L_HI(net109));
 sg13g2_tiehi \simon1.lfsr_capture[16]$_SDFFE_PN0P__110  (.L_HI(net110));
 sg13g2_tiehi \simon1.lfsr_capture[17]$_SDFFE_PN0P__111  (.L_HI(net111));
 sg13g2_tiehi \simon1.lfsr_capture[18]$_SDFFE_PN0P__112  (.L_HI(net112));
 sg13g2_tiehi \simon1.lfsr_capture[19]$_SDFFE_PN0P__113  (.L_HI(net113));
 sg13g2_tiehi \simon1.lfsr_capture[1]$_SDFFE_PN0P__114  (.L_HI(net114));
 sg13g2_tiehi \simon1.lfsr_capture[20]$_SDFFE_PN0P__115  (.L_HI(net115));
 sg13g2_tiehi \simon1.lfsr_capture[21]$_SDFFE_PN0P__116  (.L_HI(net116));
 sg13g2_tiehi \simon1.lfsr_capture[22]$_SDFFE_PN0P__117  (.L_HI(net117));
 sg13g2_tiehi \simon1.lfsr_capture[23]$_SDFFE_PN0P__118  (.L_HI(net118));
 sg13g2_tiehi \simon1.lfsr_capture[24]$_SDFFE_PN0P__119  (.L_HI(net119));
 sg13g2_tiehi \simon1.lfsr_capture[25]$_SDFFE_PN0P__120  (.L_HI(net120));
 sg13g2_tiehi \simon1.lfsr_capture[26]$_SDFFE_PN0P__121  (.L_HI(net121));
 sg13g2_tiehi \simon1.lfsr_capture[27]$_SDFFE_PN0P__122  (.L_HI(net122));
 sg13g2_tiehi \simon1.lfsr_capture[28]$_SDFFE_PN0P__123  (.L_HI(net123));
 sg13g2_tiehi \simon1.lfsr_capture[29]$_SDFFE_PN0P__124  (.L_HI(net124));
 sg13g2_tiehi \simon1.lfsr_capture[2]$_SDFFE_PN0P__125  (.L_HI(net125));
 sg13g2_tiehi \simon1.lfsr_capture[30]$_SDFFE_PN0P__126  (.L_HI(net126));
 sg13g2_tiehi \simon1.lfsr_capture[31]$_SDFFE_PN0P__127  (.L_HI(net127));
 sg13g2_tiehi \simon1.lfsr_capture[3]$_SDFFE_PN0P__128  (.L_HI(net128));
 sg13g2_tiehi \simon1.lfsr_capture[4]$_SDFFE_PN0P__129  (.L_HI(net129));
 sg13g2_tiehi \simon1.lfsr_capture[5]$_SDFFE_PN0P__130  (.L_HI(net130));
 sg13g2_tiehi \simon1.lfsr_capture[6]$_SDFFE_PN0P__131  (.L_HI(net131));
 sg13g2_tiehi \simon1.lfsr_capture[7]$_SDFFE_PN0P__132  (.L_HI(net132));
 sg13g2_tiehi \simon1.lfsr_capture[8]$_SDFFE_PN0P__133  (.L_HI(net133));
 sg13g2_tiehi \simon1.lfsr_capture[9]$_SDFFE_PN0P__134  (.L_HI(net134));
 sg13g2_tiehi \simon1.lfsr_cycles[0]$_SDFF_PN0__135  (.L_HI(net135));
 sg13g2_tiehi \simon1.lfsr_cycles[1]$_SDFF_PN0__136  (.L_HI(net136));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[0]$_SDFFE_PP0P__137  (.L_HI(net137));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[10]$_SDFFE_PP0P__138  (.L_HI(net138));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[11]$_SDFFE_PP1P__139  (.L_HI(net139));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[12]$_SDFFE_PP1P__140  (.L_HI(net140));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[13]$_SDFFE_PP1P__141  (.L_HI(net141));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[14]$_SDFFE_PP1P__142  (.L_HI(net142));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[15]$_SDFFE_PP1P__143  (.L_HI(net143));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[16]$_SDFFE_PP0P__144  (.L_HI(net144));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[17]$_SDFFE_PP0P__145  (.L_HI(net145));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[18]$_SDFFE_PP0P__146  (.L_HI(net146));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[19]$_SDFFE_PP1P__147  (.L_HI(net147));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[1]$_SDFFE_PP1P__148  (.L_HI(net148));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[20]$_SDFFE_PP0P__149  (.L_HI(net149));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[21]$_SDFFE_PP0P__150  (.L_HI(net150));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[22]$_SDFFE_PP1P__151  (.L_HI(net151));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[23]$_SDFFE_PP0P__152  (.L_HI(net152));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[24]$_SDFFE_PP0P__153  (.L_HI(net153));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[25]$_SDFFE_PP0P__154  (.L_HI(net154));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[26]$_SDFFE_PP0P__155  (.L_HI(net155));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[27]$_SDFFE_PP0P__156  (.L_HI(net156));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[28]$_SDFFE_PP0P__157  (.L_HI(net157));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[29]$_SDFFE_PP1P__158  (.L_HI(net158));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[2]$_SDFFE_PP0P__159  (.L_HI(net159));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[30]$_SDFFE_PP0P__160  (.L_HI(net160));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[31]$_SDFFE_PP0P__161  (.L_HI(net161));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[3]$_SDFFE_PP1P__162  (.L_HI(net162));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[4]$_SDFFE_PP1P__163  (.L_HI(net163));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[5]$_SDFFE_PP1P__164  (.L_HI(net164));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[6]$_SDFFE_PP1P__165  (.L_HI(net165));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[7]$_SDFFE_PP1P__166  (.L_HI(net166));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[8]$_SDFFE_PP0P__167  (.L_HI(net167));
 sg13g2_tiehi \simon1.lfsr_inst.lfsr_out[9]$_SDFFE_PP1P__168  (.L_HI(net168));
 sg13g2_tiehi \simon1.lfsr_rewind$_SDFF_PN0__169  (.L_HI(net169));
 sg13g2_tiehi \simon1.lfsr_stopped$_SDFFE_PN0P__170  (.L_HI(net170));
 sg13g2_tiehi \simon1.millis_counter[0]$_SDFF_PN0__171  (.L_HI(net171));
 sg13g2_tiehi \simon1.millis_counter[1]$_SDFF_PN0__172  (.L_HI(net172));
 sg13g2_tiehi \simon1.millis_counter[2]$_SDFF_PN0__173  (.L_HI(net173));
 sg13g2_tiehi \simon1.millis_counter[3]$_SDFF_PN0__174  (.L_HI(net174));
 sg13g2_tiehi \simon1.millis_counter[4]$_SDFF_PN0__175  (.L_HI(net175));
 sg13g2_tiehi \simon1.millis_counter[5]$_SDFF_PN0__176  (.L_HI(net176));
 sg13g2_tiehi \simon1.millis_counter[6]$_SDFF_PN0__177  (.L_HI(net177));
 sg13g2_tiehi \simon1.millis_counter[7]$_SDFF_PN0__178  (.L_HI(net178));
 sg13g2_tiehi \simon1.millis_counter[8]$_SDFF_PN0__179  (.L_HI(net179));
 sg13g2_tiehi \simon1.millis_counter[9]$_SDFF_PN0__180  (.L_HI(net180));
 sg13g2_tiehi \simon1.prev_btn[0]$_SDFFE_PN0P__181  (.L_HI(net181));
 sg13g2_tiehi \simon1.prev_btn[1]$_SDFFE_PN0P__182  (.L_HI(net182));
 sg13g2_tiehi \simon1.prev_btn[2]$_SDFFE_PN0P__183  (.L_HI(net183));
 sg13g2_tiehi \simon1.prev_btn[3]$_SDFFE_PN0P__184  (.L_HI(net184));
 sg13g2_tiehi \simon1.score_ena$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \simon1.score_inc$_SDFF_PN0__186  (.L_HI(net186));
 sg13g2_tiehi \simon1.score_inst.active_digit$_SDFF_PP0__187  (.L_HI(net187));
 sg13g2_tiehi \simon1.score_inst.digits[0]$_DFF_P__188  (.L_HI(net188));
 sg13g2_tiehi \simon1.score_inst.digits[1]$_DFF_P__189  (.L_HI(net189));
 sg13g2_tiehi \simon1.score_inst.ones[0]$_SDFFE_PP0P__190  (.L_HI(net190));
 sg13g2_tiehi \simon1.score_inst.ones[1]$_SDFFE_PP0P__191  (.L_HI(net191));
 sg13g2_tiehi \simon1.score_inst.ones[2]$_SDFFE_PP0P__192  (.L_HI(net192));
 sg13g2_tiehi \simon1.score_inst.ones[3]$_SDFFE_PP0P__193  (.L_HI(net193));
 sg13g2_tiehi \simon1.score_inst.segments[0]$_DFF_P__194  (.L_HI(net194));
 sg13g2_tiehi \simon1.score_inst.segments[1]$_DFF_P__195  (.L_HI(net195));
 sg13g2_tiehi \simon1.score_inst.segments[2]$_DFF_P__196  (.L_HI(net196));
 sg13g2_tiehi \simon1.score_inst.segments[3]$_DFF_P__197  (.L_HI(net197));
 sg13g2_tiehi \simon1.score_inst.segments[4]$_DFF_P__198  (.L_HI(net198));
 sg13g2_tiehi \simon1.score_inst.segments[5]$_DFF_P__199  (.L_HI(net199));
 sg13g2_tiehi \simon1.score_inst.segments[6]$_DFF_P__200  (.L_HI(net200));
 sg13g2_tiehi \simon1.score_inst.tens[0]$_SDFFE_PP0P__201  (.L_HI(net201));
 sg13g2_tiehi \simon1.score_inst.tens[1]$_SDFFE_PP0P__202  (.L_HI(net202));
 sg13g2_tiehi \simon1.score_inst.tens[2]$_SDFFE_PP0P__203  (.L_HI(net203));
 sg13g2_tiehi \simon1.score_inst.tens[3]$_SDFFE_PP0P__204  (.L_HI(net204));
 sg13g2_tiehi \simon1.score_rst$_SDFF_PN0__205  (.L_HI(net205));
 sg13g2_tiehi \simon1.seq_counter[0]$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \simon1.seq_counter[1]$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_tiehi \simon1.seq_counter[2]$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \simon1.seq_counter[3]$_SDFFE_PN0P__209  (.L_HI(net209));
 sg13g2_tiehi \simon1.seq_counter[4]$_SDFFE_PN0P__210  (.L_HI(net210));
 sg13g2_tiehi \simon1.seq_counter[5]$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \simon1.seq_counter[6]$_SDFFE_PN0P__212  (.L_HI(net212));
 sg13g2_tiehi \simon1.seq_length[0]$_SDFFE_PN0P__213  (.L_HI(net213));
 sg13g2_tiehi \simon1.seq_length[1]$_SDFFE_PN0P__214  (.L_HI(net214));
 sg13g2_tiehi \simon1.seq_length[2]$_SDFFE_PN0P__215  (.L_HI(net215));
 sg13g2_tiehi \simon1.seq_length[3]$_SDFFE_PN0P__216  (.L_HI(net216));
 sg13g2_tiehi \simon1.seq_length[4]$_SDFFE_PN0P__217  (.L_HI(net217));
 sg13g2_tiehi \simon1.seq_length[5]$_SDFFE_PN0P__218  (.L_HI(net218));
 sg13g2_tiehi \simon1.seq_length[6]$_SDFFE_PN0P__219  (.L_HI(net219));
 sg13g2_tiehi \simon1.sound_freq[0]$_SDFFE_PN0P__220  (.L_HI(net220));
 sg13g2_tiehi \simon1.sound_freq[1]$_SDFFE_PN0P__221  (.L_HI(net221));
 sg13g2_tiehi \simon1.sound_freq[2]$_SDFFE_PN0P__222  (.L_HI(net222));
 sg13g2_tiehi \simon1.sound_freq[3]$_SDFFE_PN0P__223  (.L_HI(net223));
 sg13g2_tiehi \simon1.sound_freq[4]$_SDFFE_PN0P__224  (.L_HI(net224));
 sg13g2_tiehi \simon1.sound_freq[5]$_SDFFE_PN0P__225  (.L_HI(net225));
 sg13g2_tiehi \simon1.sound_freq[6]$_SDFFE_PN0P__226  (.L_HI(net226));
 sg13g2_tiehi \simon1.sound_freq[7]$_SDFFE_PN0P__227  (.L_HI(net227));
 sg13g2_tiehi \simon1.sound_freq[8]$_SDFFE_PN0P__228  (.L_HI(net228));
 sg13g2_tiehi \simon1.sound_freq[9]$_SDFFE_PN0P__229  (.L_HI(net229));
 sg13g2_tiehi \simon1.sound_gen_inst.sound$_SDFFE_PP0N__230  (.L_HI(net230));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[0]$_SDFFE_PN0N__231  (.L_HI(net231));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[10]$_SDFFE_PN0N__232  (.L_HI(net232));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[11]$_SDFFE_PN0N__233  (.L_HI(net233));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[12]$_SDFFE_PN0N__234  (.L_HI(net234));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[13]$_SDFFE_PN0N__235  (.L_HI(net235));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[14]$_SDFFE_PN0N__236  (.L_HI(net236));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[15]$_SDFFE_PN0N__237  (.L_HI(net237));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[16]$_SDFFE_PN0N__238  (.L_HI(net238));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[17]$_SDFFE_PN0N__239  (.L_HI(net239));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[18]$_SDFFE_PN0N__240  (.L_HI(net240));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[19]$_SDFFE_PN0N__241  (.L_HI(net241));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[1]$_SDFFE_PN0N__242  (.L_HI(net242));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[20]$_SDFFE_PN0N__243  (.L_HI(net243));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[21]$_SDFFE_PN0N__244  (.L_HI(net244));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[22]$_SDFFE_PN0N__245  (.L_HI(net245));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[23]$_SDFFE_PN0N__246  (.L_HI(net246));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[24]$_SDFFE_PN0N__247  (.L_HI(net247));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[25]$_SDFFE_PN0N__248  (.L_HI(net248));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[26]$_SDFFE_PN0N__249  (.L_HI(net249));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[27]$_SDFFE_PN0N__250  (.L_HI(net250));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[28]$_SDFFE_PN0N__251  (.L_HI(net251));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[29]$_SDFFE_PN0N__252  (.L_HI(net252));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[2]$_SDFFE_PN0N__253  (.L_HI(net253));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[30]$_SDFFE_PN0N__254  (.L_HI(net254));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[31]$_SDFFE_PN0N__255  (.L_HI(net255));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[3]$_SDFFE_PN0N__256  (.L_HI(net256));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[4]$_SDFFE_PN0N__257  (.L_HI(net257));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[5]$_SDFFE_PN0N__258  (.L_HI(net258));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[6]$_SDFFE_PN0N__259  (.L_HI(net259));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[7]$_SDFFE_PN0N__260  (.L_HI(net260));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[8]$_SDFFE_PN0N__261  (.L_HI(net261));
 sg13g2_tiehi \simon1.sound_gen_inst.tick_counter[9]$_SDFFE_PN0N__262  (.L_HI(net262));
 sg13g2_tiehi \simon1.state[0]$_DFF_P__263  (.L_HI(net263));
 sg13g2_tiehi \simon1.state[1]$_DFF_P__264  (.L_HI(net264));
 sg13g2_tiehi \simon1.state[2]$_DFF_P__265  (.L_HI(net265));
 sg13g2_tiehi \simon1.state[3]$_DFF_P__266  (.L_HI(net266));
 sg13g2_tiehi \simon1.state[4]$_DFF_P__267  (.L_HI(net267));
 sg13g2_tiehi \simon1.state[5]$_DFF_P__268  (.L_HI(net268));
 sg13g2_tiehi \simon1.state[6]$_DFF_P__269  (.L_HI(net269));
 sg13g2_tiehi \simon1.state[7]$_DFF_P__270  (.L_HI(net270));
 sg13g2_tiehi \simon1.state[8]$_DFF_P__271  (.L_HI(net271));
 sg13g2_tiehi \simon1.tick_counter[0]$_SDFF_PP0__272  (.L_HI(net272));
 sg13g2_tiehi \simon1.tick_counter[10]$_SDFF_PP0__273  (.L_HI(net273));
 sg13g2_tiehi \simon1.tick_counter[11]$_SDFF_PP0__274  (.L_HI(net274));
 sg13g2_tiehi \simon1.tick_counter[12]$_SDFF_PP0__275  (.L_HI(net275));
 sg13g2_tiehi \simon1.tick_counter[13]$_SDFF_PP0__276  (.L_HI(net276));
 sg13g2_tiehi \simon1.tick_counter[14]$_SDFF_PP0__277  (.L_HI(net277));
 sg13g2_tiehi \simon1.tick_counter[15]$_SDFF_PP0__278  (.L_HI(net278));
 sg13g2_tiehi \simon1.tick_counter[1]$_SDFF_PP0__279  (.L_HI(net279));
 sg13g2_tiehi \simon1.tick_counter[2]$_SDFF_PP0__280  (.L_HI(net280));
 sg13g2_tiehi \simon1.tick_counter[3]$_SDFF_PP0__281  (.L_HI(net281));
 sg13g2_tiehi \simon1.tick_counter[4]$_SDFF_PP0__282  (.L_HI(net282));
 sg13g2_tiehi \simon1.tick_counter[5]$_SDFF_PP0__283  (.L_HI(net283));
 sg13g2_tiehi \simon1.tick_counter[6]$_SDFF_PP0__284  (.L_HI(net284));
 sg13g2_tiehi \simon1.tick_counter[7]$_SDFF_PP0__285  (.L_HI(net285));
 sg13g2_tiehi \simon1.tick_counter[8]$_SDFF_PP0__286  (.L_HI(net286));
 sg13g2_tiehi \simon1.tick_counter[9]$_SDFF_PP0__287  (.L_HI(net287));
 sg13g2_tiehi \simon1.tone_sequence_counter[0]$_DFFE_PP__288  (.L_HI(net288));
 sg13g2_tiehi \simon1.tone_sequence_counter[1]$_DFFE_PP__289  (.L_HI(net289));
 sg13g2_tiehi \simon1.tone_sequence_counter[2]$_DFFE_PP__290  (.L_HI(net290));
 sg13g2_tiehi \simon1.user_input[0]$_SDFFE_PN0P__291  (.L_HI(net291));
 sg13g2_tiehi \simon1.user_input[1]$_SDFFE_PN0P__292  (.L_HI(net292));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_17__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_4 FILLER_0_119 ();
 sg13g2_fill_2 FILLER_0_123 ();
 sg13g2_decap_4 FILLER_0_134 ();
 sg13g2_fill_2 FILLER_0_142 ();
 sg13g2_fill_1 FILLER_0_144 ();
 sg13g2_fill_2 FILLER_0_160 ();
 sg13g2_fill_1 FILLER_0_162 ();
 sg13g2_fill_1 FILLER_0_187 ();
 sg13g2_fill_1 FILLER_0_218 ();
 sg13g2_fill_1 FILLER_0_224 ();
 sg13g2_fill_1 FILLER_0_261 ();
 sg13g2_fill_1 FILLER_0_296 ();
 sg13g2_fill_1 FILLER_0_323 ();
 sg13g2_fill_1 FILLER_0_350 ();
 sg13g2_fill_2 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_4 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_4 FILLER_1_119 ();
 sg13g2_fill_1 FILLER_1_321 ();
 sg13g2_fill_2 FILLER_1_331 ();
 sg13g2_fill_2 FILLER_1_343 ();
 sg13g2_fill_1 FILLER_1_350 ();
 sg13g2_fill_2 FILLER_1_381 ();
 sg13g2_fill_1 FILLER_1_383 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_4 FILLER_2_119 ();
 sg13g2_fill_1 FILLER_2_138 ();
 sg13g2_fill_1 FILLER_2_157 ();
 sg13g2_fill_1 FILLER_2_163 ();
 sg13g2_fill_1 FILLER_2_193 ();
 sg13g2_fill_2 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_209 ();
 sg13g2_decap_4 FILLER_2_216 ();
 sg13g2_fill_2 FILLER_2_220 ();
 sg13g2_fill_2 FILLER_2_262 ();
 sg13g2_fill_2 FILLER_2_269 ();
 sg13g2_fill_1 FILLER_2_277 ();
 sg13g2_fill_2 FILLER_2_372 ();
 sg13g2_fill_1 FILLER_2_374 ();
 sg13g2_fill_2 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_4 FILLER_3_35 ();
 sg13g2_fill_1 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_44 ();
 sg13g2_decap_8 FILLER_3_51 ();
 sg13g2_decap_8 FILLER_3_58 ();
 sg13g2_decap_8 FILLER_3_65 ();
 sg13g2_decap_8 FILLER_3_72 ();
 sg13g2_decap_8 FILLER_3_79 ();
 sg13g2_decap_8 FILLER_3_86 ();
 sg13g2_decap_8 FILLER_3_93 ();
 sg13g2_fill_2 FILLER_3_100 ();
 sg13g2_fill_1 FILLER_3_102 ();
 sg13g2_fill_2 FILLER_3_155 ();
 sg13g2_fill_1 FILLER_3_157 ();
 sg13g2_fill_2 FILLER_3_184 ();
 sg13g2_fill_1 FILLER_3_186 ();
 sg13g2_fill_2 FILLER_3_250 ();
 sg13g2_fill_1 FILLER_3_252 ();
 sg13g2_fill_1 FILLER_3_269 ();
 sg13g2_fill_2 FILLER_3_302 ();
 sg13g2_fill_1 FILLER_3_345 ();
 sg13g2_decap_4 FILLER_3_390 ();
 sg13g2_fill_1 FILLER_3_398 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_4 FILLER_4_28 ();
 sg13g2_fill_1 FILLER_4_32 ();
 sg13g2_fill_2 FILLER_4_105 ();
 sg13g2_fill_1 FILLER_4_107 ();
 sg13g2_decap_4 FILLER_4_120 ();
 sg13g2_fill_2 FILLER_4_124 ();
 sg13g2_fill_2 FILLER_4_136 ();
 sg13g2_fill_2 FILLER_4_143 ();
 sg13g2_fill_1 FILLER_4_150 ();
 sg13g2_fill_1 FILLER_4_156 ();
 sg13g2_fill_1 FILLER_4_162 ();
 sg13g2_fill_1 FILLER_4_193 ();
 sg13g2_fill_1 FILLER_4_198 ();
 sg13g2_fill_2 FILLER_4_203 ();
 sg13g2_fill_1 FILLER_4_205 ();
 sg13g2_decap_4 FILLER_4_211 ();
 sg13g2_fill_1 FILLER_4_215 ();
 sg13g2_fill_1 FILLER_4_334 ();
 sg13g2_fill_1 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_418 ();
 sg13g2_decap_4 FILLER_4_425 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_11 ();
 sg13g2_fill_2 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_fill_1 FILLER_5_102 ();
 sg13g2_fill_2 FILLER_5_149 ();
 sg13g2_fill_1 FILLER_5_155 ();
 sg13g2_fill_2 FILLER_5_161 ();
 sg13g2_fill_2 FILLER_5_168 ();
 sg13g2_fill_2 FILLER_5_174 ();
 sg13g2_decap_4 FILLER_5_249 ();
 sg13g2_fill_2 FILLER_5_253 ();
 sg13g2_fill_2 FILLER_5_271 ();
 sg13g2_fill_2 FILLER_5_290 ();
 sg13g2_fill_1 FILLER_5_297 ();
 sg13g2_fill_1 FILLER_5_303 ();
 sg13g2_fill_1 FILLER_5_308 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_412 ();
 sg13g2_decap_8 FILLER_5_419 ();
 sg13g2_decap_4 FILLER_5_426 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_14 ();
 sg13g2_fill_2 FILLER_6_18 ();
 sg13g2_decap_4 FILLER_6_24 ();
 sg13g2_fill_1 FILLER_6_32 ();
 sg13g2_fill_2 FILLER_6_68 ();
 sg13g2_fill_1 FILLER_6_70 ();
 sg13g2_decap_4 FILLER_6_75 ();
 sg13g2_fill_1 FILLER_6_83 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_fill_1 FILLER_6_104 ();
 sg13g2_fill_1 FILLER_6_154 ();
 sg13g2_fill_1 FILLER_6_159 ();
 sg13g2_fill_1 FILLER_6_164 ();
 sg13g2_fill_1 FILLER_6_175 ();
 sg13g2_fill_1 FILLER_6_181 ();
 sg13g2_fill_2 FILLER_6_235 ();
 sg13g2_fill_2 FILLER_6_241 ();
 sg13g2_fill_2 FILLER_6_293 ();
 sg13g2_fill_2 FILLER_6_339 ();
 sg13g2_fill_1 FILLER_6_345 ();
 sg13g2_fill_1 FILLER_6_356 ();
 sg13g2_fill_2 FILLER_6_361 ();
 sg13g2_fill_1 FILLER_6_363 ();
 sg13g2_fill_1 FILLER_6_373 ();
 sg13g2_fill_1 FILLER_6_384 ();
 sg13g2_fill_1 FILLER_6_390 ();
 sg13g2_fill_2 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_decap_4 FILLER_7_26 ();
 sg13g2_fill_1 FILLER_7_63 ();
 sg13g2_fill_2 FILLER_7_124 ();
 sg13g2_fill_1 FILLER_7_160 ();
 sg13g2_fill_1 FILLER_7_174 ();
 sg13g2_fill_2 FILLER_7_224 ();
 sg13g2_fill_2 FILLER_7_308 ();
 sg13g2_fill_2 FILLER_7_314 ();
 sg13g2_fill_1 FILLER_7_316 ();
 sg13g2_fill_2 FILLER_7_336 ();
 sg13g2_fill_1 FILLER_7_338 ();
 sg13g2_fill_2 FILLER_7_343 ();
 sg13g2_fill_2 FILLER_7_381 ();
 sg13g2_fill_1 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_414 ();
 sg13g2_decap_8 FILLER_7_421 ();
 sg13g2_fill_2 FILLER_7_428 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_4 ();
 sg13g2_fill_2 FILLER_8_51 ();
 sg13g2_fill_1 FILLER_8_53 ();
 sg13g2_fill_2 FILLER_8_92 ();
 sg13g2_fill_1 FILLER_8_94 ();
 sg13g2_fill_1 FILLER_8_198 ();
 sg13g2_fill_1 FILLER_8_204 ();
 sg13g2_fill_1 FILLER_8_210 ();
 sg13g2_fill_2 FILLER_8_237 ();
 sg13g2_fill_1 FILLER_8_243 ();
 sg13g2_fill_2 FILLER_8_277 ();
 sg13g2_fill_1 FILLER_8_279 ();
 sg13g2_decap_4 FILLER_8_302 ();
 sg13g2_fill_1 FILLER_8_306 ();
 sg13g2_fill_1 FILLER_8_321 ();
 sg13g2_fill_1 FILLER_8_327 ();
 sg13g2_fill_1 FILLER_9_12 ();
 sg13g2_fill_1 FILLER_9_25 ();
 sg13g2_fill_1 FILLER_9_30 ();
 sg13g2_fill_1 FILLER_9_39 ();
 sg13g2_fill_1 FILLER_9_50 ();
 sg13g2_fill_1 FILLER_9_55 ();
 sg13g2_fill_1 FILLER_9_80 ();
 sg13g2_fill_2 FILLER_9_136 ();
 sg13g2_fill_1 FILLER_9_179 ();
 sg13g2_fill_1 FILLER_9_190 ();
 sg13g2_fill_1 FILLER_9_196 ();
 sg13g2_fill_1 FILLER_9_201 ();
 sg13g2_fill_1 FILLER_9_207 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_228 ();
 sg13g2_fill_1 FILLER_9_260 ();
 sg13g2_fill_1 FILLER_9_271 ();
 sg13g2_fill_2 FILLER_9_313 ();
 sg13g2_fill_1 FILLER_9_325 ();
 sg13g2_fill_1 FILLER_9_352 ();
 sg13g2_fill_1 FILLER_9_362 ();
 sg13g2_fill_1 FILLER_9_378 ();
 sg13g2_fill_1 FILLER_9_384 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_fill_1 FILLER_10_107 ();
 sg13g2_fill_2 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_195 ();
 sg13g2_decap_8 FILLER_10_233 ();
 sg13g2_fill_2 FILLER_10_240 ();
 sg13g2_fill_2 FILLER_10_246 ();
 sg13g2_fill_2 FILLER_10_257 ();
 sg13g2_decap_4 FILLER_10_287 ();
 sg13g2_fill_2 FILLER_10_295 ();
 sg13g2_fill_1 FILLER_10_307 ();
 sg13g2_decap_4 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_371 ();
 sg13g2_fill_2 FILLER_10_402 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_62 ();
 sg13g2_fill_1 FILLER_11_64 ();
 sg13g2_fill_1 FILLER_11_135 ();
 sg13g2_fill_1 FILLER_11_160 ();
 sg13g2_fill_1 FILLER_11_226 ();
 sg13g2_decap_4 FILLER_11_230 ();
 sg13g2_fill_2 FILLER_11_264 ();
 sg13g2_fill_1 FILLER_11_266 ();
 sg13g2_fill_2 FILLER_11_297 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_4 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_337 ();
 sg13g2_decap_8 FILLER_11_344 ();
 sg13g2_fill_2 FILLER_11_351 ();
 sg13g2_fill_1 FILLER_11_353 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_48 ();
 sg13g2_fill_2 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_90 ();
 sg13g2_decap_4 FILLER_12_97 ();
 sg13g2_fill_2 FILLER_12_110 ();
 sg13g2_fill_2 FILLER_12_116 ();
 sg13g2_fill_1 FILLER_12_118 ();
 sg13g2_fill_1 FILLER_12_145 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_fill_1 FILLER_12_158 ();
 sg13g2_fill_1 FILLER_12_185 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_217 ();
 sg13g2_decap_4 FILLER_12_249 ();
 sg13g2_fill_2 FILLER_12_257 ();
 sg13g2_fill_2 FILLER_12_263 ();
 sg13g2_fill_1 FILLER_12_265 ();
 sg13g2_fill_2 FILLER_12_270 ();
 sg13g2_fill_1 FILLER_12_272 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_fill_1 FILLER_12_279 ();
 sg13g2_decap_4 FILLER_12_293 ();
 sg13g2_fill_1 FILLER_12_379 ();
 sg13g2_decap_4 FILLER_12_406 ();
 sg13g2_fill_2 FILLER_12_410 ();
 sg13g2_fill_2 FILLER_12_416 ();
 sg13g2_fill_1 FILLER_12_418 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_20 ();
 sg13g2_fill_1 FILLER_13_33 ();
 sg13g2_fill_1 FILLER_13_38 ();
 sg13g2_fill_1 FILLER_13_43 ();
 sg13g2_decap_8 FILLER_13_51 ();
 sg13g2_fill_2 FILLER_13_58 ();
 sg13g2_decap_4 FILLER_13_117 ();
 sg13g2_fill_1 FILLER_13_155 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_fill_2 FILLER_13_184 ();
 sg13g2_fill_1 FILLER_13_186 ();
 sg13g2_decap_4 FILLER_13_215 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_225 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_fill_1 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_252 ();
 sg13g2_fill_2 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_317 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_2 FILLER_13_327 ();
 sg13g2_fill_1 FILLER_13_337 ();
 sg13g2_fill_2 FILLER_13_358 ();
 sg13g2_fill_1 FILLER_13_360 ();
 sg13g2_fill_1 FILLER_13_374 ();
 sg13g2_decap_8 FILLER_13_383 ();
 sg13g2_decap_4 FILLER_13_390 ();
 sg13g2_fill_1 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_4 FILLER_13_424 ();
 sg13g2_fill_2 FILLER_13_428 ();
 sg13g2_fill_1 FILLER_14_26 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_fill_2 FILLER_14_126 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_fill_1 FILLER_14_169 ();
 sg13g2_fill_2 FILLER_14_192 ();
 sg13g2_fill_1 FILLER_14_194 ();
 sg13g2_fill_2 FILLER_14_200 ();
 sg13g2_fill_1 FILLER_14_202 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_fill_1 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_409 ();
 sg13g2_decap_8 FILLER_14_416 ();
 sg13g2_decap_8 FILLER_14_423 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_fill_1 FILLER_15_35 ();
 sg13g2_fill_2 FILLER_15_44 ();
 sg13g2_fill_2 FILLER_15_51 ();
 sg13g2_fill_1 FILLER_15_66 ();
 sg13g2_fill_1 FILLER_15_107 ();
 sg13g2_fill_2 FILLER_15_114 ();
 sg13g2_fill_2 FILLER_15_126 ();
 sg13g2_fill_1 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_132 ();
 sg13g2_fill_1 FILLER_15_146 ();
 sg13g2_fill_2 FILLER_15_155 ();
 sg13g2_decap_4 FILLER_15_161 ();
 sg13g2_fill_1 FILLER_15_177 ();
 sg13g2_fill_2 FILLER_15_201 ();
 sg13g2_fill_1 FILLER_15_206 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_fill_1 FILLER_15_258 ();
 sg13g2_fill_2 FILLER_15_263 ();
 sg13g2_decap_4 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_fill_2 FILLER_15_322 ();
 sg13g2_fill_1 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_329 ();
 sg13g2_fill_1 FILLER_15_334 ();
 sg13g2_fill_1 FILLER_15_343 ();
 sg13g2_fill_2 FILLER_15_353 ();
 sg13g2_fill_1 FILLER_15_355 ();
 sg13g2_fill_2 FILLER_15_370 ();
 sg13g2_fill_2 FILLER_15_394 ();
 sg13g2_fill_1 FILLER_15_396 ();
 sg13g2_fill_2 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_15_415 ();
 sg13g2_decap_8 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_fill_2 FILLER_16_133 ();
 sg13g2_fill_2 FILLER_16_197 ();
 sg13g2_fill_2 FILLER_16_220 ();
 sg13g2_fill_2 FILLER_16_228 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_263 ();
 sg13g2_fill_1 FILLER_16_268 ();
 sg13g2_fill_1 FILLER_16_274 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_346 ();
 sg13g2_fill_1 FILLER_16_348 ();
 sg13g2_fill_1 FILLER_16_374 ();
 sg13g2_decap_8 FILLER_16_404 ();
 sg13g2_decap_8 FILLER_16_411 ();
 sg13g2_decap_8 FILLER_16_418 ();
 sg13g2_decap_4 FILLER_16_425 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_fill_2 FILLER_17_33 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_44 ();
 sg13g2_decap_4 FILLER_17_50 ();
 sg13g2_fill_1 FILLER_17_91 ();
 sg13g2_fill_2 FILLER_17_99 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_206 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_236 ();
 sg13g2_fill_2 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_297 ();
 sg13g2_fill_1 FILLER_17_309 ();
 sg13g2_fill_1 FILLER_17_338 ();
 sg13g2_fill_2 FILLER_17_371 ();
 sg13g2_fill_2 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_fill_2 FILLER_18_12 ();
 sg13g2_fill_2 FILLER_18_22 ();
 sg13g2_fill_2 FILLER_18_32 ();
 sg13g2_fill_1 FILLER_18_34 ();
 sg13g2_fill_1 FILLER_18_41 ();
 sg13g2_fill_2 FILLER_18_47 ();
 sg13g2_decap_8 FILLER_18_61 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_fill_1 FILLER_18_84 ();
 sg13g2_fill_2 FILLER_18_92 ();
 sg13g2_fill_1 FILLER_18_99 ();
 sg13g2_fill_2 FILLER_18_106 ();
 sg13g2_fill_1 FILLER_18_117 ();
 sg13g2_fill_1 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_139 ();
 sg13g2_fill_1 FILLER_18_145 ();
 sg13g2_fill_2 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_fill_2 FILLER_18_245 ();
 sg13g2_fill_2 FILLER_18_252 ();
 sg13g2_fill_2 FILLER_18_270 ();
 sg13g2_fill_1 FILLER_18_272 ();
 sg13g2_fill_1 FILLER_18_281 ();
 sg13g2_fill_2 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_356 ();
 sg13g2_fill_1 FILLER_18_363 ();
 sg13g2_fill_2 FILLER_18_372 ();
 sg13g2_fill_1 FILLER_18_378 ();
 sg13g2_fill_2 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_423 ();
 sg13g2_fill_2 FILLER_19_38 ();
 sg13g2_fill_2 FILLER_19_45 ();
 sg13g2_fill_2 FILLER_19_95 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_141 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_fill_2 FILLER_19_151 ();
 sg13g2_fill_2 FILLER_19_157 ();
 sg13g2_fill_2 FILLER_19_163 ();
 sg13g2_fill_1 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_197 ();
 sg13g2_fill_2 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_259 ();
 sg13g2_fill_1 FILLER_19_265 ();
 sg13g2_fill_2 FILLER_19_270 ();
 sg13g2_fill_2 FILLER_19_276 ();
 sg13g2_fill_2 FILLER_19_283 ();
 sg13g2_fill_2 FILLER_19_330 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_fill_1 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_361 ();
 sg13g2_fill_1 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_408 ();
 sg13g2_fill_1 FILLER_19_415 ();
 sg13g2_decap_8 FILLER_19_421 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_11 ();
 sg13g2_fill_1 FILLER_20_15 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_fill_2 FILLER_20_44 ();
 sg13g2_fill_1 FILLER_20_46 ();
 sg13g2_decap_4 FILLER_20_83 ();
 sg13g2_fill_2 FILLER_20_87 ();
 sg13g2_fill_2 FILLER_20_94 ();
 sg13g2_fill_1 FILLER_20_96 ();
 sg13g2_fill_2 FILLER_20_102 ();
 sg13g2_fill_1 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_115 ();
 sg13g2_fill_1 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_200 ();
 sg13g2_fill_2 FILLER_20_206 ();
 sg13g2_fill_1 FILLER_20_213 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_fill_2 FILLER_20_232 ();
 sg13g2_fill_2 FILLER_20_262 ();
 sg13g2_fill_2 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_287 ();
 sg13g2_fill_1 FILLER_20_289 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_fill_1 FILLER_20_304 ();
 sg13g2_fill_2 FILLER_20_311 ();
 sg13g2_fill_2 FILLER_20_321 ();
 sg13g2_fill_1 FILLER_20_354 ();
 sg13g2_fill_2 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_366 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_fill_1 FILLER_20_401 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_21_45 ();
 sg13g2_fill_2 FILLER_21_52 ();
 sg13g2_fill_1 FILLER_21_64 ();
 sg13g2_fill_2 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_87 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_146 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_decap_4 FILLER_21_239 ();
 sg13g2_fill_1 FILLER_21_243 ();
 sg13g2_fill_1 FILLER_21_254 ();
 sg13g2_fill_2 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_265 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_decap_4 FILLER_21_306 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_1 FILLER_21_388 ();
 sg13g2_decap_8 FILLER_21_419 ();
 sg13g2_decap_4 FILLER_21_426 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_8 ();
 sg13g2_fill_2 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_76 ();
 sg13g2_fill_2 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_177 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_205 ();
 sg13g2_decap_4 FILLER_22_211 ();
 sg13g2_fill_2 FILLER_22_246 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_decap_4 FILLER_22_287 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_404 ();
 sg13g2_fill_2 FILLER_22_409 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_2 FILLER_23_33 ();
 sg13g2_fill_2 FILLER_23_100 ();
 sg13g2_fill_1 FILLER_23_188 ();
 sg13g2_decap_8 FILLER_23_215 ();
 sg13g2_fill_1 FILLER_23_222 ();
 sg13g2_decap_8 FILLER_23_227 ();
 sg13g2_decap_4 FILLER_23_234 ();
 sg13g2_fill_2 FILLER_23_238 ();
 sg13g2_fill_2 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_247 ();
 sg13g2_fill_2 FILLER_23_386 ();
 sg13g2_fill_1 FILLER_23_388 ();
 sg13g2_fill_2 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_2 FILLER_24_37 ();
 sg13g2_fill_1 FILLER_24_39 ();
 sg13g2_fill_1 FILLER_24_44 ();
 sg13g2_fill_1 FILLER_24_71 ();
 sg13g2_fill_1 FILLER_24_76 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_decap_8 FILLER_24_87 ();
 sg13g2_fill_1 FILLER_24_94 ();
 sg13g2_decap_4 FILLER_24_104 ();
 sg13g2_fill_1 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_fill_1 FILLER_24_128 ();
 sg13g2_decap_4 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_141 ();
 sg13g2_decap_4 FILLER_24_150 ();
 sg13g2_fill_2 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_fill_2 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_199 ();
 sg13g2_decap_4 FILLER_24_206 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_fill_1 FILLER_24_237 ();
 sg13g2_fill_1 FILLER_24_243 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_262 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_fill_1 FILLER_24_281 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_fill_1 FILLER_24_312 ();
 sg13g2_decap_4 FILLER_24_318 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_333 ();
 sg13g2_fill_2 FILLER_24_339 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_2 FILLER_24_395 ();
 sg13g2_fill_1 FILLER_24_397 ();
 sg13g2_fill_2 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_35 ();
 sg13g2_decap_4 FILLER_25_40 ();
 sg13g2_fill_2 FILLER_25_44 ();
 sg13g2_fill_2 FILLER_25_50 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_62 ();
 sg13g2_fill_2 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_74 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_121 ();
 sg13g2_fill_1 FILLER_25_148 ();
 sg13g2_fill_1 FILLER_25_154 ();
 sg13g2_fill_2 FILLER_25_159 ();
 sg13g2_fill_2 FILLER_25_217 ();
 sg13g2_fill_1 FILLER_25_219 ();
 sg13g2_decap_4 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_382 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_25_419 ();
 sg13g2_decap_4 FILLER_25_425 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_7 ();
 sg13g2_fill_1 FILLER_26_9 ();
 sg13g2_fill_1 FILLER_26_40 ();
 sg13g2_fill_2 FILLER_26_92 ();
 sg13g2_fill_2 FILLER_26_209 ();
 sg13g2_fill_2 FILLER_26_215 ();
 sg13g2_decap_4 FILLER_26_224 ();
 sg13g2_fill_2 FILLER_26_228 ();
 sg13g2_decap_4 FILLER_26_234 ();
 sg13g2_fill_2 FILLER_26_238 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_decap_4 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_298 ();
 sg13g2_fill_1 FILLER_26_307 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_2 FILLER_26_377 ();
 sg13g2_fill_1 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_18 ();
 sg13g2_decap_4 FILLER_27_29 ();
 sg13g2_fill_2 FILLER_27_84 ();
 sg13g2_fill_2 FILLER_27_111 ();
 sg13g2_fill_2 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_fill_2 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_fill_2 FILLER_27_181 ();
 sg13g2_fill_1 FILLER_27_183 ();
 sg13g2_fill_1 FILLER_27_188 ();
 sg13g2_fill_1 FILLER_27_194 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_245 ();
 sg13g2_fill_2 FILLER_27_251 ();
 sg13g2_fill_1 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_264 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_274 ();
 sg13g2_fill_1 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_fill_2 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_348 ();
 sg13g2_fill_1 FILLER_27_350 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_fill_1 FILLER_27_371 ();
 sg13g2_fill_2 FILLER_27_410 ();
 sg13g2_decap_8 FILLER_27_416 ();
 sg13g2_decap_8 FILLER_27_423 ();
 sg13g2_fill_2 FILLER_28_36 ();
 sg13g2_fill_1 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_66 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_fill_2 FILLER_28_82 ();
 sg13g2_fill_1 FILLER_28_84 ();
 sg13g2_fill_2 FILLER_28_90 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_fill_2 FILLER_28_113 ();
 sg13g2_fill_1 FILLER_28_141 ();
 sg13g2_fill_2 FILLER_28_183 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_decap_4 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_241 ();
 sg13g2_fill_1 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_273 ();
 sg13g2_fill_1 FILLER_28_300 ();
 sg13g2_fill_1 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_329 ();
 sg13g2_fill_1 FILLER_28_335 ();
 sg13g2_fill_2 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_11 ();
 sg13g2_fill_2 FILLER_29_18 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_57 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_fill_1 FILLER_29_74 ();
 sg13g2_fill_1 FILLER_29_90 ();
 sg13g2_fill_1 FILLER_29_95 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_137 ();
 sg13g2_fill_1 FILLER_29_147 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_208 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_decap_4 FILLER_29_281 ();
 sg13g2_fill_2 FILLER_29_312 ();
 sg13g2_fill_2 FILLER_29_331 ();
 sg13g2_fill_2 FILLER_29_337 ();
 sg13g2_fill_2 FILLER_29_368 ();
 sg13g2_fill_1 FILLER_29_384 ();
 sg13g2_decap_4 FILLER_29_416 ();
 sg13g2_decap_4 FILLER_29_425 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_54 ();
 sg13g2_fill_2 FILLER_30_64 ();
 sg13g2_fill_2 FILLER_30_92 ();
 sg13g2_fill_1 FILLER_30_113 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_132 ();
 sg13g2_fill_1 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_169 ();
 sg13g2_fill_2 FILLER_30_178 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_2 FILLER_30_192 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_276 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_296 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_decap_4 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_fill_2 FILLER_30_402 ();
 sg13g2_fill_1 FILLER_31_45 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_fill_1 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_178 ();
 sg13g2_fill_2 FILLER_31_188 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_276 ();
 sg13g2_fill_1 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_392 ();
 sg13g2_fill_1 FILLER_31_420 ();
 sg13g2_decap_4 FILLER_31_426 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_44 ();
 sg13g2_fill_2 FILLER_32_67 ();
 sg13g2_fill_1 FILLER_32_69 ();
 sg13g2_fill_1 FILLER_32_109 ();
 sg13g2_fill_2 FILLER_32_121 ();
 sg13g2_fill_1 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_155 ();
 sg13g2_fill_2 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_176 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_189 ();
 sg13g2_fill_2 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_218 ();
 sg13g2_fill_2 FILLER_32_224 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_decap_4 FILLER_32_240 ();
 sg13g2_fill_1 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_decap_4 FILLER_32_297 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_310 ();
 sg13g2_fill_1 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_fill_1 FILLER_32_331 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_32_367 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_fill_2 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_396 ();
 sg13g2_fill_2 FILLER_32_415 ();
 sg13g2_fill_1 FILLER_32_417 ();
 sg13g2_fill_1 FILLER_33_47 ();
 sg13g2_fill_2 FILLER_33_73 ();
 sg13g2_fill_1 FILLER_33_75 ();
 sg13g2_fill_1 FILLER_33_81 ();
 sg13g2_fill_2 FILLER_33_87 ();
 sg13g2_fill_2 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_122 ();
 sg13g2_fill_1 FILLER_33_149 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_decap_4 FILLER_33_254 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_fill_1 FILLER_33_272 ();
 sg13g2_fill_1 FILLER_33_277 ();
 sg13g2_fill_1 FILLER_33_286 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_4 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_315 ();
 sg13g2_fill_1 FILLER_33_320 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_333 ();
 sg13g2_decap_4 FILLER_33_348 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_386 ();
 sg13g2_fill_2 FILLER_34_44 ();
 sg13g2_fill_2 FILLER_34_61 ();
 sg13g2_fill_1 FILLER_34_67 ();
 sg13g2_fill_1 FILLER_34_92 ();
 sg13g2_fill_2 FILLER_34_106 ();
 sg13g2_fill_2 FILLER_34_160 ();
 sg13g2_decap_4 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_211 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_fill_1 FILLER_34_251 ();
 sg13g2_fill_1 FILLER_34_257 ();
 sg13g2_fill_2 FILLER_34_276 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_decap_4 FILLER_34_343 ();
 sg13g2_fill_2 FILLER_34_352 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_2 FILLER_35_41 ();
 sg13g2_fill_1 FILLER_35_89 ();
 sg13g2_fill_2 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_104 ();
 sg13g2_fill_2 FILLER_35_131 ();
 sg13g2_fill_2 FILLER_35_219 ();
 sg13g2_decap_4 FILLER_35_231 ();
 sg13g2_fill_2 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_245 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_decap_4 FILLER_35_308 ();
 sg13g2_fill_1 FILLER_35_321 ();
 sg13g2_fill_1 FILLER_35_327 ();
 sg13g2_fill_1 FILLER_35_332 ();
 sg13g2_fill_1 FILLER_35_341 ();
 sg13g2_fill_1 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_372 ();
 sg13g2_fill_1 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_fill_1 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_181 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_decap_4 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_232 ();
 sg13g2_fill_1 FILLER_36_238 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_fill_2 FILLER_36_310 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_344 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_fill_2 FILLER_36_376 ();
 sg13g2_fill_1 FILLER_36_383 ();
 sg13g2_fill_1 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_394 ();
 sg13g2_fill_2 FILLER_36_404 ();
 sg13g2_fill_1 FILLER_36_410 ();
 sg13g2_decap_8 FILLER_36_423 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_fill_1 FILLER_37_117 ();
 sg13g2_fill_2 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_293 ();
 sg13g2_fill_2 FILLER_37_347 ();
 sg13g2_fill_2 FILLER_37_353 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_fill_2 FILLER_37_390 ();
 sg13g2_fill_1 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_427 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_1 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_60 ();
 sg13g2_fill_2 FILLER_38_87 ();
 sg13g2_fill_1 FILLER_38_121 ();
 sg13g2_fill_2 FILLER_38_168 ();
 sg13g2_fill_2 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_302 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_fill_2 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_368 ();
 sg13g2_decap_4 FILLER_38_400 ();
endmodule
