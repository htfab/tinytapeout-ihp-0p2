module tt_um_dlmiles_muldiv8 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire clknet_0_clk;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire net168;
 wire net148;
 wire \muldiv.a0_0.GATE ;
 wire \muldiv.a0_0.Q ;
 wire \muldiv.a0_1.Q ;
 wire \muldiv.a0_2.Q ;
 wire \muldiv.a0_3.Q ;
 wire \muldiv.a0_4.Q ;
 wire \muldiv.a0_5.Q ;
 wire \muldiv.a0_6.Q ;
 wire \muldiv.a0_7.Q ;
 wire \muldiv.a1_0.GATE ;
 wire \muldiv.a1_0.Q ;
 wire \muldiv.a1_1.Q ;
 wire \muldiv.a1_2.Q ;
 wire \muldiv.a1_3.Q ;
 wire \muldiv.a1_4.Q ;
 wire \muldiv.a1_5.Q ;
 wire \muldiv.a1_6.Q ;
 wire \muldiv.a1_7.Q ;
 wire \muldiv.div2reg ;
 wire \muldiv.div8.io_edivzero ;
 wire \muldiv.negedgeReg_1.area_io_q ;
 wire \muldiv.regR[0] ;
 wire \muldiv.regR[10] ;
 wire \muldiv.regR[11] ;
 wire \muldiv.regR[12] ;
 wire \muldiv.regR[13] ;
 wire \muldiv.regR[14] ;
 wire \muldiv.regR[15] ;
 wire \muldiv.regR[1] ;
 wire \muldiv.regR[2] ;
 wire \muldiv.regR[3] ;
 wire \muldiv.regR[4] ;
 wire \muldiv.regR[5] ;
 wire \muldiv.regR[6] ;
 wire \muldiv.regR[7] ;
 wire \muldiv.regR[8] ;
 wire \muldiv.regR[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 _1806_ (.A(\muldiv.a1_0.Q ),
    .X(_1501_));
 sg13g2_inv_2 _1807_ (.Y(_1512_),
    .A(net118));
 sg13g2_buf_1 _1808_ (.A(_1512_),
    .X(_1523_));
 sg13g2_buf_2 _1809_ (.A(\muldiv.a0_0.Q ),
    .X(_1534_));
 sg13g2_inv_1 _1810_ (.Y(_1545_),
    .A(_1534_));
 sg13g2_buf_1 _1811_ (.A(_1545_),
    .X(_1556_));
 sg13g2_buf_1 _1812_ (.A(_1556_),
    .X(_1567_));
 sg13g2_buf_1 _1813_ (.A(_1567_),
    .X(_1577_));
 sg13g2_nor2_1 _1814_ (.A(net96),
    .B(net55),
    .Y(_1588_));
 sg13g2_buf_1 _1815_ (.A(uio_in[7]),
    .X(_1599_));
 sg13g2_buf_2 _1816_ (.A(\muldiv.a0_3.Q ),
    .X(_1610_));
 sg13g2_buf_1 _1817_ (.A(_1610_),
    .X(_1621_));
 sg13g2_buf_1 _1818_ (.A(net115),
    .X(_1632_));
 sg13g2_buf_1 _1819_ (.A(uio_in[6]),
    .X(_1643_));
 sg13g2_buf_8 _1820_ (.A(\muldiv.a0_7.Q ),
    .X(_1654_));
 sg13g2_and2_1 _1821_ (.A(_1643_),
    .B(_1654_),
    .X(_1665_));
 sg13g2_buf_8 _1822_ (.A(_1665_),
    .X(_1676_));
 sg13g2_buf_1 _1823_ (.A(_1676_),
    .X(_1687_));
 sg13g2_xnor2_1 _1824_ (.Y(_1698_),
    .A(net94),
    .B(net68));
 sg13g2_buf_1 _1825_ (.A(_1698_),
    .X(_1709_));
 sg13g2_buf_1 _1826_ (.A(net47),
    .X(_1720_));
 sg13g2_buf_2 _1827_ (.A(\muldiv.a0_5.Q ),
    .X(_1731_));
 sg13g2_inv_1 _1828_ (.Y(_1742_),
    .A(_1731_));
 sg13g2_buf_1 _1829_ (.A(_1742_),
    .X(_1753_));
 sg13g2_buf_1 _1830_ (.A(net68),
    .X(_1764_));
 sg13g2_xnor2_1 _1831_ (.Y(_1775_),
    .A(_1753_),
    .B(net54));
 sg13g2_buf_1 _1832_ (.A(_1643_),
    .X(_0020_));
 sg13g2_inv_1 _1833_ (.Y(_0031_),
    .A(net129));
 sg13g2_buf_1 _1834_ (.A(_0031_),
    .X(_0042_));
 sg13g2_buf_1 _1835_ (.A(_1654_),
    .X(_0053_));
 sg13g2_nand2_1 _1836_ (.Y(_0064_),
    .A(net120),
    .B(_0053_));
 sg13g2_buf_8 _1837_ (.A(\muldiv.a0_6.Q ),
    .X(_0075_));
 sg13g2_buf_1 _1838_ (.A(_0075_),
    .X(_0086_));
 sg13g2_xnor2_1 _1839_ (.Y(_0097_),
    .A(_0086_),
    .B(_1687_));
 sg13g2_buf_2 _1840_ (.A(_0097_),
    .X(_0108_));
 sg13g2_nand2_1 _1841_ (.Y(_0119_),
    .A(_0064_),
    .B(_0108_));
 sg13g2_buf_2 _1842_ (.A(_0119_),
    .X(_0130_));
 sg13g2_nor2_2 _1843_ (.A(_1775_),
    .B(_0130_),
    .Y(_0141_));
 sg13g2_buf_8 _1844_ (.A(\muldiv.a1_3.Q ),
    .X(_0152_));
 sg13g2_buf_2 _1845_ (.A(\muldiv.a1_2.Q ),
    .X(_0163_));
 sg13g2_inv_1 _1846_ (.Y(_0174_),
    .A(_0163_));
 sg13g2_buf_2 _1847_ (.A(\muldiv.a1_1.Q ),
    .X(_0185_));
 sg13g2_nor2_1 _1848_ (.A(net118),
    .B(_0185_),
    .Y(_0196_));
 sg13g2_buf_2 _1849_ (.A(\muldiv.a1_7.Q ),
    .X(_0207_));
 sg13g2_nand2_1 _1850_ (.Y(_0218_),
    .A(_1643_),
    .B(_0207_));
 sg13g2_buf_2 _1851_ (.A(_0218_),
    .X(_0229_));
 sg13g2_buf_1 _1852_ (.A(_0229_),
    .X(_0240_));
 sg13g2_a21oi_1 _1853_ (.A1(_0174_),
    .A2(_0196_),
    .Y(_0251_),
    .B1(net67));
 sg13g2_xnor2_1 _1854_ (.Y(_0262_),
    .A(net117),
    .B(_0251_));
 sg13g2_buf_2 _1855_ (.A(_0262_),
    .X(_0273_));
 sg13g2_nor2_1 _1856_ (.A(net95),
    .B(_0273_),
    .Y(_0284_));
 sg13g2_xnor2_1 _1857_ (.Y(_0295_),
    .A(\muldiv.a0_2.Q ),
    .B(_1676_));
 sg13g2_buf_1 _1858_ (.A(_0295_),
    .X(_0306_));
 sg13g2_buf_2 _1859_ (.A(\muldiv.a1_6.Q ),
    .X(_0317_));
 sg13g2_nand2b_1 _1860_ (.Y(_0328_),
    .B(_0207_),
    .A_N(_0317_));
 sg13g2_buf_2 _1861_ (.A(\muldiv.a0_1.Q ),
    .X(_0339_));
 sg13g2_buf_8 _1862_ (.A(_0339_),
    .X(_0350_));
 sg13g2_nand2_1 _1863_ (.Y(_0361_),
    .A(_1534_),
    .B(net112));
 sg13g2_buf_2 _1864_ (.A(_0361_),
    .X(_0372_));
 sg13g2_nor2_1 _1865_ (.A(_0328_),
    .B(_0372_),
    .Y(_0383_));
 sg13g2_inv_2 _1866_ (.Y(_0394_),
    .A(_1610_));
 sg13g2_buf_2 _1867_ (.A(\muldiv.a0_4.Q ),
    .X(_0405_));
 sg13g2_nor4_2 _1868_ (.A(_1654_),
    .B(_0075_),
    .C(_1731_),
    .Y(_0416_),
    .D(_0405_));
 sg13g2_and4_1 _1869_ (.A(_0075_),
    .B(_1731_),
    .C(_0405_),
    .D(_1610_),
    .X(_0427_));
 sg13g2_a22oi_1 _1870_ (.Y(_0438_),
    .B1(_0427_),
    .B2(_1676_),
    .A2(_0416_),
    .A1(_0394_));
 sg13g2_buf_2 _1871_ (.A(_0438_),
    .X(_0449_));
 sg13g2_inv_2 _1872_ (.Y(_0460_),
    .A(_0339_));
 sg13g2_nand2_1 _1873_ (.Y(_0471_),
    .A(_1545_),
    .B(net111));
 sg13g2_nand3b_1 _1874_ (.B(_0471_),
    .C(_0295_),
    .Y(_0482_),
    .A_N(_0449_));
 sg13g2_inv_1 _1875_ (.Y(_0493_),
    .A(_0317_));
 sg13g2_nor4_2 _1876_ (.A(_1501_),
    .B(_0152_),
    .C(_0163_),
    .Y(_0503_),
    .D(_0185_));
 sg13g2_buf_2 _1877_ (.A(\muldiv.a1_5.Q ),
    .X(_0514_));
 sg13g2_buf_1 _1878_ (.A(\muldiv.a1_4.Q ),
    .X(_0525_));
 sg13g2_nor2_2 _1879_ (.A(_0514_),
    .B(_0525_),
    .Y(_0536_));
 sg13g2_nand3_1 _1880_ (.B(_0503_),
    .C(_0536_),
    .A(net110),
    .Y(_0547_));
 sg13g2_inv_1 _1881_ (.Y(_0557_),
    .A(_0207_));
 sg13g2_a21oi_1 _1882_ (.A1(net129),
    .A2(_0547_),
    .Y(_0568_),
    .B1(_0557_));
 sg13g2_nand3b_1 _1883_ (.B(_1654_),
    .C(_0020_),
    .Y(_0579_),
    .A_N(net112));
 sg13g2_or2_1 _1884_ (.X(_0590_),
    .B(_0579_),
    .A(_0328_));
 sg13g2_buf_1 _1885_ (.A(_0207_),
    .X(_0601_));
 sg13g2_inv_1 _1886_ (.Y(_0611_),
    .A(_1654_));
 sg13g2_and2_1 _1887_ (.A(_1534_),
    .B(net112),
    .X(_0622_));
 sg13g2_nand4_1 _1888_ (.B(_0611_),
    .C(net110),
    .A(net109),
    .Y(_0633_),
    .D(_0622_));
 sg13g2_buf_8 _1889_ (.A(_0503_),
    .X(_0644_));
 sg13g2_nand2_1 _1890_ (.Y(_0654_),
    .A(net92),
    .B(_0536_));
 sg13g2_a21oi_1 _1891_ (.A1(_0590_),
    .A2(_0633_),
    .Y(_0665_),
    .B1(_0654_));
 sg13g2_a221oi_1 _1892_ (.B2(_0568_),
    .C1(_0665_),
    .B1(_0482_),
    .A1(_0031_),
    .Y(_0675_),
    .A2(_0383_));
 sg13g2_buf_2 _1893_ (.A(_0675_),
    .X(_0686_));
 sg13g2_a21oi_1 _1894_ (.A1(net92),
    .A2(_0536_),
    .Y(_0697_),
    .B1(_0229_));
 sg13g2_xnor2_1 _1895_ (.Y(_0707_),
    .A(net110),
    .B(_0697_));
 sg13g2_nand2_1 _1896_ (.Y(_0718_),
    .A(_1643_),
    .B(_1654_));
 sg13g2_buf_2 _1897_ (.A(_0718_),
    .X(_0728_));
 sg13g2_nor2_2 _1898_ (.A(_0350_),
    .B(_0728_),
    .Y(_0739_));
 sg13g2_nand2_1 _1899_ (.Y(_0750_),
    .A(net95),
    .B(_0739_));
 sg13g2_and3_1 _1900_ (.X(_0761_),
    .A(_1534_),
    .B(_1643_),
    .C(_1654_));
 sg13g2_nor2b_1 _1901_ (.A(_1610_),
    .B_N(_1534_),
    .Y(_0771_));
 sg13g2_a22oi_1 _1902_ (.Y(_0782_),
    .B1(_0771_),
    .B2(_0416_),
    .A2(_0761_),
    .A1(_0427_));
 sg13g2_buf_1 _1903_ (.A(_0782_),
    .X(_0793_));
 sg13g2_nand2b_1 _1904_ (.Y(_0803_),
    .B(_0295_),
    .A_N(_0793_));
 sg13g2_buf_8 _1905_ (.A(_1534_),
    .X(_0814_));
 sg13g2_xnor2_1 _1906_ (.Y(_0825_),
    .A(net111),
    .B(_1676_));
 sg13g2_buf_1 _1907_ (.A(_0825_),
    .X(_0836_));
 sg13g2_nor2b_1 _1908_ (.A(_0525_),
    .B_N(_0514_),
    .Y(_0846_));
 sg13g2_a22oi_1 _1909_ (.Y(_0856_),
    .B1(_0846_),
    .B2(net92),
    .A2(_0229_),
    .A1(_0514_));
 sg13g2_buf_1 _1910_ (.A(_0856_),
    .X(_0867_));
 sg13g2_inv_2 _1911_ (.Y(_0878_),
    .A(_0525_));
 sg13g2_nand3b_1 _1912_ (.B(_0207_),
    .C(_1643_),
    .Y(_0889_),
    .A_N(_0514_));
 sg13g2_a21o_1 _1913_ (.A2(_0503_),
    .A1(_0878_),
    .B1(_0889_),
    .X(_0899_));
 sg13g2_buf_8 _1914_ (.A(_0899_),
    .X(_0910_));
 sg13g2_nand4_1 _1915_ (.B(_0836_),
    .C(_0867_),
    .A(net107),
    .Y(_0919_),
    .D(_0910_));
 sg13g2_nand4_1 _1916_ (.B(_0750_),
    .C(_0803_),
    .A(_0707_),
    .Y(_0923_),
    .D(_0919_));
 sg13g2_buf_2 _1917_ (.A(_0923_),
    .X(_0931_));
 sg13g2_nand3_1 _1918_ (.B(_0867_),
    .C(_0910_),
    .A(net107),
    .Y(_0939_));
 sg13g2_nand2_2 _1919_ (.Y(_0948_),
    .A(net95),
    .B(_1676_));
 sg13g2_nand3b_1 _1920_ (.B(_0207_),
    .C(net129),
    .Y(_0949_),
    .A_N(_0317_));
 sg13g2_a21o_1 _1921_ (.A2(_0536_),
    .A1(net92),
    .B1(_0949_),
    .X(_0950_));
 sg13g2_buf_1 _1922_ (.A(_0317_),
    .X(_0951_));
 sg13g2_nand2_1 _1923_ (.Y(_0952_),
    .A(_0557_),
    .B(net106));
 sg13g2_nand4_1 _1924_ (.B(_0317_),
    .C(_0644_),
    .A(net129),
    .Y(_0953_),
    .D(_0536_));
 sg13g2_nand4_1 _1925_ (.B(net52),
    .C(_0952_),
    .A(_0950_),
    .Y(_0954_),
    .D(_0953_));
 sg13g2_nand3_1 _1926_ (.B(_0948_),
    .C(_0954_),
    .A(_0939_),
    .Y(_0955_));
 sg13g2_buf_1 _1927_ (.A(_0955_),
    .X(_0956_));
 sg13g2_nand3_1 _1928_ (.B(_0931_),
    .C(_0956_),
    .A(_0686_),
    .Y(_0957_));
 sg13g2_buf_1 _1929_ (.A(_0957_),
    .X(_0958_));
 sg13g2_and3_1 _1930_ (.X(_0959_),
    .A(net107),
    .B(_0867_),
    .C(_0910_));
 sg13g2_nor2_1 _1931_ (.A(net107),
    .B(_0728_),
    .Y(_0960_));
 sg13g2_nor2_1 _1932_ (.A(_0449_),
    .B(net52),
    .Y(_0961_));
 sg13g2_o21ai_1 _1933_ (.B1(_0961_),
    .Y(_0962_),
    .A1(_0959_),
    .A2(_0960_));
 sg13g2_xnor2_1 _1934_ (.Y(_0963_),
    .A(_0394_),
    .B(_1676_));
 sg13g2_buf_1 _1935_ (.A(_0963_),
    .X(_0964_));
 sg13g2_and4_1 _1936_ (.A(net129),
    .B(net114),
    .C(_0075_),
    .D(_0405_),
    .X(_0965_));
 sg13g2_a21oi_2 _1937_ (.B1(_0416_),
    .Y(_0966_),
    .A2(_0965_),
    .A1(_1731_));
 sg13g2_nor2_1 _1938_ (.A(net51),
    .B(_0966_),
    .Y(_0967_));
 sg13g2_nand4_1 _1939_ (.B(net52),
    .C(_0939_),
    .A(_0967_),
    .Y(_0968_),
    .D(_0948_));
 sg13g2_nand2_2 _1940_ (.Y(_0969_),
    .A(_0962_),
    .B(_0968_));
 sg13g2_buf_8 _1941_ (.A(net107),
    .X(_0970_));
 sg13g2_buf_1 _1942_ (.A(_0525_),
    .X(_0971_));
 sg13g2_or4_1 _1943_ (.A(_1501_),
    .B(_0152_),
    .C(_0163_),
    .D(_0185_),
    .X(_0972_));
 sg13g2_nor4_2 _1944_ (.A(_0317_),
    .B(_0514_),
    .C(_0971_),
    .Y(_0973_),
    .D(_0972_));
 sg13g2_o21ai_1 _1945_ (.B1(net109),
    .Y(_0974_),
    .A1(_0031_),
    .A2(_0973_));
 sg13g2_buf_1 _1946_ (.A(_0974_),
    .X(_0975_));
 sg13g2_nand2b_1 _1947_ (.Y(_0976_),
    .B(_0295_),
    .A_N(_0449_));
 sg13g2_a21oi_2 _1948_ (.B1(_0976_),
    .Y(_0977_),
    .A2(_0975_),
    .A1(net52));
 sg13g2_xnor2_1 _1949_ (.Y(_0978_),
    .A(net106),
    .B(_0697_));
 sg13g2_a21o_1 _1950_ (.A2(_0977_),
    .A1(net91),
    .B1(_0978_),
    .X(_0979_));
 sg13g2_buf_2 _1951_ (.A(_0979_),
    .X(_0980_));
 sg13g2_a21o_1 _1952_ (.A2(_0969_),
    .A1(_0958_),
    .B1(_0980_),
    .X(_0981_));
 sg13g2_nand3_1 _1953_ (.B(_0958_),
    .C(_0969_),
    .A(_0980_),
    .Y(_0982_));
 sg13g2_a21oi_1 _1954_ (.A1(net51),
    .A2(_0686_),
    .Y(_0983_),
    .B1(_0966_));
 sg13g2_nand2_1 _1955_ (.Y(_0984_),
    .A(net53),
    .B(_0983_));
 sg13g2_a21oi_2 _1956_ (.B1(_0984_),
    .Y(_0985_),
    .A2(_0982_),
    .A1(_0981_));
 sg13g2_buf_1 _1957_ (.A(\muldiv.a0_2.Q ),
    .X(_0986_));
 sg13g2_inv_1 _1958_ (.Y(_0987_),
    .A(net116));
 sg13g2_xnor2_1 _1959_ (.Y(_0988_),
    .A(_0987_),
    .B(_1676_));
 sg13g2_buf_2 _1960_ (.A(_0988_),
    .X(_0989_));
 sg13g2_a21oi_1 _1961_ (.A1(_0931_),
    .A2(_0956_),
    .Y(_0990_),
    .B1(_0989_));
 sg13g2_and4_1 _1962_ (.A(_0707_),
    .B(_0750_),
    .C(_0803_),
    .D(_0919_),
    .X(_0991_));
 sg13g2_and3_1 _1963_ (.X(_0992_),
    .A(_0939_),
    .B(_0948_),
    .C(_0954_));
 sg13g2_nor3_1 _1964_ (.A(_0306_),
    .B(_0991_),
    .C(_0992_),
    .Y(_0993_));
 sg13g2_nor2_1 _1965_ (.A(_0990_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_nor2_1 _1966_ (.A(_0449_),
    .B(_0686_),
    .Y(_0995_));
 sg13g2_nor2b_1 _1967_ (.A(_0994_),
    .B_N(_0995_),
    .Y(_0996_));
 sg13g2_buf_1 _1968_ (.A(_0996_),
    .X(_0997_));
 sg13g2_nand2b_1 _1969_ (.Y(_0998_),
    .B(_0306_),
    .A_N(_0686_));
 sg13g2_buf_8 _1970_ (.A(_0998_),
    .X(_0999_));
 sg13g2_nand2_1 _1971_ (.Y(_1000_),
    .A(_0989_),
    .B(_0975_));
 sg13g2_o21ai_1 _1972_ (.B1(_1000_),
    .Y(_1001_),
    .A1(_0991_),
    .A2(_0992_));
 sg13g2_buf_2 _1973_ (.A(_1001_),
    .X(_1002_));
 sg13g2_nand2_1 _1974_ (.Y(_1003_),
    .A(_0878_),
    .B(_0644_));
 sg13g2_inv_1 _1975_ (.Y(_1004_),
    .A(_0793_));
 sg13g2_nand2b_1 _1976_ (.Y(_1005_),
    .B(_0514_),
    .A_N(_0971_));
 sg13g2_nand2b_1 _1977_ (.Y(_1006_),
    .B(net112),
    .A_N(_0053_));
 sg13g2_o21ai_1 _1978_ (.B1(_1006_),
    .Y(_1007_),
    .A1(net109),
    .A2(_1005_));
 sg13g2_buf_1 _1979_ (.A(_0514_),
    .X(_1008_));
 sg13g2_nor4_1 _1980_ (.A(_1008_),
    .B(_0878_),
    .C(net92),
    .D(_0229_),
    .Y(_1009_));
 sg13g2_a21oi_1 _1981_ (.A1(net111),
    .A2(_1005_),
    .Y(_1010_),
    .B1(net129));
 sg13g2_nor4_1 _1982_ (.A(_0739_),
    .B(_1007_),
    .C(_1009_),
    .D(_1010_),
    .Y(_1011_));
 sg13g2_nand3_1 _1983_ (.B(_1004_),
    .C(_1011_),
    .A(_1003_),
    .Y(_1012_));
 sg13g2_xnor2_1 _1984_ (.Y(_1013_),
    .A(_0350_),
    .B(_1676_));
 sg13g2_buf_1 _1985_ (.A(_1013_),
    .X(_1014_));
 sg13g2_nor3_1 _1986_ (.A(_0814_),
    .B(_0728_),
    .C(_0229_),
    .Y(_1015_));
 sg13g2_nor4_1 _1987_ (.A(_1556_),
    .B(_0878_),
    .C(net92),
    .D(_0229_),
    .Y(_1016_));
 sg13g2_a21oi_1 _1988_ (.A1(_1003_),
    .A2(_1015_),
    .Y(_1017_),
    .B1(_1016_));
 sg13g2_nand4_1 _1989_ (.B(net50),
    .C(_0793_),
    .A(_1008_),
    .Y(_1018_),
    .D(_1017_));
 sg13g2_inv_1 _1990_ (.Y(_1019_),
    .A(net104));
 sg13g2_nor2_1 _1991_ (.A(net92),
    .B(_0229_),
    .Y(_1020_));
 sg13g2_o21ai_1 _1992_ (.B1(net105),
    .Y(_1021_),
    .A1(_0814_),
    .A2(net109));
 sg13g2_o21ai_1 _1993_ (.B1(_1021_),
    .Y(_1022_),
    .A1(net107),
    .A2(net68));
 sg13g2_or2_1 _1994_ (.X(_1023_),
    .B(_1022_),
    .A(_1020_));
 sg13g2_nand4_1 _1995_ (.B(net50),
    .C(_0793_),
    .A(_1019_),
    .Y(_1024_),
    .D(_1023_));
 sg13g2_nand3_1 _1996_ (.B(_1004_),
    .C(_1011_),
    .A(_1019_),
    .Y(_1025_));
 sg13g2_and4_1 _1997_ (.A(_1012_),
    .B(_1018_),
    .C(_1024_),
    .D(_1025_),
    .X(_1026_));
 sg13g2_a21o_1 _1998_ (.A2(_1002_),
    .A1(_0999_),
    .B1(_1026_),
    .X(_1027_));
 sg13g2_mux2_1 _1999_ (.A0(_1017_),
    .A1(_1023_),
    .S(_1019_),
    .X(_1028_));
 sg13g2_nand4_1 _2000_ (.B(_0999_),
    .C(_1002_),
    .A(_1014_),
    .Y(_1029_),
    .D(_1028_));
 sg13g2_nand2_1 _2001_ (.Y(_1030_),
    .A(_0989_),
    .B(_0568_));
 sg13g2_a221oi_1 _2002_ (.B2(_0968_),
    .C1(_1030_),
    .B1(_0962_),
    .A1(_0931_),
    .Y(_1031_),
    .A2(_0956_));
 sg13g2_nand2_1 _2003_ (.Y(_1032_),
    .A(_0978_),
    .B(_0989_));
 sg13g2_nand3b_1 _2004_ (.B(_1032_),
    .C(_0983_),
    .Y(_1033_),
    .A_N(_1031_));
 sg13g2_buf_1 _2005_ (.A(_1033_),
    .X(_1034_));
 sg13g2_a21oi_1 _2006_ (.A1(_1027_),
    .A2(_1029_),
    .Y(_1035_),
    .B1(_1034_));
 sg13g2_or3_1 _2007_ (.A(_0985_),
    .B(_0997_),
    .C(_1035_),
    .X(_1036_));
 sg13g2_xnor2_1 _2008_ (.Y(_1037_),
    .A(net105),
    .B(_1020_));
 sg13g2_buf_1 _2009_ (.A(_1037_),
    .X(_1038_));
 sg13g2_a21oi_1 _2010_ (.A1(net91),
    .A2(_1038_),
    .Y(_1039_),
    .B1(_0960_));
 sg13g2_and2_1 _2011_ (.A(_0867_),
    .B(_0910_),
    .X(_1040_));
 sg13g2_nand4_1 _2012_ (.B(_1040_),
    .C(_0931_),
    .A(_0686_),
    .Y(_1041_),
    .D(_0956_));
 sg13g2_and2_1 _2013_ (.A(_0989_),
    .B(_1040_),
    .X(_1042_));
 sg13g2_nand3_1 _2014_ (.B(_0956_),
    .C(_1042_),
    .A(_0931_),
    .Y(_1043_));
 sg13g2_a22oi_1 _2015_ (.Y(_1044_),
    .B1(_1042_),
    .B2(_0686_),
    .A2(_1040_),
    .A1(_0793_));
 sg13g2_nand3_1 _2016_ (.B(_1043_),
    .C(_1044_),
    .A(_1041_),
    .Y(_1045_));
 sg13g2_a221oi_1 _2017_ (.B2(_1002_),
    .C1(_0793_),
    .B1(_0999_),
    .A1(_0867_),
    .Y(_1046_),
    .A2(_0910_));
 sg13g2_or2_1 _2018_ (.X(_1047_),
    .B(_1046_),
    .A(_1045_));
 sg13g2_buf_1 _2019_ (.A(_1047_),
    .X(_1048_));
 sg13g2_nor3_1 _2020_ (.A(net52),
    .B(_1039_),
    .C(_1048_),
    .Y(_1049_));
 sg13g2_xnor2_1 _2021_ (.Y(_1050_),
    .A(_0878_),
    .B(_1020_));
 sg13g2_o21ai_1 _2022_ (.B1(_0948_),
    .Y(_1051_),
    .A1(net95),
    .A2(_1050_));
 sg13g2_buf_1 _2023_ (.A(_1051_),
    .X(_1052_));
 sg13g2_o21ai_1 _2024_ (.B1(_0995_),
    .Y(_1053_),
    .A1(_0990_),
    .A2(_0993_));
 sg13g2_buf_1 _2025_ (.A(_1053_),
    .X(_1054_));
 sg13g2_and2_1 _2026_ (.A(_1054_),
    .B(_1034_),
    .X(_1055_));
 sg13g2_nor4_1 _2027_ (.A(net50),
    .B(_1052_),
    .C(_1048_),
    .D(_1055_),
    .Y(_1056_));
 sg13g2_a21oi_1 _2028_ (.A1(_1036_),
    .A2(_1049_),
    .Y(_1057_),
    .B1(_1056_));
 sg13g2_nor3_1 _2029_ (.A(_0985_),
    .B(_0997_),
    .C(_1035_),
    .Y(_1058_));
 sg13g2_nand2_1 _2030_ (.Y(_1059_),
    .A(net52),
    .B(_1052_));
 sg13g2_nand2_1 _2031_ (.Y(_1060_),
    .A(net50),
    .B(_1039_));
 sg13g2_nor2_1 _2032_ (.A(_1045_),
    .B(_1046_),
    .Y(_1061_));
 sg13g2_a21oi_1 _2033_ (.A1(_1059_),
    .A2(_1060_),
    .Y(_1062_),
    .B1(_1061_));
 sg13g2_a21oi_1 _2034_ (.A1(_1058_),
    .A2(_1048_),
    .Y(_1063_),
    .B1(_1062_));
 sg13g2_and2_1 _2035_ (.A(_1057_),
    .B(_1063_),
    .X(_1064_));
 sg13g2_buf_2 _2036_ (.A(_1064_),
    .X(_1065_));
 sg13g2_nand2_1 _2037_ (.Y(_1066_),
    .A(net91),
    .B(_0273_));
 sg13g2_inv_1 _2038_ (.Y(_1067_),
    .A(_1066_));
 sg13g2_nand2_1 _2039_ (.Y(_1068_),
    .A(_1050_),
    .B(_1067_));
 sg13g2_a21o_1 _2040_ (.A2(_0982_),
    .A1(_0981_),
    .B1(_0984_),
    .X(_1069_));
 sg13g2_nand4_1 _2041_ (.B(_1054_),
    .C(net46),
    .A(_1069_),
    .Y(_1070_),
    .D(_1067_));
 sg13g2_nor2_1 _2042_ (.A(_1034_),
    .B(_1052_),
    .Y(_1071_));
 sg13g2_a21oi_2 _2043_ (.B1(_1035_),
    .Y(_1072_),
    .A2(_1071_),
    .A1(_1061_));
 sg13g2_mux2_1 _2044_ (.A0(_1068_),
    .A1(_1070_),
    .S(_1072_),
    .X(_1073_));
 sg13g2_buf_1 _2045_ (.A(_1073_),
    .X(_1074_));
 sg13g2_nor3_1 _2046_ (.A(_0985_),
    .B(_0997_),
    .C(_0273_),
    .Y(_1075_));
 sg13g2_o21ai_1 _2047_ (.B1(_0579_),
    .Y(_1076_),
    .A1(net68),
    .A2(_0372_));
 sg13g2_o21ai_1 _2048_ (.B1(_1076_),
    .Y(_1077_),
    .A1(_1050_),
    .A2(_0273_));
 sg13g2_a21o_1 _2049_ (.A2(_1075_),
    .A1(_1072_),
    .B1(_1077_),
    .X(_1078_));
 sg13g2_nand2_1 _2050_ (.Y(_1079_),
    .A(_1069_),
    .B(_1054_));
 sg13g2_nor2_1 _2051_ (.A(net46),
    .B(_1066_),
    .Y(_1080_));
 sg13g2_nor4_1 _2052_ (.A(net50),
    .B(_0985_),
    .C(_0997_),
    .D(_1050_),
    .Y(_1081_));
 sg13g2_buf_8 _2053_ (.A(net112),
    .X(_1082_));
 sg13g2_a21oi_1 _2054_ (.A1(net90),
    .A2(net46),
    .Y(_1083_),
    .B1(_0739_));
 sg13g2_nor2_1 _2055_ (.A(net91),
    .B(_1083_),
    .Y(_1084_));
 sg13g2_a221oi_1 _2056_ (.B2(_1072_),
    .C1(_1084_),
    .B1(_1081_),
    .A1(_1079_),
    .Y(_1085_),
    .A2(_1080_));
 sg13g2_and4_1 _2057_ (.A(_1057_),
    .B(_1063_),
    .C(_1078_),
    .D(_1085_),
    .X(_1086_));
 sg13g2_and4_1 _2058_ (.A(net53),
    .B(_1078_),
    .C(_1074_),
    .D(_1085_),
    .X(_1087_));
 sg13g2_a221oi_1 _2059_ (.B2(_1086_),
    .C1(_1087_),
    .B1(_1074_),
    .A1(net53),
    .Y(_1088_),
    .A2(_1065_));
 sg13g2_buf_2 _2060_ (.A(_1088_),
    .X(_1089_));
 sg13g2_inv_1 _2061_ (.Y(_1090_),
    .A(_0405_));
 sg13g2_xnor2_1 _2062_ (.Y(_1091_),
    .A(_1090_),
    .B(net68));
 sg13g2_buf_1 _2063_ (.A(_1091_),
    .X(_1092_));
 sg13g2_a21o_1 _2064_ (.A2(_0994_),
    .A1(_0967_),
    .B1(_0686_),
    .X(_1093_));
 sg13g2_nand2_1 _2065_ (.Y(_1094_),
    .A(net45),
    .B(_1093_));
 sg13g2_a21oi_1 _2066_ (.A1(_1069_),
    .A2(_1054_),
    .Y(_1095_),
    .B1(_0989_));
 sg13g2_nor2_1 _2067_ (.A(net53),
    .B(_1055_),
    .Y(_1096_));
 sg13g2_nand2_1 _2068_ (.Y(_1097_),
    .A(_1027_),
    .B(_1029_));
 sg13g2_a21o_1 _2069_ (.A2(_1061_),
    .A1(_1039_),
    .B1(_1097_),
    .X(_1098_));
 sg13g2_mux2_1 _2070_ (.A0(_1095_),
    .A1(_1096_),
    .S(_1098_),
    .X(_1099_));
 sg13g2_o21ai_1 _2071_ (.B1(net51),
    .Y(_1100_),
    .A1(_0980_),
    .A2(_1099_));
 sg13g2_nand2_1 _2072_ (.Y(_1101_),
    .A(_1094_),
    .B(_1100_));
 sg13g2_buf_1 _2073_ (.A(net91),
    .X(_1102_));
 sg13g2_a21oi_1 _2074_ (.A1(net66),
    .A2(_0977_),
    .Y(_1103_),
    .B1(_0978_));
 sg13g2_nand2_1 _2075_ (.Y(_1104_),
    .A(_0999_),
    .B(_1002_));
 sg13g2_nand2_1 _2076_ (.Y(_1105_),
    .A(_0969_),
    .B(_1104_));
 sg13g2_inv_1 _2077_ (.Y(_1106_),
    .A(_1105_));
 sg13g2_nor3_1 _2078_ (.A(net51),
    .B(_1103_),
    .C(_1106_),
    .Y(_1107_));
 sg13g2_nor3_1 _2079_ (.A(_0964_),
    .B(_0980_),
    .C(_1106_),
    .Y(_1108_));
 sg13g2_o21ai_1 _2080_ (.B1(net53),
    .Y(_1109_),
    .A1(_0985_),
    .A2(_0997_));
 sg13g2_or2_1 _2081_ (.X(_1110_),
    .B(_1055_),
    .A(net53));
 sg13g2_mux2_1 _2082_ (.A0(_1109_),
    .A1(_1110_),
    .S(_1098_),
    .X(_1111_));
 sg13g2_mux2_1 _2083_ (.A0(_1107_),
    .A1(_1108_),
    .S(_1111_),
    .X(_1112_));
 sg13g2_buf_1 _2084_ (.A(_1112_),
    .X(_1113_));
 sg13g2_a21oi_1 _2085_ (.A1(_0958_),
    .A2(_0969_),
    .Y(_1114_),
    .B1(_0980_));
 sg13g2_and3_1 _2086_ (.X(_1115_),
    .A(_0980_),
    .B(_0958_),
    .C(_0969_));
 sg13g2_nor3_1 _2087_ (.A(net47),
    .B(_0989_),
    .C(_0966_),
    .Y(_1116_));
 sg13g2_o21ai_1 _2088_ (.B1(_1116_),
    .Y(_1117_),
    .A1(_1114_),
    .A2(_1115_));
 sg13g2_nor2b_1 _2089_ (.A(_1093_),
    .B_N(_1117_),
    .Y(_1118_));
 sg13g2_o21ai_1 _2090_ (.B1(net53),
    .Y(_1119_),
    .A1(_1114_),
    .A2(_1115_));
 sg13g2_nand2b_1 _2091_ (.Y(_1120_),
    .B(_1032_),
    .A_N(_1031_));
 sg13g2_or4_1 _2092_ (.A(_1120_),
    .B(_1052_),
    .C(_1045_),
    .D(_1046_),
    .X(_1121_));
 sg13g2_a21o_1 _2093_ (.A2(_1029_),
    .A1(_1027_),
    .B1(_1120_),
    .X(_1122_));
 sg13g2_nand4_1 _2094_ (.B(_1119_),
    .C(_1121_),
    .A(_0967_),
    .Y(_1123_),
    .D(_1122_));
 sg13g2_buf_1 _2095_ (.A(_1731_),
    .X(_1124_));
 sg13g2_xnor2_1 _2096_ (.Y(_1125_),
    .A(_1124_),
    .B(_1687_));
 sg13g2_buf_1 _2097_ (.A(_1125_),
    .X(_1126_));
 sg13g2_nor2_1 _2098_ (.A(_0020_),
    .B(net108),
    .Y(_1127_));
 sg13g2_buf_1 _2099_ (.A(_1127_),
    .X(_1128_));
 sg13g2_inv_2 _2100_ (.Y(_1129_),
    .A(_0075_));
 sg13g2_xnor2_1 _2101_ (.Y(_1130_),
    .A(_1129_),
    .B(net68));
 sg13g2_buf_1 _2102_ (.A(_1130_),
    .X(_1131_));
 sg13g2_nor2_1 _2103_ (.A(net65),
    .B(net44),
    .Y(_1132_));
 sg13g2_nand2_1 _2104_ (.Y(_1133_),
    .A(_1126_),
    .B(_1132_));
 sg13g2_buf_2 _2105_ (.A(_1133_),
    .X(_1134_));
 sg13g2_nor2_1 _2106_ (.A(net45),
    .B(_1134_),
    .Y(_1135_));
 sg13g2_nand2_1 _2107_ (.Y(_1136_),
    .A(net51),
    .B(_1135_));
 sg13g2_a21o_1 _2108_ (.A2(_1122_),
    .A1(_1121_),
    .B1(_1136_),
    .X(_1137_));
 sg13g2_nand3_1 _2109_ (.B(_1123_),
    .C(_1137_),
    .A(_1118_),
    .Y(_1138_));
 sg13g2_buf_2 _2110_ (.A(_1138_),
    .X(_1139_));
 sg13g2_nor2_1 _2111_ (.A(net45),
    .B(_1139_),
    .Y(_1140_));
 sg13g2_a21oi_1 _2112_ (.A1(_1113_),
    .A2(_1094_),
    .Y(_1141_),
    .B1(_1140_));
 sg13g2_o21ai_1 _2113_ (.B1(_1141_),
    .Y(_1142_),
    .A1(_1089_),
    .A2(_1101_));
 sg13g2_buf_8 _2114_ (.A(_1142_),
    .X(_1143_));
 sg13g2_buf_1 _2115_ (.A(_0163_),
    .X(_1144_));
 sg13g2_nor2_1 _2116_ (.A(_0196_),
    .B(net67),
    .Y(_1145_));
 sg13g2_xnor2_1 _2117_ (.Y(_1146_),
    .A(net102),
    .B(_1145_));
 sg13g2_buf_2 _2118_ (.A(_1146_),
    .X(_1147_));
 sg13g2_and4_1 _2119_ (.A(_0141_),
    .B(_0284_),
    .C(net29),
    .D(_1147_),
    .X(_1148_));
 sg13g2_nand2_1 _2120_ (.Y(_1149_),
    .A(_1067_),
    .B(_1147_));
 sg13g2_a21oi_1 _2121_ (.A1(_0141_),
    .A2(net29),
    .Y(_1150_),
    .B1(_1149_));
 sg13g2_nand2_1 _2122_ (.Y(_1151_),
    .A(net52),
    .B(_0273_));
 sg13g2_nor3_1 _2123_ (.A(_1113_),
    .B(_1140_),
    .C(_1151_),
    .Y(_1152_));
 sg13g2_and2_1 _2124_ (.A(_1089_),
    .B(_1152_),
    .X(_1153_));
 sg13g2_inv_1 _2125_ (.Y(_1154_),
    .A(net117));
 sg13g2_buf_1 _2126_ (.A(_1154_),
    .X(_1155_));
 sg13g2_xnor2_1 _2127_ (.Y(_1156_),
    .A(net89),
    .B(_0251_));
 sg13g2_nand3_1 _2128_ (.B(_1156_),
    .C(_1076_),
    .A(_0141_),
    .Y(_1157_));
 sg13g2_nor3_1 _2129_ (.A(_1089_),
    .B(_1101_),
    .C(_1157_),
    .Y(_1158_));
 sg13g2_a21o_1 _2130_ (.A2(_1100_),
    .A1(_1094_),
    .B1(_1140_),
    .X(_1159_));
 sg13g2_a21oi_1 _2131_ (.A1(_0141_),
    .A2(_1159_),
    .Y(_1160_),
    .B1(_1151_));
 sg13g2_buf_1 _2132_ (.A(net90),
    .X(_1161_));
 sg13g2_nand3_1 _2133_ (.B(net64),
    .C(_1156_),
    .A(net69),
    .Y(_1162_));
 sg13g2_o21ai_1 _2134_ (.B1(_1147_),
    .Y(_1163_),
    .A1(net111),
    .A2(_0728_));
 sg13g2_nor2_1 _2135_ (.A(net64),
    .B(net54),
    .Y(_1164_));
 sg13g2_a21oi_1 _2136_ (.A1(net66),
    .A2(_1163_),
    .Y(_1165_),
    .B1(_1164_));
 sg13g2_nand2_1 _2137_ (.Y(_1166_),
    .A(_1162_),
    .B(_1165_));
 sg13g2_o21ai_1 _2138_ (.B1(_1166_),
    .Y(_1167_),
    .A1(_1141_),
    .A2(_1157_));
 sg13g2_or4_1 _2139_ (.A(_1153_),
    .B(_1158_),
    .C(_1160_),
    .D(_1167_),
    .X(_1168_));
 sg13g2_nor3_1 _2140_ (.A(_1148_),
    .B(_1150_),
    .C(_1168_),
    .Y(_1169_));
 sg13g2_buf_1 _2141_ (.A(_1169_),
    .X(_1170_));
 sg13g2_xnor2_1 _2142_ (.Y(_1171_),
    .A(net68),
    .B(_0273_));
 sg13g2_nand2b_1 _2143_ (.Y(_1172_),
    .B(net66),
    .A_N(_1171_));
 sg13g2_xnor2_1 _2144_ (.Y(_1173_),
    .A(net111),
    .B(_1172_));
 sg13g2_nor2_1 _2145_ (.A(_1134_),
    .B(_1173_),
    .Y(_1174_));
 sg13g2_nor2_1 _2146_ (.A(net95),
    .B(_1034_),
    .Y(_1175_));
 sg13g2_nor4_1 _2147_ (.A(net95),
    .B(_1034_),
    .C(net46),
    .D(_1048_),
    .Y(_1176_));
 sg13g2_a221oi_1 _2148_ (.B2(_1175_),
    .C1(_1176_),
    .B1(_1097_),
    .A1(net66),
    .Y(_1177_),
    .A2(_1079_));
 sg13g2_buf_1 _2149_ (.A(_1177_),
    .X(_1178_));
 sg13g2_xnor2_1 _2150_ (.Y(_1179_),
    .A(net46),
    .B(_1178_));
 sg13g2_a21o_1 _2151_ (.A2(_1174_),
    .A1(_1142_),
    .B1(_1179_),
    .X(_1180_));
 sg13g2_buf_1 _2152_ (.A(_1180_),
    .X(_1181_));
 sg13g2_nand3_1 _2153_ (.B(_1174_),
    .C(_1179_),
    .A(net29),
    .Y(_1182_));
 sg13g2_buf_2 _2154_ (.A(_1182_),
    .X(_1183_));
 sg13g2_buf_1 _2155_ (.A(net116),
    .X(_1184_));
 sg13g2_buf_1 _2156_ (.A(net101),
    .X(_1185_));
 sg13g2_nor2_1 _2157_ (.A(net88),
    .B(_0728_),
    .Y(_1186_));
 sg13g2_a21oi_1 _2158_ (.A1(_1181_),
    .A2(_1183_),
    .Y(_1187_),
    .B1(_1186_));
 sg13g2_nand2_1 _2159_ (.Y(_1188_),
    .A(_0622_),
    .B(_1156_));
 sg13g2_nand2_1 _2160_ (.Y(_1189_),
    .A(net88),
    .B(_0728_));
 sg13g2_a21oi_1 _2161_ (.A1(net111),
    .A2(_1066_),
    .Y(_1190_),
    .B1(_1189_));
 sg13g2_a21oi_1 _2162_ (.A1(_1186_),
    .A2(_1188_),
    .Y(_1191_),
    .B1(_1190_));
 sg13g2_nor2_1 _2163_ (.A(_1050_),
    .B(_1191_),
    .Y(_1192_));
 sg13g2_nor3_1 _2164_ (.A(net46),
    .B(_1178_),
    .C(_1191_),
    .Y(_1193_));
 sg13g2_a21o_1 _2165_ (.A2(_1192_),
    .A1(_1178_),
    .B1(_1193_),
    .X(_1194_));
 sg13g2_nor2_1 _2166_ (.A(net64),
    .B(_0284_),
    .Y(_1195_));
 sg13g2_nand2_1 _2167_ (.Y(_1196_),
    .A(_1185_),
    .B(net54));
 sg13g2_nor2_1 _2168_ (.A(_1185_),
    .B(_1764_),
    .Y(_1197_));
 sg13g2_o21ai_1 _2169_ (.B1(_1197_),
    .Y(_1198_),
    .A1(_0372_),
    .A2(_1156_));
 sg13g2_o21ai_1 _2170_ (.B1(_1198_),
    .Y(_1199_),
    .A1(_1195_),
    .A2(_1196_));
 sg13g2_nand2_1 _2171_ (.Y(_1200_),
    .A(net46),
    .B(_1199_));
 sg13g2_nand2b_1 _2172_ (.Y(_1201_),
    .B(_1072_),
    .A_N(_1079_));
 sg13g2_nand3b_1 _2173_ (.B(_1199_),
    .C(_1050_),
    .Y(_1202_),
    .A_N(_1201_));
 sg13g2_o21ai_1 _2174_ (.B1(_1202_),
    .Y(_1203_),
    .A1(_1178_),
    .A2(_1200_));
 sg13g2_o21ai_1 _2175_ (.B1(net64),
    .Y(_1204_),
    .A1(net54),
    .A2(_1038_));
 sg13g2_a22oi_1 _2176_ (.Y(_1205_),
    .B1(_1171_),
    .B2(net111),
    .A2(_1204_),
    .A1(net95));
 sg13g2_nand2_1 _2177_ (.Y(_1206_),
    .A(net101),
    .B(net90));
 sg13g2_o21ai_1 _2178_ (.B1(_1172_),
    .Y(_1207_),
    .A1(_0948_),
    .A2(net46));
 sg13g2_nand2b_1 _2179_ (.Y(_1208_),
    .B(_1207_),
    .A_N(_1206_));
 sg13g2_o21ai_1 _2180_ (.B1(_1208_),
    .Y(_1209_),
    .A1(net88),
    .A2(_1205_));
 sg13g2_nor4_2 _2181_ (.A(_1134_),
    .B(_1194_),
    .C(_1203_),
    .Y(_1210_),
    .D(_1209_));
 sg13g2_and2_1 _2182_ (.A(_1210_),
    .B(net29),
    .X(_1211_));
 sg13g2_buf_8 _2183_ (.A(_1211_),
    .X(_1212_));
 sg13g2_and2_1 _2184_ (.A(net51),
    .B(_1065_),
    .X(_1213_));
 sg13g2_a221oi_1 _2185_ (.B2(net29),
    .C1(net47),
    .B1(_1210_),
    .A1(_1057_),
    .Y(_1214_),
    .A2(_1063_));
 sg13g2_a21oi_1 _2186_ (.A1(_1212_),
    .A2(_1213_),
    .Y(_1215_),
    .B1(_1214_));
 sg13g2_o21ai_1 _2187_ (.B1(_1215_),
    .Y(_1216_),
    .A1(net27),
    .A2(_1187_));
 sg13g2_buf_1 _2188_ (.A(_1216_),
    .X(_1217_));
 sg13g2_nand2_1 _2189_ (.Y(_1218_),
    .A(_1181_),
    .B(_1183_));
 sg13g2_buf_1 _2190_ (.A(_1218_),
    .X(_1219_));
 sg13g2_nand3_1 _2191_ (.B(_1181_),
    .C(_1183_),
    .A(_1186_),
    .Y(_1220_));
 sg13g2_a22oi_1 _2192_ (.Y(_1221_),
    .B1(_1220_),
    .B2(_1189_),
    .A2(net25),
    .A1(net27));
 sg13g2_buf_1 _2193_ (.A(_1221_),
    .X(_1222_));
 sg13g2_buf_1 _2194_ (.A(_1775_),
    .X(_1223_));
 sg13g2_a21o_1 _2195_ (.A2(_1094_),
    .A1(_1113_),
    .B1(_1140_),
    .X(_1224_));
 sg13g2_nand4_1 _2196_ (.B(_0141_),
    .C(_1224_),
    .A(net47),
    .Y(_1225_),
    .D(_1089_));
 sg13g2_xnor2_1 _2197_ (.Y(_1226_),
    .A(_1103_),
    .B(_1111_));
 sg13g2_nand2_1 _2198_ (.Y(_1227_),
    .A(_1226_),
    .B(_1105_));
 sg13g2_and2_1 _2199_ (.A(_0141_),
    .B(_1074_),
    .X(_1228_));
 sg13g2_buf_1 _2200_ (.A(_0989_),
    .X(_1229_));
 sg13g2_nor2_1 _2201_ (.A(net43),
    .B(_1134_),
    .Y(_1230_));
 sg13g2_and4_1 _2202_ (.A(_1078_),
    .B(_1074_),
    .C(_1085_),
    .D(_1230_),
    .X(_1231_));
 sg13g2_a221oi_1 _2203_ (.B2(_1065_),
    .C1(_1231_),
    .B1(_1230_),
    .A1(_1086_),
    .Y(_1232_),
    .A2(_1228_));
 sg13g2_nor4_1 _2204_ (.A(net47),
    .B(_0980_),
    .C(_1139_),
    .D(_1099_),
    .Y(_1233_));
 sg13g2_nor4_1 _2205_ (.A(net45),
    .B(_1709_),
    .C(_0980_),
    .D(_1099_),
    .Y(_1234_));
 sg13g2_nor3_1 _2206_ (.A(net45),
    .B(_1709_),
    .C(_1139_),
    .Y(_1235_));
 sg13g2_nor3_1 _2207_ (.A(_1233_),
    .B(_1234_),
    .C(_1235_),
    .Y(_1236_));
 sg13g2_or3_1 _2208_ (.A(_1227_),
    .B(_1232_),
    .C(_1236_),
    .X(_1237_));
 sg13g2_o21ai_1 _2209_ (.B1(_1227_),
    .Y(_1238_),
    .A1(_1232_),
    .A2(_1236_));
 sg13g2_nand3_1 _2210_ (.B(_1237_),
    .C(_1238_),
    .A(_1225_),
    .Y(_1239_));
 sg13g2_buf_1 _2211_ (.A(_1239_),
    .X(_1240_));
 sg13g2_a22oi_1 _2212_ (.Y(_1241_),
    .B1(_1240_),
    .B2(net45),
    .A2(_1139_),
    .A1(net38));
 sg13g2_nor2_1 _2213_ (.A(net47),
    .B(_1226_),
    .Y(_1242_));
 sg13g2_nand3_1 _2214_ (.B(_1226_),
    .C(_1105_),
    .A(net47),
    .Y(_1243_));
 sg13g2_o21ai_1 _2215_ (.B1(_1243_),
    .Y(_1244_),
    .A1(_1089_),
    .A2(_1242_));
 sg13g2_and3_1 _2216_ (.X(_1245_),
    .A(_1118_),
    .B(_1123_),
    .C(_1137_));
 sg13g2_nand2_1 _2217_ (.Y(_1246_),
    .A(_1126_),
    .B(_1245_));
 sg13g2_a21oi_2 _2218_ (.B1(_1246_),
    .Y(_1247_),
    .A2(_1244_),
    .A1(_1132_));
 sg13g2_nor2_2 _2219_ (.A(_1241_),
    .B(_1247_),
    .Y(_1248_));
 sg13g2_nor2_1 _2220_ (.A(net69),
    .B(_1134_),
    .Y(_1249_));
 sg13g2_a21oi_1 _2221_ (.A1(_1143_),
    .A2(_1249_),
    .Y(_1250_),
    .B1(_1156_));
 sg13g2_and3_1 _2222_ (.X(_1251_),
    .A(_1156_),
    .B(_1143_),
    .C(_1249_));
 sg13g2_xnor2_1 _2223_ (.Y(_1252_),
    .A(_1764_),
    .B(_1147_));
 sg13g2_nor2_1 _2224_ (.A(net69),
    .B(_1252_),
    .Y(_1253_));
 sg13g2_xnor2_1 _2225_ (.Y(_1254_),
    .A(net64),
    .B(_1253_));
 sg13g2_nor2_1 _2226_ (.A(_0130_),
    .B(_1254_),
    .Y(_1255_));
 sg13g2_o21ai_1 _2227_ (.B1(_1255_),
    .Y(_1256_),
    .A1(_1250_),
    .A2(_1251_));
 sg13g2_or4_1 _2228_ (.A(_1217_),
    .B(_1222_),
    .C(_1248_),
    .D(_1256_),
    .X(_1257_));
 sg13g2_nor2_1 _2229_ (.A(net45),
    .B(_1240_),
    .Y(_1258_));
 sg13g2_nand2_1 _2230_ (.Y(_1259_),
    .A(net47),
    .B(_1065_));
 sg13g2_a21o_1 _2231_ (.A2(net29),
    .A1(_1210_),
    .B1(_1259_),
    .X(_1260_));
 sg13g2_buf_1 _2232_ (.A(_1260_),
    .X(_1261_));
 sg13g2_nor2_1 _2233_ (.A(net51),
    .B(_1065_),
    .Y(_1262_));
 sg13g2_nand3_1 _2234_ (.B(net29),
    .C(_1262_),
    .A(_1210_),
    .Y(_1263_));
 sg13g2_buf_1 _2235_ (.A(_1263_),
    .X(_1264_));
 sg13g2_buf_1 _2236_ (.A(_0405_),
    .X(_1265_));
 sg13g2_buf_1 _2237_ (.A(net100),
    .X(_1266_));
 sg13g2_xnor2_1 _2238_ (.Y(_1267_),
    .A(net87),
    .B(net54));
 sg13g2_nor2_1 _2239_ (.A(_1267_),
    .B(_1134_),
    .Y(_1268_));
 sg13g2_nand2_1 _2240_ (.Y(_1269_),
    .A(_1100_),
    .B(_1268_));
 sg13g2_or2_1 _2241_ (.X(_1270_),
    .B(_1113_),
    .A(_0966_));
 sg13g2_mux2_1 _2242_ (.A0(_1269_),
    .A1(_1270_),
    .S(_1089_),
    .X(_1271_));
 sg13g2_a221oi_1 _2243_ (.B2(_1113_),
    .C1(_1139_),
    .B1(_1268_),
    .A1(_1135_),
    .Y(_1272_),
    .A2(_1242_));
 sg13g2_buf_1 _2244_ (.A(_1272_),
    .X(_1273_));
 sg13g2_nand3_1 _2245_ (.B(_1271_),
    .C(_1273_),
    .A(_1126_),
    .Y(_1274_));
 sg13g2_nand3_1 _2246_ (.B(_1264_),
    .C(_1274_),
    .A(_1261_),
    .Y(_1275_));
 sg13g2_or2_1 _2247_ (.X(_1276_),
    .B(_1251_),
    .A(_1250_));
 sg13g2_buf_1 _2248_ (.A(_1276_),
    .X(_1277_));
 sg13g2_nor3_1 _2249_ (.A(_1258_),
    .B(_1275_),
    .C(_1277_),
    .Y(_1278_));
 sg13g2_o21ai_1 _2250_ (.B1(_1278_),
    .Y(_1279_),
    .A1(_1217_),
    .A2(_1222_));
 sg13g2_nor2_1 _2251_ (.A(_1277_),
    .B(_1255_),
    .Y(_1280_));
 sg13g2_buf_1 _2252_ (.A(_1267_),
    .X(_1281_));
 sg13g2_and3_1 _2253_ (.X(_1282_),
    .A(_1225_),
    .B(_1237_),
    .C(_1238_));
 sg13g2_buf_1 _2254_ (.A(_1282_),
    .X(_1283_));
 sg13g2_nand2_1 _2255_ (.Y(_1284_),
    .A(net37),
    .B(_1283_));
 sg13g2_and3_1 _2256_ (.X(_1285_),
    .A(_1261_),
    .B(_1264_),
    .C(_1274_));
 sg13g2_nand2_1 _2257_ (.Y(_1286_),
    .A(net38),
    .B(_1139_));
 sg13g2_o21ai_1 _2258_ (.B1(_1286_),
    .Y(_1287_),
    .A1(_1267_),
    .A2(_1283_));
 sg13g2_inv_1 _2259_ (.Y(_1288_),
    .A(_1247_));
 sg13g2_a221oi_1 _2260_ (.B2(_1288_),
    .C1(_1256_),
    .B1(_1287_),
    .A1(_1284_),
    .Y(_1289_),
    .A2(_1285_));
 sg13g2_nor3_1 _2261_ (.A(_1241_),
    .B(_1247_),
    .C(_1277_),
    .Y(_1290_));
 sg13g2_nor3_1 _2262_ (.A(_1280_),
    .B(_1289_),
    .C(_1290_),
    .Y(_1291_));
 sg13g2_and3_1 _2263_ (.X(_1292_),
    .A(_1257_),
    .B(_1279_),
    .C(_1291_));
 sg13g2_buf_2 _2264_ (.A(_1292_),
    .X(_1293_));
 sg13g2_nand3_1 _2265_ (.B(_1279_),
    .C(_1291_),
    .A(_1257_),
    .Y(_1294_));
 sg13g2_buf_2 _2266_ (.A(_1294_),
    .X(_1295_));
 sg13g2_nor2_1 _2267_ (.A(_1258_),
    .B(_1275_),
    .Y(_1296_));
 sg13g2_o21ai_1 _2268_ (.B1(_1296_),
    .Y(_1297_),
    .A1(_1217_),
    .A2(_1222_));
 sg13g2_buf_1 _2269_ (.A(_1297_),
    .X(_1298_));
 sg13g2_buf_1 _2270_ (.A(_1102_),
    .X(_1299_));
 sg13g2_inv_1 _2271_ (.Y(_1300_),
    .A(_0185_));
 sg13g2_buf_1 _2272_ (.A(net118),
    .X(_1301_));
 sg13g2_nor2_1 _2273_ (.A(_0042_),
    .B(_0557_),
    .Y(_1302_));
 sg13g2_buf_2 _2274_ (.A(_1302_),
    .X(_1303_));
 sg13g2_nand2_1 _2275_ (.Y(_1304_),
    .A(net99),
    .B(_1303_));
 sg13g2_xnor2_1 _2276_ (.Y(_1305_),
    .A(_1300_),
    .B(_1304_));
 sg13g2_buf_1 _2277_ (.A(_1305_),
    .X(_1306_));
 sg13g2_xnor2_1 _2278_ (.Y(_1307_),
    .A(_0130_),
    .B(_1147_));
 sg13g2_nand3_1 _2279_ (.B(net36),
    .C(_1307_),
    .A(net49),
    .Y(_1308_));
 sg13g2_nor2_1 _2280_ (.A(_0130_),
    .B(_1147_),
    .Y(_1309_));
 sg13g2_o21ai_1 _2281_ (.B1(_1076_),
    .Y(_1310_),
    .A1(net36),
    .A2(_1309_));
 sg13g2_buf_1 _2282_ (.A(_0460_),
    .X(_1311_));
 sg13g2_inv_1 _2283_ (.Y(_1312_),
    .A(_1147_));
 sg13g2_o21ai_1 _2284_ (.B1(_0579_),
    .Y(_1313_),
    .A1(net86),
    .A2(_1312_));
 sg13g2_nor2_1 _2285_ (.A(net50),
    .B(_1312_),
    .Y(_1314_));
 sg13g2_a22oi_1 _2286_ (.Y(_1315_),
    .B1(_1314_),
    .B2(_0130_),
    .A2(_1313_),
    .A1(net69));
 sg13g2_nand3_1 _2287_ (.B(_1310_),
    .C(_1315_),
    .A(_1308_),
    .Y(_1316_));
 sg13g2_nor2_1 _2288_ (.A(_1248_),
    .B(_1316_),
    .Y(_1317_));
 sg13g2_nand2_1 _2289_ (.Y(_1318_),
    .A(net23),
    .B(_1317_));
 sg13g2_or2_1 _2290_ (.X(_1319_),
    .B(_1222_),
    .A(_1217_));
 sg13g2_nor2_1 _2291_ (.A(net49),
    .B(_1313_),
    .Y(_1320_));
 sg13g2_a21oi_1 _2292_ (.A1(net50),
    .A2(_1312_),
    .Y(_1321_),
    .B1(_1320_));
 sg13g2_o21ai_1 _2293_ (.B1(_1321_),
    .Y(_1322_),
    .A1(_1165_),
    .A2(net36));
 sg13g2_and2_1 _2294_ (.A(_1296_),
    .B(_1322_),
    .X(_1323_));
 sg13g2_and2_1 _2295_ (.A(_1248_),
    .B(_1322_),
    .X(_1324_));
 sg13g2_a21oi_1 _2296_ (.A1(_1319_),
    .A2(_1323_),
    .Y(_1325_),
    .B1(_1324_));
 sg13g2_nand2_1 _2297_ (.Y(_1326_),
    .A(_1318_),
    .B(_1325_));
 sg13g2_buf_1 _2298_ (.A(net53),
    .X(_1327_));
 sg13g2_xnor2_1 _2299_ (.Y(_1328_),
    .A(net42),
    .B(_1170_));
 sg13g2_nor4_2 _2300_ (.A(_0130_),
    .B(_1219_),
    .C(_1248_),
    .Y(_1329_),
    .D(_1328_));
 sg13g2_nor2b_1 _2301_ (.A(net116),
    .B_N(_1610_),
    .Y(_1330_));
 sg13g2_buf_2 _2302_ (.A(_1330_),
    .X(_1331_));
 sg13g2_nand3_1 _2303_ (.B(_1329_),
    .C(_1331_),
    .A(net23),
    .Y(_1332_));
 sg13g2_buf_1 _2304_ (.A(_0987_),
    .X(_1333_));
 sg13g2_nor2_2 _2305_ (.A(net94),
    .B(net85),
    .Y(_1334_));
 sg13g2_nand3_1 _2306_ (.B(_1329_),
    .C(_1334_),
    .A(net23),
    .Y(_1335_));
 sg13g2_nor2_1 _2307_ (.A(_1134_),
    .B(_1139_),
    .Y(_1336_));
 sg13g2_xnor2_1 _2308_ (.Y(_1337_),
    .A(_1267_),
    .B(_1244_));
 sg13g2_nand3_1 _2309_ (.B(_1336_),
    .C(_1337_),
    .A(net42),
    .Y(_1338_));
 sg13g2_nand3_1 _2310_ (.B(_1336_),
    .C(_1337_),
    .A(net43),
    .Y(_1339_));
 sg13g2_mux2_1 _2311_ (.A0(_1338_),
    .A1(_1339_),
    .S(net27),
    .X(_1340_));
 sg13g2_nand3_1 _2312_ (.B(_1340_),
    .C(_1331_),
    .A(net25),
    .Y(_1341_));
 sg13g2_nand3_1 _2313_ (.B(_1340_),
    .C(_1334_),
    .A(net25),
    .Y(_1342_));
 sg13g2_xor2_1 _2314_ (.B(_1212_),
    .A(_1065_),
    .X(_1343_));
 sg13g2_a221oi_1 _2315_ (.B2(net42),
    .C1(_1258_),
    .B1(net25),
    .A1(net39),
    .Y(_1344_),
    .A2(_1343_));
 sg13g2_o21ai_1 _2316_ (.B1(net27),
    .Y(_1345_),
    .A1(net42),
    .A2(net25));
 sg13g2_nand2_1 _2317_ (.Y(_1346_),
    .A(_1215_),
    .B(_1283_));
 sg13g2_o21ai_1 _2318_ (.B1(net37),
    .Y(_1347_),
    .A1(_1215_),
    .A2(_1283_));
 sg13g2_a21oi_1 _2319_ (.A1(net38),
    .A2(_1139_),
    .Y(_1348_),
    .B1(_0130_));
 sg13g2_nand2_1 _2320_ (.Y(_1349_),
    .A(net42),
    .B(_1348_));
 sg13g2_nand2_1 _2321_ (.Y(_1350_),
    .A(net43),
    .B(_1348_));
 sg13g2_mux2_1 _2322_ (.A0(_1349_),
    .A1(_1350_),
    .S(net27),
    .X(_1351_));
 sg13g2_a221oi_1 _2323_ (.B2(_1347_),
    .C1(_1351_),
    .B1(_1346_),
    .A1(_1344_),
    .Y(_1352_),
    .A2(_1345_));
 sg13g2_a21o_1 _2324_ (.A2(_1342_),
    .A1(_1341_),
    .B1(_1352_),
    .X(_1353_));
 sg13g2_buf_1 _2325_ (.A(net94),
    .X(_1354_));
 sg13g2_buf_1 _2326_ (.A(net88),
    .X(_1355_));
 sg13g2_nor3_1 _2327_ (.A(_1354_),
    .B(net62),
    .C(net54),
    .Y(_1356_));
 sg13g2_nand3_1 _2328_ (.B(net62),
    .C(net54),
    .A(_1354_),
    .Y(_1357_));
 sg13g2_nor2b_1 _2329_ (.A(_1356_),
    .B_N(_1357_),
    .Y(_1358_));
 sg13g2_nand4_1 _2330_ (.B(_1335_),
    .C(_1353_),
    .A(_1332_),
    .Y(_1359_),
    .D(_1358_));
 sg13g2_a21o_1 _2331_ (.A2(_1326_),
    .A1(_1295_),
    .B1(_1359_),
    .X(_1360_));
 sg13g2_nand2_1 _2332_ (.Y(_1361_),
    .A(net23),
    .B(_1329_));
 sg13g2_nand3b_1 _2333_ (.B(_1340_),
    .C(net25),
    .Y(_1362_),
    .A_N(_1352_));
 sg13g2_buf_1 _2334_ (.A(_1362_),
    .X(_1363_));
 sg13g2_a221oi_1 _2335_ (.B2(_1319_),
    .C1(_1324_),
    .B1(_1323_),
    .A1(_1298_),
    .Y(_1364_),
    .A2(_1317_));
 sg13g2_buf_1 _2336_ (.A(_1364_),
    .X(_1365_));
 sg13g2_nand4_1 _2337_ (.B(_1363_),
    .C(_1293_),
    .A(_1361_),
    .Y(_1366_),
    .D(_1365_));
 sg13g2_buf_1 _2338_ (.A(net51),
    .X(_1367_));
 sg13g2_nand3_1 _2339_ (.B(_1293_),
    .C(_1365_),
    .A(net41),
    .Y(_1368_));
 sg13g2_nand3_1 _2340_ (.B(_1361_),
    .C(_1363_),
    .A(net41),
    .Y(_1369_));
 sg13g2_or2_1 _2341_ (.X(_1370_),
    .B(_1343_),
    .A(net37));
 sg13g2_buf_1 _2342_ (.A(net45),
    .X(_1371_));
 sg13g2_nand2_1 _2343_ (.Y(_1372_),
    .A(net35),
    .B(_1343_));
 sg13g2_nor2_1 _2344_ (.A(_0130_),
    .B(_1248_),
    .Y(_1373_));
 sg13g2_nand2_1 _2345_ (.Y(_1374_),
    .A(net27),
    .B(net25));
 sg13g2_o21ai_1 _2346_ (.B1(net42),
    .Y(_1375_),
    .A1(net27),
    .A2(net25));
 sg13g2_a21o_1 _2347_ (.A2(_1375_),
    .A1(_1374_),
    .B1(net41),
    .X(_1376_));
 sg13g2_nand3_1 _2348_ (.B(_1374_),
    .C(_1375_),
    .A(net41),
    .Y(_1377_));
 sg13g2_and4_1 _2349_ (.A(net23),
    .B(_1373_),
    .C(_1376_),
    .D(_1377_),
    .X(_1378_));
 sg13g2_buf_2 _2350_ (.A(_1378_),
    .X(_1379_));
 sg13g2_mux2_1 _2351_ (.A0(_1370_),
    .A1(_1372_),
    .S(_1379_),
    .X(_1380_));
 sg13g2_and4_1 _2352_ (.A(_1366_),
    .B(_1368_),
    .C(_1369_),
    .D(_1380_),
    .X(_1381_));
 sg13g2_xnor2_1 _2353_ (.Y(_1382_),
    .A(_1343_),
    .B(_1379_));
 sg13g2_nor2_1 _2354_ (.A(net35),
    .B(_1382_),
    .Y(_1383_));
 sg13g2_a21oi_1 _2355_ (.A1(_1360_),
    .A2(_1381_),
    .Y(_1384_),
    .B1(_1383_));
 sg13g2_buf_8 _2356_ (.A(_1384_),
    .X(_1385_));
 sg13g2_nand4_1 _2357_ (.B(_1183_),
    .C(_1261_),
    .A(_1181_),
    .Y(_1386_),
    .D(_1264_));
 sg13g2_nand3_1 _2358_ (.B(_1261_),
    .C(_1264_),
    .A(net43),
    .Y(_1387_));
 sg13g2_a21o_1 _2359_ (.A2(_1387_),
    .A1(_1386_),
    .B1(net27),
    .X(_1388_));
 sg13g2_buf_1 _2360_ (.A(_1388_),
    .X(_1389_));
 sg13g2_and4_1 _2361_ (.A(_1181_),
    .B(_1183_),
    .C(_1261_),
    .D(_1264_),
    .X(_1390_));
 sg13g2_a221oi_1 _2362_ (.B2(net43),
    .C1(_1214_),
    .B1(_1390_),
    .A1(_1212_),
    .Y(_1391_),
    .A2(_1213_));
 sg13g2_buf_1 _2363_ (.A(_1391_),
    .X(_1392_));
 sg13g2_o21ai_1 _2364_ (.B1(_1092_),
    .Y(_1393_),
    .A1(_1246_),
    .A2(_1244_));
 sg13g2_nand3_1 _2365_ (.B(_1240_),
    .C(_1393_),
    .A(_1348_),
    .Y(_1394_));
 sg13g2_nand2_1 _2366_ (.Y(_1395_),
    .A(_1132_),
    .B(_1286_));
 sg13g2_a21oi_1 _2367_ (.A1(_1395_),
    .A2(_1283_),
    .Y(_1396_),
    .B1(_1092_));
 sg13g2_o21ai_1 _2368_ (.B1(_1396_),
    .Y(_1397_),
    .A1(_1285_),
    .A2(_1394_));
 sg13g2_a21oi_1 _2369_ (.A1(_1389_),
    .A2(_1392_),
    .Y(_1398_),
    .B1(_1397_));
 sg13g2_a21oi_1 _2370_ (.A1(_1395_),
    .A2(_1283_),
    .Y(_1399_),
    .B1(net37));
 sg13g2_and4_1 _2371_ (.A(_1389_),
    .B(_1392_),
    .C(_1394_),
    .D(_1399_),
    .X(_1400_));
 sg13g2_nand2_1 _2372_ (.Y(_1401_),
    .A(net35),
    .B(_1240_));
 sg13g2_a21oi_1 _2373_ (.A1(_1389_),
    .A2(_1392_),
    .Y(_1402_),
    .B1(_1401_));
 sg13g2_and4_1 _2374_ (.A(net37),
    .B(_1240_),
    .C(_1389_),
    .D(_1392_),
    .X(_1403_));
 sg13g2_nor4_2 _2375_ (.A(_1398_),
    .B(_1400_),
    .C(_1402_),
    .Y(_1404_),
    .D(_1403_));
 sg13g2_buf_1 _2376_ (.A(_1404_),
    .X(_1405_));
 sg13g2_and2_1 _2377_ (.A(net23),
    .B(_1373_),
    .X(_1406_));
 sg13g2_buf_2 _2378_ (.A(_1406_),
    .X(_1407_));
 sg13g2_a22oi_1 _2379_ (.Y(_1408_),
    .B1(_1346_),
    .B2(_1347_),
    .A2(_1345_),
    .A1(_1344_));
 sg13g2_xnor2_1 _2380_ (.Y(_1409_),
    .A(net38),
    .B(_1408_));
 sg13g2_nand2_2 _2381_ (.Y(_1410_),
    .A(_1271_),
    .B(_1273_));
 sg13g2_a21oi_2 _2382_ (.B1(_1410_),
    .Y(_1411_),
    .A2(_1409_),
    .A1(_1407_));
 sg13g2_a22oi_1 _2383_ (.Y(_1412_),
    .B1(_1411_),
    .B2(_0108_),
    .A2(net22),
    .A1(_1126_));
 sg13g2_buf_1 _2384_ (.A(_1412_),
    .X(_1413_));
 sg13g2_nand2_1 _2385_ (.Y(_1414_),
    .A(net42),
    .B(_1365_));
 sg13g2_nand2_1 _2386_ (.Y(_1415_),
    .A(net43),
    .B(_1326_));
 sg13g2_nor2_1 _2387_ (.A(_0108_),
    .B(_1245_),
    .Y(_1416_));
 sg13g2_nor2_1 _2388_ (.A(net65),
    .B(_1416_),
    .Y(_1417_));
 sg13g2_nor3_1 _2389_ (.A(net65),
    .B(net44),
    .C(_1410_),
    .Y(_1418_));
 sg13g2_nand3_1 _2390_ (.B(_1373_),
    .C(_1408_),
    .A(net23),
    .Y(_1419_));
 sg13g2_nor2_1 _2391_ (.A(_1223_),
    .B(net65),
    .Y(_1420_));
 sg13g2_nor2b_1 _2392_ (.A(_1416_),
    .B_N(_1420_),
    .Y(_1421_));
 sg13g2_a221oi_1 _2393_ (.B2(_1419_),
    .C1(_1421_),
    .B1(_1418_),
    .A1(_1404_),
    .Y(_1422_),
    .A2(_1417_));
 sg13g2_buf_1 _2394_ (.A(_1422_),
    .X(_1423_));
 sg13g2_a221oi_1 _2395_ (.B2(_1415_),
    .C1(_1423_),
    .B1(_1414_),
    .A1(_1385_),
    .Y(_1424_),
    .A2(_1413_));
 sg13g2_buf_2 _2396_ (.A(_1424_),
    .X(_1425_));
 sg13g2_xnor2_1 _2397_ (.Y(_1426_),
    .A(_1293_),
    .B(_1425_));
 sg13g2_nand2b_1 _2398_ (.Y(_1427_),
    .B(net38),
    .A_N(_1404_));
 sg13g2_inv_1 _2399_ (.Y(_1428_),
    .A(_1416_));
 sg13g2_nor2_1 _2400_ (.A(net44),
    .B(_1410_),
    .Y(_1429_));
 sg13g2_a22oi_1 _2401_ (.Y(_1430_),
    .B1(_1429_),
    .B2(_1419_),
    .A2(_1428_),
    .A1(_1427_));
 sg13g2_buf_1 _2402_ (.A(net114),
    .X(_1431_));
 sg13g2_a221oi_1 _2403_ (.B2(net96),
    .C1(net69),
    .B1(net52),
    .A1(net120),
    .Y(_1432_),
    .A2(net84));
 sg13g2_buf_1 _2404_ (.A(_0185_),
    .X(_1433_));
 sg13g2_buf_1 _2405_ (.A(net98),
    .X(_1434_));
 sg13g2_nor2_1 _2406_ (.A(net108),
    .B(net64),
    .Y(_1435_));
 sg13g2_buf_1 _2407_ (.A(_1301_),
    .X(_1436_));
 sg13g2_a22oi_1 _2408_ (.Y(_1437_),
    .B1(_1006_),
    .B2(net82),
    .A2(_1435_),
    .A1(_1434_));
 sg13g2_buf_1 _2409_ (.A(net129),
    .X(_1438_));
 sg13g2_a21oi_1 _2410_ (.A1(net49),
    .A2(net122),
    .Y(_1439_),
    .B1(net86));
 sg13g2_a221oi_1 _2411_ (.B2(net36),
    .C1(_0739_),
    .B1(_1439_),
    .A1(net49),
    .Y(_1440_),
    .A2(_1437_));
 sg13g2_a21oi_1 _2412_ (.A1(net36),
    .A2(_1432_),
    .Y(_1441_),
    .B1(_1440_));
 sg13g2_nand2b_1 _2413_ (.Y(_1442_),
    .B(_1441_),
    .A_N(_1430_));
 sg13g2_nand2_1 _2414_ (.Y(_1443_),
    .A(net96),
    .B(_1299_));
 sg13g2_a21oi_1 _2415_ (.A1(_1443_),
    .A2(_0948_),
    .Y(_1444_),
    .B1(_1014_));
 sg13g2_nor2_1 _2416_ (.A(net36),
    .B(_1444_),
    .Y(_1445_));
 sg13g2_nor2_1 _2417_ (.A(_1440_),
    .B(_1445_),
    .Y(_1446_));
 sg13g2_nand2_1 _2418_ (.Y(_1447_),
    .A(_1413_),
    .B(_1446_));
 sg13g2_mux2_1 _2419_ (.A0(_1442_),
    .A1(_1447_),
    .S(_1385_),
    .X(_1448_));
 sg13g2_buf_2 _2420_ (.A(_1448_),
    .X(_1449_));
 sg13g2_a21o_1 _2421_ (.A2(_1409_),
    .A1(_1407_),
    .B1(_1410_),
    .X(_1450_));
 sg13g2_buf_2 _2422_ (.A(_1450_),
    .X(_1451_));
 sg13g2_nand2_1 _2423_ (.Y(_1452_),
    .A(_1126_),
    .B(net22));
 sg13g2_o21ai_1 _2424_ (.B1(_1452_),
    .Y(_1453_),
    .A1(net44),
    .A2(_1451_));
 sg13g2_nand3b_1 _2425_ (.B(_1441_),
    .C(_1453_),
    .Y(_1454_),
    .A_N(_1430_));
 sg13g2_nand2_1 _2426_ (.Y(_1455_),
    .A(_1430_),
    .B(_1446_));
 sg13g2_and2_1 _2427_ (.A(_1454_),
    .B(_1455_),
    .X(_1456_));
 sg13g2_buf_1 _2428_ (.A(_1456_),
    .X(_1457_));
 sg13g2_nand2_2 _2429_ (.Y(_1458_),
    .A(_1449_),
    .B(_1457_));
 sg13g2_a21o_1 _2430_ (.A2(_1381_),
    .A1(_1360_),
    .B1(_1383_),
    .X(_1459_));
 sg13g2_buf_2 _2431_ (.A(_1459_),
    .X(_1460_));
 sg13g2_buf_1 _2432_ (.A(net64),
    .X(_1461_));
 sg13g2_xnor2_1 _2433_ (.Y(_1462_),
    .A(net54),
    .B(net36));
 sg13g2_nor2_1 _2434_ (.A(net55),
    .B(_1462_),
    .Y(_1463_));
 sg13g2_xnor2_1 _2435_ (.Y(_1464_),
    .A(net48),
    .B(_1463_));
 sg13g2_nor2_1 _2436_ (.A(_1423_),
    .B(_1464_),
    .Y(_1465_));
 sg13g2_o21ai_1 _2437_ (.B1(_1465_),
    .Y(_1466_),
    .A1(_1460_),
    .A2(_1453_));
 sg13g2_nand2_1 _2438_ (.Y(_1467_),
    .A(net23),
    .B(_1373_));
 sg13g2_nor2_1 _2439_ (.A(net55),
    .B(_1467_),
    .Y(_1468_));
 sg13g2_xnor2_1 _2440_ (.Y(_1469_),
    .A(_1147_),
    .B(_1468_));
 sg13g2_xor2_1 _2441_ (.B(_1469_),
    .A(_1466_),
    .X(_1470_));
 sg13g2_buf_8 _2442_ (.A(_1470_),
    .X(_1471_));
 sg13g2_nand2_1 _2443_ (.Y(_1472_),
    .A(_1458_),
    .B(_1471_));
 sg13g2_o21ai_1 _2444_ (.B1(net43),
    .Y(_1473_),
    .A1(_1458_),
    .A2(_1471_));
 sg13g2_buf_1 _2445_ (.A(_1473_),
    .X(_1474_));
 sg13g2_nand2_2 _2446_ (.Y(_1475_),
    .A(_1361_),
    .B(_1363_));
 sg13g2_nand2_1 _2447_ (.Y(_1476_),
    .A(_1293_),
    .B(_1365_));
 sg13g2_nor2_1 _2448_ (.A(_1293_),
    .B(_1365_),
    .Y(_1477_));
 sg13g2_a21oi_1 _2449_ (.A1(net42),
    .A2(_1476_),
    .Y(_1478_),
    .B1(_1477_));
 sg13g2_or2_1 _2450_ (.X(_1479_),
    .B(_1478_),
    .A(net39));
 sg13g2_nand2_1 _2451_ (.Y(_1480_),
    .A(net39),
    .B(_1478_));
 sg13g2_a221oi_1 _2452_ (.B2(_1480_),
    .C1(_1423_),
    .B1(_1479_),
    .A1(_1385_),
    .Y(_1481_),
    .A2(_1413_));
 sg13g2_xor2_1 _2453_ (.B(_1481_),
    .A(_1475_),
    .X(_1482_));
 sg13g2_and2_1 _2454_ (.A(net37),
    .B(_1482_),
    .X(_1483_));
 sg13g2_a221oi_1 _2455_ (.B2(_1474_),
    .C1(_1483_),
    .B1(_1472_),
    .A1(net39),
    .Y(_1484_),
    .A2(_1426_));
 sg13g2_buf_2 _2456_ (.A(_1484_),
    .X(_1485_));
 sg13g2_xnor2_1 _2457_ (.Y(_1486_),
    .A(_1295_),
    .B(_1425_));
 sg13g2_buf_1 _2458_ (.A(_1486_),
    .X(_1487_));
 sg13g2_nand2_1 _2459_ (.Y(_1488_),
    .A(net41),
    .B(_1487_));
 sg13g2_or2_1 _2460_ (.X(_1489_),
    .B(_1482_),
    .A(net37));
 sg13g2_o21ai_1 _2461_ (.B1(_1489_),
    .Y(_1490_),
    .A1(_1488_),
    .A2(_1483_));
 sg13g2_buf_2 _2462_ (.A(_1490_),
    .X(_1491_));
 sg13g2_o21ai_1 _2463_ (.B1(_1359_),
    .Y(_1492_),
    .A1(_1475_),
    .A2(_1295_));
 sg13g2_o21ai_1 _2464_ (.B1(_1326_),
    .Y(_1493_),
    .A1(_1295_),
    .A2(_1359_));
 sg13g2_nor2_1 _2465_ (.A(net35),
    .B(_1423_),
    .Y(_1494_));
 sg13g2_and3_1 _2466_ (.X(_1495_),
    .A(_1492_),
    .B(_1493_),
    .C(_1494_));
 sg13g2_a21oi_2 _2467_ (.B1(net39),
    .Y(_1496_),
    .A2(_1476_),
    .A1(_1475_));
 sg13g2_nand2b_1 _2468_ (.Y(_1497_),
    .B(net35),
    .A_N(_1423_));
 sg13g2_nor3_1 _2469_ (.A(_1496_),
    .B(_1492_),
    .C(_1497_),
    .Y(_1498_));
 sg13g2_nor2_1 _2470_ (.A(_1495_),
    .B(_1498_),
    .Y(_1499_));
 sg13g2_nor3_1 _2471_ (.A(_1496_),
    .B(_1493_),
    .C(_1497_),
    .Y(_1500_));
 sg13g2_a21o_1 _2472_ (.A2(_1494_),
    .A1(_1496_),
    .B1(_1382_),
    .X(_1502_));
 sg13g2_nor2_1 _2473_ (.A(_1500_),
    .B(_1502_),
    .Y(_1503_));
 sg13g2_xor2_1 _2474_ (.B(_1379_),
    .A(_1343_),
    .X(_1504_));
 sg13g2_nor3_1 _2475_ (.A(_1504_),
    .B(_1413_),
    .C(_1423_),
    .Y(_1505_));
 sg13g2_a21oi_1 _2476_ (.A1(_1492_),
    .A2(_1493_),
    .Y(_1506_),
    .B1(_1496_));
 sg13g2_xnor2_1 _2477_ (.Y(_1507_),
    .A(net35),
    .B(_1506_));
 sg13g2_buf_1 _2478_ (.A(_1126_),
    .X(_1508_));
 sg13g2_a221oi_1 _2479_ (.B2(_1507_),
    .C1(net34),
    .B1(_1505_),
    .A1(_1499_),
    .Y(_1509_),
    .A2(_1503_));
 sg13g2_inv_1 _2480_ (.Y(_1510_),
    .A(_1452_));
 sg13g2_o21ai_1 _2481_ (.B1(_1427_),
    .Y(_1511_),
    .A1(_1460_),
    .A2(_1510_));
 sg13g2_nand3_1 _2482_ (.B(_1411_),
    .C(_1511_),
    .A(net44),
    .Y(_1513_));
 sg13g2_a21o_1 _2483_ (.A2(_1413_),
    .A1(_1385_),
    .B1(_1423_),
    .X(_1514_));
 sg13g2_buf_2 _2484_ (.A(_1514_),
    .X(_1515_));
 sg13g2_xnor2_1 _2485_ (.Y(_1516_),
    .A(net38),
    .B(_1385_));
 sg13g2_and2_1 _2486_ (.A(_0108_),
    .B(net22),
    .X(_1517_));
 sg13g2_o21ai_1 _2487_ (.B1(_1517_),
    .Y(_1518_),
    .A1(_1515_),
    .A2(_1516_));
 sg13g2_nand2_1 _2488_ (.Y(_1519_),
    .A(net38),
    .B(net65));
 sg13g2_a21oi_1 _2489_ (.A1(_1460_),
    .A2(_1519_),
    .Y(_1520_),
    .B1(_1420_));
 sg13g2_nand3b_1 _2490_ (.B(_1411_),
    .C(_0108_),
    .Y(_1521_),
    .A_N(_1520_));
 sg13g2_nand4_1 _2491_ (.B(_1513_),
    .C(_1518_),
    .A(_1509_),
    .Y(_1522_),
    .D(_1521_));
 sg13g2_nand2_1 _2492_ (.Y(_1524_),
    .A(net22),
    .B(_1411_));
 sg13g2_mux2_1 _2493_ (.A0(net22),
    .A1(_1524_),
    .S(_1385_),
    .X(_1525_));
 sg13g2_nor2_1 _2494_ (.A(net34),
    .B(_1524_),
    .Y(_1526_));
 sg13g2_nor2_1 _2495_ (.A(net22),
    .B(_1411_),
    .Y(_1527_));
 sg13g2_a21oi_1 _2496_ (.A1(_1460_),
    .A2(_1526_),
    .Y(_1528_),
    .B1(_1527_));
 sg13g2_o21ai_1 _2497_ (.B1(_1528_),
    .Y(_1529_),
    .A1(_1223_),
    .A2(_1525_));
 sg13g2_a21oi_1 _2498_ (.A1(_1131_),
    .A2(_1529_),
    .Y(_1530_),
    .B1(net65));
 sg13g2_or4_1 _2499_ (.A(net44),
    .B(_1405_),
    .C(_1515_),
    .D(_1516_),
    .X(_1531_));
 sg13g2_nand2_1 _2500_ (.Y(_1532_),
    .A(_1518_),
    .B(_1531_));
 sg13g2_and2_1 _2501_ (.A(_1271_),
    .B(_1273_),
    .X(_1533_));
 sg13g2_nor2_1 _2502_ (.A(net38),
    .B(_1385_),
    .Y(_1535_));
 sg13g2_nor3_1 _2503_ (.A(net65),
    .B(_0108_),
    .C(_1451_),
    .Y(_1536_));
 sg13g2_o21ai_1 _2504_ (.B1(_1536_),
    .Y(_1537_),
    .A1(net34),
    .A2(_1460_));
 sg13g2_nand2b_1 _2505_ (.Y(_1538_),
    .B(_1131_),
    .A_N(net22));
 sg13g2_o21ai_1 _2506_ (.B1(_1538_),
    .Y(_1539_),
    .A1(_1535_),
    .A2(_1537_));
 sg13g2_nor3_1 _2507_ (.A(_1410_),
    .B(_1509_),
    .C(_1539_),
    .Y(_1540_));
 sg13g2_a221oi_1 _2508_ (.B2(_1533_),
    .C1(_1540_),
    .B1(_1532_),
    .A1(_1522_),
    .Y(_1541_),
    .A2(_1530_));
 sg13g2_or3_1 _2509_ (.A(_1485_),
    .B(_1491_),
    .C(_1541_),
    .X(_1542_));
 sg13g2_buf_8 _2510_ (.A(_1542_),
    .X(_1543_));
 sg13g2_nand2_1 _2511_ (.Y(_1544_),
    .A(_1522_),
    .B(_1530_));
 sg13g2_and2_1 _2512_ (.A(_1518_),
    .B(_1531_),
    .X(_1546_));
 sg13g2_nor4_1 _2513_ (.A(_1495_),
    .B(_1498_),
    .C(_1500_),
    .D(_1502_),
    .Y(_1547_));
 sg13g2_a21o_1 _2514_ (.A2(_1505_),
    .A1(_1507_),
    .B1(_1547_),
    .X(_1548_));
 sg13g2_buf_2 _2515_ (.A(_1548_),
    .X(_1549_));
 sg13g2_nand3b_1 _2516_ (.B(_1549_),
    .C(net34),
    .Y(_1550_),
    .A_N(_1539_));
 sg13g2_a21o_1 _2517_ (.A2(_1550_),
    .A1(_1546_),
    .B1(_1410_),
    .X(_1551_));
 sg13g2_o21ai_1 _2518_ (.B1(net22),
    .Y(_1552_),
    .A1(_1128_),
    .A2(_1516_));
 sg13g2_o21ai_1 _2519_ (.B1(_1552_),
    .Y(_1553_),
    .A1(_1451_),
    .A2(_1520_));
 sg13g2_and3_1 _2520_ (.X(_1554_),
    .A(net44),
    .B(_1411_),
    .C(_1511_));
 sg13g2_a221oi_1 _2521_ (.B2(_0108_),
    .C1(_1554_),
    .B1(_1553_),
    .A1(net34),
    .Y(_1555_),
    .A2(_1549_));
 sg13g2_a21o_1 _2522_ (.A2(_1551_),
    .A1(_1544_),
    .B1(_1555_),
    .X(_1557_));
 sg13g2_buf_1 _2523_ (.A(_1557_),
    .X(_1558_));
 sg13g2_nand2_1 _2524_ (.Y(_1559_),
    .A(net19),
    .B(net20));
 sg13g2_nand2_1 _2525_ (.Y(_1560_),
    .A(_1599_),
    .B(_1559_));
 sg13g2_buf_1 _2526_ (.A(_1599_),
    .X(_1561_));
 sg13g2_nor3_2 _2527_ (.A(_1485_),
    .B(_1491_),
    .C(_1541_),
    .Y(_1562_));
 sg13g2_a21oi_2 _2528_ (.B1(_1555_),
    .Y(_1563_),
    .A2(_1551_),
    .A1(_1544_));
 sg13g2_nor2_1 _2529_ (.A(_1562_),
    .B(_1563_),
    .Y(_1564_));
 sg13g2_buf_2 _2530_ (.A(_1564_),
    .X(_1565_));
 sg13g2_nand2_1 _2531_ (.Y(_1566_),
    .A(net82),
    .B(net55));
 sg13g2_o21ai_1 _2532_ (.B1(_1566_),
    .Y(_1568_),
    .A1(_1443_),
    .A2(_1565_));
 sg13g2_and2_1 _2533_ (.A(net128),
    .B(_1568_),
    .X(_1569_));
 sg13g2_a21o_1 _2534_ (.A2(_1560_),
    .A1(_1588_),
    .B1(_1569_),
    .X(_1570_));
 sg13g2_buf_1 _2535_ (.A(uio_in[0]),
    .X(_1571_));
 sg13g2_buf_1 _2536_ (.A(net131),
    .X(_1572_));
 sg13g2_mux2_1 _2537_ (.A0(\muldiv.regR[0] ),
    .A1(_1570_),
    .S(net127),
    .X(_0004_));
 sg13g2_inv_2 _2538_ (.Y(_1573_),
    .A(_1599_));
 sg13g2_buf_1 _2539_ (.A(_1573_),
    .X(_1574_));
 sg13g2_buf_1 _2540_ (.A(net122),
    .X(_1575_));
 sg13g2_buf_1 _2541_ (.A(net109),
    .X(_1576_));
 sg13g2_buf_1 _2542_ (.A(net84),
    .X(_1578_));
 sg13g2_xor2_1 _2543_ (.B(net61),
    .A(net81),
    .X(_1579_));
 sg13g2_nand2_1 _2544_ (.Y(_1580_),
    .A(net119),
    .B(_1579_));
 sg13g2_buf_1 _2545_ (.A(_1580_),
    .X(_1581_));
 sg13g2_and3_1 _2546_ (.X(_1582_),
    .A(_1515_),
    .B(net19),
    .C(net20));
 sg13g2_buf_1 _2547_ (.A(_1582_),
    .X(_1583_));
 sg13g2_nor2_1 _2548_ (.A(_1581_),
    .B(_1583_),
    .Y(_1584_));
 sg13g2_xnor2_1 _2549_ (.Y(_1585_),
    .A(_1407_),
    .B(_1584_));
 sg13g2_buf_1 _2550_ (.A(net49),
    .X(_1586_));
 sg13g2_a21o_1 _2551_ (.A2(net112),
    .A1(net107),
    .B1(net116),
    .X(_1587_));
 sg13g2_buf_2 _2552_ (.A(_1587_),
    .X(_1589_));
 sg13g2_nand3_1 _2553_ (.B(net116),
    .C(net112),
    .A(net118),
    .Y(_1590_));
 sg13g2_mux2_1 _2554_ (.A0(_1589_),
    .A1(_1590_),
    .S(_0394_),
    .X(_1591_));
 sg13g2_nand2_1 _2555_ (.Y(_1592_),
    .A(_1512_),
    .B(net115));
 sg13g2_o21ai_1 _2556_ (.B1(_1592_),
    .Y(_1593_),
    .A1(net100),
    .A2(_1591_));
 sg13g2_nand2_1 _2557_ (.Y(_1594_),
    .A(net115),
    .B(_1589_));
 sg13g2_a21oi_2 _2558_ (.B1(_1610_),
    .Y(_1595_),
    .A2(net112),
    .A1(_0986_));
 sg13g2_nor2_1 _2559_ (.A(_1300_),
    .B(_1595_),
    .Y(_1596_));
 sg13g2_nand2_1 _2560_ (.Y(_1597_),
    .A(net118),
    .B(net100));
 sg13g2_a21oi_1 _2561_ (.A1(_1594_),
    .A2(_1596_),
    .Y(_1598_),
    .B1(_1597_));
 sg13g2_a21oi_1 _2562_ (.A1(net98),
    .A2(_1593_),
    .Y(_1600_),
    .B1(_1598_));
 sg13g2_and2_1 _2563_ (.A(net107),
    .B(_0185_),
    .X(_1601_));
 sg13g2_a22oi_1 _2564_ (.Y(_1602_),
    .B1(_1331_),
    .B2(_1601_),
    .A2(_0394_),
    .A1(net95));
 sg13g2_nor2_1 _2565_ (.A(_0986_),
    .B(_0185_),
    .Y(_1603_));
 sg13g2_o21ai_1 _2566_ (.B1(_0185_),
    .Y(_1604_),
    .A1(net91),
    .A2(net116));
 sg13g2_a221oi_1 _2567_ (.B2(_1512_),
    .C1(net111),
    .B1(_1604_),
    .A1(_0394_),
    .Y(_1605_),
    .A2(_1603_));
 sg13g2_o21ai_1 _2568_ (.B1(_1605_),
    .Y(_1606_),
    .A1(_1512_),
    .A2(_1602_));
 sg13g2_xor2_1 _2569_ (.B(net98),
    .A(_1610_),
    .X(_1607_));
 sg13g2_nand4_1 _2570_ (.B(net91),
    .C(net101),
    .A(net118),
    .Y(_1608_),
    .D(_1607_));
 sg13g2_and2_1 _2571_ (.A(_1606_),
    .B(_1608_),
    .X(_1609_));
 sg13g2_nor2_1 _2572_ (.A(net101),
    .B(_1598_),
    .Y(_1611_));
 sg13g2_nand2_1 _2573_ (.Y(_1612_),
    .A(net98),
    .B(_1593_));
 sg13g2_and3_1 _2574_ (.X(_1613_),
    .A(net85),
    .B(_1606_),
    .C(_1608_));
 sg13g2_a221oi_1 _2575_ (.B2(_1612_),
    .C1(_1613_),
    .B1(_1611_),
    .A1(_1600_),
    .Y(_1614_),
    .A2(_1609_));
 sg13g2_buf_2 _2576_ (.A(_1614_),
    .X(_1615_));
 sg13g2_a21oi_1 _2577_ (.A1(net115),
    .A2(_1589_),
    .Y(_1616_),
    .B1(net100));
 sg13g2_buf_1 _2578_ (.A(_1090_),
    .X(_1617_));
 sg13g2_o21ai_1 _2579_ (.B1(_1433_),
    .Y(_1618_),
    .A1(net80),
    .A2(_1595_));
 sg13g2_nor2_1 _2580_ (.A(_1512_),
    .B(net93),
    .Y(_1619_));
 sg13g2_o21ai_1 _2581_ (.B1(_1619_),
    .Y(_1620_),
    .A1(_1616_),
    .A2(_1618_));
 sg13g2_nand2_1 _2582_ (.Y(_1622_),
    .A(net100),
    .B(_1595_));
 sg13g2_nand4_1 _2583_ (.B(_1090_),
    .C(net115),
    .A(net99),
    .Y(_1623_),
    .D(_1589_));
 sg13g2_a21oi_1 _2584_ (.A1(_1622_),
    .A2(_1623_),
    .Y(_1624_),
    .B1(net103));
 sg13g2_nor2_1 _2585_ (.A(net99),
    .B(net80),
    .Y(_1625_));
 sg13g2_o21ai_1 _2586_ (.B1(net83),
    .Y(_1626_),
    .A1(_1624_),
    .A2(_1625_));
 sg13g2_nand2_1 _2587_ (.Y(_1627_),
    .A(_1620_),
    .B(_1626_));
 sg13g2_nand3_1 _2588_ (.B(_1615_),
    .C(_1627_),
    .A(net102),
    .Y(_1628_));
 sg13g2_buf_2 _2589_ (.A(_1628_),
    .X(_1629_));
 sg13g2_buf_1 _2590_ (.A(_0394_),
    .X(_1630_));
 sg13g2_buf_1 _2591_ (.A(_0174_),
    .X(_1631_));
 sg13g2_nor2_2 _2592_ (.A(net79),
    .B(net78),
    .Y(_1633_));
 sg13g2_o21ai_1 _2593_ (.B1(_1633_),
    .Y(_1634_),
    .A1(_1615_),
    .A2(_1627_));
 sg13g2_buf_2 _2594_ (.A(_1634_),
    .X(_1635_));
 sg13g2_nor2_1 _2595_ (.A(_1742_),
    .B(_1616_),
    .Y(_1636_));
 sg13g2_o21ai_1 _2596_ (.B1(_1742_),
    .Y(_1637_),
    .A1(_1090_),
    .A2(_1595_));
 sg13g2_nand2_1 _2597_ (.Y(_1638_),
    .A(_1433_),
    .B(_1637_));
 sg13g2_nor2_1 _2598_ (.A(_1512_),
    .B(_1129_),
    .Y(_1639_));
 sg13g2_o21ai_1 _2599_ (.B1(_1639_),
    .Y(_1640_),
    .A1(_1636_),
    .A2(_1638_));
 sg13g2_o21ai_1 _2600_ (.B1(_1090_),
    .Y(_1641_),
    .A1(_0394_),
    .A2(_0372_));
 sg13g2_a22oi_1 _2601_ (.Y(_1642_),
    .B1(net90),
    .B2(net100),
    .A2(_1621_),
    .A1(_1731_));
 sg13g2_nand2_1 _2602_ (.Y(_1644_),
    .A(_1265_),
    .B(_1621_));
 sg13g2_o21ai_1 _2603_ (.B1(_1644_),
    .Y(_1645_),
    .A1(_0987_),
    .A2(_1642_));
 sg13g2_nor3_1 _2604_ (.A(net93),
    .B(_1641_),
    .C(_1645_),
    .Y(_1646_));
 sg13g2_and3_1 _2605_ (.X(_1647_),
    .A(net99),
    .B(_1742_),
    .C(_1645_));
 sg13g2_nor2_1 _2606_ (.A(_0075_),
    .B(_1300_),
    .Y(_1648_));
 sg13g2_o21ai_1 _2607_ (.B1(_1648_),
    .Y(_1649_),
    .A1(_1646_),
    .A2(_1647_));
 sg13g2_nand3_1 _2608_ (.B(net103),
    .C(net83),
    .A(net96),
    .Y(_1650_));
 sg13g2_and3_1 _2609_ (.X(_1651_),
    .A(_1640_),
    .B(_1649_),
    .C(_1650_));
 sg13g2_buf_1 _2610_ (.A(_1651_),
    .X(_1652_));
 sg13g2_nor2_1 _2611_ (.A(net80),
    .B(net78),
    .Y(_1653_));
 sg13g2_buf_2 _2612_ (.A(_1653_),
    .X(_1655_));
 sg13g2_xnor2_1 _2613_ (.Y(_1656_),
    .A(_1652_),
    .B(_1655_));
 sg13g2_a21oi_2 _2614_ (.B1(_1656_),
    .Y(_1657_),
    .A2(_1635_),
    .A1(_1629_));
 sg13g2_and3_1 _2615_ (.X(_1658_),
    .A(_1629_),
    .B(_1635_),
    .C(_1656_));
 sg13g2_buf_1 _2616_ (.A(_1658_),
    .X(_1659_));
 sg13g2_or2_1 _2617_ (.X(_1660_),
    .B(_1659_),
    .A(_1657_));
 sg13g2_buf_1 _2618_ (.A(_1660_),
    .X(_1661_));
 sg13g2_buf_1 _2619_ (.A(_1627_),
    .X(_1662_));
 sg13g2_nor2_1 _2620_ (.A(net79),
    .B(_1154_),
    .Y(_1663_));
 sg13g2_nand2_1 _2621_ (.Y(_1664_),
    .A(net94),
    .B(net102));
 sg13g2_nand2_1 _2622_ (.Y(_1666_),
    .A(net79),
    .B(net102));
 sg13g2_mux2_1 _2623_ (.A0(_1664_),
    .A1(_1666_),
    .S(_1615_),
    .X(_1667_));
 sg13g2_buf_2 _2624_ (.A(_1667_),
    .X(_1668_));
 sg13g2_nand3_1 _2625_ (.B(_1663_),
    .C(_1668_),
    .A(net33),
    .Y(_1669_));
 sg13g2_buf_1 _2626_ (.A(net117),
    .X(_1670_));
 sg13g2_nand2_1 _2627_ (.Y(_1671_),
    .A(net94),
    .B(net97));
 sg13g2_or3_1 _2628_ (.A(net33),
    .B(_1671_),
    .C(_1668_),
    .X(_1672_));
 sg13g2_nor2_1 _2629_ (.A(_1512_),
    .B(net79),
    .Y(_1673_));
 sg13g2_nand3_1 _2630_ (.B(_1206_),
    .C(_1589_),
    .A(net98),
    .Y(_1674_));
 sg13g2_nor2b_1 _2631_ (.A(net101),
    .B_N(net118),
    .Y(_1675_));
 sg13g2_nor2b_1 _2632_ (.A(net90),
    .B_N(net116),
    .Y(_1677_));
 sg13g2_buf_1 _2633_ (.A(_1677_),
    .X(_1678_));
 sg13g2_a21oi_1 _2634_ (.A1(_0622_),
    .A2(_1675_),
    .Y(_1679_),
    .B1(_1678_));
 sg13g2_nand2_1 _2635_ (.Y(_1680_),
    .A(_1512_),
    .B(net101));
 sg13g2_o21ai_1 _2636_ (.B1(_1680_),
    .Y(_1681_),
    .A1(net115),
    .A2(_1679_));
 sg13g2_a22oi_1 _2637_ (.Y(_1682_),
    .B1(_1681_),
    .B2(net98),
    .A2(_1674_),
    .A1(_1673_));
 sg13g2_nor2b_2 _2638_ (.A(net116),
    .B_N(_1082_),
    .Y(_1683_));
 sg13g2_nand3b_1 _2639_ (.B(_1184_),
    .C(_0970_),
    .Y(_1684_),
    .A_N(net90));
 sg13g2_nand2b_1 _2640_ (.Y(_1685_),
    .B(_1684_),
    .A_N(_1683_));
 sg13g2_o21ai_1 _2641_ (.B1(_0970_),
    .Y(_1686_),
    .A1(net118),
    .A2(net98));
 sg13g2_a22oi_1 _2642_ (.Y(_1688_),
    .B1(_1686_),
    .B2(net90),
    .A2(_1685_),
    .A1(net99));
 sg13g2_nor2_1 _2643_ (.A(_1631_),
    .B(_1688_),
    .Y(_1689_));
 sg13g2_xnor2_1 _2644_ (.Y(_1690_),
    .A(_1682_),
    .B(_1689_));
 sg13g2_nand2_1 _2645_ (.Y(_1691_),
    .A(net85),
    .B(net102));
 sg13g2_nand3_1 _2646_ (.B(net102),
    .C(_1608_),
    .A(net101),
    .Y(_1692_));
 sg13g2_mux2_1 _2647_ (.A0(_1691_),
    .A1(_1692_),
    .S(_1606_),
    .X(_1693_));
 sg13g2_xor2_1 _2648_ (.B(_1693_),
    .A(_1600_),
    .X(_1694_));
 sg13g2_buf_2 _2649_ (.A(_1694_),
    .X(_1695_));
 sg13g2_a21o_1 _2650_ (.A2(_1690_),
    .A1(net91),
    .B1(_1695_),
    .X(_1696_));
 sg13g2_buf_1 _2651_ (.A(_1690_),
    .X(_1697_));
 sg13g2_and3_1 _2652_ (.X(_1699_),
    .A(net66),
    .B(_1695_),
    .C(net31));
 sg13g2_a21oi_2 _2653_ (.B1(_1699_),
    .Y(_1700_),
    .A2(_1696_),
    .A1(net90));
 sg13g2_a21oi_2 _2654_ (.B1(_1700_),
    .Y(_1701_),
    .A2(_1672_),
    .A1(_1669_));
 sg13g2_nand2_1 _2655_ (.Y(_1702_),
    .A(net101),
    .B(_1663_));
 sg13g2_or2_1 _2656_ (.X(_1703_),
    .B(_1702_),
    .A(net33));
 sg13g2_nand2b_1 _2657_ (.Y(_1704_),
    .B(_1662_),
    .A_N(_1702_));
 sg13g2_mux2_1 _2658_ (.A0(_1703_),
    .A1(_1704_),
    .S(_1668_),
    .X(_1705_));
 sg13g2_o21ai_1 _2659_ (.B1(_1705_),
    .Y(_1706_),
    .A1(_1700_),
    .A2(_1702_));
 sg13g2_buf_1 _2660_ (.A(_1706_),
    .X(_1707_));
 sg13g2_nor3_2 _2661_ (.A(_1661_),
    .B(_1701_),
    .C(_1707_),
    .Y(_1708_));
 sg13g2_and4_1 _2662_ (.A(net85),
    .B(_1620_),
    .C(_1626_),
    .D(_1668_),
    .X(_1710_));
 sg13g2_nand2_1 _2663_ (.Y(_1711_),
    .A(net85),
    .B(_1627_));
 sg13g2_nor2_1 _2664_ (.A(_1668_),
    .B(_1711_),
    .Y(_1712_));
 sg13g2_or4_1 _2665_ (.A(net89),
    .B(_1700_),
    .C(_1710_),
    .D(_1712_),
    .X(_1713_));
 sg13g2_buf_1 _2666_ (.A(_1713_),
    .X(_1714_));
 sg13g2_xnor2_1 _2667_ (.Y(_1715_),
    .A(_1662_),
    .B(_1668_));
 sg13g2_nor2_1 _2668_ (.A(net85),
    .B(_1155_),
    .Y(_1716_));
 sg13g2_nand2_1 _2669_ (.Y(_1717_),
    .A(_1715_),
    .B(_1716_));
 sg13g2_and3_1 _2670_ (.X(_1718_),
    .A(_1671_),
    .B(_1714_),
    .C(_1717_));
 sg13g2_buf_2 _2671_ (.A(_1718_),
    .X(_1719_));
 sg13g2_nand3_1 _2672_ (.B(_1649_),
    .C(_1650_),
    .A(_1640_),
    .Y(_1721_));
 sg13g2_buf_1 _2673_ (.A(_1721_),
    .X(_1722_));
 sg13g2_a22oi_1 _2674_ (.Y(_1723_),
    .B1(_1722_),
    .B2(_1655_),
    .A2(_1633_),
    .A1(net33));
 sg13g2_nand2_1 _2675_ (.Y(_1724_),
    .A(_1615_),
    .B(_1633_));
 sg13g2_o21ai_1 _2676_ (.B1(_1129_),
    .Y(_1725_),
    .A1(net93),
    .A2(_1616_));
 sg13g2_a21oi_1 _2677_ (.A1(_0075_),
    .A2(_1637_),
    .Y(_1726_),
    .B1(_1300_));
 sg13g2_nand2_1 _2678_ (.Y(_1727_),
    .A(net99),
    .B(net114));
 sg13g2_a21oi_1 _2679_ (.A1(_1725_),
    .A2(_1726_),
    .Y(_1728_),
    .B1(_1727_));
 sg13g2_a21o_1 _2680_ (.A2(_1589_),
    .A1(net115),
    .B1(_1265_),
    .X(_1729_));
 sg13g2_nand2_1 _2681_ (.Y(_1730_),
    .A(_1124_),
    .B(_1729_));
 sg13g2_nand3_1 _2682_ (.B(net108),
    .C(_1648_),
    .A(net99),
    .Y(_1732_));
 sg13g2_nor2_1 _2683_ (.A(net99),
    .B(_1129_),
    .Y(_1733_));
 sg13g2_nor2b_1 _2684_ (.A(net114),
    .B_N(net98),
    .Y(_1734_));
 sg13g2_and2_1 _2685_ (.A(_0075_),
    .B(_1734_),
    .X(_1735_));
 sg13g2_a21o_1 _2686_ (.A2(_1082_),
    .A1(_1184_),
    .B1(net115),
    .X(_1736_));
 sg13g2_a21oi_1 _2687_ (.A1(net100),
    .A2(_1736_),
    .Y(_1737_),
    .B1(net103));
 sg13g2_a22oi_1 _2688_ (.Y(_1738_),
    .B1(_1735_),
    .B2(_1737_),
    .A2(_1733_),
    .A1(net83));
 sg13g2_o21ai_1 _2689_ (.B1(_1738_),
    .Y(_1739_),
    .A1(_1730_),
    .A2(_1732_));
 sg13g2_nor2_1 _2690_ (.A(net93),
    .B(net78),
    .Y(_1740_));
 sg13g2_o21ai_1 _2691_ (.B1(_1740_),
    .Y(_1741_),
    .A1(_1728_),
    .A2(_1739_));
 sg13g2_or3_1 _2692_ (.A(_1728_),
    .B(_1739_),
    .C(_1740_),
    .X(_1743_));
 sg13g2_nand2_1 _2693_ (.Y(_1744_),
    .A(net100),
    .B(net117));
 sg13g2_a21oi_1 _2694_ (.A1(_1741_),
    .A2(_1743_),
    .Y(_1745_),
    .B1(_1744_));
 sg13g2_nand4_1 _2695_ (.B(_1723_),
    .C(_1724_),
    .A(_1629_),
    .Y(_1746_),
    .D(_1745_));
 sg13g2_nand2_1 _2696_ (.Y(_1747_),
    .A(net87),
    .B(net102));
 sg13g2_and3_1 _2697_ (.X(_1748_),
    .A(_1744_),
    .B(_1741_),
    .C(_1743_));
 sg13g2_buf_1 _2698_ (.A(_1748_),
    .X(_1749_));
 sg13g2_nand4_1 _2699_ (.B(_1635_),
    .C(_1747_),
    .A(_1629_),
    .Y(_1750_),
    .D(_1749_));
 sg13g2_nor2_1 _2700_ (.A(net80),
    .B(net89),
    .Y(_1751_));
 sg13g2_and2_1 _2701_ (.A(_1741_),
    .B(_1743_),
    .X(_1752_));
 sg13g2_buf_1 _2702_ (.A(_1752_),
    .X(_1754_));
 sg13g2_or4_1 _2703_ (.A(_1635_),
    .B(_1652_),
    .C(_1751_),
    .D(_1754_),
    .X(_1755_));
 sg13g2_nor2_1 _2704_ (.A(_1722_),
    .B(_1751_),
    .Y(_1756_));
 sg13g2_nand4_1 _2705_ (.B(_1635_),
    .C(_1754_),
    .A(_1629_),
    .Y(_1757_),
    .D(_1756_));
 sg13g2_nand4_1 _2706_ (.B(_1750_),
    .C(_1755_),
    .A(_1746_),
    .Y(_1758_),
    .D(_1757_));
 sg13g2_nor2_1 _2707_ (.A(_1722_),
    .B(_1655_),
    .Y(_1759_));
 sg13g2_o21ai_1 _2708_ (.B1(_1759_),
    .Y(_1760_),
    .A1(_1745_),
    .A2(_1749_));
 sg13g2_or3_1 _2709_ (.A(_1759_),
    .B(_1745_),
    .C(_1749_),
    .X(_1761_));
 sg13g2_nor2_1 _2710_ (.A(_1722_),
    .B(_1747_),
    .Y(_1762_));
 sg13g2_nor2_1 _2711_ (.A(_1652_),
    .B(_1655_),
    .Y(_1763_));
 sg13g2_a21o_1 _2712_ (.A2(_1762_),
    .A1(_1635_),
    .B1(_1763_),
    .X(_1765_));
 sg13g2_a22oi_1 _2713_ (.Y(_1766_),
    .B1(_1765_),
    .B2(_1629_),
    .A2(_1761_),
    .A1(_1760_));
 sg13g2_nor2_1 _2714_ (.A(_1758_),
    .B(_1766_),
    .Y(_1767_));
 sg13g2_or3_1 _2715_ (.A(_1708_),
    .B(_1719_),
    .C(_1767_),
    .X(_1768_));
 sg13g2_buf_1 _2716_ (.A(_1768_),
    .X(_1769_));
 sg13g2_o21ai_1 _2717_ (.B1(_1767_),
    .Y(_1770_),
    .A1(_1708_),
    .A2(_1719_));
 sg13g2_buf_1 _2718_ (.A(_1770_),
    .X(_1771_));
 sg13g2_and2_1 _2719_ (.A(_1769_),
    .B(_1771_),
    .X(_1772_));
 sg13g2_buf_1 _2720_ (.A(_1772_),
    .X(_1773_));
 sg13g2_buf_1 _2721_ (.A(net105),
    .X(_1774_));
 sg13g2_a21oi_1 _2722_ (.A1(net66),
    .A2(net31),
    .Y(_1776_),
    .B1(_1695_));
 sg13g2_nor2_1 _2723_ (.A(net88),
    .B(_1155_),
    .Y(_1777_));
 sg13g2_a22oi_1 _2724_ (.Y(_1778_),
    .B1(_1777_),
    .B2(_1699_),
    .A2(_1716_),
    .A1(_1776_));
 sg13g2_buf_1 _2725_ (.A(_1778_),
    .X(_1779_));
 sg13g2_nand2_1 _2726_ (.Y(_1780_),
    .A(net117),
    .B(_1678_));
 sg13g2_a21oi_1 _2727_ (.A1(net66),
    .A2(net31),
    .Y(_1781_),
    .B1(_1780_));
 sg13g2_and2_1 _2728_ (.A(net117),
    .B(_1683_),
    .X(_1782_));
 sg13g2_and3_1 _2729_ (.X(_1783_),
    .A(net66),
    .B(net31),
    .C(_1782_));
 sg13g2_nor2_1 _2730_ (.A(_1695_),
    .B(_1780_),
    .Y(_1784_));
 sg13g2_and2_1 _2731_ (.A(_1695_),
    .B(_1782_),
    .X(_1785_));
 sg13g2_nor4_2 _2732_ (.A(_1781_),
    .B(_1783_),
    .C(_1784_),
    .Y(_0021_),
    .D(_1785_));
 sg13g2_and3_1 _2733_ (.X(_0022_),
    .A(_1715_),
    .B(_1779_),
    .C(_0021_));
 sg13g2_buf_1 _2734_ (.A(_0022_),
    .X(_0023_));
 sg13g2_a21oi_2 _2735_ (.B1(_1715_),
    .Y(_0024_),
    .A2(_0021_),
    .A1(_1779_));
 sg13g2_nand2_1 _2736_ (.Y(_0025_),
    .A(net64),
    .B(net117));
 sg13g2_nand2_1 _2737_ (.Y(_0026_),
    .A(_0460_),
    .B(net117));
 sg13g2_mux2_1 _2738_ (.A0(_0025_),
    .A1(_0026_),
    .S(net31),
    .X(_0027_));
 sg13g2_xor2_1 _2739_ (.B(_0027_),
    .A(_1695_),
    .X(_0028_));
 sg13g2_nor2_1 _2740_ (.A(net69),
    .B(_0028_),
    .Y(_0029_));
 sg13g2_nor3_1 _2741_ (.A(_0023_),
    .B(_0024_),
    .C(_0029_),
    .Y(_0030_));
 sg13g2_o21ai_1 _2742_ (.B1(_0029_),
    .Y(_0032_),
    .A1(_0023_),
    .A2(_0024_));
 sg13g2_o21ai_1 _2743_ (.B1(_0032_),
    .Y(_0033_),
    .A1(net86),
    .A2(_0030_));
 sg13g2_buf_2 _2744_ (.A(_0033_),
    .X(_0034_));
 sg13g2_or3_1 _2745_ (.A(_1657_),
    .B(_1659_),
    .C(_1671_),
    .X(_0035_));
 sg13g2_o21ai_1 _2746_ (.B1(_1671_),
    .Y(_0036_),
    .A1(_1657_),
    .A2(_1659_));
 sg13g2_and4_1 _2747_ (.A(_1714_),
    .B(_1717_),
    .C(_0035_),
    .D(_0036_),
    .X(_0037_));
 sg13g2_buf_1 _2748_ (.A(_0037_),
    .X(_0038_));
 sg13g2_a22oi_1 _2749_ (.Y(_0039_),
    .B1(_0035_),
    .B2(_0036_),
    .A2(_1717_),
    .A1(_1714_));
 sg13g2_nor2_2 _2750_ (.A(_0038_),
    .B(_0039_),
    .Y(_0040_));
 sg13g2_nand4_1 _2751_ (.B(_1774_),
    .C(_0034_),
    .A(_1630_),
    .Y(_0041_),
    .D(_0040_));
 sg13g2_nand3_1 _2752_ (.B(_1334_),
    .C(_0034_),
    .A(net77),
    .Y(_0043_));
 sg13g2_nand2_1 _2753_ (.Y(_0044_),
    .A(net94),
    .B(net77));
 sg13g2_or3_1 _2754_ (.A(_0034_),
    .B(_0040_),
    .C(_0044_),
    .X(_0045_));
 sg13g2_and4_1 _2755_ (.A(_1773_),
    .B(_0041_),
    .C(_0043_),
    .D(_0045_),
    .X(_0046_));
 sg13g2_nand2_1 _2756_ (.Y(_0047_),
    .A(net77),
    .B(_1331_));
 sg13g2_nor2_1 _2757_ (.A(_0034_),
    .B(_0047_),
    .Y(_0048_));
 sg13g2_and3_1 _2758_ (.X(_0049_),
    .A(net77),
    .B(_1334_),
    .C(_0040_));
 sg13g2_nor2_1 _2759_ (.A(_0040_),
    .B(_0047_),
    .Y(_0050_));
 sg13g2_nor3_1 _2760_ (.A(_0048_),
    .B(_0049_),
    .C(_0050_),
    .Y(_0051_));
 sg13g2_a21oi_1 _2761_ (.A1(_1769_),
    .A2(_1771_),
    .Y(_0052_),
    .B1(_0044_));
 sg13g2_nand2_1 _2762_ (.Y(_0054_),
    .A(_1630_),
    .B(net77));
 sg13g2_a21oi_1 _2763_ (.A1(_1769_),
    .A2(_1771_),
    .Y(_0055_),
    .B1(_0054_));
 sg13g2_o21ai_1 _2764_ (.B1(net85),
    .Y(_0056_),
    .A1(_0038_),
    .A2(_0039_));
 sg13g2_nor3_1 _2765_ (.A(net85),
    .B(_0038_),
    .C(_0039_),
    .Y(_0057_));
 sg13g2_a21o_1 _2766_ (.A2(_0056_),
    .A1(_0034_),
    .B1(_0057_),
    .X(_0058_));
 sg13g2_buf_1 _2767_ (.A(_0058_),
    .X(_0059_));
 sg13g2_mux2_1 _2768_ (.A0(_0052_),
    .A1(_0055_),
    .S(_0059_),
    .X(_0060_));
 sg13g2_a21o_1 _2769_ (.A2(_0051_),
    .A1(_0046_),
    .B1(_0060_),
    .X(_0061_));
 sg13g2_buf_1 _2770_ (.A(_0061_),
    .X(_0062_));
 sg13g2_nand3_1 _2771_ (.B(_1779_),
    .C(_0021_),
    .A(_1715_),
    .Y(_0063_));
 sg13g2_a21o_1 _2772_ (.A2(_0021_),
    .A1(_1779_),
    .B1(_1715_),
    .X(_0065_));
 sg13g2_nor2_1 _2773_ (.A(net86),
    .B(_0878_),
    .Y(_0066_));
 sg13g2_o21ai_1 _2774_ (.B1(_0066_),
    .Y(_0067_),
    .A1(net69),
    .A2(_0028_));
 sg13g2_xnor2_1 _2775_ (.Y(_0068_),
    .A(_1695_),
    .B(_0027_));
 sg13g2_nand4_1 _2776_ (.B(net86),
    .C(net105),
    .A(_1102_),
    .Y(_0069_),
    .D(_0068_));
 sg13g2_a22oi_1 _2777_ (.Y(_0070_),
    .B1(_0067_),
    .B2(_0069_),
    .A2(_0065_),
    .A1(_0063_));
 sg13g2_and4_1 _2778_ (.A(_0063_),
    .B(_0065_),
    .C(_0067_),
    .D(_0069_),
    .X(_0071_));
 sg13g2_nand2_1 _2779_ (.Y(_0072_),
    .A(net49),
    .B(net104));
 sg13g2_nor3_2 _2780_ (.A(_0070_),
    .B(_0071_),
    .C(_0072_),
    .Y(_0073_));
 sg13g2_nand4_1 _2781_ (.B(_1333_),
    .C(net105),
    .A(net49),
    .Y(_0074_),
    .D(_0068_));
 sg13g2_nand2_1 _2782_ (.Y(_0076_),
    .A(net105),
    .B(_1683_));
 sg13g2_a22oi_1 _2783_ (.Y(_0077_),
    .B1(_0074_),
    .B2(_0076_),
    .A2(_0065_),
    .A1(_0063_));
 sg13g2_nand2_1 _2784_ (.Y(_0078_),
    .A(net88),
    .B(net105));
 sg13g2_nor4_1 _2785_ (.A(_0023_),
    .B(_0024_),
    .C(_0029_),
    .D(_0078_),
    .Y(_0079_));
 sg13g2_nand2_1 _2786_ (.Y(_0080_),
    .A(net105),
    .B(_1678_));
 sg13g2_nor3_1 _2787_ (.A(_0023_),
    .B(_0024_),
    .C(_0080_),
    .Y(_0081_));
 sg13g2_a21oi_1 _2788_ (.A1(net49),
    .A2(_0068_),
    .Y(_0082_),
    .B1(_0080_));
 sg13g2_nor3_1 _2789_ (.A(net69),
    .B(_0028_),
    .C(_0076_),
    .Y(_0083_));
 sg13g2_or2_1 _2790_ (.X(_0084_),
    .B(_0083_),
    .A(_0082_));
 sg13g2_nor4_2 _2791_ (.A(_0077_),
    .B(_0079_),
    .C(_0081_),
    .Y(_0085_),
    .D(_0084_));
 sg13g2_xnor2_1 _2792_ (.Y(_0087_),
    .A(_0040_),
    .B(_0085_));
 sg13g2_buf_2 _2793_ (.A(_0087_),
    .X(_0088_));
 sg13g2_nand2_1 _2794_ (.Y(_0089_),
    .A(_0073_),
    .B(_0088_));
 sg13g2_o21ai_1 _2795_ (.B1(_1161_),
    .Y(_0090_),
    .A1(_0073_),
    .A2(_0088_));
 sg13g2_buf_1 _2796_ (.A(_0090_),
    .X(_0091_));
 sg13g2_nand2_1 _2797_ (.Y(_0092_),
    .A(net88),
    .B(net104));
 sg13g2_a21oi_2 _2798_ (.B1(_0092_),
    .Y(_0093_),
    .A2(_0091_),
    .A1(_0089_));
 sg13g2_a21oi_1 _2799_ (.A1(_0073_),
    .A2(_0088_),
    .Y(_0094_),
    .B1(net88));
 sg13g2_buf_1 _2800_ (.A(_1019_),
    .X(_0095_));
 sg13g2_a21o_1 _2801_ (.A2(_0094_),
    .A1(_0091_),
    .B1(net60),
    .X(_0096_));
 sg13g2_buf_1 _2802_ (.A(_0096_),
    .X(_0098_));
 sg13g2_nor2_1 _2803_ (.A(_0093_),
    .B(_0098_),
    .Y(_0099_));
 sg13g2_xnor2_1 _2804_ (.Y(_0100_),
    .A(_0062_),
    .B(_0099_));
 sg13g2_nand2_1 _2805_ (.Y(_0101_),
    .A(_1161_),
    .B(net104));
 sg13g2_xor2_1 _2806_ (.B(_0101_),
    .A(_0073_),
    .X(_0102_));
 sg13g2_nor2_1 _2807_ (.A(_1567_),
    .B(net110),
    .Y(_0103_));
 sg13g2_xor2_1 _2808_ (.B(_0085_),
    .A(_0040_),
    .X(_0104_));
 sg13g2_nand3b_1 _2809_ (.B(_0103_),
    .C(_0104_),
    .Y(_0105_),
    .A_N(_0102_));
 sg13g2_nand3_1 _2810_ (.B(_0103_),
    .C(_0102_),
    .A(_0088_),
    .Y(_0106_));
 sg13g2_nand2_1 _2811_ (.Y(_0107_),
    .A(_0105_),
    .B(_0106_));
 sg13g2_buf_2 _2812_ (.A(_0107_),
    .X(_0109_));
 sg13g2_nand2_1 _2813_ (.Y(_0110_),
    .A(_1461_),
    .B(_0951_));
 sg13g2_xor2_1 _2814_ (.B(_0110_),
    .A(_0109_),
    .X(_0111_));
 sg13g2_xnor2_1 _2815_ (.Y(_0112_),
    .A(_0100_),
    .B(_0111_));
 sg13g2_nor2_1 _2816_ (.A(_1299_),
    .B(net122),
    .Y(_0113_));
 sg13g2_a21oi_1 _2817_ (.A1(_1586_),
    .A2(_0112_),
    .Y(_0114_),
    .B1(_0113_));
 sg13g2_nor2_1 _2818_ (.A(_1661_),
    .B(_1751_),
    .Y(_0115_));
 sg13g2_nor2_1 _2819_ (.A(_1701_),
    .B(_1707_),
    .Y(_0116_));
 sg13g2_nand2_1 _2820_ (.Y(_0117_),
    .A(_1722_),
    .B(_1655_));
 sg13g2_nand3_1 _2821_ (.B(net33),
    .C(_1655_),
    .A(_1615_),
    .Y(_0118_));
 sg13g2_nand3_1 _2822_ (.B(_1633_),
    .C(_1655_),
    .A(_1615_),
    .Y(_0120_));
 sg13g2_nand3_1 _2823_ (.B(_1633_),
    .C(_1655_),
    .A(net33),
    .Y(_0121_));
 sg13g2_and4_1 _2824_ (.A(_0117_),
    .B(_0118_),
    .C(_0120_),
    .D(_0121_),
    .X(_0122_));
 sg13g2_buf_1 _2825_ (.A(_0122_),
    .X(_0123_));
 sg13g2_or2_1 _2826_ (.X(_0124_),
    .B(net33),
    .A(_1615_));
 sg13g2_nor2_1 _2827_ (.A(_1664_),
    .B(_1652_),
    .Y(_0125_));
 sg13g2_and4_1 _2828_ (.A(net102),
    .B(_1615_),
    .C(net33),
    .D(_1722_),
    .X(_0126_));
 sg13g2_a21oi_2 _2829_ (.B1(_0126_),
    .Y(_0127_),
    .A2(_0125_),
    .A1(_0124_));
 sg13g2_a21oi_1 _2830_ (.A1(_0123_),
    .A2(_0127_),
    .Y(_0128_),
    .B1(_1754_));
 sg13g2_and3_1 _2831_ (.X(_0129_),
    .A(_1754_),
    .B(_0123_),
    .C(_0127_));
 sg13g2_buf_1 _2832_ (.A(_0129_),
    .X(_0131_));
 sg13g2_nor3_1 _2833_ (.A(_1751_),
    .B(_0128_),
    .C(_0131_),
    .Y(_0132_));
 sg13g2_a221oi_1 _2834_ (.B2(_0116_),
    .C1(_0132_),
    .B1(_0115_),
    .A1(_1719_),
    .Y(_0133_),
    .A2(_1744_));
 sg13g2_buf_2 _2835_ (.A(_0133_),
    .X(_0134_));
 sg13g2_nor2_1 _2836_ (.A(_0128_),
    .B(_0131_),
    .Y(_0135_));
 sg13g2_nor4_1 _2837_ (.A(_1701_),
    .B(_1707_),
    .C(_0128_),
    .D(_0131_),
    .Y(_0136_));
 sg13g2_nor2_1 _2838_ (.A(_1657_),
    .B(_1659_),
    .Y(_0137_));
 sg13g2_a22oi_1 _2839_ (.Y(_0138_),
    .B1(_0136_),
    .B2(_0137_),
    .A2(_0135_),
    .A1(_1719_));
 sg13g2_buf_1 _2840_ (.A(_0138_),
    .X(_0139_));
 sg13g2_nand2_1 _2841_ (.Y(_0140_),
    .A(_0134_),
    .B(_0139_));
 sg13g2_nor2_1 _2842_ (.A(_1728_),
    .B(_1739_),
    .Y(_0142_));
 sg13g2_buf_1 _2843_ (.A(_0142_),
    .X(_0143_));
 sg13g2_inv_1 _2844_ (.Y(_0144_),
    .A(net32));
 sg13g2_nand3_1 _2845_ (.B(_0123_),
    .C(_0127_),
    .A(net93),
    .Y(_0145_));
 sg13g2_nand2_1 _2846_ (.Y(_0146_),
    .A(_1129_),
    .B(net83));
 sg13g2_nor2_1 _2847_ (.A(_1129_),
    .B(_1737_),
    .Y(_0147_));
 sg13g2_a22oi_1 _2848_ (.Y(_0148_),
    .B1(_0147_),
    .B2(_1734_),
    .A2(_0146_),
    .A1(net68));
 sg13g2_nand3_1 _2849_ (.B(net114),
    .C(net83),
    .A(net96),
    .Y(_0149_));
 sg13g2_o21ai_1 _2850_ (.B1(_0149_),
    .Y(_0150_),
    .A1(net96),
    .A2(_0148_));
 sg13g2_nor3_1 _2851_ (.A(net129),
    .B(_1636_),
    .C(_0146_),
    .Y(_0151_));
 sg13g2_a22oi_1 _2852_ (.Y(_0153_),
    .B1(_1637_),
    .B2(_0086_),
    .A2(_1729_),
    .A1(net103));
 sg13g2_nor3_1 _2853_ (.A(net96),
    .B(net120),
    .C(_0153_),
    .Y(_0154_));
 sg13g2_o21ai_1 _2854_ (.B1(net114),
    .Y(_0155_),
    .A1(_0151_),
    .A2(_0154_));
 sg13g2_nor2b_1 _2855_ (.A(_0150_),
    .B_N(_0155_),
    .Y(_0156_));
 sg13g2_buf_1 _2856_ (.A(_0156_),
    .X(_0157_));
 sg13g2_inv_1 _2857_ (.Y(_0158_),
    .A(_0157_));
 sg13g2_nand3_1 _2858_ (.B(_1144_),
    .C(_0158_),
    .A(net113),
    .Y(_0159_));
 sg13g2_buf_1 _2859_ (.A(_1129_),
    .X(_0160_));
 sg13g2_nand2_1 _2860_ (.Y(_0161_),
    .A(net76),
    .B(_0157_));
 sg13g2_a21oi_1 _2861_ (.A1(_0123_),
    .A2(_0127_),
    .Y(_0162_),
    .B1(net93));
 sg13g2_a221oi_1 _2862_ (.B2(_0161_),
    .C1(_0162_),
    .B1(_0159_),
    .A1(_0144_),
    .Y(_0164_),
    .A2(_0145_));
 sg13g2_nor2_1 _2863_ (.A(net113),
    .B(net78),
    .Y(_0165_));
 sg13g2_nand2_1 _2864_ (.Y(_0166_),
    .A(_0158_),
    .B(_0165_));
 sg13g2_nand2_1 _2865_ (.Y(_0167_),
    .A(net113),
    .B(_0157_));
 sg13g2_nand4_1 _2866_ (.B(_0118_),
    .C(_0120_),
    .A(_0117_),
    .Y(_0168_),
    .D(_0121_));
 sg13g2_a21o_1 _2867_ (.A2(_0125_),
    .A1(_0124_),
    .B1(_0126_),
    .X(_0169_));
 sg13g2_buf_1 _2868_ (.A(_0169_),
    .X(_0170_));
 sg13g2_buf_1 _2869_ (.A(net103),
    .X(_0171_));
 sg13g2_o21ai_1 _2870_ (.B1(net75),
    .Y(_0172_),
    .A1(_0168_),
    .A2(_0170_));
 sg13g2_a21oi_1 _2871_ (.A1(_0166_),
    .A2(_0167_),
    .Y(_0173_),
    .B1(_0172_));
 sg13g2_and4_1 _2872_ (.A(_0144_),
    .B(_0158_),
    .C(_0145_),
    .D(_0165_),
    .X(_0175_));
 sg13g2_nor3_2 _2873_ (.A(_0164_),
    .B(_0173_),
    .C(_0175_),
    .Y(_0176_));
 sg13g2_buf_1 _2874_ (.A(_0157_),
    .X(_0177_));
 sg13g2_buf_1 _2875_ (.A(net113),
    .X(_0178_));
 sg13g2_and4_1 _2876_ (.A(net74),
    .B(_0144_),
    .C(net30),
    .D(_0145_),
    .X(_0179_));
 sg13g2_a21oi_2 _2877_ (.B1(_0179_),
    .Y(_0180_),
    .A2(net30),
    .A1(net78));
 sg13g2_nand2_1 _2878_ (.Y(_0181_),
    .A(net75),
    .B(net97));
 sg13g2_a21o_1 _2879_ (.A2(_0180_),
    .A1(_0176_),
    .B1(_0181_),
    .X(_0182_));
 sg13g2_nand3_1 _2880_ (.B(_0180_),
    .C(_0181_),
    .A(_0176_),
    .Y(_0183_));
 sg13g2_nand3_1 _2881_ (.B(_0182_),
    .C(_0183_),
    .A(_0140_),
    .Y(_0184_));
 sg13g2_a21o_1 _2882_ (.A2(_0183_),
    .A1(_0182_),
    .B1(_0140_),
    .X(_0186_));
 sg13g2_nand2_1 _2883_ (.Y(_0187_),
    .A(_0184_),
    .B(_0186_));
 sg13g2_a21oi_1 _2884_ (.A1(_0034_),
    .A2(_0056_),
    .Y(_0188_),
    .B1(_0057_));
 sg13g2_or4_1 _2885_ (.A(net94),
    .B(_1708_),
    .C(_1719_),
    .D(_1767_),
    .X(_0189_));
 sg13g2_nor3_1 _2886_ (.A(_1632_),
    .B(_1758_),
    .C(_1766_),
    .Y(_0190_));
 sg13g2_o21ai_1 _2887_ (.B1(_0190_),
    .Y(_0191_),
    .A1(_1708_),
    .A2(_1719_));
 sg13g2_nand2_1 _2888_ (.Y(_0192_),
    .A(_0189_),
    .B(_0191_));
 sg13g2_nor4_1 _2889_ (.A(net87),
    .B(_0878_),
    .C(_0188_),
    .D(_0192_),
    .Y(_0193_));
 sg13g2_or3_1 _2890_ (.A(_1661_),
    .B(_1701_),
    .C(_1707_),
    .X(_0194_));
 sg13g2_nand3_1 _2891_ (.B(_1714_),
    .C(_1717_),
    .A(_1671_),
    .Y(_0195_));
 sg13g2_o21ai_1 _2892_ (.B1(_1632_),
    .Y(_0197_),
    .A1(_1758_),
    .A2(_1766_));
 sg13g2_a21oi_1 _2893_ (.A1(_0194_),
    .A2(_0195_),
    .Y(_0198_),
    .B1(_0197_));
 sg13g2_and4_1 _2894_ (.A(net94),
    .B(net97),
    .C(_0194_),
    .D(_1767_),
    .X(_0199_));
 sg13g2_nand2_1 _2895_ (.Y(_0200_),
    .A(net87),
    .B(net77));
 sg13g2_nor3_1 _2896_ (.A(_0198_),
    .B(_0199_),
    .C(_0200_),
    .Y(_0201_));
 sg13g2_a21oi_1 _2897_ (.A1(_0189_),
    .A2(_0191_),
    .Y(_0202_),
    .B1(_0200_));
 sg13g2_a21oi_1 _2898_ (.A1(_0188_),
    .A2(_0201_),
    .Y(_0203_),
    .B1(_0202_));
 sg13g2_nand4_1 _2899_ (.B(net63),
    .C(net77),
    .A(net80),
    .Y(_0204_),
    .D(_1773_));
 sg13g2_nand3b_1 _2900_ (.B(_0203_),
    .C(_0204_),
    .Y(_0205_),
    .A_N(_0193_));
 sg13g2_xnor2_1 _2901_ (.Y(_0206_),
    .A(_0187_),
    .B(_0205_));
 sg13g2_buf_2 _2902_ (.A(_0206_),
    .X(_0208_));
 sg13g2_a21oi_2 _2903_ (.B1(_0060_),
    .Y(_0209_),
    .A2(_0051_),
    .A1(_0046_));
 sg13g2_buf_1 _2904_ (.A(_0209_),
    .X(_0210_));
 sg13g2_or2_1 _2905_ (.X(_0211_),
    .B(_0071_),
    .A(_0070_));
 sg13g2_or2_1 _2906_ (.X(_0212_),
    .B(_0072_),
    .A(_0211_));
 sg13g2_buf_1 _2907_ (.A(_0212_),
    .X(_0213_));
 sg13g2_nand2_1 _2908_ (.Y(_0214_),
    .A(_0213_),
    .B(_0104_));
 sg13g2_o21ai_1 _2909_ (.B1(_0101_),
    .Y(_0215_),
    .A1(_0213_),
    .A2(_0104_));
 sg13g2_nand2_1 _2910_ (.Y(_0216_),
    .A(_0214_),
    .B(_0215_));
 sg13g2_or4_1 _2911_ (.A(net63),
    .B(net60),
    .C(net28),
    .D(_0216_),
    .X(_0217_));
 sg13g2_buf_1 _2912_ (.A(net104),
    .X(_0219_));
 sg13g2_nand4_1 _2913_ (.B(net73),
    .C(net28),
    .A(net63),
    .Y(_0220_),
    .D(_0216_));
 sg13g2_nand2_1 _2914_ (.Y(_0221_),
    .A(net73),
    .B(_1334_));
 sg13g2_nand2_1 _2915_ (.Y(_0222_),
    .A(net73),
    .B(_1331_));
 sg13g2_mux2_1 _2916_ (.A0(_0221_),
    .A1(_0222_),
    .S(net28),
    .X(_0223_));
 sg13g2_mux2_1 _2917_ (.A0(_0221_),
    .A1(_0222_),
    .S(_0216_),
    .X(_0224_));
 sg13g2_nand4_1 _2918_ (.B(_0220_),
    .C(_0223_),
    .A(_0217_),
    .Y(_0225_),
    .D(_0224_));
 sg13g2_xnor2_1 _2919_ (.Y(_0226_),
    .A(_0208_),
    .B(_0225_));
 sg13g2_buf_1 _2920_ (.A(_1333_),
    .X(_0227_));
 sg13g2_nor2_1 _2921_ (.A(net59),
    .B(net110),
    .Y(_0228_));
 sg13g2_nor4_1 _2922_ (.A(net28),
    .B(_0093_),
    .C(_0098_),
    .D(_0109_),
    .Y(_0230_));
 sg13g2_nor2_1 _2923_ (.A(net62),
    .B(_0493_),
    .Y(_0231_));
 sg13g2_nand3_1 _2924_ (.B(_0214_),
    .C(_0215_),
    .A(net62),
    .Y(_0232_));
 sg13g2_buf_1 _2925_ (.A(_0232_),
    .X(_0233_));
 sg13g2_a21oi_1 _2926_ (.A1(_0091_),
    .A2(_0094_),
    .Y(_0234_),
    .B1(net60));
 sg13g2_and4_1 _2927_ (.A(net28),
    .B(_0233_),
    .C(_0234_),
    .D(_0109_),
    .X(_0235_));
 sg13g2_a22oi_1 _2928_ (.Y(_0236_),
    .B1(_0231_),
    .B2(_0235_),
    .A2(_0230_),
    .A1(_0228_));
 sg13g2_nand2_1 _2929_ (.Y(_0237_),
    .A(net106),
    .B(_1678_));
 sg13g2_nor2_1 _2930_ (.A(_0210_),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_nor2_1 _2931_ (.A(net59),
    .B(_1019_),
    .Y(_0239_));
 sg13g2_and2_1 _2932_ (.A(net104),
    .B(_1683_),
    .X(_0241_));
 sg13g2_o21ai_1 _2933_ (.B1(_0241_),
    .Y(_0242_),
    .A1(_0073_),
    .A2(_0088_));
 sg13g2_o21ai_1 _2934_ (.B1(_0242_),
    .Y(_0243_),
    .A1(_0239_),
    .A2(_0089_));
 sg13g2_and2_1 _2935_ (.A(net104),
    .B(_1678_),
    .X(_0244_));
 sg13g2_o21ai_1 _2936_ (.B1(_0244_),
    .Y(_0245_),
    .A1(_0213_),
    .A2(_0104_));
 sg13g2_o21ai_1 _2937_ (.B1(_0245_),
    .Y(_0246_),
    .A1(_0092_),
    .A2(_0214_));
 sg13g2_nor4_1 _2938_ (.A(_0062_),
    .B(_0243_),
    .C(_0246_),
    .D(_0109_),
    .Y(_0247_));
 sg13g2_nand2_1 _2939_ (.Y(_0248_),
    .A(_0951_),
    .B(_1683_));
 sg13g2_nor4_1 _2940_ (.A(_0062_),
    .B(_0093_),
    .C(_0098_),
    .D(_0248_),
    .Y(_0249_));
 sg13g2_a221oi_1 _2941_ (.B2(_0228_),
    .C1(_0249_),
    .B1(_0247_),
    .A1(_0099_),
    .Y(_0250_),
    .A2(_0238_));
 sg13g2_a221oi_1 _2942_ (.B2(_0106_),
    .C1(net28),
    .B1(_0105_),
    .A1(_0233_),
    .Y(_0252_),
    .A2(_0234_));
 sg13g2_nor2_1 _2943_ (.A(_0210_),
    .B(_0248_),
    .Y(_0253_));
 sg13g2_nand2_1 _2944_ (.Y(_0254_),
    .A(_0233_),
    .B(_0234_));
 sg13g2_nor4_1 _2945_ (.A(_0062_),
    .B(_0243_),
    .C(_0246_),
    .D(_0237_),
    .Y(_0255_));
 sg13g2_a221oi_1 _2946_ (.B2(_0254_),
    .C1(_0255_),
    .B1(_0253_),
    .A1(_0252_),
    .Y(_0256_),
    .A2(_0231_));
 sg13g2_mux2_1 _2947_ (.A0(_0237_),
    .A1(_0248_),
    .S(_0109_),
    .X(_0257_));
 sg13g2_nand4_1 _2948_ (.B(_0250_),
    .C(_0256_),
    .A(_0236_),
    .Y(_0258_),
    .D(_0257_));
 sg13g2_xnor2_1 _2949_ (.Y(_0259_),
    .A(_0226_),
    .B(_0258_));
 sg13g2_a21o_1 _2950_ (.A2(_0114_),
    .A1(net109),
    .B1(_0259_),
    .X(_0260_));
 sg13g2_xnor2_1 _2951_ (.Y(_0261_),
    .A(net122),
    .B(net48));
 sg13g2_nor2_1 _2952_ (.A(_0557_),
    .B(_0261_),
    .Y(_0263_));
 sg13g2_and3_1 _2953_ (.X(_0264_),
    .A(net109),
    .B(_0114_),
    .C(_0259_));
 sg13g2_a21oi_2 _2954_ (.B1(_0264_),
    .Y(_0265_),
    .A2(_0263_),
    .A1(_0260_));
 sg13g2_nand2_1 _2955_ (.Y(_0266_),
    .A(net63),
    .B(net106));
 sg13g2_a21oi_1 _2956_ (.A1(net59),
    .A2(_0209_),
    .Y(_0267_),
    .B1(_0216_));
 sg13g2_nor3_1 _2957_ (.A(net59),
    .B(net60),
    .C(_0209_),
    .Y(_0268_));
 sg13g2_o21ai_1 _2958_ (.B1(_0208_),
    .Y(_0269_),
    .A1(_0267_),
    .A2(_0268_));
 sg13g2_nand2_1 _2959_ (.Y(_0270_),
    .A(net59),
    .B(_0209_));
 sg13g2_nand2_1 _2960_ (.Y(_0271_),
    .A(net63),
    .B(net104));
 sg13g2_a21oi_1 _2961_ (.A1(_0089_),
    .A2(_0091_),
    .Y(_0272_),
    .B1(_0271_));
 sg13g2_nor3_1 _2962_ (.A(net59),
    .B(_0209_),
    .C(_0271_),
    .Y(_0274_));
 sg13g2_a221oi_1 _2963_ (.B2(_0272_),
    .C1(_0274_),
    .B1(_0270_),
    .A1(net63),
    .Y(_0275_),
    .A2(_0208_));
 sg13g2_nand2_1 _2964_ (.Y(_0276_),
    .A(net87),
    .B(net73));
 sg13g2_inv_1 _2965_ (.Y(_0277_),
    .A(_0276_));
 sg13g2_nand3_1 _2966_ (.B(_0275_),
    .C(_0277_),
    .A(_0269_),
    .Y(_0278_));
 sg13g2_buf_1 _2967_ (.A(_0278_),
    .X(_0279_));
 sg13g2_nand2_1 _2968_ (.Y(_0280_),
    .A(net80),
    .B(net73));
 sg13g2_a21o_1 _2969_ (.A2(_0275_),
    .A1(_0269_),
    .B1(_0280_),
    .X(_0281_));
 sg13g2_buf_1 _2970_ (.A(_0281_),
    .X(_0282_));
 sg13g2_o21ai_1 _2971_ (.B1(_0144_),
    .Y(_0283_),
    .A1(_0168_),
    .A2(_0170_));
 sg13g2_nand2b_1 _2972_ (.Y(_0285_),
    .B(_0158_),
    .A_N(_0283_));
 sg13g2_nor2_2 _2973_ (.A(_0168_),
    .B(_0170_),
    .Y(_0286_));
 sg13g2_a221oi_1 _2974_ (.B2(net76),
    .C1(net93),
    .B1(_0177_),
    .A1(net32),
    .Y(_0287_),
    .A2(_0286_));
 sg13g2_a21oi_1 _2975_ (.A1(_0177_),
    .A2(_0283_),
    .Y(_0288_),
    .B1(net76));
 sg13g2_buf_1 _2976_ (.A(_1144_),
    .X(_0289_));
 sg13g2_o21ai_1 _2977_ (.B1(net72),
    .Y(_0290_),
    .A1(_0287_),
    .A2(_0288_));
 sg13g2_buf_1 _2978_ (.A(_0290_),
    .X(_0291_));
 sg13g2_a21o_1 _2979_ (.A2(_1725_),
    .A1(net83),
    .B1(net122),
    .X(_0292_));
 sg13g2_a22oi_1 _2980_ (.Y(_0293_),
    .B1(_0292_),
    .B2(_1301_),
    .A2(net83),
    .A1(net122));
 sg13g2_nand2b_1 _2981_ (.Y(_0294_),
    .B(net114),
    .A_N(_0293_));
 sg13g2_nand2_1 _2982_ (.Y(_0296_),
    .A(net114),
    .B(net72));
 sg13g2_xor2_1 _2983_ (.B(_0296_),
    .A(_0294_),
    .X(_0297_));
 sg13g2_a21o_1 _2984_ (.A2(_0291_),
    .A1(_0285_),
    .B1(_0297_),
    .X(_0298_));
 sg13g2_buf_1 _2985_ (.A(_0298_),
    .X(_0299_));
 sg13g2_nand3_1 _2986_ (.B(_0291_),
    .C(_0297_),
    .A(_0285_),
    .Y(_0300_));
 sg13g2_buf_1 _2987_ (.A(_0300_),
    .X(_0301_));
 sg13g2_nand2_1 _2988_ (.Y(_0302_),
    .A(_0299_),
    .B(_0301_));
 sg13g2_nand2_1 _2989_ (.Y(_0303_),
    .A(net113),
    .B(net103));
 sg13g2_nor2_1 _2990_ (.A(net113),
    .B(_1753_),
    .Y(_0304_));
 sg13g2_nand2_1 _2991_ (.Y(_0305_),
    .A(net32),
    .B(_0304_));
 sg13g2_nand2_1 _2992_ (.Y(_0307_),
    .A(net72),
    .B(_0304_));
 sg13g2_nand4_1 _2993_ (.B(net75),
    .C(net72),
    .A(net74),
    .Y(_0308_),
    .D(net32));
 sg13g2_mux4_1 _2994_ (.S0(_0286_),
    .A0(_0303_),
    .A1(_0305_),
    .A2(_0307_),
    .A3(_0308_),
    .S1(net30),
    .X(_0309_));
 sg13g2_nor2_1 _2995_ (.A(_0143_),
    .B(_0307_),
    .Y(_0310_));
 sg13g2_or2_1 _2996_ (.X(_0311_),
    .B(net32),
    .A(_0303_));
 sg13g2_nand2_1 _2997_ (.Y(_0312_),
    .A(net75),
    .B(net78));
 sg13g2_a21oi_1 _2998_ (.A1(_0311_),
    .A2(_0312_),
    .Y(_0313_),
    .B1(net30));
 sg13g2_a21oi_1 _2999_ (.A1(net30),
    .A2(_0310_),
    .Y(_0314_),
    .B1(_0313_));
 sg13g2_nor2_1 _3000_ (.A(net76),
    .B(net89),
    .Y(_0315_));
 sg13g2_nand3_1 _3001_ (.B(_0314_),
    .C(_0315_),
    .A(_0309_),
    .Y(_0316_));
 sg13g2_a21oi_1 _3002_ (.A1(_0134_),
    .A2(_0139_),
    .Y(_0318_),
    .B1(_0316_));
 sg13g2_nor4_1 _3003_ (.A(net113),
    .B(net75),
    .C(net78),
    .D(net32),
    .Y(_0319_));
 sg13g2_nor2_1 _3004_ (.A(net76),
    .B(net75),
    .Y(_0320_));
 sg13g2_nor2b_1 _3005_ (.A(net32),
    .B_N(_0320_),
    .Y(_0321_));
 sg13g2_nor3_1 _3006_ (.A(_1129_),
    .B(net103),
    .C(net78),
    .Y(_0322_));
 sg13g2_nor2_1 _3007_ (.A(net113),
    .B(net103),
    .Y(_0323_));
 sg13g2_mux4_1 _3008_ (.S0(net30),
    .A0(_0319_),
    .A1(_0321_),
    .A2(_0322_),
    .A3(_0323_),
    .S1(_0286_),
    .X(_0324_));
 sg13g2_nand2_1 _3009_ (.Y(_0325_),
    .A(net32),
    .B(_0322_));
 sg13g2_nand3_1 _3010_ (.B(net30),
    .C(_0323_),
    .A(_0143_),
    .Y(_0326_));
 sg13g2_o21ai_1 _3011_ (.B1(_0326_),
    .Y(_0327_),
    .A1(net30),
    .A2(_0325_));
 sg13g2_nor3_1 _3012_ (.A(net75),
    .B(net72),
    .C(_0158_),
    .Y(_0329_));
 sg13g2_or2_1 _3013_ (.X(_0330_),
    .B(_0329_),
    .A(_0327_));
 sg13g2_nand2_1 _3014_ (.Y(_0331_),
    .A(net76),
    .B(net97));
 sg13g2_nor3_1 _3015_ (.A(_0324_),
    .B(_0330_),
    .C(_0331_),
    .Y(_0332_));
 sg13g2_and3_1 _3016_ (.X(_0333_),
    .A(_0134_),
    .B(_0139_),
    .C(_0332_));
 sg13g2_o21ai_1 _3017_ (.B1(_0315_),
    .Y(_0334_),
    .A1(_0324_),
    .A2(_0330_));
 sg13g2_a21o_1 _3018_ (.A2(_0314_),
    .A1(_0309_),
    .B1(_0331_),
    .X(_0335_));
 sg13g2_nand2_1 _3019_ (.Y(_0336_),
    .A(_0334_),
    .B(_0335_));
 sg13g2_nor3_1 _3020_ (.A(_0318_),
    .B(_0333_),
    .C(_0336_),
    .Y(_0337_));
 sg13g2_xor2_1 _3021_ (.B(_0337_),
    .A(_0302_),
    .X(_0338_));
 sg13g2_buf_2 _3022_ (.A(_0338_),
    .X(_0340_));
 sg13g2_inv_1 _3023_ (.Y(_0341_),
    .A(_0340_));
 sg13g2_a21oi_1 _3024_ (.A1(_0176_),
    .A2(_0180_),
    .Y(_0342_),
    .B1(_0181_));
 sg13g2_and3_1 _3025_ (.X(_0343_),
    .A(_0176_),
    .B(_0180_),
    .C(_0181_));
 sg13g2_o21ai_1 _3026_ (.B1(_0140_),
    .Y(_0344_),
    .A1(_0342_),
    .A2(_0343_));
 sg13g2_nand4_1 _3027_ (.B(_0139_),
    .C(_0182_),
    .A(_0134_),
    .Y(_0345_),
    .D(_0183_));
 sg13g2_buf_1 _3028_ (.A(_0878_),
    .X(_0346_));
 sg13g2_nor2_1 _3029_ (.A(net79),
    .B(net71),
    .Y(_0347_));
 sg13g2_and3_1 _3030_ (.X(_0348_),
    .A(net77),
    .B(_1769_),
    .C(_1771_));
 sg13g2_o21ai_1 _3031_ (.B1(_0059_),
    .Y(_0349_),
    .A1(_0347_),
    .A2(_0348_));
 sg13g2_a21oi_1 _3032_ (.A1(_1773_),
    .A2(_0347_),
    .Y(_0351_),
    .B1(net87));
 sg13g2_a22oi_1 _3033_ (.Y(_0352_),
    .B1(_0349_),
    .B2(_0351_),
    .A2(_0345_),
    .A1(_0344_));
 sg13g2_nand2_1 _3034_ (.Y(_0353_),
    .A(_0059_),
    .B(_0348_));
 sg13g2_o21ai_1 _3035_ (.B1(_0347_),
    .Y(_0354_),
    .A1(_1773_),
    .A2(_0059_));
 sg13g2_a21oi_1 _3036_ (.A1(_0353_),
    .A2(_0354_),
    .Y(_0355_),
    .B1(net80));
 sg13g2_nor2_1 _3037_ (.A(net75),
    .B(net71),
    .Y(_0356_));
 sg13g2_o21ai_1 _3038_ (.B1(_0356_),
    .Y(_0357_),
    .A1(_0352_),
    .A2(_0355_));
 sg13g2_buf_1 _3039_ (.A(net93),
    .X(_0358_));
 sg13g2_or4_1 _3040_ (.A(net58),
    .B(net71),
    .C(_0352_),
    .D(_0355_),
    .X(_0359_));
 sg13g2_nand3_1 _3041_ (.B(_0357_),
    .C(_0359_),
    .A(_0341_),
    .Y(_0360_));
 sg13g2_a21o_1 _3042_ (.A2(_0359_),
    .A1(_0357_),
    .B1(_0341_),
    .X(_0362_));
 sg13g2_and2_1 _3043_ (.A(_0360_),
    .B(_0362_),
    .X(_0363_));
 sg13g2_and4_1 _3044_ (.A(_0266_),
    .B(_0279_),
    .C(_0282_),
    .D(_0363_),
    .X(_0364_));
 sg13g2_a221oi_1 _3045_ (.B2(_0282_),
    .C1(_0363_),
    .B1(_0279_),
    .A1(net63),
    .Y(_0365_),
    .A2(net106));
 sg13g2_nor2_1 _3046_ (.A(net79),
    .B(net110),
    .Y(_0366_));
 sg13g2_nand2_1 _3047_ (.Y(_0367_),
    .A(_0360_),
    .B(_0362_));
 sg13g2_and4_1 _3048_ (.A(_0366_),
    .B(_0279_),
    .C(_0282_),
    .D(_0367_),
    .X(_0368_));
 sg13g2_nand3_1 _3049_ (.B(_0360_),
    .C(_0362_),
    .A(_0366_),
    .Y(_0369_));
 sg13g2_a21oi_1 _3050_ (.A1(_0279_),
    .A2(_0282_),
    .Y(_0370_),
    .B1(_0369_));
 sg13g2_nor4_1 _3051_ (.A(_0364_),
    .B(_0365_),
    .C(_0368_),
    .D(_0370_),
    .Y(_0371_));
 sg13g2_a21oi_1 _3052_ (.A1(_0214_),
    .A2(_0215_),
    .Y(_0373_),
    .B1(net62));
 sg13g2_o21ai_1 _3053_ (.B1(_0233_),
    .Y(_0374_),
    .A1(net28),
    .A2(_0373_));
 sg13g2_xnor2_1 _3054_ (.Y(_0375_),
    .A(net79),
    .B(_0374_));
 sg13g2_nor4_1 _3055_ (.A(net86),
    .B(_0062_),
    .C(_0093_),
    .D(_0098_),
    .Y(_0376_));
 sg13g2_nor4_1 _3056_ (.A(net86),
    .B(net28),
    .C(_0243_),
    .D(_0246_),
    .Y(_0377_));
 sg13g2_nor4_2 _3057_ (.A(_0235_),
    .B(_0376_),
    .C(_0252_),
    .Y(_0378_),
    .D(_0377_));
 sg13g2_nand2_1 _3058_ (.Y(_0379_),
    .A(_1461_),
    .B(_0109_));
 sg13g2_nand2_1 _3059_ (.Y(_0380_),
    .A(net106),
    .B(_0208_));
 sg13g2_a221oi_1 _3060_ (.B2(_0379_),
    .C1(_0380_),
    .B1(_0378_),
    .A1(net73),
    .Y(_0381_),
    .A2(_0375_));
 sg13g2_and2_1 _3061_ (.A(_0217_),
    .B(_0220_),
    .X(_0382_));
 sg13g2_and2_1 _3062_ (.A(_0223_),
    .B(_0224_),
    .X(_0384_));
 sg13g2_or2_1 _3063_ (.X(_0385_),
    .B(_0208_),
    .A(net110));
 sg13g2_a221oi_1 _3064_ (.B2(_0379_),
    .C1(_0385_),
    .B1(_0378_),
    .A1(_0382_),
    .Y(_0386_),
    .A2(_0384_));
 sg13g2_nand2_1 _3065_ (.Y(_0387_),
    .A(_1355_),
    .B(net106));
 sg13g2_a21oi_1 _3066_ (.A1(_0378_),
    .A2(_0379_),
    .Y(_0388_),
    .B1(_0387_));
 sg13g2_and2_1 _3067_ (.A(_0208_),
    .B(_0228_),
    .X(_0389_));
 sg13g2_nor2_1 _3068_ (.A(_0208_),
    .B(_0387_),
    .Y(_0390_));
 sg13g2_mux2_1 _3069_ (.A0(_0389_),
    .A1(_0390_),
    .S(_0225_),
    .X(_0391_));
 sg13g2_nor4_2 _3070_ (.A(_0381_),
    .B(_0386_),
    .C(_0388_),
    .Y(_0392_),
    .D(_0391_));
 sg13g2_xor2_1 _3071_ (.B(_0392_),
    .A(_0371_),
    .X(_0393_));
 sg13g2_xor2_1 _3072_ (.B(net62),
    .A(_1438_),
    .X(_0395_));
 sg13g2_nand2_1 _3073_ (.Y(_0396_),
    .A(net109),
    .B(_0395_));
 sg13g2_o21ai_1 _3074_ (.B1(_0396_),
    .Y(_0397_),
    .A1(_0265_),
    .A2(_0393_));
 sg13g2_nand2_1 _3075_ (.Y(_0398_),
    .A(_0265_),
    .B(_0393_));
 sg13g2_nand2_1 _3076_ (.Y(_0399_),
    .A(_0397_),
    .B(_0398_));
 sg13g2_nor2_1 _3077_ (.A(_0368_),
    .B(_0370_),
    .Y(_0400_));
 sg13g2_nand3_1 _3078_ (.B(_0282_),
    .C(_0367_),
    .A(_0279_),
    .Y(_0401_));
 sg13g2_a21o_1 _3079_ (.A2(_0282_),
    .A1(_0279_),
    .B1(_0367_),
    .X(_0402_));
 sg13g2_a21o_1 _3080_ (.A2(_0402_),
    .A1(_0401_),
    .B1(_0392_),
    .X(_0403_));
 sg13g2_or2_1 _3081_ (.X(_0404_),
    .B(_0392_),
    .A(_0266_));
 sg13g2_nand3_1 _3082_ (.B(_0403_),
    .C(_0404_),
    .A(_0400_),
    .Y(_0406_));
 sg13g2_buf_1 _3083_ (.A(_0171_),
    .X(_0407_));
 sg13g2_buf_1 _3084_ (.A(_1774_),
    .X(_0408_));
 sg13g2_nor2_1 _3085_ (.A(_0198_),
    .B(_0199_),
    .Y(_0409_));
 sg13g2_o21ai_1 _3086_ (.B1(_0409_),
    .Y(_0410_),
    .A1(_0188_),
    .A2(_0192_));
 sg13g2_nand4_1 _3087_ (.B(_0184_),
    .C(_0186_),
    .A(net56),
    .Y(_0411_),
    .D(_0410_));
 sg13g2_nor4_1 _3088_ (.A(net57),
    .B(net71),
    .C(_0340_),
    .D(_0411_),
    .Y(_0412_));
 sg13g2_nor2_1 _3089_ (.A(net58),
    .B(net71),
    .Y(_0413_));
 sg13g2_nand3_1 _3090_ (.B(_0345_),
    .C(_0413_),
    .A(_0344_),
    .Y(_0414_));
 sg13g2_mux2_1 _3091_ (.A0(_0414_),
    .A1(net56),
    .S(_0340_),
    .X(_0415_));
 sg13g2_a21oi_1 _3092_ (.A1(_0184_),
    .A2(_0186_),
    .Y(_0417_),
    .B1(_0171_));
 sg13g2_a221oi_1 _3093_ (.B2(_0354_),
    .C1(net58),
    .B1(_0353_),
    .A1(_0344_),
    .Y(_0418_),
    .A2(_0345_));
 sg13g2_o21ai_1 _3094_ (.B1(_0340_),
    .Y(_0419_),
    .A1(_0417_),
    .A2(_0418_));
 sg13g2_nand3b_1 _3095_ (.B(_0415_),
    .C(_0419_),
    .Y(_0420_),
    .A_N(_0412_));
 sg13g2_a21oi_1 _3096_ (.A1(net56),
    .A2(_0410_),
    .Y(_0421_),
    .B1(net87));
 sg13g2_mux2_1 _3097_ (.A0(_0413_),
    .A1(net58),
    .S(_0340_),
    .X(_0422_));
 sg13g2_a21o_1 _3098_ (.A2(_0422_),
    .A1(_0421_),
    .B1(net60),
    .X(_0423_));
 sg13g2_a221oi_1 _3099_ (.B2(net80),
    .C1(_0423_),
    .B1(_0420_),
    .A1(_0269_),
    .Y(_0424_),
    .A2(_0275_));
 sg13g2_a21oi_1 _3100_ (.A1(_0277_),
    .A2(_0367_),
    .Y(_0425_),
    .B1(_0424_));
 sg13g2_or2_1 _3101_ (.X(_0426_),
    .B(_0411_),
    .A(_0340_));
 sg13g2_buf_1 _3102_ (.A(_0426_),
    .X(_0428_));
 sg13g2_nand2_1 _3103_ (.Y(_0429_),
    .A(net57),
    .B(net73));
 sg13g2_nand2_1 _3104_ (.Y(_0430_),
    .A(net56),
    .B(_0410_));
 sg13g2_a221oi_1 _3105_ (.B2(_0187_),
    .C1(_1617_),
    .B1(_0430_),
    .A1(net58),
    .Y(_0431_),
    .A2(_0340_));
 sg13g2_a21oi_1 _3106_ (.A1(_0340_),
    .A2(_0411_),
    .Y(_0432_),
    .B1(net58));
 sg13g2_o21ai_1 _3107_ (.B1(net56),
    .Y(_0433_),
    .A1(_0431_),
    .A2(_0432_));
 sg13g2_buf_1 _3108_ (.A(_0433_),
    .X(_0434_));
 sg13g2_nand2_1 _3109_ (.Y(_0435_),
    .A(net74),
    .B(net56));
 sg13g2_nand4_1 _3110_ (.B(_0139_),
    .C(_0176_),
    .A(_0134_),
    .Y(_0436_),
    .D(_0180_));
 sg13g2_nand3_1 _3111_ (.B(_0301_),
    .C(_0436_),
    .A(_0299_),
    .Y(_0437_));
 sg13g2_nand2_1 _3112_ (.Y(_0439_),
    .A(_0176_),
    .B(_0180_));
 sg13g2_a21oi_1 _3113_ (.A1(_0140_),
    .A2(_0439_),
    .Y(_0440_),
    .B1(net58));
 sg13g2_o21ai_1 _3114_ (.B1(_0315_),
    .Y(_0441_),
    .A1(_0437_),
    .A2(_0440_));
 sg13g2_buf_1 _3115_ (.A(_0441_),
    .X(_0442_));
 sg13g2_a21oi_1 _3116_ (.A1(_0299_),
    .A2(_0301_),
    .Y(_0443_),
    .B1(net89));
 sg13g2_a21oi_1 _3117_ (.A1(_0299_),
    .A2(_0301_),
    .Y(_0444_),
    .B1(_0436_));
 sg13g2_a21oi_1 _3118_ (.A1(_0440_),
    .A2(_0443_),
    .Y(_0445_),
    .B1(_0444_));
 sg13g2_buf_1 _3119_ (.A(_0445_),
    .X(_0446_));
 sg13g2_nand2_1 _3120_ (.Y(_0447_),
    .A(net84),
    .B(net89));
 sg13g2_nand2_1 _3121_ (.Y(_0448_),
    .A(net84),
    .B(net97));
 sg13g2_nand3_1 _3122_ (.B(_0291_),
    .C(_0294_),
    .A(_0285_),
    .Y(_0450_));
 sg13g2_xnor2_1 _3123_ (.Y(_0451_),
    .A(net72),
    .B(_0196_));
 sg13g2_a22oi_1 _3124_ (.Y(_0452_),
    .B1(_0451_),
    .B2(net122),
    .A2(_0450_),
    .A1(net72));
 sg13g2_buf_1 _3125_ (.A(_0452_),
    .X(_0453_));
 sg13g2_mux2_1 _3126_ (.A0(_0447_),
    .A1(_0448_),
    .S(_0453_),
    .X(_0454_));
 sg13g2_buf_1 _3127_ (.A(_0454_),
    .X(_0455_));
 sg13g2_and4_1 _3128_ (.A(_0435_),
    .B(_0442_),
    .C(_0446_),
    .D(_0455_),
    .X(_0456_));
 sg13g2_a221oi_1 _3129_ (.B2(_0446_),
    .C1(_0455_),
    .B1(_0442_),
    .A1(net74),
    .Y(_0457_),
    .A2(net56));
 sg13g2_xnor2_1 _3130_ (.Y(_0458_),
    .A(net97),
    .B(_0453_));
 sg13g2_a221oi_1 _3131_ (.B2(net84),
    .C1(_0435_),
    .B1(_0458_),
    .A1(_0442_),
    .Y(_0459_),
    .A2(_0446_));
 sg13g2_inv_1 _3132_ (.Y(_0461_),
    .A(_0435_));
 sg13g2_nor2_1 _3133_ (.A(net108),
    .B(net97),
    .Y(_0462_));
 sg13g2_nor2_1 _3134_ (.A(net108),
    .B(net89),
    .Y(_0463_));
 sg13g2_mux2_1 _3135_ (.A0(_0462_),
    .A1(_0463_),
    .S(_0453_),
    .X(_0464_));
 sg13g2_and4_1 _3136_ (.A(_0461_),
    .B(_0442_),
    .C(_0446_),
    .D(_0464_),
    .X(_0465_));
 sg13g2_nor4_2 _3137_ (.A(_0456_),
    .B(_0457_),
    .C(_0459_),
    .Y(_0466_),
    .D(_0465_));
 sg13g2_and4_1 _3138_ (.A(net26),
    .B(_0429_),
    .C(net24),
    .D(_0466_),
    .X(_0467_));
 sg13g2_a221oi_1 _3139_ (.B2(net24),
    .C1(_0466_),
    .B1(net26),
    .A1(net57),
    .Y(_0468_),
    .A2(net73));
 sg13g2_a21o_1 _3140_ (.A2(_0446_),
    .A1(_0442_),
    .B1(_0455_),
    .X(_0469_));
 sg13g2_buf_1 _3141_ (.A(_0469_),
    .X(_0470_));
 sg13g2_nand3_1 _3142_ (.B(_0446_),
    .C(_0455_),
    .A(_0442_),
    .Y(_0472_));
 sg13g2_buf_1 _3143_ (.A(_0472_),
    .X(_0473_));
 sg13g2_a21o_1 _3144_ (.A2(_0473_),
    .A1(_0470_),
    .B1(_0435_),
    .X(_0474_));
 sg13g2_nand3_1 _3145_ (.B(_0470_),
    .C(_0473_),
    .A(_0435_),
    .Y(_0475_));
 sg13g2_a221oi_1 _3146_ (.B2(_0475_),
    .C1(_0429_),
    .B1(_0474_),
    .A1(net26),
    .Y(_0476_),
    .A2(_0434_));
 sg13g2_nor2_1 _3147_ (.A(_0358_),
    .B(net60),
    .Y(_0477_));
 sg13g2_or4_1 _3148_ (.A(_0456_),
    .B(_0457_),
    .C(_0459_),
    .D(_0465_),
    .X(_0478_));
 sg13g2_and4_1 _3149_ (.A(net26),
    .B(_0477_),
    .C(net24),
    .D(_0478_),
    .X(_0479_));
 sg13g2_nor4_1 _3150_ (.A(_0467_),
    .B(_0468_),
    .C(_0476_),
    .D(_0479_),
    .Y(_0480_));
 sg13g2_xor2_1 _3151_ (.B(_0480_),
    .A(_0425_),
    .X(_0481_));
 sg13g2_buf_1 _3152_ (.A(net106),
    .X(_0483_));
 sg13g2_nand2_1 _3153_ (.Y(_0484_),
    .A(net87),
    .B(net70));
 sg13g2_xor2_1 _3154_ (.B(_0484_),
    .A(_0481_),
    .X(_0485_));
 sg13g2_xnor2_1 _3155_ (.Y(_0486_),
    .A(_0406_),
    .B(_0485_));
 sg13g2_xor2_1 _3156_ (.B(net63),
    .A(net122),
    .X(_0487_));
 sg13g2_nand2_1 _3157_ (.Y(_0488_),
    .A(_0601_),
    .B(_0487_));
 sg13g2_xnor2_1 _3158_ (.Y(_0489_),
    .A(_0486_),
    .B(_0488_));
 sg13g2_xnor2_1 _3159_ (.Y(_0490_),
    .A(_0399_),
    .B(_0489_));
 sg13g2_nand2_1 _3160_ (.Y(_0491_),
    .A(_1573_),
    .B(_0490_));
 sg13g2_o21ai_1 _3161_ (.B1(_0491_),
    .Y(_0492_),
    .A1(net121),
    .A2(_1585_));
 sg13g2_mux2_1 _3162_ (.A0(\muldiv.regR[10] ),
    .A1(_0492_),
    .S(net127),
    .X(_0005_));
 sg13g2_buf_1 _3163_ (.A(_1599_),
    .X(_0494_));
 sg13g2_and2_1 _3164_ (.A(_0141_),
    .B(net29),
    .X(_0495_));
 sg13g2_buf_1 _3165_ (.A(_0495_),
    .X(_0496_));
 sg13g2_a21oi_1 _3166_ (.A1(_1467_),
    .A2(_1583_),
    .Y(_0497_),
    .B1(_1581_));
 sg13g2_xnor2_1 _3167_ (.Y(_0498_),
    .A(_0496_),
    .B(_0497_));
 sg13g2_nand2_1 _3168_ (.Y(_0499_),
    .A(_0470_),
    .B(_0473_));
 sg13g2_nand3_1 _3169_ (.B(_0434_),
    .C(_0499_),
    .A(_0428_),
    .Y(_0500_));
 sg13g2_nand2_1 _3170_ (.Y(_0501_),
    .A(net74),
    .B(_0500_));
 sg13g2_a21oi_1 _3171_ (.A1(_0428_),
    .A2(net24),
    .Y(_0502_),
    .B1(_0499_));
 sg13g2_nand3_1 _3172_ (.B(net83),
    .C(_1725_),
    .A(net82),
    .Y(_0504_));
 sg13g2_nand3_1 _3173_ (.B(_0291_),
    .C(_0504_),
    .A(_0285_),
    .Y(_0505_));
 sg13g2_nor2_1 _3174_ (.A(net120),
    .B(net92),
    .Y(_0506_));
 sg13g2_a21oi_1 _3175_ (.A1(net72),
    .A2(_0505_),
    .Y(_0507_),
    .B1(_0506_));
 sg13g2_nand3_1 _3176_ (.B(_0446_),
    .C(_0507_),
    .A(_0442_),
    .Y(_0508_));
 sg13g2_o21ai_1 _3177_ (.B1(net84),
    .Y(_0509_),
    .A1(_1670_),
    .A2(_0506_));
 sg13g2_inv_1 _3178_ (.Y(_0510_),
    .A(_0509_));
 sg13g2_nand2_1 _3179_ (.Y(_0511_),
    .A(_0508_),
    .B(_0510_));
 sg13g2_o21ai_1 _3180_ (.B1(net84),
    .Y(_0512_),
    .A1(_0346_),
    .A2(_0511_));
 sg13g2_nor2b_1 _3181_ (.A(_0502_),
    .B_N(_0512_),
    .Y(_0513_));
 sg13g2_a21oi_1 _3182_ (.A1(_0508_),
    .A2(_0510_),
    .Y(_0515_),
    .B1(net108));
 sg13g2_a21o_1 _3183_ (.A2(_0500_),
    .A1(net74),
    .B1(_0502_),
    .X(_0516_));
 sg13g2_nand2_1 _3184_ (.Y(_0517_),
    .A(_0346_),
    .B(_0511_));
 sg13g2_inv_1 _3185_ (.Y(_0518_),
    .A(_0517_));
 sg13g2_a221oi_1 _3186_ (.B2(_0516_),
    .C1(_0518_),
    .B1(_0515_),
    .A1(_0501_),
    .Y(_0519_),
    .A2(_0513_));
 sg13g2_buf_2 _3187_ (.A(_0519_),
    .X(_0520_));
 sg13g2_nor2_1 _3188_ (.A(net76),
    .B(net60),
    .Y(_0521_));
 sg13g2_nor2_1 _3189_ (.A(_0178_),
    .B(net60),
    .Y(_0522_));
 sg13g2_a21oi_1 _3190_ (.A1(net26),
    .A2(net24),
    .Y(_0523_),
    .B1(_0466_));
 sg13g2_and3_1 _3191_ (.X(_0524_),
    .A(net26),
    .B(net24),
    .C(_0466_));
 sg13g2_nor2_1 _3192_ (.A(_0523_),
    .B(_0524_),
    .Y(_0526_));
 sg13g2_a21oi_1 _3193_ (.A1(_0277_),
    .A2(_0367_),
    .Y(_0527_),
    .B1(net57));
 sg13g2_inv_1 _3194_ (.Y(_0528_),
    .A(_0424_));
 sg13g2_nor3_1 _3195_ (.A(net57),
    .B(_0523_),
    .C(_0524_),
    .Y(_0529_));
 sg13g2_a221oi_1 _3196_ (.B2(_0528_),
    .C1(_0529_),
    .B1(_0527_),
    .A1(_0425_),
    .Y(_0530_),
    .A2(_0526_));
 sg13g2_buf_2 _3197_ (.A(_0530_),
    .X(_0531_));
 sg13g2_mux2_1 _3198_ (.A0(_0521_),
    .A1(_0522_),
    .S(_0531_),
    .X(_0532_));
 sg13g2_buf_1 _3199_ (.A(_0532_),
    .X(_0533_));
 sg13g2_xor2_1 _3200_ (.B(_0533_),
    .A(_0520_),
    .X(_0534_));
 sg13g2_nand2_1 _3201_ (.Y(_0535_),
    .A(_0358_),
    .B(net70));
 sg13g2_nand2_1 _3202_ (.Y(_0537_),
    .A(net57),
    .B(_0483_));
 sg13g2_nand2b_1 _3203_ (.Y(_0538_),
    .B(_1617_),
    .A_N(_0481_));
 sg13g2_and2_1 _3204_ (.A(_1266_),
    .B(_0481_),
    .X(_0539_));
 sg13g2_a21oi_1 _3205_ (.A1(_0406_),
    .A2(_0538_),
    .Y(_0540_),
    .B1(_0539_));
 sg13g2_mux2_1 _3206_ (.A0(_0535_),
    .A1(_0537_),
    .S(_0540_),
    .X(_0541_));
 sg13g2_xnor2_1 _3207_ (.Y(_0542_),
    .A(_0534_),
    .B(_0541_));
 sg13g2_xor2_1 _3208_ (.B(_1266_),
    .A(net119),
    .X(_0543_));
 sg13g2_nand2_1 _3209_ (.Y(_0544_),
    .A(_0601_),
    .B(_0543_));
 sg13g2_inv_1 _3210_ (.Y(_0545_),
    .A(_0544_));
 sg13g2_nand3_1 _3211_ (.B(_0398_),
    .C(_0486_),
    .A(_0397_),
    .Y(_0546_));
 sg13g2_a21oi_1 _3212_ (.A1(_0397_),
    .A2(_0398_),
    .Y(_0548_),
    .B1(_0486_));
 sg13g2_a21oi_1 _3213_ (.A1(_0488_),
    .A2(_0546_),
    .Y(_0549_),
    .B1(_0548_));
 sg13g2_xnor2_1 _3214_ (.Y(_0550_),
    .A(_0545_),
    .B(_0549_));
 sg13g2_xnor2_1 _3215_ (.Y(_0551_),
    .A(_0542_),
    .B(_0550_));
 sg13g2_nor2_1 _3216_ (.A(_1561_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_a21o_1 _3217_ (.A2(_0498_),
    .A1(net126),
    .B1(_0552_),
    .X(_0553_));
 sg13g2_buf_1 _3218_ (.A(net131),
    .X(_0554_));
 sg13g2_nor2_1 _3219_ (.A(net125),
    .B(\muldiv.regR[11] ),
    .Y(_0555_));
 sg13g2_a21oi_1 _3220_ (.A1(net127),
    .A2(_0553_),
    .Y(_0006_),
    .B1(_0555_));
 sg13g2_nor2_1 _3221_ (.A(_0496_),
    .B(_1407_),
    .Y(_0556_));
 sg13g2_a21oi_1 _3222_ (.A1(_1583_),
    .A2(_0556_),
    .Y(_0558_),
    .B1(_1581_));
 sg13g2_xnor2_1 _3223_ (.Y(_0559_),
    .A(_1201_),
    .B(_0558_));
 sg13g2_nand2_1 _3224_ (.Y(_0560_),
    .A(_0488_),
    .B(_0544_));
 sg13g2_inv_1 _3225_ (.Y(_0561_),
    .A(_0560_));
 sg13g2_nor2_1 _3226_ (.A(_0486_),
    .B(_0560_),
    .Y(_0562_));
 sg13g2_a221oi_1 _3227_ (.B2(_0399_),
    .C1(_0562_),
    .B1(_0561_),
    .A1(_0544_),
    .Y(_0563_),
    .A2(_0548_));
 sg13g2_a22oi_1 _3228_ (.Y(_0564_),
    .B1(_0563_),
    .B2(_0542_),
    .A2(_0549_),
    .A1(_0545_));
 sg13g2_xor2_1 _3229_ (.B(net57),
    .A(net119),
    .X(_0565_));
 sg13g2_nand2_1 _3230_ (.Y(_0566_),
    .A(net81),
    .B(_0565_));
 sg13g2_nand2_1 _3231_ (.Y(_0567_),
    .A(net74),
    .B(net70));
 sg13g2_o21ai_1 _3232_ (.B1(_0521_),
    .Y(_0569_),
    .A1(_0520_),
    .A2(_0531_));
 sg13g2_nand2b_1 _3233_ (.Y(_0570_),
    .B(_0512_),
    .A_N(_0502_));
 sg13g2_nand3_1 _3234_ (.B(_0502_),
    .C(_0511_),
    .A(net84),
    .Y(_0571_));
 sg13g2_and4_1 _3235_ (.A(_0219_),
    .B(_0570_),
    .C(_0517_),
    .D(_0571_),
    .X(_0572_));
 sg13g2_nand2_1 _3236_ (.Y(_0573_),
    .A(_1431_),
    .B(_0095_));
 sg13g2_nand2_1 _3237_ (.Y(_0574_),
    .A(_1431_),
    .B(_0219_));
 sg13g2_nand2_1 _3238_ (.Y(_0575_),
    .A(_0408_),
    .B(_0972_));
 sg13g2_nand3_1 _3239_ (.B(_1003_),
    .C(_0575_),
    .A(_1438_),
    .Y(_0576_));
 sg13g2_a22oi_1 _3240_ (.Y(_0577_),
    .B1(_0508_),
    .B2(_0510_),
    .A2(_0473_),
    .A1(_0470_));
 sg13g2_nand4_1 _3241_ (.B(net26),
    .C(net24),
    .A(_0576_),
    .Y(_0578_),
    .D(_0577_));
 sg13g2_and2_1 _3242_ (.A(net76),
    .B(_0576_),
    .X(_0580_));
 sg13g2_nand4_1 _3243_ (.B(net24),
    .C(_0511_),
    .A(net26),
    .Y(_0581_),
    .D(_0580_));
 sg13g2_a22oi_1 _3244_ (.Y(_0582_),
    .B1(_0577_),
    .B2(_0580_),
    .A2(_0576_),
    .A1(net71));
 sg13g2_nand3_1 _3245_ (.B(_0581_),
    .C(_0582_),
    .A(_0578_),
    .Y(_0583_));
 sg13g2_mux2_1 _3246_ (.A0(_0573_),
    .A1(_0574_),
    .S(_0583_),
    .X(_0584_));
 sg13g2_a21oi_1 _3247_ (.A1(_0531_),
    .A2(_0572_),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_and2_1 _3248_ (.A(_0521_),
    .B(_0584_),
    .X(_0586_));
 sg13g2_or2_1 _3249_ (.X(_0587_),
    .B(_0531_),
    .A(_0520_));
 sg13g2_and3_1 _3250_ (.X(_0588_),
    .A(_0531_),
    .B(_0584_),
    .C(_0572_));
 sg13g2_a221oi_1 _3251_ (.B2(_0587_),
    .C1(_0588_),
    .B1(_0586_),
    .A1(_0569_),
    .Y(_0589_),
    .A2(_0585_));
 sg13g2_xor2_1 _3252_ (.B(_0589_),
    .A(_0567_),
    .X(_0591_));
 sg13g2_or2_1 _3253_ (.X(_0592_),
    .B(_0591_),
    .A(_0566_));
 sg13g2_nand2b_1 _3254_ (.Y(_0593_),
    .B(_0591_),
    .A_N(_0566_));
 sg13g2_nor2_1 _3255_ (.A(_0407_),
    .B(_0520_),
    .Y(_0594_));
 sg13g2_and2_1 _3256_ (.A(net58),
    .B(_0520_),
    .X(_0595_));
 sg13g2_mux2_1 _3257_ (.A0(_0594_),
    .A1(_0595_),
    .S(_0533_),
    .X(_0596_));
 sg13g2_nand2_1 _3258_ (.Y(_0597_),
    .A(_0407_),
    .B(_0520_));
 sg13g2_nand2b_1 _3259_ (.Y(_0598_),
    .B(net57),
    .A_N(_0520_));
 sg13g2_mux2_1 _3260_ (.A0(_0597_),
    .A1(_0598_),
    .S(_0533_),
    .X(_0599_));
 sg13g2_o21ai_1 _3261_ (.B1(_0599_),
    .Y(_0600_),
    .A1(_0540_),
    .A2(_0596_));
 sg13g2_nand2_1 _3262_ (.Y(_0602_),
    .A(net70),
    .B(_0600_));
 sg13g2_mux2_1 _3263_ (.A0(_0592_),
    .A1(_0593_),
    .S(_0602_),
    .X(_0603_));
 sg13g2_a221oi_1 _3264_ (.B2(net70),
    .C1(_0591_),
    .B1(_0600_),
    .A1(net81),
    .Y(_0604_),
    .A2(_0565_));
 sg13g2_nand4_1 _3265_ (.B(_0566_),
    .C(_0600_),
    .A(net70),
    .Y(_0605_),
    .D(_0591_));
 sg13g2_nor2b_1 _3266_ (.A(_0604_),
    .B_N(_0605_),
    .Y(_0606_));
 sg13g2_and2_1 _3267_ (.A(_0603_),
    .B(_0606_),
    .X(_0607_));
 sg13g2_xnor2_1 _3268_ (.Y(_0608_),
    .A(_0564_),
    .B(_0607_));
 sg13g2_nand2_1 _3269_ (.Y(_0609_),
    .A(_1573_),
    .B(_0608_));
 sg13g2_o21ai_1 _3270_ (.B1(_0609_),
    .Y(_0610_),
    .A1(_1574_),
    .A2(_0559_));
 sg13g2_mux2_1 _3271_ (.A0(\muldiv.regR[12] ),
    .A1(_0610_),
    .S(net127),
    .X(_0007_));
 sg13g2_nand2_1 _3272_ (.Y(_0612_),
    .A(_0967_),
    .B(_1104_));
 sg13g2_nor3_1 _3273_ (.A(_1201_),
    .B(_0496_),
    .C(_1407_),
    .Y(_0613_));
 sg13g2_and4_1 _3274_ (.A(_1515_),
    .B(_1542_),
    .C(_1557_),
    .D(_0613_),
    .X(_0614_));
 sg13g2_buf_8 _3275_ (.A(_0614_),
    .X(_0615_));
 sg13g2_nor2_1 _3276_ (.A(_1581_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_xnor2_1 _3277_ (.Y(_0617_),
    .A(_0612_),
    .B(_0616_));
 sg13g2_and4_1 _3278_ (.A(_0570_),
    .B(_0517_),
    .C(_0531_),
    .D(_0571_),
    .X(_0618_));
 sg13g2_o21ai_1 _3279_ (.B1(_0587_),
    .Y(_0619_),
    .A1(_0178_),
    .A2(_0618_));
 sg13g2_nor2_1 _3280_ (.A(_0583_),
    .B(_0574_),
    .Y(_0620_));
 sg13g2_a21oi_1 _3281_ (.A1(net119),
    .A2(_0654_),
    .Y(_0621_),
    .B1(_0620_));
 sg13g2_o21ai_1 _3282_ (.B1(_0621_),
    .Y(_0623_),
    .A1(_0095_),
    .A2(_0619_));
 sg13g2_and2_1 _3283_ (.A(_0599_),
    .B(_0589_),
    .X(_0624_));
 sg13g2_or2_1 _3284_ (.X(_0625_),
    .B(_0596_),
    .A(_0540_));
 sg13g2_a22oi_1 _3285_ (.Y(_0626_),
    .B1(_0624_),
    .B2(_0625_),
    .A2(_0589_),
    .A1(_0567_));
 sg13g2_buf_1 _3286_ (.A(_0626_),
    .X(_0627_));
 sg13g2_and2_1 _3287_ (.A(_0160_),
    .B(_0599_),
    .X(_0628_));
 sg13g2_a22oi_1 _3288_ (.Y(_0629_),
    .B1(_0625_),
    .B2(_0628_),
    .A2(net110),
    .A1(_0160_));
 sg13g2_buf_1 _3289_ (.A(_0629_),
    .X(_0630_));
 sg13g2_and4_1 _3290_ (.A(net61),
    .B(_0623_),
    .C(_0627_),
    .D(_0630_),
    .X(_0631_));
 sg13g2_nand3b_1 _3291_ (.B(net70),
    .C(net61),
    .Y(_0632_),
    .A_N(_0623_));
 sg13g2_a21oi_1 _3292_ (.A1(_0627_),
    .A2(_0630_),
    .Y(_0634_),
    .B1(_0632_));
 sg13g2_and3_1 _3293_ (.X(_0635_),
    .A(net61),
    .B(_0493_),
    .C(_0623_));
 sg13g2_and4_1 _3294_ (.A(net108),
    .B(net70),
    .C(_0627_),
    .D(_0630_),
    .X(_0636_));
 sg13g2_nor4_2 _3295_ (.A(_0631_),
    .B(_0634_),
    .C(_0635_),
    .Y(_0637_),
    .D(_0636_));
 sg13g2_xor2_1 _3296_ (.B(net74),
    .A(net119),
    .X(_0638_));
 sg13g2_and2_1 _3297_ (.A(net81),
    .B(_0638_),
    .X(_0639_));
 sg13g2_nand2b_1 _3298_ (.Y(_0640_),
    .B(_0605_),
    .A_N(_0604_));
 sg13g2_o21ai_1 _3299_ (.B1(_0603_),
    .Y(_0641_),
    .A1(_0564_),
    .A2(_0640_));
 sg13g2_nor2_1 _3300_ (.A(_0639_),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_nand2_1 _3301_ (.Y(_0643_),
    .A(_0639_),
    .B(_0641_));
 sg13g2_nand2b_1 _3302_ (.Y(_0645_),
    .B(_0643_),
    .A_N(_0642_));
 sg13g2_xnor2_1 _3303_ (.Y(_0646_),
    .A(_0637_),
    .B(_0645_));
 sg13g2_nor2_1 _3304_ (.A(net128),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_a21o_1 _3305_ (.A2(_0617_),
    .A1(net126),
    .B1(_0647_),
    .X(_0648_));
 sg13g2_mux2_1 _3306_ (.A0(\muldiv.regR[13] ),
    .A1(_0648_),
    .S(net127),
    .X(_0008_));
 sg13g2_a21oi_1 _3307_ (.A1(_0637_),
    .A2(_0643_),
    .Y(_0649_),
    .B1(_0642_));
 sg13g2_a221oi_1 _3308_ (.B2(_0630_),
    .C1(_0623_),
    .B1(_0627_),
    .A1(net119),
    .Y(_0650_),
    .A2(_0547_));
 sg13g2_nor2_1 _3309_ (.A(net120),
    .B(_0973_),
    .Y(_0651_));
 sg13g2_o21ai_1 _3310_ (.B1(net61),
    .Y(_0652_),
    .A1(_0483_),
    .A2(_0651_));
 sg13g2_nor2_1 _3311_ (.A(_0650_),
    .B(_0652_),
    .Y(_0653_));
 sg13g2_nor2_1 _3312_ (.A(net120),
    .B(_1578_),
    .Y(_0655_));
 sg13g2_o21ai_1 _3313_ (.B1(net81),
    .Y(_0656_),
    .A1(_1128_),
    .A2(_0655_));
 sg13g2_xnor2_1 _3314_ (.Y(_0657_),
    .A(_0653_),
    .B(_0656_));
 sg13g2_xnor2_1 _3315_ (.Y(_0658_),
    .A(_0649_),
    .B(_0657_));
 sg13g2_nand2_1 _3316_ (.Y(_0659_),
    .A(net121),
    .B(_0658_));
 sg13g2_nand2_1 _3317_ (.Y(_0660_),
    .A(net125),
    .B(_0659_));
 sg13g2_a21oi_1 _3318_ (.A1(_0612_),
    .A2(_0615_),
    .Y(_0661_),
    .B1(_1581_));
 sg13g2_a21oi_1 _3319_ (.A1(net48),
    .A2(_0975_),
    .Y(_0662_),
    .B1(_0739_));
 sg13g2_nand2_1 _3320_ (.Y(_0663_),
    .A(net55),
    .B(_0662_));
 sg13g2_o21ai_1 _3321_ (.B1(_0663_),
    .Y(_0664_),
    .A1(_1577_),
    .A2(_0978_));
 sg13g2_and2_1 _3322_ (.A(_0977_),
    .B(_0664_),
    .X(_0666_));
 sg13g2_xnor2_1 _3323_ (.Y(_0667_),
    .A(_0661_),
    .B(_0666_));
 sg13g2_and2_1 _3324_ (.A(net126),
    .B(_0667_),
    .X(_0668_));
 sg13g2_inv_2 _3325_ (.Y(_0669_),
    .A(_1571_));
 sg13g2_nand2_1 _3326_ (.Y(_0670_),
    .A(net124),
    .B(\muldiv.regR[14] ));
 sg13g2_o21ai_1 _3327_ (.B1(_0670_),
    .Y(_0009_),
    .A1(_0660_),
    .A2(_0668_));
 sg13g2_nor2_1 _3328_ (.A(_1104_),
    .B(_0666_),
    .Y(_0671_));
 sg13g2_nand2_1 _3329_ (.Y(_0672_),
    .A(_0615_),
    .B(_0671_));
 sg13g2_nor2_1 _3330_ (.A(_0728_),
    .B(_0372_),
    .Y(_0673_));
 sg13g2_and2_1 _3331_ (.A(_0568_),
    .B(_0673_),
    .X(_0674_));
 sg13g2_nand2_1 _3332_ (.Y(_0676_),
    .A(_0227_),
    .B(_1164_));
 sg13g2_a21oi_1 _3333_ (.A1(net40),
    .A2(_0975_),
    .Y(_0677_),
    .B1(_0676_));
 sg13g2_a21oi_1 _3334_ (.A1(net62),
    .A2(_0674_),
    .Y(_0678_),
    .B1(_0677_));
 sg13g2_nor3_1 _3335_ (.A(_0449_),
    .B(_1581_),
    .C(_0678_),
    .Y(_0679_));
 sg13g2_a21oi_1 _3336_ (.A1(_0999_),
    .A2(_1002_),
    .Y(_0680_),
    .B1(_0449_));
 sg13g2_nor2_1 _3337_ (.A(_0449_),
    .B(_0678_),
    .Y(_0681_));
 sg13g2_a221oi_1 _3338_ (.B2(_0680_),
    .C1(_0681_),
    .B1(_0678_),
    .A1(_0977_),
    .Y(_0682_),
    .A2(_0664_));
 sg13g2_a21oi_1 _3339_ (.A1(_1575_),
    .A2(_1579_),
    .Y(_0683_),
    .B1(_0681_));
 sg13g2_a221oi_1 _3340_ (.B2(_0615_),
    .C1(_0683_),
    .B1(_0682_),
    .A1(_0672_),
    .Y(_0684_),
    .A2(_0679_));
 sg13g2_a21oi_1 _3341_ (.A1(net81),
    .A2(net61),
    .Y(_0685_),
    .B1(net119));
 sg13g2_and3_1 _3342_ (.X(_0687_),
    .A(_0637_),
    .B(_0643_),
    .C(_0685_));
 sg13g2_nor2_1 _3343_ (.A(net119),
    .B(_0653_),
    .Y(_0688_));
 sg13g2_and3_1 _3344_ (.X(_0689_),
    .A(_0637_),
    .B(_0643_),
    .C(_0688_));
 sg13g2_o21ai_1 _3345_ (.B1(net120),
    .Y(_0690_),
    .A1(_0557_),
    .A2(net108));
 sg13g2_nor2_1 _3346_ (.A(_0653_),
    .B(_0690_),
    .Y(_0691_));
 sg13g2_o21ai_1 _3347_ (.B1(net120),
    .Y(_0692_),
    .A1(_0650_),
    .A2(_0652_));
 sg13g2_a221oi_1 _3348_ (.B2(_0692_),
    .C1(_0641_),
    .B1(_0690_),
    .A1(_1576_),
    .Y(_0693_),
    .A2(_0638_));
 sg13g2_or2_1 _3349_ (.X(_0694_),
    .B(_0693_),
    .A(_0691_));
 sg13g2_nor2_1 _3350_ (.A(_1576_),
    .B(net61),
    .Y(_0695_));
 sg13g2_a21oi_1 _3351_ (.A1(net61),
    .A2(_0973_),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_and2_1 _3352_ (.A(_0637_),
    .B(_0696_),
    .X(_0698_));
 sg13g2_a221oi_1 _3353_ (.B2(_0643_),
    .C1(_0042_),
    .B1(_0698_),
    .A1(_0642_),
    .Y(_0699_),
    .A2(_0696_));
 sg13g2_nor4_2 _3354_ (.A(_0687_),
    .B(_0689_),
    .C(_0694_),
    .Y(_0700_),
    .D(_0699_));
 sg13g2_mux2_1 _3355_ (.A0(_0684_),
    .A1(_0700_),
    .S(net121),
    .X(_0701_));
 sg13g2_mux2_1 _3356_ (.A0(\muldiv.regR[15] ),
    .A1(_0701_),
    .S(net127),
    .X(_0010_));
 sg13g2_inv_1 _3357_ (.Y(_0702_),
    .A(_1304_));
 sg13g2_o21ai_1 _3358_ (.B1(_0471_),
    .Y(_0703_),
    .A1(_1562_),
    .A2(_1563_));
 sg13g2_nor2_1 _3359_ (.A(_1578_),
    .B(net48),
    .Y(_0704_));
 sg13g2_nor2b_1 _3360_ (.A(net67),
    .B_N(_0704_),
    .Y(_0705_));
 sg13g2_a21oi_1 _3361_ (.A1(net48),
    .A2(_1304_),
    .Y(_0706_),
    .B1(net40));
 sg13g2_nor2_1 _3362_ (.A(_0372_),
    .B(_1579_),
    .Y(_0708_));
 sg13g2_a21oi_1 _3363_ (.A1(_0557_),
    .A2(_0739_),
    .Y(_0709_),
    .B1(_0708_));
 sg13g2_nor2_1 _3364_ (.A(net82),
    .B(_0709_),
    .Y(_0710_));
 sg13g2_nor2_1 _3365_ (.A(net82),
    .B(_0372_),
    .Y(_0711_));
 sg13g2_a21oi_1 _3366_ (.A1(net82),
    .A2(_1311_),
    .Y(_0712_),
    .B1(_0711_));
 sg13g2_o21ai_1 _3367_ (.B1(net82),
    .Y(_0713_),
    .A1(_0673_),
    .A2(_0704_));
 sg13g2_o21ai_1 _3368_ (.B1(_0713_),
    .Y(_0714_),
    .A1(_1575_),
    .A2(_0712_));
 sg13g2_nor4_1 _3369_ (.A(_0705_),
    .B(_0706_),
    .C(_0710_),
    .D(_0714_),
    .Y(_0715_));
 sg13g2_a22oi_1 _3370_ (.Y(_0716_),
    .B1(_0715_),
    .B2(_1559_),
    .A2(_0703_),
    .A1(_0702_));
 sg13g2_nor2_1 _3371_ (.A(_1577_),
    .B(_1515_),
    .Y(_0717_));
 sg13g2_xor2_1 _3372_ (.B(_0717_),
    .A(net36),
    .X(_0719_));
 sg13g2_xor2_1 _3373_ (.B(_0719_),
    .A(_0716_),
    .X(_0720_));
 sg13g2_nand2_1 _3374_ (.Y(_0721_),
    .A(_1436_),
    .B(net48));
 sg13g2_xor2_1 _3375_ (.B(_0721_),
    .A(_1601_),
    .X(_0722_));
 sg13g2_nor2_1 _3376_ (.A(net128),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_a21o_1 _3377_ (.A2(_0720_),
    .A1(net126),
    .B1(_0723_),
    .X(_0724_));
 sg13g2_mux2_1 _3378_ (.A0(\muldiv.regR[1] ),
    .A1(_0724_),
    .S(net127),
    .X(_0011_));
 sg13g2_a21o_1 _3379_ (.A2(_1457_),
    .A1(_1449_),
    .B1(net43),
    .X(_0725_));
 sg13g2_nand3_1 _3380_ (.B(_1449_),
    .C(_1457_),
    .A(_1229_),
    .Y(_0726_));
 sg13g2_and2_1 _3381_ (.A(_0725_),
    .B(_0726_),
    .X(_0727_));
 sg13g2_a21oi_1 _3382_ (.A1(net19),
    .A2(net20),
    .Y(_0729_),
    .B1(_0727_));
 sg13g2_xnor2_1 _3383_ (.Y(_0730_),
    .A(net50),
    .B(_1306_));
 sg13g2_xnor2_1 _3384_ (.Y(_0731_),
    .A(_1515_),
    .B(_0730_));
 sg13g2_xor2_1 _3385_ (.B(_1434_),
    .A(net48),
    .X(_0732_));
 sg13g2_nor3_1 _3386_ (.A(_1436_),
    .B(net40),
    .C(_0732_),
    .Y(_0733_));
 sg13g2_a21o_1 _3387_ (.A2(_0731_),
    .A1(_1588_),
    .B1(_0733_),
    .X(_0734_));
 sg13g2_buf_1 _3388_ (.A(_0734_),
    .X(_0735_));
 sg13g2_nor2_1 _3389_ (.A(net67),
    .B(_0735_),
    .Y(_0736_));
 sg13g2_nand2_1 _3390_ (.Y(_0737_),
    .A(_0729_),
    .B(_0736_));
 sg13g2_or2_1 _3391_ (.X(_0738_),
    .B(_0729_),
    .A(_1303_));
 sg13g2_xnor2_1 _3392_ (.Y(_0740_),
    .A(_1466_),
    .B(_1469_));
 sg13g2_buf_1 _3393_ (.A(_0740_),
    .X(_0741_));
 sg13g2_a21o_1 _3394_ (.A2(_0738_),
    .A1(_0737_),
    .B1(net21),
    .X(_0742_));
 sg13g2_nand2_1 _3395_ (.Y(_0743_),
    .A(_0727_),
    .B(_0735_));
 sg13g2_and2_1 _3396_ (.A(net96),
    .B(_0719_),
    .X(_0744_));
 sg13g2_buf_1 _3397_ (.A(_0744_),
    .X(_0745_));
 sg13g2_nand3_1 _3398_ (.B(net20),
    .C(_0745_),
    .A(net19),
    .Y(_0746_));
 sg13g2_o21ai_1 _3399_ (.B1(_0746_),
    .Y(_0747_),
    .A1(_1565_),
    .A2(_0743_));
 sg13g2_nor2_1 _3400_ (.A(net67),
    .B(_0741_),
    .Y(_0748_));
 sg13g2_nor2_1 _3401_ (.A(net67),
    .B(_1471_),
    .Y(_0749_));
 sg13g2_or2_1 _3402_ (.X(_0751_),
    .B(_0735_),
    .A(_0727_));
 sg13g2_a22oi_1 _3403_ (.Y(_0752_),
    .B1(_0743_),
    .B2(_0751_),
    .A2(net20),
    .A1(net19));
 sg13g2_a21oi_1 _3404_ (.A1(_1565_),
    .A2(_0745_),
    .Y(_0753_),
    .B1(_0752_));
 sg13g2_nor2_1 _3405_ (.A(_1303_),
    .B(_1471_),
    .Y(_0754_));
 sg13g2_a21o_1 _3406_ (.A2(_0754_),
    .A1(_0729_),
    .B1(_1573_),
    .X(_0755_));
 sg13g2_a221oi_1 _3407_ (.B2(_0753_),
    .C1(_0755_),
    .B1(_0749_),
    .A1(_0747_),
    .Y(_0756_),
    .A2(_0748_));
 sg13g2_xnor2_1 _3408_ (.Y(_0757_),
    .A(_1355_),
    .B(_0289_));
 sg13g2_nor2_1 _3409_ (.A(net40),
    .B(net59),
    .Y(_0758_));
 sg13g2_nor2_1 _3410_ (.A(_1311_),
    .B(_1300_),
    .Y(_0759_));
 sg13g2_a22oi_1 _3411_ (.Y(_0760_),
    .B1(_0758_),
    .B2(_0759_),
    .A2(_0757_),
    .A1(net40));
 sg13g2_nor2_1 _3412_ (.A(_1523_),
    .B(_0760_),
    .Y(_0762_));
 sg13g2_nand2_1 _3413_ (.Y(_0763_),
    .A(net55),
    .B(net59));
 sg13g2_o21ai_1 _3414_ (.B1(_1523_),
    .Y(_0764_),
    .A1(net55),
    .A2(_1631_));
 sg13g2_a21oi_1 _3415_ (.A1(_0763_),
    .A2(_0764_),
    .Y(_0765_),
    .B1(_0759_));
 sg13g2_nand3_1 _3416_ (.B(_0289_),
    .C(_0759_),
    .A(net40),
    .Y(_0766_));
 sg13g2_o21ai_1 _3417_ (.B1(_1573_),
    .Y(_0767_),
    .A1(net82),
    .A2(_0766_));
 sg13g2_nor3_1 _3418_ (.A(_0762_),
    .B(_0765_),
    .C(_0767_),
    .Y(_0768_));
 sg13g2_a21o_1 _3419_ (.A2(_0756_),
    .A1(_0742_),
    .B1(_0768_),
    .X(_0769_));
 sg13g2_mux2_1 _3420_ (.A0(\muldiv.regR[2] ),
    .A1(_0769_),
    .S(_1572_),
    .X(_0012_));
 sg13g2_nand3_1 _3421_ (.B(_0725_),
    .C(_0726_),
    .A(net21),
    .Y(_0770_));
 sg13g2_a21o_1 _3422_ (.A2(_0726_),
    .A1(_0725_),
    .B1(net21),
    .X(_0772_));
 sg13g2_nand3_1 _3423_ (.B(_0770_),
    .C(_0772_),
    .A(_0735_),
    .Y(_0773_));
 sg13g2_nor3_1 _3424_ (.A(net39),
    .B(_1458_),
    .C(_1471_),
    .Y(_0774_));
 sg13g2_and2_1 _3425_ (.A(_1449_),
    .B(_1457_),
    .X(_0775_));
 sg13g2_buf_1 _3426_ (.A(_0775_),
    .X(_0776_));
 sg13g2_nor3_1 _3427_ (.A(net41),
    .B(_0776_),
    .C(net21),
    .Y(_0777_));
 sg13g2_nor2_1 _3428_ (.A(net39),
    .B(_1229_),
    .Y(_0778_));
 sg13g2_nor2_1 _3429_ (.A(net41),
    .B(_1327_),
    .Y(_0779_));
 sg13g2_mux2_1 _3430_ (.A0(_0778_),
    .A1(_0779_),
    .S(_1471_),
    .X(_0780_));
 sg13g2_mux2_1 _3431_ (.A0(_0778_),
    .A1(_0779_),
    .S(_1458_),
    .X(_0781_));
 sg13g2_nor4_2 _3432_ (.A(_0774_),
    .B(_0777_),
    .C(_0780_),
    .Y(_0783_),
    .D(_0781_));
 sg13g2_nand3_1 _3433_ (.B(_0773_),
    .C(_0783_),
    .A(_1303_),
    .Y(_0784_));
 sg13g2_a21oi_1 _3434_ (.A1(net19),
    .A2(net20),
    .Y(_0785_),
    .B1(_0784_));
 sg13g2_a21o_1 _3435_ (.A2(_0745_),
    .A1(_1471_),
    .B1(net67),
    .X(_0786_));
 sg13g2_nor3_1 _3436_ (.A(_1562_),
    .B(_1563_),
    .C(_0786_),
    .Y(_0787_));
 sg13g2_a221oi_1 _3437_ (.B2(_1303_),
    .C1(_0783_),
    .B1(_0773_),
    .A1(net19),
    .Y(_0788_),
    .A2(net20));
 sg13g2_or3_1 _3438_ (.A(_0785_),
    .B(_0787_),
    .C(_0788_),
    .X(_0789_));
 sg13g2_xnor2_1 _3439_ (.Y(_0790_),
    .A(_1487_),
    .B(_0789_));
 sg13g2_nand2_1 _3440_ (.Y(_0791_),
    .A(net40),
    .B(net97));
 sg13g2_xor2_1 _3441_ (.B(_0791_),
    .A(net31),
    .X(_0792_));
 sg13g2_nor2_1 _3442_ (.A(net128),
    .B(_0792_),
    .Y(_0794_));
 sg13g2_a21oi_1 _3443_ (.A1(net126),
    .A2(_0790_),
    .Y(_0795_),
    .B1(_0794_));
 sg13g2_nor2_1 _3444_ (.A(net125),
    .B(\muldiv.regR[3] ),
    .Y(_0796_));
 sg13g2_a21oi_1 _3445_ (.A1(_1572_),
    .A2(_0795_),
    .Y(_0013_),
    .B1(_0796_));
 sg13g2_xnor2_1 _3446_ (.Y(_0797_),
    .A(net67),
    .B(_1482_));
 sg13g2_nor2_1 _3447_ (.A(_1367_),
    .B(_1293_),
    .Y(_0798_));
 sg13g2_nor2_1 _3448_ (.A(_1367_),
    .B(_1295_),
    .Y(_0799_));
 sg13g2_mux2_1 _3449_ (.A0(_0798_),
    .A1(_0799_),
    .S(_1425_),
    .X(_0800_));
 sg13g2_nor2_1 _3450_ (.A(net37),
    .B(_0800_),
    .Y(_0801_));
 sg13g2_nand2_1 _3451_ (.Y(_0802_),
    .A(_1472_),
    .B(_1474_));
 sg13g2_a221oi_1 _3452_ (.B2(net41),
    .C1(net35),
    .B1(_1487_),
    .A1(_1458_),
    .Y(_0804_),
    .A2(_1471_));
 sg13g2_nor2_1 _3453_ (.A(_1720_),
    .B(_1295_),
    .Y(_0805_));
 sg13g2_nor2_1 _3454_ (.A(_1720_),
    .B(_1293_),
    .Y(_0806_));
 sg13g2_mux2_1 _3455_ (.A0(_0805_),
    .A1(_0806_),
    .S(_1425_),
    .X(_0807_));
 sg13g2_mux2_1 _3456_ (.A0(_0800_),
    .A1(_0807_),
    .S(net35),
    .X(_0808_));
 sg13g2_a21o_1 _3457_ (.A2(_0804_),
    .A1(_1474_),
    .B1(_0808_),
    .X(_0809_));
 sg13g2_a221oi_1 _3458_ (.B2(_0802_),
    .C1(_0809_),
    .B1(_0801_),
    .A1(_1543_),
    .Y(_0810_),
    .A2(_1558_));
 sg13g2_xnor2_1 _3459_ (.Y(_0811_),
    .A(_0797_),
    .B(_0810_));
 sg13g2_nand3_1 _3460_ (.B(_0745_),
    .C(_0748_),
    .A(_1487_),
    .Y(_0812_));
 sg13g2_inv_1 _3461_ (.Y(_0813_),
    .A(_0812_));
 sg13g2_or2_1 _3462_ (.X(_0815_),
    .B(_0783_),
    .A(_1487_));
 sg13g2_nand2_1 _3463_ (.Y(_0816_),
    .A(_1487_),
    .B(_0783_));
 sg13g2_or2_1 _3464_ (.X(_0817_),
    .B(_0773_),
    .A(_0240_));
 sg13g2_a221oi_1 _3465_ (.B2(_0816_),
    .C1(_0817_),
    .B1(_0815_),
    .A1(_1543_),
    .Y(_0818_),
    .A2(_1558_));
 sg13g2_a21oi_1 _3466_ (.A1(_1565_),
    .A2(_0813_),
    .Y(_0819_),
    .B1(_0818_));
 sg13g2_inv_1 _3467_ (.Y(_0820_),
    .A(_0797_));
 sg13g2_nor2_1 _3468_ (.A(_0776_),
    .B(net21),
    .Y(_0821_));
 sg13g2_a21oi_1 _3469_ (.A1(_0776_),
    .A2(net21),
    .Y(_0822_),
    .B1(_1327_));
 sg13g2_o21ai_1 _3470_ (.B1(_0801_),
    .Y(_0823_),
    .A1(_0821_),
    .A2(_0822_));
 sg13g2_a21oi_1 _3471_ (.A1(_1474_),
    .A2(_0804_),
    .Y(_0824_),
    .B1(_0808_));
 sg13g2_nand3_1 _3472_ (.B(_0823_),
    .C(_0824_),
    .A(_0820_),
    .Y(_0826_));
 sg13g2_a21o_1 _3473_ (.A2(_0824_),
    .A1(_0823_),
    .B1(_0820_),
    .X(_0827_));
 sg13g2_a221oi_1 _3474_ (.B2(_0827_),
    .C1(_0817_),
    .B1(_0826_),
    .A1(_0815_),
    .Y(_0828_),
    .A2(_0816_));
 sg13g2_nor4_1 _3475_ (.A(_1562_),
    .B(_1563_),
    .C(_0820_),
    .D(_0812_),
    .Y(_0829_));
 sg13g2_a21o_1 _3476_ (.A2(_0828_),
    .A1(_1559_),
    .B1(_0829_),
    .X(_0830_));
 sg13g2_buf_1 _3477_ (.A(_0830_),
    .X(_0831_));
 sg13g2_a21oi_1 _3478_ (.A1(_0811_),
    .A2(_0819_),
    .Y(_0832_),
    .B1(_0831_));
 sg13g2_nand3_1 _3479_ (.B(_1670_),
    .C(net31),
    .A(net71),
    .Y(_0833_));
 sg13g2_o21ai_1 _3480_ (.B1(_0833_),
    .Y(_0834_),
    .A1(net71),
    .A2(net31));
 sg13g2_a21o_1 _3481_ (.A2(_1697_),
    .A1(net48),
    .B1(net89),
    .X(_0835_));
 sg13g2_a22oi_1 _3482_ (.Y(_0837_),
    .B1(_0835_),
    .B2(net56),
    .A2(_0834_),
    .A1(net86));
 sg13g2_o21ai_1 _3483_ (.B1(net40),
    .Y(_0838_),
    .A1(_0408_),
    .A2(_1697_));
 sg13g2_nand2b_1 _3484_ (.Y(_0839_),
    .B(_0838_),
    .A_N(_0025_));
 sg13g2_o21ai_1 _3485_ (.B1(_0839_),
    .Y(_0840_),
    .A1(net55),
    .A2(_0837_));
 sg13g2_xnor2_1 _3486_ (.Y(_0841_),
    .A(_1695_),
    .B(_0840_));
 sg13g2_nor2_1 _3487_ (.A(net128),
    .B(_0841_),
    .Y(_0842_));
 sg13g2_a21o_1 _3488_ (.A2(_0832_),
    .A1(net126),
    .B1(_0842_),
    .X(_0843_));
 sg13g2_mux2_1 _3489_ (.A0(\muldiv.regR[4] ),
    .A1(_0843_),
    .S(net125),
    .X(_0014_));
 sg13g2_o21ai_1 _3490_ (.B1(_1508_),
    .Y(_0844_),
    .A1(_1485_),
    .A2(_1491_));
 sg13g2_or3_1 _3491_ (.A(_1508_),
    .B(_1485_),
    .C(_1491_),
    .X(_0845_));
 sg13g2_a22oi_1 _3492_ (.Y(_0847_),
    .B1(_0844_),
    .B2(_0845_),
    .A2(net20),
    .A1(net19));
 sg13g2_xnor2_1 _3493_ (.Y(_0848_),
    .A(_1303_),
    .B(_1549_));
 sg13g2_xnor2_1 _3494_ (.Y(_0849_),
    .A(_0847_),
    .B(_0848_));
 sg13g2_xnor2_1 _3495_ (.Y(_0850_),
    .A(_0831_),
    .B(_0849_));
 sg13g2_nand2_1 _3496_ (.Y(_0851_),
    .A(_0211_),
    .B(_0072_));
 sg13g2_a21oi_1 _3497_ (.A1(_0213_),
    .A2(_0851_),
    .Y(_0852_),
    .B1(net128));
 sg13g2_a21oi_1 _3498_ (.A1(net126),
    .A2(_0850_),
    .Y(_0853_),
    .B1(_0852_));
 sg13g2_mux2_1 _3499_ (.A0(\muldiv.regR[5] ),
    .A1(_0853_),
    .S(net125),
    .X(_0015_));
 sg13g2_o21ai_1 _3500_ (.B1(net21),
    .Y(_0854_),
    .A1(_1197_),
    .A2(_0776_));
 sg13g2_inv_1 _3501_ (.Y(_0855_),
    .A(_1196_));
 sg13g2_nand2_1 _3502_ (.Y(_0857_),
    .A(_0227_),
    .B(_0728_));
 sg13g2_nand2_1 _3503_ (.Y(_0858_),
    .A(_1460_),
    .B(_1442_));
 sg13g2_nand2_1 _3504_ (.Y(_0859_),
    .A(_1385_),
    .B(_1447_));
 sg13g2_nand2_1 _3505_ (.Y(_0860_),
    .A(_1454_),
    .B(_1455_));
 sg13g2_a221oi_1 _3506_ (.B2(_0859_),
    .C1(_0860_),
    .B1(_0858_),
    .A1(_1196_),
    .Y(_0861_),
    .A2(_0857_));
 sg13g2_a221oi_1 _3507_ (.B2(net39),
    .C1(_0861_),
    .B1(_1426_),
    .A1(_0855_),
    .Y(_0862_),
    .A2(net21));
 sg13g2_inv_1 _3508_ (.Y(_0863_),
    .A(_1482_));
 sg13g2_nand2b_1 _3509_ (.Y(_0864_),
    .B(_1549_),
    .A_N(_0807_));
 sg13g2_a221oi_1 _3510_ (.B2(_1371_),
    .C1(_0864_),
    .B1(_0863_),
    .A1(_0854_),
    .Y(_0865_),
    .A2(_0862_));
 sg13g2_nand2b_1 _3511_ (.Y(_0866_),
    .B(net34),
    .A_N(_0807_));
 sg13g2_a221oi_1 _3512_ (.B2(_1371_),
    .C1(_0866_),
    .B1(_0863_),
    .A1(_0854_),
    .Y(_0868_),
    .A2(_0862_));
 sg13g2_nand2_1 _3513_ (.Y(_0869_),
    .A(net34),
    .B(_1549_));
 sg13g2_nand3_1 _3514_ (.B(_1482_),
    .C(_1549_),
    .A(_1281_),
    .Y(_0870_));
 sg13g2_nand3_1 _3515_ (.B(net34),
    .C(_1482_),
    .A(_1281_),
    .Y(_0871_));
 sg13g2_nand3_1 _3516_ (.B(_0870_),
    .C(_0871_),
    .A(_0869_),
    .Y(_0872_));
 sg13g2_nor3_1 _3517_ (.A(_0865_),
    .B(_0868_),
    .C(_0872_),
    .Y(_0873_));
 sg13g2_xnor2_1 _3518_ (.Y(_0874_),
    .A(net44),
    .B(_0873_));
 sg13g2_nor2_1 _3519_ (.A(_1515_),
    .B(_1516_),
    .Y(_0875_));
 sg13g2_xnor2_1 _3520_ (.Y(_0876_),
    .A(_1405_),
    .B(_0875_));
 sg13g2_xnor2_1 _3521_ (.Y(_0877_),
    .A(_1303_),
    .B(_0876_));
 sg13g2_o21ai_1 _3522_ (.B1(_0877_),
    .Y(_0879_),
    .A1(_1565_),
    .A2(_0874_));
 sg13g2_or3_1 _3523_ (.A(_1565_),
    .B(_0877_),
    .C(_0874_),
    .X(_0880_));
 sg13g2_buf_1 _3524_ (.A(_0880_),
    .X(_0881_));
 sg13g2_a22oi_1 _3525_ (.Y(_0882_),
    .B1(_0879_),
    .B2(_0881_),
    .A2(_0849_),
    .A1(_0831_));
 sg13g2_and4_1 _3526_ (.A(_0831_),
    .B(_0849_),
    .C(_0879_),
    .D(_0881_),
    .X(_0883_));
 sg13g2_nor3_1 _3527_ (.A(net121),
    .B(_0882_),
    .C(_0883_),
    .Y(_0884_));
 sg13g2_xnor2_1 _3528_ (.Y(_0885_),
    .A(_0088_),
    .B(_0102_));
 sg13g2_nor2_1 _3529_ (.A(_0103_),
    .B(_0885_),
    .Y(_0886_));
 sg13g2_o21ai_1 _3530_ (.B1(_1573_),
    .Y(_0887_),
    .A1(_0109_),
    .A2(_0886_));
 sg13g2_nand2_1 _3531_ (.Y(_0888_),
    .A(net125),
    .B(_0887_));
 sg13g2_nand2_1 _3532_ (.Y(_0890_),
    .A(net124),
    .B(\muldiv.regR[6] ));
 sg13g2_o21ai_1 _3533_ (.B1(_0890_),
    .Y(_0016_),
    .A1(_0884_),
    .A2(_0888_));
 sg13g2_o21ai_1 _3534_ (.B1(_1546_),
    .Y(_0891_),
    .A1(_1539_),
    .A2(_0873_));
 sg13g2_xnor2_1 _3535_ (.Y(_0892_),
    .A(_0108_),
    .B(_1511_));
 sg13g2_nor2_1 _3536_ (.A(_1451_),
    .B(_0892_),
    .Y(_0893_));
 sg13g2_a21oi_1 _3537_ (.A1(_0891_),
    .A2(_0893_),
    .Y(_0894_),
    .B1(_0240_));
 sg13g2_nor2_1 _3538_ (.A(_0064_),
    .B(_1451_),
    .Y(_0895_));
 sg13g2_nor4_1 _3539_ (.A(_1303_),
    .B(net65),
    .C(_1451_),
    .D(_0892_),
    .Y(_0896_));
 sg13g2_mux2_1 _3540_ (.A0(_0895_),
    .A1(_0896_),
    .S(_0891_),
    .X(_0897_));
 sg13g2_o21ai_1 _3541_ (.B1(net128),
    .Y(_0898_),
    .A1(_0894_),
    .A2(_0897_));
 sg13g2_or3_1 _3542_ (.A(_1573_),
    .B(_0894_),
    .C(_0897_),
    .X(_0900_));
 sg13g2_or2_1 _3543_ (.X(_0901_),
    .B(_0848_),
    .A(_0847_));
 sg13g2_nand2_1 _3544_ (.Y(_0902_),
    .A(_0847_),
    .B(_0848_));
 sg13g2_a21oi_1 _3545_ (.A1(_1559_),
    .A2(_0828_),
    .Y(_0903_),
    .B1(_0829_));
 sg13g2_a221oi_1 _3546_ (.B2(_0881_),
    .C1(_0903_),
    .B1(_0879_),
    .A1(_0901_),
    .Y(_0904_),
    .A2(_0902_));
 sg13g2_mux2_1 _3547_ (.A0(_0898_),
    .A1(_0900_),
    .S(_0904_),
    .X(_0905_));
 sg13g2_nand2_1 _3548_ (.Y(_0906_),
    .A(_1586_),
    .B(net81));
 sg13g2_xor2_1 _3549_ (.B(_0906_),
    .A(_0112_),
    .X(_0907_));
 sg13g2_a21oi_1 _3550_ (.A1(net121),
    .A2(_0907_),
    .Y(_0908_),
    .B1(net124));
 sg13g2_nor2_1 _3551_ (.A(net131),
    .B(\muldiv.regR[7] ),
    .Y(_0909_));
 sg13g2_a21oi_1 _3552_ (.A1(_0905_),
    .A2(_0908_),
    .Y(_0017_),
    .B1(_0909_));
 sg13g2_nand2_1 _3553_ (.Y(_0911_),
    .A(net81),
    .B(_0114_));
 sg13g2_xnor2_1 _3554_ (.Y(_0912_),
    .A(_0911_),
    .B(_0263_));
 sg13g2_xnor2_1 _3555_ (.Y(_0913_),
    .A(_0259_),
    .B(_0912_));
 sg13g2_o21ai_1 _3556_ (.B1(_1560_),
    .Y(_0914_),
    .A1(_0494_),
    .A2(_0913_));
 sg13g2_mux2_1 _3557_ (.A0(\muldiv.regR[8] ),
    .A1(_0914_),
    .S(net125),
    .X(_0018_));
 sg13g2_nor2_1 _3558_ (.A(_1565_),
    .B(_1581_),
    .Y(_0915_));
 sg13g2_xor2_1 _3559_ (.B(_0915_),
    .A(_1515_),
    .X(_0916_));
 sg13g2_xor2_1 _3560_ (.B(_0393_),
    .A(_0396_),
    .X(_0917_));
 sg13g2_xnor2_1 _3561_ (.Y(_0918_),
    .A(_0265_),
    .B(_0917_));
 sg13g2_nor2_1 _3562_ (.A(_1561_),
    .B(_0918_),
    .Y(_0920_));
 sg13g2_a21oi_1 _3563_ (.A1(_0494_),
    .A2(_0916_),
    .Y(_0921_),
    .B1(_0920_));
 sg13g2_mux2_1 _3564_ (.A0(\muldiv.regR[9] ),
    .A1(_0921_),
    .S(_0554_),
    .X(_0019_));
 sg13g2_and2_1 _3565_ (.A(_0000_),
    .B(net132),
    .X(_0002_));
 sg13g2_nand2b_1 _3566_ (.Y(_0003_),
    .B(net133),
    .A_N(\muldiv.div2reg ));
 sg13g2_nor2b_2 _3567_ (.A(\muldiv.div2reg ),
    .B_N(\muldiv.negedgeReg_1.area_io_q ),
    .Y(\muldiv.a0_0.GATE ));
 sg13g2_nor2b_2 _3568_ (.A(\muldiv.negedgeReg_1.area_io_q ),
    .B_N(\muldiv.div2reg ),
    .Y(\muldiv.a1_0.GATE ));
 sg13g2_nand2_1 _3569_ (.Y(_0922_),
    .A(net79),
    .B(_0416_));
 sg13g2_nor4_1 _3570_ (.A(net62),
    .B(_1574_),
    .C(_0922_),
    .D(_0471_),
    .Y(\muldiv.div8.io_edivzero ));
 sg13g2_buf_1 _3571_ (.A(uio_in[3]),
    .X(_0924_));
 sg13g2_buf_1 _3572_ (.A(net130),
    .X(_0925_));
 sg13g2_mux4_1 _3573_ (.S0(_0554_),
    .A0(_1570_),
    .A1(_0914_),
    .A2(\muldiv.regR[0] ),
    .A3(\muldiv.regR[8] ),
    .S1(net123),
    .X(net11));
 sg13g2_mux4_1 _3574_ (.S0(net131),
    .A0(_0724_),
    .A1(_0921_),
    .A2(\muldiv.regR[1] ),
    .A3(\muldiv.regR[9] ),
    .S1(net123),
    .X(net12));
 sg13g2_mux4_1 _3575_ (.S0(_0669_),
    .A0(_0492_),
    .A1(_0769_),
    .A2(\muldiv.regR[10] ),
    .A3(\muldiv.regR[2] ),
    .S1(net123),
    .X(net13));
 sg13g2_nor2_1 _3576_ (.A(net131),
    .B(net123),
    .Y(_0926_));
 sg13g2_nor2_1 _3577_ (.A(net124),
    .B(net123),
    .Y(_0927_));
 sg13g2_nand2_1 _3578_ (.Y(_0928_),
    .A(net124),
    .B(net130));
 sg13g2_nand3b_1 _3579_ (.B(_0924_),
    .C(net131),
    .Y(_0929_),
    .A_N(\muldiv.regR[11] ));
 sg13g2_o21ai_1 _3580_ (.B1(_0929_),
    .Y(_0930_),
    .A1(\muldiv.regR[3] ),
    .A2(_0928_));
 sg13g2_a221oi_1 _3581_ (.B2(_0553_),
    .C1(_0930_),
    .B1(_0927_),
    .A1(_0795_),
    .Y(net14),
    .A2(_0926_));
 sg13g2_mux4_1 _3582_ (.S0(_0669_),
    .A0(_0610_),
    .A1(_0843_),
    .A2(\muldiv.regR[12] ),
    .A3(\muldiv.regR[4] ),
    .S1(_0925_),
    .X(net15));
 sg13g2_mux4_1 _3583_ (.S0(net124),
    .A0(_0648_),
    .A1(_0853_),
    .A2(\muldiv.regR[13] ),
    .A3(\muldiv.regR[5] ),
    .S1(_0925_),
    .X(net16));
 sg13g2_nand2_1 _3584_ (.Y(_0932_),
    .A(\muldiv.regR[14] ),
    .B(net130));
 sg13g2_nor2_1 _3585_ (.A(net131),
    .B(\muldiv.regR[6] ),
    .Y(_0933_));
 sg13g2_a22oi_1 _3586_ (.Y(_0934_),
    .B1(_0933_),
    .B2(net130),
    .A2(_0932_),
    .A1(net131));
 sg13g2_inv_1 _3587_ (.Y(_0935_),
    .A(_0934_));
 sg13g2_a21o_1 _3588_ (.A2(_0667_),
    .A1(net126),
    .B1(net123),
    .X(_0936_));
 sg13g2_or2_1 _3589_ (.X(_0937_),
    .B(_0887_),
    .A(net130));
 sg13g2_a22oi_1 _3590_ (.Y(_0938_),
    .B1(_0934_),
    .B2(_0937_),
    .A2(_0659_),
    .A1(net125));
 sg13g2_a221oi_1 _3591_ (.B2(_0936_),
    .C1(_0938_),
    .B1(_0935_),
    .A1(_0884_),
    .Y(net17),
    .A2(_0926_));
 sg13g2_mux2_1 _3592_ (.A0(_0700_),
    .A1(_0907_),
    .S(net124),
    .X(_0940_));
 sg13g2_nor2_1 _3593_ (.A(net121),
    .B(net124),
    .Y(_0941_));
 sg13g2_a221oi_1 _3594_ (.B2(_0684_),
    .C1(net123),
    .B1(_0941_),
    .A1(net121),
    .Y(_0942_),
    .A2(_0940_));
 sg13g2_nor2_1 _3595_ (.A(net128),
    .B(net130),
    .Y(_0943_));
 sg13g2_nor2_1 _3596_ (.A(net121),
    .B(net130),
    .Y(_0944_));
 sg13g2_and2_1 _3597_ (.A(\muldiv.regR[15] ),
    .B(net130),
    .X(_0945_));
 sg13g2_a221oi_1 _3598_ (.B2(_0684_),
    .C1(_0945_),
    .B1(_0944_),
    .A1(_0700_),
    .Y(_0946_),
    .A2(_0943_));
 sg13g2_and2_1 _3599_ (.A(net123),
    .B(_0909_),
    .X(_0947_));
 sg13g2_a221oi_1 _3600_ (.B2(net127),
    .C1(_0947_),
    .B1(_0946_),
    .A1(_0905_),
    .Y(net18),
    .A2(_0942_));
 sg13g2_inv_1 _1805__1 (.Y(net168),
    .A(clknet_2_1__leaf_clk));
 sg13g2_tiehi _3607__148 (.L_HI(net148));
 sg13g2_buf_1 _3603_ (.A(net135),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3604_ (.A(net136),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3605_ (.A(net137),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3606_ (.A(net138),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3607_ (.A(net148),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3608_ (.A(net149),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3609_ (.A(net139),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3610_ (.A(net140),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3611_ (.A(net141),
    .X(uio_out[0]));
 sg13g2_buf_1 _3612_ (.A(net142),
    .X(uio_out[1]));
 sg13g2_buf_1 _3613_ (.A(net143),
    .X(uio_out[2]));
 sg13g2_buf_1 _3614_ (.A(net144),
    .X(uio_out[3]));
 sg13g2_buf_1 _3615_ (.A(net145),
    .X(uio_out[4]));
 sg13g2_buf_1 _3616_ (.A(\muldiv.div8.io_edivzero ),
    .X(net10));
 sg13g2_buf_1 _3617_ (.A(net146),
    .X(uio_out[6]));
 sg13g2_buf_1 _3618_ (.A(net147),
    .X(uio_out[7]));
 sg13g2_dlhrq_1 \muldiv.a0_0.genblk1.dlhrq_1  (.D(net2),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net133),
    .Q(\muldiv.a0_0.Q ));
 sg13g2_dlhrq_1 \muldiv.a0_1.genblk1.dlhrq_1  (.D(net3),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net133),
    .Q(\muldiv.a0_1.Q ));
 sg13g2_dlhrq_1 \muldiv.a0_2.genblk1.dlhrq_1  (.D(net4),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net133),
    .Q(\muldiv.a0_2.Q ));
 sg13g2_dlhrq_1 \muldiv.a0_3.genblk1.dlhrq_1  (.D(net5),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net134),
    .Q(\muldiv.a0_3.Q ));
 sg13g2_dlhrq_1 \muldiv.a0_4.genblk1.dlhrq_1  (.D(net6),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net132),
    .Q(\muldiv.a0_4.Q ));
 sg13g2_dlhrq_1 \muldiv.a0_5.genblk1.dlhrq_1  (.D(net7),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net132),
    .Q(\muldiv.a0_5.Q ));
 sg13g2_dlhrq_1 \muldiv.a0_6.genblk1.dlhrq_1  (.D(net8),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net132),
    .Q(\muldiv.a0_6.Q ));
 sg13g2_dlhrq_1 \muldiv.a0_7.genblk1.dlhrq_1  (.D(net9),
    .GATE(\muldiv.a0_0.GATE ),
    .RESET_B(net132),
    .Q(\muldiv.a0_7.Q ));
 sg13g2_dlhrq_1 \muldiv.a1_0.genblk1.dlhrq_1  (.D(net2),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net133),
    .Q(\muldiv.a1_0.Q ));
 sg13g2_dlhrq_1 \muldiv.a1_1.genblk1.dlhrq_1  (.D(net3),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net133),
    .Q(\muldiv.a1_1.Q ));
 sg13g2_dlhrq_1 \muldiv.a1_2.genblk1.dlhrq_1  (.D(net4),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net133),
    .Q(\muldiv.a1_2.Q ));
 sg13g2_dlhrq_1 \muldiv.a1_3.genblk1.dlhrq_1  (.D(net5),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net133),
    .Q(\muldiv.a1_3.Q ));
 sg13g2_dlhrq_1 \muldiv.a1_4.genblk1.dlhrq_1  (.D(net6),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net132),
    .Q(\muldiv.a1_4.Q ));
 sg13g2_dlhrq_1 \muldiv.a1_5.genblk1.dlhrq_1  (.D(net7),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net132),
    .Q(\muldiv.a1_5.Q ));
 sg13g2_dlhrq_1 \muldiv.a1_6.genblk1.dlhrq_1  (.D(net8),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net132),
    .Q(\muldiv.a1_6.Q ));
 sg13g2_dlhrq_1 \muldiv.a1_7.genblk1.dlhrq_1  (.D(net9),
    .GATE(\muldiv.a1_0.GATE ),
    .RESET_B(net134),
    .Q(\muldiv.a1_7.Q ));
 sg13g2_dfrbp_1 \muldiv.div2reg$_SDFF_PN0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net150),
    .D(_0002_),
    .Q_N(_0000_),
    .Q(\muldiv.div2reg ));
 sg13g2_dfrbp_1 \muldiv.negedgeReg_1.area_io_q$_SDFF_NN1_  (.CLK(net168),
    .RESET_B(net151),
    .D(_0003_),
    .Q_N(_1802_),
    .Q(\muldiv.negedgeReg_1.area_io_q ));
 sg13g2_dfrbp_1 \muldiv.regR[0]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net152),
    .D(_0004_),
    .Q_N(_1801_),
    .Q(\muldiv.regR[0] ));
 sg13g2_dfrbp_1 \muldiv.regR[10]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net153),
    .D(_0005_),
    .Q_N(_1800_),
    .Q(\muldiv.regR[10] ));
 sg13g2_dfrbp_1 \muldiv.regR[11]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net154),
    .D(_0006_),
    .Q_N(_1799_),
    .Q(\muldiv.regR[11] ));
 sg13g2_dfrbp_1 \muldiv.regR[12]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net155),
    .D(_0007_),
    .Q_N(_1798_),
    .Q(\muldiv.regR[12] ));
 sg13g2_dfrbp_1 \muldiv.regR[13]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net156),
    .D(_0008_),
    .Q_N(_1797_),
    .Q(\muldiv.regR[13] ));
 sg13g2_dfrbp_1 \muldiv.regR[14]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net157),
    .D(_0009_),
    .Q_N(_1796_),
    .Q(\muldiv.regR[14] ));
 sg13g2_dfrbp_1 \muldiv.regR[15]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net158),
    .D(_0010_),
    .Q_N(_1795_),
    .Q(\muldiv.regR[15] ));
 sg13g2_dfrbp_1 \muldiv.regR[1]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net159),
    .D(_0011_),
    .Q_N(_1794_),
    .Q(\muldiv.regR[1] ));
 sg13g2_dfrbp_1 \muldiv.regR[2]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net160),
    .D(_0012_),
    .Q_N(_1793_),
    .Q(\muldiv.regR[2] ));
 sg13g2_dfrbp_1 \muldiv.regR[3]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net161),
    .D(_0013_),
    .Q_N(_1792_),
    .Q(\muldiv.regR[3] ));
 sg13g2_dfrbp_1 \muldiv.regR[4]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net162),
    .D(_0014_),
    .Q_N(_1791_),
    .Q(\muldiv.regR[4] ));
 sg13g2_dfrbp_1 \muldiv.regR[5]$_DFFE_PP_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net163),
    .D(_0015_),
    .Q_N(_1790_),
    .Q(\muldiv.regR[5] ));
 sg13g2_dfrbp_1 \muldiv.regR[6]$_DFFE_PP_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net164),
    .D(_0016_),
    .Q_N(_1789_),
    .Q(\muldiv.regR[6] ));
 sg13g2_dfrbp_1 \muldiv.regR[7]$_DFFE_PP_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net165),
    .D(_0017_),
    .Q_N(_1788_),
    .Q(\muldiv.regR[7] ));
 sg13g2_dfrbp_1 \muldiv.regR[8]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net166),
    .D(_0018_),
    .Q_N(_1787_),
    .Q(\muldiv.regR[8] ));
 sg13g2_dfrbp_1 \muldiv.regR[9]$_DFFE_PP_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net167),
    .D(_0019_),
    .Q_N(_1786_),
    .Q(\muldiv.regR[9] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[5]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout19 (.A(_1543_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_1558_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_0741_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1405_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_1298_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0434_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1219_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0428_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1170_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0210_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1143_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0177_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1697_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0143_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1662_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1508_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1371_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1306_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1281_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1223_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1720_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1586_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1367_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1327_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1229_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1131_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1092_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1038_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1709_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1461_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1299_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1014_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0964_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0836_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0306_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1764_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1577_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0408_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0407_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0358_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0227_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0095_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1578_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1355_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1354_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1161_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1128_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1102_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0240_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1687_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1567_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0483_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0346_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0289_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0219_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0178_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0171_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0160_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1774_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1631_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1630_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1617_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1576_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1436_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1434_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1431_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1333_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1311_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1266_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1185_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1155_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1082_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0970_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0644_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1753_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_1632_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_1556_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_1523_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1670_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1433_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_1301_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1265_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_1184_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_1144_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_1124_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_1008_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_0971_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_0951_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_0814_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_0611_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_0601_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_0493_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0460_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0350_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0086_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0053_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_1621_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0986_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0152_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_1501_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_1575_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0042_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_1574_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_1438_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_0925_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_0669_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_0554_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_0494_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_1572_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_1561_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_0020_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_0924_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_1571_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(net134),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_1 fanout134 (.A(net1),
    .X(net134));
 sg13g2_tielo _3603__135 (.L_LO(net135));
 sg13g2_tielo _3604__136 (.L_LO(net136));
 sg13g2_tielo _3605__137 (.L_LO(net137));
 sg13g2_tielo _3606__138 (.L_LO(net138));
 sg13g2_tielo _3609__139 (.L_LO(net139));
 sg13g2_tielo _3610__140 (.L_LO(net140));
 sg13g2_tielo _3611__141 (.L_LO(net141));
 sg13g2_tielo _3612__142 (.L_LO(net142));
 sg13g2_tielo _3613__143 (.L_LO(net143));
 sg13g2_tielo _3614__144 (.L_LO(net144));
 sg13g2_tielo _3615__145 (.L_LO(net145));
 sg13g2_tielo _3617__146 (.L_LO(net146));
 sg13g2_tielo _3618__147 (.L_LO(net147));
 sg13g2_tiehi _3608__149 (.L_HI(net149));
 sg13g2_tiehi \muldiv.div2reg$_SDFF_PN0__150  (.L_HI(net150));
 sg13g2_tiehi \muldiv.negedgeReg_1.area_io_q$_SDFF_NN1__151  (.L_HI(net151));
 sg13g2_tiehi \muldiv.regR[0]$_DFFE_PP__152  (.L_HI(net152));
 sg13g2_tiehi \muldiv.regR[10]$_DFFE_PP__153  (.L_HI(net153));
 sg13g2_tiehi \muldiv.regR[11]$_DFFE_PP__154  (.L_HI(net154));
 sg13g2_tiehi \muldiv.regR[12]$_DFFE_PP__155  (.L_HI(net155));
 sg13g2_tiehi \muldiv.regR[13]$_DFFE_PP__156  (.L_HI(net156));
 sg13g2_tiehi \muldiv.regR[14]$_DFFE_PP__157  (.L_HI(net157));
 sg13g2_tiehi \muldiv.regR[15]$_DFFE_PP__158  (.L_HI(net158));
 sg13g2_tiehi \muldiv.regR[1]$_DFFE_PP__159  (.L_HI(net159));
 sg13g2_tiehi \muldiv.regR[2]$_DFFE_PP__160  (.L_HI(net160));
 sg13g2_tiehi \muldiv.regR[3]$_DFFE_PP__161  (.L_HI(net161));
 sg13g2_tiehi \muldiv.regR[4]$_DFFE_PP__162  (.L_HI(net162));
 sg13g2_tiehi \muldiv.regR[5]$_DFFE_PP__163  (.L_HI(net163));
 sg13g2_tiehi \muldiv.regR[6]$_DFFE_PP__164  (.L_HI(net164));
 sg13g2_tiehi \muldiv.regR[7]$_DFFE_PP__165  (.L_HI(net165));
 sg13g2_tiehi \muldiv.regR[8]$_DFFE_PP__166  (.L_HI(net166));
 sg13g2_tiehi \muldiv.regR[9]$_DFFE_PP__167  (.L_HI(net167));
 sg13g2_buf_1 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_1 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_1 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_1 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_fill_2 FILLER_0_77 ();
 sg13g2_decap_4 FILLER_0_89 ();
 sg13g2_decap_4 FILLER_0_105 ();
 sg13g2_fill_2 FILLER_0_109 ();
 sg13g2_fill_2 FILLER_0_119 ();
 sg13g2_fill_2 FILLER_0_130 ();
 sg13g2_fill_2 FILLER_0_149 ();
 sg13g2_fill_2 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_fill_1 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_185 ();
 sg13g2_fill_1 FILLER_0_192 ();
 sg13g2_fill_2 FILLER_0_208 ();
 sg13g2_decap_4 FILLER_0_214 ();
 sg13g2_fill_1 FILLER_0_218 ();
 sg13g2_fill_2 FILLER_0_223 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_decap_8 FILLER_0_237 ();
 sg13g2_fill_2 FILLER_0_244 ();
 sg13g2_decap_4 FILLER_0_262 ();
 sg13g2_fill_2 FILLER_0_266 ();
 sg13g2_decap_4 FILLER_0_272 ();
 sg13g2_fill_2 FILLER_0_276 ();
 sg13g2_decap_4 FILLER_0_281 ();
 sg13g2_fill_1 FILLER_0_300 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_fill_1 FILLER_0_313 ();
 sg13g2_fill_2 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_4 FILLER_0_343 ();
 sg13g2_fill_1 FILLER_0_347 ();
 sg13g2_fill_1 FILLER_0_352 ();
 sg13g2_fill_2 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_2 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_55 ();
 sg13g2_decap_8 FILLER_1_62 ();
 sg13g2_fill_1 FILLER_1_69 ();
 sg13g2_fill_2 FILLER_1_85 ();
 sg13g2_fill_1 FILLER_1_120 ();
 sg13g2_fill_1 FILLER_1_135 ();
 sg13g2_fill_1 FILLER_1_157 ();
 sg13g2_fill_1 FILLER_1_170 ();
 sg13g2_fill_2 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_fill_1 FILLER_1_189 ();
 sg13g2_fill_1 FILLER_1_196 ();
 sg13g2_fill_2 FILLER_1_207 ();
 sg13g2_fill_1 FILLER_1_238 ();
 sg13g2_fill_2 FILLER_1_263 ();
 sg13g2_fill_1 FILLER_1_265 ();
 sg13g2_fill_1 FILLER_1_275 ();
 sg13g2_fill_1 FILLER_1_284 ();
 sg13g2_fill_1 FILLER_1_305 ();
 sg13g2_fill_2 FILLER_1_314 ();
 sg13g2_decap_4 FILLER_1_336 ();
 sg13g2_fill_2 FILLER_1_340 ();
 sg13g2_fill_2 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_8 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_1_414 ();
 sg13g2_decap_8 FILLER_1_421 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_4 FILLER_2_14 ();
 sg13g2_fill_2 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_27 ();
 sg13g2_decap_8 FILLER_2_34 ();
 sg13g2_decap_4 FILLER_2_41 ();
 sg13g2_fill_2 FILLER_2_59 ();
 sg13g2_fill_2 FILLER_2_65 ();
 sg13g2_fill_1 FILLER_2_67 ();
 sg13g2_fill_1 FILLER_2_73 ();
 sg13g2_fill_2 FILLER_2_79 ();
 sg13g2_fill_1 FILLER_2_81 ();
 sg13g2_fill_2 FILLER_2_95 ();
 sg13g2_fill_1 FILLER_2_108 ();
 sg13g2_fill_1 FILLER_2_114 ();
 sg13g2_fill_2 FILLER_2_119 ();
 sg13g2_fill_1 FILLER_2_125 ();
 sg13g2_fill_2 FILLER_2_130 ();
 sg13g2_fill_1 FILLER_2_145 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_180 ();
 sg13g2_fill_2 FILLER_2_187 ();
 sg13g2_fill_1 FILLER_2_193 ();
 sg13g2_fill_2 FILLER_2_198 ();
 sg13g2_fill_2 FILLER_2_204 ();
 sg13g2_fill_2 FILLER_2_214 ();
 sg13g2_fill_1 FILLER_2_216 ();
 sg13g2_fill_1 FILLER_2_238 ();
 sg13g2_fill_2 FILLER_2_243 ();
 sg13g2_decap_4 FILLER_2_249 ();
 sg13g2_fill_2 FILLER_2_253 ();
 sg13g2_decap_4 FILLER_2_259 ();
 sg13g2_fill_1 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_275 ();
 sg13g2_decap_8 FILLER_2_282 ();
 sg13g2_decap_4 FILLER_2_289 ();
 sg13g2_fill_1 FILLER_2_293 ();
 sg13g2_decap_8 FILLER_2_337 ();
 sg13g2_fill_2 FILLER_2_344 ();
 sg13g2_fill_1 FILLER_2_358 ();
 sg13g2_fill_1 FILLER_2_368 ();
 sg13g2_decap_4 FILLER_2_377 ();
 sg13g2_decap_4 FILLER_2_390 ();
 sg13g2_fill_1 FILLER_2_394 ();
 sg13g2_fill_2 FILLER_2_405 ();
 sg13g2_fill_2 FILLER_2_411 ();
 sg13g2_fill_1 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_14 ();
 sg13g2_fill_2 FILLER_3_20 ();
 sg13g2_fill_1 FILLER_3_22 ();
 sg13g2_decap_4 FILLER_3_31 ();
 sg13g2_fill_2 FILLER_3_35 ();
 sg13g2_fill_1 FILLER_3_52 ();
 sg13g2_fill_2 FILLER_3_57 ();
 sg13g2_fill_2 FILLER_3_64 ();
 sg13g2_fill_2 FILLER_3_70 ();
 sg13g2_fill_1 FILLER_3_72 ();
 sg13g2_fill_2 FILLER_3_80 ();
 sg13g2_decap_8 FILLER_3_87 ();
 sg13g2_decap_4 FILLER_3_94 ();
 sg13g2_decap_4 FILLER_3_103 ();
 sg13g2_fill_2 FILLER_3_107 ();
 sg13g2_fill_1 FILLER_3_136 ();
 sg13g2_fill_1 FILLER_3_142 ();
 sg13g2_fill_1 FILLER_3_148 ();
 sg13g2_fill_2 FILLER_3_154 ();
 sg13g2_fill_2 FILLER_3_164 ();
 sg13g2_fill_1 FILLER_3_166 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_fill_2 FILLER_3_179 ();
 sg13g2_decap_4 FILLER_3_186 ();
 sg13g2_decap_4 FILLER_3_207 ();
 sg13g2_decap_4 FILLER_3_215 ();
 sg13g2_fill_2 FILLER_3_230 ();
 sg13g2_fill_1 FILLER_3_237 ();
 sg13g2_fill_1 FILLER_3_249 ();
 sg13g2_decap_4 FILLER_3_300 ();
 sg13g2_fill_1 FILLER_3_313 ();
 sg13g2_fill_1 FILLER_3_323 ();
 sg13g2_fill_1 FILLER_3_328 ();
 sg13g2_decap_4 FILLER_3_337 ();
 sg13g2_fill_2 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_4 FILLER_3_366 ();
 sg13g2_fill_2 FILLER_3_370 ();
 sg13g2_fill_1 FILLER_3_388 ();
 sg13g2_fill_1 FILLER_3_394 ();
 sg13g2_fill_2 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_fill_2 FILLER_3_419 ();
 sg13g2_fill_1 FILLER_3_421 ();
 sg13g2_decap_4 FILLER_3_426 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_4 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_15 ();
 sg13g2_fill_2 FILLER_4_22 ();
 sg13g2_fill_2 FILLER_4_36 ();
 sg13g2_fill_1 FILLER_4_38 ();
 sg13g2_fill_1 FILLER_4_45 ();
 sg13g2_fill_2 FILLER_4_50 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_fill_1 FILLER_4_86 ();
 sg13g2_fill_1 FILLER_4_96 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_fill_2 FILLER_4_117 ();
 sg13g2_fill_1 FILLER_4_119 ();
 sg13g2_decap_4 FILLER_4_129 ();
 sg13g2_decap_8 FILLER_4_138 ();
 sg13g2_decap_8 FILLER_4_145 ();
 sg13g2_fill_2 FILLER_4_152 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_fill_2 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_205 ();
 sg13g2_decap_8 FILLER_4_212 ();
 sg13g2_decap_4 FILLER_4_219 ();
 sg13g2_fill_1 FILLER_4_223 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_decap_4 FILLER_4_260 ();
 sg13g2_fill_2 FILLER_4_274 ();
 sg13g2_fill_1 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_fill_2 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_293 ();
 sg13g2_decap_8 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_307 ();
 sg13g2_fill_2 FILLER_4_314 ();
 sg13g2_fill_1 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_4 FILLER_4_357 ();
 sg13g2_fill_2 FILLER_4_361 ();
 sg13g2_fill_2 FILLER_4_377 ();
 sg13g2_fill_1 FILLER_4_384 ();
 sg13g2_fill_2 FILLER_4_402 ();
 sg13g2_fill_1 FILLER_4_404 ();
 sg13g2_fill_2 FILLER_4_418 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_4 ();
 sg13g2_decap_4 FILLER_5_15 ();
 sg13g2_decap_4 FILLER_5_23 ();
 sg13g2_fill_1 FILLER_5_32 ();
 sg13g2_fill_1 FILLER_5_53 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_fill_1 FILLER_5_78 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_fill_1 FILLER_5_108 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_125 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_fill_2 FILLER_5_137 ();
 sg13g2_fill_1 FILLER_5_139 ();
 sg13g2_decap_8 FILLER_5_162 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_fill_2 FILLER_5_183 ();
 sg13g2_fill_1 FILLER_5_185 ();
 sg13g2_decap_8 FILLER_5_191 ();
 sg13g2_decap_4 FILLER_5_198 ();
 sg13g2_fill_2 FILLER_5_202 ();
 sg13g2_decap_8 FILLER_5_213 ();
 sg13g2_fill_2 FILLER_5_220 ();
 sg13g2_fill_2 FILLER_5_235 ();
 sg13g2_fill_2 FILLER_5_243 ();
 sg13g2_fill_2 FILLER_5_250 ();
 sg13g2_fill_1 FILLER_5_252 ();
 sg13g2_fill_1 FILLER_5_261 ();
 sg13g2_fill_2 FILLER_5_267 ();
 sg13g2_fill_1 FILLER_5_269 ();
 sg13g2_decap_4 FILLER_5_282 ();
 sg13g2_fill_1 FILLER_5_286 ();
 sg13g2_fill_2 FILLER_5_295 ();
 sg13g2_fill_1 FILLER_5_313 ();
 sg13g2_fill_1 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_fill_1 FILLER_5_346 ();
 sg13g2_decap_4 FILLER_5_354 ();
 sg13g2_fill_2 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_fill_2 FILLER_5_389 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_4 FILLER_5_424 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_7 ();
 sg13g2_decap_4 FILLER_6_19 ();
 sg13g2_decap_8 FILLER_6_27 ();
 sg13g2_fill_1 FILLER_6_34 ();
 sg13g2_fill_1 FILLER_6_40 ();
 sg13g2_fill_1 FILLER_6_49 ();
 sg13g2_fill_1 FILLER_6_59 ();
 sg13g2_decap_8 FILLER_6_66 ();
 sg13g2_fill_2 FILLER_6_73 ();
 sg13g2_fill_1 FILLER_6_75 ();
 sg13g2_fill_2 FILLER_6_91 ();
 sg13g2_fill_1 FILLER_6_106 ();
 sg13g2_fill_1 FILLER_6_137 ();
 sg13g2_fill_2 FILLER_6_162 ();
 sg13g2_fill_1 FILLER_6_164 ();
 sg13g2_fill_2 FILLER_6_219 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_fill_2 FILLER_6_241 ();
 sg13g2_decap_4 FILLER_6_247 ();
 sg13g2_decap_4 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_fill_2 FILLER_6_312 ();
 sg13g2_fill_1 FILLER_6_318 ();
 sg13g2_fill_1 FILLER_6_335 ();
 sg13g2_fill_2 FILLER_6_359 ();
 sg13g2_fill_1 FILLER_6_361 ();
 sg13g2_fill_1 FILLER_6_367 ();
 sg13g2_fill_2 FILLER_6_373 ();
 sg13g2_decap_4 FILLER_6_380 ();
 sg13g2_fill_1 FILLER_6_384 ();
 sg13g2_fill_1 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_7 ();
 sg13g2_fill_2 FILLER_7_26 ();
 sg13g2_fill_1 FILLER_7_32 ();
 sg13g2_fill_2 FILLER_7_40 ();
 sg13g2_fill_1 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_51 ();
 sg13g2_decap_4 FILLER_7_59 ();
 sg13g2_fill_2 FILLER_7_67 ();
 sg13g2_fill_2 FILLER_7_83 ();
 sg13g2_fill_1 FILLER_7_85 ();
 sg13g2_decap_8 FILLER_7_90 ();
 sg13g2_decap_8 FILLER_7_97 ();
 sg13g2_decap_4 FILLER_7_109 ();
 sg13g2_fill_2 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_131 ();
 sg13g2_fill_1 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_148 ();
 sg13g2_decap_8 FILLER_7_155 ();
 sg13g2_decap_8 FILLER_7_162 ();
 sg13g2_decap_4 FILLER_7_169 ();
 sg13g2_fill_2 FILLER_7_173 ();
 sg13g2_decap_4 FILLER_7_180 ();
 sg13g2_decap_4 FILLER_7_193 ();
 sg13g2_fill_2 FILLER_7_206 ();
 sg13g2_fill_1 FILLER_7_208 ();
 sg13g2_decap_4 FILLER_7_226 ();
 sg13g2_decap_4 FILLER_7_237 ();
 sg13g2_fill_2 FILLER_7_241 ();
 sg13g2_decap_4 FILLER_7_247 ();
 sg13g2_fill_2 FILLER_7_251 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_fill_2 FILLER_7_265 ();
 sg13g2_fill_1 FILLER_7_267 ();
 sg13g2_decap_4 FILLER_7_272 ();
 sg13g2_fill_1 FILLER_7_276 ();
 sg13g2_fill_1 FILLER_7_300 ();
 sg13g2_fill_1 FILLER_7_306 ();
 sg13g2_fill_1 FILLER_7_322 ();
 sg13g2_fill_2 FILLER_7_341 ();
 sg13g2_fill_1 FILLER_7_343 ();
 sg13g2_fill_1 FILLER_7_348 ();
 sg13g2_fill_2 FILLER_7_354 ();
 sg13g2_decap_4 FILLER_7_368 ();
 sg13g2_decap_4 FILLER_7_384 ();
 sg13g2_fill_2 FILLER_7_388 ();
 sg13g2_fill_2 FILLER_7_405 ();
 sg13g2_fill_1 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_7_416 ();
 sg13g2_decap_8 FILLER_7_423 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_decap_4 FILLER_8_39 ();
 sg13g2_fill_2 FILLER_8_43 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_fill_1 FILLER_8_67 ();
 sg13g2_fill_1 FILLER_8_91 ();
 sg13g2_decap_4 FILLER_8_96 ();
 sg13g2_decap_4 FILLER_8_108 ();
 sg13g2_fill_1 FILLER_8_112 ();
 sg13g2_decap_4 FILLER_8_121 ();
 sg13g2_fill_2 FILLER_8_125 ();
 sg13g2_fill_1 FILLER_8_153 ();
 sg13g2_fill_2 FILLER_8_158 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_171 ();
 sg13g2_decap_4 FILLER_8_180 ();
 sg13g2_fill_1 FILLER_8_184 ();
 sg13g2_decap_4 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_197 ();
 sg13g2_fill_2 FILLER_8_227 ();
 sg13g2_fill_2 FILLER_8_238 ();
 sg13g2_fill_1 FILLER_8_240 ();
 sg13g2_fill_1 FILLER_8_260 ();
 sg13g2_fill_1 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_275 ();
 sg13g2_decap_8 FILLER_8_282 ();
 sg13g2_fill_1 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_316 ();
 sg13g2_fill_2 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_359 ();
 sg13g2_decap_4 FILLER_8_364 ();
 sg13g2_fill_1 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_fill_2 FILLER_8_389 ();
 sg13g2_fill_1 FILLER_8_391 ();
 sg13g2_fill_1 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_405 ();
 sg13g2_fill_1 FILLER_8_412 ();
 sg13g2_fill_1 FILLER_8_418 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_9 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_21 ();
 sg13g2_fill_1 FILLER_9_23 ();
 sg13g2_fill_2 FILLER_9_54 ();
 sg13g2_fill_1 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_67 ();
 sg13g2_decap_4 FILLER_9_78 ();
 sg13g2_fill_1 FILLER_9_82 ();
 sg13g2_fill_1 FILLER_9_88 ();
 sg13g2_fill_1 FILLER_9_106 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_127 ();
 sg13g2_decap_8 FILLER_9_142 ();
 sg13g2_decap_8 FILLER_9_149 ();
 sg13g2_decap_8 FILLER_9_156 ();
 sg13g2_fill_2 FILLER_9_163 ();
 sg13g2_decap_4 FILLER_9_171 ();
 sg13g2_fill_2 FILLER_9_197 ();
 sg13g2_fill_1 FILLER_9_199 ();
 sg13g2_fill_2 FILLER_9_209 ();
 sg13g2_fill_1 FILLER_9_211 ();
 sg13g2_decap_8 FILLER_9_216 ();
 sg13g2_decap_8 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_230 ();
 sg13g2_decap_4 FILLER_9_239 ();
 sg13g2_fill_1 FILLER_9_243 ();
 sg13g2_decap_4 FILLER_9_248 ();
 sg13g2_fill_2 FILLER_9_256 ();
 sg13g2_fill_1 FILLER_9_258 ();
 sg13g2_fill_2 FILLER_9_264 ();
 sg13g2_fill_1 FILLER_9_266 ();
 sg13g2_fill_2 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_310 ();
 sg13g2_decap_4 FILLER_9_317 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_fill_2 FILLER_9_327 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_fill_1 FILLER_9_339 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_4 FILLER_9_382 ();
 sg13g2_fill_2 FILLER_9_386 ();
 sg13g2_fill_2 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_402 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_412 ();
 sg13g2_fill_1 FILLER_9_419 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_23 ();
 sg13g2_decap_8 FILLER_10_30 ();
 sg13g2_decap_8 FILLER_10_37 ();
 sg13g2_decap_8 FILLER_10_44 ();
 sg13g2_decap_4 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_55 ();
 sg13g2_fill_2 FILLER_10_65 ();
 sg13g2_fill_1 FILLER_10_67 ();
 sg13g2_fill_1 FILLER_10_73 ();
 sg13g2_fill_1 FILLER_10_80 ();
 sg13g2_decap_8 FILLER_10_85 ();
 sg13g2_decap_4 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_100 ();
 sg13g2_decap_4 FILLER_10_143 ();
 sg13g2_fill_1 FILLER_10_151 ();
 sg13g2_decap_4 FILLER_10_157 ();
 sg13g2_decap_4 FILLER_10_168 ();
 sg13g2_fill_1 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_197 ();
 sg13g2_decap_4 FILLER_10_204 ();
 sg13g2_fill_2 FILLER_10_208 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_fill_2 FILLER_10_226 ();
 sg13g2_fill_1 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_250 ();
 sg13g2_fill_2 FILLER_10_260 ();
 sg13g2_fill_1 FILLER_10_262 ();
 sg13g2_decap_8 FILLER_10_276 ();
 sg13g2_fill_1 FILLER_10_292 ();
 sg13g2_fill_2 FILLER_10_325 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_decap_4 FILLER_10_343 ();
 sg13g2_decap_4 FILLER_10_352 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_4 FILLER_10_379 ();
 sg13g2_fill_2 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_fill_1 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_11 ();
 sg13g2_fill_1 FILLER_11_18 ();
 sg13g2_fill_2 FILLER_11_27 ();
 sg13g2_fill_2 FILLER_11_33 ();
 sg13g2_decap_4 FILLER_11_40 ();
 sg13g2_decap_4 FILLER_11_52 ();
 sg13g2_fill_2 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_66 ();
 sg13g2_fill_2 FILLER_11_80 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_fill_1 FILLER_11_87 ();
 sg13g2_fill_2 FILLER_11_93 ();
 sg13g2_fill_2 FILLER_11_113 ();
 sg13g2_fill_2 FILLER_11_130 ();
 sg13g2_fill_1 FILLER_11_132 ();
 sg13g2_decap_8 FILLER_11_145 ();
 sg13g2_fill_2 FILLER_11_152 ();
 sg13g2_fill_1 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_201 ();
 sg13g2_decap_4 FILLER_11_208 ();
 sg13g2_fill_2 FILLER_11_212 ();
 sg13g2_decap_4 FILLER_11_218 ();
 sg13g2_fill_1 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_257 ();
 sg13g2_fill_1 FILLER_11_263 ();
 sg13g2_fill_1 FILLER_11_269 ();
 sg13g2_fill_1 FILLER_11_284 ();
 sg13g2_fill_2 FILLER_11_290 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_fill_1 FILLER_11_311 ();
 sg13g2_fill_1 FILLER_11_320 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_fill_1 FILLER_11_345 ();
 sg13g2_decap_8 FILLER_11_352 ();
 sg13g2_decap_4 FILLER_11_367 ();
 sg13g2_fill_2 FILLER_11_371 ();
 sg13g2_fill_1 FILLER_11_380 ();
 sg13g2_fill_2 FILLER_11_397 ();
 sg13g2_decap_8 FILLER_11_404 ();
 sg13g2_fill_2 FILLER_11_411 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_2 FILLER_12_28 ();
 sg13g2_fill_2 FILLER_12_35 ();
 sg13g2_fill_2 FILLER_12_44 ();
 sg13g2_fill_1 FILLER_12_46 ();
 sg13g2_fill_2 FILLER_12_55 ();
 sg13g2_fill_1 FILLER_12_57 ();
 sg13g2_fill_2 FILLER_12_62 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_fill_2 FILLER_12_91 ();
 sg13g2_fill_1 FILLER_12_113 ();
 sg13g2_decap_8 FILLER_12_139 ();
 sg13g2_decap_8 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_173 ();
 sg13g2_fill_1 FILLER_12_180 ();
 sg13g2_fill_1 FILLER_12_186 ();
 sg13g2_fill_1 FILLER_12_192 ();
 sg13g2_decap_4 FILLER_12_202 ();
 sg13g2_fill_1 FILLER_12_212 ();
 sg13g2_fill_2 FILLER_12_221 ();
 sg13g2_fill_1 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_243 ();
 sg13g2_decap_4 FILLER_12_265 ();
 sg13g2_fill_2 FILLER_12_269 ();
 sg13g2_fill_1 FILLER_12_291 ();
 sg13g2_fill_1 FILLER_12_301 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_fill_1 FILLER_12_319 ();
 sg13g2_fill_2 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_336 ();
 sg13g2_fill_1 FILLER_12_338 ();
 sg13g2_fill_2 FILLER_12_359 ();
 sg13g2_fill_1 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_4 FILLER_12_382 ();
 sg13g2_decap_4 FILLER_12_398 ();
 sg13g2_decap_8 FILLER_12_409 ();
 sg13g2_decap_4 FILLER_12_424 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_15 ();
 sg13g2_fill_2 FILLER_13_31 ();
 sg13g2_decap_8 FILLER_13_57 ();
 sg13g2_decap_8 FILLER_13_64 ();
 sg13g2_fill_2 FILLER_13_71 ();
 sg13g2_fill_1 FILLER_13_73 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_fill_1 FILLER_13_97 ();
 sg13g2_fill_1 FILLER_13_103 ();
 sg13g2_fill_2 FILLER_13_109 ();
 sg13g2_fill_2 FILLER_13_115 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_1 FILLER_13_128 ();
 sg13g2_decap_4 FILLER_13_144 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_fill_1 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_205 ();
 sg13g2_decap_8 FILLER_13_212 ();
 sg13g2_decap_8 FILLER_13_219 ();
 sg13g2_fill_2 FILLER_13_226 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_decap_4 FILLER_13_248 ();
 sg13g2_fill_1 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_257 ();
 sg13g2_decap_8 FILLER_13_264 ();
 sg13g2_decap_8 FILLER_13_271 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_decap_8 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_299 ();
 sg13g2_decap_8 FILLER_13_306 ();
 sg13g2_decap_8 FILLER_13_313 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_2 FILLER_13_325 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_decap_4 FILLER_13_354 ();
 sg13g2_fill_2 FILLER_13_358 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_fill_2 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_fill_1 FILLER_13_392 ();
 sg13g2_fill_2 FILLER_13_403 ();
 sg13g2_fill_1 FILLER_13_419 ();
 sg13g2_decap_4 FILLER_13_425 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_9 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_18 ();
 sg13g2_fill_1 FILLER_14_24 ();
 sg13g2_fill_2 FILLER_14_37 ();
 sg13g2_fill_1 FILLER_14_44 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_64 ();
 sg13g2_fill_2 FILLER_14_77 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_fill_2 FILLER_14_88 ();
 sg13g2_fill_1 FILLER_14_90 ();
 sg13g2_fill_1 FILLER_14_95 ();
 sg13g2_fill_1 FILLER_14_99 ();
 sg13g2_fill_2 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_109 ();
 sg13g2_decap_4 FILLER_14_114 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_decap_4 FILLER_14_145 ();
 sg13g2_fill_1 FILLER_14_149 ();
 sg13g2_fill_2 FILLER_14_154 ();
 sg13g2_fill_1 FILLER_14_156 ();
 sg13g2_decap_4 FILLER_14_185 ();
 sg13g2_fill_2 FILLER_14_189 ();
 sg13g2_fill_2 FILLER_14_204 ();
 sg13g2_fill_2 FILLER_14_224 ();
 sg13g2_fill_1 FILLER_14_226 ();
 sg13g2_decap_4 FILLER_14_236 ();
 sg13g2_fill_2 FILLER_14_253 ();
 sg13g2_fill_1 FILLER_14_255 ();
 sg13g2_decap_4 FILLER_14_292 ();
 sg13g2_fill_2 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_4 FILLER_14_315 ();
 sg13g2_decap_4 FILLER_14_323 ();
 sg13g2_fill_2 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_4 FILLER_14_361 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_decap_4 FILLER_14_397 ();
 sg13g2_fill_1 FILLER_14_416 ();
 sg13g2_decap_4 FILLER_14_425 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_14 ();
 sg13g2_fill_2 FILLER_15_35 ();
 sg13g2_fill_1 FILLER_15_37 ();
 sg13g2_decap_4 FILLER_15_42 ();
 sg13g2_fill_1 FILLER_15_69 ();
 sg13g2_fill_1 FILLER_15_77 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_fill_2 FILLER_15_101 ();
 sg13g2_decap_4 FILLER_15_125 ();
 sg13g2_fill_2 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_158 ();
 sg13g2_fill_1 FILLER_15_160 ();
 sg13g2_fill_1 FILLER_15_169 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_decap_8 FILLER_15_180 ();
 sg13g2_fill_1 FILLER_15_187 ();
 sg13g2_fill_1 FILLER_15_192 ();
 sg13g2_fill_1 FILLER_15_212 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_decap_4 FILLER_15_232 ();
 sg13g2_fill_1 FILLER_15_236 ();
 sg13g2_fill_2 FILLER_15_249 ();
 sg13g2_decap_4 FILLER_15_263 ();
 sg13g2_fill_2 FILLER_15_267 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_281 ();
 sg13g2_fill_2 FILLER_15_286 ();
 sg13g2_fill_1 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_299 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_decap_4 FILLER_15_351 ();
 sg13g2_fill_2 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_fill_2 FILLER_15_397 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_4 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_2 FILLER_16_23 ();
 sg13g2_fill_1 FILLER_16_25 ();
 sg13g2_fill_2 FILLER_16_44 ();
 sg13g2_fill_1 FILLER_16_46 ();
 sg13g2_fill_2 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_64 ();
 sg13g2_fill_2 FILLER_16_98 ();
 sg13g2_fill_1 FILLER_16_100 ();
 sg13g2_decap_4 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_fill_1 FILLER_16_125 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_fill_2 FILLER_16_165 ();
 sg13g2_fill_1 FILLER_16_167 ();
 sg13g2_fill_2 FILLER_16_181 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_fill_2 FILLER_16_202 ();
 sg13g2_fill_1 FILLER_16_204 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_fill_1 FILLER_16_244 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_fill_1 FILLER_16_258 ();
 sg13g2_fill_2 FILLER_16_280 ();
 sg13g2_fill_1 FILLER_16_282 ();
 sg13g2_decap_4 FILLER_16_288 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_2 FILLER_16_311 ();
 sg13g2_fill_1 FILLER_16_313 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_fill_1 FILLER_16_344 ();
 sg13g2_fill_2 FILLER_16_350 ();
 sg13g2_fill_2 FILLER_16_371 ();
 sg13g2_fill_1 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_1 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_418 ();
 sg13g2_decap_4 FILLER_16_425 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_19 ();
 sg13g2_decap_4 FILLER_17_71 ();
 sg13g2_fill_2 FILLER_17_75 ();
 sg13g2_decap_8 FILLER_17_82 ();
 sg13g2_decap_4 FILLER_17_89 ();
 sg13g2_fill_1 FILLER_17_101 ();
 sg13g2_fill_2 FILLER_17_107 ();
 sg13g2_decap_4 FILLER_17_129 ();
 sg13g2_fill_2 FILLER_17_133 ();
 sg13g2_decap_4 FILLER_17_163 ();
 sg13g2_decap_4 FILLER_17_172 ();
 sg13g2_fill_2 FILLER_17_176 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_fill_1 FILLER_17_184 ();
 sg13g2_decap_8 FILLER_17_190 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_decap_4 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_fill_2 FILLER_17_265 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_fill_1 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_283 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_316 ();
 sg13g2_fill_2 FILLER_17_328 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_4 FILLER_17_351 ();
 sg13g2_fill_1 FILLER_17_355 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_4 FILLER_17_379 ();
 sg13g2_fill_1 FILLER_17_383 ();
 sg13g2_fill_2 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_416 ();
 sg13g2_decap_8 FILLER_17_422 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_27 ();
 sg13g2_decap_8 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_71 ();
 sg13g2_decap_4 FILLER_18_78 ();
 sg13g2_decap_8 FILLER_18_87 ();
 sg13g2_decap_8 FILLER_18_94 ();
 sg13g2_decap_4 FILLER_18_101 ();
 sg13g2_fill_2 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_111 ();
 sg13g2_decap_8 FILLER_18_118 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_148 ();
 sg13g2_fill_1 FILLER_18_155 ();
 sg13g2_decap_4 FILLER_18_170 ();
 sg13g2_decap_8 FILLER_18_188 ();
 sg13g2_fill_1 FILLER_18_195 ();
 sg13g2_fill_1 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_222 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_232 ();
 sg13g2_decap_4 FILLER_18_239 ();
 sg13g2_fill_2 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_260 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_4 FILLER_18_273 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_332 ();
 sg13g2_fill_1 FILLER_18_337 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_fill_2 FILLER_18_375 ();
 sg13g2_fill_2 FILLER_18_381 ();
 sg13g2_fill_1 FILLER_18_387 ();
 sg13g2_fill_1 FILLER_18_411 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_decap_4 FILLER_18_424 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_17 ();
 sg13g2_fill_1 FILLER_19_43 ();
 sg13g2_fill_2 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_63 ();
 sg13g2_fill_2 FILLER_19_76 ();
 sg13g2_fill_1 FILLER_19_83 ();
 sg13g2_decap_4 FILLER_19_88 ();
 sg13g2_fill_1 FILLER_19_92 ();
 sg13g2_decap_4 FILLER_19_97 ();
 sg13g2_fill_2 FILLER_19_101 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_decap_4 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_192 ();
 sg13g2_fill_1 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_210 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_224 ();
 sg13g2_fill_2 FILLER_19_230 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_fill_1 FILLER_19_308 ();
 sg13g2_decap_4 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_fill_2 FILLER_19_327 ();
 sg13g2_fill_1 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_334 ();
 sg13g2_fill_2 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_348 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_389 ();
 sg13g2_decap_4 FILLER_19_408 ();
 sg13g2_fill_2 FILLER_19_412 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_14 ();
 sg13g2_decap_4 FILLER_20_29 ();
 sg13g2_fill_1 FILLER_20_41 ();
 sg13g2_fill_1 FILLER_20_59 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_4 FILLER_20_81 ();
 sg13g2_fill_1 FILLER_20_85 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_fill_1 FILLER_20_127 ();
 sg13g2_decap_4 FILLER_20_146 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_decap_4 FILLER_20_164 ();
 sg13g2_fill_2 FILLER_20_168 ();
 sg13g2_fill_2 FILLER_20_192 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_1 FILLER_20_244 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_decap_4 FILLER_20_255 ();
 sg13g2_decap_4 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_270 ();
 sg13g2_fill_2 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_296 ();
 sg13g2_fill_1 FILLER_20_312 ();
 sg13g2_decap_4 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_decap_4 FILLER_20_366 ();
 sg13g2_fill_1 FILLER_20_370 ();
 sg13g2_fill_1 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_4 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_418 ();
 sg13g2_decap_4 FILLER_20_425 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_16 ();
 sg13g2_fill_1 FILLER_21_31 ();
 sg13g2_fill_2 FILLER_21_53 ();
 sg13g2_fill_2 FILLER_21_59 ();
 sg13g2_fill_1 FILLER_21_61 ();
 sg13g2_fill_1 FILLER_21_72 ();
 sg13g2_fill_2 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_decap_4 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_122 ();
 sg13g2_fill_2 FILLER_21_128 ();
 sg13g2_fill_1 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_146 ();
 sg13g2_decap_8 FILLER_21_153 ();
 sg13g2_fill_1 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_206 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_decap_4 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_2 FILLER_21_246 ();
 sg13g2_fill_1 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_287 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_1 FILLER_21_298 ();
 sg13g2_fill_1 FILLER_21_304 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_4 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_fill_2 FILLER_21_346 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_fill_2 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_19 ();
 sg13g2_fill_1 FILLER_22_21 ();
 sg13g2_decap_4 FILLER_22_31 ();
 sg13g2_fill_1 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_59 ();
 sg13g2_decap_8 FILLER_22_66 ();
 sg13g2_decap_8 FILLER_22_73 ();
 sg13g2_fill_2 FILLER_22_80 ();
 sg13g2_fill_1 FILLER_22_102 ();
 sg13g2_fill_2 FILLER_22_118 ();
 sg13g2_fill_2 FILLER_22_125 ();
 sg13g2_fill_1 FILLER_22_132 ();
 sg13g2_fill_1 FILLER_22_138 ();
 sg13g2_decap_8 FILLER_22_143 ();
 sg13g2_decap_8 FILLER_22_150 ();
 sg13g2_decap_8 FILLER_22_157 ();
 sg13g2_fill_2 FILLER_22_164 ();
 sg13g2_fill_1 FILLER_22_166 ();
 sg13g2_decap_4 FILLER_22_204 ();
 sg13g2_fill_2 FILLER_22_208 ();
 sg13g2_decap_4 FILLER_22_219 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_fill_1 FILLER_22_236 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_4 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_fill_1 FILLER_22_328 ();
 sg13g2_fill_1 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_339 ();
 sg13g2_fill_2 FILLER_22_346 ();
 sg13g2_decap_4 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_35 ();
 sg13g2_fill_1 FILLER_23_44 ();
 sg13g2_fill_2 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_71 ();
 sg13g2_fill_1 FILLER_23_78 ();
 sg13g2_fill_2 FILLER_23_93 ();
 sg13g2_fill_1 FILLER_23_99 ();
 sg13g2_fill_2 FILLER_23_107 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_fill_1 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_128 ();
 sg13g2_fill_1 FILLER_23_139 ();
 sg13g2_fill_1 FILLER_23_149 ();
 sg13g2_decap_8 FILLER_23_163 ();
 sg13g2_fill_2 FILLER_23_170 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_fill_1 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_201 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_decap_8 FILLER_23_251 ();
 sg13g2_fill_1 FILLER_23_263 ();
 sg13g2_decap_4 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_280 ();
 sg13g2_fill_1 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_296 ();
 sg13g2_decap_8 FILLER_23_303 ();
 sg13g2_fill_2 FILLER_23_326 ();
 sg13g2_fill_1 FILLER_23_328 ();
 sg13g2_decap_4 FILLER_23_387 ();
 sg13g2_fill_1 FILLER_23_391 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_fill_2 FILLER_24_32 ();
 sg13g2_decap_4 FILLER_24_46 ();
 sg13g2_fill_2 FILLER_24_58 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_71 ();
 sg13g2_fill_2 FILLER_24_78 ();
 sg13g2_decap_8 FILLER_24_101 ();
 sg13g2_fill_2 FILLER_24_118 ();
 sg13g2_decap_8 FILLER_24_139 ();
 sg13g2_fill_2 FILLER_24_146 ();
 sg13g2_decap_8 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_160 ();
 sg13g2_decap_8 FILLER_24_167 ();
 sg13g2_fill_2 FILLER_24_174 ();
 sg13g2_decap_8 FILLER_24_190 ();
 sg13g2_fill_2 FILLER_24_197 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_4 FILLER_24_236 ();
 sg13g2_fill_2 FILLER_24_240 ();
 sg13g2_decap_4 FILLER_24_258 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_278 ();
 sg13g2_fill_2 FILLER_24_283 ();
 sg13g2_decap_8 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_295 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_decap_8 FILLER_24_306 ();
 sg13g2_fill_2 FILLER_24_313 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_331 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_fill_2 FILLER_24_396 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_decap_4 FILLER_25_31 ();
 sg13g2_fill_2 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_76 ();
 sg13g2_fill_1 FILLER_25_88 ();
 sg13g2_fill_1 FILLER_25_94 ();
 sg13g2_fill_1 FILLER_25_112 ();
 sg13g2_fill_2 FILLER_25_117 ();
 sg13g2_decap_4 FILLER_25_123 ();
 sg13g2_decap_4 FILLER_25_135 ();
 sg13g2_decap_4 FILLER_25_144 ();
 sg13g2_fill_2 FILLER_25_148 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_4 FILLER_25_169 ();
 sg13g2_decap_8 FILLER_25_194 ();
 sg13g2_fill_2 FILLER_25_201 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_226 ();
 sg13g2_decap_8 FILLER_25_233 ();
 sg13g2_decap_4 FILLER_25_240 ();
 sg13g2_fill_1 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_decap_4 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_329 ();
 sg13g2_fill_2 FILLER_25_358 ();
 sg13g2_fill_2 FILLER_25_364 ();
 sg13g2_fill_1 FILLER_25_366 ();
 sg13g2_fill_2 FILLER_25_372 ();
 sg13g2_fill_1 FILLER_25_374 ();
 sg13g2_fill_2 FILLER_25_380 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_2 FILLER_25_412 ();
 sg13g2_fill_1 FILLER_25_414 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_27 ();
 sg13g2_fill_2 FILLER_26_33 ();
 sg13g2_fill_1 FILLER_26_35 ();
 sg13g2_fill_1 FILLER_26_40 ();
 sg13g2_fill_2 FILLER_26_51 ();
 sg13g2_decap_8 FILLER_26_71 ();
 sg13g2_fill_1 FILLER_26_78 ();
 sg13g2_fill_1 FILLER_26_85 ();
 sg13g2_decap_4 FILLER_26_91 ();
 sg13g2_fill_2 FILLER_26_122 ();
 sg13g2_fill_1 FILLER_26_124 ();
 sg13g2_fill_2 FILLER_26_129 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_4 FILLER_26_144 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_decap_4 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_233 ();
 sg13g2_fill_1 FILLER_26_240 ();
 sg13g2_decap_4 FILLER_26_254 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_decap_4 FILLER_26_281 ();
 sg13g2_decap_8 FILLER_26_299 ();
 sg13g2_decap_4 FILLER_26_306 ();
 sg13g2_fill_2 FILLER_26_323 ();
 sg13g2_fill_1 FILLER_26_325 ();
 sg13g2_decap_4 FILLER_26_330 ();
 sg13g2_fill_2 FILLER_26_334 ();
 sg13g2_decap_4 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_348 ();
 sg13g2_fill_1 FILLER_26_355 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_4 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_1 FILLER_26_407 ();
 sg13g2_decap_4 FILLER_26_426 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_33 ();
 sg13g2_decap_8 FILLER_27_40 ();
 sg13g2_fill_2 FILLER_27_47 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_54 ();
 sg13g2_fill_1 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_62 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_fill_1 FILLER_27_85 ();
 sg13g2_fill_2 FILLER_27_93 ();
 sg13g2_decap_8 FILLER_27_103 ();
 sg13g2_fill_2 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_116 ();
 sg13g2_decap_4 FILLER_27_138 ();
 sg13g2_decap_8 FILLER_27_146 ();
 sg13g2_fill_2 FILLER_27_153 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_decap_8 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_decap_4 FILLER_27_176 ();
 sg13g2_decap_4 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_195 ();
 sg13g2_decap_8 FILLER_27_202 ();
 sg13g2_fill_2 FILLER_27_209 ();
 sg13g2_fill_2 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_235 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_fill_1 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_258 ();
 sg13g2_decap_4 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_269 ();
 sg13g2_fill_1 FILLER_27_276 ();
 sg13g2_fill_2 FILLER_27_281 ();
 sg13g2_decap_8 FILLER_27_290 ();
 sg13g2_fill_2 FILLER_27_297 ();
 sg13g2_fill_2 FILLER_27_323 ();
 sg13g2_fill_2 FILLER_27_333 ();
 sg13g2_decap_4 FILLER_27_345 ();
 sg13g2_fill_2 FILLER_27_349 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_fill_2 FILLER_27_385 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_24 ();
 sg13g2_fill_2 FILLER_28_34 ();
 sg13g2_fill_1 FILLER_28_36 ();
 sg13g2_decap_4 FILLER_28_57 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_101 ();
 sg13g2_decap_8 FILLER_28_107 ();
 sg13g2_fill_2 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_fill_1 FILLER_28_225 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_281 ();
 sg13g2_decap_8 FILLER_28_304 ();
 sg13g2_decap_4 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_fill_2 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_2 FILLER_28_392 ();
 sg13g2_fill_1 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_23 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_decap_4 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_72 ();
 sg13g2_decap_4 FILLER_29_79 ();
 sg13g2_fill_2 FILLER_29_109 ();
 sg13g2_decap_4 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_123 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_fill_2 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_152 ();
 sg13g2_decap_4 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_170 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_217 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_241 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_decap_8 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_260 ();
 sg13g2_decap_8 FILLER_29_267 ();
 sg13g2_decap_4 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_286 ();
 sg13g2_fill_2 FILLER_29_293 ();
 sg13g2_decap_4 FILLER_29_309 ();
 sg13g2_fill_2 FILLER_29_313 ();
 sg13g2_decap_4 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_328 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_1 FILLER_29_344 ();
 sg13g2_decap_4 FILLER_29_357 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_366 ();
 sg13g2_decap_8 FILLER_29_373 ();
 sg13g2_fill_2 FILLER_29_380 ();
 sg13g2_fill_2 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_409 ();
 sg13g2_fill_2 FILLER_29_415 ();
 sg13g2_fill_1 FILLER_29_417 ();
 sg13g2_decap_4 FILLER_29_425 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_decap_8 FILLER_30_30 ();
 sg13g2_decap_4 FILLER_30_62 ();
 sg13g2_fill_2 FILLER_30_71 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_1 FILLER_30_87 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_109 ();
 sg13g2_fill_1 FILLER_30_118 ();
 sg13g2_fill_1 FILLER_30_127 ();
 sg13g2_decap_4 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_137 ();
 sg13g2_fill_2 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_2 FILLER_30_207 ();
 sg13g2_fill_2 FILLER_30_214 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_decap_8 FILLER_30_248 ();
 sg13g2_fill_1 FILLER_30_255 ();
 sg13g2_decap_8 FILLER_30_269 ();
 sg13g2_decap_4 FILLER_30_276 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_decap_8 FILLER_30_292 ();
 sg13g2_decap_8 FILLER_30_299 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_2 FILLER_30_339 ();
 sg13g2_fill_1 FILLER_30_341 ();
 sg13g2_decap_4 FILLER_30_347 ();
 sg13g2_fill_2 FILLER_30_351 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_384 ();
 sg13g2_fill_2 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_17 ();
 sg13g2_decap_8 FILLER_31_24 ();
 sg13g2_decap_4 FILLER_31_31 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_51 ();
 sg13g2_fill_2 FILLER_31_58 ();
 sg13g2_decap_8 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_96 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_fill_2 FILLER_31_111 ();
 sg13g2_fill_1 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_119 ();
 sg13g2_fill_2 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_126 ();
 sg13g2_decap_4 FILLER_31_131 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_151 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_172 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_decap_4 FILLER_31_212 ();
 sg13g2_fill_2 FILLER_31_216 ();
 sg13g2_fill_2 FILLER_31_230 ();
 sg13g2_decap_4 FILLER_31_261 ();
 sg13g2_fill_1 FILLER_31_285 ();
 sg13g2_decap_8 FILLER_31_290 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_fill_2 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_decap_4 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_328 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_377 ();
 sg13g2_fill_1 FILLER_31_384 ();
 sg13g2_decap_4 FILLER_31_395 ();
 sg13g2_fill_1 FILLER_31_399 ();
 sg13g2_decap_4 FILLER_31_426 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_17 ();
 sg13g2_fill_1 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_57 ();
 sg13g2_decap_4 FILLER_32_72 ();
 sg13g2_fill_2 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_86 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_121 ();
 sg13g2_decap_4 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_2 FILLER_32_139 ();
 sg13g2_decap_8 FILLER_32_146 ();
 sg13g2_decap_8 FILLER_32_153 ();
 sg13g2_decap_4 FILLER_32_160 ();
 sg13g2_fill_2 FILLER_32_164 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_4 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_decap_4 FILLER_32_253 ();
 sg13g2_decap_4 FILLER_32_263 ();
 sg13g2_fill_1 FILLER_32_275 ();
 sg13g2_decap_4 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_284 ();
 sg13g2_fill_2 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_fill_2 FILLER_32_318 ();
 sg13g2_decap_8 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_331 ();
 sg13g2_fill_2 FILLER_32_355 ();
 sg13g2_fill_2 FILLER_32_369 ();
 sg13g2_fill_2 FILLER_32_377 ();
 sg13g2_fill_1 FILLER_32_379 ();
 sg13g2_fill_2 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_403 ();
 sg13g2_fill_2 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_32_414 ();
 sg13g2_decap_8 FILLER_32_421 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_16 ();
 sg13g2_fill_1 FILLER_33_48 ();
 sg13g2_fill_2 FILLER_33_54 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_74 ();
 sg13g2_fill_2 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_83 ();
 sg13g2_fill_2 FILLER_33_93 ();
 sg13g2_decap_4 FILLER_33_114 ();
 sg13g2_decap_4 FILLER_33_130 ();
 sg13g2_decap_8 FILLER_33_138 ();
 sg13g2_decap_4 FILLER_33_145 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_decap_4 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_decap_8 FILLER_33_187 ();
 sg13g2_decap_8 FILLER_33_194 ();
 sg13g2_decap_8 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_decap_8 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_254 ();
 sg13g2_decap_4 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_291 ();
 sg13g2_decap_8 FILLER_33_297 ();
 sg13g2_decap_8 FILLER_33_304 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_decap_8 FILLER_33_376 ();
 sg13g2_decap_4 FILLER_33_383 ();
 sg13g2_fill_2 FILLER_33_387 ();
 sg13g2_decap_4 FILLER_33_399 ();
 sg13g2_fill_1 FILLER_33_403 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_12 ();
 sg13g2_fill_2 FILLER_34_26 ();
 sg13g2_fill_1 FILLER_34_37 ();
 sg13g2_fill_1 FILLER_34_45 ();
 sg13g2_fill_2 FILLER_34_51 ();
 sg13g2_fill_2 FILLER_34_57 ();
 sg13g2_fill_2 FILLER_34_65 ();
 sg13g2_decap_8 FILLER_34_72 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_90 ();
 sg13g2_fill_1 FILLER_34_92 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_fill_1 FILLER_34_100 ();
 sg13g2_fill_1 FILLER_34_114 ();
 sg13g2_decap_8 FILLER_34_129 ();
 sg13g2_decap_4 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_decap_8 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_fill_2 FILLER_34_219 ();
 sg13g2_fill_2 FILLER_34_225 ();
 sg13g2_decap_4 FILLER_34_255 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_300 ();
 sg13g2_decap_8 FILLER_34_318 ();
 sg13g2_decap_8 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_decap_4 FILLER_34_425 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_8 ();
 sg13g2_fill_1 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_23 ();
 sg13g2_fill_1 FILLER_35_30 ();
 sg13g2_fill_2 FILLER_35_36 ();
 sg13g2_fill_1 FILLER_35_38 ();
 sg13g2_fill_2 FILLER_35_45 ();
 sg13g2_fill_1 FILLER_35_47 ();
 sg13g2_fill_2 FILLER_35_54 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_fill_1 FILLER_35_104 ();
 sg13g2_fill_1 FILLER_35_109 ();
 sg13g2_decap_8 FILLER_35_114 ();
 sg13g2_decap_4 FILLER_35_121 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_187 ();
 sg13g2_decap_4 FILLER_35_193 ();
 sg13g2_decap_8 FILLER_35_230 ();
 sg13g2_decap_4 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_241 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_decap_4 FILLER_35_289 ();
 sg13g2_fill_1 FILLER_35_293 ();
 sg13g2_decap_8 FILLER_35_298 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_fill_1 FILLER_35_343 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_2 FILLER_35_378 ();
 sg13g2_fill_2 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_9 ();
 sg13g2_fill_2 FILLER_36_30 ();
 sg13g2_decap_4 FILLER_36_79 ();
 sg13g2_fill_2 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_109 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_149 ();
 sg13g2_decap_4 FILLER_36_155 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_decap_4 FILLER_36_173 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_fill_2 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_4 FILLER_36_225 ();
 sg13g2_fill_2 FILLER_36_229 ();
 sg13g2_decap_8 FILLER_36_236 ();
 sg13g2_decap_4 FILLER_36_243 ();
 sg13g2_fill_2 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_2 FILLER_36_288 ();
 sg13g2_decap_8 FILLER_36_297 ();
 sg13g2_decap_8 FILLER_36_304 ();
 sg13g2_decap_8 FILLER_36_311 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_decap_4 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_374 ();
 sg13g2_fill_2 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_30 ();
 sg13g2_fill_2 FILLER_37_35 ();
 sg13g2_fill_1 FILLER_37_37 ();
 sg13g2_fill_2 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_44 ();
 sg13g2_decap_4 FILLER_37_50 ();
 sg13g2_fill_2 FILLER_37_54 ();
 sg13g2_fill_1 FILLER_37_85 ();
 sg13g2_decap_4 FILLER_37_93 ();
 sg13g2_fill_1 FILLER_37_97 ();
 sg13g2_decap_4 FILLER_37_106 ();
 sg13g2_fill_2 FILLER_37_110 ();
 sg13g2_fill_2 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_118 ();
 sg13g2_decap_8 FILLER_37_124 ();
 sg13g2_fill_2 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_148 ();
 sg13g2_decap_8 FILLER_37_155 ();
 sg13g2_decap_8 FILLER_37_162 ();
 sg13g2_fill_2 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_171 ();
 sg13g2_decap_4 FILLER_37_191 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_decap_4 FILLER_37_237 ();
 sg13g2_fill_2 FILLER_37_241 ();
 sg13g2_fill_1 FILLER_37_253 ();
 sg13g2_fill_2 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_296 ();
 sg13g2_decap_8 FILLER_37_302 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_366 ();
 sg13g2_fill_1 FILLER_37_368 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_78 ();
 sg13g2_fill_2 FILLER_38_82 ();
 sg13g2_fill_1 FILLER_38_113 ();
 sg13g2_decap_4 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_4 FILLER_38_208 ();
 sg13g2_decap_4 FILLER_38_225 ();
 sg13g2_decap_8 FILLER_38_237 ();
 sg13g2_decap_4 FILLER_38_256 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_314 ();
 sg13g2_decap_8 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_1 FILLER_38_423 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
