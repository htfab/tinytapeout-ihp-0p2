module tt_um_ravenslofty_chess (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire clknet_leaf_0_clk;
 wire net313;
 wire \b.gen_square[0].sq.color ;
 wire \b.gen_square[0].sq.mask ;
 wire \b.gen_square[0].sq.piece[0] ;
 wire \b.gen_square[0].sq.piece[1] ;
 wire \b.gen_square[0].sq.piece[2] ;
 wire \b.gen_square[0].sq.state_mode[0] ;
 wire \b.gen_square[0].sq.state_mode[1] ;
 wire \b.gen_square[0].sq.state_mode[2] ;
 wire \b.gen_square[0].sq.write_bus[0] ;
 wire \b.gen_square[0].sq.write_bus[1] ;
 wire \b.gen_square[0].sq.write_bus[2] ;
 wire \b.gen_square[0].sq.write_bus[3] ;
 wire \b.gen_square[0].sq.wtm ;
 wire \b.gen_square[10].sq.color ;
 wire \b.gen_square[10].sq.mask ;
 wire \b.gen_square[10].sq.piece[0] ;
 wire \b.gen_square[10].sq.piece[1] ;
 wire \b.gen_square[10].sq.piece[2] ;
 wire \b.gen_square[11].sq.color ;
 wire \b.gen_square[11].sq.mask ;
 wire \b.gen_square[11].sq.piece[0] ;
 wire \b.gen_square[11].sq.piece[1] ;
 wire \b.gen_square[11].sq.piece[2] ;
 wire \b.gen_square[12].sq.color ;
 wire \b.gen_square[12].sq.mask ;
 wire \b.gen_square[12].sq.piece[0] ;
 wire \b.gen_square[12].sq.piece[1] ;
 wire \b.gen_square[12].sq.piece[2] ;
 wire \b.gen_square[13].sq.color ;
 wire \b.gen_square[13].sq.mask ;
 wire \b.gen_square[13].sq.piece[0] ;
 wire \b.gen_square[13].sq.piece[1] ;
 wire \b.gen_square[13].sq.piece[2] ;
 wire \b.gen_square[14].sq.color ;
 wire \b.gen_square[14].sq.mask ;
 wire \b.gen_square[14].sq.piece[0] ;
 wire \b.gen_square[14].sq.piece[1] ;
 wire \b.gen_square[14].sq.piece[2] ;
 wire \b.gen_square[15].sq.color ;
 wire \b.gen_square[15].sq.mask ;
 wire \b.gen_square[15].sq.piece[0] ;
 wire \b.gen_square[15].sq.piece[1] ;
 wire \b.gen_square[15].sq.piece[2] ;
 wire \b.gen_square[16].sq.color ;
 wire \b.gen_square[16].sq.mask ;
 wire \b.gen_square[16].sq.piece[0] ;
 wire \b.gen_square[16].sq.piece[1] ;
 wire \b.gen_square[16].sq.piece[2] ;
 wire \b.gen_square[17].sq.color ;
 wire \b.gen_square[17].sq.mask ;
 wire \b.gen_square[17].sq.piece[0] ;
 wire \b.gen_square[17].sq.piece[1] ;
 wire \b.gen_square[17].sq.piece[2] ;
 wire \b.gen_square[18].sq.color ;
 wire \b.gen_square[18].sq.mask ;
 wire \b.gen_square[18].sq.piece[0] ;
 wire \b.gen_square[18].sq.piece[1] ;
 wire \b.gen_square[18].sq.piece[2] ;
 wire \b.gen_square[19].sq.color ;
 wire \b.gen_square[19].sq.mask ;
 wire \b.gen_square[19].sq.piece[0] ;
 wire \b.gen_square[19].sq.piece[1] ;
 wire \b.gen_square[19].sq.piece[2] ;
 wire \b.gen_square[1].sq.color ;
 wire \b.gen_square[1].sq.mask ;
 wire \b.gen_square[1].sq.piece[0] ;
 wire \b.gen_square[1].sq.piece[1] ;
 wire \b.gen_square[1].sq.piece[2] ;
 wire \b.gen_square[20].sq.color ;
 wire \b.gen_square[20].sq.mask ;
 wire \b.gen_square[20].sq.piece[0] ;
 wire \b.gen_square[20].sq.piece[1] ;
 wire \b.gen_square[20].sq.piece[2] ;
 wire \b.gen_square[21].sq.color ;
 wire \b.gen_square[21].sq.mask ;
 wire \b.gen_square[21].sq.piece[0] ;
 wire \b.gen_square[21].sq.piece[1] ;
 wire \b.gen_square[21].sq.piece[2] ;
 wire \b.gen_square[22].sq.color ;
 wire \b.gen_square[22].sq.mask ;
 wire \b.gen_square[22].sq.piece[0] ;
 wire \b.gen_square[22].sq.piece[1] ;
 wire \b.gen_square[22].sq.piece[2] ;
 wire \b.gen_square[23].sq.color ;
 wire \b.gen_square[23].sq.mask ;
 wire \b.gen_square[23].sq.piece[0] ;
 wire \b.gen_square[23].sq.piece[1] ;
 wire \b.gen_square[23].sq.piece[2] ;
 wire \b.gen_square[24].sq.color ;
 wire \b.gen_square[24].sq.mask ;
 wire \b.gen_square[24].sq.piece[0] ;
 wire \b.gen_square[24].sq.piece[1] ;
 wire \b.gen_square[24].sq.piece[2] ;
 wire \b.gen_square[25].sq.color ;
 wire \b.gen_square[25].sq.mask ;
 wire \b.gen_square[25].sq.piece[0] ;
 wire \b.gen_square[25].sq.piece[1] ;
 wire \b.gen_square[25].sq.piece[2] ;
 wire \b.gen_square[26].sq.color ;
 wire \b.gen_square[26].sq.mask ;
 wire \b.gen_square[26].sq.piece[0] ;
 wire \b.gen_square[26].sq.piece[1] ;
 wire \b.gen_square[26].sq.piece[2] ;
 wire \b.gen_square[27].sq.color ;
 wire \b.gen_square[27].sq.mask ;
 wire \b.gen_square[27].sq.piece[0] ;
 wire \b.gen_square[27].sq.piece[1] ;
 wire \b.gen_square[27].sq.piece[2] ;
 wire \b.gen_square[28].sq.color ;
 wire \b.gen_square[28].sq.mask ;
 wire \b.gen_square[28].sq.piece[0] ;
 wire \b.gen_square[28].sq.piece[1] ;
 wire \b.gen_square[28].sq.piece[2] ;
 wire \b.gen_square[29].sq.color ;
 wire \b.gen_square[29].sq.mask ;
 wire \b.gen_square[29].sq.piece[0] ;
 wire \b.gen_square[29].sq.piece[1] ;
 wire \b.gen_square[29].sq.piece[2] ;
 wire \b.gen_square[2].sq.color ;
 wire \b.gen_square[2].sq.mask ;
 wire \b.gen_square[2].sq.piece[0] ;
 wire \b.gen_square[2].sq.piece[1] ;
 wire \b.gen_square[2].sq.piece[2] ;
 wire \b.gen_square[30].sq.color ;
 wire \b.gen_square[30].sq.mask ;
 wire \b.gen_square[30].sq.piece[0] ;
 wire \b.gen_square[30].sq.piece[1] ;
 wire \b.gen_square[30].sq.piece[2] ;
 wire \b.gen_square[31].sq.color ;
 wire \b.gen_square[31].sq.mask ;
 wire \b.gen_square[31].sq.piece[0] ;
 wire \b.gen_square[31].sq.piece[1] ;
 wire \b.gen_square[31].sq.piece[2] ;
 wire \b.gen_square[32].sq.color ;
 wire \b.gen_square[32].sq.mask ;
 wire \b.gen_square[32].sq.piece[0] ;
 wire \b.gen_square[32].sq.piece[1] ;
 wire \b.gen_square[32].sq.piece[2] ;
 wire \b.gen_square[33].sq.color ;
 wire \b.gen_square[33].sq.mask ;
 wire \b.gen_square[33].sq.piece[0] ;
 wire \b.gen_square[33].sq.piece[1] ;
 wire \b.gen_square[33].sq.piece[2] ;
 wire \b.gen_square[34].sq.color ;
 wire \b.gen_square[34].sq.mask ;
 wire \b.gen_square[34].sq.piece[0] ;
 wire \b.gen_square[34].sq.piece[1] ;
 wire \b.gen_square[34].sq.piece[2] ;
 wire \b.gen_square[35].sq.color ;
 wire \b.gen_square[35].sq.mask ;
 wire \b.gen_square[35].sq.piece[0] ;
 wire \b.gen_square[35].sq.piece[1] ;
 wire \b.gen_square[35].sq.piece[2] ;
 wire \b.gen_square[36].sq.color ;
 wire \b.gen_square[36].sq.mask ;
 wire \b.gen_square[36].sq.piece[0] ;
 wire \b.gen_square[36].sq.piece[1] ;
 wire \b.gen_square[36].sq.piece[2] ;
 wire \b.gen_square[37].sq.color ;
 wire \b.gen_square[37].sq.mask ;
 wire \b.gen_square[37].sq.piece[0] ;
 wire \b.gen_square[37].sq.piece[1] ;
 wire \b.gen_square[37].sq.piece[2] ;
 wire \b.gen_square[38].sq.color ;
 wire \b.gen_square[38].sq.mask ;
 wire \b.gen_square[38].sq.piece[0] ;
 wire \b.gen_square[38].sq.piece[1] ;
 wire \b.gen_square[38].sq.piece[2] ;
 wire \b.gen_square[39].sq.color ;
 wire \b.gen_square[39].sq.mask ;
 wire \b.gen_square[39].sq.piece[0] ;
 wire \b.gen_square[39].sq.piece[1] ;
 wire \b.gen_square[39].sq.piece[2] ;
 wire \b.gen_square[3].sq.color ;
 wire \b.gen_square[3].sq.mask ;
 wire \b.gen_square[3].sq.piece[0] ;
 wire \b.gen_square[3].sq.piece[1] ;
 wire \b.gen_square[3].sq.piece[2] ;
 wire \b.gen_square[40].sq.color ;
 wire \b.gen_square[40].sq.mask ;
 wire \b.gen_square[40].sq.piece[0] ;
 wire \b.gen_square[40].sq.piece[1] ;
 wire \b.gen_square[40].sq.piece[2] ;
 wire \b.gen_square[41].sq.color ;
 wire \b.gen_square[41].sq.mask ;
 wire \b.gen_square[41].sq.piece[0] ;
 wire \b.gen_square[41].sq.piece[1] ;
 wire \b.gen_square[41].sq.piece[2] ;
 wire \b.gen_square[42].sq.color ;
 wire \b.gen_square[42].sq.mask ;
 wire \b.gen_square[42].sq.piece[0] ;
 wire \b.gen_square[42].sq.piece[1] ;
 wire \b.gen_square[42].sq.piece[2] ;
 wire \b.gen_square[43].sq.color ;
 wire \b.gen_square[43].sq.mask ;
 wire \b.gen_square[43].sq.piece[0] ;
 wire \b.gen_square[43].sq.piece[1] ;
 wire \b.gen_square[43].sq.piece[2] ;
 wire \b.gen_square[44].sq.color ;
 wire \b.gen_square[44].sq.mask ;
 wire \b.gen_square[44].sq.piece[0] ;
 wire \b.gen_square[44].sq.piece[1] ;
 wire \b.gen_square[44].sq.piece[2] ;
 wire \b.gen_square[45].sq.color ;
 wire \b.gen_square[45].sq.mask ;
 wire \b.gen_square[45].sq.piece[0] ;
 wire \b.gen_square[45].sq.piece[1] ;
 wire \b.gen_square[45].sq.piece[2] ;
 wire \b.gen_square[46].sq.color ;
 wire \b.gen_square[46].sq.mask ;
 wire \b.gen_square[46].sq.piece[0] ;
 wire \b.gen_square[46].sq.piece[1] ;
 wire \b.gen_square[46].sq.piece[2] ;
 wire \b.gen_square[47].sq.color ;
 wire \b.gen_square[47].sq.mask ;
 wire \b.gen_square[47].sq.piece[0] ;
 wire \b.gen_square[47].sq.piece[1] ;
 wire \b.gen_square[47].sq.piece[2] ;
 wire \b.gen_square[48].sq.color ;
 wire \b.gen_square[48].sq.mask ;
 wire \b.gen_square[48].sq.piece[0] ;
 wire \b.gen_square[48].sq.piece[1] ;
 wire \b.gen_square[48].sq.piece[2] ;
 wire \b.gen_square[49].sq.color ;
 wire \b.gen_square[49].sq.mask ;
 wire \b.gen_square[49].sq.piece[0] ;
 wire \b.gen_square[49].sq.piece[1] ;
 wire \b.gen_square[49].sq.piece[2] ;
 wire \b.gen_square[4].sq.color ;
 wire \b.gen_square[4].sq.mask ;
 wire \b.gen_square[4].sq.piece[0] ;
 wire \b.gen_square[4].sq.piece[1] ;
 wire \b.gen_square[4].sq.piece[2] ;
 wire \b.gen_square[50].sq.color ;
 wire \b.gen_square[50].sq.mask ;
 wire \b.gen_square[50].sq.piece[0] ;
 wire \b.gen_square[50].sq.piece[1] ;
 wire \b.gen_square[50].sq.piece[2] ;
 wire \b.gen_square[51].sq.color ;
 wire \b.gen_square[51].sq.mask ;
 wire \b.gen_square[51].sq.piece[0] ;
 wire \b.gen_square[51].sq.piece[1] ;
 wire \b.gen_square[51].sq.piece[2] ;
 wire \b.gen_square[52].sq.color ;
 wire \b.gen_square[52].sq.mask ;
 wire \b.gen_square[52].sq.piece[0] ;
 wire \b.gen_square[52].sq.piece[1] ;
 wire \b.gen_square[52].sq.piece[2] ;
 wire \b.gen_square[53].sq.color ;
 wire \b.gen_square[53].sq.mask ;
 wire \b.gen_square[53].sq.piece[0] ;
 wire \b.gen_square[53].sq.piece[1] ;
 wire \b.gen_square[53].sq.piece[2] ;
 wire \b.gen_square[54].sq.color ;
 wire \b.gen_square[54].sq.mask ;
 wire \b.gen_square[54].sq.piece[0] ;
 wire \b.gen_square[54].sq.piece[1] ;
 wire \b.gen_square[54].sq.piece[2] ;
 wire \b.gen_square[55].sq.color ;
 wire \b.gen_square[55].sq.mask ;
 wire \b.gen_square[55].sq.piece[0] ;
 wire \b.gen_square[55].sq.piece[1] ;
 wire \b.gen_square[55].sq.piece[2] ;
 wire \b.gen_square[56].sq.color ;
 wire \b.gen_square[56].sq.mask ;
 wire \b.gen_square[56].sq.piece[0] ;
 wire \b.gen_square[56].sq.piece[1] ;
 wire \b.gen_square[56].sq.piece[2] ;
 wire \b.gen_square[57].sq.color ;
 wire \b.gen_square[57].sq.mask ;
 wire \b.gen_square[57].sq.piece[0] ;
 wire \b.gen_square[57].sq.piece[1] ;
 wire \b.gen_square[57].sq.piece[2] ;
 wire \b.gen_square[58].sq.color ;
 wire \b.gen_square[58].sq.mask ;
 wire \b.gen_square[58].sq.piece[0] ;
 wire \b.gen_square[58].sq.piece[1] ;
 wire \b.gen_square[58].sq.piece[2] ;
 wire \b.gen_square[59].sq.color ;
 wire \b.gen_square[59].sq.mask ;
 wire \b.gen_square[59].sq.piece[0] ;
 wire \b.gen_square[59].sq.piece[1] ;
 wire \b.gen_square[59].sq.piece[2] ;
 wire \b.gen_square[5].sq.color ;
 wire \b.gen_square[5].sq.mask ;
 wire \b.gen_square[5].sq.piece[0] ;
 wire \b.gen_square[5].sq.piece[1] ;
 wire \b.gen_square[5].sq.piece[2] ;
 wire \b.gen_square[60].sq.color ;
 wire \b.gen_square[60].sq.mask ;
 wire \b.gen_square[60].sq.piece[0] ;
 wire \b.gen_square[60].sq.piece[1] ;
 wire \b.gen_square[60].sq.piece[2] ;
 wire \b.gen_square[61].sq.color ;
 wire \b.gen_square[61].sq.mask ;
 wire \b.gen_square[61].sq.piece[0] ;
 wire \b.gen_square[61].sq.piece[1] ;
 wire \b.gen_square[61].sq.piece[2] ;
 wire \b.gen_square[62].sq.color ;
 wire \b.gen_square[62].sq.mask ;
 wire \b.gen_square[62].sq.piece[0] ;
 wire \b.gen_square[62].sq.piece[1] ;
 wire \b.gen_square[62].sq.piece[2] ;
 wire \b.gen_square[63].sq.color ;
 wire \b.gen_square[63].sq.mask ;
 wire \b.gen_square[63].sq.piece[0] ;
 wire \b.gen_square[63].sq.piece[1] ;
 wire \b.gen_square[63].sq.piece[2] ;
 wire \b.gen_square[6].sq.color ;
 wire \b.gen_square[6].sq.mask ;
 wire \b.gen_square[6].sq.piece[0] ;
 wire \b.gen_square[6].sq.piece[1] ;
 wire \b.gen_square[6].sq.piece[2] ;
 wire \b.gen_square[7].sq.color ;
 wire \b.gen_square[7].sq.mask ;
 wire \b.gen_square[7].sq.piece[0] ;
 wire \b.gen_square[7].sq.piece[1] ;
 wire \b.gen_square[7].sq.piece[2] ;
 wire \b.gen_square[8].sq.color ;
 wire \b.gen_square[8].sq.mask ;
 wire \b.gen_square[8].sq.piece[0] ;
 wire \b.gen_square[8].sq.piece[1] ;
 wire \b.gen_square[8].sq.piece[2] ;
 wire \b.gen_square[9].sq.color ;
 wire \b.gen_square[9].sq.mask ;
 wire \b.gen_square[9].sq.piece[0] ;
 wire \b.gen_square[9].sq.piece[1] ;
 wire \b.gen_square[9].sq.piece[2] ;
 wire \b.ss1[0] ;
 wire \b.ss1[1] ;
 wire \b.ss1[2] ;
 wire \b.ss1[3] ;
 wire \b.ss1[4] ;
 wire \b.ss1[5] ;
 wire \data_in[0] ;
 wire \data_in[1] ;
 wire \data_in[2] ;
 wire \data_in[3] ;
 wire data_in_valid;
 wire \data_out[0] ;
 wire \data_out[1] ;
 wire \data_out[2] ;
 wire \data_out[3] ;
 wire data_out_valid;
 wire \mask_mode[1] ;
 wire \mask_mode[2] ;
 wire \mask_mode[3] ;
 wire \spi.bit_count ;
 wire \spi.sck_r0 ;
 wire \spi.sdi_r[0] ;
 wire \spi.sdi_r[1] ;
 wire \spi.sdi_r[2] ;
 wire \spi.sdi_r[3] ;
 wire \ss2[0] ;
 wire \ss2[1] ;
 wire \ss2[2] ;
 wire \ss2[3] ;
 wire \ss2[4] ;
 wire \ss2[5] ;
 wire \state[0] ;
 wire \state[10] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire \state[7] ;
 wire \state[8] ;
 wire \state[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_buf_2 _12133_ (.A(data_in_valid),
    .X(_00772_));
 sg13g2_buf_1 _12134_ (.A(\state[1] ),
    .X(_00783_));
 sg13g2_inv_1 _12135_ (.Y(_00794_),
    .A(_00783_));
 sg13g2_buf_2 _12136_ (.A(\data_in[0] ),
    .X(_00805_));
 sg13g2_buf_1 _12137_ (.A(\data_in[1] ),
    .X(_00816_));
 sg13g2_nand2_1 _12138_ (.Y(_00827_),
    .A(_00805_),
    .B(_00816_));
 sg13g2_inv_1 _12139_ (.Y(_00838_),
    .A(_00827_));
 sg13g2_buf_1 _12140_ (.A(\state[0] ),
    .X(_00849_));
 sg13g2_nand2_1 _12141_ (.Y(_00860_),
    .A(_00772_),
    .B(_00849_));
 sg13g2_inv_1 _12142_ (.Y(_00871_),
    .A(_00860_));
 sg13g2_buf_1 _12143_ (.A(_00871_),
    .X(_00882_));
 sg13g2_buf_1 _12144_ (.A(\data_in[2] ),
    .X(_00893_));
 sg13g2_buf_1 _12145_ (.A(\data_in[3] ),
    .X(_00904_));
 sg13g2_inv_1 _12146_ (.Y(_00915_),
    .A(_00904_));
 sg13g2_nor2_1 _12147_ (.A(_00893_),
    .B(_00915_),
    .Y(_00926_));
 sg13g2_nand3_1 _12148_ (.B(net184),
    .C(_00926_),
    .A(_00838_),
    .Y(_00937_));
 sg13g2_o21ai_1 _12149_ (.B1(_00937_),
    .Y(_00005_),
    .A1(_00772_),
    .A2(_00794_));
 sg13g2_inv_1 _12150_ (.Y(_00958_),
    .A(\state[2] ));
 sg13g2_inv_1 _12151_ (.Y(_00969_),
    .A(\spi.sck_r0 ));
 sg13g2_nand2_1 _12152_ (.Y(_00980_),
    .A(_00969_),
    .B(net3));
 sg13g2_inv_1 _12153_ (.Y(_00991_),
    .A(_00980_));
 sg13g2_inv_1 _12154_ (.Y(_01002_),
    .A(net2));
 sg13g2_buf_2 _12155_ (.A(net243),
    .X(_01013_));
 sg13g2_nand4_1 _12156_ (.B(data_out_valid),
    .C(_01002_),
    .A(_00991_),
    .Y(_01024_),
    .D(_01013_));
 sg13g2_buf_2 _12157_ (.A(_01024_),
    .X(_01035_));
 sg13g2_nor2_1 _12158_ (.A(_00958_),
    .B(_01035_),
    .Y(_01046_));
 sg13g2_buf_1 _12159_ (.A(_01046_),
    .X(_01057_));
 sg13g2_buf_1 _12160_ (.A(_01057_),
    .X(_00000_));
 sg13g2_buf_1 _12161_ (.A(\state[5] ),
    .X(_01078_));
 sg13g2_nor3_1 _12162_ (.A(\state[2] ),
    .B(_00849_),
    .C(_01078_),
    .Y(_01089_));
 sg13g2_inv_1 _12163_ (.Y(_01100_),
    .A(_00772_));
 sg13g2_nand2_1 _12164_ (.Y(_01111_),
    .A(_01100_),
    .B(_00849_));
 sg13g2_nand2_1 _12165_ (.Y(_01122_),
    .A(_01100_),
    .B(_01078_));
 sg13g2_nand3_1 _12166_ (.B(_01122_),
    .C(_00958_),
    .A(_01111_),
    .Y(_01133_));
 sg13g2_o21ai_1 _12167_ (.B1(\mask_mode[2] ),
    .Y(_01144_),
    .A1(_01089_),
    .A2(_01133_));
 sg13g2_inv_1 _12168_ (.Y(_01155_),
    .A(_00805_));
 sg13g2_nor2_1 _12169_ (.A(_00816_),
    .B(_01155_),
    .Y(_01166_));
 sg13g2_nand3_1 _12170_ (.B(net184),
    .C(_01166_),
    .A(_00926_),
    .Y(_01177_));
 sg13g2_nand3b_1 _12171_ (.B(_01144_),
    .C(_01177_),
    .Y(_00002_),
    .A_N(_00000_));
 sg13g2_inv_2 _12172_ (.Y(_01198_),
    .A(_01035_));
 sg13g2_nor2_1 _12173_ (.A(_00958_),
    .B(_01198_),
    .Y(_01209_));
 sg13g2_buf_1 _12174_ (.A(\mask_mode[1] ),
    .X(_01220_));
 sg13g2_buf_1 _12175_ (.A(_01220_),
    .X(_01231_));
 sg13g2_o21ai_1 _12176_ (.B1(_01231_),
    .Y(_01242_),
    .A1(_01089_),
    .A2(_01209_));
 sg13g2_nand2_1 _12177_ (.Y(_01253_),
    .A(_01111_),
    .B(_01122_));
 sg13g2_inv_1 _12178_ (.Y(_01264_),
    .A(_00068_));
 sg13g2_nand2_1 _12179_ (.Y(_01275_),
    .A(_01253_),
    .B(_01264_));
 sg13g2_nand2_1 _12180_ (.Y(_01286_),
    .A(_00893_),
    .B(_00904_));
 sg13g2_inv_1 _12181_ (.Y(_01297_),
    .A(_01286_));
 sg13g2_nor2_1 _12182_ (.A(_00805_),
    .B(_00816_),
    .Y(_01308_));
 sg13g2_nand3_1 _12183_ (.B(_01297_),
    .C(_01308_),
    .A(net184),
    .Y(_01319_));
 sg13g2_nand3_1 _12184_ (.B(_01275_),
    .C(_01319_),
    .A(_01242_),
    .Y(_00001_));
 sg13g2_inv_1 _12185_ (.Y(_01340_),
    .A(\state[9] ));
 sg13g2_buf_1 _12186_ (.A(\state[8] ),
    .X(_01351_));
 sg13g2_nor2_1 _12187_ (.A(_00783_),
    .B(_01078_),
    .Y(_01362_));
 sg13g2_inv_1 _12188_ (.Y(_01373_),
    .A(_01362_));
 sg13g2_nor2_1 _12189_ (.A(_01351_),
    .B(_01373_),
    .Y(_01384_));
 sg13g2_nand2_1 _12190_ (.Y(_01395_),
    .A(_01035_),
    .B(_01384_));
 sg13g2_inv_1 _12191_ (.Y(_01406_),
    .A(_00849_));
 sg13g2_nor2_1 _12192_ (.A(_00067_),
    .B(_01406_),
    .Y(_01417_));
 sg13g2_nand3_1 _12193_ (.B(_01297_),
    .C(_01417_),
    .A(_00838_),
    .Y(_01428_));
 sg13g2_o21ai_1 _12194_ (.B1(_01428_),
    .Y(_00010_),
    .A1(_01340_),
    .A2(_01395_));
 sg13g2_nor2_1 _12195_ (.A(\state[6] ),
    .B(\state[9] ),
    .Y(_01449_));
 sg13g2_nand2_1 _12196_ (.Y(_01460_),
    .A(_01198_),
    .B(_01384_));
 sg13g2_nand2_1 _12197_ (.Y(_01471_),
    .A(_01035_),
    .B(\state[10] ));
 sg13g2_o21ai_1 _12198_ (.B1(_01471_),
    .Y(_00004_),
    .A1(_01449_),
    .A2(_01460_));
 sg13g2_nor2_1 _12199_ (.A(_00893_),
    .B(_00904_),
    .Y(_01492_));
 sg13g2_nand3_1 _12200_ (.B(net184),
    .C(_01492_),
    .A(_00838_),
    .Y(_01503_));
 sg13g2_nand2_1 _12201_ (.Y(_01514_),
    .A(_01100_),
    .B(\state[3] ));
 sg13g2_nand2_1 _12202_ (.Y(_00006_),
    .A(_01503_),
    .B(_01514_));
 sg13g2_inv_1 _12203_ (.Y(_01535_),
    .A(\state[4] ));
 sg13g2_inv_1 _12204_ (.Y(_01546_),
    .A(_00816_));
 sg13g2_nor3_1 _12205_ (.A(_00805_),
    .B(_01546_),
    .C(_01286_),
    .Y(_01557_));
 sg13g2_nand2_1 _12206_ (.Y(_01568_),
    .A(_01557_),
    .B(_00882_));
 sg13g2_o21ai_1 _12207_ (.B1(_01568_),
    .Y(_00007_),
    .A1(_01535_),
    .A2(_01198_));
 sg13g2_nand3_1 _12208_ (.B(_01166_),
    .C(_01492_),
    .A(net184),
    .Y(_01589_));
 sg13g2_nand2_1 _12209_ (.Y(_00008_),
    .A(_01589_),
    .B(_01122_));
 sg13g2_inv_1 _12210_ (.Y(_01610_),
    .A(\state[6] ));
 sg13g2_nand3_1 _12211_ (.B(_01297_),
    .C(_01166_),
    .A(net184),
    .Y(_01621_));
 sg13g2_o21ai_1 _12212_ (.B1(_01621_),
    .Y(_00009_),
    .A1(_01610_),
    .A2(_01395_));
 sg13g2_buf_2 _12213_ (.A(\mask_mode[3] ),
    .X(_01642_));
 sg13g2_inv_2 _12214_ (.Y(_01653_),
    .A(_01642_));
 sg13g2_buf_1 _12215_ (.A(_01653_),
    .X(_01664_));
 sg13g2_nor3_1 _12216_ (.A(_01089_),
    .B(_01253_),
    .C(_01209_),
    .Y(_01675_));
 sg13g2_nand3_1 _12217_ (.B(_00926_),
    .C(_01308_),
    .A(_00882_),
    .Y(_01686_));
 sg13g2_o21ai_1 _12218_ (.B1(_01686_),
    .Y(_00003_),
    .A1(net209),
    .A2(_01675_));
 sg13g2_nor2b_1 _12219_ (.A(_00980_),
    .B_N(\spi.bit_count ),
    .Y(_00011_));
 sg13g2_inv_1 _12220_ (.Y(_01717_),
    .A(\state[3] ));
 sg13g2_nand2_1 _12221_ (.Y(_01728_),
    .A(_01100_),
    .B(_01351_));
 sg13g2_o21ai_1 _12222_ (.B1(_01728_),
    .Y(_00340_),
    .A1(_01717_),
    .A2(_01100_));
 sg13g2_a21o_1 _12223_ (.A2(_01198_),
    .A1(\state[4] ),
    .B1(_01209_),
    .X(_00341_));
 sg13g2_buf_1 _12224_ (.A(\b.gen_square[0].sq.color ),
    .X(_01759_));
 sg13g2_inv_1 _12225_ (.Y(_01770_),
    .A(_01759_));
 sg13g2_buf_8 _12226_ (.A(\b.ss1[5] ),
    .X(_01781_));
 sg13g2_buf_8 _12227_ (.A(\b.ss1[4] ),
    .X(_01792_));
 sg13g2_nor2_1 _12228_ (.A(_01781_),
    .B(_01792_),
    .Y(_01803_));
 sg13g2_buf_8 _12229_ (.A(_01803_),
    .X(_01814_));
 sg13g2_inv_2 _12230_ (.Y(_01825_),
    .A(_01814_));
 sg13g2_buf_1 _12231_ (.A(_01825_),
    .X(_01836_));
 sg13g2_buf_8 _12232_ (.A(\b.ss1[3] ),
    .X(_01847_));
 sg13g2_buf_8 _12233_ (.A(\b.ss1[2] ),
    .X(_01858_));
 sg13g2_nor2_1 _12234_ (.A(_01847_),
    .B(_01858_),
    .Y(_01869_));
 sg13g2_buf_2 _12235_ (.A(_01869_),
    .X(_01880_));
 sg13g2_buf_8 _12236_ (.A(\b.ss1[0] ),
    .X(_01891_));
 sg13g2_buf_8 _12237_ (.A(\b.ss1[1] ),
    .X(_01902_));
 sg13g2_nor2_2 _12238_ (.A(_01891_),
    .B(_01902_),
    .Y(_01913_));
 sg13g2_nand2_2 _12239_ (.Y(_01924_),
    .A(_01880_),
    .B(_01913_));
 sg13g2_nor2_1 _12240_ (.A(net171),
    .B(_01924_),
    .Y(_01935_));
 sg13g2_buf_2 _12241_ (.A(\b.gen_square[0].sq.state_mode[2] ),
    .X(_01946_));
 sg13g2_inv_2 _12242_ (.Y(_01957_),
    .A(_01946_));
 sg13g2_buf_8 _12243_ (.A(\b.gen_square[0].sq.state_mode[0] ),
    .X(_01968_));
 sg13g2_buf_8 _12244_ (.A(\b.gen_square[0].sq.state_mode[1] ),
    .X(_01979_));
 sg13g2_inv_4 _12245_ (.A(_01979_),
    .Y(_01990_));
 sg13g2_nor2_1 _12246_ (.A(_01968_),
    .B(_01990_),
    .Y(_02001_));
 sg13g2_buf_8 _12247_ (.A(_02001_),
    .X(_02012_));
 sg13g2_inv_4 _12248_ (.A(net183),
    .Y(_02023_));
 sg13g2_buf_1 _12249_ (.A(_02023_),
    .X(_02034_));
 sg13g2_buf_1 _12250_ (.A(_02034_),
    .X(_02045_));
 sg13g2_buf_1 _12251_ (.A(net137),
    .X(_02056_));
 sg13g2_buf_1 _12252_ (.A(net120),
    .X(_02067_));
 sg13g2_buf_1 _12253_ (.A(net103),
    .X(_02078_));
 sg13g2_buf_1 _12254_ (.A(net93),
    .X(_02089_));
 sg13g2_buf_1 _12255_ (.A(net83),
    .X(_02100_));
 sg13g2_buf_1 _12256_ (.A(net72),
    .X(_02111_));
 sg13g2_buf_1 _12257_ (.A(net63),
    .X(_02122_));
 sg13g2_nor2_1 _12258_ (.A(_01957_),
    .B(net48),
    .Y(_02133_));
 sg13g2_buf_1 _12259_ (.A(_02133_),
    .X(_02144_));
 sg13g2_buf_1 _12260_ (.A(net24),
    .X(_02155_));
 sg13g2_nand2_1 _12261_ (.Y(_02166_),
    .A(_01935_),
    .B(net20));
 sg13g2_buf_2 _12262_ (.A(_02166_),
    .X(_02177_));
 sg13g2_buf_2 _12263_ (.A(\b.gen_square[0].sq.write_bus[3] ),
    .X(_02188_));
 sg13g2_buf_1 _12264_ (.A(_02188_),
    .X(_02199_));
 sg13g2_nor2_1 _12265_ (.A(net228),
    .B(_02177_),
    .Y(_02210_));
 sg13g2_a21oi_1 _12266_ (.A1(_01770_),
    .A2(_02177_),
    .Y(_00342_),
    .B1(_02210_));
 sg13g2_inv_1 _12267_ (.Y(_02231_),
    .A(_00080_));
 sg13g2_buf_1 _12268_ (.A(_02231_),
    .X(_02242_));
 sg13g2_buf_1 _12269_ (.A(net227),
    .X(_02253_));
 sg13g2_nand2_1 _12270_ (.Y(_02264_),
    .A(_02177_),
    .B(_00081_));
 sg13g2_o21ai_1 _12271_ (.B1(_02264_),
    .Y(_00343_),
    .A1(net208),
    .A2(_02177_));
 sg13g2_inv_1 _12272_ (.Y(_02285_),
    .A(_00079_));
 sg13g2_buf_1 _12273_ (.A(_02285_),
    .X(_02296_));
 sg13g2_buf_1 _12274_ (.A(net226),
    .X(_02307_));
 sg13g2_nand2_1 _12275_ (.Y(_02318_),
    .A(_02177_),
    .B(_00082_));
 sg13g2_o21ai_1 _12276_ (.B1(_02318_),
    .Y(_00344_),
    .A1(net207),
    .A2(_02177_));
 sg13g2_inv_1 _12277_ (.Y(_02339_),
    .A(_00078_));
 sg13g2_buf_1 _12278_ (.A(_02339_),
    .X(_02350_));
 sg13g2_buf_1 _12279_ (.A(net225),
    .X(_02361_));
 sg13g2_nand2_1 _12280_ (.Y(_02372_),
    .A(_02177_),
    .B(_00083_));
 sg13g2_o21ai_1 _12281_ (.B1(_02372_),
    .Y(_00345_),
    .A1(net206),
    .A2(_02177_));
 sg13g2_inv_1 _12282_ (.Y(_02393_),
    .A(\b.gen_square[10].sq.color ));
 sg13g2_inv_2 _12283_ (.Y(_02404_),
    .A(_01858_));
 sg13g2_nand2_1 _12284_ (.Y(_02415_),
    .A(_02404_),
    .B(_01847_));
 sg13g2_inv_1 _12285_ (.Y(_02426_),
    .A(_01891_));
 sg13g2_nand2_1 _12286_ (.Y(_02437_),
    .A(_02426_),
    .B(_01902_));
 sg13g2_nor2_1 _12287_ (.A(_02415_),
    .B(_02437_),
    .Y(_02448_));
 sg13g2_buf_2 _12288_ (.A(_02448_),
    .X(_02459_));
 sg13g2_nand2_1 _12289_ (.Y(_02470_),
    .A(_02459_),
    .B(_01814_));
 sg13g2_inv_1 _12290_ (.Y(_02481_),
    .A(_02470_));
 sg13g2_nand2_1 _12291_ (.Y(_02492_),
    .A(_02481_),
    .B(net20));
 sg13g2_buf_2 _12292_ (.A(_02492_),
    .X(_02503_));
 sg13g2_nor2_1 _12293_ (.A(_02199_),
    .B(_02503_),
    .Y(_02514_));
 sg13g2_a21oi_1 _12294_ (.A1(_02393_),
    .A2(_02503_),
    .Y(_00346_),
    .B1(_02514_));
 sg13g2_nand2_1 _12295_ (.Y(_02535_),
    .A(_02503_),
    .B(_00084_));
 sg13g2_o21ai_1 _12296_ (.B1(_02535_),
    .Y(_00347_),
    .A1(net208),
    .A2(_02503_));
 sg13g2_nand2_1 _12297_ (.Y(_02556_),
    .A(_02503_),
    .B(_00085_));
 sg13g2_o21ai_1 _12298_ (.B1(_02556_),
    .Y(_00348_),
    .A1(net207),
    .A2(_02503_));
 sg13g2_nand2_1 _12299_ (.Y(_02577_),
    .A(_02503_),
    .B(_00086_));
 sg13g2_o21ai_1 _12300_ (.B1(_02577_),
    .Y(_00349_),
    .A1(net206),
    .A2(_02503_));
 sg13g2_inv_1 _12301_ (.Y(_02598_),
    .A(\b.gen_square[11].sq.color ));
 sg13g2_nand2_1 _12302_ (.Y(_02609_),
    .A(_01891_),
    .B(_01902_));
 sg13g2_nor2_1 _12303_ (.A(_02609_),
    .B(_02415_),
    .Y(_02620_));
 sg13g2_inv_2 _12304_ (.Y(_02631_),
    .A(_02620_));
 sg13g2_nor2_2 _12305_ (.A(net171),
    .B(_02631_),
    .Y(_02642_));
 sg13g2_nand2_1 _12306_ (.Y(_02653_),
    .A(_02642_),
    .B(net20));
 sg13g2_buf_2 _12307_ (.A(_02653_),
    .X(_02664_));
 sg13g2_nor2_1 _12308_ (.A(_02199_),
    .B(_02664_),
    .Y(_02675_));
 sg13g2_a21oi_1 _12309_ (.A1(_02598_),
    .A2(_02664_),
    .Y(_00350_),
    .B1(_02675_));
 sg13g2_nand2_1 _12310_ (.Y(_02696_),
    .A(_02664_),
    .B(_00087_));
 sg13g2_o21ai_1 _12311_ (.B1(_02696_),
    .Y(_00351_),
    .A1(net208),
    .A2(_02664_));
 sg13g2_nand2_1 _12312_ (.Y(_02717_),
    .A(_02664_),
    .B(_00088_));
 sg13g2_o21ai_1 _12313_ (.B1(_02717_),
    .Y(_00352_),
    .A1(net207),
    .A2(_02664_));
 sg13g2_nand2_1 _12314_ (.Y(_02738_),
    .A(_02664_),
    .B(_00089_));
 sg13g2_o21ai_1 _12315_ (.B1(_02738_),
    .Y(_00353_),
    .A1(net206),
    .A2(_02664_));
 sg13g2_inv_2 _12316_ (.Y(_02759_),
    .A(_02188_));
 sg13g2_inv_1 _12317_ (.Y(_02770_),
    .A(net24));
 sg13g2_nand2_1 _12318_ (.Y(_02781_),
    .A(_01847_),
    .B(_01858_));
 sg13g2_inv_2 _12319_ (.Y(_02792_),
    .A(_02781_));
 sg13g2_nand2_2 _12320_ (.Y(_02803_),
    .A(_02792_),
    .B(_01913_));
 sg13g2_nor2_1 _12321_ (.A(_01836_),
    .B(_02803_),
    .Y(_02814_));
 sg13g2_inv_1 _12322_ (.Y(_02824_),
    .A(_02814_));
 sg13g2_nor2_1 _12323_ (.A(_02770_),
    .B(_02824_),
    .Y(_02835_));
 sg13g2_buf_2 _12324_ (.A(_02835_),
    .X(_02846_));
 sg13g2_nor2_1 _12325_ (.A(\b.gen_square[12].sq.color ),
    .B(_02846_),
    .Y(_02857_));
 sg13g2_a21oi_1 _12326_ (.A1(_02759_),
    .A2(_02846_),
    .Y(_00354_),
    .B1(_02857_));
 sg13g2_nor2_1 _12327_ (.A(_00090_),
    .B(_02846_),
    .Y(_02877_));
 sg13g2_a21oi_1 _12328_ (.A1(net208),
    .A2(_02846_),
    .Y(_00355_),
    .B1(_02877_));
 sg13g2_nor2_1 _12329_ (.A(_00091_),
    .B(_02846_),
    .Y(_02897_));
 sg13g2_a21oi_1 _12330_ (.A1(net207),
    .A2(_02846_),
    .Y(_00356_),
    .B1(_02897_));
 sg13g2_nor2_1 _12331_ (.A(_00092_),
    .B(_02846_),
    .Y(_02918_));
 sg13g2_a21oi_1 _12332_ (.A1(net206),
    .A2(_02846_),
    .Y(_00357_),
    .B1(_02918_));
 sg13g2_inv_1 _12333_ (.Y(_02939_),
    .A(\b.gen_square[13].sq.color ));
 sg13g2_inv_4 _12334_ (.A(_01902_),
    .Y(_02950_));
 sg13g2_nand2_1 _12335_ (.Y(_02961_),
    .A(_02950_),
    .B(_01891_));
 sg13g2_nor2_1 _12336_ (.A(_02781_),
    .B(_02961_),
    .Y(_02972_));
 sg13g2_inv_2 _12337_ (.Y(_02983_),
    .A(_02972_));
 sg13g2_nor2_2 _12338_ (.A(_01825_),
    .B(_02983_),
    .Y(_02994_));
 sg13g2_nand2_1 _12339_ (.Y(_03003_),
    .A(_02994_),
    .B(net20));
 sg13g2_buf_2 _12340_ (.A(_03003_),
    .X(_03011_));
 sg13g2_nor2_1 _12341_ (.A(net228),
    .B(_03011_),
    .Y(_03016_));
 sg13g2_a21oi_1 _12342_ (.A1(_02939_),
    .A2(_03011_),
    .Y(_00358_),
    .B1(_03016_));
 sg13g2_nand2_1 _12343_ (.Y(_03033_),
    .A(_03011_),
    .B(_00093_));
 sg13g2_o21ai_1 _12344_ (.B1(_03033_),
    .Y(_00359_),
    .A1(net208),
    .A2(_03011_));
 sg13g2_nand2_1 _12345_ (.Y(_03046_),
    .A(_03011_),
    .B(_00094_));
 sg13g2_o21ai_1 _12346_ (.B1(_03046_),
    .Y(_00360_),
    .A1(net207),
    .A2(_03011_));
 sg13g2_nand2_1 _12347_ (.Y(_03060_),
    .A(_03011_),
    .B(_00095_));
 sg13g2_o21ai_1 _12348_ (.B1(_03060_),
    .Y(_00361_),
    .A1(net206),
    .A2(_03011_));
 sg13g2_inv_1 _12349_ (.Y(_03080_),
    .A(\b.gen_square[14].sq.color ));
 sg13g2_nor2_1 _12350_ (.A(_01891_),
    .B(_02950_),
    .Y(_03090_));
 sg13g2_nand2_1 _12351_ (.Y(_03100_),
    .A(_02792_),
    .B(_03090_));
 sg13g2_buf_2 _12352_ (.A(_03100_),
    .X(_03110_));
 sg13g2_nor2_2 _12353_ (.A(_01825_),
    .B(_03110_),
    .Y(_03119_));
 sg13g2_nand2_1 _12354_ (.Y(_03129_),
    .A(_03119_),
    .B(_02155_));
 sg13g2_buf_2 _12355_ (.A(_03129_),
    .X(_03139_));
 sg13g2_nor2_1 _12356_ (.A(net228),
    .B(_03139_),
    .Y(_03148_));
 sg13g2_a21oi_1 _12357_ (.A1(_03080_),
    .A2(_03139_),
    .Y(_00362_),
    .B1(_03148_));
 sg13g2_nand2_1 _12358_ (.Y(_03167_),
    .A(_03139_),
    .B(_00096_));
 sg13g2_o21ai_1 _12359_ (.B1(_03167_),
    .Y(_00363_),
    .A1(net208),
    .A2(_03139_));
 sg13g2_nand2_1 _12360_ (.Y(_03186_),
    .A(_03139_),
    .B(_00097_));
 sg13g2_o21ai_1 _12361_ (.B1(_03186_),
    .Y(_00364_),
    .A1(_02307_),
    .A2(_03139_));
 sg13g2_nand2_1 _12362_ (.Y(_03204_),
    .A(_03139_),
    .B(_00098_));
 sg13g2_o21ai_1 _12363_ (.B1(_03204_),
    .Y(_00365_),
    .A1(net206),
    .A2(_03139_));
 sg13g2_buf_2 _12364_ (.A(\b.gen_square[15].sq.color ),
    .X(_03221_));
 sg13g2_inv_1 _12365_ (.Y(_03231_),
    .A(_03221_));
 sg13g2_inv_1 _12366_ (.Y(_03241_),
    .A(_02609_));
 sg13g2_nand2_2 _12367_ (.Y(_03250_),
    .A(_03241_),
    .B(_02792_));
 sg13g2_nor2_1 _12368_ (.A(net171),
    .B(_03250_),
    .Y(_03260_));
 sg13g2_nand2_1 _12369_ (.Y(_03269_),
    .A(_03260_),
    .B(net20));
 sg13g2_buf_2 _12370_ (.A(_03269_),
    .X(_03279_));
 sg13g2_nor2_1 _12371_ (.A(net228),
    .B(_03279_),
    .Y(_03289_));
 sg13g2_a21oi_1 _12372_ (.A1(_03231_),
    .A2(_03279_),
    .Y(_00366_),
    .B1(_03289_));
 sg13g2_nand2_1 _12373_ (.Y(_03307_),
    .A(_03279_),
    .B(_00099_));
 sg13g2_o21ai_1 _12374_ (.B1(_03307_),
    .Y(_00367_),
    .A1(_02253_),
    .A2(_03279_));
 sg13g2_nand2_1 _12375_ (.Y(_03326_),
    .A(_03279_),
    .B(_00100_));
 sg13g2_o21ai_1 _12376_ (.B1(_03326_),
    .Y(_00368_),
    .A1(_02307_),
    .A2(_03279_));
 sg13g2_nand2_1 _12377_ (.Y(_03343_),
    .A(_03279_),
    .B(_00101_));
 sg13g2_o21ai_1 _12378_ (.B1(_03343_),
    .Y(_00369_),
    .A1(_02361_),
    .A2(_03279_));
 sg13g2_inv_1 _12379_ (.Y(_03362_),
    .A(\b.gen_square[16].sq.color ));
 sg13g2_inv_4 _12380_ (.A(_01792_),
    .Y(_03371_));
 sg13g2_nor2_1 _12381_ (.A(_01781_),
    .B(_03371_),
    .Y(_03381_));
 sg13g2_buf_8 _12382_ (.A(_03381_),
    .X(_03390_));
 sg13g2_inv_4 _12383_ (.A(net182),
    .Y(_03400_));
 sg13g2_nor2_1 _12384_ (.A(_03400_),
    .B(_01924_),
    .Y(_03409_));
 sg13g2_nand2_1 _12385_ (.Y(_03419_),
    .A(_03409_),
    .B(net20));
 sg13g2_buf_2 _12386_ (.A(_03419_),
    .X(_03429_));
 sg13g2_nor2_1 _12387_ (.A(net228),
    .B(_03429_),
    .Y(_03438_));
 sg13g2_a21oi_1 _12388_ (.A1(_03362_),
    .A2(_03429_),
    .Y(_00370_),
    .B1(_03438_));
 sg13g2_nand2_1 _12389_ (.Y(_03456_),
    .A(_03429_),
    .B(_00102_));
 sg13g2_o21ai_1 _12390_ (.B1(_03456_),
    .Y(_00371_),
    .A1(net208),
    .A2(_03429_));
 sg13g2_nand2_1 _12391_ (.Y(_03475_),
    .A(_03429_),
    .B(_00103_));
 sg13g2_o21ai_1 _12392_ (.B1(_03475_),
    .Y(_00372_),
    .A1(net207),
    .A2(_03429_));
 sg13g2_nand2_1 _12393_ (.Y(_03493_),
    .A(_03429_),
    .B(_00104_));
 sg13g2_o21ai_1 _12394_ (.B1(_03493_),
    .Y(_00373_),
    .A1(net206),
    .A2(_03429_));
 sg13g2_inv_1 _12395_ (.Y(_03512_),
    .A(\b.gen_square[17].sq.color ));
 sg13g2_buf_2 _12396_ (.A(_03400_),
    .X(_03521_));
 sg13g2_nor2_1 _12397_ (.A(_01902_),
    .B(_02426_),
    .Y(_03526_));
 sg13g2_nand2_2 _12398_ (.Y(_03527_),
    .A(_03526_),
    .B(_01880_));
 sg13g2_nor2_1 _12399_ (.A(net153),
    .B(_03527_),
    .Y(_03528_));
 sg13g2_nand2_1 _12400_ (.Y(_03529_),
    .A(_03528_),
    .B(net20));
 sg13g2_buf_2 _12401_ (.A(_03529_),
    .X(_03530_));
 sg13g2_nor2_1 _12402_ (.A(net228),
    .B(_03530_),
    .Y(_03531_));
 sg13g2_a21oi_1 _12403_ (.A1(_03512_),
    .A2(_03530_),
    .Y(_00374_),
    .B1(_03531_));
 sg13g2_nand2_1 _12404_ (.Y(_03532_),
    .A(_03530_),
    .B(_00105_));
 sg13g2_o21ai_1 _12405_ (.B1(_03532_),
    .Y(_00375_),
    .A1(net208),
    .A2(_03530_));
 sg13g2_nand2_1 _12406_ (.Y(_03533_),
    .A(_03530_),
    .B(_00106_));
 sg13g2_o21ai_1 _12407_ (.B1(_03533_),
    .Y(_00376_),
    .A1(net207),
    .A2(_03530_));
 sg13g2_nand2_1 _12408_ (.Y(_03534_),
    .A(_03530_),
    .B(_00107_));
 sg13g2_o21ai_1 _12409_ (.B1(_03534_),
    .Y(_00377_),
    .A1(net206),
    .A2(_03530_));
 sg13g2_inv_1 _12410_ (.Y(_03535_),
    .A(\b.gen_square[18].sq.color ));
 sg13g2_nand2_2 _12411_ (.Y(_03536_),
    .A(_03090_),
    .B(_01880_));
 sg13g2_nor2_1 _12412_ (.A(net153),
    .B(_03536_),
    .Y(_03537_));
 sg13g2_buf_1 _12413_ (.A(net24),
    .X(_03538_));
 sg13g2_nand2_1 _12414_ (.Y(_03539_),
    .A(_03537_),
    .B(net19));
 sg13g2_buf_2 _12415_ (.A(_03539_),
    .X(_03540_));
 sg13g2_nor2_1 _12416_ (.A(net228),
    .B(_03540_),
    .Y(_03541_));
 sg13g2_a21oi_1 _12417_ (.A1(_03535_),
    .A2(_03540_),
    .Y(_00378_),
    .B1(_03541_));
 sg13g2_buf_1 _12418_ (.A(net227),
    .X(_03542_));
 sg13g2_nand2_1 _12419_ (.Y(_03543_),
    .A(_03540_),
    .B(_00108_));
 sg13g2_o21ai_1 _12420_ (.B1(_03543_),
    .Y(_00379_),
    .A1(net205),
    .A2(_03540_));
 sg13g2_buf_1 _12421_ (.A(net226),
    .X(_03544_));
 sg13g2_nand2_1 _12422_ (.Y(_03545_),
    .A(_03540_),
    .B(_00109_));
 sg13g2_o21ai_1 _12423_ (.B1(_03545_),
    .Y(_00380_),
    .A1(net204),
    .A2(_03540_));
 sg13g2_buf_1 _12424_ (.A(net225),
    .X(_03546_));
 sg13g2_nand2_1 _12425_ (.Y(_03547_),
    .A(_03540_),
    .B(_00110_));
 sg13g2_o21ai_1 _12426_ (.B1(_03547_),
    .Y(_00381_),
    .A1(net203),
    .A2(_03540_));
 sg13g2_inv_1 _12427_ (.Y(_03548_),
    .A(\b.gen_square[19].sq.color ));
 sg13g2_nand2_2 _12428_ (.Y(_03549_),
    .A(_03241_),
    .B(_01880_));
 sg13g2_nor2_2 _12429_ (.A(_03521_),
    .B(_03549_),
    .Y(_03550_));
 sg13g2_nand2_1 _12430_ (.Y(_03551_),
    .A(_03550_),
    .B(_03538_));
 sg13g2_buf_2 _12431_ (.A(_03551_),
    .X(_03552_));
 sg13g2_nor2_1 _12432_ (.A(net228),
    .B(_03552_),
    .Y(_03553_));
 sg13g2_a21oi_1 _12433_ (.A1(_03548_),
    .A2(_03552_),
    .Y(_00382_),
    .B1(_03553_));
 sg13g2_nand2_1 _12434_ (.Y(_03554_),
    .A(_03552_),
    .B(_00111_));
 sg13g2_o21ai_1 _12435_ (.B1(_03554_),
    .Y(_00383_),
    .A1(net205),
    .A2(_03552_));
 sg13g2_nand2_1 _12436_ (.Y(_03555_),
    .A(_03552_),
    .B(_00112_));
 sg13g2_o21ai_1 _12437_ (.B1(_03555_),
    .Y(_00384_),
    .A1(net204),
    .A2(_03552_));
 sg13g2_nand2_1 _12438_ (.Y(_03556_),
    .A(_03552_),
    .B(_00113_));
 sg13g2_o21ai_1 _12439_ (.B1(_03556_),
    .Y(_00385_),
    .A1(net203),
    .A2(_03552_));
 sg13g2_buf_1 _12440_ (.A(\b.gen_square[1].sq.color ),
    .X(_03557_));
 sg13g2_inv_1 _12441_ (.Y(_03558_),
    .A(_03557_));
 sg13g2_nor2_1 _12442_ (.A(net171),
    .B(_03527_),
    .Y(_03559_));
 sg13g2_nand2_1 _12443_ (.Y(_03560_),
    .A(_03559_),
    .B(net19));
 sg13g2_buf_2 _12444_ (.A(_03560_),
    .X(_03561_));
 sg13g2_buf_1 _12445_ (.A(_02188_),
    .X(_03562_));
 sg13g2_nor2_1 _12446_ (.A(net224),
    .B(_03561_),
    .Y(_03563_));
 sg13g2_a21oi_1 _12447_ (.A1(_03558_),
    .A2(_03561_),
    .Y(_00386_),
    .B1(_03563_));
 sg13g2_nand2_1 _12448_ (.Y(_03564_),
    .A(_03561_),
    .B(_00114_));
 sg13g2_o21ai_1 _12449_ (.B1(_03564_),
    .Y(_00387_),
    .A1(net205),
    .A2(_03561_));
 sg13g2_nand2_1 _12450_ (.Y(_03565_),
    .A(_03561_),
    .B(_00115_));
 sg13g2_o21ai_1 _12451_ (.B1(_03565_),
    .Y(_00388_),
    .A1(net204),
    .A2(_03561_));
 sg13g2_nand2_1 _12452_ (.Y(_03566_),
    .A(_03561_),
    .B(_00116_));
 sg13g2_o21ai_1 _12453_ (.B1(_03566_),
    .Y(_00389_),
    .A1(net203),
    .A2(_03561_));
 sg13g2_inv_1 _12454_ (.Y(_03567_),
    .A(\b.gen_square[20].sq.color ));
 sg13g2_inv_4 _12455_ (.A(_01847_),
    .Y(_03568_));
 sg13g2_nand2_1 _12456_ (.Y(_03569_),
    .A(_03568_),
    .B(_01858_));
 sg13g2_nor2b_1 _12457_ (.A(_03569_),
    .B_N(_01913_),
    .Y(_03570_));
 sg13g2_inv_2 _12458_ (.Y(_03571_),
    .A(_03570_));
 sg13g2_nor2_2 _12459_ (.A(net153),
    .B(_03571_),
    .Y(_03572_));
 sg13g2_nand2_1 _12460_ (.Y(_03573_),
    .A(_03572_),
    .B(net19));
 sg13g2_buf_2 _12461_ (.A(_03573_),
    .X(_03574_));
 sg13g2_nor2_1 _12462_ (.A(net224),
    .B(_03574_),
    .Y(_03575_));
 sg13g2_a21oi_1 _12463_ (.A1(_03567_),
    .A2(_03574_),
    .Y(_00390_),
    .B1(_03575_));
 sg13g2_nand2_1 _12464_ (.Y(_03576_),
    .A(_03574_),
    .B(_00117_));
 sg13g2_o21ai_1 _12465_ (.B1(_03576_),
    .Y(_00391_),
    .A1(net205),
    .A2(_03574_));
 sg13g2_nand2_1 _12466_ (.Y(_03577_),
    .A(_03574_),
    .B(_00118_));
 sg13g2_o21ai_1 _12467_ (.B1(_03577_),
    .Y(_00392_),
    .A1(net204),
    .A2(_03574_));
 sg13g2_nand2_1 _12468_ (.Y(_03578_),
    .A(_03574_),
    .B(_00119_));
 sg13g2_o21ai_1 _12469_ (.B1(_03578_),
    .Y(_00393_),
    .A1(net203),
    .A2(_03574_));
 sg13g2_inv_1 _12470_ (.Y(_03579_),
    .A(\b.gen_square[21].sq.color ));
 sg13g2_nor2_1 _12471_ (.A(_02961_),
    .B(_03569_),
    .Y(_03580_));
 sg13g2_buf_8 _12472_ (.A(_03580_),
    .X(_03581_));
 sg13g2_nand2_1 _12473_ (.Y(_03582_),
    .A(_03581_),
    .B(_03390_));
 sg13g2_inv_1 _12474_ (.Y(_03583_),
    .A(_03582_));
 sg13g2_nand2_1 _12475_ (.Y(_03584_),
    .A(_03583_),
    .B(_03538_));
 sg13g2_buf_2 _12476_ (.A(_03584_),
    .X(_03585_));
 sg13g2_nor2_1 _12477_ (.A(net224),
    .B(_03585_),
    .Y(_03586_));
 sg13g2_a21oi_1 _12478_ (.A1(_03579_),
    .A2(_03585_),
    .Y(_00394_),
    .B1(_03586_));
 sg13g2_nand2_1 _12479_ (.Y(_03587_),
    .A(_03585_),
    .B(_00120_));
 sg13g2_o21ai_1 _12480_ (.B1(_03587_),
    .Y(_00395_),
    .A1(net205),
    .A2(_03585_));
 sg13g2_nand2_1 _12481_ (.Y(_03588_),
    .A(_03585_),
    .B(_00121_));
 sg13g2_o21ai_1 _12482_ (.B1(_03588_),
    .Y(_00396_),
    .A1(net204),
    .A2(_03585_));
 sg13g2_nand2_1 _12483_ (.Y(_03589_),
    .A(_03585_),
    .B(_00122_));
 sg13g2_o21ai_1 _12484_ (.B1(_03589_),
    .Y(_00397_),
    .A1(net203),
    .A2(_03585_));
 sg13g2_inv_1 _12485_ (.Y(_03590_),
    .A(\b.gen_square[22].sq.color ));
 sg13g2_nor2_1 _12486_ (.A(_02437_),
    .B(_03569_),
    .Y(_03591_));
 sg13g2_buf_8 _12487_ (.A(_03591_),
    .X(_03592_));
 sg13g2_nand2_1 _12488_ (.Y(_03593_),
    .A(_03592_),
    .B(net182));
 sg13g2_inv_1 _12489_ (.Y(_03594_),
    .A(_03593_));
 sg13g2_nand2_1 _12490_ (.Y(_03595_),
    .A(_03594_),
    .B(net19));
 sg13g2_buf_2 _12491_ (.A(_03595_),
    .X(_03596_));
 sg13g2_nor2_1 _12492_ (.A(_03562_),
    .B(_03596_),
    .Y(_03597_));
 sg13g2_a21oi_1 _12493_ (.A1(_03590_),
    .A2(_03596_),
    .Y(_00398_),
    .B1(_03597_));
 sg13g2_nand2_1 _12494_ (.Y(_03598_),
    .A(_03596_),
    .B(_00123_));
 sg13g2_o21ai_1 _12495_ (.B1(_03598_),
    .Y(_00399_),
    .A1(_03542_),
    .A2(_03596_));
 sg13g2_nand2_1 _12496_ (.Y(_03599_),
    .A(_03596_),
    .B(_00124_));
 sg13g2_o21ai_1 _12497_ (.B1(_03599_),
    .Y(_00400_),
    .A1(_03544_),
    .A2(_03596_));
 sg13g2_nand2_1 _12498_ (.Y(_03600_),
    .A(_03596_),
    .B(_00125_));
 sg13g2_o21ai_1 _12499_ (.B1(_03600_),
    .Y(_00401_),
    .A1(_03546_),
    .A2(_03596_));
 sg13g2_inv_1 _12500_ (.Y(_03601_),
    .A(\b.gen_square[23].sq.color ));
 sg13g2_buf_1 _12501_ (.A(net24),
    .X(_03602_));
 sg13g2_nor2_1 _12502_ (.A(_02609_),
    .B(_03569_),
    .Y(_03603_));
 sg13g2_buf_8 _12503_ (.A(_03603_),
    .X(_03604_));
 sg13g2_nand3_1 _12504_ (.B(net182),
    .C(_03604_),
    .A(net18),
    .Y(_03605_));
 sg13g2_buf_2 _12505_ (.A(_03605_),
    .X(_03606_));
 sg13g2_nor2_1 _12506_ (.A(_03562_),
    .B(_03606_),
    .Y(_03607_));
 sg13g2_a21oi_1 _12507_ (.A1(_03601_),
    .A2(_03606_),
    .Y(_00402_),
    .B1(_03607_));
 sg13g2_nand2_1 _12508_ (.Y(_03608_),
    .A(_03606_),
    .B(_00126_));
 sg13g2_o21ai_1 _12509_ (.B1(_03608_),
    .Y(_00403_),
    .A1(_03542_),
    .A2(_03606_));
 sg13g2_nand2_1 _12510_ (.Y(_03609_),
    .A(_03606_),
    .B(_00127_));
 sg13g2_o21ai_1 _12511_ (.B1(_03609_),
    .Y(_00404_),
    .A1(_03544_),
    .A2(_03606_));
 sg13g2_nand2_1 _12512_ (.Y(_03610_),
    .A(_03606_),
    .B(_00128_));
 sg13g2_o21ai_1 _12513_ (.B1(_03610_),
    .Y(_00405_),
    .A1(_03546_),
    .A2(_03606_));
 sg13g2_inv_1 _12514_ (.Y(_03611_),
    .A(\b.gen_square[24].sq.color ));
 sg13g2_nor2_1 _12515_ (.A(_01858_),
    .B(_03568_),
    .Y(_03612_));
 sg13g2_nand2_2 _12516_ (.Y(_03613_),
    .A(_03612_),
    .B(_01913_));
 sg13g2_nor2_1 _12517_ (.A(net153),
    .B(_03613_),
    .Y(_03614_));
 sg13g2_nand2_1 _12518_ (.Y(_03615_),
    .A(_03614_),
    .B(net19));
 sg13g2_buf_2 _12519_ (.A(_03615_),
    .X(_03616_));
 sg13g2_nor2_1 _12520_ (.A(net224),
    .B(_03616_),
    .Y(_03617_));
 sg13g2_a21oi_1 _12521_ (.A1(_03611_),
    .A2(_03616_),
    .Y(_00406_),
    .B1(_03617_));
 sg13g2_nand2_1 _12522_ (.Y(_03618_),
    .A(_03616_),
    .B(_00129_));
 sg13g2_o21ai_1 _12523_ (.B1(_03618_),
    .Y(_00407_),
    .A1(net205),
    .A2(_03616_));
 sg13g2_nand2_1 _12524_ (.Y(_03619_),
    .A(_03616_),
    .B(_00130_));
 sg13g2_o21ai_1 _12525_ (.B1(_03619_),
    .Y(_00408_),
    .A1(net204),
    .A2(_03616_));
 sg13g2_nand2_1 _12526_ (.Y(_03620_),
    .A(_03616_),
    .B(_00131_));
 sg13g2_o21ai_1 _12527_ (.B1(_03620_),
    .Y(_00409_),
    .A1(net203),
    .A2(_03616_));
 sg13g2_inv_1 _12528_ (.Y(_03621_),
    .A(\b.gen_square[25].sq.color ));
 sg13g2_nor2_1 _12529_ (.A(_02415_),
    .B(_02961_),
    .Y(_03622_));
 sg13g2_buf_2 _12530_ (.A(_03622_),
    .X(_03623_));
 sg13g2_nand2_1 _12531_ (.Y(_03624_),
    .A(_03623_),
    .B(net182));
 sg13g2_inv_1 _12532_ (.Y(_03625_),
    .A(_03624_));
 sg13g2_nand2_1 _12533_ (.Y(_03626_),
    .A(_03625_),
    .B(net19));
 sg13g2_buf_2 _12534_ (.A(_03626_),
    .X(_03627_));
 sg13g2_nor2_1 _12535_ (.A(net224),
    .B(_03627_),
    .Y(_03628_));
 sg13g2_a21oi_1 _12536_ (.A1(_03621_),
    .A2(_03627_),
    .Y(_00410_),
    .B1(_03628_));
 sg13g2_nand2_1 _12537_ (.Y(_03629_),
    .A(_03627_),
    .B(_00132_));
 sg13g2_o21ai_1 _12538_ (.B1(_03629_),
    .Y(_00411_),
    .A1(net205),
    .A2(_03627_));
 sg13g2_nand2_1 _12539_ (.Y(_03630_),
    .A(_03627_),
    .B(_00133_));
 sg13g2_o21ai_1 _12540_ (.B1(_03630_),
    .Y(_00412_),
    .A1(net204),
    .A2(_03627_));
 sg13g2_nand2_1 _12541_ (.Y(_03631_),
    .A(_03627_),
    .B(_00134_));
 sg13g2_o21ai_1 _12542_ (.B1(_03631_),
    .Y(_00413_),
    .A1(net203),
    .A2(_03627_));
 sg13g2_inv_1 _12543_ (.Y(_03632_),
    .A(\b.gen_square[26].sq.color ));
 sg13g2_nand3_1 _12544_ (.B(_02459_),
    .C(net182),
    .A(net18),
    .Y(_03633_));
 sg13g2_buf_2 _12545_ (.A(_03633_),
    .X(_03634_));
 sg13g2_nor2_1 _12546_ (.A(net224),
    .B(_03634_),
    .Y(_03635_));
 sg13g2_a21oi_1 _12547_ (.A1(_03632_),
    .A2(_03634_),
    .Y(_00414_),
    .B1(_03635_));
 sg13g2_nand2_1 _12548_ (.Y(_03636_),
    .A(_03634_),
    .B(_00135_));
 sg13g2_o21ai_1 _12549_ (.B1(_03636_),
    .Y(_00415_),
    .A1(net205),
    .A2(_03634_));
 sg13g2_nand2_1 _12550_ (.Y(_03637_),
    .A(_03634_),
    .B(_00136_));
 sg13g2_o21ai_1 _12551_ (.B1(_03637_),
    .Y(_00416_),
    .A1(net204),
    .A2(_03634_));
 sg13g2_nand2_1 _12552_ (.Y(_03638_),
    .A(_03634_),
    .B(_00137_));
 sg13g2_o21ai_1 _12553_ (.B1(_03638_),
    .Y(_00417_),
    .A1(net203),
    .A2(_03634_));
 sg13g2_inv_1 _12554_ (.Y(_03639_),
    .A(\b.gen_square[27].sq.color ));
 sg13g2_nor2_1 _12555_ (.A(net153),
    .B(_02631_),
    .Y(_03640_));
 sg13g2_nand2_1 _12556_ (.Y(_03641_),
    .A(_03640_),
    .B(net19));
 sg13g2_buf_2 _12557_ (.A(_03641_),
    .X(_03642_));
 sg13g2_nor2_1 _12558_ (.A(net224),
    .B(_03642_),
    .Y(_03643_));
 sg13g2_a21oi_1 _12559_ (.A1(_03639_),
    .A2(_03642_),
    .Y(_00418_),
    .B1(_03643_));
 sg13g2_buf_1 _12560_ (.A(net227),
    .X(_03644_));
 sg13g2_nand2_1 _12561_ (.Y(_03645_),
    .A(_03642_),
    .B(_00138_));
 sg13g2_o21ai_1 _12562_ (.B1(_03645_),
    .Y(_00419_),
    .A1(net202),
    .A2(_03642_));
 sg13g2_buf_1 _12563_ (.A(net226),
    .X(_03646_));
 sg13g2_nand2_1 _12564_ (.Y(_03647_),
    .A(_03642_),
    .B(_00139_));
 sg13g2_o21ai_1 _12565_ (.B1(_03647_),
    .Y(_00420_),
    .A1(net201),
    .A2(_03642_));
 sg13g2_buf_1 _12566_ (.A(net225),
    .X(_03648_));
 sg13g2_nand2_1 _12567_ (.Y(_03649_),
    .A(_03642_),
    .B(_00140_));
 sg13g2_o21ai_1 _12568_ (.B1(_03649_),
    .Y(_00421_),
    .A1(net200),
    .A2(_03642_));
 sg13g2_inv_1 _12569_ (.Y(_03650_),
    .A(\b.gen_square[28].sq.color ));
 sg13g2_nor2_2 _12570_ (.A(_03521_),
    .B(_02803_),
    .Y(_03651_));
 sg13g2_nand2_1 _12571_ (.Y(_03652_),
    .A(_03651_),
    .B(net19));
 sg13g2_buf_2 _12572_ (.A(_03652_),
    .X(_03653_));
 sg13g2_nor2_1 _12573_ (.A(net224),
    .B(_03653_),
    .Y(_03654_));
 sg13g2_a21oi_1 _12574_ (.A1(_03650_),
    .A2(_03653_),
    .Y(_00422_),
    .B1(_03654_));
 sg13g2_nand2_1 _12575_ (.Y(_03655_),
    .A(_03653_),
    .B(_00141_));
 sg13g2_o21ai_1 _12576_ (.B1(_03655_),
    .Y(_00423_),
    .A1(net202),
    .A2(_03653_));
 sg13g2_nand2_1 _12577_ (.Y(_03656_),
    .A(_03653_),
    .B(_00142_));
 sg13g2_o21ai_1 _12578_ (.B1(_03656_),
    .Y(_00424_),
    .A1(net201),
    .A2(_03653_));
 sg13g2_nand2_1 _12579_ (.Y(_03657_),
    .A(_03653_),
    .B(_00143_));
 sg13g2_o21ai_1 _12580_ (.B1(_03657_),
    .Y(_00425_),
    .A1(net200),
    .A2(_03653_));
 sg13g2_inv_1 _12581_ (.Y(_03658_),
    .A(\b.gen_square[29].sq.color ));
 sg13g2_nor2_2 _12582_ (.A(net153),
    .B(_02983_),
    .Y(_03659_));
 sg13g2_buf_1 _12583_ (.A(net24),
    .X(_03660_));
 sg13g2_nand2_1 _12584_ (.Y(_03661_),
    .A(_03659_),
    .B(net17));
 sg13g2_buf_2 _12585_ (.A(_03661_),
    .X(_03662_));
 sg13g2_buf_1 _12586_ (.A(_02188_),
    .X(_03663_));
 sg13g2_nor2_1 _12587_ (.A(net223),
    .B(_03662_),
    .Y(_03664_));
 sg13g2_a21oi_1 _12588_ (.A1(_03658_),
    .A2(_03662_),
    .Y(_00426_),
    .B1(_03664_));
 sg13g2_nand2_1 _12589_ (.Y(_03665_),
    .A(_03662_),
    .B(_00144_));
 sg13g2_o21ai_1 _12590_ (.B1(_03665_),
    .Y(_00427_),
    .A1(net202),
    .A2(_03662_));
 sg13g2_nand2_1 _12591_ (.Y(_03666_),
    .A(_03662_),
    .B(_00145_));
 sg13g2_o21ai_1 _12592_ (.B1(_03666_),
    .Y(_00428_),
    .A1(net201),
    .A2(_03662_));
 sg13g2_nand2_1 _12593_ (.Y(_03667_),
    .A(_03662_),
    .B(_00146_));
 sg13g2_o21ai_1 _12594_ (.B1(_03667_),
    .Y(_00429_),
    .A1(net200),
    .A2(_03662_));
 sg13g2_buf_1 _12595_ (.A(\b.gen_square[2].sq.color ),
    .X(_03668_));
 sg13g2_inv_1 _12596_ (.Y(_03669_),
    .A(_03668_));
 sg13g2_nor2_1 _12597_ (.A(net171),
    .B(_03536_),
    .Y(_03670_));
 sg13g2_nand2_1 _12598_ (.Y(_03671_),
    .A(_03670_),
    .B(_03660_));
 sg13g2_buf_2 _12599_ (.A(_03671_),
    .X(_03672_));
 sg13g2_nor2_1 _12600_ (.A(_03663_),
    .B(_03672_),
    .Y(_03673_));
 sg13g2_a21oi_1 _12601_ (.A1(_03669_),
    .A2(_03672_),
    .Y(_00430_),
    .B1(_03673_));
 sg13g2_nand2_1 _12602_ (.Y(_03674_),
    .A(_03672_),
    .B(_00147_));
 sg13g2_o21ai_1 _12603_ (.B1(_03674_),
    .Y(_00431_),
    .A1(_03644_),
    .A2(_03672_));
 sg13g2_nand2_1 _12604_ (.Y(_03675_),
    .A(_03672_),
    .B(_00148_));
 sg13g2_o21ai_1 _12605_ (.B1(_03675_),
    .Y(_00432_),
    .A1(_03646_),
    .A2(_03672_));
 sg13g2_nand2_1 _12606_ (.Y(_03676_),
    .A(_03672_),
    .B(_00149_));
 sg13g2_o21ai_1 _12607_ (.B1(_03676_),
    .Y(_00433_),
    .A1(_03648_),
    .A2(_03672_));
 sg13g2_inv_1 _12608_ (.Y(_03677_),
    .A(\b.gen_square[30].sq.color ));
 sg13g2_nor2_1 _12609_ (.A(net153),
    .B(_03110_),
    .Y(_03678_));
 sg13g2_nand2_1 _12610_ (.Y(_03679_),
    .A(_03678_),
    .B(_03660_));
 sg13g2_buf_2 _12611_ (.A(_03679_),
    .X(_03680_));
 sg13g2_nor2_1 _12612_ (.A(net223),
    .B(_03680_),
    .Y(_03681_));
 sg13g2_a21oi_1 _12613_ (.A1(_03677_),
    .A2(_03680_),
    .Y(_00434_),
    .B1(_03681_));
 sg13g2_nand2_1 _12614_ (.Y(_03682_),
    .A(_03680_),
    .B(_00150_));
 sg13g2_o21ai_1 _12615_ (.B1(_03682_),
    .Y(_00435_),
    .A1(_03644_),
    .A2(_03680_));
 sg13g2_nand2_1 _12616_ (.Y(_03683_),
    .A(_03680_),
    .B(_00151_));
 sg13g2_o21ai_1 _12617_ (.B1(_03683_),
    .Y(_00436_),
    .A1(_03646_),
    .A2(_03680_));
 sg13g2_nand2_1 _12618_ (.Y(_03684_),
    .A(_03680_),
    .B(_00152_));
 sg13g2_o21ai_1 _12619_ (.B1(_03684_),
    .Y(_00437_),
    .A1(_03648_),
    .A2(_03680_));
 sg13g2_inv_1 _12620_ (.Y(_03685_),
    .A(\b.gen_square[31].sq.color ));
 sg13g2_nor2_1 _12621_ (.A(net153),
    .B(_03250_),
    .Y(_03686_));
 sg13g2_nand2_1 _12622_ (.Y(_03687_),
    .A(_03686_),
    .B(net17));
 sg13g2_buf_2 _12623_ (.A(_03687_),
    .X(_03688_));
 sg13g2_nor2_1 _12624_ (.A(net223),
    .B(_03688_),
    .Y(_03689_));
 sg13g2_a21oi_1 _12625_ (.A1(_03685_),
    .A2(_03688_),
    .Y(_00438_),
    .B1(_03689_));
 sg13g2_nand2_1 _12626_ (.Y(_03690_),
    .A(_03688_),
    .B(_00153_));
 sg13g2_o21ai_1 _12627_ (.B1(_03690_),
    .Y(_00439_),
    .A1(net202),
    .A2(_03688_));
 sg13g2_nand2_1 _12628_ (.Y(_03691_),
    .A(_03688_),
    .B(_00154_));
 sg13g2_o21ai_1 _12629_ (.B1(_03691_),
    .Y(_00440_),
    .A1(net201),
    .A2(_03688_));
 sg13g2_nand2_1 _12630_ (.Y(_03692_),
    .A(_03688_),
    .B(_00155_));
 sg13g2_o21ai_1 _12631_ (.B1(_03692_),
    .Y(_00441_),
    .A1(net200),
    .A2(_03688_));
 sg13g2_inv_1 _12632_ (.Y(_03693_),
    .A(\b.gen_square[32].sq.color ));
 sg13g2_inv_2 _12633_ (.Y(_03694_),
    .A(_01781_));
 sg13g2_nor2_2 _12634_ (.A(_01792_),
    .B(_03694_),
    .Y(_03695_));
 sg13g2_inv_4 _12635_ (.A(_03695_),
    .Y(_03696_));
 sg13g2_buf_8 _12636_ (.A(_03696_),
    .X(_03697_));
 sg13g2_nor2_1 _12637_ (.A(net170),
    .B(_01924_),
    .Y(_03698_));
 sg13g2_nand2_1 _12638_ (.Y(_03699_),
    .A(_03698_),
    .B(net17));
 sg13g2_buf_2 _12639_ (.A(_03699_),
    .X(_03700_));
 sg13g2_nor2_1 _12640_ (.A(net223),
    .B(_03700_),
    .Y(_03701_));
 sg13g2_a21oi_1 _12641_ (.A1(_03693_),
    .A2(_03700_),
    .Y(_00442_),
    .B1(_03701_));
 sg13g2_nand2_1 _12642_ (.Y(_03702_),
    .A(_03700_),
    .B(_00156_));
 sg13g2_o21ai_1 _12643_ (.B1(_03702_),
    .Y(_00443_),
    .A1(net202),
    .A2(_03700_));
 sg13g2_nand2_1 _12644_ (.Y(_03703_),
    .A(_03700_),
    .B(_00157_));
 sg13g2_o21ai_1 _12645_ (.B1(_03703_),
    .Y(_00444_),
    .A1(net201),
    .A2(_03700_));
 sg13g2_nand2_1 _12646_ (.Y(_03704_),
    .A(_03700_),
    .B(_00158_));
 sg13g2_o21ai_1 _12647_ (.B1(_03704_),
    .Y(_00445_),
    .A1(net200),
    .A2(_03700_));
 sg13g2_inv_1 _12648_ (.Y(_03705_),
    .A(\b.gen_square[33].sq.color ));
 sg13g2_nor2_1 _12649_ (.A(_03696_),
    .B(_03527_),
    .Y(_03706_));
 sg13g2_nand2_1 _12650_ (.Y(_03707_),
    .A(_03706_),
    .B(net17));
 sg13g2_buf_2 _12651_ (.A(_03707_),
    .X(_03708_));
 sg13g2_nor2_1 _12652_ (.A(net223),
    .B(_03708_),
    .Y(_03709_));
 sg13g2_a21oi_1 _12653_ (.A1(_03705_),
    .A2(_03708_),
    .Y(_00446_),
    .B1(_03709_));
 sg13g2_nand2_1 _12654_ (.Y(_03710_),
    .A(_03708_),
    .B(_00159_));
 sg13g2_o21ai_1 _12655_ (.B1(_03710_),
    .Y(_00447_),
    .A1(net202),
    .A2(_03708_));
 sg13g2_nand2_1 _12656_ (.Y(_03711_),
    .A(_03708_),
    .B(_00160_));
 sg13g2_o21ai_1 _12657_ (.B1(_03711_),
    .Y(_00448_),
    .A1(net201),
    .A2(_03708_));
 sg13g2_nand2_1 _12658_ (.Y(_03712_),
    .A(_03708_),
    .B(_00161_));
 sg13g2_o21ai_1 _12659_ (.B1(_03712_),
    .Y(_00449_),
    .A1(net200),
    .A2(_03708_));
 sg13g2_inv_1 _12660_ (.Y(_03713_),
    .A(\b.gen_square[34].sq.color ));
 sg13g2_nor2_1 _12661_ (.A(net170),
    .B(_03536_),
    .Y(_03714_));
 sg13g2_nand2_1 _12662_ (.Y(_03715_),
    .A(_03714_),
    .B(net17));
 sg13g2_buf_2 _12663_ (.A(_03715_),
    .X(_03716_));
 sg13g2_nor2_1 _12664_ (.A(net223),
    .B(_03716_),
    .Y(_03717_));
 sg13g2_a21oi_1 _12665_ (.A1(_03713_),
    .A2(_03716_),
    .Y(_00450_),
    .B1(_03717_));
 sg13g2_nand2_1 _12666_ (.Y(_03718_),
    .A(_03716_),
    .B(_00162_));
 sg13g2_o21ai_1 _12667_ (.B1(_03718_),
    .Y(_00451_),
    .A1(net202),
    .A2(_03716_));
 sg13g2_nand2_1 _12668_ (.Y(_03719_),
    .A(_03716_),
    .B(_00163_));
 sg13g2_o21ai_1 _12669_ (.B1(_03719_),
    .Y(_00452_),
    .A1(net201),
    .A2(_03716_));
 sg13g2_nand2_1 _12670_ (.Y(_03720_),
    .A(_03716_),
    .B(_00164_));
 sg13g2_o21ai_1 _12671_ (.B1(_03720_),
    .Y(_00453_),
    .A1(net200),
    .A2(_03716_));
 sg13g2_inv_1 _12672_ (.Y(_03721_),
    .A(\b.gen_square[35].sq.color ));
 sg13g2_nor2_1 _12673_ (.A(net170),
    .B(_03549_),
    .Y(_03722_));
 sg13g2_nand2_1 _12674_ (.Y(_03723_),
    .A(_03722_),
    .B(net17));
 sg13g2_buf_2 _12675_ (.A(_03723_),
    .X(_03724_));
 sg13g2_nor2_1 _12676_ (.A(net223),
    .B(_03724_),
    .Y(_03725_));
 sg13g2_a21oi_1 _12677_ (.A1(_03721_),
    .A2(_03724_),
    .Y(_00454_),
    .B1(_03725_));
 sg13g2_nand2_1 _12678_ (.Y(_03726_),
    .A(_03724_),
    .B(_00165_));
 sg13g2_o21ai_1 _12679_ (.B1(_03726_),
    .Y(_00455_),
    .A1(net202),
    .A2(_03724_));
 sg13g2_nand2_1 _12680_ (.Y(_03727_),
    .A(_03724_),
    .B(_00166_));
 sg13g2_o21ai_1 _12681_ (.B1(_03727_),
    .Y(_00456_),
    .A1(net201),
    .A2(_03724_));
 sg13g2_nand2_1 _12682_ (.Y(_03728_),
    .A(_03724_),
    .B(_00167_));
 sg13g2_o21ai_1 _12683_ (.B1(_03728_),
    .Y(_00457_),
    .A1(net200),
    .A2(_03724_));
 sg13g2_inv_1 _12684_ (.Y(_03729_),
    .A(\b.gen_square[36].sq.color ));
 sg13g2_nor2_2 _12685_ (.A(_03697_),
    .B(_03571_),
    .Y(_03730_));
 sg13g2_nand2_1 _12686_ (.Y(_03731_),
    .A(_03730_),
    .B(net17));
 sg13g2_buf_2 _12687_ (.A(_03731_),
    .X(_03732_));
 sg13g2_nor2_1 _12688_ (.A(_03663_),
    .B(_03732_),
    .Y(_03733_));
 sg13g2_a21oi_1 _12689_ (.A1(_03729_),
    .A2(_03732_),
    .Y(_00458_),
    .B1(_03733_));
 sg13g2_buf_1 _12690_ (.A(net227),
    .X(_03734_));
 sg13g2_nand2_1 _12691_ (.Y(_03735_),
    .A(_03732_),
    .B(_00168_));
 sg13g2_o21ai_1 _12692_ (.B1(_03735_),
    .Y(_00459_),
    .A1(net199),
    .A2(_03732_));
 sg13g2_buf_1 _12693_ (.A(net226),
    .X(_03736_));
 sg13g2_nand2_1 _12694_ (.Y(_03737_),
    .A(_03732_),
    .B(_00169_));
 sg13g2_o21ai_1 _12695_ (.B1(_03737_),
    .Y(_00460_),
    .A1(net198),
    .A2(_03732_));
 sg13g2_buf_1 _12696_ (.A(net225),
    .X(_03738_));
 sg13g2_nand2_1 _12697_ (.Y(_03739_),
    .A(_03732_),
    .B(_00170_));
 sg13g2_o21ai_1 _12698_ (.B1(_03739_),
    .Y(_00461_),
    .A1(net197),
    .A2(_03732_));
 sg13g2_inv_1 _12699_ (.Y(_03740_),
    .A(\b.gen_square[37].sq.color ));
 sg13g2_nand2_1 _12700_ (.Y(_03741_),
    .A(_03581_),
    .B(_03695_));
 sg13g2_inv_1 _12701_ (.Y(_03742_),
    .A(_03741_));
 sg13g2_nand2_1 _12702_ (.Y(_03743_),
    .A(_03742_),
    .B(net17));
 sg13g2_buf_2 _12703_ (.A(_03743_),
    .X(_03744_));
 sg13g2_nor2_1 _12704_ (.A(net223),
    .B(_03744_),
    .Y(_03745_));
 sg13g2_a21oi_1 _12705_ (.A1(_03740_),
    .A2(_03744_),
    .Y(_00462_),
    .B1(_03745_));
 sg13g2_nand2_1 _12706_ (.Y(_03746_),
    .A(_03744_),
    .B(_00171_));
 sg13g2_o21ai_1 _12707_ (.B1(_03746_),
    .Y(_00463_),
    .A1(net199),
    .A2(_03744_));
 sg13g2_nand2_1 _12708_ (.Y(_03747_),
    .A(_03744_),
    .B(_00172_));
 sg13g2_o21ai_1 _12709_ (.B1(_03747_),
    .Y(_00464_),
    .A1(net198),
    .A2(_03744_));
 sg13g2_nand2_1 _12710_ (.Y(_03748_),
    .A(_03744_),
    .B(_00173_));
 sg13g2_o21ai_1 _12711_ (.B1(_03748_),
    .Y(_00465_),
    .A1(net197),
    .A2(_03744_));
 sg13g2_inv_1 _12712_ (.Y(_03749_),
    .A(\b.gen_square[38].sq.color ));
 sg13g2_nand2_1 _12713_ (.Y(_03750_),
    .A(_03592_),
    .B(_03695_));
 sg13g2_inv_1 _12714_ (.Y(_03751_),
    .A(_03750_));
 sg13g2_buf_1 _12715_ (.A(net24),
    .X(_03752_));
 sg13g2_nand2_1 _12716_ (.Y(_03753_),
    .A(_03751_),
    .B(net16));
 sg13g2_buf_2 _12717_ (.A(_03753_),
    .X(_03754_));
 sg13g2_buf_1 _12718_ (.A(_02188_),
    .X(_03755_));
 sg13g2_nor2_1 _12719_ (.A(net222),
    .B(_03754_),
    .Y(_03756_));
 sg13g2_a21oi_1 _12720_ (.A1(_03749_),
    .A2(_03754_),
    .Y(_00466_),
    .B1(_03756_));
 sg13g2_nand2_1 _12721_ (.Y(_03757_),
    .A(_03754_),
    .B(_00174_));
 sg13g2_o21ai_1 _12722_ (.B1(_03757_),
    .Y(_00467_),
    .A1(net199),
    .A2(_03754_));
 sg13g2_nand2_1 _12723_ (.Y(_03758_),
    .A(_03754_),
    .B(_00175_));
 sg13g2_o21ai_1 _12724_ (.B1(_03758_),
    .Y(_00468_),
    .A1(net198),
    .A2(_03754_));
 sg13g2_nand2_1 _12725_ (.Y(_03759_),
    .A(_03754_),
    .B(_00176_));
 sg13g2_o21ai_1 _12726_ (.B1(_03759_),
    .Y(_00469_),
    .A1(net197),
    .A2(_03754_));
 sg13g2_buf_1 _12727_ (.A(\b.gen_square[39].sq.color ),
    .X(_03760_));
 sg13g2_inv_1 _12728_ (.Y(_03761_),
    .A(_03760_));
 sg13g2_inv_1 _12729_ (.Y(_03762_),
    .A(_03604_));
 sg13g2_nor2_1 _12730_ (.A(net170),
    .B(_03762_),
    .Y(_03763_));
 sg13g2_nand2_1 _12731_ (.Y(_03764_),
    .A(_03763_),
    .B(net16));
 sg13g2_buf_2 _12732_ (.A(_03764_),
    .X(_03765_));
 sg13g2_nor2_1 _12733_ (.A(net222),
    .B(_03765_),
    .Y(_03766_));
 sg13g2_a21oi_1 _12734_ (.A1(_03761_),
    .A2(_03765_),
    .Y(_00470_),
    .B1(_03766_));
 sg13g2_nand2_1 _12735_ (.Y(_03767_),
    .A(_03765_),
    .B(_00177_));
 sg13g2_o21ai_1 _12736_ (.B1(_03767_),
    .Y(_00471_),
    .A1(_03734_),
    .A2(_03765_));
 sg13g2_nand2_1 _12737_ (.Y(_03768_),
    .A(_03765_),
    .B(_00178_));
 sg13g2_o21ai_1 _12738_ (.B1(_03768_),
    .Y(_00472_),
    .A1(_03736_),
    .A2(_03765_));
 sg13g2_nand2_1 _12739_ (.Y(_03769_),
    .A(_03765_),
    .B(_00179_));
 sg13g2_o21ai_1 _12740_ (.B1(_03769_),
    .Y(_00473_),
    .A1(_03738_),
    .A2(_03765_));
 sg13g2_nor2_1 _12741_ (.A(_01836_),
    .B(_03549_),
    .Y(_03770_));
 sg13g2_inv_1 _12742_ (.Y(_03771_),
    .A(_03770_));
 sg13g2_nor2_1 _12743_ (.A(_02770_),
    .B(_03771_),
    .Y(_03772_));
 sg13g2_buf_2 _12744_ (.A(_03772_),
    .X(_03773_));
 sg13g2_nor2_1 _12745_ (.A(\b.gen_square[3].sq.color ),
    .B(_03773_),
    .Y(_03774_));
 sg13g2_a21oi_1 _12746_ (.A1(_02759_),
    .A2(_03773_),
    .Y(_00474_),
    .B1(_03774_));
 sg13g2_nor2_1 _12747_ (.A(_00180_),
    .B(_03773_),
    .Y(_03775_));
 sg13g2_a21oi_1 _12748_ (.A1(_02253_),
    .A2(_03773_),
    .Y(_00475_),
    .B1(_03775_));
 sg13g2_nor2_1 _12749_ (.A(_00181_),
    .B(_03773_),
    .Y(_03776_));
 sg13g2_a21oi_1 _12750_ (.A1(net207),
    .A2(_03773_),
    .Y(_00476_),
    .B1(_03776_));
 sg13g2_nor2_1 _12751_ (.A(_00182_),
    .B(_03773_),
    .Y(_03777_));
 sg13g2_a21oi_1 _12752_ (.A1(_02361_),
    .A2(_03773_),
    .Y(_00477_),
    .B1(_03777_));
 sg13g2_inv_1 _12753_ (.Y(_03778_),
    .A(\b.gen_square[40].sq.color ));
 sg13g2_nor2_1 _12754_ (.A(net170),
    .B(_03613_),
    .Y(_03779_));
 sg13g2_nand2_1 _12755_ (.Y(_03780_),
    .A(_03779_),
    .B(net16));
 sg13g2_buf_2 _12756_ (.A(_03780_),
    .X(_03781_));
 sg13g2_nor2_1 _12757_ (.A(net222),
    .B(_03781_),
    .Y(_03782_));
 sg13g2_a21oi_1 _12758_ (.A1(_03778_),
    .A2(_03781_),
    .Y(_00478_),
    .B1(_03782_));
 sg13g2_nand2_1 _12759_ (.Y(_03783_),
    .A(_03781_),
    .B(_00183_));
 sg13g2_o21ai_1 _12760_ (.B1(_03783_),
    .Y(_00479_),
    .A1(net199),
    .A2(_03781_));
 sg13g2_nand2_1 _12761_ (.Y(_03784_),
    .A(_03781_),
    .B(_00184_));
 sg13g2_o21ai_1 _12762_ (.B1(_03784_),
    .Y(_00480_),
    .A1(net198),
    .A2(_03781_));
 sg13g2_nand2_1 _12763_ (.Y(_03785_),
    .A(_03781_),
    .B(_00185_));
 sg13g2_o21ai_1 _12764_ (.B1(_03785_),
    .Y(_00481_),
    .A1(net197),
    .A2(_03781_));
 sg13g2_inv_1 _12765_ (.Y(_03786_),
    .A(\b.gen_square[41].sq.color ));
 sg13g2_nand2_1 _12766_ (.Y(_03787_),
    .A(_03623_),
    .B(_03695_));
 sg13g2_inv_2 _12767_ (.Y(_03788_),
    .A(_03787_));
 sg13g2_nand2_1 _12768_ (.Y(_03789_),
    .A(_03788_),
    .B(net16));
 sg13g2_buf_2 _12769_ (.A(_03789_),
    .X(_03790_));
 sg13g2_nor2_1 _12770_ (.A(net222),
    .B(_03790_),
    .Y(_03791_));
 sg13g2_a21oi_1 _12771_ (.A1(_03786_),
    .A2(_03790_),
    .Y(_00482_),
    .B1(_03791_));
 sg13g2_nand2_1 _12772_ (.Y(_03792_),
    .A(_03790_),
    .B(_00186_));
 sg13g2_o21ai_1 _12773_ (.B1(_03792_),
    .Y(_00483_),
    .A1(net199),
    .A2(_03790_));
 sg13g2_nand2_1 _12774_ (.Y(_03793_),
    .A(_03790_),
    .B(_00187_));
 sg13g2_o21ai_1 _12775_ (.B1(_03793_),
    .Y(_00484_),
    .A1(net198),
    .A2(_03790_));
 sg13g2_nand2_1 _12776_ (.Y(_03794_),
    .A(_03790_),
    .B(_00188_));
 sg13g2_o21ai_1 _12777_ (.B1(_03794_),
    .Y(_00485_),
    .A1(net197),
    .A2(_03790_));
 sg13g2_inv_1 _12778_ (.Y(_03795_),
    .A(\b.gen_square[42].sq.color ));
 sg13g2_nand2_1 _12779_ (.Y(_03796_),
    .A(_02459_),
    .B(_03695_));
 sg13g2_inv_1 _12780_ (.Y(_03797_),
    .A(_03796_));
 sg13g2_nand2_1 _12781_ (.Y(_03798_),
    .A(_03797_),
    .B(net16));
 sg13g2_buf_2 _12782_ (.A(_03798_),
    .X(_03799_));
 sg13g2_nor2_1 _12783_ (.A(net222),
    .B(_03799_),
    .Y(_03800_));
 sg13g2_a21oi_1 _12784_ (.A1(_03795_),
    .A2(_03799_),
    .Y(_00486_),
    .B1(_03800_));
 sg13g2_nand2_1 _12785_ (.Y(_03801_),
    .A(_03799_),
    .B(_00189_));
 sg13g2_o21ai_1 _12786_ (.B1(_03801_),
    .Y(_00487_),
    .A1(net199),
    .A2(_03799_));
 sg13g2_nand2_1 _12787_ (.Y(_03802_),
    .A(_03799_),
    .B(_00190_));
 sg13g2_o21ai_1 _12788_ (.B1(_03802_),
    .Y(_00488_),
    .A1(net198),
    .A2(_03799_));
 sg13g2_nand2_1 _12789_ (.Y(_03803_),
    .A(_03799_),
    .B(_00191_));
 sg13g2_o21ai_1 _12790_ (.B1(_03803_),
    .Y(_00489_),
    .A1(net197),
    .A2(_03799_));
 sg13g2_inv_1 _12791_ (.Y(_03804_),
    .A(\b.gen_square[43].sq.color ));
 sg13g2_nor2_1 _12792_ (.A(net170),
    .B(_02631_),
    .Y(_03805_));
 sg13g2_nand2_1 _12793_ (.Y(_03806_),
    .A(_03805_),
    .B(net16));
 sg13g2_buf_2 _12794_ (.A(_03806_),
    .X(_03807_));
 sg13g2_nor2_1 _12795_ (.A(net222),
    .B(_03807_),
    .Y(_03808_));
 sg13g2_a21oi_1 _12796_ (.A1(_03804_),
    .A2(_03807_),
    .Y(_00490_),
    .B1(_03808_));
 sg13g2_nand2_1 _12797_ (.Y(_03809_),
    .A(_03807_),
    .B(_00192_));
 sg13g2_o21ai_1 _12798_ (.B1(_03809_),
    .Y(_00491_),
    .A1(net199),
    .A2(_03807_));
 sg13g2_nand2_1 _12799_ (.Y(_03810_),
    .A(_03807_),
    .B(_00193_));
 sg13g2_o21ai_1 _12800_ (.B1(_03810_),
    .Y(_00492_),
    .A1(net198),
    .A2(_03807_));
 sg13g2_nand2_1 _12801_ (.Y(_03811_),
    .A(_03807_),
    .B(_00194_));
 sg13g2_o21ai_1 _12802_ (.B1(_03811_),
    .Y(_00493_),
    .A1(net197),
    .A2(_03807_));
 sg13g2_inv_1 _12803_ (.Y(_03812_),
    .A(\b.gen_square[44].sq.color ));
 sg13g2_nor2_2 _12804_ (.A(_03696_),
    .B(_02803_),
    .Y(_03813_));
 sg13g2_nand2_1 _12805_ (.Y(_03814_),
    .A(_03813_),
    .B(net16));
 sg13g2_buf_2 _12806_ (.A(_03814_),
    .X(_03815_));
 sg13g2_nor2_1 _12807_ (.A(net222),
    .B(_03815_),
    .Y(_03816_));
 sg13g2_a21oi_1 _12808_ (.A1(_03812_),
    .A2(_03815_),
    .Y(_00494_),
    .B1(_03816_));
 sg13g2_nand2_1 _12809_ (.Y(_03817_),
    .A(_03815_),
    .B(_00195_));
 sg13g2_o21ai_1 _12810_ (.B1(_03817_),
    .Y(_00495_),
    .A1(net199),
    .A2(_03815_));
 sg13g2_nand2_1 _12811_ (.Y(_03818_),
    .A(_03815_),
    .B(_00196_));
 sg13g2_o21ai_1 _12812_ (.B1(_03818_),
    .Y(_00496_),
    .A1(net198),
    .A2(_03815_));
 sg13g2_nand2_1 _12813_ (.Y(_03819_),
    .A(_03815_),
    .B(_00197_));
 sg13g2_o21ai_1 _12814_ (.B1(_03819_),
    .Y(_00497_),
    .A1(net197),
    .A2(_03815_));
 sg13g2_inv_1 _12815_ (.Y(_03820_),
    .A(\b.gen_square[45].sq.color ));
 sg13g2_nor2_2 _12816_ (.A(net170),
    .B(_02983_),
    .Y(_03821_));
 sg13g2_nand2_1 _12817_ (.Y(_03822_),
    .A(_03821_),
    .B(net16));
 sg13g2_buf_2 _12818_ (.A(_03822_),
    .X(_03823_));
 sg13g2_nor2_1 _12819_ (.A(net222),
    .B(_03823_),
    .Y(_03824_));
 sg13g2_a21oi_1 _12820_ (.A1(_03820_),
    .A2(_03823_),
    .Y(_00498_),
    .B1(_03824_));
 sg13g2_nand2_1 _12821_ (.Y(_03825_),
    .A(_03823_),
    .B(_00198_));
 sg13g2_o21ai_1 _12822_ (.B1(_03825_),
    .Y(_00499_),
    .A1(_03734_),
    .A2(_03823_));
 sg13g2_nand2_1 _12823_ (.Y(_03826_),
    .A(_03823_),
    .B(_00199_));
 sg13g2_o21ai_1 _12824_ (.B1(_03826_),
    .Y(_00500_),
    .A1(_03736_),
    .A2(_03823_));
 sg13g2_nand2_1 _12825_ (.Y(_03827_),
    .A(_03823_),
    .B(_00200_));
 sg13g2_o21ai_1 _12826_ (.B1(_03827_),
    .Y(_00501_),
    .A1(_03738_),
    .A2(_03823_));
 sg13g2_inv_1 _12827_ (.Y(_03828_),
    .A(\b.gen_square[46].sq.color ));
 sg13g2_nor2_1 _12828_ (.A(_03697_),
    .B(_03110_),
    .Y(_03829_));
 sg13g2_nand2_1 _12829_ (.Y(_03830_),
    .A(_03829_),
    .B(_03752_));
 sg13g2_buf_2 _12830_ (.A(_03830_),
    .X(_03831_));
 sg13g2_nor2_1 _12831_ (.A(_03755_),
    .B(_03831_),
    .Y(_03832_));
 sg13g2_a21oi_1 _12832_ (.A1(_03828_),
    .A2(_03831_),
    .Y(_00502_),
    .B1(_03832_));
 sg13g2_buf_1 _12833_ (.A(net227),
    .X(_03833_));
 sg13g2_nand2_1 _12834_ (.Y(_03834_),
    .A(_03831_),
    .B(_00201_));
 sg13g2_o21ai_1 _12835_ (.B1(_03834_),
    .Y(_00503_),
    .A1(_03833_),
    .A2(_03831_));
 sg13g2_buf_1 _12836_ (.A(net226),
    .X(_03835_));
 sg13g2_nand2_1 _12837_ (.Y(_03836_),
    .A(_03831_),
    .B(_00202_));
 sg13g2_o21ai_1 _12838_ (.B1(_03836_),
    .Y(_00504_),
    .A1(_03835_),
    .A2(_03831_));
 sg13g2_buf_1 _12839_ (.A(net225),
    .X(_03837_));
 sg13g2_nand2_1 _12840_ (.Y(_03838_),
    .A(_03831_),
    .B(_00203_));
 sg13g2_o21ai_1 _12841_ (.B1(_03838_),
    .Y(_00505_),
    .A1(_03837_),
    .A2(_03831_));
 sg13g2_inv_1 _12842_ (.Y(_03839_),
    .A(\b.gen_square[47].sq.color ));
 sg13g2_nor2_1 _12843_ (.A(net170),
    .B(_03250_),
    .Y(_03840_));
 sg13g2_nand2_1 _12844_ (.Y(_03841_),
    .A(_03840_),
    .B(_03752_));
 sg13g2_buf_2 _12845_ (.A(_03841_),
    .X(_03842_));
 sg13g2_nor2_1 _12846_ (.A(_03755_),
    .B(_03842_),
    .Y(_03843_));
 sg13g2_a21oi_1 _12847_ (.A1(_03839_),
    .A2(_03842_),
    .Y(_00506_),
    .B1(_03843_));
 sg13g2_nand2_1 _12848_ (.Y(_03844_),
    .A(_03842_),
    .B(_00204_));
 sg13g2_o21ai_1 _12849_ (.B1(_03844_),
    .Y(_00507_),
    .A1(net196),
    .A2(_03842_));
 sg13g2_nand2_1 _12850_ (.Y(_03845_),
    .A(_03842_),
    .B(_00205_));
 sg13g2_o21ai_1 _12851_ (.B1(_03845_),
    .Y(_00508_),
    .A1(net195),
    .A2(_03842_));
 sg13g2_nand2_1 _12852_ (.Y(_03846_),
    .A(_03842_),
    .B(_00206_));
 sg13g2_o21ai_1 _12853_ (.B1(_03846_),
    .Y(_00509_),
    .A1(net194),
    .A2(_03842_));
 sg13g2_inv_1 _12854_ (.Y(_03847_),
    .A(\b.gen_square[48].sq.color ));
 sg13g2_nand2_1 _12855_ (.Y(_03848_),
    .A(_01781_),
    .B(_01792_));
 sg13g2_buf_2 _12856_ (.A(_03848_),
    .X(_03849_));
 sg13g2_nor2_1 _12857_ (.A(_03849_),
    .B(_01924_),
    .Y(_03850_));
 sg13g2_buf_1 _12858_ (.A(net24),
    .X(_03851_));
 sg13g2_nand2_1 _12859_ (.Y(_03852_),
    .A(_03850_),
    .B(net15));
 sg13g2_buf_2 _12860_ (.A(_03852_),
    .X(_03853_));
 sg13g2_buf_1 _12861_ (.A(_02188_),
    .X(_03854_));
 sg13g2_nor2_1 _12862_ (.A(net221),
    .B(_03853_),
    .Y(_03855_));
 sg13g2_a21oi_1 _12863_ (.A1(_03847_),
    .A2(_03853_),
    .Y(_00510_),
    .B1(_03855_));
 sg13g2_nand2_1 _12864_ (.Y(_03856_),
    .A(_03853_),
    .B(_00207_));
 sg13g2_o21ai_1 _12865_ (.B1(_03856_),
    .Y(_00511_),
    .A1(net196),
    .A2(_03853_));
 sg13g2_nand2_1 _12866_ (.Y(_03857_),
    .A(_03853_),
    .B(_00208_));
 sg13g2_o21ai_1 _12867_ (.B1(_03857_),
    .Y(_00512_),
    .A1(net195),
    .A2(_03853_));
 sg13g2_nand2_1 _12868_ (.Y(_03858_),
    .A(_03853_),
    .B(_00209_));
 sg13g2_o21ai_1 _12869_ (.B1(_03858_),
    .Y(_00513_),
    .A1(net194),
    .A2(_03853_));
 sg13g2_inv_1 _12870_ (.Y(_03859_),
    .A(\b.gen_square[49].sq.color ));
 sg13g2_nor2_1 _12871_ (.A(_03849_),
    .B(_03527_),
    .Y(_03860_));
 sg13g2_nand2_1 _12872_ (.Y(_03861_),
    .A(_03860_),
    .B(net15));
 sg13g2_buf_2 _12873_ (.A(_03861_),
    .X(_03862_));
 sg13g2_nor2_1 _12874_ (.A(net221),
    .B(_03862_),
    .Y(_03863_));
 sg13g2_a21oi_1 _12875_ (.A1(_03859_),
    .A2(_03862_),
    .Y(_00514_),
    .B1(_03863_));
 sg13g2_nand2_1 _12876_ (.Y(_03864_),
    .A(_03862_),
    .B(_00210_));
 sg13g2_o21ai_1 _12877_ (.B1(_03864_),
    .Y(_00515_),
    .A1(net196),
    .A2(_03862_));
 sg13g2_nand2_1 _12878_ (.Y(_03865_),
    .A(_03862_),
    .B(_00211_));
 sg13g2_o21ai_1 _12879_ (.B1(_03865_),
    .Y(_00516_),
    .A1(net195),
    .A2(_03862_));
 sg13g2_nand2_1 _12880_ (.Y(_03866_),
    .A(_03862_),
    .B(_00212_));
 sg13g2_o21ai_1 _12881_ (.B1(_03866_),
    .Y(_00517_),
    .A1(net194),
    .A2(_03862_));
 sg13g2_nor2_1 _12882_ (.A(net171),
    .B(_03571_),
    .Y(_03867_));
 sg13g2_nand2_1 _12883_ (.Y(_03868_),
    .A(_03867_),
    .B(net20));
 sg13g2_buf_2 _12884_ (.A(_03868_),
    .X(_03869_));
 sg13g2_buf_1 _12885_ (.A(\b.gen_square[4].sq.color ),
    .X(_03870_));
 sg13g2_nand2_1 _12886_ (.Y(_03871_),
    .A(_03869_),
    .B(_03870_));
 sg13g2_o21ai_1 _12887_ (.B1(_03871_),
    .Y(_00518_),
    .A1(_02759_),
    .A2(_03869_));
 sg13g2_nand2_1 _12888_ (.Y(_03872_),
    .A(_03869_),
    .B(_00213_));
 sg13g2_o21ai_1 _12889_ (.B1(_03872_),
    .Y(_00519_),
    .A1(_03833_),
    .A2(_03869_));
 sg13g2_nand2_1 _12890_ (.Y(_03873_),
    .A(_03869_),
    .B(_00214_));
 sg13g2_o21ai_1 _12891_ (.B1(_03873_),
    .Y(_00520_),
    .A1(_03835_),
    .A2(_03869_));
 sg13g2_nand2_1 _12892_ (.Y(_03874_),
    .A(_03869_),
    .B(_00215_));
 sg13g2_o21ai_1 _12893_ (.B1(_03874_),
    .Y(_00521_),
    .A1(_03837_),
    .A2(_03869_));
 sg13g2_inv_1 _12894_ (.Y(_03875_),
    .A(\b.gen_square[50].sq.color ));
 sg13g2_buf_8 _12895_ (.A(_03849_),
    .X(_03876_));
 sg13g2_nor2_2 _12896_ (.A(net181),
    .B(_03536_),
    .Y(_03877_));
 sg13g2_nand2_1 _12897_ (.Y(_03878_),
    .A(_03877_),
    .B(net15));
 sg13g2_buf_2 _12898_ (.A(_03878_),
    .X(_03879_));
 sg13g2_nor2_1 _12899_ (.A(net221),
    .B(_03879_),
    .Y(_03880_));
 sg13g2_a21oi_1 _12900_ (.A1(_03875_),
    .A2(_03879_),
    .Y(_00522_),
    .B1(_03880_));
 sg13g2_nand2_1 _12901_ (.Y(_03881_),
    .A(_03879_),
    .B(_00216_));
 sg13g2_o21ai_1 _12902_ (.B1(_03881_),
    .Y(_00523_),
    .A1(net196),
    .A2(_03879_));
 sg13g2_nand2_1 _12903_ (.Y(_03882_),
    .A(_03879_),
    .B(_00217_));
 sg13g2_o21ai_1 _12904_ (.B1(_03882_),
    .Y(_00524_),
    .A1(net195),
    .A2(_03879_));
 sg13g2_nand2_1 _12905_ (.Y(_03883_),
    .A(_03879_),
    .B(_00218_));
 sg13g2_o21ai_1 _12906_ (.B1(_03883_),
    .Y(_00525_),
    .A1(net194),
    .A2(_03879_));
 sg13g2_inv_1 _12907_ (.Y(_03884_),
    .A(\b.gen_square[51].sq.color ));
 sg13g2_nor2_1 _12908_ (.A(net181),
    .B(_03549_),
    .Y(_03885_));
 sg13g2_nand2_1 _12909_ (.Y(_03886_),
    .A(_03885_),
    .B(net15));
 sg13g2_buf_2 _12910_ (.A(_03886_),
    .X(_03887_));
 sg13g2_nor2_1 _12911_ (.A(net221),
    .B(_03887_),
    .Y(_03888_));
 sg13g2_a21oi_1 _12912_ (.A1(_03884_),
    .A2(_03887_),
    .Y(_00526_),
    .B1(_03888_));
 sg13g2_nand2_1 _12913_ (.Y(_03889_),
    .A(_03887_),
    .B(_00219_));
 sg13g2_o21ai_1 _12914_ (.B1(_03889_),
    .Y(_00527_),
    .A1(net196),
    .A2(_03887_));
 sg13g2_nand2_1 _12915_ (.Y(_03890_),
    .A(_03887_),
    .B(_00220_));
 sg13g2_o21ai_1 _12916_ (.B1(_03890_),
    .Y(_00528_),
    .A1(net195),
    .A2(_03887_));
 sg13g2_nand2_1 _12917_ (.Y(_03891_),
    .A(_03887_),
    .B(_00221_));
 sg13g2_o21ai_1 _12918_ (.B1(_03891_),
    .Y(_00529_),
    .A1(net194),
    .A2(_03887_));
 sg13g2_inv_1 _12919_ (.Y(_03892_),
    .A(\b.gen_square[52].sq.color ));
 sg13g2_nor2_2 _12920_ (.A(net181),
    .B(_03571_),
    .Y(_03893_));
 sg13g2_nand2_1 _12921_ (.Y(_03894_),
    .A(_03893_),
    .B(net15));
 sg13g2_buf_2 _12922_ (.A(_03894_),
    .X(_03895_));
 sg13g2_nor2_1 _12923_ (.A(net221),
    .B(_03895_),
    .Y(_03896_));
 sg13g2_a21oi_1 _12924_ (.A1(_03892_),
    .A2(_03895_),
    .Y(_00530_),
    .B1(_03896_));
 sg13g2_nand2_1 _12925_ (.Y(_03897_),
    .A(_03895_),
    .B(_00222_));
 sg13g2_o21ai_1 _12926_ (.B1(_03897_),
    .Y(_00531_),
    .A1(net196),
    .A2(_03895_));
 sg13g2_nand2_1 _12927_ (.Y(_03898_),
    .A(_03895_),
    .B(_00223_));
 sg13g2_o21ai_1 _12928_ (.B1(_03898_),
    .Y(_00532_),
    .A1(net195),
    .A2(_03895_));
 sg13g2_nand2_1 _12929_ (.Y(_03899_),
    .A(_03895_),
    .B(_00224_));
 sg13g2_o21ai_1 _12930_ (.B1(_03899_),
    .Y(_00533_),
    .A1(net194),
    .A2(_03895_));
 sg13g2_inv_1 _12931_ (.Y(_03900_),
    .A(\b.gen_square[53].sq.color ));
 sg13g2_inv_2 _12932_ (.Y(_03901_),
    .A(_03849_));
 sg13g2_buf_8 _12933_ (.A(_03901_),
    .X(_03902_));
 sg13g2_nand3_1 _12934_ (.B(_03581_),
    .C(net169),
    .A(net18),
    .Y(_03903_));
 sg13g2_buf_2 _12935_ (.A(_03903_),
    .X(_03904_));
 sg13g2_nor2_1 _12936_ (.A(_03854_),
    .B(_03904_),
    .Y(_03905_));
 sg13g2_a21oi_1 _12937_ (.A1(_03900_),
    .A2(_03904_),
    .Y(_00534_),
    .B1(_03905_));
 sg13g2_nand2_1 _12938_ (.Y(_03906_),
    .A(_03904_),
    .B(_00225_));
 sg13g2_o21ai_1 _12939_ (.B1(_03906_),
    .Y(_00535_),
    .A1(net196),
    .A2(_03904_));
 sg13g2_nand2_1 _12940_ (.Y(_03907_),
    .A(_03904_),
    .B(_00226_));
 sg13g2_o21ai_1 _12941_ (.B1(_03907_),
    .Y(_00536_),
    .A1(net195),
    .A2(_03904_));
 sg13g2_nand2_1 _12942_ (.Y(_03908_),
    .A(_03904_),
    .B(_00227_));
 sg13g2_o21ai_1 _12943_ (.B1(_03908_),
    .Y(_00537_),
    .A1(net194),
    .A2(_03904_));
 sg13g2_inv_1 _12944_ (.Y(_03909_),
    .A(\b.gen_square[54].sq.color ));
 sg13g2_nand3_1 _12945_ (.B(_03592_),
    .C(net169),
    .A(net18),
    .Y(_03910_));
 sg13g2_buf_2 _12946_ (.A(_03910_),
    .X(_03911_));
 sg13g2_nor2_1 _12947_ (.A(_03854_),
    .B(_03911_),
    .Y(_03912_));
 sg13g2_a21oi_1 _12948_ (.A1(_03909_),
    .A2(_03911_),
    .Y(_00538_),
    .B1(_03912_));
 sg13g2_nand2_1 _12949_ (.Y(_03913_),
    .A(_03911_),
    .B(_00228_));
 sg13g2_o21ai_1 _12950_ (.B1(_03913_),
    .Y(_00539_),
    .A1(net196),
    .A2(_03911_));
 sg13g2_nand2_1 _12951_ (.Y(_03914_),
    .A(_03911_),
    .B(_00229_));
 sg13g2_o21ai_1 _12952_ (.B1(_03914_),
    .Y(_00540_),
    .A1(net195),
    .A2(_03911_));
 sg13g2_nand2_1 _12953_ (.Y(_03915_),
    .A(_03911_),
    .B(_00230_));
 sg13g2_o21ai_1 _12954_ (.B1(_03915_),
    .Y(_00541_),
    .A1(net194),
    .A2(_03911_));
 sg13g2_inv_1 _12955_ (.Y(_03916_),
    .A(\b.gen_square[55].sq.color ));
 sg13g2_nor2_1 _12956_ (.A(net181),
    .B(_03762_),
    .Y(_03917_));
 sg13g2_nand2_1 _12957_ (.Y(_03918_),
    .A(_03917_),
    .B(_03851_));
 sg13g2_buf_2 _12958_ (.A(_03918_),
    .X(_03919_));
 sg13g2_nor2_1 _12959_ (.A(net221),
    .B(_03919_),
    .Y(_03920_));
 sg13g2_a21oi_1 _12960_ (.A1(_03916_),
    .A2(_03919_),
    .Y(_00542_),
    .B1(_03920_));
 sg13g2_buf_1 _12961_ (.A(_02231_),
    .X(_03921_));
 sg13g2_nand2_1 _12962_ (.Y(_03922_),
    .A(_03919_),
    .B(_00231_));
 sg13g2_o21ai_1 _12963_ (.B1(_03922_),
    .Y(_00543_),
    .A1(net220),
    .A2(_03919_));
 sg13g2_buf_1 _12964_ (.A(_02285_),
    .X(_03923_));
 sg13g2_nand2_1 _12965_ (.Y(_03924_),
    .A(_03919_),
    .B(_00232_));
 sg13g2_o21ai_1 _12966_ (.B1(_03924_),
    .Y(_00544_),
    .A1(net219),
    .A2(_03919_));
 sg13g2_buf_1 _12967_ (.A(_02339_),
    .X(_03925_));
 sg13g2_nand2_1 _12968_ (.Y(_03926_),
    .A(_03919_),
    .B(_00233_));
 sg13g2_o21ai_1 _12969_ (.B1(_03926_),
    .Y(_00545_),
    .A1(net218),
    .A2(_03919_));
 sg13g2_nor2_1 _12970_ (.A(net181),
    .B(_03613_),
    .Y(_03927_));
 sg13g2_nand2_1 _12971_ (.Y(_03928_),
    .A(_03927_),
    .B(_02155_));
 sg13g2_buf_2 _12972_ (.A(_03928_),
    .X(_03929_));
 sg13g2_nand2_1 _12973_ (.Y(_03930_),
    .A(_03929_),
    .B(\b.gen_square[56].sq.color ));
 sg13g2_o21ai_1 _12974_ (.B1(_03930_),
    .Y(_00546_),
    .A1(_02759_),
    .A2(_03929_));
 sg13g2_nand2_1 _12975_ (.Y(_03931_),
    .A(_03929_),
    .B(_00234_));
 sg13g2_o21ai_1 _12976_ (.B1(_03931_),
    .Y(_00547_),
    .A1(net220),
    .A2(_03929_));
 sg13g2_nand2_1 _12977_ (.Y(_03932_),
    .A(_03929_),
    .B(_00235_));
 sg13g2_o21ai_1 _12978_ (.B1(_03932_),
    .Y(_00548_),
    .A1(net219),
    .A2(_03929_));
 sg13g2_nand2_1 _12979_ (.Y(_03933_),
    .A(_03929_),
    .B(_00236_));
 sg13g2_o21ai_1 _12980_ (.B1(_03933_),
    .Y(_00549_),
    .A1(net218),
    .A2(_03929_));
 sg13g2_inv_1 _12981_ (.Y(_03934_),
    .A(\b.gen_square[57].sq.color ));
 sg13g2_nand3_1 _12982_ (.B(_03623_),
    .C(net169),
    .A(net24),
    .Y(_03935_));
 sg13g2_buf_2 _12983_ (.A(_03935_),
    .X(_03936_));
 sg13g2_nor2_1 _12984_ (.A(net221),
    .B(_03936_),
    .Y(_03937_));
 sg13g2_a21oi_1 _12985_ (.A1(_03934_),
    .A2(_03936_),
    .Y(_00550_),
    .B1(_03937_));
 sg13g2_nand2_1 _12986_ (.Y(_03938_),
    .A(_03936_),
    .B(_00237_));
 sg13g2_o21ai_1 _12987_ (.B1(_03938_),
    .Y(_00551_),
    .A1(net220),
    .A2(_03936_));
 sg13g2_nand2_1 _12988_ (.Y(_03939_),
    .A(_03936_),
    .B(_00238_));
 sg13g2_o21ai_1 _12989_ (.B1(_03939_),
    .Y(_00552_),
    .A1(net219),
    .A2(_03936_));
 sg13g2_nand2_1 _12990_ (.Y(_03940_),
    .A(_03936_),
    .B(_00239_));
 sg13g2_o21ai_1 _12991_ (.B1(_03940_),
    .Y(_00553_),
    .A1(net218),
    .A2(_03936_));
 sg13g2_inv_1 _12992_ (.Y(_03941_),
    .A(\b.gen_square[58].sq.color ));
 sg13g2_nand2_1 _12993_ (.Y(_03942_),
    .A(_02459_),
    .B(net169));
 sg13g2_inv_1 _12994_ (.Y(_03943_),
    .A(_03942_));
 sg13g2_nand2_1 _12995_ (.Y(_03944_),
    .A(_03943_),
    .B(net15));
 sg13g2_buf_2 _12996_ (.A(_03944_),
    .X(_03945_));
 sg13g2_nor2_1 _12997_ (.A(net221),
    .B(_03945_),
    .Y(_03946_));
 sg13g2_a21oi_1 _12998_ (.A1(_03941_),
    .A2(_03945_),
    .Y(_00554_),
    .B1(_03946_));
 sg13g2_nand2_1 _12999_ (.Y(_03947_),
    .A(_03945_),
    .B(_00240_));
 sg13g2_o21ai_1 _13000_ (.B1(_03947_),
    .Y(_00555_),
    .A1(net220),
    .A2(_03945_));
 sg13g2_nand2_1 _13001_ (.Y(_03948_),
    .A(_03945_),
    .B(_00241_));
 sg13g2_o21ai_1 _13002_ (.B1(_03948_),
    .Y(_00556_),
    .A1(net219),
    .A2(_03945_));
 sg13g2_nand2_1 _13003_ (.Y(_03949_),
    .A(_03945_),
    .B(_00242_));
 sg13g2_o21ai_1 _13004_ (.B1(_03949_),
    .Y(_00557_),
    .A1(net218),
    .A2(_03945_));
 sg13g2_inv_1 _13005_ (.Y(_03950_),
    .A(\b.gen_square[59].sq.color ));
 sg13g2_nor2_1 _13006_ (.A(net181),
    .B(_02631_),
    .Y(_03951_));
 sg13g2_nand2_1 _13007_ (.Y(_03952_),
    .A(_03951_),
    .B(net15));
 sg13g2_buf_2 _13008_ (.A(_03952_),
    .X(_03953_));
 sg13g2_buf_1 _13009_ (.A(_02188_),
    .X(_03954_));
 sg13g2_nor2_1 _13010_ (.A(net217),
    .B(_03953_),
    .Y(_03955_));
 sg13g2_a21oi_1 _13011_ (.A1(_03950_),
    .A2(_03953_),
    .Y(_00558_),
    .B1(_03955_));
 sg13g2_nand2_1 _13012_ (.Y(_03956_),
    .A(_03953_),
    .B(_00243_));
 sg13g2_o21ai_1 _13013_ (.B1(_03956_),
    .Y(_00559_),
    .A1(net220),
    .A2(_03953_));
 sg13g2_nand2_1 _13014_ (.Y(_03957_),
    .A(_03953_),
    .B(_00244_));
 sg13g2_o21ai_1 _13015_ (.B1(_03957_),
    .Y(_00560_),
    .A1(net219),
    .A2(_03953_));
 sg13g2_nand2_1 _13016_ (.Y(_03958_),
    .A(_03953_),
    .B(_00245_));
 sg13g2_o21ai_1 _13017_ (.B1(_03958_),
    .Y(_00561_),
    .A1(net218),
    .A2(_03953_));
 sg13g2_inv_1 _13018_ (.Y(_03959_),
    .A(\b.gen_square[5].sq.color ));
 sg13g2_nand2_1 _13019_ (.Y(_03960_),
    .A(_03581_),
    .B(_01814_));
 sg13g2_inv_1 _13020_ (.Y(_03961_),
    .A(_03960_));
 sg13g2_nand2_1 _13021_ (.Y(_03962_),
    .A(_03961_),
    .B(_03851_));
 sg13g2_buf_2 _13022_ (.A(_03962_),
    .X(_03963_));
 sg13g2_nor2_1 _13023_ (.A(net217),
    .B(_03963_),
    .Y(_03964_));
 sg13g2_a21oi_1 _13024_ (.A1(_03959_),
    .A2(_03963_),
    .Y(_00562_),
    .B1(_03964_));
 sg13g2_nand2_1 _13025_ (.Y(_03965_),
    .A(_03963_),
    .B(_00246_));
 sg13g2_o21ai_1 _13026_ (.B1(_03965_),
    .Y(_00563_),
    .A1(_03921_),
    .A2(_03963_));
 sg13g2_nand2_1 _13027_ (.Y(_03966_),
    .A(_03963_),
    .B(_00247_));
 sg13g2_o21ai_1 _13028_ (.B1(_03966_),
    .Y(_00564_),
    .A1(_03923_),
    .A2(_03963_));
 sg13g2_nand2_1 _13029_ (.Y(_03967_),
    .A(_03963_),
    .B(_00248_));
 sg13g2_o21ai_1 _13030_ (.B1(_03967_),
    .Y(_00565_),
    .A1(_03925_),
    .A2(_03963_));
 sg13g2_inv_1 _13031_ (.Y(_03968_),
    .A(\b.gen_square[60].sq.color ));
 sg13g2_nor2_1 _13032_ (.A(net181),
    .B(_02803_),
    .Y(_03969_));
 sg13g2_nand2_1 _13033_ (.Y(_03970_),
    .A(_03969_),
    .B(net15));
 sg13g2_buf_2 _13034_ (.A(_03970_),
    .X(_03971_));
 sg13g2_nor2_1 _13035_ (.A(net217),
    .B(_03971_),
    .Y(_03972_));
 sg13g2_a21oi_1 _13036_ (.A1(_03968_),
    .A2(_03971_),
    .Y(_00566_),
    .B1(_03972_));
 sg13g2_nand2_1 _13037_ (.Y(_03973_),
    .A(_03971_),
    .B(_00249_));
 sg13g2_o21ai_1 _13038_ (.B1(_03973_),
    .Y(_00567_),
    .A1(net220),
    .A2(_03971_));
 sg13g2_nand2_1 _13039_ (.Y(_03974_),
    .A(_03971_),
    .B(_00250_));
 sg13g2_o21ai_1 _13040_ (.B1(_03974_),
    .Y(_00568_),
    .A1(net219),
    .A2(_03971_));
 sg13g2_nand2_1 _13041_ (.Y(_03975_),
    .A(_03971_),
    .B(_00251_));
 sg13g2_o21ai_1 _13042_ (.B1(_03975_),
    .Y(_00569_),
    .A1(net218),
    .A2(_03971_));
 sg13g2_inv_1 _13043_ (.Y(_03976_),
    .A(\b.gen_square[61].sq.color ));
 sg13g2_nor2_1 _13044_ (.A(net181),
    .B(_02983_),
    .Y(_03977_));
 sg13g2_nand2_1 _13045_ (.Y(_03978_),
    .A(_03977_),
    .B(net18));
 sg13g2_buf_2 _13046_ (.A(_03978_),
    .X(_03979_));
 sg13g2_nor2_1 _13047_ (.A(net217),
    .B(_03979_),
    .Y(_03980_));
 sg13g2_a21oi_1 _13048_ (.A1(_03976_),
    .A2(_03979_),
    .Y(_00570_),
    .B1(_03980_));
 sg13g2_nand2_1 _13049_ (.Y(_03981_),
    .A(_03979_),
    .B(_00252_));
 sg13g2_o21ai_1 _13050_ (.B1(_03981_),
    .Y(_00571_),
    .A1(net220),
    .A2(_03979_));
 sg13g2_nand2_1 _13051_ (.Y(_03982_),
    .A(_03979_),
    .B(_00253_));
 sg13g2_o21ai_1 _13052_ (.B1(_03982_),
    .Y(_00572_),
    .A1(net219),
    .A2(_03979_));
 sg13g2_nand2_1 _13053_ (.Y(_03983_),
    .A(_03979_),
    .B(_00254_));
 sg13g2_o21ai_1 _13054_ (.B1(_03983_),
    .Y(_00573_),
    .A1(net218),
    .A2(_03979_));
 sg13g2_buf_1 _13055_ (.A(\b.gen_square[62].sq.color ),
    .X(_03984_));
 sg13g2_inv_1 _13056_ (.Y(_03985_),
    .A(_03984_));
 sg13g2_nor2_1 _13057_ (.A(_03876_),
    .B(_03110_),
    .Y(_03986_));
 sg13g2_nand2_1 _13058_ (.Y(_03987_),
    .A(_03986_),
    .B(net18));
 sg13g2_buf_2 _13059_ (.A(_03987_),
    .X(_03988_));
 sg13g2_nor2_1 _13060_ (.A(net217),
    .B(_03988_),
    .Y(_03989_));
 sg13g2_a21oi_1 _13061_ (.A1(_03985_),
    .A2(_03988_),
    .Y(_00574_),
    .B1(_03989_));
 sg13g2_nand2_1 _13062_ (.Y(_03990_),
    .A(_03988_),
    .B(_00255_));
 sg13g2_o21ai_1 _13063_ (.B1(_03990_),
    .Y(_00575_),
    .A1(net220),
    .A2(_03988_));
 sg13g2_nand2_1 _13064_ (.Y(_03991_),
    .A(_03988_),
    .B(_00256_));
 sg13g2_o21ai_1 _13065_ (.B1(_03991_),
    .Y(_00576_),
    .A1(net219),
    .A2(_03988_));
 sg13g2_nand2_1 _13066_ (.Y(_03992_),
    .A(_03988_),
    .B(_00257_));
 sg13g2_o21ai_1 _13067_ (.B1(_03992_),
    .Y(_00577_),
    .A1(net218),
    .A2(_03988_));
 sg13g2_inv_1 _13068_ (.Y(_03993_),
    .A(\b.gen_square[63].sq.color ));
 sg13g2_nor2_1 _13069_ (.A(_03876_),
    .B(_03250_),
    .Y(_03994_));
 sg13g2_nand2_1 _13070_ (.Y(_03995_),
    .A(_03994_),
    .B(net18));
 sg13g2_buf_2 _13071_ (.A(_03995_),
    .X(_03996_));
 sg13g2_nor2_1 _13072_ (.A(net217),
    .B(_03996_),
    .Y(_03997_));
 sg13g2_a21oi_1 _13073_ (.A1(_03993_),
    .A2(_03996_),
    .Y(_00578_),
    .B1(_03997_));
 sg13g2_nand2_1 _13074_ (.Y(_03998_),
    .A(_03996_),
    .B(_00258_));
 sg13g2_o21ai_1 _13075_ (.B1(_03998_),
    .Y(_00579_),
    .A1(_03921_),
    .A2(_03996_));
 sg13g2_nand2_1 _13076_ (.Y(_03999_),
    .A(_03996_),
    .B(_00259_));
 sg13g2_o21ai_1 _13077_ (.B1(_03999_),
    .Y(_00580_),
    .A1(_03923_),
    .A2(_03996_));
 sg13g2_nand2_1 _13078_ (.Y(_04000_),
    .A(_03996_),
    .B(_00260_));
 sg13g2_o21ai_1 _13079_ (.B1(_04000_),
    .Y(_00581_),
    .A1(_03925_),
    .A2(_03996_));
 sg13g2_buf_2 _13080_ (.A(\b.gen_square[6].sq.color ),
    .X(_04001_));
 sg13g2_inv_1 _13081_ (.Y(_04002_),
    .A(_04001_));
 sg13g2_nand3_1 _13082_ (.B(_01814_),
    .C(_03592_),
    .A(_02144_),
    .Y(_04003_));
 sg13g2_buf_2 _13083_ (.A(_04003_),
    .X(_04004_));
 sg13g2_nor2_1 _13084_ (.A(net217),
    .B(_04004_),
    .Y(_04005_));
 sg13g2_a21oi_1 _13085_ (.A1(_04002_),
    .A2(_04004_),
    .Y(_00582_),
    .B1(_04005_));
 sg13g2_nand2_1 _13086_ (.Y(_04006_),
    .A(_04004_),
    .B(_00261_));
 sg13g2_o21ai_1 _13087_ (.B1(_04006_),
    .Y(_00583_),
    .A1(net227),
    .A2(_04004_));
 sg13g2_nand2_1 _13088_ (.Y(_04007_),
    .A(_04004_),
    .B(_00262_));
 sg13g2_o21ai_1 _13089_ (.B1(_04007_),
    .Y(_00584_),
    .A1(net226),
    .A2(_04004_));
 sg13g2_nand2_1 _13090_ (.Y(_04008_),
    .A(_04004_),
    .B(_00263_));
 sg13g2_o21ai_1 _13091_ (.B1(_04008_),
    .Y(_00585_),
    .A1(net225),
    .A2(_04004_));
 sg13g2_buf_8 _13092_ (.A(\b.gen_square[7].sq.color ),
    .X(_04009_));
 sg13g2_inv_1 _13093_ (.Y(_04010_),
    .A(_04009_));
 sg13g2_nor2_1 _13094_ (.A(net171),
    .B(_03762_),
    .Y(_04011_));
 sg13g2_nand2_1 _13095_ (.Y(_04012_),
    .A(_04011_),
    .B(net18));
 sg13g2_buf_2 _13096_ (.A(_04012_),
    .X(_04013_));
 sg13g2_nor2_1 _13097_ (.A(net217),
    .B(_04013_),
    .Y(_04014_));
 sg13g2_a21oi_1 _13098_ (.A1(_04010_),
    .A2(_04013_),
    .Y(_00586_),
    .B1(_04014_));
 sg13g2_nand2_1 _13099_ (.Y(_04015_),
    .A(_04013_),
    .B(_00264_));
 sg13g2_o21ai_1 _13100_ (.B1(_04015_),
    .Y(_00587_),
    .A1(net227),
    .A2(_04013_));
 sg13g2_nand2_1 _13101_ (.Y(_04016_),
    .A(_04013_),
    .B(_00265_));
 sg13g2_o21ai_1 _13102_ (.B1(_04016_),
    .Y(_00588_),
    .A1(net226),
    .A2(_04013_));
 sg13g2_nand2_1 _13103_ (.Y(_04017_),
    .A(_04013_),
    .B(_00266_));
 sg13g2_o21ai_1 _13104_ (.B1(_04017_),
    .Y(_00589_),
    .A1(net225),
    .A2(_04013_));
 sg13g2_inv_1 _13105_ (.Y(_04018_),
    .A(\b.gen_square[8].sq.color ));
 sg13g2_nor2_1 _13106_ (.A(net171),
    .B(_03613_),
    .Y(_04019_));
 sg13g2_nand2_1 _13107_ (.Y(_04020_),
    .A(_04019_),
    .B(_03602_));
 sg13g2_buf_2 _13108_ (.A(_04020_),
    .X(_04021_));
 sg13g2_nor2_1 _13109_ (.A(_03954_),
    .B(_04021_),
    .Y(_04022_));
 sg13g2_a21oi_1 _13110_ (.A1(_04018_),
    .A2(_04021_),
    .Y(_00590_),
    .B1(_04022_));
 sg13g2_nand2_1 _13111_ (.Y(_04023_),
    .A(_04021_),
    .B(_00267_));
 sg13g2_o21ai_1 _13112_ (.B1(_04023_),
    .Y(_00591_),
    .A1(net227),
    .A2(_04021_));
 sg13g2_nand2_1 _13113_ (.Y(_04024_),
    .A(_04021_),
    .B(_00268_));
 sg13g2_o21ai_1 _13114_ (.B1(_04024_),
    .Y(_00592_),
    .A1(net226),
    .A2(_04021_));
 sg13g2_nand2_1 _13115_ (.Y(_04025_),
    .A(_04021_),
    .B(_00269_));
 sg13g2_o21ai_1 _13116_ (.B1(_04025_),
    .Y(_00593_),
    .A1(net225),
    .A2(_04021_));
 sg13g2_inv_1 _13117_ (.Y(_04026_),
    .A(\b.gen_square[9].sq.color ));
 sg13g2_nand2_1 _13118_ (.Y(_04027_),
    .A(_03623_),
    .B(_01814_));
 sg13g2_inv_1 _13119_ (.Y(_04028_),
    .A(_04027_));
 sg13g2_nand2_1 _13120_ (.Y(_04029_),
    .A(_04028_),
    .B(_03602_));
 sg13g2_buf_2 _13121_ (.A(_04029_),
    .X(_04030_));
 sg13g2_nor2_1 _13122_ (.A(_03954_),
    .B(_04030_),
    .Y(_04031_));
 sg13g2_a21oi_1 _13123_ (.A1(_04026_),
    .A2(_04030_),
    .Y(_00594_),
    .B1(_04031_));
 sg13g2_nand2_1 _13124_ (.Y(_04032_),
    .A(_04030_),
    .B(_00270_));
 sg13g2_o21ai_1 _13125_ (.B1(_04032_),
    .Y(_00595_),
    .A1(_02242_),
    .A2(_04030_));
 sg13g2_nand2_1 _13126_ (.Y(_04033_),
    .A(_04030_),
    .B(_00271_));
 sg13g2_o21ai_1 _13127_ (.B1(_04033_),
    .Y(_00596_),
    .A1(_02296_),
    .A2(_04030_));
 sg13g2_nand2_1 _13128_ (.Y(_04034_),
    .A(_04030_),
    .B(_00272_));
 sg13g2_o21ai_1 _13129_ (.B1(_04034_),
    .Y(_00597_),
    .A1(_02350_),
    .A2(_04030_));
 sg13g2_buf_8 _13130_ (.A(\b.gen_square[0].sq.wtm ),
    .X(_04035_));
 sg13g2_buf_8 _13131_ (.A(_04035_),
    .X(_04036_));
 sg13g2_xnor2_1 _13132_ (.Y(_04037_),
    .A(net216),
    .B(\b.gen_square[54].sq.color ));
 sg13g2_buf_1 _13133_ (.A(_04037_),
    .X(_04038_));
 sg13g2_buf_8 _13134_ (.A(net216),
    .X(_04039_));
 sg13g2_xnor2_1 _13135_ (.Y(_04040_),
    .A(net193),
    .B(\b.gen_square[45].sq.color ));
 sg13g2_buf_2 _13136_ (.A(_04040_),
    .X(_04041_));
 sg13g2_inv_1 _13137_ (.Y(_04042_),
    .A(_04041_));
 sg13g2_nor3_1 _13138_ (.A(_01968_),
    .B(_01979_),
    .C(_01946_),
    .Y(_04043_));
 sg13g2_buf_2 _13139_ (.A(_04043_),
    .X(_04044_));
 sg13g2_inv_4 _13140_ (.A(_01968_),
    .Y(_04045_));
 sg13g2_buf_8 _13141_ (.A(_04045_),
    .X(_04046_));
 sg13g2_nor3_2 _13142_ (.A(_01979_),
    .B(_01946_),
    .C(net192),
    .Y(_04047_));
 sg13g2_buf_8 _13143_ (.A(_04047_),
    .X(_04048_));
 sg13g2_nor2_1 _13144_ (.A(_04044_),
    .B(net168),
    .Y(_04049_));
 sg13g2_buf_8 _13145_ (.A(_04049_),
    .X(_04050_));
 sg13g2_buf_8 _13146_ (.A(_04050_),
    .X(_04051_));
 sg13g2_nor2_1 _13147_ (.A(_04042_),
    .B(net119),
    .Y(_04052_));
 sg13g2_buf_1 _13148_ (.A(\b.gen_square[45].sq.piece[1] ),
    .X(_04053_));
 sg13g2_inv_1 _13149_ (.Y(_04054_),
    .A(_04053_));
 sg13g2_buf_2 _13150_ (.A(\b.gen_square[45].sq.piece[2] ),
    .X(_04055_));
 sg13g2_buf_2 _13151_ (.A(\b.gen_square[45].sq.piece[0] ),
    .X(_04056_));
 sg13g2_nand3_1 _13152_ (.B(_04055_),
    .C(_04056_),
    .A(_04054_),
    .Y(_04057_));
 sg13g2_buf_1 _13153_ (.A(_04057_),
    .X(_04058_));
 sg13g2_inv_1 _13154_ (.Y(_04059_),
    .A(_04058_));
 sg13g2_nor2_1 _13155_ (.A(_04058_),
    .B(_04041_),
    .Y(_04060_));
 sg13g2_buf_8 _13156_ (.A(net168),
    .X(_04061_));
 sg13g2_nor3_1 _13157_ (.A(_01968_),
    .B(_01946_),
    .C(_01990_),
    .Y(_04062_));
 sg13g2_buf_8 _13158_ (.A(_04062_),
    .X(_04063_));
 sg13g2_buf_8 _13159_ (.A(_04063_),
    .X(_04064_));
 sg13g2_buf_8 _13160_ (.A(net167),
    .X(_04065_));
 sg13g2_a22oi_1 _13161_ (.Y(_04066_),
    .B1(net151),
    .B2(_03821_),
    .A2(net152),
    .A1(_04060_));
 sg13g2_buf_1 _13162_ (.A(_04066_),
    .X(_04067_));
 sg13g2_inv_1 _13163_ (.Y(_04068_),
    .A(_04067_));
 sg13g2_a21oi_1 _13164_ (.A1(_04052_),
    .A2(_04059_),
    .Y(_04069_),
    .B1(_04068_));
 sg13g2_buf_1 _13165_ (.A(\b.gen_square[31].sq.piece[1] ),
    .X(_04070_));
 sg13g2_inv_1 _13166_ (.Y(_04071_),
    .A(_04070_));
 sg13g2_buf_1 _13167_ (.A(\b.gen_square[31].sq.piece[2] ),
    .X(_04072_));
 sg13g2_buf_1 _13168_ (.A(\b.gen_square[31].sq.piece[0] ),
    .X(_04073_));
 sg13g2_nand3_1 _13169_ (.B(_04072_),
    .C(_04073_),
    .A(_04071_),
    .Y(_04074_));
 sg13g2_buf_1 _13170_ (.A(_04074_),
    .X(_04075_));
 sg13g2_buf_8 _13171_ (.A(net193),
    .X(_04076_));
 sg13g2_buf_8 _13172_ (.A(net179),
    .X(_04077_));
 sg13g2_buf_8 _13173_ (.A(net166),
    .X(_04078_));
 sg13g2_buf_8 _13174_ (.A(net150),
    .X(_04079_));
 sg13g2_xnor2_1 _13175_ (.Y(_04080_),
    .A(net136),
    .B(\b.gen_square[31].sq.color ));
 sg13g2_buf_1 _13176_ (.A(_04080_),
    .X(_04081_));
 sg13g2_nor2_1 _13177_ (.A(_04075_),
    .B(_04081_),
    .Y(_04082_));
 sg13g2_buf_8 _13178_ (.A(net152),
    .X(_04083_));
 sg13g2_buf_8 _13179_ (.A(net135),
    .X(_04084_));
 sg13g2_buf_8 _13180_ (.A(net118),
    .X(_04085_));
 sg13g2_buf_8 _13181_ (.A(net102),
    .X(_04086_));
 sg13g2_buf_8 _13182_ (.A(net151),
    .X(_04087_));
 sg13g2_buf_8 _13183_ (.A(net134),
    .X(_04088_));
 sg13g2_buf_8 _13184_ (.A(net117),
    .X(_04089_));
 sg13g2_buf_8 _13185_ (.A(net101),
    .X(_04090_));
 sg13g2_a22oi_1 _13186_ (.Y(_04091_),
    .B1(net91),
    .B2(_03686_),
    .A2(net92),
    .A1(_04082_));
 sg13g2_buf_1 _13187_ (.A(_04091_),
    .X(_04092_));
 sg13g2_inv_1 _13188_ (.Y(_04093_),
    .A(_04072_));
 sg13g2_nand2_1 _13189_ (.Y(_04094_),
    .A(_04070_),
    .B(_04073_));
 sg13g2_nor2_2 _13190_ (.A(_04093_),
    .B(_04094_),
    .Y(_04095_));
 sg13g2_nand2_1 _13191_ (.Y(_04096_),
    .A(_04092_),
    .B(_04095_));
 sg13g2_nand2_1 _13192_ (.Y(_04097_),
    .A(_04096_),
    .B(\b.gen_square[31].sq.color ));
 sg13g2_buf_2 _13193_ (.A(_04097_),
    .X(_04098_));
 sg13g2_buf_1 _13194_ (.A(\b.gen_square[38].sq.piece[2] ),
    .X(_04099_));
 sg13g2_inv_1 _13195_ (.Y(_04100_),
    .A(_04099_));
 sg13g2_buf_1 _13196_ (.A(\b.gen_square[38].sq.piece[1] ),
    .X(_04101_));
 sg13g2_buf_2 _13197_ (.A(\b.gen_square[38].sq.piece[0] ),
    .X(_04102_));
 sg13g2_nand2_1 _13198_ (.Y(_04103_),
    .A(_04101_),
    .B(_04102_));
 sg13g2_nor2_1 _13199_ (.A(_04100_),
    .B(_04103_),
    .Y(_04104_));
 sg13g2_inv_1 _13200_ (.Y(_04105_),
    .A(_04104_));
 sg13g2_inv_1 _13201_ (.Y(_04106_),
    .A(_04101_));
 sg13g2_nand3_1 _13202_ (.B(_04099_),
    .C(_04102_),
    .A(_04106_),
    .Y(_04107_));
 sg13g2_buf_1 _13203_ (.A(_04107_),
    .X(_04108_));
 sg13g2_xnor2_1 _13204_ (.Y(_04109_),
    .A(net150),
    .B(\b.gen_square[38].sq.color ));
 sg13g2_buf_2 _13205_ (.A(_04109_),
    .X(_04110_));
 sg13g2_nor2_1 _13206_ (.A(_04108_),
    .B(_04110_),
    .Y(_04111_));
 sg13g2_a22oi_1 _13207_ (.Y(_04112_),
    .B1(net101),
    .B2(_03751_),
    .A2(net102),
    .A1(_04111_));
 sg13g2_buf_2 _13208_ (.A(_04112_),
    .X(_04113_));
 sg13g2_inv_4 _13209_ (.A(_04113_),
    .Y(_04114_));
 sg13g2_nor2_1 _13210_ (.A(_04105_),
    .B(_04114_),
    .Y(_04115_));
 sg13g2_buf_8 _13211_ (.A(_04115_),
    .X(_04116_));
 sg13g2_buf_1 _13212_ (.A(_04116_),
    .X(_04117_));
 sg13g2_inv_1 _13213_ (.Y(_04118_),
    .A(_00035_));
 sg13g2_nor2_1 _13214_ (.A(_04118_),
    .B(_04116_),
    .Y(_04119_));
 sg13g2_buf_8 _13215_ (.A(_04119_),
    .X(_04120_));
 sg13g2_a21oi_2 _13216_ (.B1(_04120_),
    .Y(_04121_),
    .A2(net34),
    .A1(_04098_));
 sg13g2_inv_1 _13217_ (.Y(_04122_),
    .A(_04121_));
 sg13g2_inv_1 _13218_ (.Y(_04123_),
    .A(_04055_));
 sg13g2_nand2_1 _13219_ (.Y(_04124_),
    .A(_04053_),
    .B(_04056_));
 sg13g2_nor2_1 _13220_ (.A(_04123_),
    .B(_04124_),
    .Y(_04125_));
 sg13g2_nand2_1 _13221_ (.Y(_04126_),
    .A(_04067_),
    .B(_04125_));
 sg13g2_buf_2 _13222_ (.A(_04126_),
    .X(_04127_));
 sg13g2_inv_2 _13223_ (.Y(_04128_),
    .A(_04127_));
 sg13g2_buf_1 _13224_ (.A(_04128_),
    .X(_04129_));
 sg13g2_nand2_1 _13225_ (.Y(_04130_),
    .A(_04127_),
    .B(_00072_));
 sg13g2_inv_1 _13226_ (.Y(_04131_),
    .A(_04130_));
 sg13g2_a21oi_1 _13227_ (.A1(_04122_),
    .A2(net71),
    .Y(_04132_),
    .B1(_04131_));
 sg13g2_nor2_1 _13228_ (.A(_04069_),
    .B(_04132_),
    .Y(_04133_));
 sg13g2_buf_2 _13229_ (.A(_04133_),
    .X(_04134_));
 sg13g2_buf_1 _13230_ (.A(\b.gen_square[30].sq.piece[2] ),
    .X(_04135_));
 sg13g2_inv_1 _13231_ (.Y(_04136_),
    .A(_04135_));
 sg13g2_buf_2 _13232_ (.A(\b.gen_square[30].sq.piece[0] ),
    .X(_04137_));
 sg13g2_nand2_1 _13233_ (.Y(_04138_),
    .A(\b.gen_square[30].sq.piece[1] ),
    .B(_04137_));
 sg13g2_nor2_1 _13234_ (.A(_04136_),
    .B(_04138_),
    .Y(_04139_));
 sg13g2_inv_1 _13235_ (.Y(_04140_),
    .A(_04139_));
 sg13g2_inv_4 _13236_ (.A(net167),
    .Y(_04141_));
 sg13g2_inv_1 _13237_ (.Y(_04142_),
    .A(_03110_));
 sg13g2_nand2_1 _13238_ (.Y(_04143_),
    .A(_04142_),
    .B(net182));
 sg13g2_inv_1 _13239_ (.Y(_04144_),
    .A(\b.gen_square[30].sq.piece[1] ));
 sg13g2_nand3_1 _13240_ (.B(_04135_),
    .C(_04137_),
    .A(_04144_),
    .Y(_04145_));
 sg13g2_buf_1 _13241_ (.A(_04145_),
    .X(_04146_));
 sg13g2_xnor2_1 _13242_ (.Y(_04147_),
    .A(net136),
    .B(\b.gen_square[30].sq.color ));
 sg13g2_buf_2 _13243_ (.A(_04147_),
    .X(_04148_));
 sg13g2_nor2_1 _13244_ (.A(_04146_),
    .B(_04148_),
    .Y(_04149_));
 sg13g2_nand2_1 _13245_ (.Y(_04150_),
    .A(_04149_),
    .B(net92));
 sg13g2_o21ai_1 _13246_ (.B1(_04150_),
    .Y(_04151_),
    .A1(net149),
    .A2(_04143_));
 sg13g2_nor2_1 _13247_ (.A(_04140_),
    .B(_04151_),
    .Y(_04152_));
 sg13g2_buf_8 _13248_ (.A(_04152_),
    .X(_04153_));
 sg13g2_buf_1 _13249_ (.A(_04153_),
    .X(_04154_));
 sg13g2_inv_1 _13250_ (.Y(_04155_),
    .A(net33));
 sg13g2_buf_2 _13251_ (.A(\b.gen_square[6].sq.piece[2] ),
    .X(_04156_));
 sg13g2_inv_1 _13252_ (.Y(_04157_),
    .A(_04156_));
 sg13g2_buf_2 _13253_ (.A(\b.gen_square[6].sq.piece[1] ),
    .X(_04158_));
 sg13g2_buf_2 _13254_ (.A(\b.gen_square[6].sq.piece[0] ),
    .X(_04159_));
 sg13g2_nand2_1 _13255_ (.Y(_04160_),
    .A(_04158_),
    .B(_04159_));
 sg13g2_nor2_1 _13256_ (.A(_04157_),
    .B(_04160_),
    .Y(_04161_));
 sg13g2_inv_1 _13257_ (.Y(_04162_),
    .A(_04161_));
 sg13g2_inv_1 _13258_ (.Y(_04163_),
    .A(_04158_));
 sg13g2_nand3_1 _13259_ (.B(_04156_),
    .C(_04159_),
    .A(_04163_),
    .Y(_04164_));
 sg13g2_buf_2 _13260_ (.A(_04164_),
    .X(_04165_));
 sg13g2_xnor2_1 _13261_ (.Y(_04166_),
    .A(_04036_),
    .B(_04001_));
 sg13g2_buf_2 _13262_ (.A(_04166_),
    .X(_04167_));
 sg13g2_nor2_1 _13263_ (.A(_04165_),
    .B(_04167_),
    .Y(_04168_));
 sg13g2_nand2_1 _13264_ (.Y(_04169_),
    .A(_04168_),
    .B(_04048_));
 sg13g2_nand3_1 _13265_ (.B(net167),
    .C(_01814_),
    .A(_03592_),
    .Y(_04170_));
 sg13g2_nand2_1 _13266_ (.Y(_04171_),
    .A(_04169_),
    .B(_04170_));
 sg13g2_nor2_1 _13267_ (.A(_04162_),
    .B(_04171_),
    .Y(_04172_));
 sg13g2_buf_2 _13268_ (.A(_04172_),
    .X(_04173_));
 sg13g2_inv_2 _13269_ (.Y(_04174_),
    .A(_04173_));
 sg13g2_nand2_1 _13270_ (.Y(_04175_),
    .A(_04174_),
    .B(_04001_));
 sg13g2_buf_2 _13271_ (.A(_04175_),
    .X(_04176_));
 sg13g2_buf_2 _13272_ (.A(\b.gen_square[14].sq.piece[2] ),
    .X(_04177_));
 sg13g2_inv_1 _13273_ (.Y(_04178_),
    .A(_04177_));
 sg13g2_buf_1 _13274_ (.A(\b.gen_square[14].sq.piece[1] ),
    .X(_04179_));
 sg13g2_buf_2 _13275_ (.A(\b.gen_square[14].sq.piece[0] ),
    .X(_04180_));
 sg13g2_nand2_1 _13276_ (.Y(_04181_),
    .A(_04179_),
    .B(_04180_));
 sg13g2_nor2_1 _13277_ (.A(_04178_),
    .B(_04181_),
    .Y(_04182_));
 sg13g2_inv_1 _13278_ (.Y(_04183_),
    .A(_04182_));
 sg13g2_nand2_1 _13279_ (.Y(_04184_),
    .A(_03119_),
    .B(_04064_));
 sg13g2_inv_2 _13280_ (.Y(_04185_),
    .A(_04179_));
 sg13g2_nand3_1 _13281_ (.B(_04177_),
    .C(_04180_),
    .A(_04185_),
    .Y(_04186_));
 sg13g2_buf_1 _13282_ (.A(_04186_),
    .X(_04187_));
 sg13g2_xnor2_1 _13283_ (.Y(_04188_),
    .A(_04036_),
    .B(\b.gen_square[14].sq.color ));
 sg13g2_buf_2 _13284_ (.A(_04188_),
    .X(_04189_));
 sg13g2_nor2_1 _13285_ (.A(_04187_),
    .B(_04189_),
    .Y(_04190_));
 sg13g2_nand2_1 _13286_ (.Y(_04191_),
    .A(_04190_),
    .B(_04048_));
 sg13g2_nand2_1 _13287_ (.Y(_04192_),
    .A(_04184_),
    .B(_04191_));
 sg13g2_nor2_1 _13288_ (.A(_04183_),
    .B(_04192_),
    .Y(_04193_));
 sg13g2_buf_1 _13289_ (.A(_04193_),
    .X(_04194_));
 sg13g2_inv_2 _13290_ (.Y(_04195_),
    .A(net90));
 sg13g2_nand2_1 _13291_ (.Y(_04196_),
    .A(_04195_),
    .B(_00038_));
 sg13g2_inv_2 _13292_ (.Y(_04197_),
    .A(_04196_));
 sg13g2_a21oi_2 _13293_ (.B1(_04197_),
    .Y(_04198_),
    .A2(net90),
    .A1(_04176_));
 sg13g2_inv_1 _13294_ (.Y(_04199_),
    .A(_04198_));
 sg13g2_buf_1 _13295_ (.A(\b.gen_square[22].sq.piece[2] ),
    .X(_04200_));
 sg13g2_inv_1 _13296_ (.Y(_04201_),
    .A(_04200_));
 sg13g2_buf_1 _13297_ (.A(\b.gen_square[22].sq.piece[1] ),
    .X(_04202_));
 sg13g2_buf_2 _13298_ (.A(\b.gen_square[22].sq.piece[0] ),
    .X(_04203_));
 sg13g2_nand2_1 _13299_ (.Y(_04204_),
    .A(_04202_),
    .B(_04203_));
 sg13g2_nor2_1 _13300_ (.A(_04201_),
    .B(_04204_),
    .Y(_04205_));
 sg13g2_inv_1 _13301_ (.Y(_04206_),
    .A(_04205_));
 sg13g2_inv_1 _13302_ (.Y(_04207_),
    .A(_04202_));
 sg13g2_nand3_1 _13303_ (.B(_04200_),
    .C(_04203_),
    .A(_04207_),
    .Y(_04208_));
 sg13g2_buf_1 _13304_ (.A(_04208_),
    .X(_04209_));
 sg13g2_xnor2_1 _13305_ (.Y(_04210_),
    .A(net150),
    .B(\b.gen_square[22].sq.color ));
 sg13g2_buf_1 _13306_ (.A(_04210_),
    .X(_04211_));
 sg13g2_nor2_1 _13307_ (.A(_04209_),
    .B(net116),
    .Y(_04212_));
 sg13g2_nand2_1 _13308_ (.Y(_04213_),
    .A(_04212_),
    .B(net102));
 sg13g2_o21ai_1 _13309_ (.B1(_04213_),
    .Y(_04214_),
    .A1(_03593_),
    .A2(net149));
 sg13g2_nor2_1 _13310_ (.A(_04206_),
    .B(_04214_),
    .Y(_04215_));
 sg13g2_buf_1 _13311_ (.A(_04215_),
    .X(_04216_));
 sg13g2_buf_1 _13312_ (.A(net62),
    .X(_04217_));
 sg13g2_inv_1 _13313_ (.Y(_04218_),
    .A(_00037_));
 sg13g2_nor2_1 _13314_ (.A(_04218_),
    .B(net62),
    .Y(_04219_));
 sg13g2_buf_2 _13315_ (.A(_04219_),
    .X(_04220_));
 sg13g2_a21oi_1 _13316_ (.A1(_04199_),
    .A2(_04217_),
    .Y(_04221_),
    .B1(_04220_));
 sg13g2_inv_1 _13317_ (.Y(_04222_),
    .A(_00036_));
 sg13g2_nor2_1 _13318_ (.A(_04222_),
    .B(_04153_),
    .Y(_04223_));
 sg13g2_buf_8 _13319_ (.A(_04223_),
    .X(_04224_));
 sg13g2_inv_1 _13320_ (.Y(_04225_),
    .A(_04224_));
 sg13g2_o21ai_1 _13321_ (.B1(_04225_),
    .Y(_04226_),
    .A1(_04155_),
    .A2(_04221_));
 sg13g2_a21oi_1 _13322_ (.A1(_04226_),
    .A2(net34),
    .Y(_04227_),
    .B1(_04120_));
 sg13g2_inv_1 _13323_ (.Y(_04228_),
    .A(_04227_));
 sg13g2_buf_1 _13324_ (.A(\b.gen_square[46].sq.piece[2] ),
    .X(_04229_));
 sg13g2_inv_1 _13325_ (.Y(_04230_),
    .A(_04229_));
 sg13g2_buf_1 _13326_ (.A(\b.gen_square[46].sq.piece[1] ),
    .X(_04231_));
 sg13g2_buf_1 _13327_ (.A(\b.gen_square[46].sq.piece[0] ),
    .X(_04232_));
 sg13g2_nand2_1 _13328_ (.Y(_04233_),
    .A(_04231_),
    .B(_04232_));
 sg13g2_nor2_1 _13329_ (.A(_04230_),
    .B(_04233_),
    .Y(_04234_));
 sg13g2_inv_1 _13330_ (.Y(_04235_),
    .A(_04234_));
 sg13g2_nand2_1 _13331_ (.Y(_04236_),
    .A(_03829_),
    .B(net151));
 sg13g2_inv_1 _13332_ (.Y(_04237_),
    .A(_04231_));
 sg13g2_nand3_1 _13333_ (.B(_04229_),
    .C(_04232_),
    .A(_04237_),
    .Y(_04238_));
 sg13g2_buf_1 _13334_ (.A(_04238_),
    .X(_04239_));
 sg13g2_xnor2_1 _13335_ (.Y(_04240_),
    .A(net193),
    .B(\b.gen_square[46].sq.color ));
 sg13g2_buf_1 _13336_ (.A(_04240_),
    .X(_04241_));
 sg13g2_nor2_1 _13337_ (.A(_04239_),
    .B(net165),
    .Y(_04242_));
 sg13g2_buf_8 _13338_ (.A(net168),
    .X(_04243_));
 sg13g2_nand2_1 _13339_ (.Y(_04244_),
    .A(_04242_),
    .B(net148));
 sg13g2_nand2_1 _13340_ (.Y(_04245_),
    .A(_04236_),
    .B(_04244_));
 sg13g2_nor2_1 _13341_ (.A(_04235_),
    .B(_04245_),
    .Y(_04246_));
 sg13g2_buf_2 _13342_ (.A(_04246_),
    .X(_04247_));
 sg13g2_buf_1 _13343_ (.A(_04247_),
    .X(_04248_));
 sg13g2_inv_4 _13344_ (.A(_04247_),
    .Y(_04249_));
 sg13g2_nand2_1 _13345_ (.Y(_04250_),
    .A(_04249_),
    .B(_00070_));
 sg13g2_inv_1 _13346_ (.Y(_04251_),
    .A(_04250_));
 sg13g2_a21oi_1 _13347_ (.A1(_04228_),
    .A2(net82),
    .Y(_04252_),
    .B1(_04251_));
 sg13g2_buf_1 _13348_ (.A(net90),
    .X(_04253_));
 sg13g2_nand3_1 _13349_ (.B(_01957_),
    .C(_01968_),
    .A(_01990_),
    .Y(_04254_));
 sg13g2_buf_2 _13350_ (.A(_04254_),
    .X(_04255_));
 sg13g2_nor3_1 _13351_ (.A(_04165_),
    .B(_04167_),
    .C(_04255_),
    .Y(_04256_));
 sg13g2_inv_1 _13352_ (.Y(_04257_),
    .A(_04170_));
 sg13g2_nor2_1 _13353_ (.A(_04256_),
    .B(_04257_),
    .Y(_04258_));
 sg13g2_nor2_1 _13354_ (.A(_01968_),
    .B(_01979_),
    .Y(_04259_));
 sg13g2_nand2_1 _13355_ (.Y(_04260_),
    .A(_04259_),
    .B(_01957_));
 sg13g2_buf_8 _13356_ (.A(_04260_),
    .X(_04261_));
 sg13g2_nand2_1 _13357_ (.Y(_04262_),
    .A(_04255_),
    .B(_04261_));
 sg13g2_buf_8 _13358_ (.A(_04262_),
    .X(_04263_));
 sg13g2_nand3_1 _13359_ (.B(_04158_),
    .C(_04159_),
    .A(_04157_),
    .Y(_04264_));
 sg13g2_nor2_1 _13360_ (.A(_04158_),
    .B(_04159_),
    .Y(_04265_));
 sg13g2_nand2_1 _13361_ (.Y(_04266_),
    .A(_04265_),
    .B(_04156_));
 sg13g2_nand2_1 _13362_ (.Y(_04267_),
    .A(_04264_),
    .B(_04266_));
 sg13g2_nand3_1 _13363_ (.B(_04267_),
    .C(_04167_),
    .A(net147),
    .Y(_04268_));
 sg13g2_nand2_1 _13364_ (.Y(_04269_),
    .A(_04258_),
    .B(_04268_));
 sg13g2_inv_1 _13365_ (.Y(_04270_),
    .A(_04269_));
 sg13g2_inv_1 _13366_ (.Y(_04271_),
    .A(_04192_));
 sg13g2_inv_1 _13367_ (.Y(_04272_),
    .A(_04189_));
 sg13g2_nor2_1 _13368_ (.A(_04272_),
    .B(_04051_),
    .Y(_04273_));
 sg13g2_nor2_1 _13369_ (.A(_04177_),
    .B(_04181_),
    .Y(_04274_));
 sg13g2_nor2_1 _13370_ (.A(_04179_),
    .B(_04180_),
    .Y(_04275_));
 sg13g2_nand2_1 _13371_ (.Y(_04276_),
    .A(_04275_),
    .B(_04177_));
 sg13g2_nand2b_1 _13372_ (.Y(_04277_),
    .B(_04276_),
    .A_N(_04274_));
 sg13g2_nand2_1 _13373_ (.Y(_04278_),
    .A(_04273_),
    .B(_04277_));
 sg13g2_nand3_1 _13374_ (.B(_04183_),
    .C(_04278_),
    .A(_04271_),
    .Y(_04279_));
 sg13g2_inv_1 _13375_ (.Y(_04280_),
    .A(_04279_));
 sg13g2_a21oi_2 _13376_ (.B1(_04280_),
    .Y(_04281_),
    .A2(_04270_),
    .A1(net81));
 sg13g2_inv_1 _13377_ (.Y(_04282_),
    .A(_04281_));
 sg13g2_a22oi_1 _13378_ (.Y(_04283_),
    .B1(net91),
    .B2(_03594_),
    .A2(net92),
    .A1(_04212_));
 sg13g2_inv_1 _13379_ (.Y(_04284_),
    .A(net116));
 sg13g2_buf_8 _13380_ (.A(net119),
    .X(_04285_));
 sg13g2_buf_8 _13381_ (.A(net100),
    .X(_04286_));
 sg13g2_buf_8 _13382_ (.A(net89),
    .X(_04287_));
 sg13g2_nor2_1 _13383_ (.A(_04284_),
    .B(net80),
    .Y(_04288_));
 sg13g2_nor2_1 _13384_ (.A(_04200_),
    .B(_04204_),
    .Y(_04289_));
 sg13g2_nor2_1 _13385_ (.A(_04202_),
    .B(_04203_),
    .Y(_04290_));
 sg13g2_nand2_1 _13386_ (.Y(_04291_),
    .A(_04290_),
    .B(_04200_));
 sg13g2_nand2b_1 _13387_ (.Y(_04292_),
    .B(_04291_),
    .A_N(_04289_));
 sg13g2_nand2_1 _13388_ (.Y(_04293_),
    .A(_04288_),
    .B(_04292_));
 sg13g2_nand3_1 _13389_ (.B(_04206_),
    .C(_04293_),
    .A(_04283_),
    .Y(_04294_));
 sg13g2_inv_2 _13390_ (.Y(_04295_),
    .A(_04294_));
 sg13g2_a21oi_1 _13391_ (.A1(_04282_),
    .A2(net47),
    .Y(_04296_),
    .B1(_04295_));
 sg13g2_inv_1 _13392_ (.Y(_04297_),
    .A(_04296_));
 sg13g2_a22oi_1 _13393_ (.Y(_04298_),
    .B1(_03678_),
    .B2(net91),
    .A2(net92),
    .A1(_04149_));
 sg13g2_inv_1 _13394_ (.Y(_04299_),
    .A(_04148_));
 sg13g2_buf_8 _13395_ (.A(net80),
    .X(_04300_));
 sg13g2_nor2_1 _13396_ (.A(_04299_),
    .B(net70),
    .Y(_04301_));
 sg13g2_inv_1 _13397_ (.Y(_04302_),
    .A(_04138_));
 sg13g2_nand2_1 _13398_ (.Y(_04303_),
    .A(_04302_),
    .B(_04136_));
 sg13g2_nor2_1 _13399_ (.A(\b.gen_square[30].sq.piece[1] ),
    .B(_04137_),
    .Y(_04304_));
 sg13g2_nand2_1 _13400_ (.Y(_04305_),
    .A(_04304_),
    .B(_04135_));
 sg13g2_nand2_1 _13401_ (.Y(_04306_),
    .A(_04303_),
    .B(_04305_));
 sg13g2_nand2_1 _13402_ (.Y(_04307_),
    .A(_04301_),
    .B(_04306_));
 sg13g2_nand2_1 _13403_ (.Y(_04308_),
    .A(_04298_),
    .B(_04307_));
 sg13g2_nor2_1 _13404_ (.A(_04139_),
    .B(_04308_),
    .Y(_04309_));
 sg13g2_a21oi_1 _13405_ (.A1(_04297_),
    .A2(net33),
    .Y(_04310_),
    .B1(_04309_));
 sg13g2_inv_1 _13406_ (.Y(_04311_),
    .A(_04310_));
 sg13g2_inv_1 _13407_ (.Y(_04312_),
    .A(_04110_));
 sg13g2_buf_8 _13408_ (.A(net89),
    .X(_04313_));
 sg13g2_nor2_1 _13409_ (.A(_04312_),
    .B(net79),
    .Y(_04314_));
 sg13g2_nor2_1 _13410_ (.A(_04099_),
    .B(_04103_),
    .Y(_04315_));
 sg13g2_inv_1 _13411_ (.Y(_04316_),
    .A(_04315_));
 sg13g2_nor2_1 _13412_ (.A(_04101_),
    .B(_04102_),
    .Y(_04317_));
 sg13g2_nand2_1 _13413_ (.Y(_04318_),
    .A(_04317_),
    .B(_04099_));
 sg13g2_nand2_1 _13414_ (.Y(_04319_),
    .A(_04316_),
    .B(_04318_));
 sg13g2_nand2_1 _13415_ (.Y(_04320_),
    .A(_04113_),
    .B(_04105_));
 sg13g2_a21oi_1 _13416_ (.A1(_04314_),
    .A2(_04319_),
    .Y(_04321_),
    .B1(_04320_));
 sg13g2_a21oi_1 _13417_ (.A1(_04311_),
    .A2(net34),
    .Y(_04322_),
    .B1(_04321_));
 sg13g2_inv_1 _13418_ (.Y(_04323_),
    .A(_04322_));
 sg13g2_inv_1 _13419_ (.Y(_04324_),
    .A(_04245_));
 sg13g2_inv_1 _13420_ (.Y(_04325_),
    .A(net165));
 sg13g2_nor2_1 _13421_ (.A(_04325_),
    .B(net119),
    .Y(_04326_));
 sg13g2_nor2_1 _13422_ (.A(_04229_),
    .B(_04233_),
    .Y(_04327_));
 sg13g2_nor2_1 _13423_ (.A(_04231_),
    .B(_04232_),
    .Y(_04328_));
 sg13g2_nand2_1 _13424_ (.Y(_04329_),
    .A(_04328_),
    .B(_04229_));
 sg13g2_nand2b_1 _13425_ (.Y(_04330_),
    .B(_04329_),
    .A_N(_04327_));
 sg13g2_nand2_1 _13426_ (.Y(_04331_),
    .A(_04326_),
    .B(_04330_));
 sg13g2_nand3_1 _13427_ (.B(_04235_),
    .C(_04331_),
    .A(_04324_),
    .Y(_04332_));
 sg13g2_inv_1 _13428_ (.Y(_04333_),
    .A(_04332_));
 sg13g2_a21oi_1 _13429_ (.A1(_04323_),
    .A2(net82),
    .Y(_04334_),
    .B1(_04333_));
 sg13g2_inv_1 _13430_ (.Y(_04335_),
    .A(_04334_));
 sg13g2_buf_2 _13431_ (.A(\b.gen_square[55].sq.piece[1] ),
    .X(_04336_));
 sg13g2_buf_2 _13432_ (.A(\b.gen_square[55].sq.piece[2] ),
    .X(_04337_));
 sg13g2_inv_1 _13433_ (.Y(_04338_),
    .A(_04337_));
 sg13g2_buf_1 _13434_ (.A(\b.gen_square[55].sq.piece[0] ),
    .X(_04339_));
 sg13g2_inv_1 _13435_ (.Y(_04340_),
    .A(_04339_));
 sg13g2_nor3_2 _13436_ (.A(_04336_),
    .B(_04338_),
    .C(_04340_),
    .Y(_04341_));
 sg13g2_xor2_1 _13437_ (.B(\b.gen_square[55].sq.color ),
    .A(net179),
    .X(_04342_));
 sg13g2_buf_2 _13438_ (.A(_04342_),
    .X(_04343_));
 sg13g2_nand3_1 _13439_ (.B(_04343_),
    .C(net148),
    .A(_04341_),
    .Y(_04344_));
 sg13g2_nand3_1 _13440_ (.B(net167),
    .C(net169),
    .A(_03604_),
    .Y(_04345_));
 sg13g2_nand2_1 _13441_ (.Y(_04346_),
    .A(_04344_),
    .B(_04345_));
 sg13g2_buf_8 _13442_ (.A(net70),
    .X(_04347_));
 sg13g2_buf_8 _13443_ (.A(net61),
    .X(_04348_));
 sg13g2_nand2_1 _13444_ (.Y(_04349_),
    .A(_04336_),
    .B(_04339_));
 sg13g2_nor2_1 _13445_ (.A(_04337_),
    .B(_04349_),
    .Y(_04350_));
 sg13g2_nor2_1 _13446_ (.A(_04336_),
    .B(_04339_),
    .Y(_04351_));
 sg13g2_nand2_1 _13447_ (.Y(_04352_),
    .A(_04351_),
    .B(_04337_));
 sg13g2_inv_1 _13448_ (.Y(_04353_),
    .A(_04352_));
 sg13g2_nor2_1 _13449_ (.A(_04350_),
    .B(_04353_),
    .Y(_04354_));
 sg13g2_nor3_1 _13450_ (.A(_04343_),
    .B(net46),
    .C(_04354_),
    .Y(_04355_));
 sg13g2_nor2_1 _13451_ (.A(_04346_),
    .B(_04355_),
    .Y(_04356_));
 sg13g2_inv_1 _13452_ (.Y(_04357_),
    .A(_04356_));
 sg13g2_nand2_1 _13453_ (.Y(_04358_),
    .A(_04357_),
    .B(_03916_));
 sg13g2_o21ai_1 _13454_ (.B1(_04358_),
    .Y(_04359_),
    .A1(_04252_),
    .A2(_04335_));
 sg13g2_xnor2_1 _13455_ (.Y(_04360_),
    .A(net136),
    .B(\b.gen_square[61].sq.color ));
 sg13g2_buf_2 _13456_ (.A(_04360_),
    .X(_04361_));
 sg13g2_inv_1 _13457_ (.Y(_04362_),
    .A(_04361_));
 sg13g2_buf_1 _13458_ (.A(\b.gen_square[61].sq.piece[1] ),
    .X(_04363_));
 sg13g2_buf_1 _13459_ (.A(\b.gen_square[61].sq.piece[2] ),
    .X(_04364_));
 sg13g2_inv_1 _13460_ (.Y(_04365_),
    .A(_04364_));
 sg13g2_buf_1 _13461_ (.A(\b.gen_square[61].sq.piece[0] ),
    .X(_04366_));
 sg13g2_inv_1 _13462_ (.Y(_04367_),
    .A(_04366_));
 sg13g2_nor3_1 _13463_ (.A(_04363_),
    .B(_04365_),
    .C(_04367_),
    .Y(_04368_));
 sg13g2_inv_1 _13464_ (.Y(_04369_),
    .A(_04368_));
 sg13g2_buf_1 _13465_ (.A(net46),
    .X(_04370_));
 sg13g2_nor3_1 _13466_ (.A(_04362_),
    .B(_04369_),
    .C(net32),
    .Y(_04371_));
 sg13g2_nor2_1 _13467_ (.A(_04361_),
    .B(_04369_),
    .Y(_04372_));
 sg13g2_a22oi_1 _13468_ (.Y(_04373_),
    .B1(net92),
    .B2(_04372_),
    .A2(net91),
    .A1(_03977_));
 sg13g2_inv_2 _13469_ (.Y(_04374_),
    .A(_04373_));
 sg13g2_nor2_1 _13470_ (.A(_04371_),
    .B(_04374_),
    .Y(_04375_));
 sg13g2_buf_1 _13471_ (.A(_04375_),
    .X(_04376_));
 sg13g2_nand2_1 _13472_ (.Y(_04377_),
    .A(_04363_),
    .B(_04366_));
 sg13g2_nor2_2 _13473_ (.A(_04365_),
    .B(_04377_),
    .Y(_04378_));
 sg13g2_nor2b_1 _13474_ (.A(_04374_),
    .B_N(_04378_),
    .Y(_04379_));
 sg13g2_buf_2 _13475_ (.A(_04379_),
    .X(_04380_));
 sg13g2_nor2_1 _13476_ (.A(_03976_),
    .B(_04380_),
    .Y(_04381_));
 sg13g2_buf_2 _13477_ (.A(_04381_),
    .X(_04382_));
 sg13g2_nor2_1 _13478_ (.A(_04376_),
    .B(_04382_),
    .Y(_04383_));
 sg13g2_buf_1 _13479_ (.A(\b.gen_square[47].sq.piece[1] ),
    .X(_04384_));
 sg13g2_buf_1 _13480_ (.A(\b.gen_square[47].sq.piece[2] ),
    .X(_04385_));
 sg13g2_inv_1 _13481_ (.Y(_04386_),
    .A(_04385_));
 sg13g2_buf_2 _13482_ (.A(\b.gen_square[47].sq.piece[0] ),
    .X(_04387_));
 sg13g2_inv_1 _13483_ (.Y(_04388_),
    .A(_04387_));
 sg13g2_nor3_1 _13484_ (.A(_04384_),
    .B(_04386_),
    .C(_04388_),
    .Y(_04389_));
 sg13g2_xnor2_1 _13485_ (.Y(_04390_),
    .A(net150),
    .B(\b.gen_square[47].sq.color ));
 sg13g2_buf_2 _13486_ (.A(_04390_),
    .X(_04391_));
 sg13g2_inv_2 _13487_ (.Y(_04392_),
    .A(_04391_));
 sg13g2_nor2_1 _13488_ (.A(_04392_),
    .B(net32),
    .Y(_04393_));
 sg13g2_inv_1 _13489_ (.Y(_04394_),
    .A(_04389_));
 sg13g2_nor2_1 _13490_ (.A(_04391_),
    .B(_04394_),
    .Y(_04395_));
 sg13g2_inv_1 _13491_ (.Y(_04396_),
    .A(_03840_));
 sg13g2_nor2_1 _13492_ (.A(net149),
    .B(_04396_),
    .Y(_04397_));
 sg13g2_a21oi_1 _13493_ (.A1(net102),
    .A2(_04395_),
    .Y(_04398_),
    .B1(_04397_));
 sg13g2_inv_2 _13494_ (.Y(_04399_),
    .A(_04398_));
 sg13g2_a21oi_1 _13495_ (.A1(_04389_),
    .A2(_04393_),
    .Y(_04400_),
    .B1(_04399_));
 sg13g2_buf_1 _13496_ (.A(_04400_),
    .X(_04401_));
 sg13g2_nand2_1 _13497_ (.Y(_04402_),
    .A(_04384_),
    .B(_04387_));
 sg13g2_nor2_1 _13498_ (.A(_04386_),
    .B(_04402_),
    .Y(_04403_));
 sg13g2_inv_1 _13499_ (.Y(_04404_),
    .A(_04403_));
 sg13g2_nor2_1 _13500_ (.A(_04404_),
    .B(_04399_),
    .Y(_04405_));
 sg13g2_buf_2 _13501_ (.A(_04405_),
    .X(_04406_));
 sg13g2_nor2_2 _13502_ (.A(_03839_),
    .B(_04406_),
    .Y(_04407_));
 sg13g2_nor2_2 _13503_ (.A(_04401_),
    .B(_04407_),
    .Y(_04408_));
 sg13g2_nor2_1 _13504_ (.A(_04383_),
    .B(_04408_),
    .Y(_04409_));
 sg13g2_buf_1 _13505_ (.A(\b.gen_square[63].sq.piece[1] ),
    .X(_04410_));
 sg13g2_inv_1 _13506_ (.Y(_04411_),
    .A(_04410_));
 sg13g2_buf_1 _13507_ (.A(\b.gen_square[63].sq.piece[2] ),
    .X(_04412_));
 sg13g2_buf_2 _13508_ (.A(\b.gen_square[63].sq.piece[0] ),
    .X(_04413_));
 sg13g2_nand3_1 _13509_ (.B(_04412_),
    .C(_04413_),
    .A(_04411_),
    .Y(_04414_));
 sg13g2_buf_2 _13510_ (.A(_04414_),
    .X(_04415_));
 sg13g2_xnor2_1 _13511_ (.Y(_04416_),
    .A(net193),
    .B(\b.gen_square[63].sq.color ));
 sg13g2_nor2_1 _13512_ (.A(_04415_),
    .B(_04416_),
    .Y(_04417_));
 sg13g2_nand2_1 _13513_ (.Y(_04418_),
    .A(_04417_),
    .B(net148));
 sg13g2_nor2_1 _13514_ (.A(_02609_),
    .B(_02781_),
    .Y(_04419_));
 sg13g2_nand3_1 _13515_ (.B(net151),
    .C(net169),
    .A(_04419_),
    .Y(_04420_));
 sg13g2_inv_1 _13516_ (.Y(_04421_),
    .A(_04412_));
 sg13g2_nand2_1 _13517_ (.Y(_04422_),
    .A(_04410_),
    .B(_04413_));
 sg13g2_nor2_2 _13518_ (.A(_04421_),
    .B(_04422_),
    .Y(_04423_));
 sg13g2_nand3_1 _13519_ (.B(_04420_),
    .C(_04423_),
    .A(_04418_),
    .Y(_04424_));
 sg13g2_nand2b_1 _13520_ (.Y(_04425_),
    .B(_04424_),
    .A_N(_00033_));
 sg13g2_buf_2 _13521_ (.A(_04425_),
    .X(_04426_));
 sg13g2_inv_2 _13522_ (.Y(_04427_),
    .A(_04416_));
 sg13g2_nor3_1 _13523_ (.A(_04427_),
    .B(_04415_),
    .C(_04370_),
    .Y(_04428_));
 sg13g2_nand2_2 _13524_ (.Y(_04429_),
    .A(_04418_),
    .B(_04420_));
 sg13g2_inv_2 _13525_ (.Y(_04430_),
    .A(_04429_));
 sg13g2_nand2b_1 _13526_ (.Y(_04431_),
    .B(_04430_),
    .A_N(_04428_));
 sg13g2_nand2_1 _13527_ (.Y(_04432_),
    .A(_04426_),
    .B(_04431_));
 sg13g2_nor2_1 _13528_ (.A(_04343_),
    .B(net32),
    .Y(_04433_));
 sg13g2_a21oi_1 _13529_ (.A1(_04341_),
    .A2(_04433_),
    .Y(_04434_),
    .B1(_04346_));
 sg13g2_buf_1 _13530_ (.A(_04434_),
    .X(_04435_));
 sg13g2_nor2_1 _13531_ (.A(_04338_),
    .B(_04349_),
    .Y(_04436_));
 sg13g2_nand3_1 _13532_ (.B(_04345_),
    .C(_04436_),
    .A(_04344_),
    .Y(_04437_));
 sg13g2_buf_1 _13533_ (.A(_04437_),
    .X(_04438_));
 sg13g2_nand2_1 _13534_ (.Y(_04439_),
    .A(_04438_),
    .B(\b.gen_square[55].sq.color ));
 sg13g2_buf_1 _13535_ (.A(_04439_),
    .X(_04440_));
 sg13g2_inv_1 _13536_ (.Y(_04441_),
    .A(_04440_));
 sg13g2_nor2_1 _13537_ (.A(_04435_),
    .B(_04441_),
    .Y(_04442_));
 sg13g2_buf_2 _13538_ (.A(\b.gen_square[62].sq.piece[1] ),
    .X(_04443_));
 sg13g2_inv_1 _13539_ (.Y(_04444_),
    .A(_04443_));
 sg13g2_buf_2 _13540_ (.A(\b.gen_square[62].sq.piece[2] ),
    .X(_04445_));
 sg13g2_buf_2 _13541_ (.A(\b.gen_square[62].sq.piece[0] ),
    .X(_04446_));
 sg13g2_nand3_1 _13542_ (.B(_04445_),
    .C(_04446_),
    .A(_04444_),
    .Y(_04447_));
 sg13g2_buf_1 _13543_ (.A(_04447_),
    .X(_04448_));
 sg13g2_inv_1 _13544_ (.Y(_04449_),
    .A(_04448_));
 sg13g2_xnor2_1 _13545_ (.Y(_04450_),
    .A(net193),
    .B(_03984_));
 sg13g2_buf_1 _13546_ (.A(_04450_),
    .X(_04451_));
 sg13g2_inv_2 _13547_ (.Y(_04452_),
    .A(_04451_));
 sg13g2_nor2_1 _13548_ (.A(_04452_),
    .B(net46),
    .Y(_04453_));
 sg13g2_nand2_1 _13549_ (.Y(_04454_),
    .A(_03986_),
    .B(net151));
 sg13g2_nor2_1 _13550_ (.A(_04448_),
    .B(_04451_),
    .Y(_04455_));
 sg13g2_nand2_1 _13551_ (.Y(_04456_),
    .A(_04455_),
    .B(net148));
 sg13g2_nand2_1 _13552_ (.Y(_04457_),
    .A(_04454_),
    .B(_04456_));
 sg13g2_a21oi_1 _13553_ (.A1(_04449_),
    .A2(_04453_),
    .Y(_04458_),
    .B1(_04457_));
 sg13g2_buf_1 _13554_ (.A(_04458_),
    .X(_04459_));
 sg13g2_inv_1 _13555_ (.Y(_04460_),
    .A(_04445_));
 sg13g2_nand2_1 _13556_ (.Y(_04461_),
    .A(_04443_),
    .B(_04446_));
 sg13g2_nor2_2 _13557_ (.A(_04460_),
    .B(_04461_),
    .Y(_04462_));
 sg13g2_nand3_1 _13558_ (.B(_04456_),
    .C(_04462_),
    .A(_04454_),
    .Y(_04463_));
 sg13g2_buf_1 _13559_ (.A(_04463_),
    .X(_04464_));
 sg13g2_nand2_2 _13560_ (.Y(_04465_),
    .A(_04464_),
    .B(_03984_));
 sg13g2_inv_4 _13561_ (.A(_04465_),
    .Y(_04466_));
 sg13g2_nor2_1 _13562_ (.A(_04459_),
    .B(_04466_),
    .Y(_04467_));
 sg13g2_nor2_1 _13563_ (.A(_04442_),
    .B(_04467_),
    .Y(_04468_));
 sg13g2_nand3_1 _13564_ (.B(_04432_),
    .C(_04468_),
    .A(_04409_),
    .Y(_04469_));
 sg13g2_and3_1 _13565_ (.X(_04470_),
    .A(_04365_),
    .B(_04367_),
    .C(_04363_));
 sg13g2_inv_1 _13566_ (.Y(_04471_),
    .A(_04470_));
 sg13g2_nor2_1 _13567_ (.A(_04363_),
    .B(_04366_),
    .Y(_04472_));
 sg13g2_inv_1 _13568_ (.Y(_04473_),
    .A(_04472_));
 sg13g2_nor2_1 _13569_ (.A(_04365_),
    .B(_04473_),
    .Y(_04474_));
 sg13g2_inv_1 _13570_ (.Y(_04475_),
    .A(_04474_));
 sg13g2_a21oi_1 _13571_ (.A1(_04471_),
    .A2(_04475_),
    .Y(_04476_),
    .B1(net70));
 sg13g2_a21oi_1 _13572_ (.A1(_04361_),
    .A2(_04476_),
    .Y(_04477_),
    .B1(_04374_));
 sg13g2_buf_2 _13573_ (.A(_04477_),
    .X(_04478_));
 sg13g2_nor2_1 _13574_ (.A(_04478_),
    .B(_04382_),
    .Y(_04479_));
 sg13g2_inv_8 _13575_ (.Y(_04480_),
    .A(_04407_));
 sg13g2_nor2_1 _13576_ (.A(_04384_),
    .B(_04387_),
    .Y(_04481_));
 sg13g2_inv_1 _13577_ (.Y(_04482_),
    .A(_04481_));
 sg13g2_nor2_1 _13578_ (.A(_04386_),
    .B(_04482_),
    .Y(_04483_));
 sg13g2_and3_1 _13579_ (.X(_04484_),
    .A(_04386_),
    .B(_04388_),
    .C(_04384_));
 sg13g2_buf_2 _13580_ (.A(net147),
    .X(_04485_));
 sg13g2_o21ai_1 _13581_ (.B1(_04485_),
    .Y(_04486_),
    .A1(_04483_),
    .A2(_04484_));
 sg13g2_o21ai_1 _13582_ (.B1(_04398_),
    .Y(_04487_),
    .A1(_04392_),
    .A2(_04486_));
 sg13g2_nand2_1 _13583_ (.Y(_04488_),
    .A(_04480_),
    .B(_04487_));
 sg13g2_nand2b_1 _13584_ (.Y(_04489_),
    .B(_04488_),
    .A_N(_04479_));
 sg13g2_inv_1 _13585_ (.Y(_04490_),
    .A(_04457_));
 sg13g2_nor2_1 _13586_ (.A(_04443_),
    .B(_04446_),
    .Y(_04491_));
 sg13g2_nand2_1 _13587_ (.Y(_04492_),
    .A(_04491_),
    .B(_04445_));
 sg13g2_o21ai_1 _13588_ (.B1(_04492_),
    .Y(_04493_),
    .A1(_04445_),
    .A2(_04461_));
 sg13g2_nand2_1 _13589_ (.Y(_04494_),
    .A(_04453_),
    .B(_04493_));
 sg13g2_nand2_1 _13590_ (.Y(_04495_),
    .A(_04490_),
    .B(_04494_));
 sg13g2_inv_1 _13591_ (.Y(_04496_),
    .A(_04495_));
 sg13g2_nor2_1 _13592_ (.A(_03984_),
    .B(_04496_),
    .Y(_04497_));
 sg13g2_nor3_1 _13593_ (.A(_04412_),
    .B(_04413_),
    .C(_04411_),
    .Y(_04498_));
 sg13g2_nor2_1 _13594_ (.A(_04410_),
    .B(_04413_),
    .Y(_04499_));
 sg13g2_inv_1 _13595_ (.Y(_04500_),
    .A(_04499_));
 sg13g2_nor2_1 _13596_ (.A(_04421_),
    .B(_04500_),
    .Y(_04501_));
 sg13g2_nor2_1 _13597_ (.A(_04498_),
    .B(_04501_),
    .Y(_04502_));
 sg13g2_nor3_1 _13598_ (.A(_04427_),
    .B(_04050_),
    .C(_04502_),
    .Y(_04503_));
 sg13g2_nor2_1 _13599_ (.A(_04429_),
    .B(_04503_),
    .Y(_04504_));
 sg13g2_nand2b_1 _13600_ (.Y(_04505_),
    .B(_04426_),
    .A_N(_04504_));
 sg13g2_nand2b_1 _13601_ (.Y(_04506_),
    .B(_04505_),
    .A_N(_04497_));
 sg13g2_inv_1 _13602_ (.Y(_04507_),
    .A(_00029_));
 sg13g2_buf_1 _13603_ (.A(_04485_),
    .X(_04508_));
 sg13g2_buf_1 _13604_ (.A(net115),
    .X(_04509_));
 sg13g2_buf_2 _13605_ (.A(net99),
    .X(_04510_));
 sg13g2_buf_1 _13606_ (.A(net88),
    .X(_04511_));
 sg13g2_xnor2_1 _13607_ (.Y(_04512_),
    .A(net193),
    .B(\b.gen_square[44].sq.color ));
 sg13g2_buf_8 _13608_ (.A(_04512_),
    .X(_04513_));
 sg13g2_buf_2 _13609_ (.A(\b.gen_square[44].sq.piece[2] ),
    .X(_04514_));
 sg13g2_inv_1 _13610_ (.Y(_04515_),
    .A(_04514_));
 sg13g2_inv_1 _13611_ (.Y(_04516_),
    .A(\b.gen_square[44].sq.piece[1] ));
 sg13g2_buf_2 _13612_ (.A(\b.gen_square[44].sq.piece[0] ),
    .X(_04517_));
 sg13g2_nand4_1 _13613_ (.B(_04515_),
    .C(_04516_),
    .A(_04513_),
    .Y(_04518_),
    .D(_04517_));
 sg13g2_inv_1 _13614_ (.Y(_04519_),
    .A(_04518_));
 sg13g2_nand3_1 _13615_ (.B(_04514_),
    .C(_04517_),
    .A(_04516_),
    .Y(_04520_));
 sg13g2_buf_2 _13616_ (.A(_04520_),
    .X(_04521_));
 sg13g2_nor2_1 _13617_ (.A(_04521_),
    .B(_04513_),
    .Y(_04522_));
 sg13g2_a22oi_1 _13618_ (.Y(_04523_),
    .B1(_03813_),
    .B2(net167),
    .A2(net148),
    .A1(_04522_));
 sg13g2_buf_1 _13619_ (.A(_04523_),
    .X(_04524_));
 sg13g2_inv_1 _13620_ (.Y(_04525_),
    .A(_04524_));
 sg13g2_a21oi_1 _13621_ (.A1(net78),
    .A2(_04519_),
    .Y(_04526_),
    .B1(_04525_));
 sg13g2_nor2_1 _13622_ (.A(_04507_),
    .B(_04526_),
    .Y(_04527_));
 sg13g2_buf_2 _13623_ (.A(_04527_),
    .X(_04528_));
 sg13g2_inv_1 _13624_ (.Y(_04529_),
    .A(_00044_));
 sg13g2_buf_1 _13625_ (.A(_04511_),
    .X(_04530_));
 sg13g2_xnor2_1 _13626_ (.Y(_04531_),
    .A(net193),
    .B(\b.gen_square[37].sq.color ));
 sg13g2_buf_1 _13627_ (.A(_04531_),
    .X(_04532_));
 sg13g2_buf_2 _13628_ (.A(\b.gen_square[37].sq.piece[2] ),
    .X(_04533_));
 sg13g2_buf_1 _13629_ (.A(\b.gen_square[37].sq.piece[1] ),
    .X(_04534_));
 sg13g2_buf_1 _13630_ (.A(\b.gen_square[37].sq.piece[0] ),
    .X(_04535_));
 sg13g2_inv_1 _13631_ (.Y(_04536_),
    .A(_04535_));
 sg13g2_nor3_1 _13632_ (.A(_04533_),
    .B(_04534_),
    .C(_04536_),
    .Y(_04537_));
 sg13g2_nand2_1 _13633_ (.Y(_04538_),
    .A(net164),
    .B(_04537_));
 sg13g2_inv_1 _13634_ (.Y(_04539_),
    .A(_04538_));
 sg13g2_inv_1 _13635_ (.Y(_04540_),
    .A(_04534_));
 sg13g2_nand3_1 _13636_ (.B(_04533_),
    .C(_04535_),
    .A(_04540_),
    .Y(_04541_));
 sg13g2_buf_1 _13637_ (.A(_04541_),
    .X(_04542_));
 sg13g2_nor2_1 _13638_ (.A(_04542_),
    .B(net164),
    .Y(_04543_));
 sg13g2_a22oi_1 _13639_ (.Y(_04544_),
    .B1(_04065_),
    .B2(_03742_),
    .A2(net148),
    .A1(_04543_));
 sg13g2_buf_2 _13640_ (.A(_04544_),
    .X(_04545_));
 sg13g2_inv_4 _13641_ (.A(_04545_),
    .Y(_04546_));
 sg13g2_a21oi_1 _13642_ (.A1(net69),
    .A2(_04539_),
    .Y(_04547_),
    .B1(_04546_));
 sg13g2_nor2_2 _13643_ (.A(_04529_),
    .B(_04547_),
    .Y(_04548_));
 sg13g2_inv_1 _13644_ (.Y(_04549_),
    .A(_00023_));
 sg13g2_buf_1 _13645_ (.A(net69),
    .X(_04550_));
 sg13g2_xnor2_1 _13646_ (.Y(_04551_),
    .A(net136),
    .B(\b.gen_square[60].sq.color ));
 sg13g2_buf_2 _13647_ (.A(_04551_),
    .X(_04552_));
 sg13g2_buf_2 _13648_ (.A(\b.gen_square[60].sq.piece[2] ),
    .X(_04553_));
 sg13g2_buf_1 _13649_ (.A(\b.gen_square[60].sq.piece[1] ),
    .X(_04554_));
 sg13g2_buf_2 _13650_ (.A(\b.gen_square[60].sq.piece[0] ),
    .X(_04555_));
 sg13g2_inv_1 _13651_ (.Y(_04556_),
    .A(_04555_));
 sg13g2_nor3_1 _13652_ (.A(_04553_),
    .B(_04554_),
    .C(_04556_),
    .Y(_04557_));
 sg13g2_nand2_1 _13653_ (.Y(_04558_),
    .A(_04552_),
    .B(_04557_));
 sg13g2_inv_1 _13654_ (.Y(_04559_),
    .A(_04558_));
 sg13g2_inv_1 _13655_ (.Y(_04560_),
    .A(_04553_));
 sg13g2_nor3_1 _13656_ (.A(_04554_),
    .B(_04560_),
    .C(_04556_),
    .Y(_04561_));
 sg13g2_inv_1 _13657_ (.Y(_04562_),
    .A(_04561_));
 sg13g2_nor2_1 _13658_ (.A(_04552_),
    .B(_04562_),
    .Y(_04563_));
 sg13g2_a22oi_1 _13659_ (.Y(_04564_),
    .B1(net92),
    .B2(_04563_),
    .A2(net91),
    .A1(_03969_));
 sg13g2_inv_2 _13660_ (.Y(_04565_),
    .A(_04564_));
 sg13g2_a21oi_1 _13661_ (.A1(net60),
    .A2(_04559_),
    .Y(_04566_),
    .B1(_04565_));
 sg13g2_nor2_1 _13662_ (.A(_04549_),
    .B(_04566_),
    .Y(_04567_));
 sg13g2_inv_1 _13663_ (.Y(_04568_),
    .A(_00016_));
 sg13g2_xnor2_1 _13664_ (.Y(_04569_),
    .A(net136),
    .B(_03760_));
 sg13g2_buf_2 _13665_ (.A(_04569_),
    .X(_04570_));
 sg13g2_buf_1 _13666_ (.A(\b.gen_square[39].sq.piece[2] ),
    .X(_04571_));
 sg13g2_buf_1 _13667_ (.A(\b.gen_square[39].sq.piece[1] ),
    .X(_04572_));
 sg13g2_buf_1 _13668_ (.A(\b.gen_square[39].sq.piece[0] ),
    .X(_04573_));
 sg13g2_inv_1 _13669_ (.Y(_04574_),
    .A(_04573_));
 sg13g2_nor3_1 _13670_ (.A(_04571_),
    .B(_04572_),
    .C(_04574_),
    .Y(_04575_));
 sg13g2_nand2_1 _13671_ (.Y(_04576_),
    .A(_04570_),
    .B(_04575_));
 sg13g2_inv_1 _13672_ (.Y(_04577_),
    .A(_04576_));
 sg13g2_inv_1 _13673_ (.Y(_04578_),
    .A(_04572_));
 sg13g2_nand3_1 _13674_ (.B(_04571_),
    .C(_04573_),
    .A(_04578_),
    .Y(_04579_));
 sg13g2_buf_1 _13675_ (.A(_04579_),
    .X(_04580_));
 sg13g2_nor2_1 _13676_ (.A(_04580_),
    .B(_04570_),
    .Y(_04581_));
 sg13g2_a22oi_1 _13677_ (.Y(_04582_),
    .B1(net91),
    .B2(_03763_),
    .A2(net92),
    .A1(_04581_));
 sg13g2_inv_1 _13678_ (.Y(_04583_),
    .A(_04582_));
 sg13g2_a21oi_1 _13679_ (.A1(_04550_),
    .A2(_04577_),
    .Y(_04584_),
    .B1(_04583_));
 sg13g2_nor2_2 _13680_ (.A(_04568_),
    .B(_04584_),
    .Y(_04585_));
 sg13g2_or4_1 _13681_ (.A(_04528_),
    .B(_04548_),
    .C(_04567_),
    .D(_04585_),
    .X(_04586_));
 sg13g2_nor3_1 _13682_ (.A(_04489_),
    .B(_04506_),
    .C(_04586_),
    .Y(_04587_));
 sg13g2_nand2b_1 _13683_ (.Y(_04588_),
    .B(_04587_),
    .A_N(_04469_));
 sg13g2_buf_2 _13684_ (.A(\b.gen_square[48].sq.piece[2] ),
    .X(_04589_));
 sg13g2_inv_1 _13685_ (.Y(_04590_),
    .A(_04589_));
 sg13g2_buf_2 _13686_ (.A(\b.gen_square[48].sq.piece[1] ),
    .X(_04591_));
 sg13g2_buf_2 _13687_ (.A(\b.gen_square[48].sq.piece[0] ),
    .X(_04592_));
 sg13g2_nand2_1 _13688_ (.Y(_04593_),
    .A(_04591_),
    .B(_04592_));
 sg13g2_nor2_1 _13689_ (.A(_04590_),
    .B(_04593_),
    .Y(_04594_));
 sg13g2_inv_1 _13690_ (.Y(_04595_),
    .A(_04594_));
 sg13g2_inv_1 _13691_ (.Y(_04596_),
    .A(_04591_));
 sg13g2_nand3_1 _13692_ (.B(_04589_),
    .C(_04592_),
    .A(_04596_),
    .Y(_04597_));
 sg13g2_buf_1 _13693_ (.A(_04597_),
    .X(_04598_));
 sg13g2_xnor2_1 _13694_ (.Y(_04599_),
    .A(net216),
    .B(\b.gen_square[48].sq.color ));
 sg13g2_buf_8 _13695_ (.A(_04599_),
    .X(_04600_));
 sg13g2_nor2_1 _13696_ (.A(_04598_),
    .B(_04600_),
    .Y(_04601_));
 sg13g2_nand2_1 _13697_ (.Y(_04602_),
    .A(_04601_),
    .B(net168));
 sg13g2_nand2_1 _13698_ (.Y(_04603_),
    .A(_03850_),
    .B(net167));
 sg13g2_nand2_1 _13699_ (.Y(_04604_),
    .A(_04602_),
    .B(_04603_));
 sg13g2_nor2_1 _13700_ (.A(_04595_),
    .B(_04604_),
    .Y(_04605_));
 sg13g2_buf_2 _13701_ (.A(_04605_),
    .X(_04606_));
 sg13g2_nor2_1 _13702_ (.A(_03847_),
    .B(_04606_),
    .Y(_04607_));
 sg13g2_inv_1 _13703_ (.Y(_04608_),
    .A(_04607_));
 sg13g2_buf_1 _13704_ (.A(\b.gen_square[49].sq.piece[2] ),
    .X(_04609_));
 sg13g2_inv_1 _13705_ (.Y(_04610_),
    .A(_04609_));
 sg13g2_buf_2 _13706_ (.A(\b.gen_square[49].sq.piece[1] ),
    .X(_04611_));
 sg13g2_buf_1 _13707_ (.A(\b.gen_square[49].sq.piece[0] ),
    .X(_04612_));
 sg13g2_nand2_1 _13708_ (.Y(_04613_),
    .A(_04611_),
    .B(_04612_));
 sg13g2_nor2_1 _13709_ (.A(_04610_),
    .B(_04613_),
    .Y(_04614_));
 sg13g2_inv_1 _13710_ (.Y(_04615_),
    .A(_04614_));
 sg13g2_nand2_1 _13711_ (.Y(_04616_),
    .A(_03860_),
    .B(_04063_));
 sg13g2_inv_1 _13712_ (.Y(_04617_),
    .A(_04612_));
 sg13g2_nor3_1 _13713_ (.A(_04611_),
    .B(_04610_),
    .C(_04617_),
    .Y(_04618_));
 sg13g2_buf_2 _13714_ (.A(_04618_),
    .X(_04619_));
 sg13g2_xor2_1 _13715_ (.B(\b.gen_square[49].sq.color ),
    .A(net216),
    .X(_04620_));
 sg13g2_buf_2 _13716_ (.A(_04620_),
    .X(_04621_));
 sg13g2_nand3_1 _13717_ (.B(_04621_),
    .C(_04047_),
    .A(_04619_),
    .Y(_04622_));
 sg13g2_nand2_1 _13718_ (.Y(_04623_),
    .A(_04616_),
    .B(_04622_));
 sg13g2_nor2_1 _13719_ (.A(_04615_),
    .B(_04623_),
    .Y(_04624_));
 sg13g2_buf_8 _13720_ (.A(_04624_),
    .X(_04625_));
 sg13g2_buf_1 _13721_ (.A(_04625_),
    .X(_04626_));
 sg13g2_inv_4 _13722_ (.A(_04625_),
    .Y(_04627_));
 sg13g2_nand2_1 _13723_ (.Y(_04628_),
    .A(_04627_),
    .B(_00056_));
 sg13g2_inv_1 _13724_ (.Y(_04629_),
    .A(_04628_));
 sg13g2_a21oi_1 _13725_ (.A1(_04608_),
    .A2(net87),
    .Y(_04630_),
    .B1(_04629_));
 sg13g2_inv_1 _13726_ (.Y(_04631_),
    .A(_04630_));
 sg13g2_buf_2 _13727_ (.A(\b.gen_square[50].sq.piece[2] ),
    .X(_04632_));
 sg13g2_inv_1 _13728_ (.Y(_04633_),
    .A(_04632_));
 sg13g2_buf_1 _13729_ (.A(\b.gen_square[50].sq.piece[1] ),
    .X(_04634_));
 sg13g2_buf_1 _13730_ (.A(\b.gen_square[50].sq.piece[0] ),
    .X(_04635_));
 sg13g2_nand2_1 _13731_ (.Y(_04636_),
    .A(_04634_),
    .B(_04635_));
 sg13g2_nor2_1 _13732_ (.A(_04633_),
    .B(_04636_),
    .Y(_04637_));
 sg13g2_inv_1 _13733_ (.Y(_04638_),
    .A(_04637_));
 sg13g2_inv_1 _13734_ (.Y(_04639_),
    .A(_04634_));
 sg13g2_nand3_1 _13735_ (.B(_04632_),
    .C(_04635_),
    .A(_04639_),
    .Y(_04640_));
 sg13g2_buf_8 _13736_ (.A(_04640_),
    .X(_04641_));
 sg13g2_buf_8 _13737_ (.A(net179),
    .X(_04642_));
 sg13g2_xnor2_1 _13738_ (.Y(_04643_),
    .A(net163),
    .B(\b.gen_square[50].sq.color ));
 sg13g2_buf_8 _13739_ (.A(_04643_),
    .X(_04644_));
 sg13g2_nor2_1 _13740_ (.A(_04641_),
    .B(_04644_),
    .Y(_04645_));
 sg13g2_a22oi_1 _13741_ (.Y(_04646_),
    .B1(_03877_),
    .B2(net117),
    .A2(net135),
    .A1(_04645_));
 sg13g2_buf_1 _13742_ (.A(_04646_),
    .X(_04647_));
 sg13g2_inv_4 _13743_ (.A(_04647_),
    .Y(_04648_));
 sg13g2_nor2_1 _13744_ (.A(_04638_),
    .B(_04648_),
    .Y(_04649_));
 sg13g2_buf_8 _13745_ (.A(_04649_),
    .X(_04650_));
 sg13g2_buf_1 _13746_ (.A(_04650_),
    .X(_04651_));
 sg13g2_inv_1 _13747_ (.Y(_04652_),
    .A(_00049_));
 sg13g2_nor2_1 _13748_ (.A(_04652_),
    .B(_04650_),
    .Y(_04653_));
 sg13g2_buf_8 _13749_ (.A(_04653_),
    .X(_04654_));
 sg13g2_a21oi_1 _13750_ (.A1(_04631_),
    .A2(net45),
    .Y(_04655_),
    .B1(_04654_));
 sg13g2_inv_1 _13751_ (.Y(_04656_),
    .A(_04655_));
 sg13g2_buf_2 _13752_ (.A(\b.gen_square[51].sq.piece[2] ),
    .X(_04657_));
 sg13g2_inv_1 _13753_ (.Y(_04658_),
    .A(_04657_));
 sg13g2_buf_1 _13754_ (.A(\b.gen_square[51].sq.piece[1] ),
    .X(_04659_));
 sg13g2_buf_1 _13755_ (.A(\b.gen_square[51].sq.piece[0] ),
    .X(_04660_));
 sg13g2_nand2_1 _13756_ (.Y(_04661_),
    .A(_04659_),
    .B(_04660_));
 sg13g2_nor2_1 _13757_ (.A(_04658_),
    .B(_04661_),
    .Y(_04662_));
 sg13g2_inv_1 _13758_ (.Y(_04663_),
    .A(_04662_));
 sg13g2_xnor2_1 _13759_ (.Y(_04664_),
    .A(net150),
    .B(\b.gen_square[51].sq.color ));
 sg13g2_buf_2 _13760_ (.A(_04664_),
    .X(_04665_));
 sg13g2_inv_1 _13761_ (.Y(_04666_),
    .A(_04660_));
 sg13g2_nor3_2 _13762_ (.A(_04659_),
    .B(_04658_),
    .C(_04666_),
    .Y(_04667_));
 sg13g2_inv_1 _13763_ (.Y(_04668_),
    .A(_04667_));
 sg13g2_nor2_1 _13764_ (.A(_04665_),
    .B(_04668_),
    .Y(_04669_));
 sg13g2_a22oi_1 _13765_ (.Y(_04670_),
    .B1(net102),
    .B2(_04669_),
    .A2(net101),
    .A1(_03885_));
 sg13g2_buf_1 _13766_ (.A(_04670_),
    .X(_04671_));
 sg13g2_inv_2 _13767_ (.Y(_04672_),
    .A(_04671_));
 sg13g2_nor2_1 _13768_ (.A(_04663_),
    .B(_04672_),
    .Y(_04673_));
 sg13g2_buf_1 _13769_ (.A(_04673_),
    .X(_04674_));
 sg13g2_buf_1 _13770_ (.A(net44),
    .X(_04675_));
 sg13g2_inv_1 _13771_ (.Y(_04676_),
    .A(_00040_));
 sg13g2_nor2_1 _13772_ (.A(_04676_),
    .B(net44),
    .Y(_04677_));
 sg13g2_buf_2 _13773_ (.A(_04677_),
    .X(_04678_));
 sg13g2_a21oi_1 _13774_ (.A1(_04656_),
    .A2(_04675_),
    .Y(_04679_),
    .B1(_04678_));
 sg13g2_inv_1 _13775_ (.Y(_04680_),
    .A(_04679_));
 sg13g2_buf_2 _13776_ (.A(\b.gen_square[52].sq.piece[2] ),
    .X(_04681_));
 sg13g2_inv_1 _13777_ (.Y(_04682_),
    .A(_04681_));
 sg13g2_buf_1 _13778_ (.A(\b.gen_square[52].sq.piece[1] ),
    .X(_04683_));
 sg13g2_buf_1 _13779_ (.A(\b.gen_square[52].sq.piece[0] ),
    .X(_04684_));
 sg13g2_nand2_1 _13780_ (.Y(_04685_),
    .A(_04683_),
    .B(_04684_));
 sg13g2_nor2_1 _13781_ (.A(_04682_),
    .B(_04685_),
    .Y(_04686_));
 sg13g2_inv_1 _13782_ (.Y(_04687_),
    .A(_04686_));
 sg13g2_xnor2_1 _13783_ (.Y(_04688_),
    .A(net136),
    .B(\b.gen_square[52].sq.color ));
 sg13g2_buf_2 _13784_ (.A(_04688_),
    .X(_04689_));
 sg13g2_inv_1 _13785_ (.Y(_04690_),
    .A(_04684_));
 sg13g2_nor3_2 _13786_ (.A(_04683_),
    .B(_04682_),
    .C(_04690_),
    .Y(_04691_));
 sg13g2_inv_1 _13787_ (.Y(_04692_),
    .A(_04691_));
 sg13g2_nor2_1 _13788_ (.A(_04689_),
    .B(_04692_),
    .Y(_04693_));
 sg13g2_a22oi_1 _13789_ (.Y(_04694_),
    .B1(net91),
    .B2(_03893_),
    .A2(net102),
    .A1(_04693_));
 sg13g2_buf_1 _13790_ (.A(_04694_),
    .X(_04695_));
 sg13g2_inv_2 _13791_ (.Y(_04696_),
    .A(_04695_));
 sg13g2_nor2_1 _13792_ (.A(_04687_),
    .B(_04696_),
    .Y(_04697_));
 sg13g2_buf_1 _13793_ (.A(_04697_),
    .X(_04698_));
 sg13g2_buf_1 _13794_ (.A(net30),
    .X(_04699_));
 sg13g2_inv_1 _13795_ (.Y(_04700_),
    .A(_00028_));
 sg13g2_nor2_1 _13796_ (.A(_04700_),
    .B(net30),
    .Y(_04701_));
 sg13g2_buf_2 _13797_ (.A(_04701_),
    .X(_04702_));
 sg13g2_a21oi_1 _13798_ (.A1(_04680_),
    .A2(_04699_),
    .Y(_04703_),
    .B1(_04702_));
 sg13g2_inv_1 _13799_ (.Y(_04704_),
    .A(_04703_));
 sg13g2_buf_2 _13800_ (.A(\b.gen_square[53].sq.piece[2] ),
    .X(_04705_));
 sg13g2_inv_1 _13801_ (.Y(_04706_),
    .A(_04705_));
 sg13g2_buf_2 _13802_ (.A(\b.gen_square[53].sq.piece[1] ),
    .X(_04707_));
 sg13g2_buf_2 _13803_ (.A(\b.gen_square[53].sq.piece[0] ),
    .X(_04708_));
 sg13g2_nand2_1 _13804_ (.Y(_04709_),
    .A(_04707_),
    .B(_04708_));
 sg13g2_nor2_2 _13805_ (.A(_04706_),
    .B(_04709_),
    .Y(_04710_));
 sg13g2_inv_2 _13806_ (.Y(_04711_),
    .A(_04710_));
 sg13g2_nand2_1 _13807_ (.Y(_04712_),
    .A(_03581_),
    .B(_03902_));
 sg13g2_inv_1 _13808_ (.Y(_04713_),
    .A(_04707_));
 sg13g2_nand3_1 _13809_ (.B(_04705_),
    .C(_04708_),
    .A(_04713_),
    .Y(_04714_));
 sg13g2_buf_1 _13810_ (.A(_04714_),
    .X(_04715_));
 sg13g2_xnor2_1 _13811_ (.Y(_04716_),
    .A(net216),
    .B(\b.gen_square[53].sq.color ));
 sg13g2_buf_1 _13812_ (.A(_04716_),
    .X(_04717_));
 sg13g2_nor2_1 _13813_ (.A(_04715_),
    .B(net178),
    .Y(_04718_));
 sg13g2_nand2_1 _13814_ (.Y(_04719_),
    .A(_04718_),
    .B(net168));
 sg13g2_o21ai_1 _13815_ (.B1(_04719_),
    .Y(_04720_),
    .A1(_04712_),
    .A2(net149));
 sg13g2_buf_2 _13816_ (.A(_04720_),
    .X(_04721_));
 sg13g2_nor2_1 _13817_ (.A(_04711_),
    .B(_04721_),
    .Y(_04722_));
 sg13g2_buf_8 _13818_ (.A(_04722_),
    .X(_04723_));
 sg13g2_buf_1 _13819_ (.A(_04723_),
    .X(_04724_));
 sg13g2_inv_4 _13820_ (.A(_04721_),
    .Y(_04725_));
 sg13g2_nand2_1 _13821_ (.Y(_04726_),
    .A(_04725_),
    .B(_04710_));
 sg13g2_nand2_1 _13822_ (.Y(_04727_),
    .A(_04726_),
    .B(_00071_));
 sg13g2_inv_1 _13823_ (.Y(_04728_),
    .A(_04727_));
 sg13g2_a21oi_1 _13824_ (.A1(_04704_),
    .A2(_04724_),
    .Y(_04729_),
    .B1(_04728_));
 sg13g2_inv_1 _13825_ (.Y(_04730_),
    .A(_04729_));
 sg13g2_inv_1 _13826_ (.Y(_04731_),
    .A(_04604_));
 sg13g2_inv_1 _13827_ (.Y(_04732_),
    .A(_04600_));
 sg13g2_nor2_1 _13828_ (.A(_04732_),
    .B(_04050_),
    .Y(_04733_));
 sg13g2_nand3_1 _13829_ (.B(_04591_),
    .C(_04592_),
    .A(_04590_),
    .Y(_04734_));
 sg13g2_nor2_1 _13830_ (.A(_04591_),
    .B(_04592_),
    .Y(_04735_));
 sg13g2_nand2_1 _13831_ (.Y(_04736_),
    .A(_04735_),
    .B(_04589_));
 sg13g2_nand2_1 _13832_ (.Y(_04737_),
    .A(_04734_),
    .B(_04736_));
 sg13g2_nand2_1 _13833_ (.Y(_04738_),
    .A(_04733_),
    .B(_04737_));
 sg13g2_nand2_1 _13834_ (.Y(_04739_),
    .A(_04731_),
    .B(_04738_));
 sg13g2_inv_1 _13835_ (.Y(_04740_),
    .A(_04739_));
 sg13g2_nand3_1 _13836_ (.B(_03526_),
    .C(_01880_),
    .A(net169),
    .Y(_04741_));
 sg13g2_nor2_1 _13837_ (.A(net149),
    .B(_04741_),
    .Y(_04742_));
 sg13g2_nand2_1 _13838_ (.Y(_04743_),
    .A(_04619_),
    .B(_04621_));
 sg13g2_nor2_1 _13839_ (.A(_04255_),
    .B(_04743_),
    .Y(_04744_));
 sg13g2_nor2_1 _13840_ (.A(_04742_),
    .B(_04744_),
    .Y(_04745_));
 sg13g2_nor2_1 _13841_ (.A(_04621_),
    .B(_04050_),
    .Y(_04746_));
 sg13g2_inv_1 _13842_ (.Y(_04747_),
    .A(_04613_));
 sg13g2_nand2_1 _13843_ (.Y(_04748_),
    .A(_04747_),
    .B(_04610_));
 sg13g2_nor2_1 _13844_ (.A(_04611_),
    .B(_04612_),
    .Y(_04749_));
 sg13g2_nand2_1 _13845_ (.Y(_04750_),
    .A(_04749_),
    .B(_04609_));
 sg13g2_nand2_1 _13846_ (.Y(_04751_),
    .A(_04748_),
    .B(_04750_));
 sg13g2_nand2_1 _13847_ (.Y(_04752_),
    .A(_04746_),
    .B(_04751_));
 sg13g2_nand3_1 _13848_ (.B(_04752_),
    .C(_04615_),
    .A(_04745_),
    .Y(_04753_));
 sg13g2_inv_1 _13849_ (.Y(_04754_),
    .A(_04753_));
 sg13g2_a21oi_1 _13850_ (.A1(_04740_),
    .A2(net87),
    .Y(_04755_),
    .B1(_04754_));
 sg13g2_inv_1 _13851_ (.Y(_04756_),
    .A(_04755_));
 sg13g2_inv_1 _13852_ (.Y(_04757_),
    .A(_04644_));
 sg13g2_nor2_1 _13853_ (.A(_04757_),
    .B(net89),
    .Y(_04758_));
 sg13g2_nor2_1 _13854_ (.A(_04632_),
    .B(_04636_),
    .Y(_04759_));
 sg13g2_nor2_1 _13855_ (.A(_04634_),
    .B(_04635_),
    .Y(_04760_));
 sg13g2_nand2_1 _13856_ (.Y(_04761_),
    .A(_04760_),
    .B(_04632_));
 sg13g2_nand2b_1 _13857_ (.Y(_04762_),
    .B(_04761_),
    .A_N(_04759_));
 sg13g2_nand2_1 _13858_ (.Y(_04763_),
    .A(_04758_),
    .B(_04762_));
 sg13g2_nand3_1 _13859_ (.B(_04763_),
    .C(_04638_),
    .A(_04647_),
    .Y(_04764_));
 sg13g2_inv_1 _13860_ (.Y(_04765_),
    .A(_04764_));
 sg13g2_a21oi_1 _13861_ (.A1(_04756_),
    .A2(net45),
    .Y(_04766_),
    .B1(_04765_));
 sg13g2_inv_1 _13862_ (.Y(_04767_),
    .A(_04766_));
 sg13g2_inv_1 _13863_ (.Y(_04768_),
    .A(_04665_));
 sg13g2_nor2_1 _13864_ (.A(_04768_),
    .B(net70),
    .Y(_04769_));
 sg13g2_nor2_1 _13865_ (.A(_04657_),
    .B(_04661_),
    .Y(_04770_));
 sg13g2_nor2_1 _13866_ (.A(_04659_),
    .B(_04660_),
    .Y(_04771_));
 sg13g2_nand2_1 _13867_ (.Y(_04772_),
    .A(_04771_),
    .B(_04657_));
 sg13g2_nand2b_1 _13868_ (.Y(_04773_),
    .B(_04772_),
    .A_N(_04770_));
 sg13g2_nand2_1 _13869_ (.Y(_04774_),
    .A(_04769_),
    .B(_04773_));
 sg13g2_nand3_1 _13870_ (.B(_04663_),
    .C(_04774_),
    .A(_04671_),
    .Y(_04775_));
 sg13g2_inv_1 _13871_ (.Y(_04776_),
    .A(_04775_));
 sg13g2_a21oi_1 _13872_ (.A1(_04767_),
    .A2(_04675_),
    .Y(_04777_),
    .B1(_04776_));
 sg13g2_inv_1 _13873_ (.Y(_04778_),
    .A(_04777_));
 sg13g2_inv_1 _13874_ (.Y(_04779_),
    .A(_04689_));
 sg13g2_nor2_1 _13875_ (.A(_04779_),
    .B(net80),
    .Y(_04780_));
 sg13g2_nor2_1 _13876_ (.A(_04681_),
    .B(_04685_),
    .Y(_04781_));
 sg13g2_nor2_1 _13877_ (.A(_04683_),
    .B(_04684_),
    .Y(_04782_));
 sg13g2_nand2_1 _13878_ (.Y(_04783_),
    .A(_04782_),
    .B(_04681_));
 sg13g2_nand2b_1 _13879_ (.Y(_04784_),
    .B(_04783_),
    .A_N(_04781_));
 sg13g2_nand2_1 _13880_ (.Y(_04785_),
    .A(_04780_),
    .B(_04784_));
 sg13g2_nand3_1 _13881_ (.B(_04687_),
    .C(_04785_),
    .A(_04695_),
    .Y(_04786_));
 sg13g2_inv_1 _13882_ (.Y(_04787_),
    .A(_04786_));
 sg13g2_a21oi_1 _13883_ (.A1(_04778_),
    .A2(net23),
    .Y(_04788_),
    .B1(_04787_));
 sg13g2_inv_1 _13884_ (.Y(_04789_),
    .A(_04788_));
 sg13g2_nand2_1 _13885_ (.Y(_04790_),
    .A(net147),
    .B(net178));
 sg13g2_nor2_1 _13886_ (.A(_04707_),
    .B(_04708_),
    .Y(_04791_));
 sg13g2_nor2_1 _13887_ (.A(_04705_),
    .B(_04709_),
    .Y(_04792_));
 sg13g2_a21oi_1 _13888_ (.A1(_04705_),
    .A2(_04791_),
    .Y(_04793_),
    .B1(_04792_));
 sg13g2_nor2_1 _13889_ (.A(_04710_),
    .B(_04721_),
    .Y(_04794_));
 sg13g2_o21ai_1 _13890_ (.B1(_04794_),
    .Y(_04795_),
    .A1(_04790_),
    .A2(_04793_));
 sg13g2_inv_1 _13891_ (.Y(_04796_),
    .A(_04795_));
 sg13g2_a21oi_2 _13892_ (.B1(_04796_),
    .Y(_04797_),
    .A2(net77),
    .A1(_04789_));
 sg13g2_buf_2 _13893_ (.A(\b.gen_square[18].sq.piece[2] ),
    .X(_04798_));
 sg13g2_inv_1 _13894_ (.Y(_04799_),
    .A(_04798_));
 sg13g2_buf_1 _13895_ (.A(\b.gen_square[18].sq.piece[1] ),
    .X(_04800_));
 sg13g2_buf_1 _13896_ (.A(\b.gen_square[18].sq.piece[0] ),
    .X(_04801_));
 sg13g2_nand2_1 _13897_ (.Y(_04802_),
    .A(_04800_),
    .B(_04801_));
 sg13g2_nor2_1 _13898_ (.A(_04799_),
    .B(_04802_),
    .Y(_04803_));
 sg13g2_inv_1 _13899_ (.Y(_04804_),
    .A(_04803_));
 sg13g2_xnor2_1 _13900_ (.Y(_04805_),
    .A(net166),
    .B(\b.gen_square[18].sq.color ));
 sg13g2_buf_2 _13901_ (.A(_04805_),
    .X(_04806_));
 sg13g2_inv_1 _13902_ (.Y(_04807_),
    .A(_04801_));
 sg13g2_nor3_2 _13903_ (.A(_04800_),
    .B(_04799_),
    .C(_04807_),
    .Y(_04808_));
 sg13g2_inv_1 _13904_ (.Y(_04809_),
    .A(_04808_));
 sg13g2_nor2_1 _13905_ (.A(_04806_),
    .B(_04809_),
    .Y(_04810_));
 sg13g2_a22oi_1 _13906_ (.Y(_04811_),
    .B1(net118),
    .B2(_04810_),
    .A2(net101),
    .A1(_03537_));
 sg13g2_buf_1 _13907_ (.A(_04811_),
    .X(_04812_));
 sg13g2_inv_2 _13908_ (.Y(_04813_),
    .A(_04812_));
 sg13g2_nor2_1 _13909_ (.A(_04804_),
    .B(_04813_),
    .Y(_04814_));
 sg13g2_buf_2 _13910_ (.A(_04814_),
    .X(_04815_));
 sg13g2_inv_1 _13911_ (.Y(_04816_),
    .A(_04815_));
 sg13g2_buf_2 _13912_ (.A(\b.gen_square[9].sq.piece[2] ),
    .X(_04817_));
 sg13g2_inv_1 _13913_ (.Y(_04818_),
    .A(_04817_));
 sg13g2_buf_1 _13914_ (.A(\b.gen_square[9].sq.piece[1] ),
    .X(_04819_));
 sg13g2_buf_1 _13915_ (.A(\b.gen_square[9].sq.piece[0] ),
    .X(_04820_));
 sg13g2_nand2_1 _13916_ (.Y(_04821_),
    .A(_04819_),
    .B(_04820_));
 sg13g2_nor2_1 _13917_ (.A(_04818_),
    .B(_04821_),
    .Y(_04822_));
 sg13g2_inv_2 _13918_ (.Y(_04823_),
    .A(_04822_));
 sg13g2_xnor2_1 _13919_ (.Y(_04824_),
    .A(net166),
    .B(\b.gen_square[9].sq.color ));
 sg13g2_buf_1 _13920_ (.A(_04824_),
    .X(_04825_));
 sg13g2_inv_1 _13921_ (.Y(_04826_),
    .A(_04820_));
 sg13g2_nor3_2 _13922_ (.A(_04819_),
    .B(_04818_),
    .C(_04826_),
    .Y(_04827_));
 sg13g2_inv_1 _13923_ (.Y(_04828_),
    .A(_04827_));
 sg13g2_nor2_1 _13924_ (.A(net132),
    .B(_04828_),
    .Y(_04829_));
 sg13g2_a22oi_1 _13925_ (.Y(_04830_),
    .B1(net118),
    .B2(_04829_),
    .A2(net117),
    .A1(_04028_));
 sg13g2_buf_1 _13926_ (.A(_04830_),
    .X(_04831_));
 sg13g2_inv_2 _13927_ (.Y(_04832_),
    .A(_04831_));
 sg13g2_nor2_2 _13928_ (.A(_04823_),
    .B(_04832_),
    .Y(_04833_));
 sg13g2_buf_8 _13929_ (.A(_04833_),
    .X(_04834_));
 sg13g2_buf_1 _13930_ (.A(_04834_),
    .X(_04835_));
 sg13g2_buf_1 _13931_ (.A(\b.gen_square[0].sq.piece[2] ),
    .X(_04836_));
 sg13g2_inv_2 _13932_ (.Y(_04837_),
    .A(_04836_));
 sg13g2_buf_1 _13933_ (.A(\b.gen_square[0].sq.piece[1] ),
    .X(_04838_));
 sg13g2_buf_1 _13934_ (.A(\b.gen_square[0].sq.piece[0] ),
    .X(_04839_));
 sg13g2_nand2_1 _13935_ (.Y(_04840_),
    .A(_04838_),
    .B(_04839_));
 sg13g2_nor2_1 _13936_ (.A(_04837_),
    .B(_04840_),
    .Y(_04841_));
 sg13g2_xnor2_1 _13937_ (.Y(_04842_),
    .A(net163),
    .B(_01759_));
 sg13g2_buf_8 _13938_ (.A(_04842_),
    .X(_04843_));
 sg13g2_nand2b_1 _13939_ (.Y(_04844_),
    .B(net131),
    .A_N(_04841_));
 sg13g2_nor2_1 _13940_ (.A(net80),
    .B(_04844_),
    .Y(_04845_));
 sg13g2_nor2_1 _13941_ (.A(_04838_),
    .B(_04839_),
    .Y(_04846_));
 sg13g2_inv_2 _13942_ (.Y(_04847_),
    .A(_04846_));
 sg13g2_inv_1 _13943_ (.Y(_04848_),
    .A(_04839_));
 sg13g2_nand3_1 _13944_ (.B(_04848_),
    .C(_04838_),
    .A(_04837_),
    .Y(_04849_));
 sg13g2_o21ai_1 _13945_ (.B1(_04849_),
    .Y(_04850_),
    .A1(_04837_),
    .A2(_04847_));
 sg13g2_inv_1 _13946_ (.Y(_04851_),
    .A(_04838_));
 sg13g2_nand3_1 _13947_ (.B(_04836_),
    .C(_04839_),
    .A(_04851_),
    .Y(_04852_));
 sg13g2_buf_1 _13948_ (.A(_04852_),
    .X(_04853_));
 sg13g2_nor2_1 _13949_ (.A(_04853_),
    .B(net131),
    .Y(_04854_));
 sg13g2_a22oi_1 _13950_ (.Y(_04855_),
    .B1(net135),
    .B2(_04854_),
    .A2(net117),
    .A1(_01935_));
 sg13g2_buf_1 _13951_ (.A(_04855_),
    .X(_04856_));
 sg13g2_inv_1 _13952_ (.Y(_04857_),
    .A(_04856_));
 sg13g2_a21oi_1 _13953_ (.A1(_04845_),
    .A2(_04850_),
    .Y(_04858_),
    .B1(_04857_));
 sg13g2_nor2_1 _13954_ (.A(_04819_),
    .B(_04820_),
    .Y(_04859_));
 sg13g2_nand2_1 _13955_ (.Y(_04860_),
    .A(_04859_),
    .B(_04817_));
 sg13g2_inv_1 _13956_ (.Y(_04861_),
    .A(_04860_));
 sg13g2_and3_1 _13957_ (.X(_04862_),
    .A(_04818_),
    .B(_04826_),
    .C(_04819_));
 sg13g2_inv_1 _13958_ (.Y(_04863_),
    .A(net132));
 sg13g2_nor2_1 _13959_ (.A(_04863_),
    .B(net80),
    .Y(_04864_));
 sg13g2_o21ai_1 _13960_ (.B1(_04864_),
    .Y(_04865_),
    .A1(_04861_),
    .A2(_04862_));
 sg13g2_nand3_1 _13961_ (.B(_04823_),
    .C(_04865_),
    .A(_04831_),
    .Y(_04866_));
 sg13g2_inv_1 _13962_ (.Y(_04867_),
    .A(_04866_));
 sg13g2_a21oi_1 _13963_ (.A1(net43),
    .A2(_04858_),
    .Y(_04868_),
    .B1(_04867_));
 sg13g2_nor2_1 _13964_ (.A(_04800_),
    .B(_04801_),
    .Y(_04869_));
 sg13g2_nand2_1 _13965_ (.Y(_04870_),
    .A(_04869_),
    .B(_04798_));
 sg13g2_nand3_1 _13966_ (.B(_04807_),
    .C(_04800_),
    .A(_04799_),
    .Y(_04871_));
 sg13g2_inv_1 _13967_ (.Y(_04872_),
    .A(_04806_));
 sg13g2_nor2_1 _13968_ (.A(_04872_),
    .B(net89),
    .Y(_04873_));
 sg13g2_inv_1 _13969_ (.Y(_04874_),
    .A(_04873_));
 sg13g2_a21o_1 _13970_ (.A2(_04871_),
    .A1(_04870_),
    .B1(_04874_),
    .X(_04875_));
 sg13g2_nand3_1 _13971_ (.B(_04812_),
    .C(_04804_),
    .A(_04875_),
    .Y(_04876_));
 sg13g2_buf_1 _13972_ (.A(_04876_),
    .X(_04877_));
 sg13g2_o21ai_1 _13973_ (.B1(_04877_),
    .Y(_04878_),
    .A1(_04816_),
    .A2(_04868_));
 sg13g2_buf_1 _13974_ (.A(\b.gen_square[27].sq.piece[2] ),
    .X(_04879_));
 sg13g2_inv_1 _13975_ (.Y(_04880_),
    .A(_04879_));
 sg13g2_buf_2 _13976_ (.A(\b.gen_square[27].sq.piece[1] ),
    .X(_04881_));
 sg13g2_buf_1 _13977_ (.A(\b.gen_square[27].sq.piece[0] ),
    .X(_04882_));
 sg13g2_nand2_1 _13978_ (.Y(_04883_),
    .A(_04881_),
    .B(_04882_));
 sg13g2_nor2_1 _13979_ (.A(_04880_),
    .B(_04883_),
    .Y(_04884_));
 sg13g2_inv_1 _13980_ (.Y(_04885_),
    .A(_04884_));
 sg13g2_xnor2_1 _13981_ (.Y(_04886_),
    .A(net166),
    .B(\b.gen_square[27].sq.color ));
 sg13g2_buf_8 _13982_ (.A(_04886_),
    .X(_04887_));
 sg13g2_inv_1 _13983_ (.Y(_04888_),
    .A(_04882_));
 sg13g2_nor3_2 _13984_ (.A(_04881_),
    .B(_04880_),
    .C(_04888_),
    .Y(_04889_));
 sg13g2_inv_1 _13985_ (.Y(_04890_),
    .A(_04889_));
 sg13g2_nor2_1 _13986_ (.A(_04887_),
    .B(_04890_),
    .Y(_04891_));
 sg13g2_inv_1 _13987_ (.Y(_04892_),
    .A(_03640_));
 sg13g2_nor2_1 _13988_ (.A(net149),
    .B(_04892_),
    .Y(_04893_));
 sg13g2_a21oi_2 _13989_ (.B1(_04893_),
    .Y(_04894_),
    .A2(_04891_),
    .A1(net118));
 sg13g2_inv_2 _13990_ (.Y(_04895_),
    .A(_04894_));
 sg13g2_nor2_1 _13991_ (.A(_04885_),
    .B(_04895_),
    .Y(_04896_));
 sg13g2_buf_2 _13992_ (.A(_04896_),
    .X(_04897_));
 sg13g2_buf_1 _13993_ (.A(_04897_),
    .X(_04898_));
 sg13g2_and3_1 _13994_ (.X(_04899_),
    .A(_04880_),
    .B(_04888_),
    .C(_04881_));
 sg13g2_nor2_1 _13995_ (.A(_04881_),
    .B(_04882_),
    .Y(_04900_));
 sg13g2_nand2_1 _13996_ (.Y(_04901_),
    .A(_04900_),
    .B(_04879_));
 sg13g2_nand2b_1 _13997_ (.Y(_04902_),
    .B(_04901_),
    .A_N(_04899_));
 sg13g2_inv_1 _13998_ (.Y(_04903_),
    .A(_04887_));
 sg13g2_nor2_1 _13999_ (.A(_04903_),
    .B(net89),
    .Y(_04904_));
 sg13g2_nand2_1 _14000_ (.Y(_04905_),
    .A(_04902_),
    .B(_04904_));
 sg13g2_nand3_1 _14001_ (.B(_04885_),
    .C(_04905_),
    .A(_04894_),
    .Y(_04906_));
 sg13g2_inv_1 _14002_ (.Y(_04907_),
    .A(_04906_));
 sg13g2_a21oi_1 _14003_ (.A1(_04878_),
    .A2(net42),
    .Y(_04908_),
    .B1(_04907_));
 sg13g2_inv_1 _14004_ (.Y(_04909_),
    .A(_04908_));
 sg13g2_buf_1 _14005_ (.A(\b.gen_square[36].sq.piece[2] ),
    .X(_04910_));
 sg13g2_inv_1 _14006_ (.Y(_04911_),
    .A(_04910_));
 sg13g2_buf_1 _14007_ (.A(\b.gen_square[36].sq.piece[1] ),
    .X(_04912_));
 sg13g2_buf_2 _14008_ (.A(\b.gen_square[36].sq.piece[0] ),
    .X(_04913_));
 sg13g2_nand2_1 _14009_ (.Y(_04914_),
    .A(_04912_),
    .B(_04913_));
 sg13g2_nor2_1 _14010_ (.A(_04911_),
    .B(_04914_),
    .Y(_04915_));
 sg13g2_inv_1 _14011_ (.Y(_04916_),
    .A(_04915_));
 sg13g2_xnor2_1 _14012_ (.Y(_04917_),
    .A(net179),
    .B(\b.gen_square[36].sq.color ));
 sg13g2_buf_1 _14013_ (.A(_04917_),
    .X(_04918_));
 sg13g2_inv_1 _14014_ (.Y(_04919_),
    .A(_04913_));
 sg13g2_nor3_1 _14015_ (.A(_04912_),
    .B(_04911_),
    .C(_04919_),
    .Y(_04920_));
 sg13g2_inv_1 _14016_ (.Y(_04921_),
    .A(_04920_));
 sg13g2_nor2_1 _14017_ (.A(net146),
    .B(_04921_),
    .Y(_04922_));
 sg13g2_a22oi_1 _14018_ (.Y(_04923_),
    .B1(net134),
    .B2(_03730_),
    .A2(net152),
    .A1(_04922_));
 sg13g2_buf_2 _14019_ (.A(_04923_),
    .X(_04924_));
 sg13g2_inv_4 _14020_ (.A(_04924_),
    .Y(_04925_));
 sg13g2_nor2_1 _14021_ (.A(_04916_),
    .B(_04925_),
    .Y(_04926_));
 sg13g2_buf_2 _14022_ (.A(_04926_),
    .X(_04927_));
 sg13g2_buf_8 _14023_ (.A(_04927_),
    .X(_04928_));
 sg13g2_inv_1 _14024_ (.Y(_04929_),
    .A(net146));
 sg13g2_nor2_1 _14025_ (.A(_04929_),
    .B(net100),
    .Y(_04930_));
 sg13g2_nand3_1 _14026_ (.B(_04919_),
    .C(_04912_),
    .A(_04911_),
    .Y(_04931_));
 sg13g2_nor2_1 _14027_ (.A(_04912_),
    .B(_04913_),
    .Y(_04932_));
 sg13g2_nand2_1 _14028_ (.Y(_04933_),
    .A(_04932_),
    .B(_04910_));
 sg13g2_nand2_1 _14029_ (.Y(_04934_),
    .A(_04931_),
    .B(_04933_));
 sg13g2_nand2_1 _14030_ (.Y(_04935_),
    .A(_04930_),
    .B(_04934_));
 sg13g2_nand3_1 _14031_ (.B(_04916_),
    .C(_04935_),
    .A(_04924_),
    .Y(_04936_));
 sg13g2_buf_1 _14032_ (.A(_04936_),
    .X(_04937_));
 sg13g2_inv_1 _14033_ (.Y(_04938_),
    .A(_04937_));
 sg13g2_a21oi_1 _14034_ (.A1(_04909_),
    .A2(net58),
    .Y(_04939_),
    .B1(_04938_));
 sg13g2_inv_1 _14035_ (.Y(_04940_),
    .A(_04939_));
 sg13g2_nor3_1 _14036_ (.A(_04055_),
    .B(_04056_),
    .C(_04054_),
    .Y(_04941_));
 sg13g2_nor2_1 _14037_ (.A(_04053_),
    .B(_04056_),
    .Y(_04942_));
 sg13g2_nand2_1 _14038_ (.Y(_04943_),
    .A(_04942_),
    .B(_04055_));
 sg13g2_nand2b_1 _14039_ (.Y(_04944_),
    .B(_04943_),
    .A_N(_04941_));
 sg13g2_nand2_1 _14040_ (.Y(_04945_),
    .A(_04052_),
    .B(_04944_));
 sg13g2_inv_1 _14041_ (.Y(_04946_),
    .A(_04125_));
 sg13g2_nand3_1 _14042_ (.B(_04945_),
    .C(_04946_),
    .A(_04067_),
    .Y(_04947_));
 sg13g2_buf_1 _14043_ (.A(_04947_),
    .X(_04948_));
 sg13g2_inv_1 _14044_ (.Y(_04949_),
    .A(_04948_));
 sg13g2_a21oi_2 _14045_ (.B1(_04949_),
    .Y(_04950_),
    .A2(net71),
    .A1(_04940_));
 sg13g2_nand2_1 _14046_ (.Y(_04951_),
    .A(_04856_),
    .B(_04841_));
 sg13g2_nand2_1 _14047_ (.Y(_04952_),
    .A(_04951_),
    .B(_01759_));
 sg13g2_buf_2 _14048_ (.A(_04952_),
    .X(_04953_));
 sg13g2_inv_1 _14049_ (.Y(_04954_),
    .A(_00076_));
 sg13g2_nor2_1 _14050_ (.A(_04954_),
    .B(_04833_),
    .Y(_04955_));
 sg13g2_buf_2 _14051_ (.A(_04955_),
    .X(_04956_));
 sg13g2_a21oi_2 _14052_ (.B1(_04956_),
    .Y(_04957_),
    .A2(_04833_),
    .A1(_04953_));
 sg13g2_inv_2 _14053_ (.Y(_04958_),
    .A(_04957_));
 sg13g2_buf_1 _14054_ (.A(_04815_),
    .X(_04959_));
 sg13g2_inv_1 _14055_ (.Y(_04960_),
    .A(_00075_));
 sg13g2_nor2_1 _14056_ (.A(_04960_),
    .B(_04815_),
    .Y(_04961_));
 sg13g2_buf_2 _14057_ (.A(_04961_),
    .X(_04962_));
 sg13g2_a21oi_1 _14058_ (.A1(_04958_),
    .A2(net29),
    .Y(_04963_),
    .B1(_04962_));
 sg13g2_inv_1 _14059_ (.Y(_04964_),
    .A(_04963_));
 sg13g2_inv_1 _14060_ (.Y(_04965_),
    .A(_00074_));
 sg13g2_nor2_1 _14061_ (.A(_04965_),
    .B(_04897_),
    .Y(_04966_));
 sg13g2_buf_2 _14062_ (.A(_04966_),
    .X(_04967_));
 sg13g2_a21oi_1 _14063_ (.A1(_04964_),
    .A2(_04898_),
    .Y(_04968_),
    .B1(_04967_));
 sg13g2_inv_1 _14064_ (.Y(_04969_),
    .A(_04968_));
 sg13g2_inv_1 _14065_ (.Y(_04970_),
    .A(_00073_));
 sg13g2_nor2_1 _14066_ (.A(_04970_),
    .B(_04927_),
    .Y(_04971_));
 sg13g2_buf_2 _14067_ (.A(_04971_),
    .X(_04972_));
 sg13g2_a21oi_1 _14068_ (.A1(_04969_),
    .A2(net58),
    .Y(_04973_),
    .B1(_04972_));
 sg13g2_inv_1 _14069_ (.Y(_04974_),
    .A(_04973_));
 sg13g2_a21oi_1 _14070_ (.A1(_04974_),
    .A2(_04129_),
    .Y(_04975_),
    .B1(_04131_));
 sg13g2_inv_1 _14071_ (.Y(_04976_),
    .A(_04975_));
 sg13g2_a22oi_1 _14072_ (.Y(_04977_),
    .B1(_04950_),
    .B2(_04976_),
    .A2(_04797_),
    .A1(_04730_));
 sg13g2_inv_1 _14073_ (.Y(_04978_),
    .A(_04239_));
 sg13g2_a21oi_2 _14074_ (.B1(_04245_),
    .Y(_04979_),
    .A2(_04978_),
    .A1(_04326_));
 sg13g2_inv_1 _14075_ (.Y(_04980_),
    .A(_04571_));
 sg13g2_nand2_1 _14076_ (.Y(_04981_),
    .A(_04572_),
    .B(_04573_));
 sg13g2_nor2_1 _14077_ (.A(_04980_),
    .B(_04981_),
    .Y(_04982_));
 sg13g2_nand2_1 _14078_ (.Y(_04983_),
    .A(_04582_),
    .B(_04982_));
 sg13g2_nand2_1 _14079_ (.Y(_04984_),
    .A(_04983_),
    .B(_03760_));
 sg13g2_buf_2 _14080_ (.A(_04984_),
    .X(_04985_));
 sg13g2_a21oi_1 _14081_ (.A1(_04985_),
    .A2(net82),
    .Y(_04986_),
    .B1(_04251_));
 sg13g2_nor2_1 _14082_ (.A(_04979_),
    .B(_04986_),
    .Y(_04987_));
 sg13g2_buf_1 _14083_ (.A(_04987_),
    .X(_04988_));
 sg13g2_o21ai_1 _14084_ (.B1(_04725_),
    .Y(_04989_),
    .A1(_04715_),
    .A2(_04790_));
 sg13g2_inv_1 _14085_ (.Y(_04990_),
    .A(_04989_));
 sg13g2_nand2_1 _14086_ (.Y(_04991_),
    .A(_04554_),
    .B(_04555_));
 sg13g2_nor2_1 _14087_ (.A(_04560_),
    .B(_04991_),
    .Y(_04992_));
 sg13g2_inv_1 _14088_ (.Y(_04993_),
    .A(_04992_));
 sg13g2_nor2_1 _14089_ (.A(_04993_),
    .B(_04565_),
    .Y(_04994_));
 sg13g2_buf_2 _14090_ (.A(_04994_),
    .X(_04995_));
 sg13g2_nor2_2 _14091_ (.A(_03968_),
    .B(_04995_),
    .Y(_04996_));
 sg13g2_inv_4 _14092_ (.A(_04996_),
    .Y(_04997_));
 sg13g2_a21oi_2 _14093_ (.B1(_04728_),
    .Y(_04998_),
    .A2(net77),
    .A1(_04997_));
 sg13g2_nor2_2 _14094_ (.A(_04990_),
    .B(_04998_),
    .Y(_04999_));
 sg13g2_nor2_1 _14095_ (.A(_04988_),
    .B(_04999_),
    .Y(_05000_));
 sg13g2_nand2_1 _14096_ (.Y(_05001_),
    .A(_04977_),
    .B(_05000_));
 sg13g2_nor4_1 _14097_ (.A(_04134_),
    .B(_04359_),
    .C(_04588_),
    .D(_05001_),
    .Y(_05002_));
 sg13g2_inv_1 _14098_ (.Y(_05003_),
    .A(_04487_));
 sg13g2_nor2_1 _14099_ (.A(_05003_),
    .B(_04480_),
    .Y(_05004_));
 sg13g2_nor2_1 _14100_ (.A(_04435_),
    .B(_04440_),
    .Y(_05005_));
 sg13g2_nor2_1 _14101_ (.A(_04401_),
    .B(_04480_),
    .Y(_05006_));
 sg13g2_nor2_1 _14102_ (.A(_05005_),
    .B(_05006_),
    .Y(_05007_));
 sg13g2_nor2_1 _14103_ (.A(_04459_),
    .B(_04465_),
    .Y(_05008_));
 sg13g2_inv_2 _14104_ (.Y(_05009_),
    .A(_04382_));
 sg13g2_nor2_1 _14105_ (.A(_04376_),
    .B(_05009_),
    .Y(_05010_));
 sg13g2_nor2_1 _14106_ (.A(_05008_),
    .B(_05010_),
    .Y(_05011_));
 sg13g2_nand2_1 _14107_ (.Y(_05012_),
    .A(_05007_),
    .B(_05011_));
 sg13g2_nor2_1 _14108_ (.A(_04478_),
    .B(_05009_),
    .Y(_05013_));
 sg13g2_nor2_1 _14109_ (.A(_03812_),
    .B(_04526_),
    .Y(_05014_));
 sg13g2_buf_1 _14110_ (.A(_05014_),
    .X(_05015_));
 sg13g2_nor2_1 _14111_ (.A(_03968_),
    .B(_04566_),
    .Y(_05016_));
 sg13g2_nor2_1 _14112_ (.A(_03761_),
    .B(_04584_),
    .Y(_05017_));
 sg13g2_nor2_1 _14113_ (.A(_03740_),
    .B(_04547_),
    .Y(_05018_));
 sg13g2_buf_2 _14114_ (.A(_05018_),
    .X(_05019_));
 sg13g2_or2_1 _14115_ (.X(_05020_),
    .B(_05019_),
    .A(_05017_));
 sg13g2_nor3_1 _14116_ (.A(_05015_),
    .B(_05016_),
    .C(_05020_),
    .Y(_05021_));
 sg13g2_nand2b_1 _14117_ (.Y(_05022_),
    .B(_05021_),
    .A_N(_05013_));
 sg13g2_inv_1 _14118_ (.Y(_05023_),
    .A(_04950_));
 sg13g2_a21oi_2 _14119_ (.B1(_03993_),
    .Y(_05024_),
    .A2(_04423_),
    .A1(_04430_));
 sg13g2_nand2b_1 _14120_ (.Y(_05025_),
    .B(_05024_),
    .A_N(_04504_));
 sg13g2_o21ai_1 _14121_ (.B1(_05025_),
    .Y(_05026_),
    .A1(_05023_),
    .A2(_04976_));
 sg13g2_nor4_1 _14122_ (.A(_05004_),
    .B(_05012_),
    .C(_05022_),
    .D(_05026_),
    .Y(_05027_));
 sg13g2_nand2_1 _14123_ (.Y(_05028_),
    .A(_04495_),
    .B(_03984_));
 sg13g2_o21ai_1 _14124_ (.B1(_05028_),
    .Y(_05029_),
    .A1(_04356_),
    .A2(_04440_));
 sg13g2_a221oi_1 _14125_ (.B2(_04797_),
    .C1(_05029_),
    .B1(_04729_),
    .A1(_04334_),
    .Y(_05030_),
    .A2(_04252_));
 sg13g2_buf_2 _14126_ (.A(\b.gen_square[54].sq.piece[2] ),
    .X(_05031_));
 sg13g2_inv_1 _14127_ (.Y(_05032_),
    .A(_05031_));
 sg13g2_buf_1 _14128_ (.A(\b.gen_square[54].sq.piece[1] ),
    .X(_05033_));
 sg13g2_buf_2 _14129_ (.A(\b.gen_square[54].sq.piece[0] ),
    .X(_05034_));
 sg13g2_nand2_1 _14130_ (.Y(_05035_),
    .A(_05033_),
    .B(_05034_));
 sg13g2_nor2_1 _14131_ (.A(_05032_),
    .B(_05035_),
    .Y(_05036_));
 sg13g2_inv_1 _14132_ (.Y(_05037_),
    .A(_05036_));
 sg13g2_inv_1 _14133_ (.Y(_05038_),
    .A(_05033_));
 sg13g2_nand3_1 _14134_ (.B(_05031_),
    .C(_05034_),
    .A(_05038_),
    .Y(_05039_));
 sg13g2_buf_2 _14135_ (.A(_05039_),
    .X(_05040_));
 sg13g2_nor2_1 _14136_ (.A(_05040_),
    .B(net180),
    .Y(_05041_));
 sg13g2_nand2_1 _14137_ (.Y(_05042_),
    .A(_05041_),
    .B(net168));
 sg13g2_nand3_1 _14138_ (.B(_04063_),
    .C(_03901_),
    .A(_03592_),
    .Y(_05043_));
 sg13g2_nand2_1 _14139_ (.Y(_05044_),
    .A(_05042_),
    .B(_05043_));
 sg13g2_nor2_1 _14140_ (.A(_05037_),
    .B(_05044_),
    .Y(_05045_));
 sg13g2_buf_8 _14141_ (.A(_05045_),
    .X(_05046_));
 sg13g2_nand2_1 _14142_ (.Y(_05047_),
    .A(_04426_),
    .B(net98));
 sg13g2_inv_2 _14143_ (.Y(_05048_),
    .A(_05046_));
 sg13g2_nand2_1 _14144_ (.Y(_05049_),
    .A(_05048_),
    .B(_00034_));
 sg13g2_nand2_1 _14145_ (.Y(_05050_),
    .A(_05047_),
    .B(_05049_));
 sg13g2_nand2_1 _14146_ (.Y(_05051_),
    .A(_05050_),
    .B(_04128_));
 sg13g2_nand2_1 _14147_ (.Y(_05052_),
    .A(_05051_),
    .B(_04130_));
 sg13g2_nor2_1 _14148_ (.A(_04069_),
    .B(_05052_),
    .Y(_05053_));
 sg13g2_buf_2 _14149_ (.A(_05053_),
    .X(_05054_));
 sg13g2_inv_1 _14150_ (.Y(_05055_),
    .A(_05054_));
 sg13g2_nand2_1 _14151_ (.Y(_05056_),
    .A(_05024_),
    .B(_04431_));
 sg13g2_inv_1 _14152_ (.Y(_05057_),
    .A(_00039_));
 sg13g2_nand2_1 _14153_ (.Y(_05058_),
    .A(_04438_),
    .B(_05057_));
 sg13g2_nand2_1 _14154_ (.Y(_05059_),
    .A(_05058_),
    .B(_04247_));
 sg13g2_nand2_1 _14155_ (.Y(_05060_),
    .A(_05059_),
    .B(_04250_));
 sg13g2_nor2_1 _14156_ (.A(_04979_),
    .B(_05060_),
    .Y(_05061_));
 sg13g2_buf_1 _14157_ (.A(_05061_),
    .X(_05062_));
 sg13g2_inv_1 _14158_ (.Y(_05063_),
    .A(_00021_));
 sg13g2_nand2_2 _14159_ (.Y(_05064_),
    .A(_04464_),
    .B(_05063_));
 sg13g2_nand2_1 _14160_ (.Y(_05065_),
    .A(_05064_),
    .B(_04723_));
 sg13g2_nand2_1 _14161_ (.Y(_05066_),
    .A(_04727_),
    .B(_05065_));
 sg13g2_nor2_2 _14162_ (.A(_04990_),
    .B(_05066_),
    .Y(_05067_));
 sg13g2_nor2_1 _14163_ (.A(_05062_),
    .B(_05067_),
    .Y(_05068_));
 sg13g2_and3_1 _14164_ (.X(_05069_),
    .A(_05055_),
    .B(_05056_),
    .C(_05068_));
 sg13g2_and3_1 _14165_ (.X(_05070_),
    .A(_05027_),
    .B(_05030_),
    .C(_05069_));
 sg13g2_nor3_1 _14166_ (.A(net180),
    .B(_05002_),
    .C(_05070_),
    .Y(_05071_));
 sg13g2_buf_1 _14167_ (.A(_01968_),
    .X(_05072_));
 sg13g2_buf_1 _14168_ (.A(net215),
    .X(_05073_));
 sg13g2_buf_1 _14169_ (.A(net191),
    .X(_05074_));
 sg13g2_buf_1 _14170_ (.A(net177),
    .X(_05075_));
 sg13g2_buf_1 _14171_ (.A(_05075_),
    .X(_05076_));
 sg13g2_buf_1 _14172_ (.A(_05076_),
    .X(_05077_));
 sg13g2_buf_1 _14173_ (.A(net130),
    .X(_05078_));
 sg13g2_buf_1 _14174_ (.A(net114),
    .X(_05079_));
 sg13g2_nand2_1 _14175_ (.Y(_05080_),
    .A(_05071_),
    .B(net97));
 sg13g2_nand2_1 _14176_ (.Y(_05081_),
    .A(_05070_),
    .B(_05002_));
 sg13g2_buf_1 _14177_ (.A(_04044_),
    .X(_05082_));
 sg13g2_buf_1 _14178_ (.A(net176),
    .X(_05083_));
 sg13g2_buf_1 _14179_ (.A(net161),
    .X(_05084_));
 sg13g2_buf_1 _14180_ (.A(_05084_),
    .X(_05085_));
 sg13g2_buf_1 _14181_ (.A(net129),
    .X(_05086_));
 sg13g2_buf_1 _14182_ (.A(net113),
    .X(_05087_));
 sg13g2_buf_1 _14183_ (.A(net96),
    .X(_05088_));
 sg13g2_buf_1 _14184_ (.A(net86),
    .X(_05089_));
 sg13g2_buf_1 _14185_ (.A(net76),
    .X(_05090_));
 sg13g2_buf_1 _14186_ (.A(net68),
    .X(_05091_));
 sg13g2_buf_1 _14187_ (.A(net57),
    .X(_05092_));
 sg13g2_inv_1 _14188_ (.Y(_05093_),
    .A(net180));
 sg13g2_nand3_1 _14189_ (.B(net41),
    .C(_05093_),
    .A(_05081_),
    .Y(_05094_));
 sg13g2_nand2_1 _14190_ (.Y(_05095_),
    .A(_05080_),
    .B(_05094_));
 sg13g2_nand2_1 _14191_ (.Y(_05096_),
    .A(_05080_),
    .B(_05036_));
 sg13g2_nor2_1 _14192_ (.A(_05033_),
    .B(_05034_),
    .Y(_05097_));
 sg13g2_nand2b_1 _14193_ (.Y(_05098_),
    .B(_05035_),
    .A_N(_05097_));
 sg13g2_nand3_1 _14194_ (.B(_05096_),
    .C(_05098_),
    .A(_05095_),
    .Y(_05099_));
 sg13g2_a221oi_1 _14195_ (.B2(_04797_),
    .C1(_04359_),
    .B1(_04730_),
    .A1(_03985_),
    .Y(_05100_),
    .A2(_04495_));
 sg13g2_a21oi_1 _14196_ (.A1(_05100_),
    .A2(_05030_),
    .Y(_05101_),
    .B1(_05093_));
 sg13g2_inv_1 _14197_ (.Y(_05102_),
    .A(_05101_));
 sg13g2_nand4_1 _14198_ (.B(_05003_),
    .C(_04478_),
    .A(_05025_),
    .Y(_05103_),
    .D(_04505_));
 sg13g2_o21ai_1 _14199_ (.B1(net180),
    .Y(_05104_),
    .A1(_05103_),
    .A2(_04950_));
 sg13g2_nand2_1 _14200_ (.Y(_05105_),
    .A(_05097_),
    .B(_05031_));
 sg13g2_a21o_1 _14201_ (.A2(_05104_),
    .A1(_05102_),
    .B1(_05105_),
    .X(_05106_));
 sg13g2_nand4_1 _14202_ (.B(_05032_),
    .C(_05033_),
    .A(_05101_),
    .Y(_05107_),
    .D(_05034_));
 sg13g2_buf_1 _14203_ (.A(net183),
    .X(_05108_));
 sg13g2_buf_1 _14204_ (.A(net160),
    .X(_05109_));
 sg13g2_buf_1 _14205_ (.A(net143),
    .X(_05110_));
 sg13g2_buf_1 _14206_ (.A(net128),
    .X(_05111_));
 sg13g2_buf_1 _14207_ (.A(net112),
    .X(_05112_));
 sg13g2_buf_1 _14208_ (.A(_05112_),
    .X(_05113_));
 sg13g2_buf_1 _14209_ (.A(net85),
    .X(_05114_));
 sg13g2_buf_1 _14210_ (.A(net75),
    .X(_05115_));
 sg13g2_buf_1 _14211_ (.A(net67),
    .X(_05116_));
 sg13g2_nand2_1 _14212_ (.Y(_05117_),
    .A(_05040_),
    .B(net56));
 sg13g2_a21o_1 _14213_ (.A2(_05107_),
    .A1(_05106_),
    .B1(_05117_),
    .X(_05118_));
 sg13g2_nand2_1 _14214_ (.Y(_05119_),
    .A(_05099_),
    .B(_05118_));
 sg13g2_buf_1 _14215_ (.A(\b.gen_square[54].sq.mask ),
    .X(_05120_));
 sg13g2_nand2_1 _14216_ (.Y(_05121_),
    .A(_05119_),
    .B(_05120_));
 sg13g2_inv_1 _14217_ (.Y(_05122_),
    .A(_05121_));
 sg13g2_nor2_1 _14218_ (.A(net93),
    .B(_04619_),
    .Y(_05123_));
 sg13g2_inv_1 _14219_ (.Y(_05124_),
    .A(_04621_));
 sg13g2_nor3_1 _14220_ (.A(_04609_),
    .B(_04611_),
    .C(_04617_),
    .Y(_05125_));
 sg13g2_nand2_1 _14221_ (.Y(_05126_),
    .A(_05124_),
    .B(_05125_));
 sg13g2_inv_1 _14222_ (.Y(_05127_),
    .A(_00042_));
 sg13g2_xnor2_1 _14223_ (.Y(_05128_),
    .A(net150),
    .B(\b.gen_square[34].sq.color ));
 sg13g2_buf_2 _14224_ (.A(_05128_),
    .X(_05129_));
 sg13g2_buf_2 _14225_ (.A(\b.gen_square[34].sq.piece[2] ),
    .X(_05130_));
 sg13g2_buf_1 _14226_ (.A(\b.gen_square[34].sq.piece[1] ),
    .X(_05131_));
 sg13g2_buf_1 _14227_ (.A(\b.gen_square[34].sq.piece[0] ),
    .X(_05132_));
 sg13g2_inv_1 _14228_ (.Y(_05133_),
    .A(_05132_));
 sg13g2_nor3_1 _14229_ (.A(_05130_),
    .B(_05131_),
    .C(_05133_),
    .Y(_05134_));
 sg13g2_nand2_1 _14230_ (.Y(_05135_),
    .A(_05129_),
    .B(_05134_));
 sg13g2_inv_1 _14231_ (.Y(_05136_),
    .A(_05135_));
 sg13g2_inv_1 _14232_ (.Y(_05137_),
    .A(_05130_));
 sg13g2_nor3_2 _14233_ (.A(_05131_),
    .B(_05137_),
    .C(_05133_),
    .Y(_05138_));
 sg13g2_inv_1 _14234_ (.Y(_05139_),
    .A(_05138_));
 sg13g2_nor2_1 _14235_ (.A(_05129_),
    .B(_05139_),
    .Y(_05140_));
 sg13g2_a22oi_1 _14236_ (.Y(_05141_),
    .B1(net102),
    .B2(_05140_),
    .A2(net101),
    .A1(_03714_));
 sg13g2_buf_1 _14237_ (.A(_05141_),
    .X(_05142_));
 sg13g2_inv_2 _14238_ (.Y(_05143_),
    .A(_05142_));
 sg13g2_a21oi_1 _14239_ (.A1(net99),
    .A2(_05136_),
    .Y(_05144_),
    .B1(_05143_));
 sg13g2_nor2_1 _14240_ (.A(_05127_),
    .B(_05144_),
    .Y(_05145_));
 sg13g2_buf_2 _14241_ (.A(_05145_),
    .X(_05146_));
 sg13g2_inv_1 _14242_ (.Y(_05147_),
    .A(_00058_));
 sg13g2_xnor2_1 _14243_ (.Y(_05148_),
    .A(net163),
    .B(\b.gen_square[32].sq.color ));
 sg13g2_buf_8 _14244_ (.A(_05148_),
    .X(_05149_));
 sg13g2_buf_1 _14245_ (.A(\b.gen_square[32].sq.piece[2] ),
    .X(_05150_));
 sg13g2_buf_1 _14246_ (.A(\b.gen_square[32].sq.piece[1] ),
    .X(_05151_));
 sg13g2_buf_1 _14247_ (.A(\b.gen_square[32].sq.piece[0] ),
    .X(_05152_));
 sg13g2_inv_1 _14248_ (.Y(_05153_),
    .A(_05152_));
 sg13g2_nor3_1 _14249_ (.A(_05150_),
    .B(_05151_),
    .C(_05153_),
    .Y(_05154_));
 sg13g2_nand2_1 _14250_ (.Y(_05155_),
    .A(_05149_),
    .B(_05154_));
 sg13g2_inv_1 _14251_ (.Y(_05156_),
    .A(_05155_));
 sg13g2_inv_1 _14252_ (.Y(_05157_),
    .A(_05150_));
 sg13g2_nor3_2 _14253_ (.A(_05151_),
    .B(_05157_),
    .C(_05153_),
    .Y(_05158_));
 sg13g2_nor2b_1 _14254_ (.A(_05149_),
    .B_N(_05158_),
    .Y(_05159_));
 sg13g2_a22oi_1 _14255_ (.Y(_05160_),
    .B1(net135),
    .B2(_05159_),
    .A2(net134),
    .A1(_03698_));
 sg13g2_inv_4 _14256_ (.A(_05160_),
    .Y(_05161_));
 sg13g2_a21oi_1 _14257_ (.A1(net99),
    .A2(_05156_),
    .Y(_05162_),
    .B1(_05161_));
 sg13g2_nor2_1 _14258_ (.A(_05147_),
    .B(_05162_),
    .Y(_05163_));
 sg13g2_nor2_1 _14259_ (.A(_05146_),
    .B(_05163_),
    .Y(_05164_));
 sg13g2_inv_1 _14260_ (.Y(_05165_),
    .A(_00041_));
 sg13g2_xnor2_1 _14261_ (.Y(_05166_),
    .A(net136),
    .B(\b.gen_square[43].sq.color ));
 sg13g2_buf_1 _14262_ (.A(_05166_),
    .X(_05167_));
 sg13g2_buf_2 _14263_ (.A(\b.gen_square[43].sq.piece[2] ),
    .X(_05168_));
 sg13g2_buf_1 _14264_ (.A(\b.gen_square[43].sq.piece[1] ),
    .X(_05169_));
 sg13g2_buf_2 _14265_ (.A(\b.gen_square[43].sq.piece[0] ),
    .X(_05170_));
 sg13g2_inv_1 _14266_ (.Y(_05171_),
    .A(_05170_));
 sg13g2_nor3_1 _14267_ (.A(_05168_),
    .B(_05169_),
    .C(_05171_),
    .Y(_05172_));
 sg13g2_nand2_1 _14268_ (.Y(_05173_),
    .A(net94),
    .B(_05172_));
 sg13g2_inv_1 _14269_ (.Y(_05174_),
    .A(_05173_));
 sg13g2_inv_1 _14270_ (.Y(_05175_),
    .A(_05168_));
 sg13g2_nor3_2 _14271_ (.A(_05169_),
    .B(_05175_),
    .C(_05171_),
    .Y(_05176_));
 sg13g2_inv_1 _14272_ (.Y(_05177_),
    .A(_05176_));
 sg13g2_nor2_1 _14273_ (.A(net94),
    .B(_05177_),
    .Y(_05178_));
 sg13g2_a22oi_1 _14274_ (.Y(_05179_),
    .B1(net92),
    .B2(_05178_),
    .A2(net91),
    .A1(_03805_));
 sg13g2_buf_2 _14275_ (.A(_05179_),
    .X(_05180_));
 sg13g2_inv_4 _14276_ (.A(_05180_),
    .Y(_05181_));
 sg13g2_a21oi_1 _14277_ (.A1(net88),
    .A2(_05174_),
    .Y(_05182_),
    .B1(_05181_));
 sg13g2_nor2_2 _14278_ (.A(_05165_),
    .B(_05182_),
    .Y(_05183_));
 sg13g2_inv_1 _14279_ (.Y(_05184_),
    .A(_05183_));
 sg13g2_inv_1 _14280_ (.Y(_05185_),
    .A(_00024_));
 sg13g2_xnor2_1 _14281_ (.Y(_05186_),
    .A(net150),
    .B(\b.gen_square[59].sq.color ));
 sg13g2_buf_2 _14282_ (.A(_05186_),
    .X(_05187_));
 sg13g2_buf_1 _14283_ (.A(\b.gen_square[59].sq.piece[2] ),
    .X(_05188_));
 sg13g2_buf_1 _14284_ (.A(\b.gen_square[59].sq.piece[1] ),
    .X(_05189_));
 sg13g2_buf_1 _14285_ (.A(\b.gen_square[59].sq.piece[0] ),
    .X(_05190_));
 sg13g2_inv_1 _14286_ (.Y(_05191_),
    .A(_05190_));
 sg13g2_nor3_1 _14287_ (.A(_05188_),
    .B(_05189_),
    .C(_05191_),
    .Y(_05192_));
 sg13g2_nand2_1 _14288_ (.Y(_05193_),
    .A(_05187_),
    .B(_05192_));
 sg13g2_inv_1 _14289_ (.Y(_05194_),
    .A(_05193_));
 sg13g2_inv_1 _14290_ (.Y(_05195_),
    .A(_05188_));
 sg13g2_nor3_2 _14291_ (.A(_05189_),
    .B(_05195_),
    .C(_05191_),
    .Y(_05196_));
 sg13g2_nor2b_1 _14292_ (.A(_05187_),
    .B_N(_05196_),
    .Y(_05197_));
 sg13g2_a22oi_1 _14293_ (.Y(_05198_),
    .B1(net102),
    .B2(_05197_),
    .A2(net101),
    .A1(_03951_));
 sg13g2_inv_2 _14294_ (.Y(_05199_),
    .A(_05198_));
 sg13g2_a21oi_1 _14295_ (.A1(net69),
    .A2(_05194_),
    .Y(_05200_),
    .B1(_05199_));
 sg13g2_nor2_1 _14296_ (.A(_05185_),
    .B(_05200_),
    .Y(_05201_));
 sg13g2_inv_1 _14297_ (.Y(_05202_),
    .A(_05201_));
 sg13g2_nand3_1 _14298_ (.B(_05184_),
    .C(_05202_),
    .A(_05164_),
    .Y(_05203_));
 sg13g2_nor2_1 _14299_ (.A(_03693_),
    .B(_05162_),
    .Y(_05204_));
 sg13g2_nor2_1 _14300_ (.A(_03713_),
    .B(_05144_),
    .Y(_05205_));
 sg13g2_inv_1 _14301_ (.Y(_05206_),
    .A(_05205_));
 sg13g2_nand2b_1 _14302_ (.Y(_05207_),
    .B(_05206_),
    .A_N(_05204_));
 sg13g2_nor2_2 _14303_ (.A(_03804_),
    .B(_05182_),
    .Y(_05208_));
 sg13g2_nor2_1 _14304_ (.A(_03950_),
    .B(_05200_),
    .Y(_05209_));
 sg13g2_nor2_1 _14305_ (.A(_05208_),
    .B(_05209_),
    .Y(_05210_));
 sg13g2_nor2b_1 _14306_ (.A(_05207_),
    .B_N(_05210_),
    .Y(_05211_));
 sg13g2_nor2b_1 _14307_ (.A(_05203_),
    .B_N(_05211_),
    .Y(_05212_));
 sg13g2_xnor2_1 _14308_ (.Y(_05213_),
    .A(net150),
    .B(\b.gen_square[58].sq.color ));
 sg13g2_buf_8 _14309_ (.A(_05213_),
    .X(_05214_));
 sg13g2_buf_1 _14310_ (.A(\b.gen_square[58].sq.piece[1] ),
    .X(_05215_));
 sg13g2_buf_2 _14311_ (.A(\b.gen_square[58].sq.piece[0] ),
    .X(_05216_));
 sg13g2_nor2_1 _14312_ (.A(_05215_),
    .B(_05216_),
    .Y(_05217_));
 sg13g2_buf_1 _14313_ (.A(\b.gen_square[58].sq.piece[2] ),
    .X(_05218_));
 sg13g2_nand2_1 _14314_ (.Y(_05219_),
    .A(_05217_),
    .B(_05218_));
 sg13g2_inv_1 _14315_ (.Y(_05220_),
    .A(_05218_));
 sg13g2_inv_1 _14316_ (.Y(_05221_),
    .A(_05216_));
 sg13g2_nand3_1 _14317_ (.B(_05221_),
    .C(_05215_),
    .A(_05220_),
    .Y(_05222_));
 sg13g2_a21oi_1 _14318_ (.A1(_05219_),
    .A2(_05222_),
    .Y(_05223_),
    .B1(net32));
 sg13g2_inv_1 _14319_ (.Y(_05224_),
    .A(_05215_));
 sg13g2_nand3_1 _14320_ (.B(_05218_),
    .C(_05216_),
    .A(_05224_),
    .Y(_05225_));
 sg13g2_buf_1 _14321_ (.A(_05225_),
    .X(_05226_));
 sg13g2_nor2_1 _14322_ (.A(_05226_),
    .B(_05214_),
    .Y(_05227_));
 sg13g2_a22oi_1 _14323_ (.Y(_05228_),
    .B1(net101),
    .B2(_03943_),
    .A2(net118),
    .A1(_05227_));
 sg13g2_buf_1 _14324_ (.A(_05228_),
    .X(_05229_));
 sg13g2_inv_1 _14325_ (.Y(_05230_),
    .A(_05229_));
 sg13g2_a21oi_2 _14326_ (.B1(_05230_),
    .Y(_05231_),
    .A2(_05223_),
    .A1(_05214_));
 sg13g2_xnor2_1 _14327_ (.Y(_05232_),
    .A(net179),
    .B(\b.gen_square[40].sq.color ));
 sg13g2_buf_8 _14328_ (.A(_05232_),
    .X(_05233_));
 sg13g2_buf_1 _14329_ (.A(\b.gen_square[40].sq.piece[2] ),
    .X(_05234_));
 sg13g2_inv_1 _14330_ (.Y(_05235_),
    .A(_05234_));
 sg13g2_buf_1 _14331_ (.A(\b.gen_square[40].sq.piece[1] ),
    .X(_05236_));
 sg13g2_buf_2 _14332_ (.A(\b.gen_square[40].sq.piece[0] ),
    .X(_05237_));
 sg13g2_nor2_1 _14333_ (.A(_05236_),
    .B(_05237_),
    .Y(_05238_));
 sg13g2_inv_1 _14334_ (.Y(_05239_),
    .A(_05238_));
 sg13g2_nor2_1 _14335_ (.A(_05235_),
    .B(_05239_),
    .Y(_05240_));
 sg13g2_inv_1 _14336_ (.Y(_05241_),
    .A(_05240_));
 sg13g2_inv_1 _14337_ (.Y(_05242_),
    .A(_05237_));
 sg13g2_nand3_1 _14338_ (.B(_05242_),
    .C(_05236_),
    .A(_05235_),
    .Y(_05243_));
 sg13g2_a21oi_1 _14339_ (.A1(_05241_),
    .A2(_05243_),
    .Y(_05244_),
    .B1(net46));
 sg13g2_inv_1 _14340_ (.Y(_05245_),
    .A(_05236_));
 sg13g2_nand3_1 _14341_ (.B(_05234_),
    .C(_05237_),
    .A(_05245_),
    .Y(_05246_));
 sg13g2_buf_1 _14342_ (.A(_05246_),
    .X(_05247_));
 sg13g2_nor2_1 _14343_ (.A(_05247_),
    .B(_05233_),
    .Y(_05248_));
 sg13g2_a22oi_1 _14344_ (.Y(_05249_),
    .B1(_03779_),
    .B2(net134),
    .A2(net152),
    .A1(_05248_));
 sg13g2_inv_2 _14345_ (.Y(_05250_),
    .A(_05249_));
 sg13g2_a21oi_1 _14346_ (.A1(_05233_),
    .A2(_05244_),
    .Y(_05251_),
    .B1(_05250_));
 sg13g2_buf_2 _14347_ (.A(_05251_),
    .X(_05252_));
 sg13g2_buf_1 _14348_ (.A(\b.gen_square[56].sq.piece[1] ),
    .X(_05253_));
 sg13g2_buf_2 _14349_ (.A(\b.gen_square[56].sq.piece[0] ),
    .X(_05254_));
 sg13g2_nor2_1 _14350_ (.A(_05253_),
    .B(_05254_),
    .Y(_05255_));
 sg13g2_buf_1 _14351_ (.A(\b.gen_square[56].sq.piece[2] ),
    .X(_05256_));
 sg13g2_nand2_1 _14352_ (.Y(_05257_),
    .A(_05255_),
    .B(_05256_));
 sg13g2_inv_1 _14353_ (.Y(_05258_),
    .A(_05253_));
 sg13g2_nor3_1 _14354_ (.A(_05256_),
    .B(_05254_),
    .C(_05258_),
    .Y(_05259_));
 sg13g2_inv_1 _14355_ (.Y(_05260_),
    .A(_05259_));
 sg13g2_a21oi_1 _14356_ (.A1(_05257_),
    .A2(_05260_),
    .Y(_05261_),
    .B1(net46));
 sg13g2_xnor2_1 _14357_ (.Y(_05262_),
    .A(net216),
    .B(\b.gen_square[56].sq.color ));
 sg13g2_buf_2 _14358_ (.A(_05262_),
    .X(_05263_));
 sg13g2_nand2_1 _14359_ (.Y(_05264_),
    .A(_03927_),
    .B(net167));
 sg13g2_nand3_1 _14360_ (.B(_05256_),
    .C(_05254_),
    .A(_05258_),
    .Y(_05265_));
 sg13g2_buf_2 _14361_ (.A(_05265_),
    .X(_05266_));
 sg13g2_nor2_1 _14362_ (.A(_05266_),
    .B(_05263_),
    .Y(_05267_));
 sg13g2_nand2_1 _14363_ (.Y(_05268_),
    .A(_05267_),
    .B(net148));
 sg13g2_nand2_2 _14364_ (.Y(_05269_),
    .A(_05264_),
    .B(_05268_));
 sg13g2_a21oi_2 _14365_ (.B1(_05269_),
    .Y(_05270_),
    .A2(_05263_),
    .A1(_05261_));
 sg13g2_nand3_1 _14366_ (.B(_05252_),
    .C(_05270_),
    .A(_05231_),
    .Y(_05271_));
 sg13g2_buf_2 _14367_ (.A(\b.gen_square[21].sq.piece[2] ),
    .X(_05272_));
 sg13g2_inv_2 _14368_ (.Y(_05273_),
    .A(_05272_));
 sg13g2_buf_1 _14369_ (.A(\b.gen_square[21].sq.piece[1] ),
    .X(_05274_));
 sg13g2_buf_1 _14370_ (.A(\b.gen_square[21].sq.piece[0] ),
    .X(_05275_));
 sg13g2_nand2_1 _14371_ (.Y(_05276_),
    .A(_05274_),
    .B(_05275_));
 sg13g2_nor2_1 _14372_ (.A(_05273_),
    .B(_05276_),
    .Y(_05277_));
 sg13g2_inv_1 _14373_ (.Y(_05278_),
    .A(_05277_));
 sg13g2_xnor2_1 _14374_ (.Y(_05279_),
    .A(_04078_),
    .B(\b.gen_square[21].sq.color ));
 sg13g2_buf_2 _14375_ (.A(_05279_),
    .X(_05280_));
 sg13g2_inv_1 _14376_ (.Y(_05281_),
    .A(_05275_));
 sg13g2_nor3_2 _14377_ (.A(_05274_),
    .B(_05273_),
    .C(_05281_),
    .Y(_05282_));
 sg13g2_inv_1 _14378_ (.Y(_05283_),
    .A(_05282_));
 sg13g2_nor2_1 _14379_ (.A(_05280_),
    .B(_05283_),
    .Y(_05284_));
 sg13g2_a22oi_1 _14380_ (.Y(_05285_),
    .B1(_04085_),
    .B2(_05284_),
    .A2(net101),
    .A1(_03583_));
 sg13g2_buf_2 _14381_ (.A(_05285_),
    .X(_05286_));
 sg13g2_inv_4 _14382_ (.A(_05286_),
    .Y(_05287_));
 sg13g2_nor2_1 _14383_ (.A(_05278_),
    .B(_05287_),
    .Y(_05288_));
 sg13g2_buf_2 _14384_ (.A(_05288_),
    .X(_05289_));
 sg13g2_inv_2 _14385_ (.Y(_05290_),
    .A(_05289_));
 sg13g2_buf_1 _14386_ (.A(\b.gen_square[7].sq.piece[2] ),
    .X(_05291_));
 sg13g2_buf_1 _14387_ (.A(\b.gen_square[7].sq.piece[0] ),
    .X(_05292_));
 sg13g2_buf_1 _14388_ (.A(\b.gen_square[7].sq.piece[1] ),
    .X(_05293_));
 sg13g2_inv_1 _14389_ (.Y(_05294_),
    .A(_05293_));
 sg13g2_nor3_1 _14390_ (.A(_05291_),
    .B(_05292_),
    .C(_05294_),
    .Y(_05295_));
 sg13g2_inv_2 _14391_ (.Y(_05296_),
    .A(_05291_));
 sg13g2_nor2_1 _14392_ (.A(_05293_),
    .B(_05292_),
    .Y(_05297_));
 sg13g2_inv_1 _14393_ (.Y(_05298_),
    .A(_05297_));
 sg13g2_nor2_2 _14394_ (.A(_05296_),
    .B(_05298_),
    .Y(_05299_));
 sg13g2_nor2_1 _14395_ (.A(_05295_),
    .B(_05299_),
    .Y(_05300_));
 sg13g2_xnor2_1 _14396_ (.Y(_05301_),
    .A(net179),
    .B(_04009_));
 sg13g2_buf_2 _14397_ (.A(_05301_),
    .X(_05302_));
 sg13g2_nand2_1 _14398_ (.Y(_05303_),
    .A(net147),
    .B(_05302_));
 sg13g2_nand3_1 _14399_ (.B(_05291_),
    .C(_05292_),
    .A(_05294_),
    .Y(_05304_));
 sg13g2_buf_1 _14400_ (.A(_05304_),
    .X(_05305_));
 sg13g2_nor2_1 _14401_ (.A(_05305_),
    .B(_05302_),
    .Y(_05306_));
 sg13g2_nand2_1 _14402_ (.Y(_05307_),
    .A(_05306_),
    .B(_04061_));
 sg13g2_nand3_1 _14403_ (.B(net151),
    .C(_01814_),
    .A(_03604_),
    .Y(_05308_));
 sg13g2_nand2_1 _14404_ (.Y(_05309_),
    .A(_05307_),
    .B(_05308_));
 sg13g2_inv_1 _14405_ (.Y(_05310_),
    .A(_05309_));
 sg13g2_o21ai_1 _14406_ (.B1(_05310_),
    .Y(_05311_),
    .A1(_05300_),
    .A2(_05303_));
 sg13g2_inv_1 _14407_ (.Y(_05312_),
    .A(_05311_));
 sg13g2_nor3_1 _14408_ (.A(_04177_),
    .B(_04180_),
    .C(_04185_),
    .Y(_05313_));
 sg13g2_nand2b_1 _14409_ (.Y(_05314_),
    .B(_04276_),
    .A_N(_05313_));
 sg13g2_nand2_1 _14410_ (.Y(_05315_),
    .A(_04273_),
    .B(_05314_));
 sg13g2_nand3_1 _14411_ (.B(_04183_),
    .C(_05315_),
    .A(_04271_),
    .Y(_05316_));
 sg13g2_inv_1 _14412_ (.Y(_05317_),
    .A(_05316_));
 sg13g2_a21oi_1 _14413_ (.A1(_05312_),
    .A2(net81),
    .Y(_05318_),
    .B1(_05317_));
 sg13g2_inv_1 _14414_ (.Y(_05319_),
    .A(_05280_));
 sg13g2_nor2_1 _14415_ (.A(_05319_),
    .B(net70),
    .Y(_05320_));
 sg13g2_and3_1 _14416_ (.X(_05321_),
    .A(_05273_),
    .B(_05281_),
    .C(_05274_));
 sg13g2_inv_1 _14417_ (.Y(_05322_),
    .A(_05321_));
 sg13g2_nor2_1 _14418_ (.A(_05274_),
    .B(_05275_),
    .Y(_05323_));
 sg13g2_nand2_1 _14419_ (.Y(_05324_),
    .A(_05323_),
    .B(_05272_));
 sg13g2_nand2_1 _14420_ (.Y(_05325_),
    .A(_05322_),
    .B(_05324_));
 sg13g2_nand2_1 _14421_ (.Y(_05326_),
    .A(_05320_),
    .B(_05325_));
 sg13g2_nand3_1 _14422_ (.B(_05278_),
    .C(_05326_),
    .A(_05286_),
    .Y(_05327_));
 sg13g2_o21ai_1 _14423_ (.B1(_05327_),
    .Y(_05328_),
    .A1(_05290_),
    .A2(_05318_));
 sg13g2_buf_1 _14424_ (.A(\b.gen_square[28].sq.piece[2] ),
    .X(_05329_));
 sg13g2_inv_1 _14425_ (.Y(_05330_),
    .A(_05329_));
 sg13g2_buf_1 _14426_ (.A(\b.gen_square[28].sq.piece[1] ),
    .X(_05331_));
 sg13g2_buf_1 _14427_ (.A(\b.gen_square[28].sq.piece[0] ),
    .X(_05332_));
 sg13g2_nand2_1 _14428_ (.Y(_05333_),
    .A(_05331_),
    .B(_05332_));
 sg13g2_nor2_1 _14429_ (.A(_05330_),
    .B(_05333_),
    .Y(_05334_));
 sg13g2_inv_1 _14430_ (.Y(_05335_),
    .A(_05334_));
 sg13g2_xnor2_1 _14431_ (.Y(_05336_),
    .A(net163),
    .B(\b.gen_square[28].sq.color ));
 sg13g2_buf_2 _14432_ (.A(_05336_),
    .X(_05337_));
 sg13g2_inv_1 _14433_ (.Y(_05338_),
    .A(_05332_));
 sg13g2_nor3_1 _14434_ (.A(_05331_),
    .B(_05330_),
    .C(_05338_),
    .Y(_05339_));
 sg13g2_inv_1 _14435_ (.Y(_05340_),
    .A(_05339_));
 sg13g2_nor2_1 _14436_ (.A(_05337_),
    .B(_05340_),
    .Y(_05341_));
 sg13g2_a22oi_1 _14437_ (.Y(_05342_),
    .B1(net135),
    .B2(_05341_),
    .A2(net134),
    .A1(_03651_));
 sg13g2_buf_1 _14438_ (.A(_05342_),
    .X(_05343_));
 sg13g2_inv_4 _14439_ (.A(_05343_),
    .Y(_05344_));
 sg13g2_nor2_1 _14440_ (.A(_05335_),
    .B(_05344_),
    .Y(_05345_));
 sg13g2_buf_1 _14441_ (.A(_05345_),
    .X(_05346_));
 sg13g2_buf_1 _14442_ (.A(net55),
    .X(_05347_));
 sg13g2_and3_1 _14443_ (.X(_05348_),
    .A(_05330_),
    .B(_05338_),
    .C(_05331_));
 sg13g2_nor2_1 _14444_ (.A(_05331_),
    .B(_05332_),
    .Y(_05349_));
 sg13g2_nand2_1 _14445_ (.Y(_05350_),
    .A(_05349_),
    .B(_05329_));
 sg13g2_nand2b_1 _14446_ (.Y(_05351_),
    .B(_05350_),
    .A_N(_05348_));
 sg13g2_inv_1 _14447_ (.Y(_05352_),
    .A(_05337_));
 sg13g2_nor2_1 _14448_ (.A(_05352_),
    .B(net89),
    .Y(_05353_));
 sg13g2_nand2_1 _14449_ (.Y(_05354_),
    .A(_05351_),
    .B(_05353_));
 sg13g2_nand3_1 _14450_ (.B(_05335_),
    .C(_05354_),
    .A(_05343_),
    .Y(_05355_));
 sg13g2_buf_1 _14451_ (.A(_05355_),
    .X(_05356_));
 sg13g2_inv_1 _14452_ (.Y(_05357_),
    .A(_05356_));
 sg13g2_a21oi_1 _14453_ (.A1(_05328_),
    .A2(net40),
    .Y(_05358_),
    .B1(_05357_));
 sg13g2_inv_1 _14454_ (.Y(_05359_),
    .A(_05358_));
 sg13g2_buf_1 _14455_ (.A(\b.gen_square[35].sq.piece[2] ),
    .X(_05360_));
 sg13g2_inv_1 _14456_ (.Y(_05361_),
    .A(_05360_));
 sg13g2_buf_1 _14457_ (.A(\b.gen_square[35].sq.piece[1] ),
    .X(_05362_));
 sg13g2_buf_1 _14458_ (.A(\b.gen_square[35].sq.piece[0] ),
    .X(_05363_));
 sg13g2_nand2_1 _14459_ (.Y(_05364_),
    .A(_05362_),
    .B(_05363_));
 sg13g2_nor2_1 _14460_ (.A(_05361_),
    .B(_05364_),
    .Y(_05365_));
 sg13g2_inv_1 _14461_ (.Y(_05366_),
    .A(_05365_));
 sg13g2_xnor2_1 _14462_ (.Y(_05367_),
    .A(net179),
    .B(\b.gen_square[35].sq.color ));
 sg13g2_buf_8 _14463_ (.A(_05367_),
    .X(_05368_));
 sg13g2_inv_1 _14464_ (.Y(_05369_),
    .A(_05363_));
 sg13g2_nor3_2 _14465_ (.A(_05362_),
    .B(_05361_),
    .C(_05369_),
    .Y(_05370_));
 sg13g2_inv_1 _14466_ (.Y(_05371_),
    .A(_05370_));
 sg13g2_nor2_1 _14467_ (.A(_05368_),
    .B(_05371_),
    .Y(_05372_));
 sg13g2_a22oi_1 _14468_ (.Y(_05373_),
    .B1(net152),
    .B2(_05372_),
    .A2(net151),
    .A1(_03722_));
 sg13g2_buf_2 _14469_ (.A(_05373_),
    .X(_05374_));
 sg13g2_inv_4 _14470_ (.A(_05374_),
    .Y(_05375_));
 sg13g2_nor2_1 _14471_ (.A(_05366_),
    .B(_05375_),
    .Y(_05376_));
 sg13g2_buf_8 _14472_ (.A(_05376_),
    .X(_05377_));
 sg13g2_buf_1 _14473_ (.A(_05377_),
    .X(_05378_));
 sg13g2_inv_1 _14474_ (.Y(_05379_),
    .A(_05368_));
 sg13g2_nor2_1 _14475_ (.A(_05379_),
    .B(net100),
    .Y(_05380_));
 sg13g2_nand3_1 _14476_ (.B(_05369_),
    .C(_05362_),
    .A(_05361_),
    .Y(_05381_));
 sg13g2_nor2_1 _14477_ (.A(_05362_),
    .B(_05363_),
    .Y(_05382_));
 sg13g2_nand2_1 _14478_ (.Y(_05383_),
    .A(_05382_),
    .B(_05360_));
 sg13g2_nand2_1 _14479_ (.Y(_05384_),
    .A(_05381_),
    .B(_05383_));
 sg13g2_nand2_1 _14480_ (.Y(_05385_),
    .A(_05380_),
    .B(_05384_));
 sg13g2_nand3_1 _14481_ (.B(_05366_),
    .C(_05385_),
    .A(_05374_),
    .Y(_05386_));
 sg13g2_inv_1 _14482_ (.Y(_05387_),
    .A(_05386_));
 sg13g2_a21oi_1 _14483_ (.A1(_05359_),
    .A2(net54),
    .Y(_05388_),
    .B1(_05387_));
 sg13g2_inv_1 _14484_ (.Y(_05389_),
    .A(_05388_));
 sg13g2_buf_2 _14485_ (.A(\b.gen_square[42].sq.piece[2] ),
    .X(_05390_));
 sg13g2_inv_2 _14486_ (.Y(_05391_),
    .A(_05390_));
 sg13g2_buf_1 _14487_ (.A(\b.gen_square[42].sq.piece[1] ),
    .X(_05392_));
 sg13g2_buf_2 _14488_ (.A(\b.gen_square[42].sq.piece[0] ),
    .X(_05393_));
 sg13g2_nand2_1 _14489_ (.Y(_05394_),
    .A(_05392_),
    .B(_05393_));
 sg13g2_nor2_1 _14490_ (.A(_05391_),
    .B(_05394_),
    .Y(_05395_));
 sg13g2_inv_1 _14491_ (.Y(_05396_),
    .A(_05395_));
 sg13g2_xnor2_1 _14492_ (.Y(_05397_),
    .A(net166),
    .B(\b.gen_square[42].sq.color ));
 sg13g2_buf_2 _14493_ (.A(_05397_),
    .X(_05398_));
 sg13g2_inv_2 _14494_ (.Y(_05399_),
    .A(_05393_));
 sg13g2_nor3_2 _14495_ (.A(_05392_),
    .B(_05391_),
    .C(_05399_),
    .Y(_05400_));
 sg13g2_inv_2 _14496_ (.Y(_05401_),
    .A(_05400_));
 sg13g2_nor2_1 _14497_ (.A(_05398_),
    .B(_05401_),
    .Y(_05402_));
 sg13g2_a22oi_1 _14498_ (.Y(_05403_),
    .B1(net135),
    .B2(_05402_),
    .A2(net117),
    .A1(_03797_));
 sg13g2_buf_2 _14499_ (.A(_05403_),
    .X(_05404_));
 sg13g2_inv_4 _14500_ (.A(_05404_),
    .Y(_05405_));
 sg13g2_nor2_1 _14501_ (.A(_05396_),
    .B(_05405_),
    .Y(_05406_));
 sg13g2_buf_1 _14502_ (.A(_05406_),
    .X(_05407_));
 sg13g2_buf_1 _14503_ (.A(_05407_),
    .X(_05408_));
 sg13g2_inv_1 _14504_ (.Y(_05409_),
    .A(_05398_));
 sg13g2_nor2_1 _14505_ (.A(_05409_),
    .B(net79),
    .Y(_05410_));
 sg13g2_nand3_1 _14506_ (.B(_05399_),
    .C(_05392_),
    .A(_05391_),
    .Y(_05411_));
 sg13g2_nor2_1 _14507_ (.A(_05392_),
    .B(_05393_),
    .Y(_05412_));
 sg13g2_nand2_1 _14508_ (.Y(_05413_),
    .A(_05412_),
    .B(_05390_));
 sg13g2_nand2_1 _14509_ (.Y(_05414_),
    .A(_05411_),
    .B(_05413_));
 sg13g2_nand2_1 _14510_ (.Y(_05415_),
    .A(_05410_),
    .B(_05414_));
 sg13g2_nand3_1 _14511_ (.B(_05396_),
    .C(_05415_),
    .A(_05404_),
    .Y(_05416_));
 sg13g2_inv_1 _14512_ (.Y(_05417_),
    .A(_05416_));
 sg13g2_a21oi_1 _14513_ (.A1(_05389_),
    .A2(_05408_),
    .Y(_05418_),
    .B1(_05417_));
 sg13g2_o21ai_1 _14514_ (.B1(_05124_),
    .Y(_05419_),
    .A1(_05271_),
    .A2(_05418_));
 sg13g2_and3_1 _14515_ (.X(_05420_),
    .A(_04610_),
    .B(_04617_),
    .C(_04611_));
 sg13g2_nand2b_1 _14516_ (.Y(_05421_),
    .B(_05420_),
    .A_N(_05419_));
 sg13g2_o21ai_1 _14517_ (.B1(_05421_),
    .Y(_05422_),
    .A1(_05126_),
    .A2(_05212_));
 sg13g2_xnor2_1 _14518_ (.Y(_05423_),
    .A(_04609_),
    .B(_04749_));
 sg13g2_a21oi_1 _14519_ (.A1(_05410_),
    .A2(_05400_),
    .Y(_05424_),
    .B1(_05405_));
 sg13g2_inv_1 _14520_ (.Y(_05425_),
    .A(_05256_));
 sg13g2_nand2_1 _14521_ (.Y(_05426_),
    .A(_05253_),
    .B(_05254_));
 sg13g2_nor2_1 _14522_ (.A(_05425_),
    .B(_05426_),
    .Y(_05427_));
 sg13g2_nand3_1 _14523_ (.B(_05268_),
    .C(_05427_),
    .A(_05264_),
    .Y(_05428_));
 sg13g2_inv_1 _14524_ (.Y(_05429_),
    .A(_00027_));
 sg13g2_nand2_1 _14525_ (.Y(_05430_),
    .A(_05428_),
    .B(_05429_));
 sg13g2_buf_2 _14526_ (.A(_05430_),
    .X(_05431_));
 sg13g2_a21oi_1 _14527_ (.A1(_05431_),
    .A2(_04625_),
    .Y(_05432_),
    .B1(_04629_));
 sg13g2_inv_1 _14528_ (.Y(_05433_),
    .A(_05432_));
 sg13g2_inv_1 _14529_ (.Y(_05434_),
    .A(_00050_));
 sg13g2_nor2_1 _14530_ (.A(_05434_),
    .B(_05407_),
    .Y(_05435_));
 sg13g2_buf_8 _14531_ (.A(_05435_),
    .X(_05436_));
 sg13g2_a21oi_1 _14532_ (.A1(_05433_),
    .A2(net39),
    .Y(_05437_),
    .B1(_05436_));
 sg13g2_nor2_1 _14533_ (.A(_05424_),
    .B(_05437_),
    .Y(_05438_));
 sg13g2_buf_2 _14534_ (.A(_05438_),
    .X(_05439_));
 sg13g2_inv_2 _14535_ (.Y(_05440_),
    .A(_05439_));
 sg13g2_inv_1 _14536_ (.Y(_05441_),
    .A(_05263_));
 sg13g2_nor3_1 _14537_ (.A(_05441_),
    .B(_05266_),
    .C(net32),
    .Y(_05442_));
 sg13g2_nor2_1 _14538_ (.A(_05442_),
    .B(_05269_),
    .Y(_05443_));
 sg13g2_inv_1 _14539_ (.Y(_05444_),
    .A(_05431_));
 sg13g2_nor2_1 _14540_ (.A(_05443_),
    .B(_05444_),
    .Y(_05445_));
 sg13g2_buf_1 _14541_ (.A(\b.gen_square[57].sq.piece[1] ),
    .X(_05446_));
 sg13g2_inv_1 _14542_ (.Y(_05447_),
    .A(_05446_));
 sg13g2_buf_2 _14543_ (.A(\b.gen_square[57].sq.piece[2] ),
    .X(_05448_));
 sg13g2_buf_2 _14544_ (.A(\b.gen_square[57].sq.piece[0] ),
    .X(_05449_));
 sg13g2_nand3_1 _14545_ (.B(_05448_),
    .C(_05449_),
    .A(_05447_),
    .Y(_05450_));
 sg13g2_buf_2 _14546_ (.A(_05450_),
    .X(_05451_));
 sg13g2_xnor2_1 _14547_ (.Y(_05452_),
    .A(net216),
    .B(\b.gen_square[57].sq.color ));
 sg13g2_buf_2 _14548_ (.A(_05452_),
    .X(_05453_));
 sg13g2_nor2_1 _14549_ (.A(_05451_),
    .B(_05453_),
    .Y(_05454_));
 sg13g2_nand2_1 _14550_ (.Y(_05455_),
    .A(_05454_),
    .B(net168));
 sg13g2_nand3_1 _14551_ (.B(_04063_),
    .C(_03901_),
    .A(_03623_),
    .Y(_05456_));
 sg13g2_inv_1 _14552_ (.Y(_05457_),
    .A(_05448_));
 sg13g2_nand2_1 _14553_ (.Y(_05458_),
    .A(_05446_),
    .B(_05449_));
 sg13g2_nor2_2 _14554_ (.A(_05457_),
    .B(_05458_),
    .Y(_05459_));
 sg13g2_nand3_1 _14555_ (.B(_05456_),
    .C(_05459_),
    .A(_05455_),
    .Y(_05460_));
 sg13g2_inv_1 _14556_ (.Y(_05461_),
    .A(_00026_));
 sg13g2_nand2_1 _14557_ (.Y(_05462_),
    .A(_05460_),
    .B(_05461_));
 sg13g2_buf_1 _14558_ (.A(_05462_),
    .X(_05463_));
 sg13g2_inv_1 _14559_ (.Y(_05464_),
    .A(_05463_));
 sg13g2_nand2_1 _14560_ (.Y(_05465_),
    .A(net147),
    .B(_05453_));
 sg13g2_nand2_1 _14561_ (.Y(_05466_),
    .A(_05455_),
    .B(_05456_));
 sg13g2_inv_1 _14562_ (.Y(_05467_),
    .A(_05466_));
 sg13g2_o21ai_1 _14563_ (.B1(_05467_),
    .Y(_05468_),
    .A1(_05451_),
    .A2(_05465_));
 sg13g2_inv_1 _14564_ (.Y(_05469_),
    .A(_05468_));
 sg13g2_nor2_1 _14565_ (.A(_05464_),
    .B(_05469_),
    .Y(_05470_));
 sg13g2_nor2_1 _14566_ (.A(_05445_),
    .B(_05470_),
    .Y(_05471_));
 sg13g2_nor2b_1 _14567_ (.A(_05203_),
    .B_N(_05471_),
    .Y(_05472_));
 sg13g2_nand3_1 _14568_ (.B(_05446_),
    .C(_05449_),
    .A(_05457_),
    .Y(_05473_));
 sg13g2_nor2_1 _14569_ (.A(_05446_),
    .B(_05449_),
    .Y(_05474_));
 sg13g2_nand2_1 _14570_ (.Y(_05475_),
    .A(_05474_),
    .B(_05448_));
 sg13g2_nand2_1 _14571_ (.Y(_05476_),
    .A(_05473_),
    .B(_05475_));
 sg13g2_nor2b_1 _14572_ (.A(_05465_),
    .B_N(_05476_),
    .Y(_05477_));
 sg13g2_nor2_1 _14573_ (.A(_05477_),
    .B(_05466_),
    .Y(_05478_));
 sg13g2_nor2_1 _14574_ (.A(_05461_),
    .B(_05478_),
    .Y(_05479_));
 sg13g2_nor2_1 _14575_ (.A(_05270_),
    .B(_05444_),
    .Y(_05480_));
 sg13g2_inv_1 _14576_ (.Y(_05481_),
    .A(_05226_));
 sg13g2_inv_2 _14577_ (.Y(_05482_),
    .A(_05214_));
 sg13g2_nor2_1 _14578_ (.A(_05482_),
    .B(net89),
    .Y(_05483_));
 sg13g2_a21oi_2 _14579_ (.B1(_05230_),
    .Y(_05484_),
    .A2(_05483_),
    .A1(_05481_));
 sg13g2_nand2_2 _14580_ (.Y(_05485_),
    .A(_05215_),
    .B(_05216_));
 sg13g2_nor2_2 _14581_ (.A(_05220_),
    .B(_05485_),
    .Y(_05486_));
 sg13g2_nand2_1 _14582_ (.Y(_05487_),
    .A(_05229_),
    .B(_05486_));
 sg13g2_inv_1 _14583_ (.Y(_05488_),
    .A(_00025_));
 sg13g2_nand2_1 _14584_ (.Y(_05489_),
    .A(_05487_),
    .B(_05488_));
 sg13g2_buf_2 _14585_ (.A(_05489_),
    .X(_05490_));
 sg13g2_inv_1 _14586_ (.Y(_05491_),
    .A(_05490_));
 sg13g2_nor2_2 _14587_ (.A(_05484_),
    .B(_05491_),
    .Y(_05492_));
 sg13g2_nor2_1 _14588_ (.A(_05231_),
    .B(_05491_),
    .Y(_05493_));
 sg13g2_nor4_1 _14589_ (.A(_05479_),
    .B(_05480_),
    .C(_05492_),
    .D(_05493_),
    .Y(_05494_));
 sg13g2_nand2_1 _14590_ (.Y(_05495_),
    .A(_05236_),
    .B(_05237_));
 sg13g2_nor2_1 _14591_ (.A(_05235_),
    .B(_05495_),
    .Y(_05496_));
 sg13g2_nand2_1 _14592_ (.Y(_05497_),
    .A(_05249_),
    .B(_05496_));
 sg13g2_inv_1 _14593_ (.Y(_05498_),
    .A(_00062_));
 sg13g2_nand2_1 _14594_ (.Y(_05499_),
    .A(_05497_),
    .B(_05498_));
 sg13g2_buf_2 _14595_ (.A(_05499_),
    .X(_05500_));
 sg13g2_inv_1 _14596_ (.Y(_05501_),
    .A(_05500_));
 sg13g2_nor2_1 _14597_ (.A(_05252_),
    .B(_05501_),
    .Y(_05502_));
 sg13g2_nor2_1 _14598_ (.A(\b.gen_square[48].sq.color ),
    .B(_04740_),
    .Y(_05503_));
 sg13g2_inv_1 _14599_ (.Y(_05504_),
    .A(_04598_));
 sg13g2_a21oi_1 _14600_ (.A1(_05504_),
    .A2(_04733_),
    .Y(_05505_),
    .B1(_04604_));
 sg13g2_buf_1 _14601_ (.A(_05505_),
    .X(_05506_));
 sg13g2_nor2_1 _14602_ (.A(_05506_),
    .B(_04607_),
    .Y(_05507_));
 sg13g2_inv_2 _14603_ (.Y(_05508_),
    .A(_05233_));
 sg13g2_nor3_1 _14604_ (.A(_05508_),
    .B(_05247_),
    .C(net46),
    .Y(_05509_));
 sg13g2_nor2_2 _14605_ (.A(_05509_),
    .B(_05250_),
    .Y(_05510_));
 sg13g2_nor2_1 _14606_ (.A(_05510_),
    .B(_05501_),
    .Y(_05511_));
 sg13g2_inv_1 _14607_ (.Y(_05512_),
    .A(_05511_));
 sg13g2_nand2b_1 _14608_ (.Y(_05513_),
    .B(_05512_),
    .A_N(_05507_));
 sg13g2_nor3_1 _14609_ (.A(_05502_),
    .B(_05503_),
    .C(_05513_),
    .Y(_05514_));
 sg13g2_nand4_1 _14610_ (.B(_05472_),
    .C(_05494_),
    .A(_05440_),
    .Y(_05515_),
    .D(_05514_));
 sg13g2_inv_1 _14611_ (.Y(_05516_),
    .A(_05418_));
 sg13g2_nand2_1 _14612_ (.Y(_05517_),
    .A(_05293_),
    .B(_05292_));
 sg13g2_nor2_1 _14613_ (.A(_05296_),
    .B(_05517_),
    .Y(_05518_));
 sg13g2_nand3_1 _14614_ (.B(_05308_),
    .C(_05518_),
    .A(_05307_),
    .Y(_05519_));
 sg13g2_buf_1 _14615_ (.A(_05519_),
    .X(_05520_));
 sg13g2_inv_1 _14616_ (.Y(_05521_),
    .A(_00020_));
 sg13g2_nand2_1 _14617_ (.Y(_05522_),
    .A(_05520_),
    .B(_05521_));
 sg13g2_a21oi_1 _14618_ (.A1(_05522_),
    .A2(net90),
    .Y(_05523_),
    .B1(_04197_));
 sg13g2_inv_1 _14619_ (.Y(_05524_),
    .A(_05523_));
 sg13g2_inv_1 _14620_ (.Y(_05525_),
    .A(_00046_));
 sg13g2_nor2_1 _14621_ (.A(_05525_),
    .B(_05289_),
    .Y(_05526_));
 sg13g2_buf_1 _14622_ (.A(_05526_),
    .X(_05527_));
 sg13g2_a21oi_1 _14623_ (.A1(_05524_),
    .A2(_05289_),
    .Y(_05528_),
    .B1(_05527_));
 sg13g2_inv_1 _14624_ (.Y(_05529_),
    .A(_05528_));
 sg13g2_inv_1 _14625_ (.Y(_05530_),
    .A(_00052_));
 sg13g2_nor2_1 _14626_ (.A(_05530_),
    .B(net55),
    .Y(_05531_));
 sg13g2_buf_2 _14627_ (.A(_05531_),
    .X(_05532_));
 sg13g2_a21oi_1 _14628_ (.A1(_05529_),
    .A2(net40),
    .Y(_05533_),
    .B1(_05532_));
 sg13g2_inv_1 _14629_ (.Y(_05534_),
    .A(_05533_));
 sg13g2_inv_1 _14630_ (.Y(_05535_),
    .A(_00030_));
 sg13g2_nor2_1 _14631_ (.A(_05535_),
    .B(_05377_),
    .Y(_05536_));
 sg13g2_buf_2 _14632_ (.A(_05536_),
    .X(_05537_));
 sg13g2_a21oi_1 _14633_ (.A1(_05534_),
    .A2(net54),
    .Y(_05538_),
    .B1(_05537_));
 sg13g2_inv_1 _14634_ (.Y(_05539_),
    .A(_05538_));
 sg13g2_a21oi_1 _14635_ (.A1(_05539_),
    .A2(net39),
    .Y(_05540_),
    .B1(_05436_));
 sg13g2_inv_1 _14636_ (.Y(_05541_),
    .A(_04641_));
 sg13g2_a21oi_1 _14637_ (.A1(_04758_),
    .A2(_05541_),
    .Y(_05542_),
    .B1(_04648_));
 sg13g2_buf_2 _14638_ (.A(_05542_),
    .X(_05543_));
 sg13g2_a21oi_1 _14639_ (.A1(_04650_),
    .A2(_05463_),
    .Y(_05544_),
    .B1(_04654_));
 sg13g2_nor2_1 _14640_ (.A(_05543_),
    .B(_05544_),
    .Y(_05545_));
 sg13g2_buf_2 _14641_ (.A(_05545_),
    .X(_05546_));
 sg13g2_buf_1 _14642_ (.A(\b.gen_square[41].sq.piece[1] ),
    .X(_05547_));
 sg13g2_inv_1 _14643_ (.Y(_05548_),
    .A(_05547_));
 sg13g2_buf_2 _14644_ (.A(\b.gen_square[41].sq.piece[2] ),
    .X(_05549_));
 sg13g2_buf_2 _14645_ (.A(\b.gen_square[41].sq.piece[0] ),
    .X(_05550_));
 sg13g2_nand3_1 _14646_ (.B(_05549_),
    .C(_05550_),
    .A(_05548_),
    .Y(_05551_));
 sg13g2_buf_1 _14647_ (.A(_05551_),
    .X(_05552_));
 sg13g2_inv_1 _14648_ (.Y(_05553_),
    .A(_05552_));
 sg13g2_xnor2_1 _14649_ (.Y(_05554_),
    .A(_04035_),
    .B(\b.gen_square[41].sq.color ));
 sg13g2_buf_1 _14650_ (.A(_05554_),
    .X(_05555_));
 sg13g2_inv_1 _14651_ (.Y(_05556_),
    .A(net190));
 sg13g2_nor2_1 _14652_ (.A(_05556_),
    .B(net119),
    .Y(_05557_));
 sg13g2_nor2_1 _14653_ (.A(_05552_),
    .B(_05555_),
    .Y(_05558_));
 sg13g2_a22oi_1 _14654_ (.Y(_05559_),
    .B1(_04063_),
    .B2(_03788_),
    .A2(_04047_),
    .A1(_05558_));
 sg13g2_buf_2 _14655_ (.A(_05559_),
    .X(_05560_));
 sg13g2_inv_4 _14656_ (.A(_05560_),
    .Y(_05561_));
 sg13g2_a21oi_2 _14657_ (.B1(_05561_),
    .Y(_05562_),
    .A2(_05557_),
    .A1(_05553_));
 sg13g2_inv_1 _14658_ (.Y(_05563_),
    .A(_05549_));
 sg13g2_nand2_1 _14659_ (.Y(_05564_),
    .A(_05547_),
    .B(_05550_));
 sg13g2_nor2_1 _14660_ (.A(_05563_),
    .B(_05564_),
    .Y(_05565_));
 sg13g2_inv_1 _14661_ (.Y(_05566_),
    .A(_05565_));
 sg13g2_nor2_1 _14662_ (.A(_05566_),
    .B(_05561_),
    .Y(_05567_));
 sg13g2_buf_8 _14663_ (.A(_05567_),
    .X(_05568_));
 sg13g2_inv_1 _14664_ (.Y(_05569_),
    .A(_00057_));
 sg13g2_nor2_1 _14665_ (.A(_05569_),
    .B(_05568_),
    .Y(_05570_));
 sg13g2_buf_8 _14666_ (.A(_05570_),
    .X(_05571_));
 sg13g2_a21oi_2 _14667_ (.B1(_05571_),
    .Y(_05572_),
    .A2(_05568_),
    .A1(_04608_));
 sg13g2_nor2_2 _14668_ (.A(_05562_),
    .B(_05572_),
    .Y(_05573_));
 sg13g2_nor2_1 _14669_ (.A(_05546_),
    .B(_05573_),
    .Y(_05574_));
 sg13g2_o21ai_1 _14670_ (.B1(_05574_),
    .Y(_05575_),
    .A1(_05516_),
    .A2(_05540_));
 sg13g2_xnor2_1 _14671_ (.Y(_05576_),
    .A(net163),
    .B(\b.gen_square[17].sq.color ));
 sg13g2_buf_2 _14672_ (.A(_05576_),
    .X(_05577_));
 sg13g2_buf_1 _14673_ (.A(\b.gen_square[17].sq.piece[1] ),
    .X(_05578_));
 sg13g2_buf_1 _14674_ (.A(\b.gen_square[17].sq.piece[2] ),
    .X(_05579_));
 sg13g2_buf_1 _14675_ (.A(\b.gen_square[17].sq.piece[0] ),
    .X(_05580_));
 sg13g2_nand3b_1 _14676_ (.B(_05579_),
    .C(_05580_),
    .Y(_05581_),
    .A_N(_05578_));
 sg13g2_buf_2 _14677_ (.A(_05581_),
    .X(_05582_));
 sg13g2_nor2_1 _14678_ (.A(_05577_),
    .B(_05582_),
    .Y(_05583_));
 sg13g2_a22oi_1 _14679_ (.Y(_05584_),
    .B1(net135),
    .B2(_05583_),
    .A2(net117),
    .A1(_03528_));
 sg13g2_buf_1 _14680_ (.A(_05584_),
    .X(_05585_));
 sg13g2_inv_1 _14681_ (.Y(_05586_),
    .A(_05579_));
 sg13g2_nand2_1 _14682_ (.Y(_05587_),
    .A(_05578_),
    .B(_05580_));
 sg13g2_nor2_1 _14683_ (.A(_05586_),
    .B(_05587_),
    .Y(_05588_));
 sg13g2_nand2_1 _14684_ (.Y(_05589_),
    .A(_05585_),
    .B(_05588_));
 sg13g2_buf_2 _14685_ (.A(_05589_),
    .X(_05590_));
 sg13g2_buf_2 _14686_ (.A(\b.gen_square[1].sq.piece[2] ),
    .X(_05591_));
 sg13g2_buf_1 _14687_ (.A(\b.gen_square[1].sq.piece[1] ),
    .X(_05592_));
 sg13g2_buf_1 _14688_ (.A(\b.gen_square[1].sq.piece[0] ),
    .X(_05593_));
 sg13g2_nand2_1 _14689_ (.Y(_05594_),
    .A(_05592_),
    .B(_05593_));
 sg13g2_nor2_1 _14690_ (.A(_05591_),
    .B(_05594_),
    .Y(_05595_));
 sg13g2_inv_1 _14691_ (.Y(_05596_),
    .A(_05591_));
 sg13g2_nor2_1 _14692_ (.A(_05592_),
    .B(_05593_),
    .Y(_05597_));
 sg13g2_inv_1 _14693_ (.Y(_05598_),
    .A(_05597_));
 sg13g2_nor2_1 _14694_ (.A(_05596_),
    .B(_05598_),
    .Y(_05599_));
 sg13g2_nor2_1 _14695_ (.A(_05595_),
    .B(_05599_),
    .Y(_05600_));
 sg13g2_xnor2_1 _14696_ (.Y(_05601_),
    .A(net163),
    .B(_03557_));
 sg13g2_buf_8 _14697_ (.A(_05601_),
    .X(_05602_));
 sg13g2_inv_1 _14698_ (.Y(_05603_),
    .A(_05602_));
 sg13g2_nor2_1 _14699_ (.A(_05603_),
    .B(net89),
    .Y(_05604_));
 sg13g2_inv_1 _14700_ (.Y(_05605_),
    .A(_05604_));
 sg13g2_nor2_1 _14701_ (.A(_05600_),
    .B(_05605_),
    .Y(_05606_));
 sg13g2_inv_1 _14702_ (.Y(_05607_),
    .A(_05593_));
 sg13g2_nor3_2 _14703_ (.A(_05592_),
    .B(_05596_),
    .C(_05607_),
    .Y(_05608_));
 sg13g2_nor2b_1 _14704_ (.A(_05602_),
    .B_N(_05608_),
    .Y(_05609_));
 sg13g2_a22oi_1 _14705_ (.Y(_05610_),
    .B1(net135),
    .B2(_05609_),
    .A2(net134),
    .A1(_03559_));
 sg13g2_inv_2 _14706_ (.Y(_05611_),
    .A(_05610_));
 sg13g2_nor2_1 _14707_ (.A(_05606_),
    .B(_05611_),
    .Y(_05612_));
 sg13g2_nor2_1 _14708_ (.A(_04817_),
    .B(_04821_),
    .Y(_05613_));
 sg13g2_o21ai_1 _14709_ (.B1(_04864_),
    .Y(_05614_),
    .A1(_04861_),
    .A2(_05613_));
 sg13g2_nand3_1 _14710_ (.B(_04823_),
    .C(_05614_),
    .A(_04831_),
    .Y(_05615_));
 sg13g2_inv_1 _14711_ (.Y(_05616_),
    .A(_05615_));
 sg13g2_a21oi_1 _14712_ (.A1(net43),
    .A2(_05612_),
    .Y(_05617_),
    .B1(_05616_));
 sg13g2_nor2_1 _14713_ (.A(_05578_),
    .B(_05580_),
    .Y(_05618_));
 sg13g2_inv_1 _14714_ (.Y(_05619_),
    .A(_05618_));
 sg13g2_nor2_1 _14715_ (.A(_05586_),
    .B(_05619_),
    .Y(_05620_));
 sg13g2_nor2_1 _14716_ (.A(_05579_),
    .B(_05587_),
    .Y(_05621_));
 sg13g2_inv_1 _14717_ (.Y(_05622_),
    .A(_05577_));
 sg13g2_nor2_1 _14718_ (.A(_05622_),
    .B(net79),
    .Y(_05623_));
 sg13g2_o21ai_1 _14719_ (.B1(_05623_),
    .Y(_05624_),
    .A1(_05620_),
    .A2(_05621_));
 sg13g2_inv_1 _14720_ (.Y(_05625_),
    .A(_05588_));
 sg13g2_nand3_1 _14721_ (.B(_05624_),
    .C(_05625_),
    .A(_05585_),
    .Y(_05626_));
 sg13g2_buf_1 _14722_ (.A(_05626_),
    .X(_05627_));
 sg13g2_o21ai_1 _14723_ (.B1(_05627_),
    .Y(_05628_),
    .A1(_05590_),
    .A2(_05617_));
 sg13g2_buf_1 _14724_ (.A(\b.gen_square[25].sq.piece[2] ),
    .X(_05629_));
 sg13g2_inv_1 _14725_ (.Y(_05630_),
    .A(_05629_));
 sg13g2_buf_1 _14726_ (.A(\b.gen_square[25].sq.piece[1] ),
    .X(_05631_));
 sg13g2_buf_1 _14727_ (.A(\b.gen_square[25].sq.piece[0] ),
    .X(_05632_));
 sg13g2_nand2_1 _14728_ (.Y(_05633_),
    .A(_05631_),
    .B(_05632_));
 sg13g2_nor2_1 _14729_ (.A(_05630_),
    .B(_05633_),
    .Y(_05634_));
 sg13g2_inv_1 _14730_ (.Y(_05635_),
    .A(_05634_));
 sg13g2_xnor2_1 _14731_ (.Y(_05636_),
    .A(net179),
    .B(\b.gen_square[25].sq.color ));
 sg13g2_buf_2 _14732_ (.A(_05636_),
    .X(_05637_));
 sg13g2_inv_1 _14733_ (.Y(_05638_),
    .A(_05632_));
 sg13g2_nor3_1 _14734_ (.A(_05631_),
    .B(_05630_),
    .C(_05638_),
    .Y(_05639_));
 sg13g2_inv_1 _14735_ (.Y(_05640_),
    .A(_05639_));
 sg13g2_nor2_1 _14736_ (.A(_05637_),
    .B(_05640_),
    .Y(_05641_));
 sg13g2_a22oi_1 _14737_ (.Y(_05642_),
    .B1(net152),
    .B2(_05641_),
    .A2(net134),
    .A1(_03625_));
 sg13g2_buf_1 _14738_ (.A(_05642_),
    .X(_05643_));
 sg13g2_inv_1 _14739_ (.Y(_05644_),
    .A(_05643_));
 sg13g2_nor2_1 _14740_ (.A(_05635_),
    .B(_05644_),
    .Y(_05645_));
 sg13g2_buf_2 _14741_ (.A(_05645_),
    .X(_05646_));
 sg13g2_buf_1 _14742_ (.A(_05646_),
    .X(_05647_));
 sg13g2_nor2_1 _14743_ (.A(_05631_),
    .B(_05632_),
    .Y(_05648_));
 sg13g2_inv_1 _14744_ (.Y(_05649_),
    .A(_05648_));
 sg13g2_nor2_2 _14745_ (.A(_05630_),
    .B(_05649_),
    .Y(_05650_));
 sg13g2_nor2_1 _14746_ (.A(_05629_),
    .B(_05633_),
    .Y(_05651_));
 sg13g2_inv_1 _14747_ (.Y(_05652_),
    .A(_05637_));
 sg13g2_nor2_1 _14748_ (.A(_05652_),
    .B(_04286_),
    .Y(_05653_));
 sg13g2_o21ai_1 _14749_ (.B1(_05653_),
    .Y(_05654_),
    .A1(_05650_),
    .A2(_05651_));
 sg13g2_nand3_1 _14750_ (.B(_05635_),
    .C(_05654_),
    .A(_05643_),
    .Y(_05655_));
 sg13g2_buf_1 _14751_ (.A(_05655_),
    .X(_05656_));
 sg13g2_inv_1 _14752_ (.Y(_05657_),
    .A(_05656_));
 sg13g2_a21oi_1 _14753_ (.A1(_05628_),
    .A2(net53),
    .Y(_05658_),
    .B1(_05657_));
 sg13g2_inv_1 _14754_ (.Y(_05659_),
    .A(_05658_));
 sg13g2_buf_2 _14755_ (.A(\b.gen_square[33].sq.piece[2] ),
    .X(_05660_));
 sg13g2_inv_2 _14756_ (.Y(_05661_),
    .A(_05660_));
 sg13g2_buf_2 _14757_ (.A(\b.gen_square[33].sq.piece[1] ),
    .X(_05662_));
 sg13g2_buf_1 _14758_ (.A(\b.gen_square[33].sq.piece[0] ),
    .X(_05663_));
 sg13g2_nand2_1 _14759_ (.Y(_05664_),
    .A(_05662_),
    .B(_05663_));
 sg13g2_nor2_1 _14760_ (.A(_05661_),
    .B(_05664_),
    .Y(_05665_));
 sg13g2_inv_2 _14761_ (.Y(_05666_),
    .A(_05665_));
 sg13g2_xnor2_1 _14762_ (.Y(_05667_),
    .A(net216),
    .B(\b.gen_square[33].sq.color ));
 sg13g2_buf_8 _14763_ (.A(_05667_),
    .X(_05668_));
 sg13g2_inv_2 _14764_ (.Y(_05669_),
    .A(_05663_));
 sg13g2_nor3_1 _14765_ (.A(_05662_),
    .B(_05661_),
    .C(_05669_),
    .Y(_05670_));
 sg13g2_inv_1 _14766_ (.Y(_05671_),
    .A(_05670_));
 sg13g2_nor2_1 _14767_ (.A(_05668_),
    .B(_05671_),
    .Y(_05672_));
 sg13g2_a22oi_1 _14768_ (.Y(_05673_),
    .B1(net168),
    .B2(_05672_),
    .A2(net167),
    .A1(_03706_));
 sg13g2_buf_2 _14769_ (.A(_05673_),
    .X(_05674_));
 sg13g2_inv_4 _14770_ (.A(_05674_),
    .Y(_05675_));
 sg13g2_nor2_1 _14771_ (.A(_05666_),
    .B(_05675_),
    .Y(_05676_));
 sg13g2_buf_8 _14772_ (.A(_05676_),
    .X(_05677_));
 sg13g2_buf_1 _14773_ (.A(_05677_),
    .X(_05678_));
 sg13g2_inv_1 _14774_ (.Y(_05679_),
    .A(_05668_));
 sg13g2_nor2_1 _14775_ (.A(_05679_),
    .B(net100),
    .Y(_05680_));
 sg13g2_nor2_1 _14776_ (.A(_05660_),
    .B(_05664_),
    .Y(_05681_));
 sg13g2_nor2_1 _14777_ (.A(_05662_),
    .B(_05663_),
    .Y(_05682_));
 sg13g2_nand2_1 _14778_ (.Y(_05683_),
    .A(_05682_),
    .B(_05660_));
 sg13g2_nand2b_1 _14779_ (.Y(_05684_),
    .B(_05683_),
    .A_N(_05681_));
 sg13g2_nand2_1 _14780_ (.Y(_05685_),
    .A(_05680_),
    .B(_05684_));
 sg13g2_nand3_1 _14781_ (.B(_05666_),
    .C(_05685_),
    .A(_05674_),
    .Y(_05686_));
 sg13g2_buf_1 _14782_ (.A(_05686_),
    .X(_05687_));
 sg13g2_inv_1 _14783_ (.Y(_05688_),
    .A(_05687_));
 sg13g2_a21oi_2 _14784_ (.B1(_05688_),
    .Y(_05689_),
    .A2(net74),
    .A1(_05659_));
 sg13g2_inv_1 _14785_ (.Y(_05690_),
    .A(_05689_));
 sg13g2_buf_1 _14786_ (.A(_05568_),
    .X(_05691_));
 sg13g2_nor2_1 _14787_ (.A(_05549_),
    .B(_05564_),
    .Y(_05692_));
 sg13g2_nor2_1 _14788_ (.A(_05547_),
    .B(_05550_),
    .Y(_05693_));
 sg13g2_nand2_1 _14789_ (.Y(_05694_),
    .A(_05693_),
    .B(_05549_));
 sg13g2_nand2b_1 _14790_ (.Y(_05695_),
    .B(_05694_),
    .A_N(_05692_));
 sg13g2_nand2_1 _14791_ (.Y(_05696_),
    .A(_05557_),
    .B(_05695_));
 sg13g2_nand3_1 _14792_ (.B(_05566_),
    .C(_05696_),
    .A(_05560_),
    .Y(_05697_));
 sg13g2_inv_1 _14793_ (.Y(_05698_),
    .A(_05697_));
 sg13g2_a21oi_1 _14794_ (.A1(_05690_),
    .A2(net52),
    .Y(_05699_),
    .B1(_05698_));
 sg13g2_inv_1 _14795_ (.Y(_05700_),
    .A(_05699_));
 sg13g2_nor2_2 _14796_ (.A(_05596_),
    .B(_05594_),
    .Y(_05701_));
 sg13g2_inv_1 _14797_ (.Y(_05702_),
    .A(_05701_));
 sg13g2_nor2_1 _14798_ (.A(_05702_),
    .B(_05611_),
    .Y(_05703_));
 sg13g2_buf_2 _14799_ (.A(_05703_),
    .X(_05704_));
 sg13g2_nor2_1 _14800_ (.A(_03558_),
    .B(_05704_),
    .Y(_05705_));
 sg13g2_inv_2 _14801_ (.Y(_05706_),
    .A(_05705_));
 sg13g2_a21oi_1 _14802_ (.A1(_05706_),
    .A2(net43),
    .Y(_05707_),
    .B1(_04956_));
 sg13g2_inv_1 _14803_ (.Y(_05708_),
    .A(_05707_));
 sg13g2_inv_2 _14804_ (.Y(_05709_),
    .A(_05590_));
 sg13g2_buf_8 _14805_ (.A(_05709_),
    .X(_05710_));
 sg13g2_nand2_1 _14806_ (.Y(_05711_),
    .A(_05590_),
    .B(_00032_));
 sg13g2_buf_2 _14807_ (.A(_05711_),
    .X(_05712_));
 sg13g2_inv_4 _14808_ (.A(_05712_),
    .Y(_05713_));
 sg13g2_a21oi_2 _14809_ (.B1(_05713_),
    .Y(_05714_),
    .A2(net38),
    .A1(_05708_));
 sg13g2_inv_1 _14810_ (.Y(_05715_),
    .A(_05714_));
 sg13g2_inv_1 _14811_ (.Y(_05716_),
    .A(_00043_));
 sg13g2_nor2_1 _14812_ (.A(_05716_),
    .B(_05646_),
    .Y(_05717_));
 sg13g2_buf_8 _14813_ (.A(_05717_),
    .X(_05718_));
 sg13g2_a21oi_2 _14814_ (.B1(_05718_),
    .Y(_05719_),
    .A2(net53),
    .A1(_05715_));
 sg13g2_inv_1 _14815_ (.Y(_05720_),
    .A(_05719_));
 sg13g2_inv_1 _14816_ (.Y(_05721_),
    .A(_00051_));
 sg13g2_nor2_1 _14817_ (.A(_05721_),
    .B(_05677_),
    .Y(_05722_));
 sg13g2_buf_2 _14818_ (.A(_05722_),
    .X(_05723_));
 sg13g2_a21oi_1 _14819_ (.A1(_05720_),
    .A2(net74),
    .Y(_05724_),
    .B1(_05723_));
 sg13g2_inv_1 _14820_ (.Y(_05725_),
    .A(_05724_));
 sg13g2_a21oi_1 _14821_ (.A1(_05725_),
    .A2(net52),
    .Y(_05726_),
    .B1(_05571_));
 sg13g2_buf_1 _14822_ (.A(net98),
    .X(_05727_));
 sg13g2_inv_1 _14823_ (.Y(_05728_),
    .A(_05049_));
 sg13g2_a21oi_1 _14824_ (.A1(_05058_),
    .A2(net84),
    .Y(_05729_),
    .B1(_05728_));
 sg13g2_inv_1 _14825_ (.Y(_05730_),
    .A(_05729_));
 sg13g2_a21oi_1 _14826_ (.A1(_05730_),
    .A2(net77),
    .Y(_05731_),
    .B1(_04728_));
 sg13g2_inv_1 _14827_ (.Y(_05732_),
    .A(_05731_));
 sg13g2_a21oi_1 _14828_ (.A1(_05732_),
    .A2(net30),
    .Y(_05733_),
    .B1(_04702_));
 sg13g2_inv_1 _14829_ (.Y(_05734_),
    .A(_05733_));
 sg13g2_a21oi_1 _14830_ (.A1(_05734_),
    .A2(_04674_),
    .Y(_05735_),
    .B1(_04678_));
 sg13g2_inv_1 _14831_ (.Y(_05736_),
    .A(_05735_));
 sg13g2_a21oi_1 _14832_ (.A1(_05736_),
    .A2(net45),
    .Y(_05737_),
    .B1(_04654_));
 sg13g2_inv_1 _14833_ (.Y(_05738_),
    .A(_05737_));
 sg13g2_nand2_1 _14834_ (.Y(_05739_),
    .A(net147),
    .B(net180));
 sg13g2_o21ai_1 _14835_ (.B1(_05105_),
    .Y(_05740_),
    .A1(_05031_),
    .A2(_05035_));
 sg13g2_nor2b_1 _14836_ (.A(_05739_),
    .B_N(_05740_),
    .Y(_05741_));
 sg13g2_inv_1 _14837_ (.Y(_05742_),
    .A(_05044_));
 sg13g2_nand3b_1 _14838_ (.B(_05742_),
    .C(_05037_),
    .Y(_05743_),
    .A_N(_05741_));
 sg13g2_inv_1 _14839_ (.Y(_05744_),
    .A(_05743_));
 sg13g2_a21oi_1 _14840_ (.A1(net98),
    .A2(_04356_),
    .Y(_05745_),
    .B1(_05744_));
 sg13g2_inv_1 _14841_ (.Y(_05746_),
    .A(_05745_));
 sg13g2_a21oi_1 _14842_ (.A1(_05746_),
    .A2(_04723_),
    .Y(_05747_),
    .B1(_04796_));
 sg13g2_inv_1 _14843_ (.Y(_05748_),
    .A(_05747_));
 sg13g2_a21oi_1 _14844_ (.A1(_05748_),
    .A2(net30),
    .Y(_05749_),
    .B1(_04787_));
 sg13g2_inv_1 _14845_ (.Y(_05750_),
    .A(_05749_));
 sg13g2_a21oi_1 _14846_ (.A1(_05750_),
    .A2(net44),
    .Y(_05751_),
    .B1(_04776_));
 sg13g2_inv_1 _14847_ (.Y(_05752_),
    .A(_05751_));
 sg13g2_a21oi_1 _14848_ (.A1(_05752_),
    .A2(net45),
    .Y(_05753_),
    .B1(_04765_));
 sg13g2_nand2_1 _14849_ (.Y(_05754_),
    .A(_05738_),
    .B(_05753_));
 sg13g2_o21ai_1 _14850_ (.B1(_05754_),
    .Y(_05755_),
    .A1(_05700_),
    .A2(_05726_));
 sg13g2_nor3_1 _14851_ (.A(_05515_),
    .B(_05575_),
    .C(_05755_),
    .Y(_05756_));
 sg13g2_inv_1 _14852_ (.Y(_05757_),
    .A(_05407_));
 sg13g2_a21oi_1 _14853_ (.A1(_05490_),
    .A2(_04650_),
    .Y(_05758_),
    .B1(_04654_));
 sg13g2_inv_1 _14854_ (.Y(_05759_),
    .A(_05436_));
 sg13g2_o21ai_1 _14855_ (.B1(_05759_),
    .Y(_05760_),
    .A1(_05757_),
    .A2(_05758_));
 sg13g2_buf_1 _14856_ (.A(_05760_),
    .X(_05761_));
 sg13g2_nor2_1 _14857_ (.A(_05424_),
    .B(_05761_),
    .Y(_05762_));
 sg13g2_buf_2 _14858_ (.A(_05762_),
    .X(_05763_));
 sg13g2_inv_1 _14859_ (.Y(_05764_),
    .A(_05763_));
 sg13g2_nor2_1 _14860_ (.A(_05490_),
    .B(_05484_),
    .Y(_05765_));
 sg13g2_inv_1 _14861_ (.Y(_05766_),
    .A(_05765_));
 sg13g2_inv_1 _14862_ (.Y(_05767_),
    .A(_05544_));
 sg13g2_nor2_2 _14863_ (.A(_05543_),
    .B(_05767_),
    .Y(_05768_));
 sg13g2_a21oi_1 _14864_ (.A1(_05500_),
    .A2(_05568_),
    .Y(_05769_),
    .B1(_05571_));
 sg13g2_inv_1 _14865_ (.Y(_05770_),
    .A(_05769_));
 sg13g2_nor2_1 _14866_ (.A(_05562_),
    .B(_05770_),
    .Y(_05771_));
 sg13g2_nor2_1 _14867_ (.A(_05768_),
    .B(_05771_),
    .Y(_05772_));
 sg13g2_nand3_1 _14868_ (.B(_05766_),
    .C(_05772_),
    .A(_05764_),
    .Y(_05773_));
 sg13g2_nand2_1 _14869_ (.Y(_05774_),
    .A(_05540_),
    .B(_05418_));
 sg13g2_nor2_1 _14870_ (.A(_05270_),
    .B(_05431_),
    .Y(_05775_));
 sg13g2_nor2_1 _14871_ (.A(_05506_),
    .B(_04608_),
    .Y(_05776_));
 sg13g2_nor2_1 _14872_ (.A(_05490_),
    .B(_05231_),
    .Y(_05777_));
 sg13g2_nor3_1 _14873_ (.A(_05775_),
    .B(_05776_),
    .C(_05777_),
    .Y(_05778_));
 sg13g2_nor2_1 _14874_ (.A(_05510_),
    .B(_05500_),
    .Y(_05779_));
 sg13g2_nor2_1 _14875_ (.A(_05500_),
    .B(_05252_),
    .Y(_05780_));
 sg13g2_nor2_1 _14876_ (.A(_05443_),
    .B(_05431_),
    .Y(_05781_));
 sg13g2_nor2_1 _14877_ (.A(_05463_),
    .B(_05469_),
    .Y(_05782_));
 sg13g2_nor2_1 _14878_ (.A(_05781_),
    .B(_05782_),
    .Y(_05783_));
 sg13g2_inv_1 _14879_ (.Y(_05784_),
    .A(_05783_));
 sg13g2_nor3_1 _14880_ (.A(_05779_),
    .B(_05780_),
    .C(_05784_),
    .Y(_05785_));
 sg13g2_nand4_1 _14881_ (.B(_05211_),
    .C(_05778_),
    .A(_05774_),
    .Y(_05786_),
    .D(_05785_));
 sg13g2_inv_1 _14882_ (.Y(_05787_),
    .A(_05753_));
 sg13g2_nor2_1 _14883_ (.A(_05738_),
    .B(_05787_),
    .Y(_05788_));
 sg13g2_nor2_1 _14884_ (.A(_00026_),
    .B(_05478_),
    .Y(_05789_));
 sg13g2_nor2_1 _14885_ (.A(_03847_),
    .B(_04740_),
    .Y(_05790_));
 sg13g2_nor2b_1 _14886_ (.A(_05700_),
    .B_N(_05726_),
    .Y(_05791_));
 sg13g2_nor4_1 _14887_ (.A(_05788_),
    .B(_05789_),
    .C(_05790_),
    .D(_05791_),
    .Y(_05792_));
 sg13g2_inv_1 _14888_ (.Y(_05793_),
    .A(_05792_));
 sg13g2_nor3_1 _14889_ (.A(_05773_),
    .B(_05786_),
    .C(_05793_),
    .Y(_05794_));
 sg13g2_nor3_1 _14890_ (.A(_05124_),
    .B(_05756_),
    .C(_05794_),
    .Y(_05795_));
 sg13g2_nand2_1 _14891_ (.Y(_05796_),
    .A(_05795_),
    .B(net162));
 sg13g2_nand2_1 _14892_ (.Y(_05797_),
    .A(_05794_),
    .B(_05756_));
 sg13g2_nand3_1 _14893_ (.B(net96),
    .C(_04621_),
    .A(_05797_),
    .Y(_05798_));
 sg13g2_nand2_1 _14894_ (.Y(_05799_),
    .A(_05796_),
    .B(_05798_));
 sg13g2_a22oi_1 _14895_ (.Y(_05800_),
    .B1(_05423_),
    .B2(_05799_),
    .A2(_05422_),
    .A1(_05123_));
 sg13g2_nor3_1 _14896_ (.A(_05479_),
    .B(_05503_),
    .C(_05755_),
    .Y(_05801_));
 sg13g2_a21oi_1 _14897_ (.A1(_05792_),
    .A2(_05801_),
    .Y(_05802_),
    .B1(_04621_));
 sg13g2_inv_1 _14898_ (.Y(_05803_),
    .A(_05802_));
 sg13g2_a21o_1 _14899_ (.A2(_05419_),
    .A1(_05803_),
    .B1(_04750_),
    .X(_05804_));
 sg13g2_o21ai_1 _14900_ (.B1(_05804_),
    .Y(_05805_),
    .A1(_04748_),
    .A2(_05803_));
 sg13g2_nand2_1 _14901_ (.Y(_05806_),
    .A(_05805_),
    .B(net95));
 sg13g2_nand2_1 _14902_ (.Y(_05807_),
    .A(_05800_),
    .B(_05806_));
 sg13g2_buf_1 _14903_ (.A(\b.gen_square[49].sq.mask ),
    .X(_05808_));
 sg13g2_nand2_1 _14904_ (.Y(_05809_),
    .A(_05807_),
    .B(_05808_));
 sg13g2_nor2_1 _14905_ (.A(net103),
    .B(_05504_),
    .Y(_05810_));
 sg13g2_nor3_1 _14906_ (.A(_05660_),
    .B(_05662_),
    .C(_05669_),
    .Y(_05811_));
 sg13g2_nand2_1 _14907_ (.Y(_05812_),
    .A(_05668_),
    .B(_05811_));
 sg13g2_inv_1 _14908_ (.Y(_05813_),
    .A(_05812_));
 sg13g2_a21oi_1 _14909_ (.A1(_04509_),
    .A2(_05813_),
    .Y(_05814_),
    .B1(_05675_));
 sg13g2_nor2_2 _14910_ (.A(_03705_),
    .B(_05814_),
    .Y(_05815_));
 sg13g2_nor3_1 _14911_ (.A(_05390_),
    .B(_05392_),
    .C(_05399_),
    .Y(_05816_));
 sg13g2_nand2_1 _14912_ (.Y(_05817_),
    .A(_05398_),
    .B(_05816_));
 sg13g2_inv_1 _14913_ (.Y(_05818_),
    .A(_05817_));
 sg13g2_a21oi_1 _14914_ (.A1(net99),
    .A2(_05818_),
    .Y(_05819_),
    .B1(_05405_));
 sg13g2_nand4_1 _14915_ (.B(_05220_),
    .C(_05224_),
    .A(_05214_),
    .Y(_05820_),
    .D(_05216_));
 sg13g2_inv_1 _14916_ (.Y(_05821_),
    .A(_05820_));
 sg13g2_a21oi_1 _14917_ (.A1(net78),
    .A2(_05821_),
    .Y(_05822_),
    .B1(_05230_));
 sg13g2_nor2_1 _14918_ (.A(_03941_),
    .B(_05822_),
    .Y(_05823_));
 sg13g2_inv_1 _14919_ (.Y(_05824_),
    .A(_05823_));
 sg13g2_o21ai_1 _14920_ (.B1(_05824_),
    .Y(_05825_),
    .A1(_03795_),
    .A2(_05819_));
 sg13g2_nor2_1 _14921_ (.A(_05815_),
    .B(_05825_),
    .Y(_05826_));
 sg13g2_nor2_1 _14922_ (.A(_05721_),
    .B(_05814_),
    .Y(_05827_));
 sg13g2_buf_2 _14923_ (.A(_05827_),
    .X(_05828_));
 sg13g2_nor2_1 _14924_ (.A(_05434_),
    .B(_05819_),
    .Y(_05829_));
 sg13g2_inv_1 _14925_ (.Y(_05830_),
    .A(_05829_));
 sg13g2_nor2_1 _14926_ (.A(_05488_),
    .B(_05822_),
    .Y(_05831_));
 sg13g2_inv_1 _14927_ (.Y(_05832_),
    .A(_05831_));
 sg13g2_nand2_2 _14928_ (.Y(_05833_),
    .A(_05830_),
    .B(_05832_));
 sg13g2_nor2_1 _14929_ (.A(_05828_),
    .B(_05833_),
    .Y(_05834_));
 sg13g2_inv_1 _14930_ (.Y(_05835_),
    .A(_04592_));
 sg13g2_nor3_1 _14931_ (.A(_04589_),
    .B(_04591_),
    .C(_05835_),
    .Y(_05836_));
 sg13g2_nand2_1 _14932_ (.Y(_05837_),
    .A(_04600_),
    .B(_05836_));
 sg13g2_a21oi_1 _14933_ (.A1(_05826_),
    .A2(_05834_),
    .Y(_05838_),
    .B1(_05837_));
 sg13g2_nand3_1 _14934_ (.B(_05835_),
    .C(_04591_),
    .A(_04590_),
    .Y(_05839_));
 sg13g2_nand2_1 _14935_ (.Y(_05840_),
    .A(_05131_),
    .B(_05132_));
 sg13g2_nor2_1 _14936_ (.A(_05137_),
    .B(_05840_),
    .Y(_05841_));
 sg13g2_inv_1 _14937_ (.Y(_05842_),
    .A(_05841_));
 sg13g2_nor2_1 _14938_ (.A(_05842_),
    .B(_05143_),
    .Y(_05843_));
 sg13g2_buf_2 _14939_ (.A(_05843_),
    .X(_05844_));
 sg13g2_inv_1 _14940_ (.Y(_05845_),
    .A(_05844_));
 sg13g2_buf_2 _14941_ (.A(\b.gen_square[20].sq.piece[2] ),
    .X(_05846_));
 sg13g2_inv_1 _14942_ (.Y(_05847_),
    .A(_05846_));
 sg13g2_buf_1 _14943_ (.A(\b.gen_square[20].sq.piece[1] ),
    .X(_05848_));
 sg13g2_buf_2 _14944_ (.A(\b.gen_square[20].sq.piece[0] ),
    .X(_05849_));
 sg13g2_nand2_1 _14945_ (.Y(_05850_),
    .A(_05848_),
    .B(_05849_));
 sg13g2_nor2_1 _14946_ (.A(_05847_),
    .B(_05850_),
    .Y(_05851_));
 sg13g2_inv_1 _14947_ (.Y(_05852_),
    .A(_05851_));
 sg13g2_xnor2_1 _14948_ (.Y(_05853_),
    .A(_04079_),
    .B(\b.gen_square[20].sq.color ));
 sg13g2_buf_2 _14949_ (.A(_05853_),
    .X(_05854_));
 sg13g2_inv_1 _14950_ (.Y(_05855_),
    .A(_05849_));
 sg13g2_nor3_2 _14951_ (.A(_05848_),
    .B(_05847_),
    .C(_05855_),
    .Y(_05856_));
 sg13g2_inv_1 _14952_ (.Y(_05857_),
    .A(_05856_));
 sg13g2_nor2_1 _14953_ (.A(_05854_),
    .B(_05857_),
    .Y(_05858_));
 sg13g2_a22oi_1 _14954_ (.Y(_05859_),
    .B1(_04090_),
    .B2(_03572_),
    .A2(_04086_),
    .A1(_05858_));
 sg13g2_buf_1 _14955_ (.A(_05859_),
    .X(_05860_));
 sg13g2_inv_1 _14956_ (.Y(_05861_),
    .A(_05860_));
 sg13g2_nor2_1 _14957_ (.A(_05852_),
    .B(_05861_),
    .Y(_05862_));
 sg13g2_buf_2 _14958_ (.A(_05862_),
    .X(_05863_));
 sg13g2_inv_2 _14959_ (.Y(_05864_),
    .A(_05863_));
 sg13g2_inv_1 _14960_ (.Y(_05865_),
    .A(_04167_));
 sg13g2_nor2_1 _14961_ (.A(_05865_),
    .B(_04348_),
    .Y(_05866_));
 sg13g2_inv_1 _14962_ (.Y(_05867_),
    .A(_05866_));
 sg13g2_nor2_1 _14963_ (.A(_04159_),
    .B(_04163_),
    .Y(_05868_));
 sg13g2_inv_1 _14964_ (.Y(_05869_),
    .A(_04266_));
 sg13g2_a21oi_1 _14965_ (.A1(_04157_),
    .A2(_05868_),
    .Y(_05870_),
    .B1(_05869_));
 sg13g2_o21ai_1 _14966_ (.B1(_04258_),
    .Y(_05871_),
    .A1(_05867_),
    .A2(_05870_));
 sg13g2_inv_1 _14967_ (.Y(_05872_),
    .A(_05871_));
 sg13g2_buf_2 _14968_ (.A(\b.gen_square[13].sq.piece[2] ),
    .X(_05873_));
 sg13g2_inv_1 _14969_ (.Y(_05874_),
    .A(_05873_));
 sg13g2_buf_1 _14970_ (.A(\b.gen_square[13].sq.piece[1] ),
    .X(_05875_));
 sg13g2_buf_2 _14971_ (.A(\b.gen_square[13].sq.piece[0] ),
    .X(_05876_));
 sg13g2_nand2_1 _14972_ (.Y(_05877_),
    .A(_05875_),
    .B(_05876_));
 sg13g2_nor2_1 _14973_ (.A(_05874_),
    .B(_05877_),
    .Y(_05878_));
 sg13g2_inv_1 _14974_ (.Y(_05879_),
    .A(_05878_));
 sg13g2_inv_1 _14975_ (.Y(_05880_),
    .A(_05875_));
 sg13g2_nand3_1 _14976_ (.B(_05873_),
    .C(_05876_),
    .A(_05880_),
    .Y(_05881_));
 sg13g2_buf_2 _14977_ (.A(_05881_),
    .X(_05882_));
 sg13g2_xnor2_1 _14978_ (.Y(_05883_),
    .A(_04039_),
    .B(\b.gen_square[13].sq.color ));
 sg13g2_buf_2 _14979_ (.A(_05883_),
    .X(_05884_));
 sg13g2_nor2_1 _14980_ (.A(_05882_),
    .B(_05884_),
    .Y(_05885_));
 sg13g2_a22oi_1 _14981_ (.Y(_05886_),
    .B1(_04064_),
    .B2(_02994_),
    .A2(_04243_),
    .A1(_05885_));
 sg13g2_buf_1 _14982_ (.A(_05886_),
    .X(_05887_));
 sg13g2_inv_4 _14983_ (.A(_05887_),
    .Y(_05888_));
 sg13g2_nor2_1 _14984_ (.A(_05879_),
    .B(_05888_),
    .Y(_05889_));
 sg13g2_buf_1 _14985_ (.A(_05889_),
    .X(_05890_));
 sg13g2_inv_1 _14986_ (.Y(_05891_),
    .A(_05884_));
 sg13g2_nor2_1 _14987_ (.A(_05891_),
    .B(_04051_),
    .Y(_05892_));
 sg13g2_nor3_1 _14988_ (.A(_05873_),
    .B(_05876_),
    .C(_05880_),
    .Y(_05893_));
 sg13g2_nor2_1 _14989_ (.A(_05875_),
    .B(_05876_),
    .Y(_05894_));
 sg13g2_nand2_1 _14990_ (.Y(_05895_),
    .A(_05894_),
    .B(_05873_));
 sg13g2_nand2b_1 _14991_ (.Y(_05896_),
    .B(_05895_),
    .A_N(_05893_));
 sg13g2_nand2_1 _14992_ (.Y(_05897_),
    .A(_05892_),
    .B(_05896_));
 sg13g2_nand3_1 _14993_ (.B(_05879_),
    .C(_05897_),
    .A(_05887_),
    .Y(_05898_));
 sg13g2_inv_1 _14994_ (.Y(_05899_),
    .A(_05898_));
 sg13g2_a21oi_1 _14995_ (.A1(_05872_),
    .A2(net73),
    .Y(_05900_),
    .B1(_05899_));
 sg13g2_nor2_1 _14996_ (.A(_05848_),
    .B(_05849_),
    .Y(_05901_));
 sg13g2_nand2_1 _14997_ (.Y(_05902_),
    .A(_05901_),
    .B(_05846_));
 sg13g2_and3_1 _14998_ (.X(_05903_),
    .A(_05847_),
    .B(_05855_),
    .C(_05848_));
 sg13g2_inv_1 _14999_ (.Y(_05904_),
    .A(_05903_));
 sg13g2_inv_1 _15000_ (.Y(_05905_),
    .A(_05854_));
 sg13g2_nor2_1 _15001_ (.A(_05905_),
    .B(_04300_),
    .Y(_05906_));
 sg13g2_inv_1 _15002_ (.Y(_05907_),
    .A(_05906_));
 sg13g2_a21o_1 _15003_ (.A2(_05904_),
    .A1(_05902_),
    .B1(_05907_),
    .X(_05908_));
 sg13g2_nand3_1 _15004_ (.B(_05860_),
    .C(_05852_),
    .A(_05908_),
    .Y(_05909_));
 sg13g2_buf_1 _15005_ (.A(_05909_),
    .X(_05910_));
 sg13g2_o21ai_1 _15006_ (.B1(_05910_),
    .Y(_05911_),
    .A1(_05864_),
    .A2(_05900_));
 sg13g2_buf_1 _15007_ (.A(_05911_),
    .X(_05912_));
 sg13g2_a21oi_2 _15008_ (.B1(_04907_),
    .Y(_05913_),
    .A2(net42),
    .A1(_05912_));
 sg13g2_nor2_1 _15009_ (.A(_05131_),
    .B(_05132_),
    .Y(_05914_));
 sg13g2_inv_1 _15010_ (.Y(_05915_),
    .A(_05914_));
 sg13g2_nor2_1 _15011_ (.A(_05137_),
    .B(_05915_),
    .Y(_05916_));
 sg13g2_and3_1 _15012_ (.X(_05917_),
    .A(_05137_),
    .B(_05133_),
    .C(_05131_));
 sg13g2_inv_1 _15013_ (.Y(_05918_),
    .A(_05129_));
 sg13g2_nor2_1 _15014_ (.A(_05918_),
    .B(net70),
    .Y(_05919_));
 sg13g2_o21ai_1 _15015_ (.B1(_05919_),
    .Y(_05920_),
    .A1(_05916_),
    .A2(_05917_));
 sg13g2_nand3_1 _15016_ (.B(_05920_),
    .C(_05842_),
    .A(_05142_),
    .Y(_05921_));
 sg13g2_buf_1 _15017_ (.A(_05921_),
    .X(_05922_));
 sg13g2_o21ai_1 _15018_ (.B1(_05922_),
    .Y(_05923_),
    .A1(_05845_),
    .A2(_05913_));
 sg13g2_nor3_1 _15019_ (.A(_05549_),
    .B(_05550_),
    .C(_05548_),
    .Y(_05924_));
 sg13g2_nand2b_1 _15020_ (.Y(_05925_),
    .B(_05694_),
    .A_N(_05924_));
 sg13g2_nand2_1 _15021_ (.Y(_05926_),
    .A(_05557_),
    .B(_05925_));
 sg13g2_nand3_1 _15022_ (.B(_05566_),
    .C(_05926_),
    .A(_05560_),
    .Y(_05927_));
 sg13g2_inv_1 _15023_ (.Y(_05928_),
    .A(_05927_));
 sg13g2_a21oi_1 _15024_ (.A1(_05923_),
    .A2(net52),
    .Y(_05929_),
    .B1(_05928_));
 sg13g2_inv_1 _15025_ (.Y(_05930_),
    .A(_05929_));
 sg13g2_inv_1 _15026_ (.Y(_05931_),
    .A(_05449_));
 sg13g2_nand3_1 _15027_ (.B(_05931_),
    .C(_05446_),
    .A(_05457_),
    .Y(_05932_));
 sg13g2_a21oi_1 _15028_ (.A1(_05475_),
    .A2(_05932_),
    .Y(_05933_),
    .B1(net32));
 sg13g2_a21oi_2 _15029_ (.B1(_05466_),
    .Y(_05934_),
    .A2(_05453_),
    .A1(_05933_));
 sg13g2_a21oi_1 _15030_ (.A1(_05930_),
    .A2(_05934_),
    .Y(_05935_),
    .B1(_04732_));
 sg13g2_nand2b_1 _15031_ (.Y(_05936_),
    .B(_05935_),
    .A_N(_05839_));
 sg13g2_nand2b_1 _15032_ (.Y(_05937_),
    .B(_05936_),
    .A_N(_05838_));
 sg13g2_xnor2_1 _15033_ (.Y(_05938_),
    .A(_04589_),
    .B(_04735_));
 sg13g2_inv_1 _15034_ (.Y(_05939_),
    .A(_05573_));
 sg13g2_a21oi_1 _15035_ (.A1(_04746_),
    .A2(_04619_),
    .Y(_05940_),
    .B1(_04623_));
 sg13g2_buf_1 _15036_ (.A(_05940_),
    .X(_05941_));
 sg13g2_nand2_1 _15037_ (.Y(_05942_),
    .A(_05463_),
    .B(_04625_));
 sg13g2_nand2_1 _15038_ (.Y(_05943_),
    .A(_05942_),
    .B(_04628_));
 sg13g2_inv_1 _15039_ (.Y(_05944_),
    .A(_05943_));
 sg13g2_nor2_2 _15040_ (.A(_05941_),
    .B(_05944_),
    .Y(_05945_));
 sg13g2_inv_1 _15041_ (.Y(_05946_),
    .A(_05945_));
 sg13g2_nand4_1 _15042_ (.B(_05946_),
    .C(_05512_),
    .A(_05939_),
    .Y(_05947_),
    .D(_05471_));
 sg13g2_inv_1 _15043_ (.Y(_05948_),
    .A(_00047_));
 sg13g2_nor2_1 _15044_ (.A(_05948_),
    .B(net73),
    .Y(_05949_));
 sg13g2_buf_2 _15045_ (.A(_05949_),
    .X(_05950_));
 sg13g2_a21oi_1 _15046_ (.A1(_04176_),
    .A2(net73),
    .Y(_05951_),
    .B1(_05950_));
 sg13g2_inv_1 _15047_ (.Y(_05952_),
    .A(_05951_));
 sg13g2_buf_1 _15048_ (.A(_05863_),
    .X(_05953_));
 sg13g2_inv_1 _15049_ (.Y(_05954_),
    .A(_00053_));
 sg13g2_nor2_1 _15050_ (.A(_05954_),
    .B(_05863_),
    .Y(_05955_));
 sg13g2_buf_2 _15051_ (.A(_05955_),
    .X(_05956_));
 sg13g2_a21oi_1 _15052_ (.A1(_05952_),
    .A2(net22),
    .Y(_05957_),
    .B1(_05956_));
 sg13g2_inv_1 _15053_ (.Y(_05958_),
    .A(_05957_));
 sg13g2_a21oi_2 _15054_ (.B1(_04967_),
    .Y(_05959_),
    .A2(net42),
    .A1(_05958_));
 sg13g2_inv_1 _15055_ (.Y(_05960_),
    .A(_05959_));
 sg13g2_buf_2 _15056_ (.A(_05844_),
    .X(_05961_));
 sg13g2_nor2_1 _15057_ (.A(_05127_),
    .B(_05844_),
    .Y(_05962_));
 sg13g2_buf_2 _15058_ (.A(_05962_),
    .X(_05963_));
 sg13g2_a21oi_2 _15059_ (.B1(_05963_),
    .Y(_05964_),
    .A2(net28),
    .A1(_05960_));
 sg13g2_inv_1 _15060_ (.Y(_05965_),
    .A(_05964_));
 sg13g2_a21oi_1 _15061_ (.A1(_05965_),
    .A2(_05691_),
    .Y(_05966_),
    .B1(_05571_));
 sg13g2_nor2_1 _15062_ (.A(_05934_),
    .B(_05464_),
    .Y(_05967_));
 sg13g2_nor3_1 _15063_ (.A(_05828_),
    .B(_05967_),
    .C(_05833_),
    .Y(_05968_));
 sg13g2_o21ai_1 _15064_ (.B1(_05968_),
    .Y(_05969_),
    .A1(_05930_),
    .A2(_05966_));
 sg13g2_a21oi_1 _15065_ (.A1(_05738_),
    .A2(_04626_),
    .Y(_05970_),
    .B1(_04629_));
 sg13g2_a21oi_1 _15066_ (.A1(_05787_),
    .A2(net87),
    .Y(_05971_),
    .B1(_04754_));
 sg13g2_nand2b_1 _15067_ (.Y(_05972_),
    .B(_05971_),
    .A_N(_05970_));
 sg13g2_nand3_1 _15068_ (.B(_05253_),
    .C(_05254_),
    .A(_05425_),
    .Y(_05973_));
 sg13g2_nand2_1 _15069_ (.Y(_05974_),
    .A(_05973_),
    .B(_05257_));
 sg13g2_nand2_1 _15070_ (.Y(_05975_),
    .A(net147),
    .B(_05974_));
 sg13g2_nor2_1 _15071_ (.A(_05441_),
    .B(_05975_),
    .Y(_05976_));
 sg13g2_nor2_2 _15072_ (.A(_05976_),
    .B(_05269_),
    .Y(_05977_));
 sg13g2_nand2b_1 _15073_ (.Y(_05978_),
    .B(_05431_),
    .A_N(_05977_));
 sg13g2_buf_1 _15074_ (.A(\b.gen_square[8].sq.piece[2] ),
    .X(_05979_));
 sg13g2_inv_1 _15075_ (.Y(_05980_),
    .A(_05979_));
 sg13g2_buf_1 _15076_ (.A(\b.gen_square[8].sq.piece[1] ),
    .X(_05981_));
 sg13g2_buf_1 _15077_ (.A(\b.gen_square[8].sq.piece[0] ),
    .X(_05982_));
 sg13g2_nand2_1 _15078_ (.Y(_05983_),
    .A(_05981_),
    .B(_05982_));
 sg13g2_nor2_2 _15079_ (.A(_05980_),
    .B(_05983_),
    .Y(_05984_));
 sg13g2_inv_1 _15080_ (.Y(_05985_),
    .A(_05984_));
 sg13g2_inv_1 _15081_ (.Y(_05986_),
    .A(_05981_));
 sg13g2_nand3_1 _15082_ (.B(_05979_),
    .C(_05982_),
    .A(_05986_),
    .Y(_05987_));
 sg13g2_buf_1 _15083_ (.A(_05987_),
    .X(_05988_));
 sg13g2_xnor2_1 _15084_ (.Y(_05989_),
    .A(net166),
    .B(\b.gen_square[8].sq.color ));
 sg13g2_buf_8 _15085_ (.A(_05989_),
    .X(_05990_));
 sg13g2_nor2_1 _15086_ (.A(_05988_),
    .B(_05990_),
    .Y(_05991_));
 sg13g2_a22oi_1 _15087_ (.Y(_05992_),
    .B1(_04019_),
    .B2(_04089_),
    .A2(net118),
    .A1(_05991_));
 sg13g2_inv_2 _15088_ (.Y(_05993_),
    .A(_05992_));
 sg13g2_nor2_1 _15089_ (.A(_05985_),
    .B(_05993_),
    .Y(_05994_));
 sg13g2_buf_2 _15090_ (.A(_05994_),
    .X(_05995_));
 sg13g2_nor2_1 _15091_ (.A(_04836_),
    .B(_04840_),
    .Y(_05996_));
 sg13g2_nor2_1 _15092_ (.A(_04837_),
    .B(_04847_),
    .Y(_05997_));
 sg13g2_nor2_1 _15093_ (.A(_05996_),
    .B(_05997_),
    .Y(_05998_));
 sg13g2_inv_1 _15094_ (.Y(_05999_),
    .A(_05998_));
 sg13g2_a21oi_2 _15095_ (.B1(_04857_),
    .Y(_06000_),
    .A2(_04845_),
    .A1(_05999_));
 sg13g2_inv_1 _15096_ (.Y(_06001_),
    .A(_05990_));
 sg13g2_nor2_1 _15097_ (.A(_05979_),
    .B(_05983_),
    .Y(_06002_));
 sg13g2_nor2_1 _15098_ (.A(_05981_),
    .B(_05982_),
    .Y(_06003_));
 sg13g2_inv_1 _15099_ (.Y(_06004_),
    .A(_06003_));
 sg13g2_nor2_1 _15100_ (.A(_05980_),
    .B(_06004_),
    .Y(_06005_));
 sg13g2_nor2_1 _15101_ (.A(_06002_),
    .B(_06005_),
    .Y(_06006_));
 sg13g2_nor3_1 _15102_ (.A(_06001_),
    .B(net80),
    .C(_06006_),
    .Y(_06007_));
 sg13g2_nor2_2 _15103_ (.A(_06007_),
    .B(_05993_),
    .Y(_06008_));
 sg13g2_inv_1 _15104_ (.Y(_06009_),
    .A(_06008_));
 sg13g2_nor2_1 _15105_ (.A(_05984_),
    .B(_06009_),
    .Y(_06010_));
 sg13g2_a21oi_1 _15106_ (.A1(_05995_),
    .A2(_06000_),
    .Y(_06011_),
    .B1(_06010_));
 sg13g2_inv_1 _15107_ (.Y(_06012_),
    .A(_06011_));
 sg13g2_buf_2 _15108_ (.A(\b.gen_square[16].sq.piece[2] ),
    .X(_06013_));
 sg13g2_inv_1 _15109_ (.Y(_06014_),
    .A(_06013_));
 sg13g2_buf_1 _15110_ (.A(\b.gen_square[16].sq.piece[1] ),
    .X(_06015_));
 sg13g2_buf_2 _15111_ (.A(\b.gen_square[16].sq.piece[0] ),
    .X(_06016_));
 sg13g2_nand2_1 _15112_ (.Y(_06017_),
    .A(_06015_),
    .B(_06016_));
 sg13g2_nor2_1 _15113_ (.A(_06014_),
    .B(_06017_),
    .Y(_06018_));
 sg13g2_inv_1 _15114_ (.Y(_06019_),
    .A(_06018_));
 sg13g2_xnor2_1 _15115_ (.Y(_06020_),
    .A(_04076_),
    .B(\b.gen_square[16].sq.color ));
 sg13g2_buf_2 _15116_ (.A(_06020_),
    .X(_06021_));
 sg13g2_inv_8 _15117_ (.Y(_06022_),
    .A(_06021_));
 sg13g2_inv_1 _15118_ (.Y(_06023_),
    .A(_06016_));
 sg13g2_nor3_2 _15119_ (.A(_06015_),
    .B(_06014_),
    .C(_06023_),
    .Y(_06024_));
 sg13g2_nand2_1 _15120_ (.Y(_06025_),
    .A(_06022_),
    .B(_06024_));
 sg13g2_nand2_1 _15121_ (.Y(_06026_),
    .A(_03409_),
    .B(net134));
 sg13g2_o21ai_1 _15122_ (.B1(_06026_),
    .Y(_06027_),
    .A1(_04255_),
    .A2(_06025_));
 sg13g2_buf_2 _15123_ (.A(_06027_),
    .X(_06028_));
 sg13g2_nor2_1 _15124_ (.A(_06019_),
    .B(_06028_),
    .Y(_06029_));
 sg13g2_buf_2 _15125_ (.A(_06029_),
    .X(_06030_));
 sg13g2_nor2_1 _15126_ (.A(_06013_),
    .B(_06017_),
    .Y(_06031_));
 sg13g2_nor2_1 _15127_ (.A(_06015_),
    .B(_06016_),
    .Y(_06032_));
 sg13g2_inv_1 _15128_ (.Y(_06033_),
    .A(_06032_));
 sg13g2_nor2_1 _15129_ (.A(_06014_),
    .B(_06033_),
    .Y(_06034_));
 sg13g2_nor2_1 _15130_ (.A(_06031_),
    .B(_06034_),
    .Y(_06035_));
 sg13g2_nor3_1 _15131_ (.A(_06022_),
    .B(net80),
    .C(_06035_),
    .Y(_06036_));
 sg13g2_nor2_1 _15132_ (.A(_06036_),
    .B(_06028_),
    .Y(_06037_));
 sg13g2_inv_1 _15133_ (.Y(_06038_),
    .A(_06037_));
 sg13g2_nor2_1 _15134_ (.A(_06018_),
    .B(_06038_),
    .Y(_06039_));
 sg13g2_a21oi_1 _15135_ (.A1(_06012_),
    .A2(_06030_),
    .Y(_06040_),
    .B1(_06039_));
 sg13g2_inv_2 _15136_ (.Y(_06041_),
    .A(_06040_));
 sg13g2_inv_1 _15137_ (.Y(_06042_),
    .A(_03614_));
 sg13g2_inv_1 _15138_ (.Y(_06043_),
    .A(\b.gen_square[24].sq.piece[1] ));
 sg13g2_buf_1 _15139_ (.A(\b.gen_square[24].sq.piece[2] ),
    .X(_06044_));
 sg13g2_buf_2 _15140_ (.A(\b.gen_square[24].sq.piece[0] ),
    .X(_06045_));
 sg13g2_nand3_1 _15141_ (.B(_06044_),
    .C(_06045_),
    .A(_06043_),
    .Y(_06046_));
 sg13g2_buf_1 _15142_ (.A(_06046_),
    .X(_06047_));
 sg13g2_xnor2_1 _15143_ (.Y(_06048_),
    .A(net163),
    .B(\b.gen_square[24].sq.color ));
 sg13g2_buf_2 _15144_ (.A(_06048_),
    .X(_06049_));
 sg13g2_nor2_1 _15145_ (.A(_06047_),
    .B(_06049_),
    .Y(_06050_));
 sg13g2_nand2_1 _15146_ (.Y(_06051_),
    .A(_06050_),
    .B(net152));
 sg13g2_o21ai_1 _15147_ (.B1(_06051_),
    .Y(_06052_),
    .A1(net149),
    .A2(_06042_));
 sg13g2_buf_1 _15148_ (.A(_06052_),
    .X(_06053_));
 sg13g2_inv_1 _15149_ (.Y(_06054_),
    .A(_06044_));
 sg13g2_nand2_1 _15150_ (.Y(_06055_),
    .A(\b.gen_square[24].sq.piece[1] ),
    .B(_06045_));
 sg13g2_nor2_2 _15151_ (.A(_06054_),
    .B(_06055_),
    .Y(_06056_));
 sg13g2_nor2b_1 _15152_ (.A(_06053_),
    .B_N(_06056_),
    .Y(_06057_));
 sg13g2_buf_2 _15153_ (.A(_06057_),
    .X(_06058_));
 sg13g2_nor2_1 _15154_ (.A(\b.gen_square[24].sq.piece[1] ),
    .B(_06045_),
    .Y(_06059_));
 sg13g2_inv_1 _15155_ (.Y(_06060_),
    .A(_06059_));
 sg13g2_nor2_1 _15156_ (.A(_06054_),
    .B(_06060_),
    .Y(_06061_));
 sg13g2_inv_1 _15157_ (.Y(_06062_),
    .A(_06061_));
 sg13g2_nor2_1 _15158_ (.A(_06044_),
    .B(_06055_),
    .Y(_06063_));
 sg13g2_inv_1 _15159_ (.Y(_06064_),
    .A(_06063_));
 sg13g2_inv_2 _15160_ (.Y(_06065_),
    .A(_06049_));
 sg13g2_nor2_1 _15161_ (.A(_06065_),
    .B(net100),
    .Y(_06066_));
 sg13g2_inv_1 _15162_ (.Y(_06067_),
    .A(_06066_));
 sg13g2_a21oi_1 _15163_ (.A1(_06062_),
    .A2(_06064_),
    .Y(_06068_),
    .B1(_06067_));
 sg13g2_nor2_1 _15164_ (.A(_06053_),
    .B(_06068_),
    .Y(_06069_));
 sg13g2_inv_2 _15165_ (.Y(_06070_),
    .A(_06069_));
 sg13g2_nor2_1 _15166_ (.A(_06056_),
    .B(_06070_),
    .Y(_06071_));
 sg13g2_a21oi_1 _15167_ (.A1(_06041_),
    .A2(_06058_),
    .Y(_06072_),
    .B1(_06071_));
 sg13g2_inv_1 _15168_ (.Y(_06073_),
    .A(_06072_));
 sg13g2_nand2_1 _15169_ (.Y(_06074_),
    .A(_05151_),
    .B(_05152_));
 sg13g2_nor2_2 _15170_ (.A(_05157_),
    .B(_06074_),
    .Y(_06075_));
 sg13g2_inv_1 _15171_ (.Y(_06076_),
    .A(_06075_));
 sg13g2_nor2_2 _15172_ (.A(_06076_),
    .B(_05161_),
    .Y(_06077_));
 sg13g2_nor2_1 _15173_ (.A(_05151_),
    .B(_05152_),
    .Y(_06078_));
 sg13g2_inv_1 _15174_ (.Y(_06079_),
    .A(_06078_));
 sg13g2_nor2_1 _15175_ (.A(_05157_),
    .B(_06079_),
    .Y(_06080_));
 sg13g2_inv_1 _15176_ (.Y(_06081_),
    .A(_06080_));
 sg13g2_nor2_1 _15177_ (.A(_05150_),
    .B(_06074_),
    .Y(_06082_));
 sg13g2_inv_1 _15178_ (.Y(_06083_),
    .A(_06082_));
 sg13g2_inv_4 _15179_ (.A(_05149_),
    .Y(_06084_));
 sg13g2_nor2_1 _15180_ (.A(_06084_),
    .B(_04050_),
    .Y(_06085_));
 sg13g2_inv_1 _15181_ (.Y(_06086_),
    .A(_06085_));
 sg13g2_a21oi_1 _15182_ (.A1(_06081_),
    .A2(_06083_),
    .Y(_06087_),
    .B1(_06086_));
 sg13g2_nor2_1 _15183_ (.A(_06087_),
    .B(_05161_),
    .Y(_06088_));
 sg13g2_inv_2 _15184_ (.Y(_06089_),
    .A(_06088_));
 sg13g2_nor2_1 _15185_ (.A(_06075_),
    .B(_06089_),
    .Y(_06090_));
 sg13g2_a21oi_1 _15186_ (.A1(_06073_),
    .A2(_06077_),
    .Y(_06091_),
    .B1(_06090_));
 sg13g2_inv_1 _15187_ (.Y(_06092_),
    .A(_06091_));
 sg13g2_inv_2 _15188_ (.Y(_06093_),
    .A(_05497_));
 sg13g2_inv_1 _15189_ (.Y(_06094_),
    .A(_05495_));
 sg13g2_a21oi_1 _15190_ (.A1(_05235_),
    .A2(_06094_),
    .Y(_06095_),
    .B1(_05240_));
 sg13g2_nor3_1 _15191_ (.A(net119),
    .B(_05508_),
    .C(_06095_),
    .Y(_06096_));
 sg13g2_nor2_1 _15192_ (.A(_06096_),
    .B(_05250_),
    .Y(_06097_));
 sg13g2_inv_1 _15193_ (.Y(_06098_),
    .A(_05496_));
 sg13g2_nand2_1 _15194_ (.Y(_06099_),
    .A(_06097_),
    .B(_06098_));
 sg13g2_inv_1 _15195_ (.Y(_06100_),
    .A(_06099_));
 sg13g2_a21oi_1 _15196_ (.A1(_06092_),
    .A2(_06093_),
    .Y(_06101_),
    .B1(_06100_));
 sg13g2_inv_1 _15197_ (.Y(_06102_),
    .A(_00066_));
 sg13g2_nor2_1 _15198_ (.A(_06102_),
    .B(_05995_),
    .Y(_06103_));
 sg13g2_a21oi_1 _15199_ (.A1(_04953_),
    .A2(_05995_),
    .Y(_06104_),
    .B1(_06103_));
 sg13g2_inv_2 _15200_ (.Y(_06105_),
    .A(_06104_));
 sg13g2_inv_1 _15201_ (.Y(_06106_),
    .A(_00065_));
 sg13g2_nor2_1 _15202_ (.A(_06106_),
    .B(_06030_),
    .Y(_06107_));
 sg13g2_a21oi_2 _15203_ (.B1(_06107_),
    .Y(_06108_),
    .A2(_06030_),
    .A1(_06105_));
 sg13g2_inv_2 _15204_ (.Y(_06109_),
    .A(_06108_));
 sg13g2_inv_1 _15205_ (.Y(_06110_),
    .A(_00064_));
 sg13g2_nor2_1 _15206_ (.A(_06110_),
    .B(_06058_),
    .Y(_06111_));
 sg13g2_a21oi_2 _15207_ (.B1(_06111_),
    .Y(_06112_),
    .A2(_06058_),
    .A1(_06109_));
 sg13g2_nor2_1 _15208_ (.A(_00058_),
    .B(_06077_),
    .Y(_06113_));
 sg13g2_buf_2 _15209_ (.A(_06113_),
    .X(_06114_));
 sg13g2_a21oi_1 _15210_ (.A1(_06112_),
    .A2(_06077_),
    .Y(_06115_),
    .B1(_06114_));
 sg13g2_inv_1 _15211_ (.Y(_06116_),
    .A(_06115_));
 sg13g2_a21oi_2 _15212_ (.B1(_05501_),
    .Y(_06117_),
    .A2(_06093_),
    .A1(_06116_));
 sg13g2_nand2_1 _15213_ (.Y(_06118_),
    .A(_06101_),
    .B(_06117_));
 sg13g2_nand3_1 _15214_ (.B(_05978_),
    .C(_06118_),
    .A(_05972_),
    .Y(_06119_));
 sg13g2_nor3_1 _15215_ (.A(_05947_),
    .B(_05969_),
    .C(_06119_),
    .Y(_06120_));
 sg13g2_inv_1 _15216_ (.Y(_06121_),
    .A(_05562_));
 sg13g2_a21oi_1 _15217_ (.A1(_05966_),
    .A2(_06121_),
    .Y(_06122_),
    .B1(_05784_));
 sg13g2_nor2_1 _15218_ (.A(_05941_),
    .B(_05943_),
    .Y(_06123_));
 sg13g2_inv_1 _15219_ (.Y(_06124_),
    .A(_06123_));
 sg13g2_inv_1 _15220_ (.Y(_06125_),
    .A(_05779_));
 sg13g2_nand3_1 _15221_ (.B(_06124_),
    .C(_06125_),
    .A(_06122_),
    .Y(_06126_));
 sg13g2_nor2_1 _15222_ (.A(_05934_),
    .B(_05463_),
    .Y(_06127_));
 sg13g2_a21oi_1 _15223_ (.A1(_05966_),
    .A2(_05929_),
    .Y(_06128_),
    .B1(_06127_));
 sg13g2_nand2_1 _15224_ (.Y(_06129_),
    .A(_06128_),
    .B(_05826_));
 sg13g2_inv_1 _15225_ (.Y(_06130_),
    .A(_06101_));
 sg13g2_nor2_1 _15226_ (.A(_05977_),
    .B(_05431_),
    .Y(_06131_));
 sg13g2_a21oi_1 _15227_ (.A1(_05971_),
    .A2(_05970_),
    .Y(_06132_),
    .B1(_06131_));
 sg13g2_o21ai_1 _15228_ (.B1(_06132_),
    .Y(_06133_),
    .A1(_06117_),
    .A2(_06130_));
 sg13g2_nor3_1 _15229_ (.A(_06126_),
    .B(_06129_),
    .C(_06133_),
    .Y(_06134_));
 sg13g2_nor3_1 _15230_ (.A(_04600_),
    .B(_06120_),
    .C(_06134_),
    .Y(_06135_));
 sg13g2_nand2_1 _15231_ (.Y(_06136_),
    .A(_06135_),
    .B(net162));
 sg13g2_nand2_1 _15232_ (.Y(_06137_),
    .A(_06134_),
    .B(_06120_));
 sg13g2_nand3_1 _15233_ (.B(net113),
    .C(_04732_),
    .A(_06137_),
    .Y(_06138_));
 sg13g2_nand2_1 _15234_ (.Y(_06139_),
    .A(_06136_),
    .B(_06138_));
 sg13g2_a22oi_1 _15235_ (.Y(_06140_),
    .B1(_05938_),
    .B2(_06139_),
    .A2(_05937_),
    .A1(_05810_));
 sg13g2_o21ai_1 _15236_ (.B1(_04600_),
    .Y(_06141_),
    .A1(_06119_),
    .A2(_06133_));
 sg13g2_inv_1 _15237_ (.Y(_06142_),
    .A(_05935_));
 sg13g2_a21o_1 _15238_ (.A2(_06142_),
    .A1(_06141_),
    .B1(_04736_),
    .X(_06143_));
 sg13g2_o21ai_1 _15239_ (.B1(_06143_),
    .Y(_06144_),
    .A1(_04734_),
    .A2(_06141_));
 sg13g2_nand2_1 _15240_ (.Y(_06145_),
    .A(_06144_),
    .B(net95));
 sg13g2_nand2_1 _15241_ (.Y(_06146_),
    .A(_06140_),
    .B(_06145_));
 sg13g2_buf_1 _15242_ (.A(\b.gen_square[48].sq.mask ),
    .X(_06147_));
 sg13g2_nand2_1 _15243_ (.Y(_06148_),
    .A(_06146_),
    .B(_06147_));
 sg13g2_nand2_1 _15244_ (.Y(_06149_),
    .A(_05809_),
    .B(_06148_));
 sg13g2_nand2_1 _15245_ (.Y(_06150_),
    .A(_03260_),
    .B(_04065_));
 sg13g2_buf_1 _15246_ (.A(\b.gen_square[15].sq.piece[1] ),
    .X(_06151_));
 sg13g2_inv_1 _15247_ (.Y(_06152_),
    .A(_06151_));
 sg13g2_buf_2 _15248_ (.A(\b.gen_square[15].sq.piece[2] ),
    .X(_06153_));
 sg13g2_buf_2 _15249_ (.A(\b.gen_square[15].sq.piece[0] ),
    .X(_06154_));
 sg13g2_nand3_1 _15250_ (.B(_06153_),
    .C(_06154_),
    .A(_06152_),
    .Y(_06155_));
 sg13g2_buf_1 _15251_ (.A(_06155_),
    .X(_06156_));
 sg13g2_xnor2_1 _15252_ (.Y(_06157_),
    .A(_04039_),
    .B(_03221_));
 sg13g2_buf_8 _15253_ (.A(_06157_),
    .X(_06158_));
 sg13g2_nor2_1 _15254_ (.A(_06156_),
    .B(net159),
    .Y(_06159_));
 sg13g2_nand2_1 _15255_ (.Y(_06160_),
    .A(_06159_),
    .B(_04243_));
 sg13g2_inv_1 _15256_ (.Y(_06161_),
    .A(_06153_));
 sg13g2_nand2_1 _15257_ (.Y(_06162_),
    .A(_06151_),
    .B(_06154_));
 sg13g2_nor2_1 _15258_ (.A(_06161_),
    .B(_06162_),
    .Y(_06163_));
 sg13g2_nand3_1 _15259_ (.B(_06160_),
    .C(_06163_),
    .A(_06150_),
    .Y(_06164_));
 sg13g2_buf_8 _15260_ (.A(_06164_),
    .X(_06165_));
 sg13g2_inv_1 _15261_ (.Y(_06166_),
    .A(_00019_));
 sg13g2_nand2_2 _15262_ (.Y(_06167_),
    .A(_06165_),
    .B(_06166_));
 sg13g2_a21oi_2 _15263_ (.B1(_04220_),
    .Y(_06168_),
    .A2(_06167_),
    .A1(net62));
 sg13g2_inv_1 _15264_ (.Y(_06169_),
    .A(_06168_));
 sg13g2_buf_1 _15265_ (.A(\b.gen_square[29].sq.piece[1] ),
    .X(_06170_));
 sg13g2_inv_1 _15266_ (.Y(_06171_),
    .A(_06170_));
 sg13g2_buf_2 _15267_ (.A(\b.gen_square[29].sq.piece[2] ),
    .X(_06172_));
 sg13g2_buf_2 _15268_ (.A(\b.gen_square[29].sq.piece[0] ),
    .X(_06173_));
 sg13g2_nand3_1 _15269_ (.B(_06172_),
    .C(_06173_),
    .A(_06171_),
    .Y(_06174_));
 sg13g2_buf_1 _15270_ (.A(_06174_),
    .X(_06175_));
 sg13g2_xnor2_1 _15271_ (.Y(_06176_),
    .A(_04079_),
    .B(\b.gen_square[29].sq.color ));
 sg13g2_buf_2 _15272_ (.A(_06176_),
    .X(_06177_));
 sg13g2_nor2_1 _15273_ (.A(_06175_),
    .B(_06177_),
    .Y(_06178_));
 sg13g2_a22oi_1 _15274_ (.Y(_06179_),
    .B1(_04090_),
    .B2(_03659_),
    .A2(_04086_),
    .A1(_06178_));
 sg13g2_buf_2 _15275_ (.A(_06179_),
    .X(_06180_));
 sg13g2_inv_1 _15276_ (.Y(_06181_),
    .A(_06172_));
 sg13g2_nand2_1 _15277_ (.Y(_06182_),
    .A(_06170_),
    .B(_06173_));
 sg13g2_nor2_1 _15278_ (.A(_06181_),
    .B(_06182_),
    .Y(_06183_));
 sg13g2_nand2_2 _15279_ (.Y(_06184_),
    .A(_06180_),
    .B(_06183_));
 sg13g2_inv_4 _15280_ (.A(_06184_),
    .Y(_06185_));
 sg13g2_buf_1 _15281_ (.A(_06185_),
    .X(_06186_));
 sg13g2_inv_1 _15282_ (.Y(_06187_),
    .A(_00045_));
 sg13g2_nor2_1 _15283_ (.A(_06187_),
    .B(_06185_),
    .Y(_06188_));
 sg13g2_buf_8 _15284_ (.A(_06188_),
    .X(_06189_));
 sg13g2_a21oi_1 _15285_ (.A1(_06169_),
    .A2(net27),
    .Y(_06190_),
    .B1(_06189_));
 sg13g2_inv_1 _15286_ (.Y(_06191_),
    .A(_06190_));
 sg13g2_a21oi_1 _15287_ (.A1(_06191_),
    .A2(net58),
    .Y(_06192_),
    .B1(_04972_));
 sg13g2_inv_1 _15288_ (.Y(_06193_),
    .A(_06192_));
 sg13g2_nand2_1 _15289_ (.Y(_06194_),
    .A(_05169_),
    .B(_05170_));
 sg13g2_nor2_1 _15290_ (.A(_05175_),
    .B(_06194_),
    .Y(_06195_));
 sg13g2_inv_1 _15291_ (.Y(_06196_),
    .A(_06195_));
 sg13g2_nor2_1 _15292_ (.A(_06196_),
    .B(_05181_),
    .Y(_06197_));
 sg13g2_buf_2 _15293_ (.A(_06197_),
    .X(_06198_));
 sg13g2_buf_1 _15294_ (.A(_06198_),
    .X(_06199_));
 sg13g2_nor2_1 _15295_ (.A(_05165_),
    .B(_06198_),
    .Y(_06200_));
 sg13g2_buf_2 _15296_ (.A(_06200_),
    .X(_06201_));
 sg13g2_a21oi_1 _15297_ (.A1(_06193_),
    .A2(net21),
    .Y(_06202_),
    .B1(_06201_));
 sg13g2_inv_2 _15298_ (.Y(_06203_),
    .A(_04927_));
 sg13g2_inv_1 _15299_ (.Y(_06204_),
    .A(_06154_));
 sg13g2_nand3_1 _15300_ (.B(_06204_),
    .C(_06151_),
    .A(_06161_),
    .Y(_06205_));
 sg13g2_nor2_1 _15301_ (.A(_06151_),
    .B(_06154_),
    .Y(_06206_));
 sg13g2_nand2_1 _15302_ (.Y(_06207_),
    .A(_06206_),
    .B(_06153_));
 sg13g2_nand2_1 _15303_ (.Y(_06208_),
    .A(_06205_),
    .B(_06207_));
 sg13g2_nand2_1 _15304_ (.Y(_06209_),
    .A(_04263_),
    .B(net159));
 sg13g2_inv_1 _15305_ (.Y(_06210_),
    .A(_06209_));
 sg13g2_nand2_1 _15306_ (.Y(_06211_),
    .A(_06150_),
    .B(_06160_));
 sg13g2_a21oi_2 _15307_ (.B1(_06211_),
    .Y(_06212_),
    .A2(_06210_),
    .A1(_06208_));
 sg13g2_nor3_1 _15308_ (.A(_04200_),
    .B(_04203_),
    .C(_04207_),
    .Y(_06213_));
 sg13g2_nand2b_1 _15309_ (.Y(_06214_),
    .B(_04291_),
    .A_N(_06213_));
 sg13g2_nand2_1 _15310_ (.Y(_06215_),
    .A(_04288_),
    .B(_06214_));
 sg13g2_nand3_1 _15311_ (.B(_04206_),
    .C(_06215_),
    .A(_04283_),
    .Y(_06216_));
 sg13g2_inv_1 _15312_ (.Y(_06217_),
    .A(_06216_));
 sg13g2_a21oi_1 _15313_ (.A1(net47),
    .A2(_06212_),
    .Y(_06218_),
    .B1(_06217_));
 sg13g2_inv_1 _15314_ (.Y(_06219_),
    .A(_06218_));
 sg13g2_inv_1 _15315_ (.Y(_06220_),
    .A(_06183_));
 sg13g2_inv_1 _15316_ (.Y(_06221_),
    .A(_06177_));
 sg13g2_nor2_1 _15317_ (.A(_06221_),
    .B(_04287_),
    .Y(_06222_));
 sg13g2_nor3_1 _15318_ (.A(_06172_),
    .B(_06173_),
    .C(_06171_),
    .Y(_06223_));
 sg13g2_nor2_1 _15319_ (.A(_06170_),
    .B(_06173_),
    .Y(_06224_));
 sg13g2_nand2_1 _15320_ (.Y(_06225_),
    .A(_06224_),
    .B(_06172_));
 sg13g2_nand2b_1 _15321_ (.Y(_06226_),
    .B(_06225_),
    .A_N(_06223_));
 sg13g2_nand2_1 _15322_ (.Y(_06227_),
    .A(_06222_),
    .B(_06226_));
 sg13g2_nand3_1 _15323_ (.B(_06220_),
    .C(_06227_),
    .A(_06180_),
    .Y(_06228_));
 sg13g2_inv_1 _15324_ (.Y(_06229_),
    .A(_06228_));
 sg13g2_a21oi_2 _15325_ (.B1(_06229_),
    .Y(_06230_),
    .A2(net27),
    .A1(_06219_));
 sg13g2_o21ai_1 _15326_ (.B1(_04937_),
    .Y(_06231_),
    .A1(_06203_),
    .A2(_06230_));
 sg13g2_buf_1 _15327_ (.A(_06231_),
    .X(_06232_));
 sg13g2_and3_1 _15328_ (.X(_06233_),
    .A(_05175_),
    .B(_05171_),
    .C(_05169_));
 sg13g2_nor2_1 _15329_ (.A(_05169_),
    .B(_05170_),
    .Y(_06234_));
 sg13g2_nand2_1 _15330_ (.Y(_06235_),
    .A(_06234_),
    .B(_05168_));
 sg13g2_nand2b_1 _15331_ (.Y(_06236_),
    .B(_06235_),
    .A_N(_06233_));
 sg13g2_inv_1 _15332_ (.Y(_06237_),
    .A(net94));
 sg13g2_nor2_1 _15333_ (.A(_06237_),
    .B(net70),
    .Y(_06238_));
 sg13g2_nand2_1 _15334_ (.Y(_06239_),
    .A(_06236_),
    .B(_06238_));
 sg13g2_nand3_1 _15335_ (.B(_06196_),
    .C(_06239_),
    .A(_05180_),
    .Y(_06240_));
 sg13g2_inv_1 _15336_ (.Y(_06241_),
    .A(_06240_));
 sg13g2_a21oi_1 _15337_ (.A1(_06232_),
    .A2(net21),
    .Y(_06242_),
    .B1(_06241_));
 sg13g2_inv_1 _15338_ (.Y(_06243_),
    .A(_06242_));
 sg13g2_nor2_1 _15339_ (.A(_06202_),
    .B(_06243_),
    .Y(_06244_));
 sg13g2_nor2_1 _15340_ (.A(_05967_),
    .B(_06244_),
    .Y(_06245_));
 sg13g2_inv_1 _15341_ (.Y(_06246_),
    .A(_06245_));
 sg13g2_a21oi_2 _15342_ (.B1(_04672_),
    .Y(_06247_),
    .A2(_04667_),
    .A1(_04769_));
 sg13g2_a21oi_1 _15343_ (.A1(_05490_),
    .A2(net44),
    .Y(_06248_),
    .B1(_04678_));
 sg13g2_nor2_1 _15344_ (.A(_06247_),
    .B(_06248_),
    .Y(_06249_));
 sg13g2_buf_1 _15345_ (.A(_06249_),
    .X(_06250_));
 sg13g2_inv_1 _15346_ (.Y(_06251_),
    .A(_06250_));
 sg13g2_nand2_1 _15347_ (.Y(_06252_),
    .A(_05440_),
    .B(_06251_));
 sg13g2_nor2_1 _15348_ (.A(_04756_),
    .B(_04630_),
    .Y(_06253_));
 sg13g2_inv_1 _15349_ (.Y(_06254_),
    .A(_05187_));
 sg13g2_nor2_1 _15350_ (.A(_06254_),
    .B(net70),
    .Y(_06255_));
 sg13g2_a21oi_1 _15351_ (.A1(_05196_),
    .A2(_06255_),
    .Y(_06256_),
    .B1(_05199_));
 sg13g2_buf_1 _15352_ (.A(_06256_),
    .X(_06257_));
 sg13g2_nand2_1 _15353_ (.Y(_06258_),
    .A(_05189_),
    .B(_05190_));
 sg13g2_nor2_2 _15354_ (.A(_05195_),
    .B(_06258_),
    .Y(_06259_));
 sg13g2_inv_1 _15355_ (.Y(_06260_),
    .A(_06259_));
 sg13g2_nor2_1 _15356_ (.A(_06260_),
    .B(_05199_),
    .Y(_06261_));
 sg13g2_buf_2 _15357_ (.A(_06261_),
    .X(_06262_));
 sg13g2_nor2_2 _15358_ (.A(_03950_),
    .B(_06262_),
    .Y(_06263_));
 sg13g2_nor2_1 _15359_ (.A(_06257_),
    .B(_06263_),
    .Y(_06264_));
 sg13g2_nor2_1 _15360_ (.A(_05492_),
    .B(_06264_),
    .Y(_06265_));
 sg13g2_inv_1 _15361_ (.Y(_06266_),
    .A(_05470_));
 sg13g2_and3_1 _15362_ (.X(_06267_),
    .A(_05195_),
    .B(_05191_),
    .C(_05189_));
 sg13g2_inv_1 _15363_ (.Y(_06268_),
    .A(_06267_));
 sg13g2_nor2_1 _15364_ (.A(_05189_),
    .B(_05190_),
    .Y(_06269_));
 sg13g2_inv_1 _15365_ (.Y(_06270_),
    .A(_06269_));
 sg13g2_nor2_1 _15366_ (.A(_05195_),
    .B(_06270_),
    .Y(_06271_));
 sg13g2_inv_1 _15367_ (.Y(_06272_),
    .A(_06271_));
 sg13g2_a21oi_1 _15368_ (.A1(_06268_),
    .A2(_06272_),
    .Y(_06273_),
    .B1(net46));
 sg13g2_a21oi_2 _15369_ (.B1(_05199_),
    .Y(_06274_),
    .A2(_06273_),
    .A1(_05187_));
 sg13g2_nor2_1 _15370_ (.A(_06274_),
    .B(_06263_),
    .Y(_06275_));
 sg13g2_inv_1 _15371_ (.Y(_06276_),
    .A(_06275_));
 sg13g2_o21ai_1 _15372_ (.B1(_05219_),
    .Y(_06277_),
    .A1(_05218_),
    .A2(_05485_));
 sg13g2_nand2_1 _15373_ (.Y(_06278_),
    .A(_05483_),
    .B(_06277_));
 sg13g2_nand2_1 _15374_ (.Y(_06279_),
    .A(_05229_),
    .B(_06278_));
 sg13g2_nand2_1 _15375_ (.Y(_06280_),
    .A(_06279_),
    .B(_00025_));
 sg13g2_nand4_1 _15376_ (.B(_06266_),
    .C(_06276_),
    .A(_06265_),
    .Y(_06281_),
    .D(_06280_));
 sg13g2_nand4_1 _15377_ (.B(_05425_),
    .C(_05258_),
    .A(_05263_),
    .Y(_06282_),
    .D(_05254_));
 sg13g2_inv_1 _15378_ (.Y(_06283_),
    .A(_06282_));
 sg13g2_a21oi_1 _15379_ (.A1(_06283_),
    .A2(net78),
    .Y(_06284_),
    .B1(_05269_));
 sg13g2_nor2_1 _15380_ (.A(_05429_),
    .B(_06284_),
    .Y(_06285_));
 sg13g2_nand4_1 _15381_ (.B(_05235_),
    .C(_05245_),
    .A(_05233_),
    .Y(_06286_),
    .D(_05237_));
 sg13g2_inv_1 _15382_ (.Y(_06287_),
    .A(_06286_));
 sg13g2_a21oi_1 _15383_ (.A1(net99),
    .A2(_06287_),
    .Y(_06288_),
    .B1(_05250_));
 sg13g2_nor2_2 _15384_ (.A(_05498_),
    .B(_06288_),
    .Y(_06289_));
 sg13g2_nor2_1 _15385_ (.A(_06289_),
    .B(_04528_),
    .Y(_06290_));
 sg13g2_nor3_1 _15386_ (.A(_05360_),
    .B(_05362_),
    .C(_05369_),
    .Y(_06291_));
 sg13g2_nand2_1 _15387_ (.Y(_06292_),
    .A(_05368_),
    .B(_06291_));
 sg13g2_inv_1 _15388_ (.Y(_06293_),
    .A(_06292_));
 sg13g2_a21oi_1 _15389_ (.A1(net99),
    .A2(_06293_),
    .Y(_06294_),
    .B1(_05375_));
 sg13g2_nor2_1 _15390_ (.A(_05535_),
    .B(_06294_),
    .Y(_06295_));
 sg13g2_buf_2 _15391_ (.A(_06295_),
    .X(_06296_));
 sg13g2_inv_1 _15392_ (.Y(_06297_),
    .A(_06296_));
 sg13g2_nand3b_1 _15393_ (.B(_06290_),
    .C(_06297_),
    .Y(_06298_),
    .A_N(_04567_));
 sg13g2_nor3_1 _15394_ (.A(_05828_),
    .B(_06285_),
    .C(_06298_),
    .Y(_06299_));
 sg13g2_inv_2 _15395_ (.Y(_06300_),
    .A(_06114_));
 sg13g2_a21oi_1 _15396_ (.A1(_06300_),
    .A2(net52),
    .Y(_06301_),
    .B1(_05571_));
 sg13g2_inv_1 _15397_ (.Y(_06302_),
    .A(_06301_));
 sg13g2_and3_1 _15398_ (.X(_06303_),
    .A(_05157_),
    .B(_05153_),
    .C(_05151_));
 sg13g2_o21ai_1 _15399_ (.B1(net99),
    .Y(_06304_),
    .A1(_06080_),
    .A2(_06303_));
 sg13g2_o21ai_1 _15400_ (.B1(_05160_),
    .Y(_06305_),
    .A1(_06084_),
    .A2(_06304_));
 sg13g2_inv_1 _15401_ (.Y(_06306_),
    .A(_06305_));
 sg13g2_a21oi_1 _15402_ (.A1(_06306_),
    .A2(net52),
    .Y(_06307_),
    .B1(_05928_));
 sg13g2_nand2_1 _15403_ (.Y(_06308_),
    .A(_06302_),
    .B(_06307_));
 sg13g2_nand2_1 _15404_ (.Y(_06309_),
    .A(_06299_),
    .B(_06308_));
 sg13g2_nor3_1 _15405_ (.A(_06253_),
    .B(_06281_),
    .C(_06309_),
    .Y(_06310_));
 sg13g2_a21oi_2 _15406_ (.B1(_05181_),
    .Y(_06311_),
    .A2(_06238_),
    .A1(_05176_));
 sg13g2_a21oi_2 _15407_ (.B1(_06201_),
    .Y(_06312_),
    .A2(net21),
    .A1(_05767_));
 sg13g2_nor2_2 _15408_ (.A(_06311_),
    .B(_06312_),
    .Y(_06313_));
 sg13g2_inv_1 _15409_ (.Y(_06314_),
    .A(_06313_));
 sg13g2_nand4_1 _15410_ (.B(_05946_),
    .C(_06314_),
    .A(_06310_),
    .Y(_06315_),
    .D(_05939_));
 sg13g2_buf_2 _15411_ (.A(\b.gen_square[10].sq.piece[2] ),
    .X(_06316_));
 sg13g2_inv_2 _15412_ (.Y(_06317_),
    .A(_06316_));
 sg13g2_buf_1 _15413_ (.A(\b.gen_square[10].sq.piece[1] ),
    .X(_06318_));
 sg13g2_buf_2 _15414_ (.A(\b.gen_square[10].sq.piece[0] ),
    .X(_06319_));
 sg13g2_nand2_1 _15415_ (.Y(_06320_),
    .A(_06318_),
    .B(_06319_));
 sg13g2_nor2_1 _15416_ (.A(_06317_),
    .B(_06320_),
    .Y(_06321_));
 sg13g2_inv_1 _15417_ (.Y(_06322_),
    .A(_06321_));
 sg13g2_xnor2_1 _15418_ (.Y(_06323_),
    .A(net163),
    .B(\b.gen_square[10].sq.color ));
 sg13g2_buf_2 _15419_ (.A(_06323_),
    .X(_06324_));
 sg13g2_inv_2 _15420_ (.Y(_06325_),
    .A(_06319_));
 sg13g2_nor3_2 _15421_ (.A(_06318_),
    .B(_06317_),
    .C(_06325_),
    .Y(_06326_));
 sg13g2_inv_2 _15422_ (.Y(_06327_),
    .A(_06326_));
 sg13g2_nor2_1 _15423_ (.A(_06324_),
    .B(_06327_),
    .Y(_06328_));
 sg13g2_a22oi_1 _15424_ (.Y(_06329_),
    .B1(_04083_),
    .B2(_06328_),
    .A2(net117),
    .A1(_02481_));
 sg13g2_buf_1 _15425_ (.A(_06329_),
    .X(_06330_));
 sg13g2_inv_2 _15426_ (.Y(_06331_),
    .A(_06330_));
 sg13g2_nor2_1 _15427_ (.A(_06322_),
    .B(_06331_),
    .Y(_06332_));
 sg13g2_buf_8 _15428_ (.A(_06332_),
    .X(_06333_));
 sg13g2_buf_1 _15429_ (.A(_06333_),
    .X(_06334_));
 sg13g2_xnor2_1 _15430_ (.Y(_06335_),
    .A(net166),
    .B(_03668_));
 sg13g2_buf_1 _15431_ (.A(\b.gen_square[2].sq.piece[1] ),
    .X(_06336_));
 sg13g2_buf_2 _15432_ (.A(\b.gen_square[2].sq.piece[2] ),
    .X(_06337_));
 sg13g2_inv_2 _15433_ (.Y(_06338_),
    .A(_06337_));
 sg13g2_buf_2 _15434_ (.A(\b.gen_square[2].sq.piece[0] ),
    .X(_06339_));
 sg13g2_inv_1 _15435_ (.Y(_06340_),
    .A(_06339_));
 sg13g2_nor3_1 _15436_ (.A(_06336_),
    .B(_06338_),
    .C(_06340_),
    .Y(_06341_));
 sg13g2_inv_1 _15437_ (.Y(_06342_),
    .A(_06341_));
 sg13g2_nor2_1 _15438_ (.A(_06335_),
    .B(_06342_),
    .Y(_06343_));
 sg13g2_a22oi_1 _15439_ (.Y(_06344_),
    .B1(net118),
    .B2(_06343_),
    .A2(net117),
    .A1(_03670_));
 sg13g2_buf_1 _15440_ (.A(_06344_),
    .X(_06345_));
 sg13g2_nor2_1 _15441_ (.A(_06336_),
    .B(_06339_),
    .Y(_06346_));
 sg13g2_inv_1 _15442_ (.Y(_06347_),
    .A(_06346_));
 sg13g2_nor2_1 _15443_ (.A(_06338_),
    .B(_06347_),
    .Y(_06348_));
 sg13g2_nand2_1 _15444_ (.Y(_06349_),
    .A(_06336_),
    .B(_06339_));
 sg13g2_nor2_1 _15445_ (.A(_06337_),
    .B(_06349_),
    .Y(_06350_));
 sg13g2_inv_2 _15446_ (.Y(_06351_),
    .A(_06335_));
 sg13g2_nor2_1 _15447_ (.A(_06351_),
    .B(_04286_),
    .Y(_06352_));
 sg13g2_o21ai_1 _15448_ (.B1(_06352_),
    .Y(_06353_),
    .A1(_06348_),
    .A2(_06350_));
 sg13g2_nand2_1 _15449_ (.Y(_06354_),
    .A(_06345_),
    .B(_06353_));
 sg13g2_inv_1 _15450_ (.Y(_06355_),
    .A(_06354_));
 sg13g2_inv_2 _15451_ (.Y(_06356_),
    .A(_06324_));
 sg13g2_nor2_1 _15452_ (.A(_06356_),
    .B(net79),
    .Y(_06357_));
 sg13g2_nor2_1 _15453_ (.A(_06318_),
    .B(_06319_),
    .Y(_06358_));
 sg13g2_nand2_1 _15454_ (.Y(_06359_),
    .A(_06358_),
    .B(_06316_));
 sg13g2_o21ai_1 _15455_ (.B1(_06359_),
    .Y(_06360_),
    .A1(_06316_),
    .A2(_06320_));
 sg13g2_nand2_1 _15456_ (.Y(_06361_),
    .A(_06357_),
    .B(_06360_));
 sg13g2_nand3_1 _15457_ (.B(_06361_),
    .C(_06322_),
    .A(_06330_),
    .Y(_06362_));
 sg13g2_inv_1 _15458_ (.Y(_06363_),
    .A(_06362_));
 sg13g2_a21oi_1 _15459_ (.A1(_06334_),
    .A2(_06355_),
    .Y(_06364_),
    .B1(_06363_));
 sg13g2_inv_1 _15460_ (.Y(_06365_),
    .A(_06364_));
 sg13g2_nor2_1 _15461_ (.A(_04798_),
    .B(_04802_),
    .Y(_06366_));
 sg13g2_inv_1 _15462_ (.Y(_06367_),
    .A(_06366_));
 sg13g2_a21o_1 _15463_ (.A2(_06367_),
    .A1(_04870_),
    .B1(_04874_),
    .X(_06368_));
 sg13g2_nand3_1 _15464_ (.B(_04812_),
    .C(_04804_),
    .A(_06368_),
    .Y(_06369_));
 sg13g2_inv_1 _15465_ (.Y(_06370_),
    .A(_06369_));
 sg13g2_a21oi_2 _15466_ (.B1(_06370_),
    .Y(_06371_),
    .A2(net29),
    .A1(_06365_));
 sg13g2_inv_1 _15467_ (.Y(_06372_),
    .A(_06371_));
 sg13g2_buf_2 _15468_ (.A(\b.gen_square[26].sq.piece[2] ),
    .X(_06373_));
 sg13g2_inv_1 _15469_ (.Y(_06374_),
    .A(_06373_));
 sg13g2_buf_1 _15470_ (.A(\b.gen_square[26].sq.piece[1] ),
    .X(_06375_));
 sg13g2_buf_2 _15471_ (.A(\b.gen_square[26].sq.piece[0] ),
    .X(_06376_));
 sg13g2_nand2_1 _15472_ (.Y(_06377_),
    .A(_06375_),
    .B(_06376_));
 sg13g2_nor2_1 _15473_ (.A(_06374_),
    .B(_06377_),
    .Y(_06378_));
 sg13g2_inv_1 _15474_ (.Y(_06379_),
    .A(_06378_));
 sg13g2_xnor2_1 _15475_ (.Y(_06380_),
    .A(net166),
    .B(\b.gen_square[26].sq.color ));
 sg13g2_buf_1 _15476_ (.A(_06380_),
    .X(_06381_));
 sg13g2_inv_1 _15477_ (.Y(_06382_),
    .A(_06376_));
 sg13g2_nor3_2 _15478_ (.A(_06375_),
    .B(_06374_),
    .C(_06382_),
    .Y(_06383_));
 sg13g2_inv_1 _15479_ (.Y(_06384_),
    .A(_06383_));
 sg13g2_nor2_1 _15480_ (.A(net127),
    .B(_06384_),
    .Y(_06385_));
 sg13g2_nand2_1 _15481_ (.Y(_06386_),
    .A(_02459_),
    .B(net182));
 sg13g2_nor2_1 _15482_ (.A(net149),
    .B(_06386_),
    .Y(_06387_));
 sg13g2_a21oi_2 _15483_ (.B1(_06387_),
    .Y(_06388_),
    .A2(net118),
    .A1(_06385_));
 sg13g2_inv_2 _15484_ (.Y(_06389_),
    .A(_06388_));
 sg13g2_nor2_1 _15485_ (.A(_06379_),
    .B(_06389_),
    .Y(_06390_));
 sg13g2_buf_8 _15486_ (.A(_06390_),
    .X(_06391_));
 sg13g2_buf_1 _15487_ (.A(_06391_),
    .X(_06392_));
 sg13g2_nor2_1 _15488_ (.A(_06375_),
    .B(_06376_),
    .Y(_06393_));
 sg13g2_nand2_1 _15489_ (.Y(_06394_),
    .A(_06393_),
    .B(_06373_));
 sg13g2_nor2_1 _15490_ (.A(_06373_),
    .B(_06377_),
    .Y(_06395_));
 sg13g2_inv_1 _15491_ (.Y(_06396_),
    .A(_06395_));
 sg13g2_inv_1 _15492_ (.Y(_06397_),
    .A(net127));
 sg13g2_nor2_1 _15493_ (.A(_06397_),
    .B(net100),
    .Y(_06398_));
 sg13g2_inv_1 _15494_ (.Y(_06399_),
    .A(_06398_));
 sg13g2_a21oi_1 _15495_ (.A1(_06394_),
    .A2(_06396_),
    .Y(_06400_),
    .B1(_06399_));
 sg13g2_nand3b_1 _15496_ (.B(_06388_),
    .C(_06379_),
    .Y(_06401_),
    .A_N(_06400_));
 sg13g2_inv_1 _15497_ (.Y(_06402_),
    .A(_06401_));
 sg13g2_a21oi_1 _15498_ (.A1(_06372_),
    .A2(_06392_),
    .Y(_06403_),
    .B1(_06402_));
 sg13g2_inv_1 _15499_ (.Y(_06404_),
    .A(_06403_));
 sg13g2_nor2_1 _15500_ (.A(_05130_),
    .B(_05840_),
    .Y(_06405_));
 sg13g2_o21ai_1 _15501_ (.B1(_05919_),
    .Y(_06406_),
    .A1(_05916_),
    .A2(_06405_));
 sg13g2_nand3_1 _15502_ (.B(_06406_),
    .C(_05842_),
    .A(_05142_),
    .Y(_06407_));
 sg13g2_inv_1 _15503_ (.Y(_06408_),
    .A(_06407_));
 sg13g2_a21oi_2 _15504_ (.B1(_06408_),
    .Y(_06409_),
    .A2(net28),
    .A1(_06404_));
 sg13g2_nor2_1 _15505_ (.A(_05390_),
    .B(_05394_),
    .Y(_06410_));
 sg13g2_inv_1 _15506_ (.Y(_06411_),
    .A(_06410_));
 sg13g2_nand2_1 _15507_ (.Y(_06412_),
    .A(_06411_),
    .B(_05413_));
 sg13g2_nand2_1 _15508_ (.Y(_06413_),
    .A(_05410_),
    .B(_06412_));
 sg13g2_nand3_1 _15509_ (.B(_06413_),
    .C(_05396_),
    .A(_05404_),
    .Y(_06414_));
 sg13g2_o21ai_1 _15510_ (.B1(_06414_),
    .Y(_06415_),
    .A1(_05757_),
    .A2(_06409_));
 sg13g2_buf_1 _15511_ (.A(_06415_),
    .X(_06416_));
 sg13g2_nor2_1 _15512_ (.A(_06338_),
    .B(_06349_),
    .Y(_06417_));
 sg13g2_inv_1 _15513_ (.Y(_06418_),
    .A(_06417_));
 sg13g2_inv_2 _15514_ (.Y(_06419_),
    .A(_06345_));
 sg13g2_nor2_1 _15515_ (.A(_06418_),
    .B(_06419_),
    .Y(_06420_));
 sg13g2_buf_8 _15516_ (.A(_06420_),
    .X(_06421_));
 sg13g2_nor2_2 _15517_ (.A(_03669_),
    .B(_06421_),
    .Y(_06422_));
 sg13g2_inv_4 _15518_ (.A(_06422_),
    .Y(_06423_));
 sg13g2_inv_1 _15519_ (.Y(_06424_),
    .A(_00063_));
 sg13g2_nor2_1 _15520_ (.A(_06424_),
    .B(_06333_),
    .Y(_06425_));
 sg13g2_buf_1 _15521_ (.A(_06425_),
    .X(_06426_));
 sg13g2_a21oi_1 _15522_ (.A1(_06423_),
    .A2(net37),
    .Y(_06427_),
    .B1(_06426_));
 sg13g2_inv_1 _15523_ (.Y(_06428_),
    .A(_06427_));
 sg13g2_a21oi_1 _15524_ (.A1(_06428_),
    .A2(net29),
    .Y(_06429_),
    .B1(_04962_));
 sg13g2_inv_1 _15525_ (.Y(_06430_),
    .A(_06429_));
 sg13g2_inv_1 _15526_ (.Y(_06431_),
    .A(_00031_));
 sg13g2_nor2_1 _15527_ (.A(_06431_),
    .B(_06391_),
    .Y(_06432_));
 sg13g2_buf_2 _15528_ (.A(_06432_),
    .X(_06433_));
 sg13g2_a21oi_2 _15529_ (.B1(_06433_),
    .Y(_06434_),
    .A2(_06392_),
    .A1(_06430_));
 sg13g2_inv_1 _15530_ (.Y(_06435_),
    .A(_06434_));
 sg13g2_a21oi_1 _15531_ (.A1(_06435_),
    .A2(net28),
    .Y(_06436_),
    .B1(_05963_));
 sg13g2_inv_1 _15532_ (.Y(_06437_),
    .A(_06436_));
 sg13g2_a21oi_1 _15533_ (.A1(_06437_),
    .A2(net39),
    .Y(_06438_),
    .B1(_05436_));
 sg13g2_inv_1 _15534_ (.Y(_06439_),
    .A(_06438_));
 sg13g2_nand2b_1 _15535_ (.Y(_06440_),
    .B(_06439_),
    .A_N(_06416_));
 sg13g2_o21ai_1 _15536_ (.B1(_06440_),
    .Y(_06441_),
    .A1(_05735_),
    .A2(_05752_));
 sg13g2_nor4_1 _15537_ (.A(_06246_),
    .B(_06252_),
    .C(_06315_),
    .D(_06441_),
    .Y(_06442_));
 sg13g2_inv_1 _15538_ (.Y(_06443_),
    .A(_06442_));
 sg13g2_inv_4 _15539_ (.A(_06263_),
    .Y(_06444_));
 sg13g2_nor2_1 _15540_ (.A(_06274_),
    .B(_06444_),
    .Y(_06445_));
 sg13g2_inv_1 _15541_ (.Y(_06446_),
    .A(_06202_));
 sg13g2_a21oi_1 _15542_ (.A1(_06301_),
    .A2(_06307_),
    .Y(_06447_),
    .B1(_06127_));
 sg13g2_o21ai_1 _15543_ (.B1(_06447_),
    .Y(_06448_),
    .A1(_06243_),
    .A2(_06446_));
 sg13g2_nor2_1 _15544_ (.A(_06445_),
    .B(_06448_),
    .Y(_06449_));
 sg13g2_nor2_1 _15545_ (.A(_05782_),
    .B(_05765_),
    .Y(_06450_));
 sg13g2_nand2_1 _15546_ (.Y(_06451_),
    .A(_06449_),
    .B(_06450_));
 sg13g2_inv_1 _15547_ (.Y(_06452_),
    .A(_06248_));
 sg13g2_nor2_1 _15548_ (.A(_06247_),
    .B(_06452_),
    .Y(_06453_));
 sg13g2_buf_1 _15549_ (.A(_06453_),
    .X(_06454_));
 sg13g2_nor2_1 _15550_ (.A(_06257_),
    .B(_06444_),
    .Y(_06455_));
 sg13g2_nor4_1 _15551_ (.A(_06454_),
    .B(_06123_),
    .C(_06455_),
    .D(_05763_),
    .Y(_06456_));
 sg13g2_inv_1 _15552_ (.Y(_06457_),
    .A(_06456_));
 sg13g2_nor2_1 _15553_ (.A(_06416_),
    .B(_06439_),
    .Y(_06458_));
 sg13g2_a21oi_1 _15554_ (.A1(_04630_),
    .A2(_04755_),
    .Y(_06459_),
    .B1(_06458_));
 sg13g2_a22oi_1 _15555_ (.Y(_06460_),
    .B1(_05735_),
    .B2(_05751_),
    .A2(_06279_),
    .A1(_05488_));
 sg13g2_nor2_2 _15556_ (.A(_03721_),
    .B(_06294_),
    .Y(_06461_));
 sg13g2_nand2b_1 _15557_ (.Y(_06462_),
    .B(\b.gen_square[56].sq.color ),
    .A_N(_06284_));
 sg13g2_o21ai_1 _15558_ (.B1(_06462_),
    .Y(_06463_),
    .A1(_03968_),
    .A2(_04566_));
 sg13g2_nor2_1 _15559_ (.A(_03778_),
    .B(_06288_),
    .Y(_06464_));
 sg13g2_nor2_1 _15560_ (.A(_06464_),
    .B(_05015_),
    .Y(_06465_));
 sg13g2_inv_1 _15561_ (.Y(_06466_),
    .A(_06465_));
 sg13g2_nor4_2 _15562_ (.A(_05815_),
    .B(_06461_),
    .C(_06463_),
    .Y(_06467_),
    .D(_06466_));
 sg13g2_inv_1 _15563_ (.Y(_06468_),
    .A(_06312_));
 sg13g2_nor2_1 _15564_ (.A(_06311_),
    .B(_06468_),
    .Y(_06469_));
 sg13g2_buf_2 _15565_ (.A(_06469_),
    .X(_06470_));
 sg13g2_a21oi_1 _15566_ (.A1(_06301_),
    .A2(_06121_),
    .Y(_06471_),
    .B1(_06470_));
 sg13g2_nand4_1 _15567_ (.B(_06460_),
    .C(_06467_),
    .A(_06459_),
    .Y(_06472_),
    .D(_06471_));
 sg13g2_nor3_1 _15568_ (.A(_06451_),
    .B(_06457_),
    .C(_06472_),
    .Y(_06473_));
 sg13g2_inv_1 _15569_ (.Y(_06474_),
    .A(_06473_));
 sg13g2_nor2_1 _15570_ (.A(_06443_),
    .B(_06474_),
    .Y(_06475_));
 sg13g2_inv_1 _15571_ (.Y(_06476_),
    .A(_06475_));
 sg13g2_nand3_1 _15572_ (.B(net86),
    .C(_04757_),
    .A(_06476_),
    .Y(_06477_));
 sg13g2_nand4_1 _15573_ (.B(net145),
    .C(_04757_),
    .A(_06474_),
    .Y(_06478_),
    .D(_06443_));
 sg13g2_buf_1 _15574_ (.A(_06478_),
    .X(_06479_));
 sg13g2_nand2_1 _15575_ (.Y(_06480_),
    .A(_06477_),
    .B(_06479_));
 sg13g2_xnor2_1 _15576_ (.Y(_06481_),
    .A(_04632_),
    .B(_04760_));
 sg13g2_nand3b_1 _15577_ (.B(_06274_),
    .C(_06308_),
    .Y(_06482_),
    .A_N(_06448_));
 sg13g2_o21ai_1 _15578_ (.B1(_04644_),
    .Y(_06483_),
    .A1(_06246_),
    .A2(_06482_));
 sg13g2_nor3_1 _15579_ (.A(_04632_),
    .B(_04635_),
    .C(_04639_),
    .Y(_06484_));
 sg13g2_nand2b_1 _15580_ (.Y(_06485_),
    .B(_06484_),
    .A_N(_06483_));
 sg13g2_inv_1 _15581_ (.Y(_06486_),
    .A(_04635_));
 sg13g2_nor3_1 _15582_ (.A(_04632_),
    .B(_04634_),
    .C(_06486_),
    .Y(_06487_));
 sg13g2_nand2_1 _15583_ (.Y(_06488_),
    .A(_04644_),
    .B(_06487_));
 sg13g2_a21o_1 _15584_ (.A2(_06467_),
    .A1(_06299_),
    .B1(_06488_),
    .X(_06489_));
 sg13g2_nand2_1 _15585_ (.Y(_06490_),
    .A(_04641_),
    .B(net85));
 sg13g2_a21oi_1 _15586_ (.A1(_06485_),
    .A2(_06489_),
    .Y(_06491_),
    .B1(_06490_));
 sg13g2_a21oi_1 _15587_ (.A1(_06480_),
    .A2(_06481_),
    .Y(_06492_),
    .B1(_06491_));
 sg13g2_nand2_1 _15588_ (.Y(_06493_),
    .A(_06460_),
    .B(_06280_));
 sg13g2_nor4_1 _15589_ (.A(_04755_),
    .B(_06458_),
    .C(_06493_),
    .D(_06441_),
    .Y(_06494_));
 sg13g2_nand2b_1 _15590_ (.Y(_06495_),
    .B(_04644_),
    .A_N(_06494_));
 sg13g2_a21o_1 _15591_ (.A2(_06483_),
    .A1(_06495_),
    .B1(_04761_),
    .X(_06496_));
 sg13g2_nand2b_1 _15592_ (.Y(_06497_),
    .B(_04759_),
    .A_N(_06495_));
 sg13g2_a21o_1 _15593_ (.A2(_06497_),
    .A1(_06496_),
    .B1(_06490_),
    .X(_06498_));
 sg13g2_inv_1 _15594_ (.Y(_06499_),
    .A(\b.gen_square[50].sq.mask ));
 sg13g2_a21o_1 _15595_ (.A2(_06498_),
    .A1(_06492_),
    .B1(_06499_),
    .X(_06500_));
 sg13g2_buf_1 _15596_ (.A(_06500_),
    .X(_06501_));
 sg13g2_nor2b_1 _15597_ (.A(_06149_),
    .B_N(_06501_),
    .Y(_06502_));
 sg13g2_nor2_1 _15598_ (.A(_05734_),
    .B(_05750_),
    .Y(_06503_));
 sg13g2_inv_1 _15599_ (.Y(_06504_),
    .A(_06503_));
 sg13g2_nand2_1 _15600_ (.Y(_06505_),
    .A(_05734_),
    .B(_05749_));
 sg13g2_nor2_1 _15601_ (.A(_05188_),
    .B(_06258_),
    .Y(_06506_));
 sg13g2_nor2_1 _15602_ (.A(_06506_),
    .B(_06271_),
    .Y(_06507_));
 sg13g2_inv_1 _15603_ (.Y(_06508_),
    .A(_06255_));
 sg13g2_nor2_1 _15604_ (.A(_06507_),
    .B(_06508_),
    .Y(_06509_));
 sg13g2_nor2_1 _15605_ (.A(_06509_),
    .B(_05199_),
    .Y(_06510_));
 sg13g2_nand4_1 _15606_ (.B(_06505_),
    .C(_06510_),
    .A(_06504_),
    .Y(_06511_),
    .D(_04767_));
 sg13g2_inv_1 _15607_ (.Y(_06512_),
    .A(_05377_));
 sg13g2_buf_1 _15608_ (.A(\b.gen_square[11].sq.piece[2] ),
    .X(_06513_));
 sg13g2_inv_2 _15609_ (.Y(_06514_),
    .A(_06513_));
 sg13g2_buf_1 _15610_ (.A(\b.gen_square[11].sq.piece[1] ),
    .X(_06515_));
 sg13g2_buf_2 _15611_ (.A(\b.gen_square[11].sq.piece[0] ),
    .X(_06516_));
 sg13g2_nand2_1 _15612_ (.Y(_06517_),
    .A(_06515_),
    .B(_06516_));
 sg13g2_nor2_1 _15613_ (.A(_06514_),
    .B(_06517_),
    .Y(_06518_));
 sg13g2_inv_1 _15614_ (.Y(_06519_),
    .A(_06518_));
 sg13g2_xnor2_1 _15615_ (.Y(_06520_),
    .A(_04077_),
    .B(\b.gen_square[11].sq.color ));
 sg13g2_buf_2 _15616_ (.A(_06520_),
    .X(_06521_));
 sg13g2_inv_2 _15617_ (.Y(_06522_),
    .A(_06516_));
 sg13g2_nor3_2 _15618_ (.A(_06515_),
    .B(_06514_),
    .C(_06522_),
    .Y(_06523_));
 sg13g2_nor2b_1 _15619_ (.A(_06521_),
    .B_N(_06523_),
    .Y(_06524_));
 sg13g2_a22oi_1 _15620_ (.Y(_06525_),
    .B1(_04084_),
    .B2(_06524_),
    .A2(_04088_),
    .A1(_02642_));
 sg13g2_buf_1 _15621_ (.A(_06525_),
    .X(_06526_));
 sg13g2_inv_1 _15622_ (.Y(_06527_),
    .A(_06526_));
 sg13g2_nor2_1 _15623_ (.A(_06519_),
    .B(_06527_),
    .Y(_06528_));
 sg13g2_buf_2 _15624_ (.A(_06528_),
    .X(_06529_));
 sg13g2_buf_1 _15625_ (.A(_06529_),
    .X(_06530_));
 sg13g2_buf_1 _15626_ (.A(\b.gen_square[3].sq.piece[2] ),
    .X(_06531_));
 sg13g2_inv_1 _15627_ (.Y(_06532_),
    .A(_06531_));
 sg13g2_buf_2 _15628_ (.A(\b.gen_square[3].sq.piece[0] ),
    .X(_06533_));
 sg13g2_nor2_1 _15629_ (.A(\b.gen_square[3].sq.piece[1] ),
    .B(_06533_),
    .Y(_06534_));
 sg13g2_inv_1 _15630_ (.Y(_06535_),
    .A(_06534_));
 sg13g2_nor2_1 _15631_ (.A(_06532_),
    .B(_06535_),
    .Y(_06536_));
 sg13g2_nand2_1 _15632_ (.Y(_06537_),
    .A(\b.gen_square[3].sq.piece[1] ),
    .B(_06533_));
 sg13g2_nor2_1 _15633_ (.A(_06531_),
    .B(_06537_),
    .Y(_06538_));
 sg13g2_xnor2_1 _15634_ (.Y(_06539_),
    .A(_04642_),
    .B(\b.gen_square[3].sq.color ));
 sg13g2_buf_1 _15635_ (.A(_06539_),
    .X(_06540_));
 sg13g2_inv_2 _15636_ (.Y(_06541_),
    .A(_06540_));
 sg13g2_nor2_1 _15637_ (.A(_06541_),
    .B(_04285_),
    .Y(_06542_));
 sg13g2_o21ai_1 _15638_ (.B1(_06542_),
    .Y(_06543_),
    .A1(_06536_),
    .A2(_06538_));
 sg13g2_inv_1 _15639_ (.Y(_06544_),
    .A(\b.gen_square[3].sq.piece[1] ));
 sg13g2_nand3_1 _15640_ (.B(_06531_),
    .C(_06533_),
    .A(_06544_),
    .Y(_06545_));
 sg13g2_buf_1 _15641_ (.A(_06545_),
    .X(_06546_));
 sg13g2_nor2_1 _15642_ (.A(_06546_),
    .B(_06540_),
    .Y(_06547_));
 sg13g2_a22oi_1 _15643_ (.Y(_06548_),
    .B1(_03770_),
    .B2(_04088_),
    .A2(_04083_),
    .A1(_06547_));
 sg13g2_buf_2 _15644_ (.A(_06548_),
    .X(_06549_));
 sg13g2_nand2_1 _15645_ (.Y(_06550_),
    .A(_06543_),
    .B(_06549_));
 sg13g2_inv_1 _15646_ (.Y(_06551_),
    .A(_06550_));
 sg13g2_nor2_1 _15647_ (.A(_06515_),
    .B(_06516_),
    .Y(_06552_));
 sg13g2_inv_1 _15648_ (.Y(_06553_),
    .A(_06552_));
 sg13g2_nor2_2 _15649_ (.A(_06514_),
    .B(_06553_),
    .Y(_06554_));
 sg13g2_nor2_1 _15650_ (.A(_06513_),
    .B(_06517_),
    .Y(_06555_));
 sg13g2_inv_1 _15651_ (.Y(_06556_),
    .A(_06521_));
 sg13g2_nor2_1 _15652_ (.A(_06556_),
    .B(net79),
    .Y(_06557_));
 sg13g2_o21ai_1 _15653_ (.B1(_06557_),
    .Y(_06558_),
    .A1(_06554_),
    .A2(_06555_));
 sg13g2_nand3_1 _15654_ (.B(_06519_),
    .C(_06558_),
    .A(_06526_),
    .Y(_06559_));
 sg13g2_inv_1 _15655_ (.Y(_06560_),
    .A(_06559_));
 sg13g2_a21oi_1 _15656_ (.A1(net36),
    .A2(_06551_),
    .Y(_06561_),
    .B1(_06560_));
 sg13g2_inv_1 _15657_ (.Y(_06562_),
    .A(_06561_));
 sg13g2_buf_1 _15658_ (.A(\b.gen_square[19].sq.piece[1] ),
    .X(_06563_));
 sg13g2_buf_2 _15659_ (.A(\b.gen_square[19].sq.piece[0] ),
    .X(_06564_));
 sg13g2_nand2_1 _15660_ (.Y(_06565_),
    .A(_06563_),
    .B(_06564_));
 sg13g2_buf_2 _15661_ (.A(\b.gen_square[19].sq.piece[2] ),
    .X(_06566_));
 sg13g2_nor2b_1 _15662_ (.A(_06565_),
    .B_N(_06566_),
    .Y(_06567_));
 sg13g2_inv_1 _15663_ (.Y(_06568_),
    .A(_06567_));
 sg13g2_inv_1 _15664_ (.Y(_06569_),
    .A(_06563_));
 sg13g2_nand3_1 _15665_ (.B(_06566_),
    .C(_06564_),
    .A(_06569_),
    .Y(_06570_));
 sg13g2_buf_1 _15666_ (.A(_06570_),
    .X(_06571_));
 sg13g2_xnor2_1 _15667_ (.Y(_06572_),
    .A(_04077_),
    .B(\b.gen_square[19].sq.color ));
 sg13g2_buf_8 _15668_ (.A(_06572_),
    .X(_06573_));
 sg13g2_nor2_1 _15669_ (.A(_06571_),
    .B(net126),
    .Y(_06574_));
 sg13g2_a22oi_1 _15670_ (.Y(_06575_),
    .B1(_03550_),
    .B2(_04089_),
    .A2(_04084_),
    .A1(_06574_));
 sg13g2_buf_1 _15671_ (.A(_06575_),
    .X(_06576_));
 sg13g2_inv_1 _15672_ (.Y(_06577_),
    .A(_06576_));
 sg13g2_nor2_1 _15673_ (.A(_06568_),
    .B(_06577_),
    .Y(_06578_));
 sg13g2_buf_1 _15674_ (.A(_06578_),
    .X(_06579_));
 sg13g2_buf_1 _15675_ (.A(net35),
    .X(_06580_));
 sg13g2_inv_1 _15676_ (.Y(_06581_),
    .A(net126));
 sg13g2_nor2_1 _15677_ (.A(_06581_),
    .B(_04287_),
    .Y(_06582_));
 sg13g2_nor2_1 _15678_ (.A(_06566_),
    .B(_06565_),
    .Y(_06583_));
 sg13g2_nor2_1 _15679_ (.A(_06563_),
    .B(_06564_),
    .Y(_06584_));
 sg13g2_nand2_1 _15680_ (.Y(_06585_),
    .A(_06584_),
    .B(_06566_));
 sg13g2_nand2b_1 _15681_ (.Y(_06586_),
    .B(_06585_),
    .A_N(_06583_));
 sg13g2_nand2_1 _15682_ (.Y(_06587_),
    .A(_06582_),
    .B(_06586_));
 sg13g2_nand3_1 _15683_ (.B(_06568_),
    .C(_06587_),
    .A(_06576_),
    .Y(_06588_));
 sg13g2_inv_1 _15684_ (.Y(_06589_),
    .A(_06588_));
 sg13g2_a21oi_1 _15685_ (.A1(_06562_),
    .A2(net26),
    .Y(_06590_),
    .B1(_06589_));
 sg13g2_inv_1 _15686_ (.Y(_06591_),
    .A(_06590_));
 sg13g2_o21ai_1 _15687_ (.B1(_04901_),
    .Y(_06592_),
    .A1(_04879_),
    .A2(_04883_));
 sg13g2_nand2_1 _15688_ (.Y(_06593_),
    .A(_04904_),
    .B(_06592_));
 sg13g2_nand3_1 _15689_ (.B(_04885_),
    .C(_06593_),
    .A(_04894_),
    .Y(_06594_));
 sg13g2_buf_1 _15690_ (.A(_06594_),
    .X(_06595_));
 sg13g2_inv_1 _15691_ (.Y(_06596_),
    .A(_06595_));
 sg13g2_a21oi_2 _15692_ (.B1(_06596_),
    .Y(_06597_),
    .A2(net42),
    .A1(_06591_));
 sg13g2_nor2_1 _15693_ (.A(_05360_),
    .B(_05364_),
    .Y(_06598_));
 sg13g2_inv_1 _15694_ (.Y(_06599_),
    .A(_06598_));
 sg13g2_nand2_1 _15695_ (.Y(_06600_),
    .A(_06599_),
    .B(_05383_));
 sg13g2_nand2_1 _15696_ (.Y(_06601_),
    .A(_05380_),
    .B(_06600_));
 sg13g2_nand3_1 _15697_ (.B(_05366_),
    .C(_06601_),
    .A(_05374_),
    .Y(_06602_));
 sg13g2_buf_1 _15698_ (.A(_06602_),
    .X(_06603_));
 sg13g2_o21ai_1 _15699_ (.B1(_06603_),
    .Y(_06604_),
    .A1(_06512_),
    .A2(_06597_));
 sg13g2_buf_1 _15700_ (.A(_06604_),
    .X(_06605_));
 sg13g2_nor2_1 _15701_ (.A(_05168_),
    .B(_06194_),
    .Y(_06606_));
 sg13g2_inv_1 _15702_ (.Y(_06607_),
    .A(_06606_));
 sg13g2_nand2_1 _15703_ (.Y(_06608_),
    .A(_06607_),
    .B(_06235_));
 sg13g2_nand2_1 _15704_ (.Y(_06609_),
    .A(_06238_),
    .B(_06608_));
 sg13g2_nand3_1 _15705_ (.B(_06196_),
    .C(_06609_),
    .A(_05180_),
    .Y(_06610_));
 sg13g2_inv_1 _15706_ (.Y(_06611_),
    .A(_06610_));
 sg13g2_a21oi_1 _15707_ (.A1(_06605_),
    .A2(_06199_),
    .Y(_06612_),
    .B1(_06611_));
 sg13g2_o21ai_1 _15708_ (.B1(_04665_),
    .Y(_06613_),
    .A1(_06511_),
    .A2(_06612_));
 sg13g2_nor2b_1 _15709_ (.A(_06613_),
    .B_N(_04770_),
    .Y(_06614_));
 sg13g2_inv_1 _15710_ (.Y(_06615_),
    .A(_05550_));
 sg13g2_nor3_1 _15711_ (.A(_05549_),
    .B(_05547_),
    .C(_06615_),
    .Y(_06616_));
 sg13g2_nand2_1 _15712_ (.Y(_06617_),
    .A(net190),
    .B(_06616_));
 sg13g2_inv_1 _15713_ (.Y(_06618_),
    .A(_06617_));
 sg13g2_a21oi_1 _15714_ (.A1(net88),
    .A2(_06618_),
    .Y(_06619_),
    .B1(_05561_));
 sg13g2_nor2_2 _15715_ (.A(_05569_),
    .B(_06619_),
    .Y(_06620_));
 sg13g2_nand3_1 _15716_ (.B(_04054_),
    .C(_04056_),
    .A(_04123_),
    .Y(_06621_));
 sg13g2_nor2_1 _15717_ (.A(_06621_),
    .B(_04042_),
    .Y(_06622_));
 sg13g2_a21oi_1 _15718_ (.A1(net69),
    .A2(_06622_),
    .Y(_06623_),
    .B1(_04068_));
 sg13g2_nor2b_1 _15719_ (.A(_06623_),
    .B_N(_00072_),
    .Y(_06624_));
 sg13g2_buf_2 _15720_ (.A(_06624_),
    .X(_06625_));
 sg13g2_nand4_1 _15721_ (.B(_05457_),
    .C(_05447_),
    .A(_05453_),
    .Y(_06626_),
    .D(_05449_));
 sg13g2_o21ai_1 _15722_ (.B1(_05467_),
    .Y(_06627_),
    .A1(net46),
    .A2(_06626_));
 sg13g2_inv_1 _15723_ (.Y(_06628_),
    .A(_06627_));
 sg13g2_nor2_1 _15724_ (.A(_05461_),
    .B(_06628_),
    .Y(_06629_));
 sg13g2_inv_1 _15725_ (.Y(_06630_),
    .A(_00022_));
 sg13g2_nor3_1 _15726_ (.A(_04364_),
    .B(_04363_),
    .C(_04367_),
    .Y(_06631_));
 sg13g2_nand2_1 _15727_ (.Y(_06632_),
    .A(_04361_),
    .B(_06631_));
 sg13g2_inv_1 _15728_ (.Y(_06633_),
    .A(_06632_));
 sg13g2_a21oi_1 _15729_ (.A1(net60),
    .A2(_06633_),
    .Y(_06634_),
    .B1(_04374_));
 sg13g2_nor2_1 _15730_ (.A(_06630_),
    .B(_06634_),
    .Y(_06635_));
 sg13g2_nor3_1 _15731_ (.A(_04910_),
    .B(_04912_),
    .C(_04919_),
    .Y(_06636_));
 sg13g2_nand2_1 _15732_ (.Y(_06637_),
    .A(net146),
    .B(_06636_));
 sg13g2_inv_1 _15733_ (.Y(_06638_),
    .A(_06637_));
 sg13g2_a21oi_1 _15734_ (.A1(net88),
    .A2(_06638_),
    .Y(_06639_),
    .B1(_04925_));
 sg13g2_nor2_1 _15735_ (.A(_04970_),
    .B(_06639_),
    .Y(_06640_));
 sg13g2_buf_2 _15736_ (.A(_06640_),
    .X(_06641_));
 sg13g2_nor2_1 _15737_ (.A(_05146_),
    .B(_06641_),
    .Y(_06642_));
 sg13g2_nand2b_1 _15738_ (.Y(_06643_),
    .B(_06642_),
    .A_N(_06635_));
 sg13g2_nor4_1 _15739_ (.A(_06620_),
    .B(_06625_),
    .C(_06629_),
    .D(_06643_),
    .Y(_06644_));
 sg13g2_nor2_1 _15740_ (.A(_03976_),
    .B(_06634_),
    .Y(_06645_));
 sg13g2_nor2_2 _15741_ (.A(_03729_),
    .B(_06639_),
    .Y(_06646_));
 sg13g2_nor2_1 _15742_ (.A(_06645_),
    .B(_06646_),
    .Y(_06647_));
 sg13g2_nor2_1 _15743_ (.A(_03934_),
    .B(_06628_),
    .Y(_06648_));
 sg13g2_nor2_1 _15744_ (.A(_06648_),
    .B(_05205_),
    .Y(_06649_));
 sg13g2_nor2_2 _15745_ (.A(_03820_),
    .B(_06623_),
    .Y(_06650_));
 sg13g2_nor2_2 _15746_ (.A(_03786_),
    .B(_06619_),
    .Y(_06651_));
 sg13g2_nor2_1 _15747_ (.A(_06650_),
    .B(_06651_),
    .Y(_06652_));
 sg13g2_nand3_1 _15748_ (.B(_06649_),
    .C(_06652_),
    .A(_06647_),
    .Y(_06653_));
 sg13g2_inv_1 _15749_ (.Y(_06654_),
    .A(_06653_));
 sg13g2_nor3_1 _15750_ (.A(_04657_),
    .B(_04659_),
    .C(_04666_),
    .Y(_06655_));
 sg13g2_nand2_1 _15751_ (.Y(_06656_),
    .A(_04665_),
    .B(_06655_));
 sg13g2_a21oi_1 _15752_ (.A1(_06644_),
    .A2(_06654_),
    .Y(_06657_),
    .B1(_06656_));
 sg13g2_nand3_1 _15753_ (.B(_04666_),
    .C(_04659_),
    .A(_04658_),
    .Y(_06658_));
 sg13g2_nand2_1 _15754_ (.Y(_06659_),
    .A(\b.gen_square[44].sq.piece[1] ),
    .B(_04517_));
 sg13g2_nor2_1 _15755_ (.A(_04515_),
    .B(_06659_),
    .Y(_06660_));
 sg13g2_nand2_1 _15756_ (.Y(_06661_),
    .A(_04524_),
    .B(_06660_));
 sg13g2_buf_2 _15757_ (.A(_06661_),
    .X(_06662_));
 sg13g2_xnor2_1 _15758_ (.Y(_06663_),
    .A(_04078_),
    .B(\b.gen_square[23].sq.color ));
 sg13g2_buf_2 _15759_ (.A(_06663_),
    .X(_06664_));
 sg13g2_buf_1 _15760_ (.A(\b.gen_square[23].sq.piece[1] ),
    .X(_06665_));
 sg13g2_buf_1 _15761_ (.A(\b.gen_square[23].sq.piece[0] ),
    .X(_06666_));
 sg13g2_nor2_1 _15762_ (.A(_06665_),
    .B(_06666_),
    .Y(_06667_));
 sg13g2_buf_1 _15763_ (.A(\b.gen_square[23].sq.piece[2] ),
    .X(_06668_));
 sg13g2_nand2_1 _15764_ (.Y(_06669_),
    .A(_06667_),
    .B(_06668_));
 sg13g2_inv_1 _15765_ (.Y(_06670_),
    .A(_06666_));
 sg13g2_inv_1 _15766_ (.Y(_06671_),
    .A(_06668_));
 sg13g2_nand3_1 _15767_ (.B(_06671_),
    .C(_06665_),
    .A(_06670_),
    .Y(_06672_));
 sg13g2_a21oi_1 _15768_ (.A1(_06669_),
    .A2(_06672_),
    .Y(_06673_),
    .B1(_04348_));
 sg13g2_nand2_1 _15769_ (.Y(_06674_),
    .A(_03604_),
    .B(net182));
 sg13g2_nor2_1 _15770_ (.A(_04141_),
    .B(_06674_),
    .Y(_06675_));
 sg13g2_nand3b_1 _15771_ (.B(_06666_),
    .C(_06668_),
    .Y(_06676_),
    .A_N(_06665_));
 sg13g2_buf_1 _15772_ (.A(_06676_),
    .X(_06677_));
 sg13g2_nor2_1 _15773_ (.A(_06664_),
    .B(_06677_),
    .Y(_06678_));
 sg13g2_nand2_1 _15774_ (.Y(_06679_),
    .A(_06678_),
    .B(_04085_));
 sg13g2_nand2b_1 _15775_ (.Y(_06680_),
    .B(_06679_),
    .A_N(_06675_));
 sg13g2_buf_1 _15776_ (.A(_06680_),
    .X(_06681_));
 sg13g2_a21oi_1 _15777_ (.A1(_06664_),
    .A2(_06673_),
    .Y(_06682_),
    .B1(_06681_));
 sg13g2_buf_1 _15778_ (.A(_06682_),
    .X(_06683_));
 sg13g2_nor3_1 _15779_ (.A(_04135_),
    .B(_04137_),
    .C(_04144_),
    .Y(_06684_));
 sg13g2_nand2b_1 _15780_ (.Y(_06685_),
    .B(_04305_),
    .A_N(_06684_));
 sg13g2_nand2_1 _15781_ (.Y(_06686_),
    .A(_04301_),
    .B(_06685_));
 sg13g2_nand3_1 _15782_ (.B(_06686_),
    .C(_04140_),
    .A(_04298_),
    .Y(_06687_));
 sg13g2_inv_1 _15783_ (.Y(_06688_),
    .A(_06687_));
 sg13g2_a21oi_1 _15784_ (.A1(_06683_),
    .A2(net33),
    .Y(_06689_),
    .B1(_06688_));
 sg13g2_inv_1 _15785_ (.Y(_06690_),
    .A(_06689_));
 sg13g2_inv_1 _15786_ (.Y(_06691_),
    .A(_04533_));
 sg13g2_nand2_1 _15787_ (.Y(_06692_),
    .A(_04534_),
    .B(_04535_));
 sg13g2_nor2_1 _15788_ (.A(_06691_),
    .B(_06692_),
    .Y(_06693_));
 sg13g2_inv_1 _15789_ (.Y(_06694_),
    .A(_06693_));
 sg13g2_nor2_1 _15790_ (.A(_06694_),
    .B(_04546_),
    .Y(_06695_));
 sg13g2_buf_2 _15791_ (.A(_06695_),
    .X(_06696_));
 sg13g2_buf_1 _15792_ (.A(_06696_),
    .X(_06697_));
 sg13g2_inv_1 _15793_ (.Y(_06698_),
    .A(net164));
 sg13g2_nor2_1 _15794_ (.A(_06698_),
    .B(net100),
    .Y(_06699_));
 sg13g2_nor3_1 _15795_ (.A(_04533_),
    .B(_04535_),
    .C(_04540_),
    .Y(_06700_));
 sg13g2_nor2_1 _15796_ (.A(_04534_),
    .B(_04535_),
    .Y(_06701_));
 sg13g2_nand2_1 _15797_ (.Y(_06702_),
    .A(_06701_),
    .B(_04533_));
 sg13g2_nand2b_1 _15798_ (.Y(_06703_),
    .B(_06702_),
    .A_N(_06700_));
 sg13g2_nand2_1 _15799_ (.Y(_06704_),
    .A(_06699_),
    .B(_06703_));
 sg13g2_nand3_1 _15800_ (.B(_06704_),
    .C(_06694_),
    .A(_04545_),
    .Y(_06705_));
 sg13g2_buf_1 _15801_ (.A(_06705_),
    .X(_06706_));
 sg13g2_inv_1 _15802_ (.Y(_06707_),
    .A(_06706_));
 sg13g2_a21oi_2 _15803_ (.B1(_06707_),
    .Y(_06708_),
    .A2(net50),
    .A1(_06690_));
 sg13g2_nor2_1 _15804_ (.A(\b.gen_square[44].sq.piece[1] ),
    .B(_04517_),
    .Y(_06709_));
 sg13g2_inv_1 _15805_ (.Y(_06710_),
    .A(_06709_));
 sg13g2_nor2_1 _15806_ (.A(_04515_),
    .B(_06710_),
    .Y(_06711_));
 sg13g2_nor3_1 _15807_ (.A(_04514_),
    .B(_04517_),
    .C(_04516_),
    .Y(_06712_));
 sg13g2_inv_1 _15808_ (.Y(_06713_),
    .A(_04513_));
 sg13g2_nor2_1 _15809_ (.A(_06713_),
    .B(net119),
    .Y(_06714_));
 sg13g2_o21ai_1 _15810_ (.B1(_06714_),
    .Y(_06715_),
    .A1(_06711_),
    .A2(_06712_));
 sg13g2_inv_1 _15811_ (.Y(_06716_),
    .A(_06660_));
 sg13g2_nand3_1 _15812_ (.B(_04524_),
    .C(_06716_),
    .A(_06715_),
    .Y(_06717_));
 sg13g2_buf_1 _15813_ (.A(_06717_),
    .X(_06718_));
 sg13g2_o21ai_1 _15814_ (.B1(_06718_),
    .Y(_06719_),
    .A1(_06662_),
    .A2(_06708_));
 sg13g2_inv_1 _15815_ (.Y(_06720_),
    .A(_06719_));
 sg13g2_nand2_1 _15816_ (.Y(_06721_),
    .A(_06665_),
    .B(_06666_));
 sg13g2_nor2_2 _15817_ (.A(_06671_),
    .B(_06721_),
    .Y(_06722_));
 sg13g2_nand3b_1 _15818_ (.B(_06679_),
    .C(_06722_),
    .Y(_06723_),
    .A_N(_06675_));
 sg13g2_buf_1 _15819_ (.A(_06723_),
    .X(_06724_));
 sg13g2_inv_1 _15820_ (.Y(_06725_),
    .A(_00018_));
 sg13g2_nand2_1 _15821_ (.Y(_06726_),
    .A(_06724_),
    .B(_06725_));
 sg13g2_buf_2 _15822_ (.A(_06726_),
    .X(_06727_));
 sg13g2_a21oi_2 _15823_ (.B1(_04224_),
    .Y(_06728_),
    .A2(net33),
    .A1(_06727_));
 sg13g2_inv_1 _15824_ (.Y(_06729_),
    .A(_06728_));
 sg13g2_nor2_1 _15825_ (.A(_04529_),
    .B(_06696_),
    .Y(_06730_));
 sg13g2_buf_2 _15826_ (.A(_06730_),
    .X(_06731_));
 sg13g2_a21oi_2 _15827_ (.B1(_06731_),
    .Y(_06732_),
    .A2(_06697_),
    .A1(_06729_));
 sg13g2_inv_1 _15828_ (.Y(_06733_),
    .A(_06732_));
 sg13g2_inv_4 _15829_ (.A(_06662_),
    .Y(_06734_));
 sg13g2_buf_1 _15830_ (.A(_06734_),
    .X(_06735_));
 sg13g2_nor2_1 _15831_ (.A(_04507_),
    .B(_06734_),
    .Y(_06736_));
 sg13g2_buf_8 _15832_ (.A(_06736_),
    .X(_06737_));
 sg13g2_a21oi_1 _15833_ (.A1(_06733_),
    .A2(net66),
    .Y(_06738_),
    .B1(_06737_));
 sg13g2_nand2_1 _15834_ (.Y(_06739_),
    .A(_06720_),
    .B(_06738_));
 sg13g2_inv_1 _15835_ (.Y(_06740_),
    .A(_05777_));
 sg13g2_nor2_1 _15836_ (.A(_03611_),
    .B(_06058_),
    .Y(_06741_));
 sg13g2_buf_8 _15837_ (.A(_06741_),
    .X(_06742_));
 sg13g2_inv_1 _15838_ (.Y(_06743_),
    .A(_06742_));
 sg13g2_a21oi_2 _15839_ (.B1(_05723_),
    .Y(_06744_),
    .A2(net74),
    .A1(_06743_));
 sg13g2_inv_1 _15840_ (.Y(_06745_),
    .A(_06744_));
 sg13g2_a21oi_1 _15841_ (.A1(_06745_),
    .A2(net39),
    .Y(_06746_),
    .B1(_05436_));
 sg13g2_nor3_1 _15842_ (.A(_06044_),
    .B(_06045_),
    .C(_06043_),
    .Y(_06747_));
 sg13g2_inv_1 _15843_ (.Y(_06748_),
    .A(_06747_));
 sg13g2_a21oi_1 _15844_ (.A1(_06062_),
    .A2(_06748_),
    .Y(_06749_),
    .B1(_04347_));
 sg13g2_a21oi_2 _15845_ (.B1(_06053_),
    .Y(_06750_),
    .A2(_06749_),
    .A1(_06049_));
 sg13g2_and3_1 _15846_ (.X(_06751_),
    .A(_05661_),
    .B(_05669_),
    .C(_05662_));
 sg13g2_nand2b_1 _15847_ (.Y(_06752_),
    .B(_05683_),
    .A_N(_06751_));
 sg13g2_nand2_1 _15848_ (.Y(_06753_),
    .A(_06752_),
    .B(_05680_));
 sg13g2_nand3_1 _15849_ (.B(_05666_),
    .C(_06753_),
    .A(_05674_),
    .Y(_06754_));
 sg13g2_inv_1 _15850_ (.Y(_06755_),
    .A(_06754_));
 sg13g2_a21oi_1 _15851_ (.A1(_06750_),
    .A2(_05678_),
    .Y(_06756_),
    .B1(_06755_));
 sg13g2_inv_1 _15852_ (.Y(_06757_),
    .A(_06756_));
 sg13g2_a21oi_1 _15853_ (.A1(_06757_),
    .A2(net39),
    .Y(_06758_),
    .B1(_05417_));
 sg13g2_nand2_1 _15854_ (.Y(_06759_),
    .A(_06746_),
    .B(_06758_));
 sg13g2_nor2_1 _15855_ (.A(_04554_),
    .B(_04555_),
    .Y(_06760_));
 sg13g2_inv_1 _15856_ (.Y(_06761_),
    .A(_06760_));
 sg13g2_nor2_1 _15857_ (.A(_04560_),
    .B(_06761_),
    .Y(_06762_));
 sg13g2_inv_1 _15858_ (.Y(_06763_),
    .A(_06762_));
 sg13g2_nand3_1 _15859_ (.B(_04556_),
    .C(_04554_),
    .A(_04560_),
    .Y(_06764_));
 sg13g2_a21oi_1 _15860_ (.A1(_06763_),
    .A2(_06764_),
    .Y(_06765_),
    .B1(net61));
 sg13g2_a21oi_2 _15861_ (.B1(_04565_),
    .Y(_06766_),
    .A2(_06765_),
    .A1(_04552_));
 sg13g2_nor2_1 _15862_ (.A(_06766_),
    .B(_04997_),
    .Y(_06767_));
 sg13g2_inv_1 _15863_ (.Y(_06768_),
    .A(_06767_));
 sg13g2_nand4_1 _15864_ (.B(_06740_),
    .C(_06759_),
    .A(_06739_),
    .Y(_06769_),
    .D(_06768_));
 sg13g2_inv_1 _15865_ (.Y(_06770_),
    .A(_06738_));
 sg13g2_a21oi_1 _15866_ (.A1(_06770_),
    .A2(_06720_),
    .Y(_06771_),
    .B1(_05493_));
 sg13g2_inv_1 _15867_ (.Y(_06772_),
    .A(_06758_));
 sg13g2_nor2_1 _15868_ (.A(_06772_),
    .B(_06746_),
    .Y(_06773_));
 sg13g2_inv_1 _15869_ (.Y(_06774_),
    .A(_06773_));
 sg13g2_nor2_1 _15870_ (.A(_06766_),
    .B(_04996_),
    .Y(_06775_));
 sg13g2_inv_1 _15871_ (.Y(_06776_),
    .A(_06775_));
 sg13g2_nand3_1 _15872_ (.B(_06774_),
    .C(_06776_),
    .A(_06771_),
    .Y(_06777_));
 sg13g2_o21ai_1 _15873_ (.B1(_04665_),
    .Y(_06778_),
    .A1(_06769_),
    .A2(_06777_));
 sg13g2_nor2_1 _15874_ (.A(_06658_),
    .B(_06778_),
    .Y(_06779_));
 sg13g2_a21oi_1 _15875_ (.A1(_06613_),
    .A2(_06778_),
    .Y(_06780_),
    .B1(_04772_));
 sg13g2_nor4_1 _15876_ (.A(_06614_),
    .B(_06657_),
    .C(_06779_),
    .D(_06780_),
    .Y(_06781_));
 sg13g2_nor2_1 _15877_ (.A(_04767_),
    .B(_04655_),
    .Y(_06782_));
 sg13g2_inv_1 _15878_ (.Y(_06783_),
    .A(_06510_));
 sg13g2_inv_1 _15879_ (.Y(_06784_),
    .A(_04552_));
 sg13g2_nor2_1 _15880_ (.A(_06784_),
    .B(net61),
    .Y(_06785_));
 sg13g2_a21oi_1 _15881_ (.A1(_04561_),
    .A2(_06785_),
    .Y(_06786_),
    .B1(_04565_));
 sg13g2_buf_1 _15882_ (.A(_06786_),
    .X(_06787_));
 sg13g2_inv_1 _15883_ (.Y(_06788_),
    .A(_06787_));
 sg13g2_a221oi_1 _15884_ (.B2(_06788_),
    .C1(_06775_),
    .B1(_04997_),
    .A1(_03950_),
    .Y(_06789_),
    .A2(_06783_));
 sg13g2_nand4_1 _15885_ (.B(_06774_),
    .C(_06265_),
    .A(_06644_),
    .Y(_06790_),
    .D(_06789_));
 sg13g2_nor4_1 _15886_ (.A(_05546_),
    .B(_05439_),
    .C(_06782_),
    .D(_06790_),
    .Y(_06791_));
 sg13g2_inv_1 _15887_ (.Y(_06792_),
    .A(_04521_));
 sg13g2_a21oi_2 _15888_ (.B1(_04525_),
    .Y(_06793_),
    .A2(_06792_),
    .A1(_06714_));
 sg13g2_a21oi_2 _15889_ (.B1(_06737_),
    .Y(_06794_),
    .A2(net66),
    .A1(_06452_));
 sg13g2_nor2_2 _15890_ (.A(_06793_),
    .B(_06794_),
    .Y(_06795_));
 sg13g2_inv_1 _15891_ (.Y(_06796_),
    .A(_06795_));
 sg13g2_nand4_1 _15892_ (.B(_06796_),
    .C(_06771_),
    .A(_06791_),
    .Y(_06797_),
    .D(_06505_));
 sg13g2_inv_1 _15893_ (.Y(_06798_),
    .A(\b.gen_square[3].sq.color ));
 sg13g2_nor2_1 _15894_ (.A(_06532_),
    .B(_06537_),
    .Y(_06799_));
 sg13g2_inv_1 _15895_ (.Y(_06800_),
    .A(_06799_));
 sg13g2_inv_2 _15896_ (.Y(_06801_),
    .A(_06549_));
 sg13g2_nor2_1 _15897_ (.A(_06800_),
    .B(_06801_),
    .Y(_06802_));
 sg13g2_buf_2 _15898_ (.A(_06802_),
    .X(_06803_));
 sg13g2_nor2_2 _15899_ (.A(_06798_),
    .B(_06803_),
    .Y(_06804_));
 sg13g2_inv_4 _15900_ (.A(_06804_),
    .Y(_06805_));
 sg13g2_inv_1 _15901_ (.Y(_06806_),
    .A(_00060_));
 sg13g2_nor2_1 _15902_ (.A(_06806_),
    .B(_06529_),
    .Y(_06807_));
 sg13g2_buf_2 _15903_ (.A(_06807_),
    .X(_06808_));
 sg13g2_a21oi_2 _15904_ (.B1(_06808_),
    .Y(_06809_),
    .A2(net36),
    .A1(_06805_));
 sg13g2_inv_2 _15905_ (.Y(_06810_),
    .A(_06809_));
 sg13g2_nor2b_1 _15906_ (.A(net35),
    .B_N(_00059_),
    .Y(_06811_));
 sg13g2_buf_2 _15907_ (.A(_06811_),
    .X(_06812_));
 sg13g2_a21oi_1 _15908_ (.A1(_06810_),
    .A2(net35),
    .Y(_06813_),
    .B1(_06812_));
 sg13g2_inv_1 _15909_ (.Y(_06814_),
    .A(_06813_));
 sg13g2_a21oi_1 _15910_ (.A1(_06814_),
    .A2(net42),
    .Y(_06815_),
    .B1(_04967_));
 sg13g2_inv_1 _15911_ (.Y(_06816_),
    .A(_06815_));
 sg13g2_a21oi_2 _15912_ (.B1(_05537_),
    .Y(_06817_),
    .A2(net54),
    .A1(_06816_));
 sg13g2_inv_1 _15913_ (.Y(_06818_),
    .A(_06817_));
 sg13g2_a21oi_1 _15914_ (.A1(_06818_),
    .A2(net21),
    .Y(_06819_),
    .B1(_06201_));
 sg13g2_inv_1 _15915_ (.Y(_06820_),
    .A(_06819_));
 sg13g2_nand2_1 _15916_ (.Y(_06821_),
    .A(_06820_),
    .B(_06612_));
 sg13g2_a21oi_2 _15917_ (.B1(_04696_),
    .Y(_06822_),
    .A2(_04780_),
    .A1(_04691_));
 sg13g2_a21oi_1 _15918_ (.A1(_04997_),
    .A2(net30),
    .Y(_06823_),
    .B1(_04702_));
 sg13g2_nor2_1 _15919_ (.A(_06822_),
    .B(_06823_),
    .Y(_06824_));
 sg13g2_buf_2 _15920_ (.A(_06824_),
    .X(_06825_));
 sg13g2_nor2_1 _15921_ (.A(_06825_),
    .B(_06313_),
    .Y(_06826_));
 sg13g2_nand3b_1 _15922_ (.B(_06821_),
    .C(_06826_),
    .Y(_06827_),
    .A_N(_06797_));
 sg13g2_inv_1 _15923_ (.Y(_06828_),
    .A(_06823_));
 sg13g2_nor2_1 _15924_ (.A(_06822_),
    .B(_06828_),
    .Y(_06829_));
 sg13g2_buf_2 _15925_ (.A(_06829_),
    .X(_06830_));
 sg13g2_nor2_1 _15926_ (.A(_06787_),
    .B(_04997_),
    .Y(_06831_));
 sg13g2_nor4_1 _15927_ (.A(_05768_),
    .B(_06830_),
    .C(_06831_),
    .D(_06470_),
    .Y(_06832_));
 sg13g2_inv_1 _15928_ (.Y(_06833_),
    .A(_06832_));
 sg13g2_nor2_1 _15929_ (.A(_05765_),
    .B(_06455_),
    .Y(_06834_));
 sg13g2_inv_1 _15930_ (.Y(_06835_),
    .A(_06793_));
 sg13g2_a221oi_1 _15931_ (.B2(_06835_),
    .C1(_05763_),
    .B1(_06794_),
    .A1(_06783_),
    .Y(_06836_),
    .A2(_06263_));
 sg13g2_nand4_1 _15932_ (.B(_06654_),
    .C(_06834_),
    .A(_06504_),
    .Y(_06837_),
    .D(_06836_));
 sg13g2_inv_1 _15933_ (.Y(_06838_),
    .A(_06612_));
 sg13g2_nand2_1 _15934_ (.Y(_06839_),
    .A(_04655_),
    .B(_04766_));
 sg13g2_o21ai_1 _15935_ (.B1(_06839_),
    .Y(_06840_),
    .A1(_06838_),
    .A2(_06820_));
 sg13g2_nor4_1 _15936_ (.A(_06769_),
    .B(_06833_),
    .C(_06837_),
    .D(_06840_),
    .Y(_06841_));
 sg13g2_inv_1 _15937_ (.Y(_06842_),
    .A(_06841_));
 sg13g2_nor2_1 _15938_ (.A(_06827_),
    .B(_06842_),
    .Y(_06843_));
 sg13g2_inv_1 _15939_ (.Y(_06844_),
    .A(_06843_));
 sg13g2_nand3_1 _15940_ (.B(net68),
    .C(_04768_),
    .A(_06844_),
    .Y(_06845_));
 sg13g2_nand4_1 _15941_ (.B(net130),
    .C(_04768_),
    .A(_06842_),
    .Y(_06846_),
    .D(_06827_));
 sg13g2_buf_1 _15942_ (.A(_06846_),
    .X(_06847_));
 sg13g2_nand2_1 _15943_ (.Y(_06848_),
    .A(_06845_),
    .B(_06847_));
 sg13g2_xnor2_1 _15944_ (.Y(_06849_),
    .A(_04657_),
    .B(_04771_));
 sg13g2_nand2_1 _15945_ (.Y(_06850_),
    .A(_06848_),
    .B(_06849_));
 sg13g2_o21ai_1 _15946_ (.B1(_06850_),
    .Y(_06851_),
    .A1(net72),
    .A2(_06781_));
 sg13g2_buf_1 _15947_ (.A(\b.gen_square[51].sq.mask ),
    .X(_06852_));
 sg13g2_nand2_1 _15948_ (.Y(_06853_),
    .A(_06851_),
    .B(_06852_));
 sg13g2_nand2_1 _15949_ (.Y(_06854_),
    .A(_06502_),
    .B(_06853_));
 sg13g2_inv_2 _15950_ (.Y(_06855_),
    .A(_04081_));
 sg13g2_nor2_1 _15951_ (.A(_04070_),
    .B(_04073_),
    .Y(_06856_));
 sg13g2_nand2_1 _15952_ (.Y(_06857_),
    .A(_06856_),
    .B(_04072_));
 sg13g2_nor3_1 _15953_ (.A(_04072_),
    .B(_04073_),
    .C(_04071_),
    .Y(_06858_));
 sg13g2_inv_1 _15954_ (.Y(_06859_),
    .A(_06858_));
 sg13g2_a21o_1 _15955_ (.A2(_06859_),
    .A1(_06857_),
    .B1(_04347_),
    .X(_06860_));
 sg13g2_o21ai_1 _15956_ (.B1(_04092_),
    .Y(_06861_),
    .A1(_06855_),
    .A2(_06860_));
 sg13g2_buf_1 _15957_ (.A(_06861_),
    .X(_06862_));
 sg13g2_inv_1 _15958_ (.Y(_06863_),
    .A(_06862_));
 sg13g2_nor3_1 _15959_ (.A(_04099_),
    .B(_04102_),
    .C(_04106_),
    .Y(_06864_));
 sg13g2_nand2b_1 _15960_ (.Y(_06865_),
    .B(_04318_),
    .A_N(_06864_));
 sg13g2_nand2_1 _15961_ (.Y(_06866_),
    .A(_04314_),
    .B(_06865_));
 sg13g2_nand3_1 _15962_ (.B(_06866_),
    .C(_04105_),
    .A(_04113_),
    .Y(_06867_));
 sg13g2_inv_2 _15963_ (.Y(_06868_),
    .A(_06867_));
 sg13g2_a21oi_1 _15964_ (.A1(_06863_),
    .A2(net34),
    .Y(_06869_),
    .B1(_06868_));
 sg13g2_inv_1 _15965_ (.Y(_06870_),
    .A(_06869_));
 sg13g2_a21oi_1 _15966_ (.A1(_06870_),
    .A2(net71),
    .Y(_06871_),
    .B1(_04949_));
 sg13g2_and3_1 _15967_ (.X(_06872_),
    .A(_06014_),
    .B(_06023_),
    .C(_06015_));
 sg13g2_o21ai_1 _15968_ (.B1(net133),
    .Y(_06873_),
    .A1(_06034_),
    .A2(_06872_));
 sg13g2_inv_1 _15969_ (.Y(_06874_),
    .A(_06028_));
 sg13g2_o21ai_1 _15970_ (.B1(_06874_),
    .Y(_06875_),
    .A1(_06022_),
    .A2(_06873_));
 sg13g2_inv_1 _15971_ (.Y(_06876_),
    .A(_06875_));
 sg13g2_and3_1 _15972_ (.X(_06877_),
    .A(_05630_),
    .B(_05638_),
    .C(_05631_));
 sg13g2_o21ai_1 _15973_ (.B1(_05653_),
    .Y(_06878_),
    .A1(_05650_),
    .A2(_06877_));
 sg13g2_nand3_1 _15974_ (.B(_05635_),
    .C(_06878_),
    .A(_05643_),
    .Y(_06879_));
 sg13g2_inv_1 _15975_ (.Y(_06880_),
    .A(_06879_));
 sg13g2_a21oi_1 _15976_ (.A1(_06876_),
    .A2(net53),
    .Y(_06881_),
    .B1(_06880_));
 sg13g2_inv_1 _15977_ (.Y(_06882_),
    .A(_06881_));
 sg13g2_inv_1 _15978_ (.Y(_06883_),
    .A(_05922_));
 sg13g2_a21oi_1 _15979_ (.A1(_06882_),
    .A2(net28),
    .Y(_06884_),
    .B1(_06883_));
 sg13g2_inv_1 _15980_ (.Y(_06885_),
    .A(_06884_));
 sg13g2_a21oi_1 _15981_ (.A1(_06885_),
    .A2(net21),
    .Y(_06886_),
    .B1(_06241_));
 sg13g2_nor2_1 _15982_ (.A(_03362_),
    .B(_06030_),
    .Y(_06887_));
 sg13g2_buf_8 _15983_ (.A(_06887_),
    .X(_06888_));
 sg13g2_inv_4 _15984_ (.A(_06888_),
    .Y(_06889_));
 sg13g2_a21oi_2 _15985_ (.B1(_05718_),
    .Y(_06890_),
    .A2(_05646_),
    .A1(_06889_));
 sg13g2_inv_1 _15986_ (.Y(_06891_),
    .A(_05963_));
 sg13g2_o21ai_1 _15987_ (.B1(_06891_),
    .Y(_06892_),
    .A1(_05845_),
    .A2(_06890_));
 sg13g2_buf_1 _15988_ (.A(_06892_),
    .X(_06893_));
 sg13g2_a21oi_1 _15989_ (.A1(_06893_),
    .A2(net21),
    .Y(_06894_),
    .B1(_06201_));
 sg13g2_a221oi_1 _15990_ (.B2(_06894_),
    .C1(_06445_),
    .B1(_06886_),
    .A1(_06871_),
    .Y(_06895_),
    .A2(_04132_));
 sg13g2_nor2_1 _15991_ (.A(_05054_),
    .B(_06470_),
    .Y(_06896_));
 sg13g2_nand4_1 _15992_ (.B(_04460_),
    .C(_04444_),
    .A(_04451_),
    .Y(_06897_),
    .D(_04446_));
 sg13g2_o21ai_1 _15993_ (.B1(_04490_),
    .Y(_06898_),
    .A1(net32),
    .A2(_06897_));
 sg13g2_inv_1 _15994_ (.Y(_06899_),
    .A(_06898_));
 sg13g2_nor2_1 _15995_ (.A(_03985_),
    .B(_06899_),
    .Y(_06900_));
 sg13g2_nand4_1 _15996_ (.B(_04230_),
    .C(_04237_),
    .A(net165),
    .Y(_06901_),
    .D(_04232_));
 sg13g2_inv_1 _15997_ (.Y(_06902_),
    .A(_06901_));
 sg13g2_a21oi_1 _15998_ (.A1(_06902_),
    .A2(_04550_),
    .Y(_06903_),
    .B1(_04245_));
 sg13g2_nor2_1 _15999_ (.A(_03828_),
    .B(_06903_),
    .Y(_06904_));
 sg13g2_nor2_1 _16000_ (.A(_06904_),
    .B(_05019_),
    .Y(_06905_));
 sg13g2_inv_1 _16001_ (.Y(_06906_),
    .A(_06905_));
 sg13g2_nor4_1 _16002_ (.A(_06900_),
    .B(_06461_),
    .C(_06906_),
    .D(_05825_),
    .Y(_06907_));
 sg13g2_nor2_1 _16003_ (.A(_06831_),
    .B(_06455_),
    .Y(_06908_));
 sg13g2_o21ai_1 _16004_ (.B1(_06763_),
    .Y(_06909_),
    .A1(_04553_),
    .A2(_04991_));
 sg13g2_nand2_1 _16005_ (.Y(_06910_),
    .A(_06909_),
    .B(_06785_));
 sg13g2_nand2_1 _16006_ (.Y(_06911_),
    .A(_04564_),
    .B(_06910_));
 sg13g2_a21oi_1 _16007_ (.A1(_06911_),
    .A2(_04996_),
    .Y(_06912_),
    .B1(_05013_));
 sg13g2_nand3_1 _16008_ (.B(_06908_),
    .C(_06912_),
    .A(_06907_),
    .Y(_06913_));
 sg13g2_a21oi_1 _16009_ (.A1(_05731_),
    .A2(_05747_),
    .Y(_06914_),
    .B1(_06913_));
 sg13g2_nand3_1 _16010_ (.B(_06896_),
    .C(_06914_),
    .A(_06895_),
    .Y(_06915_));
 sg13g2_xnor2_1 _16011_ (.Y(_06916_),
    .A(_04642_),
    .B(_03870_));
 sg13g2_buf_1 _16012_ (.A(\b.gen_square[4].sq.piece[1] ),
    .X(_06917_));
 sg13g2_buf_2 _16013_ (.A(\b.gen_square[4].sq.piece[2] ),
    .X(_06918_));
 sg13g2_inv_2 _16014_ (.Y(_06919_),
    .A(_06918_));
 sg13g2_buf_1 _16015_ (.A(\b.gen_square[4].sq.piece[0] ),
    .X(_06920_));
 sg13g2_inv_1 _16016_ (.Y(_06921_),
    .A(_06920_));
 sg13g2_nor3_1 _16017_ (.A(_06917_),
    .B(_06919_),
    .C(_06921_),
    .Y(_06922_));
 sg13g2_inv_2 _16018_ (.Y(_06923_),
    .A(_06922_));
 sg13g2_nor2_1 _16019_ (.A(_06916_),
    .B(_06923_),
    .Y(_06924_));
 sg13g2_a22oi_1 _16020_ (.Y(_06925_),
    .B1(_04087_),
    .B2(_03867_),
    .A2(_04061_),
    .A1(_06924_));
 sg13g2_buf_1 _16021_ (.A(_06925_),
    .X(_06926_));
 sg13g2_nor2_1 _16022_ (.A(_06917_),
    .B(_06920_),
    .Y(_06927_));
 sg13g2_inv_1 _16023_ (.Y(_06928_),
    .A(_06927_));
 sg13g2_nor2_1 _16024_ (.A(_06919_),
    .B(_06928_),
    .Y(_06929_));
 sg13g2_nand2_1 _16025_ (.Y(_06930_),
    .A(_06917_),
    .B(_06920_));
 sg13g2_nor2_1 _16026_ (.A(_06918_),
    .B(_06930_),
    .Y(_06931_));
 sg13g2_inv_2 _16027_ (.Y(_06932_),
    .A(_06916_));
 sg13g2_nor2_1 _16028_ (.A(_06932_),
    .B(_04285_),
    .Y(_06933_));
 sg13g2_o21ai_1 _16029_ (.B1(_06933_),
    .Y(_06934_),
    .A1(_06929_),
    .A2(_06931_));
 sg13g2_nand2_1 _16030_ (.Y(_06935_),
    .A(_06926_),
    .B(_06934_));
 sg13g2_inv_1 _16031_ (.Y(_06936_),
    .A(_06935_));
 sg13g2_buf_1 _16032_ (.A(\b.gen_square[12].sq.piece[2] ),
    .X(_06937_));
 sg13g2_inv_1 _16033_ (.Y(_06938_),
    .A(_06937_));
 sg13g2_buf_1 _16034_ (.A(\b.gen_square[12].sq.piece[1] ),
    .X(_06939_));
 sg13g2_buf_1 _16035_ (.A(\b.gen_square[12].sq.piece[0] ),
    .X(_06940_));
 sg13g2_nand2_1 _16036_ (.Y(_06941_),
    .A(_06939_),
    .B(_06940_));
 sg13g2_nor2_1 _16037_ (.A(_06938_),
    .B(_06941_),
    .Y(_06942_));
 sg13g2_inv_1 _16038_ (.Y(_06943_),
    .A(_06942_));
 sg13g2_xnor2_1 _16039_ (.Y(_06944_),
    .A(_04076_),
    .B(\b.gen_square[12].sq.color ));
 sg13g2_buf_2 _16040_ (.A(_06944_),
    .X(_06945_));
 sg13g2_inv_1 _16041_ (.Y(_06946_),
    .A(_06940_));
 sg13g2_nor3_2 _16042_ (.A(_06939_),
    .B(_06938_),
    .C(_06946_),
    .Y(_06947_));
 sg13g2_inv_1 _16043_ (.Y(_06948_),
    .A(_06947_));
 sg13g2_nor2_1 _16044_ (.A(_06945_),
    .B(_06948_),
    .Y(_06949_));
 sg13g2_a22oi_1 _16045_ (.Y(_06950_),
    .B1(net152),
    .B2(_06949_),
    .A2(_04087_),
    .A1(_02814_));
 sg13g2_buf_2 _16046_ (.A(_06950_),
    .X(_06951_));
 sg13g2_inv_4 _16047_ (.A(_06951_),
    .Y(_06952_));
 sg13g2_nor2_1 _16048_ (.A(_06943_),
    .B(_06952_),
    .Y(_06953_));
 sg13g2_buf_1 _16049_ (.A(_06953_),
    .X(_06954_));
 sg13g2_buf_1 _16050_ (.A(net65),
    .X(_06955_));
 sg13g2_inv_1 _16051_ (.Y(_06956_),
    .A(_06945_));
 sg13g2_nor2_1 _16052_ (.A(_06956_),
    .B(net100),
    .Y(_06957_));
 sg13g2_nor2_1 _16053_ (.A(_06937_),
    .B(_06941_),
    .Y(_06958_));
 sg13g2_nor2_1 _16054_ (.A(_06939_),
    .B(_06940_),
    .Y(_06959_));
 sg13g2_nand2_1 _16055_ (.Y(_06960_),
    .A(_06959_),
    .B(_06937_));
 sg13g2_nand2b_1 _16056_ (.Y(_06961_),
    .B(_06960_),
    .A_N(_06958_));
 sg13g2_nand2_1 _16057_ (.Y(_06962_),
    .A(_06957_),
    .B(_06961_));
 sg13g2_nand3_1 _16058_ (.B(_06943_),
    .C(_06962_),
    .A(_06951_),
    .Y(_06963_));
 sg13g2_inv_1 _16059_ (.Y(_06964_),
    .A(_06963_));
 sg13g2_a21oi_1 _16060_ (.A1(_06936_),
    .A2(net49),
    .Y(_06965_),
    .B1(_06964_));
 sg13g2_inv_1 _16061_ (.Y(_06966_),
    .A(_06965_));
 sg13g2_nor2_1 _16062_ (.A(_05846_),
    .B(_05850_),
    .Y(_06967_));
 sg13g2_inv_1 _16063_ (.Y(_06968_),
    .A(_06967_));
 sg13g2_a21oi_1 _16064_ (.A1(_05902_),
    .A2(_06968_),
    .Y(_06969_),
    .B1(_05907_));
 sg13g2_nand3b_1 _16065_ (.B(_05860_),
    .C(_05852_),
    .Y(_06970_),
    .A_N(_06969_));
 sg13g2_inv_1 _16066_ (.Y(_06971_),
    .A(_06970_));
 sg13g2_a21oi_1 _16067_ (.A1(_06966_),
    .A2(_05953_),
    .Y(_06972_),
    .B1(_06971_));
 sg13g2_inv_1 _16068_ (.Y(_06973_),
    .A(_06972_));
 sg13g2_nor2_1 _16069_ (.A(_05329_),
    .B(_05333_),
    .Y(_06974_));
 sg13g2_inv_1 _16070_ (.Y(_06975_),
    .A(_06974_));
 sg13g2_nand2_1 _16071_ (.Y(_06976_),
    .A(_06975_),
    .B(_05350_));
 sg13g2_nand2_1 _16072_ (.Y(_06977_),
    .A(_05353_),
    .B(_06976_));
 sg13g2_nand3_1 _16073_ (.B(_05335_),
    .C(_06977_),
    .A(_05343_),
    .Y(_06978_));
 sg13g2_inv_1 _16074_ (.Y(_06979_),
    .A(_06978_));
 sg13g2_a21oi_2 _16075_ (.B1(_06979_),
    .Y(_06980_),
    .A2(net40),
    .A1(_06973_));
 sg13g2_o21ai_1 _16076_ (.B1(_04933_),
    .Y(_06981_),
    .A1(_04910_),
    .A2(_04914_));
 sg13g2_nand2_1 _16077_ (.Y(_06982_),
    .A(_04930_),
    .B(_06981_));
 sg13g2_nand3_1 _16078_ (.B(_04916_),
    .C(_06982_),
    .A(_04924_),
    .Y(_06983_));
 sg13g2_buf_1 _16079_ (.A(_06983_),
    .X(_06984_));
 sg13g2_o21ai_1 _16080_ (.B1(_06984_),
    .Y(_06985_),
    .A1(_06203_),
    .A2(_06980_));
 sg13g2_buf_1 _16081_ (.A(_06985_),
    .X(_06986_));
 sg13g2_nor2_1 _16082_ (.A(_04514_),
    .B(_06659_),
    .Y(_06987_));
 sg13g2_o21ai_1 _16083_ (.B1(_06714_),
    .Y(_06988_),
    .A1(_06711_),
    .A2(_06987_));
 sg13g2_nand3_1 _16084_ (.B(_04524_),
    .C(_06716_),
    .A(_06988_),
    .Y(_06989_));
 sg13g2_inv_1 _16085_ (.Y(_06990_),
    .A(_06989_));
 sg13g2_a21oi_2 _16086_ (.B1(_06990_),
    .Y(_06991_),
    .A2(net66),
    .A1(_06986_));
 sg13g2_nor2_2 _16087_ (.A(_06919_),
    .B(_06930_),
    .Y(_06992_));
 sg13g2_inv_1 _16088_ (.Y(_06993_),
    .A(_06992_));
 sg13g2_inv_2 _16089_ (.Y(_06994_),
    .A(_06926_));
 sg13g2_nor2_1 _16090_ (.A(_06993_),
    .B(_06994_),
    .Y(_06995_));
 sg13g2_buf_2 _16091_ (.A(_06995_),
    .X(_06996_));
 sg13g2_nor2_1 _16092_ (.A(_00055_),
    .B(_06996_),
    .Y(_06997_));
 sg13g2_buf_2 _16093_ (.A(_06997_),
    .X(_06998_));
 sg13g2_inv_1 _16094_ (.Y(_06999_),
    .A(_06998_));
 sg13g2_inv_1 _16095_ (.Y(_07000_),
    .A(_00054_));
 sg13g2_nor2_1 _16096_ (.A(_07000_),
    .B(net65),
    .Y(_07001_));
 sg13g2_buf_2 _16097_ (.A(_07001_),
    .X(_07002_));
 sg13g2_a21oi_1 _16098_ (.A1(_06999_),
    .A2(net49),
    .Y(_07003_),
    .B1(_07002_));
 sg13g2_inv_1 _16099_ (.Y(_07004_),
    .A(_07003_));
 sg13g2_a21oi_1 _16100_ (.A1(_07004_),
    .A2(_05953_),
    .Y(_07005_),
    .B1(_05956_));
 sg13g2_inv_1 _16101_ (.Y(_07006_),
    .A(_07005_));
 sg13g2_a21oi_1 _16102_ (.A1(_07006_),
    .A2(net40),
    .Y(_07007_),
    .B1(_05532_));
 sg13g2_inv_1 _16103_ (.Y(_07008_),
    .A(_07007_));
 sg13g2_a21oi_1 _16104_ (.A1(_07008_),
    .A2(net58),
    .Y(_07009_),
    .B1(_04972_));
 sg13g2_inv_1 _16105_ (.Y(_07010_),
    .A(_07009_));
 sg13g2_a21oi_1 _16106_ (.A1(_07010_),
    .A2(net66),
    .Y(_07011_),
    .B1(_06737_));
 sg13g2_a22oi_1 _16107_ (.Y(_07012_),
    .B1(_06991_),
    .B2(_07011_),
    .A2(_04777_),
    .A1(_04679_));
 sg13g2_nand2_1 _16108_ (.Y(_07013_),
    .A(_05066_),
    .B(_06734_));
 sg13g2_inv_2 _16109_ (.Y(_07014_),
    .A(_06737_));
 sg13g2_nand2_1 _16110_ (.Y(_07015_),
    .A(_07013_),
    .B(_07014_));
 sg13g2_nor2_1 _16111_ (.A(_06793_),
    .B(_07015_),
    .Y(_07016_));
 sg13g2_buf_2 _16112_ (.A(_07016_),
    .X(_07017_));
 sg13g2_nor4_1 _16113_ (.A(_05067_),
    .B(_05010_),
    .C(_06454_),
    .D(_07017_),
    .Y(_07018_));
 sg13g2_nand2_1 _16114_ (.Y(_07019_),
    .A(_07012_),
    .B(_07018_));
 sg13g2_nor2_1 _16115_ (.A(_06915_),
    .B(_07019_),
    .Y(_07020_));
 sg13g2_inv_1 _16116_ (.Y(_07021_),
    .A(_07020_));
 sg13g2_inv_1 _16117_ (.Y(_07022_),
    .A(_07011_));
 sg13g2_inv_1 _16118_ (.Y(_07023_),
    .A(_04134_));
 sg13g2_nand2_1 _16119_ (.Y(_07024_),
    .A(_07023_),
    .B(_06314_));
 sg13g2_a221oi_1 _16120_ (.B2(_06991_),
    .C1(_07024_),
    .B1(_07022_),
    .A1(_05732_),
    .Y(_07025_),
    .A2(_05747_));
 sg13g2_nor2_1 _16121_ (.A(_04999_),
    .B(_06795_),
    .Y(_07026_));
 sg13g2_a21oi_1 _16122_ (.A1(_04778_),
    .A2(_06247_),
    .Y(_07027_),
    .B1(_04679_));
 sg13g2_nor2b_1 _16123_ (.A(_06903_),
    .B_N(_00070_),
    .Y(_07028_));
 sg13g2_buf_1 _16124_ (.A(_07028_),
    .X(_07029_));
 sg13g2_nor2_1 _16125_ (.A(_05063_),
    .B(_06899_),
    .Y(_07030_));
 sg13g2_nor2_1 _16126_ (.A(_07030_),
    .B(_04548_),
    .Y(_07031_));
 sg13g2_inv_1 _16127_ (.Y(_07032_),
    .A(_07031_));
 sg13g2_nor4_2 _16128_ (.A(_07029_),
    .B(_06296_),
    .C(_07032_),
    .Y(_07033_),
    .D(_05833_));
 sg13g2_inv_1 _16129_ (.Y(_07034_),
    .A(_04383_));
 sg13g2_nand2_1 _16130_ (.Y(_07035_),
    .A(_06911_),
    .B(_03968_));
 sg13g2_nor2_1 _16131_ (.A(_06787_),
    .B(_04996_),
    .Y(_07036_));
 sg13g2_nor2_1 _16132_ (.A(_07036_),
    .B(_06264_),
    .Y(_07037_));
 sg13g2_nand4_1 _16133_ (.B(_07034_),
    .C(_07035_),
    .A(_07033_),
    .Y(_07038_),
    .D(_07037_));
 sg13g2_inv_1 _16134_ (.Y(_07039_),
    .A(_06886_));
 sg13g2_inv_1 _16135_ (.Y(_07040_),
    .A(_04132_));
 sg13g2_a21oi_1 _16136_ (.A1(_07040_),
    .A2(_06871_),
    .Y(_07041_),
    .B1(_06275_));
 sg13g2_o21ai_1 _16137_ (.B1(_07041_),
    .Y(_07042_),
    .A1(_06894_),
    .A2(_07039_));
 sg13g2_nor4_1 _16138_ (.A(_04479_),
    .B(_07027_),
    .C(_07038_),
    .D(_07042_),
    .Y(_07043_));
 sg13g2_nand3_1 _16139_ (.B(_07026_),
    .C(_07043_),
    .A(_07025_),
    .Y(_07044_));
 sg13g2_nor2_1 _16140_ (.A(_07021_),
    .B(_07044_),
    .Y(_07045_));
 sg13g2_nand2_1 _16141_ (.Y(_07046_),
    .A(_04779_),
    .B(net68));
 sg13g2_nand4_1 _16142_ (.B(net114),
    .C(_04779_),
    .A(_07044_),
    .Y(_07047_),
    .D(_07021_));
 sg13g2_buf_1 _16143_ (.A(_07047_),
    .X(_07048_));
 sg13g2_o21ai_1 _16144_ (.B1(_07048_),
    .Y(_07049_),
    .A1(_07045_),
    .A2(_07046_));
 sg13g2_xnor2_1 _16145_ (.Y(_07050_),
    .A(_04681_),
    .B(_04782_));
 sg13g2_nand2_1 _16146_ (.Y(_07051_),
    .A(_06895_),
    .B(_04478_));
 sg13g2_o21ai_1 _16147_ (.B1(_04689_),
    .Y(_07052_),
    .A1(_07042_),
    .A2(_07051_));
 sg13g2_and3_1 _16148_ (.X(_07053_),
    .A(_04682_),
    .B(_04690_),
    .C(_04683_));
 sg13g2_nand2b_1 _16149_ (.Y(_07054_),
    .B(_07053_),
    .A_N(_07052_));
 sg13g2_nor3_1 _16150_ (.A(_04681_),
    .B(_04683_),
    .C(_04690_),
    .Y(_07055_));
 sg13g2_nand2_1 _16151_ (.Y(_07056_),
    .A(_04689_),
    .B(_07055_));
 sg13g2_a21o_1 _16152_ (.A2(_07033_),
    .A1(_06907_),
    .B1(_07056_),
    .X(_07057_));
 sg13g2_nand2_1 _16153_ (.Y(_07058_),
    .A(_04692_),
    .B(net67));
 sg13g2_a21oi_1 _16154_ (.A1(_07054_),
    .A2(_07057_),
    .Y(_07059_),
    .B1(_07058_));
 sg13g2_a21oi_1 _16155_ (.A1(_07049_),
    .A2(_07050_),
    .Y(_07060_),
    .B1(_07059_));
 sg13g2_inv_1 _16156_ (.Y(_07061_),
    .A(_06911_));
 sg13g2_nand3_1 _16157_ (.B(_07061_),
    .C(_05748_),
    .A(_04778_),
    .Y(_07062_));
 sg13g2_o21ai_1 _16158_ (.B1(_04689_),
    .Y(_07063_),
    .A1(_07062_),
    .A2(_06991_));
 sg13g2_a21o_1 _16159_ (.A2(_07063_),
    .A1(_07052_),
    .B1(_04783_),
    .X(_07064_));
 sg13g2_nand2b_1 _16160_ (.Y(_07065_),
    .B(_04781_),
    .A_N(_07063_));
 sg13g2_a21o_1 _16161_ (.A2(_07065_),
    .A1(_07064_),
    .B1(_07058_),
    .X(_07066_));
 sg13g2_inv_1 _16162_ (.Y(_07067_),
    .A(\b.gen_square[52].sq.mask ));
 sg13g2_a21o_1 _16163_ (.A2(_07066_),
    .A1(_07060_),
    .B1(_07067_),
    .X(_07068_));
 sg13g2_buf_1 _16164_ (.A(_07068_),
    .X(_07069_));
 sg13g2_nor2b_1 _16165_ (.A(_06854_),
    .B_N(_07069_),
    .Y(_07070_));
 sg13g2_buf_1 _16166_ (.A(net73),
    .X(_07071_));
 sg13g2_buf_1 _16167_ (.A(\b.gen_square[5].sq.piece[2] ),
    .X(_07072_));
 sg13g2_inv_2 _16168_ (.Y(_07073_),
    .A(_07072_));
 sg13g2_buf_2 _16169_ (.A(\b.gen_square[5].sq.piece[0] ),
    .X(_07074_));
 sg13g2_nand2_1 _16170_ (.Y(_07075_),
    .A(\b.gen_square[5].sq.piece[1] ),
    .B(_07074_));
 sg13g2_inv_1 _16171_ (.Y(_07076_),
    .A(_07075_));
 sg13g2_nor2_1 _16172_ (.A(\b.gen_square[5].sq.piece[1] ),
    .B(_07074_),
    .Y(_07077_));
 sg13g2_inv_1 _16173_ (.Y(_07078_),
    .A(_07077_));
 sg13g2_nor2_1 _16174_ (.A(_07073_),
    .B(_07078_),
    .Y(_07079_));
 sg13g2_a21oi_1 _16175_ (.A1(_07073_),
    .A2(_07076_),
    .Y(_07080_),
    .B1(_07079_));
 sg13g2_xnor2_1 _16176_ (.Y(_07081_),
    .A(net193),
    .B(\b.gen_square[5].sq.color ));
 sg13g2_inv_2 _16177_ (.Y(_07082_),
    .A(_07081_));
 sg13g2_nor2_1 _16178_ (.A(_07082_),
    .B(net119),
    .Y(_07083_));
 sg13g2_inv_2 _16179_ (.Y(_07084_),
    .A(_07083_));
 sg13g2_nor2_1 _16180_ (.A(_07080_),
    .B(_07084_),
    .Y(_07085_));
 sg13g2_inv_1 _16181_ (.Y(_07086_),
    .A(\b.gen_square[5].sq.piece[1] ));
 sg13g2_nand3_1 _16182_ (.B(_07072_),
    .C(_07074_),
    .A(_07086_),
    .Y(_07087_));
 sg13g2_buf_1 _16183_ (.A(_07087_),
    .X(_07088_));
 sg13g2_nor2_1 _16184_ (.A(_07088_),
    .B(_07081_),
    .Y(_07089_));
 sg13g2_a22oi_1 _16185_ (.Y(_07090_),
    .B1(net151),
    .B2(_03961_),
    .A2(net148),
    .A1(_07089_));
 sg13g2_inv_2 _16186_ (.Y(_07091_),
    .A(_07090_));
 sg13g2_nor2_1 _16187_ (.A(_07085_),
    .B(_07091_),
    .Y(_07092_));
 sg13g2_o21ai_1 _16188_ (.B1(_05895_),
    .Y(_07093_),
    .A1(_05873_),
    .A2(_05877_));
 sg13g2_nand2_1 _16189_ (.Y(_07094_),
    .A(_05892_),
    .B(_07093_));
 sg13g2_nand3_1 _16190_ (.B(_05879_),
    .C(_07094_),
    .A(_05887_),
    .Y(_07095_));
 sg13g2_buf_1 _16191_ (.A(_07095_),
    .X(_07096_));
 sg13g2_inv_1 _16192_ (.Y(_07097_),
    .A(_07096_));
 sg13g2_a21oi_1 _16193_ (.A1(net64),
    .A2(_07092_),
    .Y(_07098_),
    .B1(_07097_));
 sg13g2_inv_1 _16194_ (.Y(_07099_),
    .A(_07098_));
 sg13g2_buf_1 _16195_ (.A(_05289_),
    .X(_07100_));
 sg13g2_nor2_1 _16196_ (.A(_05272_),
    .B(_05276_),
    .Y(_07101_));
 sg13g2_inv_1 _16197_ (.Y(_07102_),
    .A(_07101_));
 sg13g2_nand2_1 _16198_ (.Y(_07103_),
    .A(_07102_),
    .B(_05324_));
 sg13g2_nand2_1 _16199_ (.Y(_07104_),
    .A(_05320_),
    .B(_07103_));
 sg13g2_nand3_1 _16200_ (.B(_05278_),
    .C(_07104_),
    .A(_05286_),
    .Y(_07105_));
 sg13g2_inv_1 _16201_ (.Y(_07106_),
    .A(_07105_));
 sg13g2_a21oi_1 _16202_ (.A1(_07099_),
    .A2(net25),
    .Y(_07107_),
    .B1(_07106_));
 sg13g2_inv_1 _16203_ (.Y(_07108_),
    .A(_07107_));
 sg13g2_nor2_1 _16204_ (.A(_06172_),
    .B(_06182_),
    .Y(_07109_));
 sg13g2_inv_1 _16205_ (.Y(_07110_),
    .A(_07109_));
 sg13g2_nand2_1 _16206_ (.Y(_07111_),
    .A(_07110_),
    .B(_06225_));
 sg13g2_nand2_1 _16207_ (.Y(_07112_),
    .A(_06222_),
    .B(_07111_));
 sg13g2_nand3_1 _16208_ (.B(_06220_),
    .C(_07112_),
    .A(_06180_),
    .Y(_07113_));
 sg13g2_inv_1 _16209_ (.Y(_07114_),
    .A(_07113_));
 sg13g2_a21oi_1 _16210_ (.A1(_07108_),
    .A2(net27),
    .Y(_07115_),
    .B1(_07114_));
 sg13g2_inv_1 _16211_ (.Y(_07116_),
    .A(_07115_));
 sg13g2_nor2_1 _16212_ (.A(_04533_),
    .B(_06692_),
    .Y(_07117_));
 sg13g2_inv_1 _16213_ (.Y(_07118_),
    .A(_07117_));
 sg13g2_nand2_1 _16214_ (.Y(_07119_),
    .A(_07118_),
    .B(_06702_));
 sg13g2_nand2_1 _16215_ (.Y(_07120_),
    .A(_06699_),
    .B(_07119_));
 sg13g2_nand3_1 _16216_ (.B(_06694_),
    .C(_07120_),
    .A(_04545_),
    .Y(_07121_));
 sg13g2_inv_1 _16217_ (.Y(_07122_),
    .A(_07121_));
 sg13g2_a21oi_2 _16218_ (.B1(_07122_),
    .Y(_07123_),
    .A2(net50),
    .A1(_07116_));
 sg13g2_o21ai_1 _16219_ (.B1(_04943_),
    .Y(_07124_),
    .A1(_04055_),
    .A2(_04124_));
 sg13g2_nand2_1 _16220_ (.Y(_07125_),
    .A(_04052_),
    .B(_07124_));
 sg13g2_nand3_1 _16221_ (.B(_04946_),
    .C(_07125_),
    .A(_04067_),
    .Y(_07126_));
 sg13g2_buf_1 _16222_ (.A(_07126_),
    .X(_07127_));
 sg13g2_o21ai_1 _16223_ (.B1(_07127_),
    .Y(_07128_),
    .A1(_04127_),
    .A2(_07123_));
 sg13g2_inv_1 _16224_ (.Y(_07129_),
    .A(_07128_));
 sg13g2_nor2_1 _16225_ (.A(_07073_),
    .B(_07075_),
    .Y(_07130_));
 sg13g2_inv_1 _16226_ (.Y(_07131_),
    .A(_07130_));
 sg13g2_nor2_1 _16227_ (.A(_07131_),
    .B(_07091_),
    .Y(_07132_));
 sg13g2_buf_1 _16228_ (.A(_07132_),
    .X(_07133_));
 sg13g2_inv_2 _16229_ (.Y(_07134_),
    .A(_07133_));
 sg13g2_inv_1 _16230_ (.Y(_07135_),
    .A(_00048_));
 sg13g2_nand2_1 _16231_ (.Y(_07136_),
    .A(_07134_),
    .B(_07135_));
 sg13g2_buf_2 _16232_ (.A(_07136_),
    .X(_07137_));
 sg13g2_a21oi_1 _16233_ (.A1(_07137_),
    .A2(net64),
    .Y(_07138_),
    .B1(_05950_));
 sg13g2_inv_1 _16234_ (.Y(_07139_),
    .A(_07138_));
 sg13g2_a21oi_1 _16235_ (.A1(_07139_),
    .A2(net25),
    .Y(_07140_),
    .B1(_05527_));
 sg13g2_inv_1 _16236_ (.Y(_07141_),
    .A(_07140_));
 sg13g2_a21oi_1 _16237_ (.A1(_07141_),
    .A2(net27),
    .Y(_07142_),
    .B1(_06189_));
 sg13g2_inv_1 _16238_ (.Y(_07143_),
    .A(_07142_));
 sg13g2_a21oi_1 _16239_ (.A1(_07143_),
    .A2(net50),
    .Y(_07144_),
    .B1(_06731_));
 sg13g2_inv_1 _16240_ (.Y(_07145_),
    .A(_07144_));
 sg13g2_a21oi_1 _16241_ (.A1(_07145_),
    .A2(net71),
    .Y(_07146_),
    .B1(_04131_));
 sg13g2_a22oi_1 _16242_ (.Y(_07147_),
    .B1(_07129_),
    .B2(_07146_),
    .A2(_04788_),
    .A1(_04703_));
 sg13g2_o21ai_1 _16243_ (.B1(_05742_),
    .Y(_07148_),
    .A1(_05040_),
    .A2(_05739_));
 sg13g2_inv_1 _16244_ (.Y(_07149_),
    .A(_07148_));
 sg13g2_nor2_2 _16245_ (.A(_07149_),
    .B(_05050_),
    .Y(_07150_));
 sg13g2_nor4_1 _16246_ (.A(_07150_),
    .B(_05008_),
    .C(_05054_),
    .D(_06830_),
    .Y(_07151_));
 sg13g2_nor2_1 _16247_ (.A(_04364_),
    .B(_04377_),
    .Y(_07152_));
 sg13g2_nor2_1 _16248_ (.A(_07152_),
    .B(_04474_),
    .Y(_07153_));
 sg13g2_nor3_1 _16249_ (.A(_04362_),
    .B(net61),
    .C(_07153_),
    .Y(_07154_));
 sg13g2_nor2_1 _16250_ (.A(_07154_),
    .B(_04374_),
    .Y(_07155_));
 sg13g2_inv_1 _16251_ (.Y(_07156_),
    .A(_07155_));
 sg13g2_nand4_1 _16252_ (.B(_04100_),
    .C(_04106_),
    .A(_04110_),
    .Y(_07157_),
    .D(_04102_));
 sg13g2_inv_1 _16253_ (.Y(_07158_),
    .A(_07157_));
 sg13g2_a21oi_1 _16254_ (.A1(net60),
    .A2(_07158_),
    .Y(_07159_),
    .B1(_04114_));
 sg13g2_nor2_1 _16255_ (.A(_03749_),
    .B(_07159_),
    .Y(_07160_));
 sg13g2_nor2_1 _16256_ (.A(_07160_),
    .B(_06646_),
    .Y(_07161_));
 sg13g2_nand4_1 _16257_ (.B(_04421_),
    .C(_04411_),
    .A(_04416_),
    .Y(_07162_),
    .D(_04413_));
 sg13g2_inv_1 _16258_ (.Y(_07163_),
    .A(_07162_));
 sg13g2_a21oi_1 _16259_ (.A1(_07163_),
    .A2(net60),
    .Y(_07164_),
    .B1(_04429_));
 sg13g2_nor2_1 _16260_ (.A(_03993_),
    .B(_07164_),
    .Y(_07165_));
 sg13g2_nor3_1 _16261_ (.A(_04385_),
    .B(_04384_),
    .C(_04388_),
    .Y(_07166_));
 sg13g2_nand2_1 _16262_ (.Y(_07167_),
    .A(_04391_),
    .B(_07166_));
 sg13g2_inv_1 _16263_ (.Y(_07168_),
    .A(_07167_));
 sg13g2_a21oi_1 _16264_ (.A1(net60),
    .A2(_07168_),
    .Y(_07169_),
    .B1(_04399_));
 sg13g2_nor2_1 _16265_ (.A(_03839_),
    .B(_07169_),
    .Y(_07170_));
 sg13g2_nor2_1 _16266_ (.A(_07165_),
    .B(_07170_),
    .Y(_07171_));
 sg13g2_and3_1 _16267_ (.X(_07172_),
    .A(_07161_),
    .B(_05210_),
    .C(_07171_));
 sg13g2_inv_1 _16268_ (.Y(_07173_),
    .A(_07172_));
 sg13g2_a221oi_1 _16269_ (.B2(_05745_),
    .C1(_07173_),
    .B1(_05729_),
    .A1(_07156_),
    .Y(_07174_),
    .A2(_04382_));
 sg13g2_nor2_1 _16270_ (.A(_05062_),
    .B(_07017_),
    .Y(_07175_));
 sg13g2_nor2_1 _16271_ (.A(_06831_),
    .B(_05010_),
    .Y(_07176_));
 sg13g2_nand3_1 _16272_ (.B(_07175_),
    .C(_07176_),
    .A(_07174_),
    .Y(_07177_));
 sg13g2_nor2_1 _16273_ (.A(_04018_),
    .B(_05995_),
    .Y(_07178_));
 sg13g2_buf_2 _16274_ (.A(_07178_),
    .X(_07179_));
 sg13g2_inv_1 _16275_ (.Y(_07180_),
    .A(_07179_));
 sg13g2_a21oi_1 _16276_ (.A1(_07180_),
    .A2(_05710_),
    .Y(_07181_),
    .B1(_05713_));
 sg13g2_inv_1 _16277_ (.Y(_07182_),
    .A(_07181_));
 sg13g2_a21oi_1 _16278_ (.A1(_07182_),
    .A2(net51),
    .Y(_07183_),
    .B1(_06433_));
 sg13g2_inv_1 _16279_ (.Y(_07184_),
    .A(_07183_));
 sg13g2_a21oi_1 _16280_ (.A1(_07184_),
    .A2(net54),
    .Y(_07185_),
    .B1(_05537_));
 sg13g2_inv_1 _16281_ (.Y(_07186_),
    .A(_07185_));
 sg13g2_a21oi_1 _16282_ (.A1(_07186_),
    .A2(net66),
    .Y(_07187_),
    .B1(_06737_));
 sg13g2_nor3_1 _16283_ (.A(_05979_),
    .B(_05982_),
    .C(_05986_),
    .Y(_07188_));
 sg13g2_o21ai_1 _16284_ (.B1(net115),
    .Y(_07189_),
    .A1(_07188_),
    .A2(_06005_));
 sg13g2_o21ai_1 _16285_ (.B1(_05992_),
    .Y(_07190_),
    .A1(_06001_),
    .A2(_07189_));
 sg13g2_inv_1 _16286_ (.Y(_07191_),
    .A(_07190_));
 sg13g2_inv_1 _16287_ (.Y(_07192_),
    .A(_05580_));
 sg13g2_and3_1 _16288_ (.X(_07193_),
    .A(_05586_),
    .B(_07192_),
    .C(_05578_));
 sg13g2_o21ai_1 _16289_ (.B1(_05623_),
    .Y(_07194_),
    .A1(_05620_),
    .A2(_07193_));
 sg13g2_nand3_1 _16290_ (.B(_07194_),
    .C(_05625_),
    .A(_05585_),
    .Y(_07195_));
 sg13g2_inv_1 _16291_ (.Y(_07196_),
    .A(_07195_));
 sg13g2_a21oi_2 _16292_ (.B1(_07196_),
    .Y(_07197_),
    .A2(net38),
    .A1(_07191_));
 sg13g2_inv_1 _16293_ (.Y(_07198_),
    .A(_07197_));
 sg13g2_nand3_1 _16294_ (.B(_06382_),
    .C(_06375_),
    .A(_06374_),
    .Y(_07199_));
 sg13g2_a21o_1 _16295_ (.A2(_07199_),
    .A1(_06394_),
    .B1(_06399_),
    .X(_07200_));
 sg13g2_nand3_1 _16296_ (.B(_06388_),
    .C(_06379_),
    .A(_07200_),
    .Y(_07201_));
 sg13g2_buf_1 _16297_ (.A(_07201_),
    .X(_07202_));
 sg13g2_inv_1 _16298_ (.Y(_07203_),
    .A(_07202_));
 sg13g2_a21oi_1 _16299_ (.A1(_07198_),
    .A2(net51),
    .Y(_07204_),
    .B1(_07203_));
 sg13g2_inv_1 _16300_ (.Y(_07205_),
    .A(_07204_));
 sg13g2_a21oi_2 _16301_ (.B1(_05387_),
    .Y(_07206_),
    .A2(net54),
    .A1(_07205_));
 sg13g2_inv_1 _16302_ (.Y(_07207_),
    .A(_07206_));
 sg13g2_inv_1 _16303_ (.Y(_07208_),
    .A(_06718_));
 sg13g2_a21oi_1 _16304_ (.A1(_07207_),
    .A2(net66),
    .Y(_07209_),
    .B1(_07208_));
 sg13g2_nand2_1 _16305_ (.Y(_07210_),
    .A(_07187_),
    .B(_07209_));
 sg13g2_inv_1 _16306_ (.Y(_07211_),
    .A(_04446_));
 sg13g2_nand3_1 _16307_ (.B(_07211_),
    .C(_04443_),
    .A(_04460_),
    .Y(_07212_));
 sg13g2_nand2_1 _16308_ (.Y(_07213_),
    .A(_07212_),
    .B(_04492_));
 sg13g2_nand2_1 _16309_ (.Y(_07214_),
    .A(net147),
    .B(_07213_));
 sg13g2_nor2_1 _16310_ (.A(_04452_),
    .B(_07214_),
    .Y(_07215_));
 sg13g2_nor2_1 _16311_ (.A(_07215_),
    .B(_04457_),
    .Y(_07216_));
 sg13g2_nand2b_1 _16312_ (.Y(_07217_),
    .B(_04466_),
    .A_N(_07216_));
 sg13g2_nor2_1 _16313_ (.A(_04572_),
    .B(_04573_),
    .Y(_07218_));
 sg13g2_inv_1 _16314_ (.Y(_07219_),
    .A(_07218_));
 sg13g2_nor2_1 _16315_ (.A(_04980_),
    .B(_07219_),
    .Y(_07220_));
 sg13g2_inv_1 _16316_ (.Y(_07221_),
    .A(_07220_));
 sg13g2_nand3_1 _16317_ (.B(_04574_),
    .C(_04572_),
    .A(_04980_),
    .Y(_07222_));
 sg13g2_a21oi_1 _16318_ (.A1(_07221_),
    .A2(_07222_),
    .Y(_07223_),
    .B1(net61));
 sg13g2_a21oi_1 _16319_ (.A1(_04570_),
    .A2(_07223_),
    .Y(_07224_),
    .B1(_04583_));
 sg13g2_buf_2 _16320_ (.A(_07224_),
    .X(_07225_));
 sg13g2_inv_1 _16321_ (.Y(_07226_),
    .A(_04232_));
 sg13g2_nand3_1 _16322_ (.B(_07226_),
    .C(_04231_),
    .A(_04230_),
    .Y(_07227_));
 sg13g2_nand2_1 _16323_ (.Y(_07228_),
    .A(_07227_),
    .B(_04329_));
 sg13g2_nand2_1 _16324_ (.Y(_07229_),
    .A(_04326_),
    .B(_07228_));
 sg13g2_nand3_1 _16325_ (.B(_07229_),
    .C(_04235_),
    .A(_04324_),
    .Y(_07230_));
 sg13g2_inv_1 _16326_ (.Y(_07231_),
    .A(_07230_));
 sg13g2_a21oi_1 _16327_ (.A1(_07225_),
    .A2(net82),
    .Y(_07232_),
    .B1(_07231_));
 sg13g2_a21oi_1 _16328_ (.A1(_07232_),
    .A2(_04986_),
    .Y(_07233_),
    .B1(_06767_));
 sg13g2_nand3_1 _16329_ (.B(_07217_),
    .C(_07233_),
    .A(_07210_),
    .Y(_07234_));
 sg13g2_nor2_1 _16330_ (.A(_07177_),
    .B(_07234_),
    .Y(_07235_));
 sg13g2_and3_1 _16331_ (.X(_07236_),
    .A(_07147_),
    .B(_07151_),
    .C(_07235_));
 sg13g2_inv_1 _16332_ (.Y(_07237_),
    .A(_07146_));
 sg13g2_a22oi_1 _16333_ (.Y(_07238_),
    .B1(_07129_),
    .B2(_07237_),
    .A2(_05745_),
    .A1(_05730_));
 sg13g2_a21oi_2 _16334_ (.B1(_05728_),
    .Y(_07239_),
    .A2(net98),
    .A1(_05064_));
 sg13g2_nor2_1 _16335_ (.A(_07149_),
    .B(_07239_),
    .Y(_07240_));
 sg13g2_buf_1 _16336_ (.A(_07240_),
    .X(_07241_));
 sg13g2_nor2_1 _16337_ (.A(_07241_),
    .B(_04134_),
    .Y(_07242_));
 sg13g2_nor2_1 _16338_ (.A(_04988_),
    .B(_06795_),
    .Y(_07243_));
 sg13g2_nor2_1 _16339_ (.A(_04789_),
    .B(_04703_),
    .Y(_07244_));
 sg13g2_nor2b_1 _16340_ (.A(_07187_),
    .B_N(_07209_),
    .Y(_07245_));
 sg13g2_nor2_2 _16341_ (.A(_04118_),
    .B(_07159_),
    .Y(_07246_));
 sg13g2_nand2b_1 _16342_ (.Y(_07247_),
    .B(_00033_),
    .A_N(_07164_));
 sg13g2_nand2_1 _16343_ (.Y(_07248_),
    .A(_05202_),
    .B(_07247_));
 sg13g2_inv_1 _16344_ (.Y(_07249_),
    .A(_00015_));
 sg13g2_nor2_1 _16345_ (.A(_07249_),
    .B(_07169_),
    .Y(_07250_));
 sg13g2_nor2_1 _16346_ (.A(_05183_),
    .B(_07250_),
    .Y(_07251_));
 sg13g2_inv_1 _16347_ (.Y(_07252_),
    .A(_07251_));
 sg13g2_nor4_1 _16348_ (.A(_07246_),
    .B(_06641_),
    .C(_07248_),
    .D(_07252_),
    .Y(_07253_));
 sg13g2_nor2_1 _16349_ (.A(_07216_),
    .B(_04466_),
    .Y(_07254_));
 sg13g2_nor2_1 _16350_ (.A(_04467_),
    .B(_07254_),
    .Y(_07255_));
 sg13g2_nor2_1 _16351_ (.A(_07036_),
    .B(_04383_),
    .Y(_07256_));
 sg13g2_and3_1 _16352_ (.X(_07257_),
    .A(_07253_),
    .B(_07255_),
    .C(_07256_));
 sg13g2_inv_1 _16353_ (.Y(_07258_),
    .A(_06825_));
 sg13g2_inv_1 _16354_ (.Y(_07259_),
    .A(_04986_));
 sg13g2_a21oi_1 _16355_ (.A1(_07259_),
    .A2(_07232_),
    .Y(_07260_),
    .B1(_06775_));
 sg13g2_nand2_1 _16356_ (.Y(_07261_),
    .A(_07156_),
    .B(_03976_));
 sg13g2_nand4_1 _16357_ (.B(_07258_),
    .C(_07260_),
    .A(_07257_),
    .Y(_07262_),
    .D(_07261_));
 sg13g2_nor3_1 _16358_ (.A(_07244_),
    .B(_07245_),
    .C(_07262_),
    .Y(_07263_));
 sg13g2_and4_1 _16359_ (.A(_07238_),
    .B(_07242_),
    .C(_07243_),
    .D(_07263_),
    .X(_07264_));
 sg13g2_nor3_1 _16360_ (.A(_04717_),
    .B(_07236_),
    .C(_07264_),
    .Y(_07265_));
 sg13g2_nand2_1 _16361_ (.Y(_07266_),
    .A(_07265_),
    .B(net114));
 sg13g2_nand2_1 _16362_ (.Y(_07267_),
    .A(_07264_),
    .B(_07236_));
 sg13g2_inv_1 _16363_ (.Y(_07268_),
    .A(net178));
 sg13g2_nand3_1 _16364_ (.B(net57),
    .C(_07268_),
    .A(_07267_),
    .Y(_07269_));
 sg13g2_nand2_1 _16365_ (.Y(_07270_),
    .A(_07266_),
    .B(_07269_));
 sg13g2_xnor2_1 _16366_ (.Y(_07271_),
    .A(_04705_),
    .B(_04791_));
 sg13g2_nand2_1 _16367_ (.Y(_07272_),
    .A(_07270_),
    .B(_07271_));
 sg13g2_inv_1 _16368_ (.Y(_07273_),
    .A(_04708_));
 sg13g2_nor3_1 _16369_ (.A(_04705_),
    .B(_04707_),
    .C(_07273_),
    .Y(_07274_));
 sg13g2_nand2_1 _16370_ (.Y(_07275_),
    .A(_04717_),
    .B(_07274_));
 sg13g2_a21oi_1 _16371_ (.A1(_07253_),
    .A2(_07172_),
    .Y(_07276_),
    .B1(_07275_));
 sg13g2_nand3_1 _16372_ (.B(_07273_),
    .C(_04707_),
    .A(_04706_),
    .Y(_07277_));
 sg13g2_nor2_1 _16373_ (.A(_07254_),
    .B(_07245_),
    .Y(_07278_));
 sg13g2_nand2_1 _16374_ (.Y(_07279_),
    .A(_07278_),
    .B(_07260_));
 sg13g2_o21ai_1 _16375_ (.B1(net178),
    .Y(_07280_),
    .A1(_07234_),
    .A2(_07279_));
 sg13g2_nor2_1 _16376_ (.A(_07277_),
    .B(_07280_),
    .Y(_07281_));
 sg13g2_inv_1 _16377_ (.Y(_07282_),
    .A(_04715_));
 sg13g2_nor2_1 _16378_ (.A(net63),
    .B(_07282_),
    .Y(_07283_));
 sg13g2_o21ai_1 _16379_ (.B1(_07283_),
    .Y(_07284_),
    .A1(_07276_),
    .A2(_07281_));
 sg13g2_nand3_1 _16380_ (.B(_07155_),
    .C(_05746_),
    .A(_04789_),
    .Y(_07285_));
 sg13g2_o21ai_1 _16381_ (.B1(net178),
    .Y(_07286_),
    .A1(_07285_),
    .A2(_07129_));
 sg13g2_nor2b_1 _16382_ (.A(_07286_),
    .B_N(_04792_),
    .Y(_07287_));
 sg13g2_nand2_1 _16383_ (.Y(_07288_),
    .A(_04791_),
    .B(_04705_));
 sg13g2_a21oi_1 _16384_ (.A1(_07280_),
    .A2(_07286_),
    .Y(_07289_),
    .B1(_07288_));
 sg13g2_o21ai_1 _16385_ (.B1(_07283_),
    .Y(_07290_),
    .A1(_07287_),
    .A2(_07289_));
 sg13g2_nand3_1 _16386_ (.B(_07284_),
    .C(_07290_),
    .A(_07272_),
    .Y(_07291_));
 sg13g2_buf_1 _16387_ (.A(\b.gen_square[53].sq.mask ),
    .X(_07292_));
 sg13g2_nand2_1 _16388_ (.Y(_07293_),
    .A(_07291_),
    .B(_07292_));
 sg13g2_nand2_1 _16389_ (.Y(_07294_),
    .A(_07070_),
    .B(_07293_));
 sg13g2_xnor2_1 _16390_ (.Y(_07295_),
    .A(_05031_),
    .B(_05097_));
 sg13g2_inv_1 _16391_ (.Y(_07296_),
    .A(_05034_));
 sg13g2_nand3_1 _16392_ (.B(_07296_),
    .C(_05033_),
    .A(_05032_),
    .Y(_07297_));
 sg13g2_or2_1 _16393_ (.X(_07298_),
    .B(_05104_),
    .A(_07297_));
 sg13g2_nand2b_1 _16394_ (.Y(_07299_),
    .B(_05021_),
    .A_N(_04586_));
 sg13g2_nand4_1 _16395_ (.B(_05032_),
    .C(_05038_),
    .A(net180),
    .Y(_07300_),
    .D(_05034_));
 sg13g2_inv_1 _16396_ (.Y(_07301_),
    .A(_07300_));
 sg13g2_nand2_1 _16397_ (.Y(_07302_),
    .A(_07299_),
    .B(_07301_));
 sg13g2_a21oi_1 _16398_ (.A1(_07298_),
    .A2(_07302_),
    .Y(_07303_),
    .B1(_05117_));
 sg13g2_a21oi_1 _16399_ (.A1(_05095_),
    .A2(_07295_),
    .Y(_07304_),
    .B1(_07303_));
 sg13g2_nand2_1 _16400_ (.Y(_07305_),
    .A(_07304_),
    .B(_05118_));
 sg13g2_nand2_1 _16401_ (.Y(_07306_),
    .A(_07305_),
    .B(_05120_));
 sg13g2_nand2_1 _16402_ (.Y(_07307_),
    .A(_07266_),
    .B(_04710_));
 sg13g2_nand2b_1 _16403_ (.Y(_07308_),
    .B(_04709_),
    .A_N(_04791_));
 sg13g2_nand3_1 _16404_ (.B(_07307_),
    .C(_07308_),
    .A(_07270_),
    .Y(_07309_));
 sg13g2_nand2_1 _16405_ (.Y(_07310_),
    .A(_07309_),
    .B(_07290_));
 sg13g2_nand2_1 _16406_ (.Y(_07311_),
    .A(_07310_),
    .B(_07292_));
 sg13g2_inv_1 _16407_ (.Y(_07312_),
    .A(_07311_));
 sg13g2_nand2_1 _16408_ (.Y(_07313_),
    .A(_07048_),
    .B(_04686_));
 sg13g2_nand2b_1 _16409_ (.Y(_07314_),
    .B(_04685_),
    .A_N(_04782_));
 sg13g2_nand3_1 _16410_ (.B(_07313_),
    .C(_07314_),
    .A(_07049_),
    .Y(_07315_));
 sg13g2_a21o_1 _16411_ (.A2(_07066_),
    .A1(_07315_),
    .B1(_07067_),
    .X(_07316_));
 sg13g2_inv_1 _16412_ (.Y(_07317_),
    .A(_07316_));
 sg13g2_nor2_1 _16413_ (.A(_04749_),
    .B(_04747_),
    .Y(_07318_));
 sg13g2_a21oi_1 _16414_ (.A1(_05796_),
    .A2(_04614_),
    .Y(_07319_),
    .B1(_07318_));
 sg13g2_a22oi_1 _16415_ (.Y(_07320_),
    .B1(_05799_),
    .B2(_07319_),
    .A2(net95),
    .A1(_05805_));
 sg13g2_nand2b_1 _16416_ (.Y(_07321_),
    .B(_05808_),
    .A_N(_07320_));
 sg13g2_inv_1 _16417_ (.Y(_07322_),
    .A(_07321_));
 sg13g2_nand2_1 _16418_ (.Y(_07323_),
    .A(_06136_),
    .B(_04594_));
 sg13g2_nand2b_1 _16419_ (.Y(_07324_),
    .B(_04593_),
    .A_N(_04735_));
 sg13g2_nand3_1 _16420_ (.B(_07323_),
    .C(_07324_),
    .A(_06139_),
    .Y(_07325_));
 sg13g2_inv_1 _16421_ (.Y(_07326_),
    .A(_06147_));
 sg13g2_a21o_1 _16422_ (.A2(_07325_),
    .A1(_06145_),
    .B1(_07326_),
    .X(_07327_));
 sg13g2_buf_1 _16423_ (.A(_07327_),
    .X(_07328_));
 sg13g2_nor2_1 _16424_ (.A(_07328_),
    .B(_07322_),
    .Y(_07329_));
 sg13g2_nand3b_1 _16425_ (.B(_05804_),
    .C(_05421_),
    .Y(_07330_),
    .A_N(_04619_));
 sg13g2_inv_1 _16426_ (.Y(_07331_),
    .A(_05773_));
 sg13g2_and2_1 _16427_ (.A(_05506_),
    .B(_05443_),
    .X(_07332_));
 sg13g2_nand4_1 _16428_ (.B(_04619_),
    .C(_05469_),
    .A(_07332_),
    .Y(_07333_),
    .D(_05510_));
 sg13g2_nor2_1 _16429_ (.A(_05492_),
    .B(_07333_),
    .Y(_07334_));
 sg13g2_nand4_1 _16430_ (.B(_05440_),
    .C(_05574_),
    .A(_07331_),
    .Y(_07335_),
    .D(_07334_));
 sg13g2_nand4_1 _16431_ (.B(net95),
    .C(_04743_),
    .A(_07330_),
    .Y(_07336_),
    .D(_07335_));
 sg13g2_o21ai_1 _16432_ (.B1(_04615_),
    .Y(_07337_),
    .A1(_04612_),
    .A2(_05124_));
 sg13g2_nand3_1 _16433_ (.B(net86),
    .C(_07337_),
    .A(_05797_),
    .Y(_07338_));
 sg13g2_nand3_1 _16434_ (.B(net145),
    .C(_04617_),
    .A(_05795_),
    .Y(_07339_));
 sg13g2_nand3_1 _16435_ (.B(_07338_),
    .C(_07339_),
    .A(_07336_),
    .Y(_07340_));
 sg13g2_nand2_1 _16436_ (.Y(_07341_),
    .A(_07340_),
    .B(_05808_));
 sg13g2_inv_1 _16437_ (.Y(_07342_),
    .A(_06148_));
 sg13g2_nor2_1 _16438_ (.A(_05809_),
    .B(_07342_),
    .Y(_07343_));
 sg13g2_a21oi_1 _16439_ (.A1(_07322_),
    .A2(_07328_),
    .Y(_07344_),
    .B1(_07343_));
 sg13g2_o21ai_1 _16440_ (.B1(_07344_),
    .Y(_07345_),
    .A1(_07329_),
    .A2(_07341_));
 sg13g2_nand3_1 _16441_ (.B(_04598_),
    .C(_05936_),
    .A(_06143_),
    .Y(_07346_));
 sg13g2_o21ai_1 _16442_ (.B1(_04600_),
    .Y(_07347_),
    .A1(_05947_),
    .A2(_06126_));
 sg13g2_nand2_1 _16443_ (.Y(_07348_),
    .A(_07347_),
    .B(_05504_));
 sg13g2_nand3_1 _16444_ (.B(net95),
    .C(_07348_),
    .A(_07346_),
    .Y(_07349_));
 sg13g2_nand2_1 _16445_ (.Y(_07350_),
    .A(_04595_),
    .B(_04600_));
 sg13g2_nand3_1 _16446_ (.B(net96),
    .C(_07350_),
    .A(_06137_),
    .Y(_07351_));
 sg13g2_a21o_1 _16447_ (.A2(_04595_),
    .A1(_04592_),
    .B1(_07351_),
    .X(_07352_));
 sg13g2_nand3_1 _16448_ (.B(net145),
    .C(_05835_),
    .A(_06135_),
    .Y(_07353_));
 sg13g2_nand3_1 _16449_ (.B(_07352_),
    .C(_07353_),
    .A(_07349_),
    .Y(_07354_));
 sg13g2_nand2_1 _16450_ (.Y(_07355_),
    .A(_07354_),
    .B(_06147_));
 sg13g2_inv_1 _16451_ (.Y(_07356_),
    .A(_07355_));
 sg13g2_nand2_1 _16452_ (.Y(_07357_),
    .A(_07344_),
    .B(_07356_));
 sg13g2_nand2_1 _16453_ (.Y(_07358_),
    .A(_07342_),
    .B(_05809_));
 sg13g2_nand3_1 _16454_ (.B(_07357_),
    .C(_07358_),
    .A(_07345_),
    .Y(_07359_));
 sg13g2_buf_2 _16455_ (.A(_07359_),
    .X(_07360_));
 sg13g2_nand2_1 _16456_ (.Y(_07361_),
    .A(_07360_),
    .B(_07328_));
 sg13g2_o21ai_1 _16457_ (.B1(_07361_),
    .Y(_07362_),
    .A1(_07322_),
    .A2(_07360_));
 sg13g2_buf_1 _16458_ (.A(_07362_),
    .X(_07363_));
 sg13g2_nand2_1 _16459_ (.Y(_07364_),
    .A(_06479_),
    .B(_04637_));
 sg13g2_nand2b_1 _16460_ (.Y(_07365_),
    .B(_04636_),
    .A_N(_04760_));
 sg13g2_nand3_1 _16461_ (.B(_07364_),
    .C(_07365_),
    .A(_06480_),
    .Y(_07366_));
 sg13g2_a21o_1 _16462_ (.A2(_06498_),
    .A1(_07366_),
    .B1(_06499_),
    .X(_07367_));
 sg13g2_inv_1 _16463_ (.Y(_07368_),
    .A(_07367_));
 sg13g2_nor2_1 _16464_ (.A(_07368_),
    .B(_07363_),
    .Y(_07369_));
 sg13g2_nand2_1 _16465_ (.Y(_07370_),
    .A(_07360_),
    .B(_07356_));
 sg13g2_o21ai_1 _16466_ (.B1(_07370_),
    .Y(_07371_),
    .A1(_07341_),
    .A2(_07360_));
 sg13g2_nand3_1 _16467_ (.B(_04641_),
    .C(_06485_),
    .A(_06496_),
    .Y(_07372_));
 sg13g2_inv_1 _16468_ (.Y(_07373_),
    .A(_05484_));
 sg13g2_nor2_1 _16469_ (.A(_07373_),
    .B(_06264_),
    .Y(_07374_));
 sg13g2_nand3_1 _16470_ (.B(_05946_),
    .C(_05469_),
    .A(_07374_),
    .Y(_07375_));
 sg13g2_nand2_1 _16471_ (.Y(_07376_),
    .A(_06311_),
    .B(_05562_));
 sg13g2_nor3_1 _16472_ (.A(_07375_),
    .B(_07376_),
    .C(_06252_),
    .Y(_07377_));
 sg13g2_nand3_1 _16473_ (.B(_06456_),
    .C(_05541_),
    .A(_07377_),
    .Y(_07378_));
 sg13g2_nor2_1 _16474_ (.A(net83),
    .B(_04645_),
    .Y(_07379_));
 sg13g2_nand3_1 _16475_ (.B(_07378_),
    .C(_07379_),
    .A(_07372_),
    .Y(_07380_));
 sg13g2_buf_1 _16476_ (.A(_04261_),
    .X(_07381_));
 sg13g2_a21oi_1 _16477_ (.A1(_04757_),
    .A2(_06486_),
    .Y(_07382_),
    .B1(_04637_));
 sg13g2_nor3_1 _16478_ (.A(net158),
    .B(_07382_),
    .C(_06475_),
    .Y(_07383_));
 sg13g2_nor2_1 _16479_ (.A(_04635_),
    .B(_06479_),
    .Y(_07384_));
 sg13g2_nor2_1 _16480_ (.A(_07383_),
    .B(_07384_),
    .Y(_07385_));
 sg13g2_a21oi_1 _16481_ (.A1(_07380_),
    .A2(_07385_),
    .Y(_07386_),
    .B1(_06499_));
 sg13g2_nand2b_1 _16482_ (.Y(_07387_),
    .B(_07386_),
    .A_N(_07371_));
 sg13g2_nor2_1 _16483_ (.A(_06149_),
    .B(_06501_),
    .Y(_07388_));
 sg13g2_a21oi_1 _16484_ (.A1(_07363_),
    .A2(_07368_),
    .Y(_07389_),
    .B1(_07388_));
 sg13g2_o21ai_1 _16485_ (.B1(_07389_),
    .Y(_07390_),
    .A1(_07369_),
    .A2(_07387_));
 sg13g2_nand2_1 _16486_ (.Y(_07391_),
    .A(_06501_),
    .B(_06149_));
 sg13g2_nand2_1 _16487_ (.Y(_07392_),
    .A(_07390_),
    .B(_07391_));
 sg13g2_buf_1 _16488_ (.A(_07392_),
    .X(_07393_));
 sg13g2_nor2_1 _16489_ (.A(_07368_),
    .B(_07393_),
    .Y(_07394_));
 sg13g2_a21oi_1 _16490_ (.A1(_07363_),
    .A2(_07393_),
    .Y(_07395_),
    .B1(_07394_));
 sg13g2_inv_1 _16491_ (.Y(_07396_),
    .A(_06502_));
 sg13g2_nand2_1 _16492_ (.Y(_07397_),
    .A(_06847_),
    .B(_04662_));
 sg13g2_nand2b_1 _16493_ (.Y(_07398_),
    .B(_04661_),
    .A_N(_04771_));
 sg13g2_nand3_1 _16494_ (.B(_07397_),
    .C(_07398_),
    .A(_06848_),
    .Y(_07399_));
 sg13g2_o21ai_1 _16495_ (.B1(net75),
    .Y(_07400_),
    .A1(_06614_),
    .A2(_06780_));
 sg13g2_inv_1 _16496_ (.Y(_07401_),
    .A(_06852_));
 sg13g2_a21o_1 _16497_ (.A2(_07400_),
    .A1(_07399_),
    .B1(_07401_),
    .X(_07402_));
 sg13g2_buf_1 _16498_ (.A(_07402_),
    .X(_07403_));
 sg13g2_mux2_1 _16499_ (.A0(_07386_),
    .A1(_07371_),
    .S(_07393_),
    .X(_07404_));
 sg13g2_inv_1 _16500_ (.Y(_07405_),
    .A(_06257_));
 sg13g2_nor4_1 _16501_ (.A(_07405_),
    .B(_07373_),
    .C(_07036_),
    .D(_05546_),
    .Y(_07406_));
 sg13g2_nor2b_1 _16502_ (.A(_06835_),
    .B_N(_05424_),
    .Y(_07407_));
 sg13g2_nand4_1 _16503_ (.B(_06826_),
    .C(_07406_),
    .A(_06832_),
    .Y(_07408_),
    .D(_07407_));
 sg13g2_o21ai_1 _16504_ (.B1(net75),
    .Y(_07409_),
    .A1(_04668_),
    .A2(_07408_));
 sg13g2_nor3_1 _16505_ (.A(_04667_),
    .B(_06779_),
    .C(_06780_),
    .Y(_07410_));
 sg13g2_nor3_1 _16506_ (.A(_04669_),
    .B(_07409_),
    .C(_07410_),
    .Y(_07411_));
 sg13g2_buf_1 _16507_ (.A(net158),
    .X(_07412_));
 sg13g2_a21oi_1 _16508_ (.A1(_04768_),
    .A2(_04666_),
    .Y(_07413_),
    .B1(_04662_));
 sg13g2_nor3_1 _16509_ (.A(net142),
    .B(_07413_),
    .C(_06843_),
    .Y(_07414_));
 sg13g2_nor2_1 _16510_ (.A(_04660_),
    .B(_06847_),
    .Y(_07415_));
 sg13g2_nor3_1 _16511_ (.A(_07411_),
    .B(_07414_),
    .C(_07415_),
    .Y(_07416_));
 sg13g2_nor2_1 _16512_ (.A(_07401_),
    .B(_07416_),
    .Y(_07417_));
 sg13g2_nand2b_1 _16513_ (.Y(_07418_),
    .B(_07417_),
    .A_N(_07404_));
 sg13g2_o21ai_1 _16514_ (.B1(_07418_),
    .Y(_07419_),
    .A1(_07403_),
    .A2(_07395_));
 sg13g2_nand2b_1 _16515_ (.Y(_07420_),
    .B(_06853_),
    .A_N(_06502_));
 sg13g2_nand2_1 _16516_ (.Y(_07421_),
    .A(_07395_),
    .B(_07403_));
 sg13g2_nand3_1 _16517_ (.B(_07420_),
    .C(_07421_),
    .A(_07419_),
    .Y(_07422_));
 sg13g2_o21ai_1 _16518_ (.B1(_07422_),
    .Y(_07423_),
    .A1(_07396_),
    .A2(_06853_));
 sg13g2_buf_1 _16519_ (.A(_07423_),
    .X(_07424_));
 sg13g2_nand2_1 _16520_ (.Y(_07425_),
    .A(_07424_),
    .B(_07403_));
 sg13g2_o21ai_1 _16521_ (.B1(_07425_),
    .Y(_07426_),
    .A1(_07395_),
    .A2(_07424_));
 sg13g2_nor2_1 _16522_ (.A(_07317_),
    .B(_07426_),
    .Y(_07427_));
 sg13g2_mux2_1 _16523_ (.A0(_07404_),
    .A1(_07417_),
    .S(_07424_),
    .X(_07428_));
 sg13g2_a21oi_1 _16524_ (.A1(_04779_),
    .A2(_04690_),
    .Y(_07429_),
    .B1(_04686_));
 sg13g2_nor3_1 _16525_ (.A(net142),
    .B(_07429_),
    .C(_07045_),
    .Y(_07430_));
 sg13g2_nor2_1 _16526_ (.A(_04684_),
    .B(_07048_),
    .Y(_07431_));
 sg13g2_nor2_1 _16527_ (.A(_07430_),
    .B(_07431_),
    .Y(_07432_));
 sg13g2_nand3_1 _16528_ (.B(_04692_),
    .C(_07054_),
    .A(_07064_),
    .Y(_07433_));
 sg13g2_inv_1 _16529_ (.Y(_07434_),
    .A(_04693_));
 sg13g2_nand4_1 _16530_ (.B(_04691_),
    .C(_06257_),
    .A(_07034_),
    .Y(_07435_),
    .D(_06787_));
 sg13g2_nor3_1 _16531_ (.A(_06250_),
    .B(_07435_),
    .C(_07024_),
    .Y(_07436_));
 sg13g2_nand4_1 _16532_ (.B(_06896_),
    .C(_07018_),
    .A(_07436_),
    .Y(_07437_),
    .D(_07026_));
 sg13g2_nand4_1 _16533_ (.B(net67),
    .C(_07434_),
    .A(_07433_),
    .Y(_07438_),
    .D(_07437_));
 sg13g2_a21oi_1 _16534_ (.A1(_07432_),
    .A2(_07438_),
    .Y(_07439_),
    .B1(_07067_));
 sg13g2_nand2b_1 _16535_ (.Y(_07440_),
    .B(_07439_),
    .A_N(_07428_));
 sg13g2_nor2_1 _16536_ (.A(_07069_),
    .B(_06854_),
    .Y(_07441_));
 sg13g2_a21oi_1 _16537_ (.A1(_07426_),
    .A2(_07317_),
    .Y(_07442_),
    .B1(_07441_));
 sg13g2_o21ai_1 _16538_ (.B1(_07442_),
    .Y(_07443_),
    .A1(_07427_),
    .A2(_07440_));
 sg13g2_nand2_1 _16539_ (.Y(_07444_),
    .A(_06854_),
    .B(_07069_));
 sg13g2_nand2_1 _16540_ (.Y(_07445_),
    .A(_07443_),
    .B(_07444_));
 sg13g2_nand2_1 _16541_ (.Y(_07446_),
    .A(_07445_),
    .B(_07426_));
 sg13g2_o21ai_1 _16542_ (.B1(_07446_),
    .Y(_07447_),
    .A1(_07317_),
    .A2(_07445_));
 sg13g2_nand2_1 _16543_ (.Y(_07448_),
    .A(_07268_),
    .B(_07273_));
 sg13g2_a21oi_1 _16544_ (.A1(_07448_),
    .A2(_04711_),
    .Y(_07449_),
    .B1(net142));
 sg13g2_nand3_1 _16545_ (.B(_07175_),
    .C(_07176_),
    .A(_07151_),
    .Y(_07450_));
 sg13g2_nor2_1 _16546_ (.A(_04467_),
    .B(_06825_),
    .Y(_07451_));
 sg13g2_nand4_1 _16547_ (.B(_07242_),
    .C(_07256_),
    .A(_07243_),
    .Y(_07452_),
    .D(_07451_));
 sg13g2_o21ai_1 _16548_ (.B1(net178),
    .Y(_07453_),
    .A1(_07450_),
    .A2(_07452_));
 sg13g2_nor3_1 _16549_ (.A(_07282_),
    .B(_07281_),
    .C(_07289_),
    .Y(_07454_));
 sg13g2_a21oi_1 _16550_ (.A1(_07282_),
    .A2(_07453_),
    .Y(_07455_),
    .B1(_07454_));
 sg13g2_a22oi_1 _16551_ (.Y(_07456_),
    .B1(net56),
    .B2(_07455_),
    .A2(_07449_),
    .A1(_07267_));
 sg13g2_o21ai_1 _16552_ (.B1(_07456_),
    .Y(_07457_),
    .A1(_04708_),
    .A2(_07266_));
 sg13g2_nand2_1 _16553_ (.Y(_07458_),
    .A(_07457_),
    .B(_07292_));
 sg13g2_mux2_1 _16554_ (.A0(_07439_),
    .A1(_07428_),
    .S(_07445_),
    .X(_07459_));
 sg13g2_nor2_1 _16555_ (.A(_07458_),
    .B(_07459_),
    .Y(_07460_));
 sg13g2_o21ai_1 _16556_ (.B1(_07460_),
    .Y(_07461_),
    .A1(_07447_),
    .A2(_07312_));
 sg13g2_nand2b_1 _16557_ (.Y(_07462_),
    .B(_07293_),
    .A_N(_07070_));
 sg13g2_nand2b_1 _16558_ (.Y(_07463_),
    .B(_07070_),
    .A_N(_07293_));
 sg13g2_nand2_1 _16559_ (.Y(_07464_),
    .A(_07447_),
    .B(_07312_));
 sg13g2_nand4_1 _16560_ (.B(_07462_),
    .C(_07463_),
    .A(_07461_),
    .Y(_07465_),
    .D(_07464_));
 sg13g2_nand2_2 _16561_ (.Y(_07466_),
    .A(_07465_),
    .B(_07462_));
 sg13g2_nand2_1 _16562_ (.Y(_07467_),
    .A(_07466_),
    .B(_07447_));
 sg13g2_o21ai_1 _16563_ (.B1(_07467_),
    .Y(_07468_),
    .A1(_07312_),
    .A2(_07466_));
 sg13g2_nor2_1 _16564_ (.A(_07306_),
    .B(_07294_),
    .Y(_07469_));
 sg13g2_a21oi_1 _16565_ (.A1(_07468_),
    .A2(_05122_),
    .Y(_07470_),
    .B1(_07469_));
 sg13g2_nand3_1 _16566_ (.B(_05040_),
    .C(_07298_),
    .A(_05106_),
    .Y(_07471_));
 sg13g2_nor3_1 _16567_ (.A(_05040_),
    .B(_05012_),
    .C(_04469_),
    .Y(_07472_));
 sg13g2_nand4_1 _16568_ (.B(_07472_),
    .C(_07023_),
    .A(_05069_),
    .Y(_07473_),
    .D(_05000_));
 sg13g2_nor2_1 _16569_ (.A(net48),
    .B(_05041_),
    .Y(_07474_));
 sg13g2_nand3_1 _16570_ (.B(_07473_),
    .C(_07474_),
    .A(_07471_),
    .Y(_07475_));
 sg13g2_nand3_1 _16571_ (.B(net97),
    .C(_07296_),
    .A(_05071_),
    .Y(_07476_));
 sg13g2_o21ai_1 _16572_ (.B1(_05037_),
    .Y(_07477_),
    .A1(_05034_),
    .A2(_04038_));
 sg13g2_nand3_1 _16573_ (.B(net41),
    .C(_07477_),
    .A(_05081_),
    .Y(_07478_));
 sg13g2_nand3_1 _16574_ (.B(_07476_),
    .C(_07478_),
    .A(_07475_),
    .Y(_07479_));
 sg13g2_nand2_1 _16575_ (.Y(_07480_),
    .A(_07479_),
    .B(_05120_));
 sg13g2_nand2_1 _16576_ (.Y(_07481_),
    .A(_07466_),
    .B(_07459_));
 sg13g2_o21ai_1 _16577_ (.B1(_07481_),
    .Y(_07482_),
    .A1(_07458_),
    .A2(_07466_));
 sg13g2_nor2_1 _16578_ (.A(_07480_),
    .B(_07482_),
    .Y(_07483_));
 sg13g2_o21ai_1 _16579_ (.B1(_07483_),
    .Y(_07484_),
    .A1(_05122_),
    .A2(_07468_));
 sg13g2_a22oi_1 _16580_ (.Y(_07485_),
    .B1(_07470_),
    .B2(_07484_),
    .A2(_07306_),
    .A1(_07294_));
 sg13g2_buf_2 _16581_ (.A(_07485_),
    .X(_07486_));
 sg13g2_nor2_1 _16582_ (.A(_07468_),
    .B(_07486_),
    .Y(_07487_));
 sg13g2_a21oi_1 _16583_ (.A1(_05122_),
    .A2(_07486_),
    .Y(_07488_),
    .B1(_07487_));
 sg13g2_o21ai_1 _16584_ (.B1(_06167_),
    .Y(_07489_),
    .A1(_06165_),
    .A2(_05522_));
 sg13g2_buf_1 _16585_ (.A(_07489_),
    .X(_07490_));
 sg13g2_inv_1 _16586_ (.Y(_07491_),
    .A(_06724_));
 sg13g2_inv_1 _16587_ (.Y(_07492_),
    .A(_06727_));
 sg13g2_a21oi_2 _16588_ (.B1(_07492_),
    .Y(_07493_),
    .A2(_07491_),
    .A1(_07490_));
 sg13g2_inv_1 _16589_ (.Y(_07494_),
    .A(_04096_));
 sg13g2_inv_1 _16590_ (.Y(_07495_),
    .A(_00017_));
 sg13g2_nor2_1 _16591_ (.A(_07495_),
    .B(_07494_),
    .Y(_07496_));
 sg13g2_a21oi_2 _16592_ (.B1(_07496_),
    .Y(_07497_),
    .A2(_07494_),
    .A1(_07493_));
 sg13g2_inv_1 _16593_ (.Y(_07498_),
    .A(_07497_));
 sg13g2_inv_1 _16594_ (.Y(_07499_),
    .A(_04983_));
 sg13g2_nor2_1 _16595_ (.A(_04568_),
    .B(_07499_),
    .Y(_07500_));
 sg13g2_a21oi_1 _16596_ (.A1(_07498_),
    .A2(_07499_),
    .Y(_07501_),
    .B1(_07500_));
 sg13g2_inv_1 _16597_ (.Y(_07502_),
    .A(_07501_));
 sg13g2_nor2_1 _16598_ (.A(_07249_),
    .B(_04406_),
    .Y(_07503_));
 sg13g2_a21oi_1 _16599_ (.A1(_07502_),
    .A2(_04406_),
    .Y(_07504_),
    .B1(_07503_));
 sg13g2_inv_1 _16600_ (.Y(_07505_),
    .A(_06165_));
 sg13g2_inv_1 _16601_ (.Y(_07506_),
    .A(_05517_));
 sg13g2_a21oi_1 _16602_ (.A1(_05296_),
    .A2(_07506_),
    .Y(_07507_),
    .B1(_05299_));
 sg13g2_nor2_1 _16603_ (.A(_07507_),
    .B(_05303_),
    .Y(_07508_));
 sg13g2_nor2_2 _16604_ (.A(_05309_),
    .B(_07508_),
    .Y(_07509_));
 sg13g2_nor2_1 _16605_ (.A(_06153_),
    .B(_06162_),
    .Y(_07510_));
 sg13g2_a21oi_1 _16606_ (.A1(_06153_),
    .A2(_06206_),
    .Y(_07511_),
    .B1(_07510_));
 sg13g2_nor2_1 _16607_ (.A(_07511_),
    .B(_06209_),
    .Y(_07512_));
 sg13g2_nor2_1 _16608_ (.A(_07512_),
    .B(_06211_),
    .Y(_07513_));
 sg13g2_inv_1 _16609_ (.Y(_07514_),
    .A(_07513_));
 sg13g2_nor2_1 _16610_ (.A(_07505_),
    .B(_07514_),
    .Y(_07515_));
 sg13g2_a21oi_1 _16611_ (.A1(_07505_),
    .A2(_07509_),
    .Y(_07516_),
    .B1(_07515_));
 sg13g2_nor2_1 _16612_ (.A(_06668_),
    .B(_06721_),
    .Y(_07517_));
 sg13g2_nand2b_1 _16613_ (.Y(_07518_),
    .B(_06669_),
    .A_N(_07517_));
 sg13g2_inv_1 _16614_ (.Y(_07519_),
    .A(_06664_));
 sg13g2_nor2_1 _16615_ (.A(_07519_),
    .B(net80),
    .Y(_07520_));
 sg13g2_a21oi_1 _16616_ (.A1(_07518_),
    .A2(_07520_),
    .Y(_07521_),
    .B1(_06681_));
 sg13g2_inv_1 _16617_ (.Y(_07522_),
    .A(_07521_));
 sg13g2_nor2_1 _16618_ (.A(_06722_),
    .B(_07522_),
    .Y(_07523_));
 sg13g2_inv_1 _16619_ (.Y(_07524_),
    .A(_07523_));
 sg13g2_o21ai_1 _16620_ (.B1(_07524_),
    .Y(_07525_),
    .A1(_06724_),
    .A2(_07516_));
 sg13g2_inv_1 _16621_ (.Y(_07526_),
    .A(_04092_));
 sg13g2_nor2_1 _16622_ (.A(_06855_),
    .B(_04300_),
    .Y(_07527_));
 sg13g2_nand3_1 _16623_ (.B(_04070_),
    .C(_04073_),
    .A(_04093_),
    .Y(_07528_));
 sg13g2_nand2_1 _16624_ (.Y(_07529_),
    .A(_07528_),
    .B(_06857_));
 sg13g2_nand2_1 _16625_ (.Y(_07530_),
    .A(_07527_),
    .B(_07529_));
 sg13g2_nor2b_1 _16626_ (.A(_07526_),
    .B_N(_07530_),
    .Y(_07531_));
 sg13g2_inv_1 _16627_ (.Y(_07532_),
    .A(_07531_));
 sg13g2_nor2_1 _16628_ (.A(_04095_),
    .B(_07532_),
    .Y(_07533_));
 sg13g2_a21oi_1 _16629_ (.A1(_07525_),
    .A2(_07494_),
    .Y(_07534_),
    .B1(_07533_));
 sg13g2_inv_2 _16630_ (.Y(_07535_),
    .A(_04570_));
 sg13g2_inv_1 _16631_ (.Y(_07536_),
    .A(_04981_));
 sg13g2_a21oi_1 _16632_ (.A1(_04980_),
    .A2(_07536_),
    .Y(_07537_),
    .B1(_07220_));
 sg13g2_nor3_1 _16633_ (.A(net61),
    .B(_07535_),
    .C(_07537_),
    .Y(_07538_));
 sg13g2_nor2_1 _16634_ (.A(_07538_),
    .B(_04583_),
    .Y(_07539_));
 sg13g2_inv_1 _16635_ (.Y(_07540_),
    .A(_07539_));
 sg13g2_nor2_1 _16636_ (.A(_04982_),
    .B(_07540_),
    .Y(_07541_));
 sg13g2_inv_1 _16637_ (.Y(_07542_),
    .A(_07541_));
 sg13g2_o21ai_1 _16638_ (.B1(_07542_),
    .Y(_07543_),
    .A1(_04983_),
    .A2(_07534_));
 sg13g2_nor2_1 _16639_ (.A(_04385_),
    .B(_04402_),
    .Y(_07544_));
 sg13g2_nor2_1 _16640_ (.A(_07544_),
    .B(_04483_),
    .Y(_07545_));
 sg13g2_nor3_1 _16641_ (.A(_04392_),
    .B(net61),
    .C(_07545_),
    .Y(_07546_));
 sg13g2_nor2_1 _16642_ (.A(_07546_),
    .B(_04399_),
    .Y(_07547_));
 sg13g2_inv_1 _16643_ (.Y(_07548_),
    .A(_07547_));
 sg13g2_nor2_1 _16644_ (.A(_04403_),
    .B(_07548_),
    .Y(_07549_));
 sg13g2_a21oi_1 _16645_ (.A1(_07543_),
    .A2(_04406_),
    .Y(_07550_),
    .B1(_07549_));
 sg13g2_inv_1 _16646_ (.Y(_07551_),
    .A(_07550_));
 sg13g2_nor2_1 _16647_ (.A(_04423_),
    .B(_04427_),
    .Y(_07552_));
 sg13g2_inv_1 _16648_ (.Y(_07553_),
    .A(_07552_));
 sg13g2_nor2_1 _16649_ (.A(_04370_),
    .B(_07553_),
    .Y(_07554_));
 sg13g2_inv_1 _16650_ (.Y(_07555_),
    .A(_04501_));
 sg13g2_o21ai_1 _16651_ (.B1(_07555_),
    .Y(_07556_),
    .A1(_04412_),
    .A2(_04422_));
 sg13g2_a21oi_2 _16652_ (.B1(_04429_),
    .Y(_07557_),
    .A2(_07556_),
    .A1(_07554_));
 sg13g2_inv_1 _16653_ (.Y(_07558_),
    .A(_04426_));
 sg13g2_nor2_1 _16654_ (.A(_07557_),
    .B(_07558_),
    .Y(_07559_));
 sg13g2_a21oi_1 _16655_ (.A1(_04730_),
    .A2(net84),
    .Y(_07560_),
    .B1(_05728_));
 sg13g2_inv_1 _16656_ (.Y(_07561_),
    .A(_04797_));
 sg13g2_a21oi_1 _16657_ (.A1(_07561_),
    .A2(net84),
    .Y(_07562_),
    .B1(_05744_));
 sg13g2_nand2b_1 _16658_ (.Y(_07563_),
    .B(_07562_),
    .A_N(_07560_));
 sg13g2_nor2b_1 _16659_ (.A(_07559_),
    .B_N(_07563_),
    .Y(_07564_));
 sg13g2_o21ai_1 _16660_ (.B1(_07564_),
    .Y(_07565_),
    .A1(_07504_),
    .A2(_07551_));
 sg13g2_inv_1 _16661_ (.Y(_07566_),
    .A(_07565_));
 sg13g2_o21ai_1 _16662_ (.B1(_05058_),
    .Y(_07567_),
    .A1(_04438_),
    .A2(_04426_));
 sg13g2_buf_1 _16663_ (.A(_07567_),
    .X(_07568_));
 sg13g2_inv_1 _16664_ (.Y(_07569_),
    .A(_07568_));
 sg13g2_a21oi_1 _16665_ (.A1(_07569_),
    .A2(_04406_),
    .Y(_07570_),
    .B1(_07503_));
 sg13g2_nor2_1 _16666_ (.A(_04401_),
    .B(_07570_),
    .Y(_07571_));
 sg13g2_nor3_1 _16667_ (.A(_06625_),
    .B(_07246_),
    .C(_06635_),
    .Y(_07572_));
 sg13g2_nand3_1 _16668_ (.B(_04432_),
    .C(_07255_),
    .A(_07572_),
    .Y(_07573_));
 sg13g2_inv_1 _16669_ (.Y(_07574_),
    .A(net55));
 sg13g2_and3_1 _16670_ (.X(_07575_),
    .A(_05596_),
    .B(_05607_),
    .C(_05592_));
 sg13g2_nor2_1 _16671_ (.A(_05599_),
    .B(_07575_),
    .Y(_07576_));
 sg13g2_o21ai_1 _16672_ (.B1(_05610_),
    .Y(_07577_),
    .A1(_05605_),
    .A2(_07576_));
 sg13g2_inv_1 _16673_ (.Y(_07578_),
    .A(_07577_));
 sg13g2_nand3_1 _16674_ (.B(_06325_),
    .C(_06318_),
    .A(_06317_),
    .Y(_07579_));
 sg13g2_nand2_1 _16675_ (.Y(_07580_),
    .A(_07579_),
    .B(_06359_));
 sg13g2_nand2_1 _16676_ (.Y(_07581_),
    .A(_06357_),
    .B(_07580_));
 sg13g2_nand3_1 _16677_ (.B(_06322_),
    .C(_07581_),
    .A(_06330_),
    .Y(_07582_));
 sg13g2_inv_1 _16678_ (.Y(_07583_),
    .A(_07582_));
 sg13g2_a21oi_1 _16679_ (.A1(_07578_),
    .A2(net37),
    .Y(_07584_),
    .B1(_07583_));
 sg13g2_inv_1 _16680_ (.Y(_07585_),
    .A(_07584_));
 sg13g2_nor3_1 _16681_ (.A(_06566_),
    .B(_06564_),
    .C(_06569_),
    .Y(_07586_));
 sg13g2_nand2b_1 _16682_ (.Y(_07587_),
    .B(_06585_),
    .A_N(_07586_));
 sg13g2_nand2_1 _16683_ (.Y(_07588_),
    .A(_06582_),
    .B(_07587_));
 sg13g2_nand3_1 _16684_ (.B(_06568_),
    .C(_07588_),
    .A(_06576_),
    .Y(_07589_));
 sg13g2_inv_1 _16685_ (.Y(_07590_),
    .A(_07589_));
 sg13g2_a21oi_1 _16686_ (.A1(_07585_),
    .A2(net26),
    .Y(_07591_),
    .B1(_07590_));
 sg13g2_o21ai_1 _16687_ (.B1(_05356_),
    .Y(_07592_),
    .A1(_07574_),
    .A2(_07591_));
 sg13g2_buf_1 _16688_ (.A(_07592_),
    .X(_07593_));
 sg13g2_a21oi_2 _16689_ (.B1(_06707_),
    .Y(_07594_),
    .A2(net50),
    .A1(_07593_));
 sg13g2_inv_1 _16690_ (.Y(_07595_),
    .A(_07594_));
 sg13g2_a21oi_1 _16691_ (.A1(_07595_),
    .A2(net82),
    .Y(_07596_),
    .B1(_07231_));
 sg13g2_inv_1 _16692_ (.Y(_07597_),
    .A(_07596_));
 sg13g2_a21oi_1 _16693_ (.A1(_05706_),
    .A2(net37),
    .Y(_07598_),
    .B1(_06426_));
 sg13g2_inv_1 _16694_ (.Y(_07599_),
    .A(_07598_));
 sg13g2_a21oi_1 _16695_ (.A1(_07599_),
    .A2(net26),
    .Y(_07600_),
    .B1(_06812_));
 sg13g2_inv_1 _16696_ (.Y(_07601_),
    .A(_07600_));
 sg13g2_a21oi_1 _16697_ (.A1(_07601_),
    .A2(_05347_),
    .Y(_07602_),
    .B1(_05532_));
 sg13g2_inv_1 _16698_ (.Y(_07603_),
    .A(_07602_));
 sg13g2_a21oi_1 _16699_ (.A1(_07603_),
    .A2(net50),
    .Y(_07604_),
    .B1(_06731_));
 sg13g2_inv_1 _16700_ (.Y(_07605_),
    .A(_07604_));
 sg13g2_a21oi_1 _16701_ (.A1(_07605_),
    .A2(net82),
    .Y(_07606_),
    .B1(_04251_));
 sg13g2_a21oi_1 _16702_ (.A1(_07597_),
    .A2(_04979_),
    .Y(_07607_),
    .B1(_07606_));
 sg13g2_nor4_1 _16703_ (.A(_07241_),
    .B(_07571_),
    .C(_07573_),
    .D(_07607_),
    .Y(_07608_));
 sg13g2_nand2_1 _16704_ (.Y(_07609_),
    .A(_07566_),
    .B(_07608_));
 sg13g2_a22oi_1 _16705_ (.Y(_07610_),
    .B1(_07562_),
    .B2(_07560_),
    .A2(_07550_),
    .A1(_07504_));
 sg13g2_inv_1 _16706_ (.Y(_07611_),
    .A(_07570_));
 sg13g2_nor2_1 _16707_ (.A(_04401_),
    .B(_07611_),
    .Y(_07612_));
 sg13g2_nor2_1 _16708_ (.A(_07150_),
    .B(_07612_),
    .Y(_07613_));
 sg13g2_nand2_1 _16709_ (.Y(_07614_),
    .A(_07610_),
    .B(_07613_));
 sg13g2_inv_1 _16710_ (.Y(_07615_),
    .A(_04459_));
 sg13g2_inv_1 _16711_ (.Y(_07616_),
    .A(_05024_));
 sg13g2_nor2_1 _16712_ (.A(_07557_),
    .B(_07616_),
    .Y(_07617_));
 sg13g2_inv_1 _16713_ (.Y(_07618_),
    .A(_07617_));
 sg13g2_nand2_1 _16714_ (.Y(_07619_),
    .A(_07618_),
    .B(_05056_));
 sg13g2_a221oi_1 _16715_ (.B2(_07596_),
    .C1(_07619_),
    .B1(_07606_),
    .A1(_07615_),
    .Y(_07620_),
    .A2(_04466_));
 sg13g2_nor2_1 _16716_ (.A(_07160_),
    .B(_06645_),
    .Y(_07621_));
 sg13g2_inv_1 _16717_ (.Y(_07622_),
    .A(_06650_));
 sg13g2_nand2_1 _16718_ (.Y(_07623_),
    .A(_07621_),
    .B(_07622_));
 sg13g2_inv_1 _16719_ (.Y(_07624_),
    .A(_07623_));
 sg13g2_nand3_1 _16720_ (.B(_07217_),
    .C(_07624_),
    .A(_07620_),
    .Y(_07625_));
 sg13g2_nor3_1 _16721_ (.A(_05062_),
    .B(_07614_),
    .C(_07625_),
    .Y(_07626_));
 sg13g2_nand2b_1 _16722_ (.Y(_07627_),
    .B(_07626_),
    .A_N(_07609_));
 sg13g2_nand3_1 _16723_ (.B(net41),
    .C(_04343_),
    .A(_07627_),
    .Y(_07628_));
 sg13g2_inv_2 _16724_ (.Y(_07629_),
    .A(_04343_));
 sg13g2_nor2_1 _16725_ (.A(net192),
    .B(_07629_),
    .Y(_07630_));
 sg13g2_nand3b_1 _16726_ (.B(_07609_),
    .C(_07630_),
    .Y(_07631_),
    .A_N(_07626_));
 sg13g2_buf_1 _16727_ (.A(_07631_),
    .X(_07632_));
 sg13g2_nand2_1 _16728_ (.Y(_07633_),
    .A(_07628_),
    .B(_07632_));
 sg13g2_nand2_1 _16729_ (.Y(_07634_),
    .A(_07632_),
    .B(_04436_));
 sg13g2_nand2b_1 _16730_ (.Y(_07635_),
    .B(_04349_),
    .A_N(_04351_));
 sg13g2_nand3_1 _16731_ (.B(_07634_),
    .C(_07635_),
    .A(_07633_),
    .Y(_07636_));
 sg13g2_inv_1 _16732_ (.Y(_07637_),
    .A(_04341_));
 sg13g2_nand2_1 _16733_ (.Y(_07638_),
    .A(_07637_),
    .B(net56));
 sg13g2_nand3_1 _16734_ (.B(_07618_),
    .C(_07610_),
    .A(_07566_),
    .Y(_07639_));
 sg13g2_a21oi_1 _16735_ (.A1(_07597_),
    .A2(_07216_),
    .Y(_07640_),
    .B1(_04343_));
 sg13g2_a21oi_1 _16736_ (.A1(_07639_),
    .A2(_07629_),
    .Y(_07641_),
    .B1(_07640_));
 sg13g2_nand2b_1 _16737_ (.Y(_07642_),
    .B(_04353_),
    .A_N(_07641_));
 sg13g2_nand3_1 _16738_ (.B(_07629_),
    .C(_04350_),
    .A(_07639_),
    .Y(_07643_));
 sg13g2_nand2_1 _16739_ (.Y(_07644_),
    .A(_07642_),
    .B(_07643_));
 sg13g2_nand2b_1 _16740_ (.Y(_07645_),
    .B(_07644_),
    .A_N(_07638_));
 sg13g2_buf_1 _16741_ (.A(\b.gen_square[55].sq.mask ),
    .X(_07646_));
 sg13g2_inv_1 _16742_ (.Y(_07647_),
    .A(_07646_));
 sg13g2_a221oi_1 _16743_ (.B2(_07645_),
    .C1(_07647_),
    .B1(_07636_),
    .A1(_01946_),
    .Y(_07648_),
    .A2(_04259_));
 sg13g2_buf_1 _16744_ (.A(_07648_),
    .X(_07649_));
 sg13g2_nand3_1 _16745_ (.B(_04340_),
    .C(_04336_),
    .A(_04338_),
    .Y(_07650_));
 sg13g2_nand2b_1 _16746_ (.Y(_07651_),
    .B(_07640_),
    .A_N(_07650_));
 sg13g2_nand3_1 _16747_ (.B(_07637_),
    .C(_07651_),
    .A(_07642_),
    .Y(_07652_));
 sg13g2_inv_1 _16748_ (.Y(_07653_),
    .A(_04979_));
 sg13g2_nand2_1 _16749_ (.Y(_07654_),
    .A(_05056_),
    .B(_04432_));
 sg13g2_nor4_1 _16750_ (.A(_07241_),
    .B(_07653_),
    .C(_07654_),
    .D(_07571_),
    .Y(_07655_));
 sg13g2_nand4_1 _16751_ (.B(_04341_),
    .C(_04459_),
    .A(_07655_),
    .Y(_07656_),
    .D(_07613_));
 sg13g2_nor2_1 _16752_ (.A(_07629_),
    .B(_07637_),
    .Y(_07657_));
 sg13g2_nor2_1 _16753_ (.A(_02122_),
    .B(_07657_),
    .Y(_07658_));
 sg13g2_nand3_1 _16754_ (.B(_07656_),
    .C(_07658_),
    .A(_07652_),
    .Y(_07659_));
 sg13g2_inv_1 _16755_ (.Y(_07660_),
    .A(_04436_));
 sg13g2_nand2_1 _16756_ (.Y(_07661_),
    .A(_07629_),
    .B(_07660_));
 sg13g2_nand3_1 _16757_ (.B(net41),
    .C(_07661_),
    .A(_07627_),
    .Y(_07662_));
 sg13g2_a21o_1 _16758_ (.A2(_07660_),
    .A1(_04339_),
    .B1(_07662_),
    .X(_07663_));
 sg13g2_nand2b_1 _16759_ (.Y(_07664_),
    .B(_04340_),
    .A_N(_07632_));
 sg13g2_nand3_1 _16760_ (.B(_07663_),
    .C(_07664_),
    .A(_07659_),
    .Y(_07665_));
 sg13g2_nand2_1 _16761_ (.Y(_07666_),
    .A(_07665_),
    .B(_07646_));
 sg13g2_nor2_1 _16762_ (.A(_07482_),
    .B(_07486_),
    .Y(_07667_));
 sg13g2_a21oi_1 _16763_ (.A1(_07480_),
    .A2(_07486_),
    .Y(_07668_),
    .B1(_07667_));
 sg13g2_nor2_1 _16764_ (.A(_07666_),
    .B(_07668_),
    .Y(_07669_));
 sg13g2_o21ai_1 _16765_ (.B1(_07669_),
    .Y(_07670_),
    .A1(_07488_),
    .A2(_07649_));
 sg13g2_nor2b_1 _16766_ (.A(_07294_),
    .B_N(_07306_),
    .Y(_07671_));
 sg13g2_nor3_1 _16767_ (.A(_04337_),
    .B(_04336_),
    .C(_04340_),
    .Y(_07672_));
 sg13g2_nand2_1 _16768_ (.Y(_07673_),
    .A(_07629_),
    .B(_07672_));
 sg13g2_a21oi_1 _16769_ (.A1(_07624_),
    .A2(_07572_),
    .Y(_07674_),
    .B1(_07673_));
 sg13g2_nand2b_1 _16770_ (.Y(_07675_),
    .B(_07651_),
    .A_N(_07674_));
 sg13g2_nor2_1 _16771_ (.A(_07675_),
    .B(_07644_),
    .Y(_07676_));
 sg13g2_nor2_1 _16772_ (.A(_04337_),
    .B(_04351_),
    .Y(_07677_));
 sg13g2_o21ai_1 _16773_ (.B1(_07633_),
    .Y(_07678_),
    .A1(_04353_),
    .A2(_07677_));
 sg13g2_o21ai_1 _16774_ (.B1(_07678_),
    .Y(_07679_),
    .A1(_07638_),
    .A2(_07676_));
 sg13g2_nand2_1 _16775_ (.Y(_07680_),
    .A(_07679_),
    .B(_07646_));
 sg13g2_inv_1 _16776_ (.Y(_07681_),
    .A(_07680_));
 sg13g2_a22oi_1 _16777_ (.Y(_07682_),
    .B1(_07649_),
    .B2(_07488_),
    .A2(_07681_),
    .A1(_07671_));
 sg13g2_nand2_1 _16778_ (.Y(_07683_),
    .A(_07670_),
    .B(_07682_));
 sg13g2_inv_1 _16779_ (.Y(_07684_),
    .A(_07671_));
 sg13g2_nand2_1 _16780_ (.Y(_07685_),
    .A(_07684_),
    .B(_07680_));
 sg13g2_nand2_2 _16781_ (.Y(_07686_),
    .A(_07683_),
    .B(_07685_));
 sg13g2_nor2_1 _16782_ (.A(_07649_),
    .B(_07686_),
    .Y(_07687_));
 sg13g2_a21oi_1 _16783_ (.A1(_07488_),
    .A2(_07686_),
    .Y(_07688_),
    .B1(_07687_));
 sg13g2_inv_1 _16784_ (.Y(_07689_),
    .A(_07688_));
 sg13g2_inv_1 _16785_ (.Y(_07690_),
    .A(_06794_));
 sg13g2_nand2_1 _16786_ (.Y(_07691_),
    .A(_06658_),
    .B(_04772_));
 sg13g2_nand2_1 _16787_ (.Y(_07692_),
    .A(_04769_),
    .B(_07691_));
 sg13g2_nand3_1 _16788_ (.B(_07692_),
    .C(_04663_),
    .A(_04671_),
    .Y(_07693_));
 sg13g2_inv_1 _16789_ (.Y(_07694_),
    .A(_07693_));
 sg13g2_a21oi_1 _16790_ (.A1(_05231_),
    .A2(net31),
    .Y(_07695_),
    .B1(_07694_));
 sg13g2_inv_1 _16791_ (.Y(_07696_),
    .A(_07695_));
 sg13g2_a21oi_2 _16792_ (.B1(_07208_),
    .Y(_07697_),
    .A2(net66),
    .A1(_07696_));
 sg13g2_nand2_1 _16793_ (.Y(_07698_),
    .A(_07690_),
    .B(_07697_));
 sg13g2_o21ai_1 _16794_ (.B1(_07698_),
    .Y(_07699_),
    .A1(_07593_),
    .A2(_07602_));
 sg13g2_inv_1 _16795_ (.Y(_07700_),
    .A(_06175_));
 sg13g2_inv_1 _16796_ (.Y(_07701_),
    .A(_06180_));
 sg13g2_a21oi_2 _16797_ (.B1(_07701_),
    .Y(_07702_),
    .A2(_06222_),
    .A1(_07700_));
 sg13g2_nor2_1 _16798_ (.A(_07702_),
    .B(_06190_),
    .Y(_07703_));
 sg13g2_buf_2 _16799_ (.A(_07703_),
    .X(_07704_));
 sg13g2_a21oi_1 _16800_ (.A1(_04920_),
    .A2(_04930_),
    .Y(_07705_),
    .B1(_04925_));
 sg13g2_nor2_1 _16801_ (.A(_07705_),
    .B(_06192_),
    .Y(_07706_));
 sg13g2_buf_1 _16802_ (.A(_07706_),
    .X(_07707_));
 sg13g2_a21oi_2 _16803_ (.B1(_05344_),
    .Y(_07708_),
    .A2(_05353_),
    .A1(_05339_));
 sg13g2_a21oi_1 _16804_ (.A1(_04098_),
    .A2(_04153_),
    .Y(_07709_),
    .B1(_04224_));
 sg13g2_inv_1 _16805_ (.Y(_07710_),
    .A(_06189_));
 sg13g2_o21ai_1 _16806_ (.B1(_07710_),
    .Y(_07711_),
    .A1(_06184_),
    .A2(_07709_));
 sg13g2_buf_2 _16807_ (.A(_07711_),
    .X(_07712_));
 sg13g2_a21oi_2 _16808_ (.B1(_05532_),
    .Y(_07713_),
    .A2(net55),
    .A1(_07712_));
 sg13g2_nor2_1 _16809_ (.A(_07708_),
    .B(_07713_),
    .Y(_07714_));
 sg13g2_buf_2 _16810_ (.A(_07714_),
    .X(_07715_));
 sg13g2_nor4_1 _16811_ (.A(_06795_),
    .B(_07704_),
    .C(_07707_),
    .D(_07715_),
    .Y(_07716_));
 sg13g2_inv_1 _16812_ (.Y(_07717_),
    .A(_04108_));
 sg13g2_a21oi_1 _16813_ (.A1(_04314_),
    .A2(_07717_),
    .Y(_07718_),
    .B1(_04114_));
 sg13g2_nor2_1 _16814_ (.A(_07718_),
    .B(_04121_),
    .Y(_07719_));
 sg13g2_buf_2 _16815_ (.A(_07719_),
    .X(_07720_));
 sg13g2_inv_1 _16816_ (.Y(_07721_),
    .A(_07720_));
 sg13g2_inv_1 _16817_ (.Y(_07722_),
    .A(_04146_));
 sg13g2_a21oi_1 _16818_ (.A1(_04301_),
    .A2(_07722_),
    .Y(_07723_),
    .B1(_04151_));
 sg13g2_nor2_2 _16819_ (.A(_07723_),
    .B(_06728_),
    .Y(_07724_));
 sg13g2_nand2_1 _16820_ (.Y(_07725_),
    .A(_04440_),
    .B(_04247_));
 sg13g2_nand2_1 _16821_ (.Y(_07726_),
    .A(_04249_),
    .B(_03828_));
 sg13g2_nand2_1 _16822_ (.Y(_07727_),
    .A(_07725_),
    .B(_07726_));
 sg13g2_inv_2 _16823_ (.Y(_07728_),
    .A(_07727_));
 sg13g2_nor2_1 _16824_ (.A(_04979_),
    .B(_07728_),
    .Y(_07729_));
 sg13g2_nor3_1 _16825_ (.A(_07724_),
    .B(_07729_),
    .C(_04134_),
    .Y(_07730_));
 sg13g2_nand3_1 _16826_ (.B(_07721_),
    .C(_07730_),
    .A(_07716_),
    .Y(_07731_));
 sg13g2_inv_1 _16827_ (.Y(_07732_),
    .A(_07056_));
 sg13g2_a21oi_1 _16828_ (.A1(net69),
    .A2(_07732_),
    .Y(_07733_),
    .B1(_04696_));
 sg13g2_nor2_1 _16829_ (.A(_04700_),
    .B(_07733_),
    .Y(_07734_));
 sg13g2_buf_2 _16830_ (.A(_07734_),
    .X(_07735_));
 sg13g2_a21oi_1 _16831_ (.A1(_07301_),
    .A2(net60),
    .Y(_07736_),
    .B1(_05044_));
 sg13g2_nor2b_2 _16832_ (.A(_07736_),
    .B_N(_00034_),
    .Y(_07737_));
 sg13g2_inv_1 _16833_ (.Y(_07738_),
    .A(_04073_));
 sg13g2_nor3_1 _16834_ (.A(_04072_),
    .B(_04070_),
    .C(_07738_),
    .Y(_07739_));
 sg13g2_nand2_1 _16835_ (.Y(_07740_),
    .A(_04081_),
    .B(_07739_));
 sg13g2_inv_1 _16836_ (.Y(_07741_),
    .A(_07740_));
 sg13g2_a21oi_1 _16837_ (.A1(net69),
    .A2(_07741_),
    .Y(_07742_),
    .B1(_07526_));
 sg13g2_nor2_1 _16838_ (.A(_07495_),
    .B(_07742_),
    .Y(_07743_));
 sg13g2_nand3_1 _16839_ (.B(_04207_),
    .C(_04203_),
    .A(_04201_),
    .Y(_07744_));
 sg13g2_nor2_1 _16840_ (.A(_07744_),
    .B(_04284_),
    .Y(_07745_));
 sg13g2_a21oi_1 _16841_ (.A1(_04511_),
    .A2(_07745_),
    .Y(_07746_),
    .B1(_04214_));
 sg13g2_nor2_2 _16842_ (.A(_04218_),
    .B(_07746_),
    .Y(_07747_));
 sg13g2_nor3_1 _16843_ (.A(_05846_),
    .B(_05848_),
    .C(_05855_),
    .Y(_07748_));
 sg13g2_nand2_1 _16844_ (.Y(_07749_),
    .A(_05854_),
    .B(_07748_));
 sg13g2_inv_1 _16845_ (.Y(_07750_),
    .A(_07749_));
 sg13g2_a21oi_1 _16846_ (.A1(net115),
    .A2(_07750_),
    .Y(_07751_),
    .B1(_05861_));
 sg13g2_nor2_2 _16847_ (.A(_05954_),
    .B(_07751_),
    .Y(_07752_));
 sg13g2_nor2_1 _16848_ (.A(_07747_),
    .B(_07752_),
    .Y(_07753_));
 sg13g2_nor3_1 _16849_ (.A(_04879_),
    .B(_04881_),
    .C(_04888_),
    .Y(_07754_));
 sg13g2_nand2_1 _16850_ (.Y(_07755_),
    .A(_04887_),
    .B(_07754_));
 sg13g2_inv_1 _16851_ (.Y(_07756_),
    .A(_07755_));
 sg13g2_a21oi_1 _16852_ (.A1(net115),
    .A2(_07756_),
    .Y(_07757_),
    .B1(_04895_));
 sg13g2_nor2_1 _16853_ (.A(_04965_),
    .B(_07757_),
    .Y(_07758_));
 sg13g2_inv_2 _16854_ (.Y(_07759_),
    .A(_07758_));
 sg13g2_nand3b_1 _16855_ (.B(_07753_),
    .C(_07759_),
    .Y(_07760_),
    .A_N(_07743_));
 sg13g2_nor4_1 _16856_ (.A(_07735_),
    .B(_07737_),
    .C(_07252_),
    .D(_07760_),
    .Y(_07761_));
 sg13g2_nor2b_1 _16857_ (.A(_04353_),
    .B_N(_07650_),
    .Y(_07762_));
 sg13g2_nor3_1 _16858_ (.A(net119),
    .B(_07661_),
    .C(_07762_),
    .Y(_07763_));
 sg13g2_nor2_1 _16859_ (.A(_04346_),
    .B(_07763_),
    .Y(_07764_));
 sg13g2_buf_2 _16860_ (.A(_07764_),
    .X(_07765_));
 sg13g2_nand2_1 _16861_ (.Y(_07766_),
    .A(_07765_),
    .B(_04247_));
 sg13g2_nand2_1 _16862_ (.Y(_07767_),
    .A(_07766_),
    .B(_07230_));
 sg13g2_inv_1 _16863_ (.Y(_07768_),
    .A(_07767_));
 sg13g2_nand2_1 _16864_ (.Y(_07769_),
    .A(_07768_),
    .B(_05060_));
 sg13g2_o21ai_1 _16865_ (.B1(_07769_),
    .Y(_07770_),
    .A1(_06728_),
    .A2(_06690_));
 sg13g2_inv_1 _16866_ (.Y(_07771_),
    .A(_07770_));
 sg13g2_nand2_1 _16867_ (.Y(_07772_),
    .A(_07761_),
    .B(_07771_));
 sg13g2_a21oi_1 _16868_ (.A1(_06088_),
    .A2(net74),
    .Y(_07773_),
    .B1(_05688_));
 sg13g2_inv_1 _16869_ (.Y(_07774_),
    .A(_07773_));
 sg13g2_a21oi_1 _16870_ (.A1(_07774_),
    .A2(net28),
    .Y(_07775_),
    .B1(_06408_));
 sg13g2_inv_1 _16871_ (.Y(_07776_),
    .A(_07775_));
 sg13g2_inv_1 _16872_ (.Y(_07777_),
    .A(_06603_));
 sg13g2_a21oi_2 _16873_ (.B1(_07777_),
    .Y(_07778_),
    .A2(net54),
    .A1(_07776_));
 sg13g2_o21ai_1 _16874_ (.B1(_06984_),
    .Y(_07779_),
    .A1(_06203_),
    .A2(_07778_));
 sg13g2_buf_1 _16875_ (.A(_07779_),
    .X(_07780_));
 sg13g2_a21oi_1 _16876_ (.A1(_06300_),
    .A2(net74),
    .Y(_07781_),
    .B1(_05723_));
 sg13g2_inv_1 _16877_ (.Y(_07782_),
    .A(_07781_));
 sg13g2_a21oi_1 _16878_ (.A1(_07782_),
    .A2(net28),
    .Y(_07783_),
    .B1(_05963_));
 sg13g2_inv_1 _16879_ (.Y(_07784_),
    .A(_07783_));
 sg13g2_a21oi_1 _16880_ (.A1(_07784_),
    .A2(_05378_),
    .Y(_07785_),
    .B1(_05537_));
 sg13g2_inv_1 _16881_ (.Y(_07786_),
    .A(_07785_));
 sg13g2_a21oi_1 _16882_ (.A1(_07786_),
    .A2(_04928_),
    .Y(_07787_),
    .B1(_04972_));
 sg13g2_a21oi_1 _16883_ (.A1(_04985_),
    .A2(_04116_),
    .Y(_07788_),
    .B1(_04120_));
 sg13g2_inv_1 _16884_ (.Y(_07789_),
    .A(_07788_));
 sg13g2_a21oi_1 _16885_ (.A1(_04116_),
    .A2(_07539_),
    .Y(_07790_),
    .B1(_04321_));
 sg13g2_a21oi_1 _16886_ (.A1(_07155_),
    .A2(_04723_),
    .Y(_07791_),
    .B1(_04796_));
 sg13g2_o21ai_1 _16887_ (.B1(_07127_),
    .Y(_07792_),
    .A1(_04127_),
    .A2(_07791_));
 sg13g2_a21oi_1 _16888_ (.A1(_05009_),
    .A2(_04723_),
    .Y(_07793_),
    .B1(_04728_));
 sg13g2_inv_1 _16889_ (.Y(_07794_),
    .A(_07793_));
 sg13g2_a21oi_1 _16890_ (.A1(_07794_),
    .A2(net71),
    .Y(_07795_),
    .B1(_04131_));
 sg13g2_nor2_1 _16891_ (.A(_07792_),
    .B(_07795_),
    .Y(_07796_));
 sg13g2_a221oi_1 _16892_ (.B2(_07115_),
    .C1(_07796_),
    .B1(_07143_),
    .A1(_07789_),
    .Y(_07797_),
    .A2(_07790_));
 sg13g2_o21ai_1 _16893_ (.B1(_07797_),
    .Y(_07798_),
    .A1(_07780_),
    .A2(_07787_));
 sg13g2_nor4_1 _16894_ (.A(_07699_),
    .B(_07731_),
    .C(_07772_),
    .D(_07798_),
    .Y(_07799_));
 sg13g2_nor2_1 _16895_ (.A(_07723_),
    .B(_06729_),
    .Y(_07800_));
 sg13g2_buf_2 _16896_ (.A(_07800_),
    .X(_07801_));
 sg13g2_nand2_1 _16897_ (.Y(_07802_),
    .A(_05060_),
    .B(_06696_));
 sg13g2_inv_2 _16898_ (.Y(_07803_),
    .A(_06731_));
 sg13g2_nand2_1 _16899_ (.Y(_07804_),
    .A(_07802_),
    .B(_07803_));
 sg13g2_nand2_1 _16900_ (.Y(_07805_),
    .A(_07804_),
    .B(net55));
 sg13g2_nand2b_1 _16901_ (.Y(_07806_),
    .B(_07805_),
    .A_N(_05532_));
 sg13g2_nor2_2 _16902_ (.A(_07708_),
    .B(_07806_),
    .Y(_07807_));
 sg13g2_nor2_1 _16903_ (.A(_07705_),
    .B(_07010_),
    .Y(_07808_));
 sg13g2_buf_2 _16904_ (.A(_07808_),
    .X(_07809_));
 sg13g2_inv_1 _16905_ (.Y(_07810_),
    .A(_07809_));
 sg13g2_nor2_1 _16906_ (.A(_07718_),
    .B(_07789_),
    .Y(_07811_));
 sg13g2_buf_2 _16907_ (.A(_07811_),
    .X(_07812_));
 sg13g2_nor2_1 _16908_ (.A(_05062_),
    .B(_07812_),
    .Y(_07813_));
 sg13g2_nor2_1 _16909_ (.A(_07702_),
    .B(_07712_),
    .Y(_07814_));
 sg13g2_buf_2 _16910_ (.A(_07814_),
    .X(_07815_));
 sg13g2_inv_1 _16911_ (.Y(_07816_),
    .A(_07815_));
 sg13g2_nand4_1 _16912_ (.B(_07813_),
    .C(_05055_),
    .A(_07810_),
    .Y(_07817_),
    .D(_07816_));
 sg13g2_nor4_1 _16913_ (.A(_07017_),
    .B(_07801_),
    .C(_07807_),
    .D(_07817_),
    .Y(_07818_));
 sg13g2_inv_1 _16914_ (.Y(_07819_),
    .A(_07593_));
 sg13g2_nand2_1 _16915_ (.Y(_07820_),
    .A(_06689_),
    .B(_06728_));
 sg13g2_o21ai_1 _16916_ (.B1(_07820_),
    .Y(_07821_),
    .A1(_07767_),
    .A2(_07727_));
 sg13g2_a221oi_1 _16917_ (.B2(_07819_),
    .C1(_07821_),
    .B1(_07602_),
    .A1(_06794_),
    .Y(_07822_),
    .A2(_07697_));
 sg13g2_inv_1 _16918_ (.Y(_07823_),
    .A(_07795_));
 sg13g2_nand2_1 _16919_ (.Y(_07824_),
    .A(_07790_),
    .B(_07788_));
 sg13g2_o21ai_1 _16920_ (.B1(_07824_),
    .Y(_07825_),
    .A1(_07792_),
    .A2(_07823_));
 sg13g2_nor2_1 _16921_ (.A(_07116_),
    .B(_07143_),
    .Y(_07826_));
 sg13g2_inv_1 _16922_ (.Y(_07827_),
    .A(_07787_));
 sg13g2_nor2_1 _16923_ (.A(_07780_),
    .B(_07827_),
    .Y(_07828_));
 sg13g2_nor3_1 _16924_ (.A(_07825_),
    .B(_07826_),
    .C(_07828_),
    .Y(_07829_));
 sg13g2_nor2_2 _16925_ (.A(_03892_),
    .B(_07733_),
    .Y(_07830_));
 sg13g2_nor2_1 _16926_ (.A(_03909_),
    .B(_07736_),
    .Y(_07831_));
 sg13g2_inv_1 _16927_ (.Y(_07832_),
    .A(_05208_));
 sg13g2_nand2b_1 _16928_ (.Y(_07833_),
    .B(_07832_),
    .A_N(_07170_));
 sg13g2_nor2_1 _16929_ (.A(_03685_),
    .B(_07742_),
    .Y(_07834_));
 sg13g2_nor2_2 _16930_ (.A(_03639_),
    .B(_07757_),
    .Y(_07835_));
 sg13g2_nor2_1 _16931_ (.A(_07834_),
    .B(_07835_),
    .Y(_07836_));
 sg13g2_nor2_2 _16932_ (.A(_03590_),
    .B(_07746_),
    .Y(_07837_));
 sg13g2_nor2_2 _16933_ (.A(_03567_),
    .B(_07751_),
    .Y(_07838_));
 sg13g2_nor2_1 _16934_ (.A(_07837_),
    .B(_07838_),
    .Y(_07839_));
 sg13g2_nand2_1 _16935_ (.Y(_07840_),
    .A(_07836_),
    .B(_07839_));
 sg13g2_nor4_1 _16936_ (.A(_07830_),
    .B(_07831_),
    .C(_07833_),
    .D(_07840_),
    .Y(_07841_));
 sg13g2_nand4_1 _16937_ (.B(_07822_),
    .C(_07829_),
    .A(_07818_),
    .Y(_07842_),
    .D(_07841_));
 sg13g2_inv_1 _16938_ (.Y(_07843_),
    .A(_07842_));
 sg13g2_nor3_1 _16939_ (.A(net164),
    .B(_07799_),
    .C(_07843_),
    .Y(_07844_));
 sg13g2_nand2_1 _16940_ (.Y(_07845_),
    .A(_07844_),
    .B(_05077_));
 sg13g2_nand2_1 _16941_ (.Y(_07846_),
    .A(_07843_),
    .B(_07799_));
 sg13g2_nand3_1 _16942_ (.B(_05089_),
    .C(_06698_),
    .A(_07846_),
    .Y(_07847_));
 sg13g2_nand2_1 _16943_ (.Y(_07848_),
    .A(_07845_),
    .B(_07847_));
 sg13g2_nand2_1 _16944_ (.Y(_07849_),
    .A(_07845_),
    .B(_06693_));
 sg13g2_nand2b_1 _16945_ (.Y(_07850_),
    .B(_06692_),
    .A_N(_06701_));
 sg13g2_nand3_1 _16946_ (.B(_07849_),
    .C(_07850_),
    .A(_07848_),
    .Y(_07851_));
 sg13g2_inv_1 _16947_ (.Y(_07852_),
    .A(_07829_));
 sg13g2_o21ai_1 _16948_ (.B1(net164),
    .Y(_07853_),
    .A1(_07798_),
    .A2(_07852_));
 sg13g2_nand2_1 _16949_ (.Y(_07854_),
    .A(_07822_),
    .B(_07771_));
 sg13g2_o21ai_1 _16950_ (.B1(net164),
    .Y(_07855_),
    .A1(_07699_),
    .A2(_07854_));
 sg13g2_a21o_1 _16951_ (.A2(_07855_),
    .A1(_07853_),
    .B1(_06702_),
    .X(_07856_));
 sg13g2_o21ai_1 _16952_ (.B1(_07856_),
    .Y(_07857_),
    .A1(_07118_),
    .A2(_07853_));
 sg13g2_nand2_1 _16953_ (.Y(_07858_),
    .A(_07857_),
    .B(net75));
 sg13g2_buf_1 _16954_ (.A(\b.gen_square[37].sq.mask ),
    .X(_07859_));
 sg13g2_inv_1 _16955_ (.Y(_07860_),
    .A(_07859_));
 sg13g2_a21o_1 _16956_ (.A2(_07858_),
    .A1(_07851_),
    .B1(_07860_),
    .X(_07861_));
 sg13g2_buf_1 _16957_ (.A(_07861_),
    .X(_07862_));
 sg13g2_nor2_1 _16958_ (.A(_02089_),
    .B(_04920_),
    .Y(_07863_));
 sg13g2_nand2b_1 _16959_ (.Y(_07864_),
    .B(_04761_),
    .A_N(_06484_));
 sg13g2_nand2_1 _16960_ (.Y(_07865_),
    .A(_04758_),
    .B(_07864_));
 sg13g2_nand3_1 _16961_ (.B(_04638_),
    .C(_07865_),
    .A(_04647_),
    .Y(_07866_));
 sg13g2_inv_1 _16962_ (.Y(_07867_),
    .A(_07866_));
 sg13g2_a21oi_1 _16963_ (.A1(_04650_),
    .A2(_05934_),
    .Y(_07868_),
    .B1(_07867_));
 sg13g2_inv_1 _16964_ (.Y(_07869_),
    .A(_07868_));
 sg13g2_a21oi_2 _16965_ (.B1(_06241_),
    .Y(_07870_),
    .A2(net21),
    .A1(_07869_));
 sg13g2_nand2_1 _16966_ (.Y(_07871_),
    .A(_04504_),
    .B(net98));
 sg13g2_nand2_1 _16967_ (.Y(_07872_),
    .A(_07297_),
    .B(_05105_));
 sg13g2_nor2b_1 _16968_ (.A(_05739_),
    .B_N(_07872_),
    .Y(_07873_));
 sg13g2_nor2_1 _16969_ (.A(_07873_),
    .B(_05044_),
    .Y(_07874_));
 sg13g2_nand2_1 _16970_ (.Y(_07875_),
    .A(_07874_),
    .B(_05037_));
 sg13g2_nand2_1 _16971_ (.Y(_07876_),
    .A(_07871_),
    .B(_07875_));
 sg13g2_nand2_1 _16972_ (.Y(_07877_),
    .A(_07876_),
    .B(_04128_));
 sg13g2_nand2_1 _16973_ (.Y(_07878_),
    .A(_07877_),
    .B(_04948_));
 sg13g2_nor2_1 _16974_ (.A(_03909_),
    .B(net98),
    .Y(_07879_));
 sg13g2_a21oi_1 _16975_ (.A1(_05024_),
    .A2(net98),
    .Y(_07880_),
    .B1(_07879_));
 sg13g2_nand2_1 _16976_ (.Y(_07881_),
    .A(_07880_),
    .B(_04128_));
 sg13g2_nand2_1 _16977_ (.Y(_07882_),
    .A(_04127_),
    .B(_03820_));
 sg13g2_nand2_1 _16978_ (.Y(_07883_),
    .A(_07881_),
    .B(_07882_));
 sg13g2_nor2_1 _16979_ (.A(_07878_),
    .B(_07883_),
    .Y(_07884_));
 sg13g2_a221oi_1 _16980_ (.B2(_06230_),
    .C1(_07884_),
    .B1(_06190_),
    .A1(_07870_),
    .Y(_07885_),
    .A2(_06312_));
 sg13g2_o21ai_1 _16981_ (.B1(_07885_),
    .Y(_07886_),
    .A1(_04909_),
    .A2(_04969_));
 sg13g2_a21oi_1 _16982_ (.A1(_05051_),
    .A2(_04130_),
    .Y(_07887_),
    .B1(_07878_));
 sg13g2_a21o_1 _16983_ (.A2(_06230_),
    .A1(_06191_),
    .B1(_07887_),
    .X(_07888_));
 sg13g2_a221oi_1 _16984_ (.B2(_04908_),
    .C1(_07888_),
    .B1(_04969_),
    .A1(_06468_),
    .Y(_07889_),
    .A2(_07870_));
 sg13g2_inv_1 _16985_ (.Y(_07890_),
    .A(_07889_));
 sg13g2_o21ai_1 _16986_ (.B1(net146),
    .Y(_07891_),
    .A1(_07886_),
    .A2(_07890_));
 sg13g2_or2_1 _16987_ (.X(_07892_),
    .B(_07891_),
    .A(_04931_));
 sg13g2_nand4_1 _16988_ (.B(_04136_),
    .C(_04144_),
    .A(_04148_),
    .Y(_07893_),
    .D(_04137_));
 sg13g2_inv_1 _16989_ (.Y(_07894_),
    .A(_07893_));
 sg13g2_a21oi_1 _16990_ (.A1(net69),
    .A2(_07894_),
    .Y(_07895_),
    .B1(_04151_));
 sg13g2_nor2_2 _16991_ (.A(_03677_),
    .B(_07895_),
    .Y(_07896_));
 sg13g2_nor3_1 _16992_ (.A(_05272_),
    .B(_05274_),
    .C(_05281_),
    .Y(_07897_));
 sg13g2_nand2_1 _16993_ (.Y(_07898_),
    .A(_05280_),
    .B(_07897_));
 sg13g2_inv_1 _16994_ (.Y(_07899_),
    .A(_07898_));
 sg13g2_a21oi_1 _16995_ (.A1(_04509_),
    .A2(_07899_),
    .Y(_07900_),
    .B1(_05287_));
 sg13g2_nor2_1 _16996_ (.A(_03579_),
    .B(_07900_),
    .Y(_07901_));
 sg13g2_buf_2 _16997_ (.A(_07901_),
    .X(_07902_));
 sg13g2_inv_1 _16998_ (.Y(_07903_),
    .A(_07275_));
 sg13g2_a21oi_1 _16999_ (.A1(net60),
    .A2(_07903_),
    .Y(_07904_),
    .B1(_04721_));
 sg13g2_nor2_2 _17000_ (.A(_03900_),
    .B(_07904_),
    .Y(_07905_));
 sg13g2_nor2_1 _17001_ (.A(_06904_),
    .B(_07905_),
    .Y(_07906_));
 sg13g2_inv_1 _17002_ (.Y(_07907_),
    .A(_07906_));
 sg13g2_nor3_1 _17003_ (.A(_07896_),
    .B(_07902_),
    .C(_07907_),
    .Y(_07908_));
 sg13g2_inv_1 _17004_ (.Y(_07909_),
    .A(_06656_));
 sg13g2_a21oi_1 _17005_ (.A1(net78),
    .A2(_07909_),
    .Y(_07910_),
    .B1(_04672_));
 sg13g2_nor2_2 _17006_ (.A(_03884_),
    .B(_07910_),
    .Y(_07911_));
 sg13g2_nor2_1 _17007_ (.A(_03795_),
    .B(_05819_),
    .Y(_07912_));
 sg13g2_nor2_1 _17008_ (.A(_07911_),
    .B(_07912_),
    .Y(_07913_));
 sg13g2_inv_1 _17009_ (.Y(_07914_),
    .A(_06564_));
 sg13g2_nor3_1 _17010_ (.A(_06566_),
    .B(_06563_),
    .C(_07914_),
    .Y(_07915_));
 sg13g2_nand2_1 _17011_ (.Y(_07916_),
    .A(net126),
    .B(_07915_));
 sg13g2_o21ai_1 _17012_ (.B1(_06576_),
    .Y(_07917_),
    .A1(net79),
    .A2(_07916_));
 sg13g2_nand2_1 _17013_ (.Y(_07918_),
    .A(_07917_),
    .B(\b.gen_square[19].sq.color ));
 sg13g2_inv_2 _17014_ (.Y(_07919_),
    .A(_07918_));
 sg13g2_nor3_1 _17015_ (.A(_06373_),
    .B(_06375_),
    .C(_06382_),
    .Y(_07920_));
 sg13g2_nand2_1 _17016_ (.Y(_07921_),
    .A(net127),
    .B(_07920_));
 sg13g2_o21ai_1 _17017_ (.B1(_06388_),
    .Y(_07922_),
    .A1(net79),
    .A2(_07921_));
 sg13g2_nand2_2 _17018_ (.Y(_07923_),
    .A(_07922_),
    .B(\b.gen_square[26].sq.color ));
 sg13g2_nor2b_1 _17019_ (.A(_07919_),
    .B_N(_07923_),
    .Y(_07924_));
 sg13g2_nand3_1 _17020_ (.B(_07913_),
    .C(_07924_),
    .A(_07908_),
    .Y(_07925_));
 sg13g2_nor2_2 _17021_ (.A(_04676_),
    .B(_07910_),
    .Y(_07926_));
 sg13g2_inv_1 _17022_ (.Y(_07927_),
    .A(_07926_));
 sg13g2_nand2_1 _17023_ (.Y(_07928_),
    .A(_05830_),
    .B(_07927_));
 sg13g2_nand2b_1 _17024_ (.Y(_07929_),
    .B(_00071_),
    .A_N(_07904_));
 sg13g2_inv_1 _17025_ (.Y(_07930_),
    .A(_07929_));
 sg13g2_nor2_1 _17026_ (.A(_07029_),
    .B(_07930_),
    .Y(_07931_));
 sg13g2_inv_1 _17027_ (.Y(_07932_),
    .A(_07931_));
 sg13g2_nor2_1 _17028_ (.A(_04222_),
    .B(_07895_),
    .Y(_07933_));
 sg13g2_buf_2 _17029_ (.A(_07933_),
    .X(_07934_));
 sg13g2_nor2_1 _17030_ (.A(_05525_),
    .B(_07900_),
    .Y(_07935_));
 sg13g2_buf_2 _17031_ (.A(_07935_),
    .X(_07936_));
 sg13g2_nor2_1 _17032_ (.A(_07934_),
    .B(_07936_),
    .Y(_07937_));
 sg13g2_nand2_2 _17033_ (.Y(_07938_),
    .A(_07922_),
    .B(_00031_));
 sg13g2_nand2_2 _17034_ (.Y(_07939_),
    .A(_07917_),
    .B(_00059_));
 sg13g2_nand3_1 _17035_ (.B(_07938_),
    .C(_07939_),
    .A(_07937_),
    .Y(_07940_));
 sg13g2_nor3_1 _17036_ (.A(_07928_),
    .B(_07932_),
    .C(_07940_),
    .Y(_07941_));
 sg13g2_nand2b_1 _17037_ (.Y(_07942_),
    .B(_07941_),
    .A_N(_07925_));
 sg13g2_nand2_1 _17038_ (.Y(_07943_),
    .A(_07942_),
    .B(_06638_));
 sg13g2_nand2_1 _17039_ (.Y(_07944_),
    .A(_07892_),
    .B(_07943_));
 sg13g2_o21ai_1 _17040_ (.B1(_04911_),
    .Y(_07945_),
    .A1(_04912_),
    .A2(_04913_));
 sg13g2_a22oi_1 _17041_ (.Y(_07946_),
    .B1(_06980_),
    .B2(_07008_),
    .A2(_07778_),
    .A1(_07786_));
 sg13g2_a21oi_1 _17042_ (.A1(_06828_),
    .A2(_06734_),
    .Y(_07947_),
    .B1(_06737_));
 sg13g2_inv_1 _17043_ (.Y(_07948_),
    .A(_07947_));
 sg13g2_a21oi_1 _17044_ (.A1(_07061_),
    .A2(net30),
    .Y(_07949_),
    .B1(_04787_));
 sg13g2_inv_1 _17045_ (.Y(_07950_),
    .A(_07949_));
 sg13g2_a21oi_1 _17046_ (.A1(_07950_),
    .A2(_06735_),
    .Y(_07951_),
    .B1(_06990_));
 sg13g2_inv_1 _17047_ (.Y(_07952_),
    .A(_06696_));
 sg13g2_o21ai_1 _17048_ (.B1(_07121_),
    .Y(_07953_),
    .A1(_07952_),
    .A2(_07790_));
 sg13g2_buf_1 _17049_ (.A(_07953_),
    .X(_07954_));
 sg13g2_o21ai_1 _17050_ (.B1(_07803_),
    .Y(_07955_),
    .A1(_07952_),
    .A2(_07788_));
 sg13g2_nor2b_1 _17051_ (.A(_07954_),
    .B_N(_07955_),
    .Y(_07956_));
 sg13g2_a21oi_1 _17052_ (.A1(_07948_),
    .A2(_07951_),
    .Y(_07957_),
    .B1(_07956_));
 sg13g2_nand2_1 _17053_ (.Y(_07958_),
    .A(_07946_),
    .B(_07957_));
 sg13g2_inv_1 _17054_ (.Y(_07959_),
    .A(_04542_));
 sg13g2_a21oi_1 _17055_ (.A1(_06699_),
    .A2(_07959_),
    .Y(_07960_),
    .B1(_04546_));
 sg13g2_nor2_1 _17056_ (.A(_07960_),
    .B(_06732_),
    .Y(_07961_));
 sg13g2_buf_1 _17057_ (.A(_07961_),
    .X(_07962_));
 sg13g2_nand2b_1 _17058_ (.Y(_07963_),
    .B(_07883_),
    .A_N(_04069_));
 sg13g2_nand2_1 _17059_ (.Y(_07964_),
    .A(_06796_),
    .B(_07963_));
 sg13g2_a21oi_2 _17060_ (.B1(_04895_),
    .Y(_07965_),
    .A2(_04904_),
    .A1(_04889_));
 sg13g2_nor2_1 _17061_ (.A(_07965_),
    .B(_05959_),
    .Y(_07966_));
 sg13g2_buf_2 _17062_ (.A(_07966_),
    .X(_07967_));
 sg13g2_nor2_1 _17063_ (.A(_06313_),
    .B(_07967_),
    .Y(_07968_));
 sg13g2_inv_1 _17064_ (.Y(_07969_),
    .A(_07968_));
 sg13g2_nor4_1 _17065_ (.A(net14),
    .B(_07704_),
    .C(_07964_),
    .D(_07969_),
    .Y(_07970_));
 sg13g2_inv_1 _17066_ (.Y(_07971_),
    .A(_07970_));
 sg13g2_a21oi_2 _17067_ (.B1(_05375_),
    .Y(_07972_),
    .A2(_05380_),
    .A1(_05370_));
 sg13g2_inv_1 _17068_ (.Y(_07973_),
    .A(_05437_));
 sg13g2_a21oi_2 _17069_ (.B1(_05537_),
    .Y(_07974_),
    .A2(net54),
    .A1(_07973_));
 sg13g2_nor2_2 _17070_ (.A(_07972_),
    .B(_07974_),
    .Y(_07975_));
 sg13g2_nor2_1 _17071_ (.A(_07715_),
    .B(_07975_),
    .Y(_07976_));
 sg13g2_nand3_1 _17072_ (.B(_07941_),
    .C(_07976_),
    .A(_07889_),
    .Y(_07977_));
 sg13g2_nor3_1 _17073_ (.A(_07958_),
    .B(_07971_),
    .C(_07977_),
    .Y(_07978_));
 sg13g2_nand2_1 _17074_ (.Y(_07979_),
    .A(_07015_),
    .B(_05377_));
 sg13g2_inv_1 _17075_ (.Y(_07980_),
    .A(_05537_));
 sg13g2_nand2_1 _17076_ (.Y(_07981_),
    .A(_07979_),
    .B(_07980_));
 sg13g2_nor2_1 _17077_ (.A(_07972_),
    .B(_07981_),
    .Y(_07982_));
 sg13g2_buf_2 _17078_ (.A(_07982_),
    .X(_07983_));
 sg13g2_nand2_1 _17079_ (.Y(_07984_),
    .A(_05052_),
    .B(_04927_));
 sg13g2_inv_1 _17080_ (.Y(_07985_),
    .A(_04972_));
 sg13g2_nand2_1 _17081_ (.Y(_07986_),
    .A(_07984_),
    .B(_07985_));
 sg13g2_nand2_1 _17082_ (.Y(_07987_),
    .A(_07986_),
    .B(_04897_));
 sg13g2_inv_1 _17083_ (.Y(_07988_),
    .A(_04967_));
 sg13g2_nand2_1 _17084_ (.Y(_07989_),
    .A(_07987_),
    .B(_07988_));
 sg13g2_nor2_2 _17085_ (.A(_07965_),
    .B(_07989_),
    .Y(_07990_));
 sg13g2_nor3_1 _17086_ (.A(_07983_),
    .B(_07807_),
    .C(_07990_),
    .Y(_07991_));
 sg13g2_nor2_1 _17087_ (.A(_07960_),
    .B(_07804_),
    .Y(_07992_));
 sg13g2_buf_2 _17088_ (.A(_07992_),
    .X(_07993_));
 sg13g2_nor3_1 _17089_ (.A(_07993_),
    .B(_07017_),
    .C(_07815_),
    .Y(_07994_));
 sg13g2_nand3_1 _17090_ (.B(_06896_),
    .C(_07994_),
    .A(_07991_),
    .Y(_07995_));
 sg13g2_nor2_1 _17091_ (.A(_07955_),
    .B(_07954_),
    .Y(_07996_));
 sg13g2_a21oi_1 _17092_ (.A1(_07007_),
    .A2(_06980_),
    .Y(_07997_),
    .B1(_07996_));
 sg13g2_a22oi_1 _17093_ (.Y(_07998_),
    .B1(_07778_),
    .B2(_07785_),
    .A2(_07951_),
    .A1(_07947_));
 sg13g2_nand2_1 _17094_ (.Y(_07999_),
    .A(_07997_),
    .B(_07998_));
 sg13g2_nor4_1 _17095_ (.A(_07925_),
    .B(_07886_),
    .C(_07995_),
    .D(_07999_),
    .Y(_08000_));
 sg13g2_nand2_1 _17096_ (.Y(_08001_),
    .A(_07978_),
    .B(_08000_));
 sg13g2_nand3_1 _17097_ (.B(_05088_),
    .C(_04929_),
    .A(_08001_),
    .Y(_08002_));
 sg13g2_nor3_1 _17098_ (.A(_04918_),
    .B(_08000_),
    .C(_07978_),
    .Y(_08003_));
 sg13g2_nand2_1 _17099_ (.Y(_08004_),
    .A(_08003_),
    .B(net145));
 sg13g2_a22oi_1 _17100_ (.Y(_08005_),
    .B1(_08002_),
    .B2(_08004_),
    .A2(_07945_),
    .A1(_04933_));
 sg13g2_a21oi_1 _17101_ (.A1(_07863_),
    .A2(_07944_),
    .Y(_08006_),
    .B1(_08005_));
 sg13g2_o21ai_1 _17102_ (.B1(net146),
    .Y(_08007_),
    .A1(_07999_),
    .A2(_07958_));
 sg13g2_nor3_1 _17103_ (.A(_04910_),
    .B(_04914_),
    .C(_08007_),
    .Y(_08008_));
 sg13g2_a21o_1 _17104_ (.A2(_08007_),
    .A1(_07891_),
    .B1(_04933_),
    .X(_08009_));
 sg13g2_nand2b_1 _17105_ (.Y(_08010_),
    .B(_08009_),
    .A_N(_08008_));
 sg13g2_nand2_1 _17106_ (.Y(_08011_),
    .A(_08010_),
    .B(_05113_));
 sg13g2_inv_1 _17107_ (.Y(_08012_),
    .A(\b.gen_square[36].sq.mask ));
 sg13g2_a21oi_1 _17108_ (.A1(_08006_),
    .A2(_08011_),
    .Y(_08013_),
    .B1(_08012_));
 sg13g2_a21oi_1 _17109_ (.A1(_05009_),
    .A2(net30),
    .Y(_08014_),
    .B1(_04702_));
 sg13g2_inv_1 _17110_ (.Y(_08015_),
    .A(_08014_));
 sg13g2_a21oi_2 _17111_ (.B1(_06201_),
    .Y(_08016_),
    .A2(_06198_),
    .A1(_08015_));
 sg13g2_nand2b_1 _17112_ (.Y(_08017_),
    .B(_04783_),
    .A_N(_07053_));
 sg13g2_nand2_1 _17113_ (.Y(_08018_),
    .A(_08017_),
    .B(_04780_));
 sg13g2_nand3_1 _17114_ (.B(_04687_),
    .C(_08018_),
    .A(_04695_),
    .Y(_08019_));
 sg13g2_inv_1 _17115_ (.Y(_08020_),
    .A(_08019_));
 sg13g2_a21oi_1 _17116_ (.A1(_04478_),
    .A2(net30),
    .Y(_08021_),
    .B1(_08020_));
 sg13g2_inv_1 _17117_ (.Y(_08022_),
    .A(_08021_));
 sg13g2_a21oi_1 _17118_ (.A1(_08022_),
    .A2(_06198_),
    .Y(_08023_),
    .B1(_06241_));
 sg13g2_a22oi_1 _17119_ (.Y(_08024_),
    .B1(_05913_),
    .B2(_05959_),
    .A2(_08023_),
    .A1(_08016_));
 sg13g2_nand2_1 _17120_ (.Y(_08025_),
    .A(_05839_),
    .B(_04736_));
 sg13g2_nand3_1 _17121_ (.B(_08025_),
    .C(_04600_),
    .A(net78),
    .Y(_08026_));
 sg13g2_nand2_1 _17122_ (.Y(_08027_),
    .A(_04731_),
    .B(_08026_));
 sg13g2_inv_1 _17123_ (.Y(_08028_),
    .A(_08027_));
 sg13g2_a21oi_1 _17124_ (.A1(_05691_),
    .A2(_08028_),
    .Y(_08029_),
    .B1(_05928_));
 sg13g2_a22oi_1 _17125_ (.Y(_08030_),
    .B1(_06881_),
    .B2(_06890_),
    .A2(_08029_),
    .A1(_05572_));
 sg13g2_nand2_1 _17126_ (.Y(_08031_),
    .A(_08024_),
    .B(_08030_));
 sg13g2_inv_1 _17127_ (.Y(_08032_),
    .A(_05126_));
 sg13g2_a21oi_1 _17128_ (.A1(net78),
    .A2(_08032_),
    .Y(_08033_),
    .B1(_04623_));
 sg13g2_nor2_1 _17129_ (.A(_03859_),
    .B(_08033_),
    .Y(_08034_));
 sg13g2_nor3_1 _17130_ (.A(_05329_),
    .B(_05331_),
    .C(_05338_),
    .Y(_08035_));
 sg13g2_nand2_1 _17131_ (.Y(_08036_),
    .A(_05337_),
    .B(_08035_));
 sg13g2_inv_1 _17132_ (.Y(_08037_),
    .A(_08036_));
 sg13g2_a21oi_1 _17133_ (.A1(net99),
    .A2(_08037_),
    .Y(_08038_),
    .B1(_05344_));
 sg13g2_nor2_1 _17134_ (.A(_03650_),
    .B(_08038_),
    .Y(_08039_));
 sg13g2_buf_2 _17135_ (.A(_08039_),
    .X(_08040_));
 sg13g2_nor3_1 _17136_ (.A(_05579_),
    .B(_05578_),
    .C(_07192_),
    .Y(_08041_));
 sg13g2_nand2_1 _17137_ (.Y(_08042_),
    .A(_05577_),
    .B(_08041_));
 sg13g2_inv_1 _17138_ (.Y(_08043_),
    .A(_08042_));
 sg13g2_inv_1 _17139_ (.Y(_08044_),
    .A(_05585_));
 sg13g2_a21oi_1 _17140_ (.A1(net133),
    .A2(_08043_),
    .Y(_08045_),
    .B1(_08044_));
 sg13g2_nor2_1 _17141_ (.A(_03512_),
    .B(_08045_),
    .Y(_08046_));
 sg13g2_nor2_1 _17142_ (.A(_07919_),
    .B(_08046_),
    .Y(_08047_));
 sg13g2_inv_1 _17143_ (.Y(_08048_),
    .A(_08047_));
 sg13g2_nand4_1 _17144_ (.B(_06054_),
    .C(_06043_),
    .A(_06049_),
    .Y(_08049_),
    .D(_06045_));
 sg13g2_inv_1 _17145_ (.Y(_08050_),
    .A(_08049_));
 sg13g2_a21oi_1 _17146_ (.A1(net133),
    .A2(_08050_),
    .Y(_08051_),
    .B1(_06053_));
 sg13g2_nor2_1 _17147_ (.A(_03611_),
    .B(_08051_),
    .Y(_08052_));
 sg13g2_nor2_1 _17148_ (.A(_08052_),
    .B(_07911_),
    .Y(_08053_));
 sg13g2_nand2_1 _17149_ (.Y(_08054_),
    .A(_08053_),
    .B(_06465_));
 sg13g2_nor4_1 _17150_ (.A(_08034_),
    .B(_08040_),
    .C(_08048_),
    .D(_08054_),
    .Y(_08055_));
 sg13g2_inv_1 _17151_ (.Y(_08056_),
    .A(_08055_));
 sg13g2_a21oi_1 _17152_ (.A1(_05670_),
    .A2(_05680_),
    .Y(_08057_),
    .B1(_05675_));
 sg13g2_a21oi_2 _17153_ (.B1(_05723_),
    .Y(_08058_),
    .A2(_05677_),
    .A1(_05500_));
 sg13g2_inv_2 _17154_ (.Y(_08059_),
    .A(_08058_));
 sg13g2_nor2_1 _17155_ (.A(_08057_),
    .B(_08059_),
    .Y(_08060_));
 sg13g2_buf_2 _17156_ (.A(_08060_),
    .X(_08061_));
 sg13g2_a21oi_2 _17157_ (.B1(_06389_),
    .Y(_08062_),
    .A2(_06383_),
    .A1(_06398_));
 sg13g2_a21oi_2 _17158_ (.B1(_06433_),
    .Y(_08063_),
    .A2(net51),
    .A1(_08059_));
 sg13g2_inv_2 _17159_ (.Y(_08064_),
    .A(_08063_));
 sg13g2_nor2_2 _17160_ (.A(_08062_),
    .B(_08064_),
    .Y(_08065_));
 sg13g2_nor4_1 _17161_ (.A(_05763_),
    .B(_08061_),
    .C(_07983_),
    .D(_08065_),
    .Y(_08066_));
 sg13g2_inv_1 _17162_ (.Y(_08067_),
    .A(_06470_));
 sg13g2_inv_1 _17163_ (.Y(_08068_),
    .A(_07990_));
 sg13g2_a21oi_1 _17164_ (.A1(_05639_),
    .A2(_05653_),
    .Y(_08069_),
    .B1(_05644_));
 sg13g2_a21oi_1 _17165_ (.A1(_06743_),
    .A2(_05646_),
    .Y(_08070_),
    .B1(_05718_));
 sg13g2_inv_1 _17166_ (.Y(_08071_),
    .A(_08070_));
 sg13g2_nor2_2 _17167_ (.A(_08069_),
    .B(_08071_),
    .Y(_08072_));
 sg13g2_a21oi_1 _17168_ (.A1(_05572_),
    .A2(_06121_),
    .Y(_08073_),
    .B1(_08072_));
 sg13g2_nand4_1 _17169_ (.B(_08067_),
    .C(_08068_),
    .A(_08066_),
    .Y(_08074_),
    .D(_08073_));
 sg13g2_inv_1 _17170_ (.Y(_08075_),
    .A(_06984_));
 sg13g2_a21oi_2 _17171_ (.B1(_08075_),
    .Y(_08076_),
    .A2(net58),
    .A1(_07954_));
 sg13g2_o21ai_1 _17172_ (.B1(_06603_),
    .Y(_08077_),
    .A1(_06512_),
    .A2(_08076_));
 sg13g2_buf_1 _17173_ (.A(_08077_),
    .X(_08078_));
 sg13g2_a21oi_2 _17174_ (.B1(_04972_),
    .Y(_08079_),
    .A2(net58),
    .A1(_07955_));
 sg13g2_o21ai_1 _17175_ (.B1(_07980_),
    .Y(_08080_),
    .A1(_06512_),
    .A2(_08079_));
 sg13g2_inv_1 _17176_ (.Y(_08081_),
    .A(_08080_));
 sg13g2_nand2b_1 _17177_ (.Y(_08082_),
    .B(_08081_),
    .A_N(_08078_));
 sg13g2_a22oi_1 _17178_ (.Y(_08083_),
    .B1(_06403_),
    .B2(_06434_),
    .A2(_07773_),
    .A1(_07781_));
 sg13g2_inv_1 _17179_ (.Y(_08084_),
    .A(_05761_));
 sg13g2_inv_4 _17180_ (.A(_04650_),
    .Y(_08085_));
 sg13g2_o21ai_1 _17181_ (.B1(_04764_),
    .Y(_08086_),
    .A1(_06279_),
    .A2(_08085_));
 sg13g2_inv_1 _17182_ (.Y(_08087_),
    .A(_06414_));
 sg13g2_a21oi_1 _17183_ (.A1(_08086_),
    .A2(_05407_),
    .Y(_08088_),
    .B1(_08087_));
 sg13g2_nand2_1 _17184_ (.Y(_08089_),
    .A(_08084_),
    .B(_08088_));
 sg13g2_nand3_1 _17185_ (.B(_08083_),
    .C(_08089_),
    .A(_08082_),
    .Y(_08090_));
 sg13g2_nor4_1 _17186_ (.A(_08031_),
    .B(_08056_),
    .C(_08074_),
    .D(_08090_),
    .Y(_08091_));
 sg13g2_nor2_1 _17187_ (.A(_08078_),
    .B(_08081_),
    .Y(_08092_));
 sg13g2_nor2_1 _17188_ (.A(_06404_),
    .B(_06434_),
    .Y(_08093_));
 sg13g2_nor2_2 _17189_ (.A(_08057_),
    .B(_08058_),
    .Y(_08094_));
 sg13g2_nor2_1 _17190_ (.A(_08062_),
    .B(_08063_),
    .Y(_08095_));
 sg13g2_buf_2 _17191_ (.A(_08095_),
    .X(_08096_));
 sg13g2_inv_1 _17192_ (.Y(_08097_),
    .A(_05572_));
 sg13g2_nand2_1 _17193_ (.Y(_08098_),
    .A(_08097_),
    .B(_08029_));
 sg13g2_o21ai_1 _17194_ (.B1(_08098_),
    .Y(_08099_),
    .A1(_06890_),
    .A2(_06882_));
 sg13g2_nor2_1 _17195_ (.A(_07774_),
    .B(_07781_),
    .Y(_08100_));
 sg13g2_nor2_1 _17196_ (.A(_08069_),
    .B(_06890_),
    .Y(_08101_));
 sg13g2_buf_2 _17197_ (.A(_08101_),
    .X(_08102_));
 sg13g2_inv_1 _17198_ (.Y(_08103_),
    .A(_08102_));
 sg13g2_nand2_1 _17199_ (.Y(_08104_),
    .A(_08103_),
    .B(_05939_));
 sg13g2_nor2_1 _17200_ (.A(_05530_),
    .B(_08038_),
    .Y(_08105_));
 sg13g2_buf_1 _17201_ (.A(_08105_),
    .X(_08106_));
 sg13g2_nand2b_1 _17202_ (.Y(_08107_),
    .B(_00064_),
    .A_N(_08051_));
 sg13g2_inv_1 _17203_ (.Y(_08108_),
    .A(_08107_));
 sg13g2_inv_1 _17204_ (.Y(_08109_),
    .A(_07939_));
 sg13g2_nand2b_1 _17205_ (.Y(_08110_),
    .B(_00032_),
    .A_N(_08045_));
 sg13g2_inv_1 _17206_ (.Y(_08111_),
    .A(_08110_));
 sg13g2_nor2_1 _17207_ (.A(_08109_),
    .B(_08111_),
    .Y(_08112_));
 sg13g2_inv_1 _17208_ (.Y(_08113_),
    .A(_08112_));
 sg13g2_nor3_1 _17209_ (.A(_08106_),
    .B(_08108_),
    .C(_08113_),
    .Y(_08114_));
 sg13g2_inv_1 _17210_ (.Y(_08115_),
    .A(_08033_));
 sg13g2_nand2_1 _17211_ (.Y(_08116_),
    .A(_08115_),
    .B(_00056_));
 sg13g2_nand4_1 _17212_ (.B(_07927_),
    .C(_08116_),
    .A(_08114_),
    .Y(_08117_),
    .D(_06290_));
 sg13g2_nor4_1 _17213_ (.A(_08099_),
    .B(_08100_),
    .C(_08104_),
    .D(_08117_),
    .Y(_08118_));
 sg13g2_nor2b_1 _17214_ (.A(_08084_),
    .B_N(_08088_),
    .Y(_08119_));
 sg13g2_inv_1 _17215_ (.Y(_08120_),
    .A(_08023_));
 sg13g2_nor2_1 _17216_ (.A(_08120_),
    .B(_08016_),
    .Y(_08121_));
 sg13g2_nor2_1 _17217_ (.A(_08119_),
    .B(_08121_),
    .Y(_08122_));
 sg13g2_nand4_1 _17218_ (.B(_06314_),
    .C(_05440_),
    .A(_08118_),
    .Y(_08123_),
    .D(_08122_));
 sg13g2_nor3_1 _17219_ (.A(_08094_),
    .B(_08096_),
    .C(_08123_),
    .Y(_08124_));
 sg13g2_nand2_1 _17220_ (.Y(_08125_),
    .A(_05960_),
    .B(_05913_));
 sg13g2_inv_1 _17221_ (.Y(_08126_),
    .A(_07967_));
 sg13g2_nand3_1 _17222_ (.B(_08125_),
    .C(_08126_),
    .A(_08124_),
    .Y(_08127_));
 sg13g2_nor4_1 _17223_ (.A(_07975_),
    .B(_08092_),
    .C(_08093_),
    .D(_08127_),
    .Y(_08128_));
 sg13g2_nor3_1 _17224_ (.A(_05129_),
    .B(_08091_),
    .C(_08128_),
    .Y(_08129_));
 sg13g2_nand2_1 _17225_ (.Y(_08130_),
    .A(_08129_),
    .B(net177));
 sg13g2_nand2_1 _17226_ (.Y(_08131_),
    .A(_08128_),
    .B(_08091_));
 sg13g2_nand3_1 _17227_ (.B(net129),
    .C(_05918_),
    .A(_08131_),
    .Y(_08132_));
 sg13g2_nand2_1 _17228_ (.Y(_08133_),
    .A(_08130_),
    .B(_08132_));
 sg13g2_xnor2_1 _17229_ (.Y(_08134_),
    .A(_05130_),
    .B(_05914_));
 sg13g2_nand2b_1 _17230_ (.Y(_08135_),
    .B(_08125_),
    .A_N(_08121_));
 sg13g2_nor3_1 _17231_ (.A(_08099_),
    .B(_08135_),
    .C(_08031_),
    .Y(_08136_));
 sg13g2_nor2_1 _17232_ (.A(_05918_),
    .B(_08136_),
    .Y(_08137_));
 sg13g2_nand2_1 _17233_ (.Y(_08138_),
    .A(_08137_),
    .B(_05917_));
 sg13g2_o21ai_1 _17234_ (.B1(_05136_),
    .Y(_08139_),
    .A1(_08056_),
    .A2(_08117_));
 sg13g2_nand2_1 _17235_ (.Y(_08140_),
    .A(_05139_),
    .B(net128));
 sg13g2_a21oi_1 _17236_ (.A1(_08138_),
    .A2(_08139_),
    .Y(_08141_),
    .B1(_08140_));
 sg13g2_a21oi_1 _17237_ (.A1(_08133_),
    .A2(_08134_),
    .Y(_08142_),
    .B1(_08141_));
 sg13g2_nor4_1 _17238_ (.A(_08093_),
    .B(_08100_),
    .C(_08119_),
    .D(_08092_),
    .Y(_08143_));
 sg13g2_inv_1 _17239_ (.Y(_08144_),
    .A(_08090_));
 sg13g2_a21oi_1 _17240_ (.A1(_08143_),
    .A2(_08144_),
    .Y(_08145_),
    .B1(_05918_));
 sg13g2_o21ai_1 _17241_ (.B1(_05916_),
    .Y(_08146_),
    .A1(_08137_),
    .A2(_08145_));
 sg13g2_nand2_1 _17242_ (.Y(_08147_),
    .A(_08145_),
    .B(_06405_));
 sg13g2_a21o_1 _17243_ (.A2(_08147_),
    .A1(_08146_),
    .B1(_08140_),
    .X(_08148_));
 sg13g2_nand2_1 _17244_ (.Y(_08149_),
    .A(_08142_),
    .B(_08148_));
 sg13g2_buf_1 _17245_ (.A(\b.gen_square[34].sq.mask ),
    .X(_08150_));
 sg13g2_nand2_1 _17246_ (.Y(_08151_),
    .A(_08149_),
    .B(_08150_));
 sg13g2_a21oi_1 _17247_ (.A1(_06274_),
    .A2(_04650_),
    .Y(_08152_),
    .B1(_07867_));
 sg13g2_inv_1 _17248_ (.Y(_08153_),
    .A(_08152_));
 sg13g2_a21oi_1 _17249_ (.A1(_08153_),
    .A2(_05568_),
    .Y(_08154_),
    .B1(_05928_));
 sg13g2_inv_1 _17250_ (.Y(_08155_),
    .A(net53));
 sg13g2_inv_1 _17251_ (.Y(_08156_),
    .A(_06933_));
 sg13g2_nor2b_1 _17252_ (.A(_06920_),
    .B_N(_06917_),
    .Y(_08157_));
 sg13g2_a21oi_1 _17253_ (.A1(_06919_),
    .A2(_08157_),
    .Y(_08158_),
    .B1(_06929_));
 sg13g2_o21ai_1 _17254_ (.B1(_06926_),
    .Y(_08159_),
    .A1(_08156_),
    .A2(_08158_));
 sg13g2_inv_1 _17255_ (.Y(_08160_),
    .A(_08159_));
 sg13g2_and3_1 _17256_ (.X(_08161_),
    .A(_06514_),
    .B(_06522_),
    .C(_06515_));
 sg13g2_buf_1 _17257_ (.A(_08161_),
    .X(_08162_));
 sg13g2_o21ai_1 _17258_ (.B1(_06557_),
    .Y(_08163_),
    .A1(_06554_),
    .A2(_08162_));
 sg13g2_nand3_1 _17259_ (.B(_06519_),
    .C(_08163_),
    .A(_06526_),
    .Y(_08164_));
 sg13g2_buf_1 _17260_ (.A(_08164_),
    .X(_08165_));
 sg13g2_inv_1 _17261_ (.Y(_08166_),
    .A(_08165_));
 sg13g2_a21oi_1 _17262_ (.A1(_08160_),
    .A2(net36),
    .Y(_08167_),
    .B1(_08166_));
 sg13g2_inv_1 _17263_ (.Y(_08168_),
    .A(_08167_));
 sg13g2_inv_1 _17264_ (.Y(_08169_),
    .A(_04877_));
 sg13g2_a21oi_2 _17265_ (.B1(_08169_),
    .Y(_08170_),
    .A2(_04959_),
    .A1(_08168_));
 sg13g2_o21ai_1 _17266_ (.B1(_06879_),
    .Y(_08171_),
    .A1(_08155_),
    .A2(_08170_));
 sg13g2_inv_1 _17267_ (.Y(_08172_),
    .A(_08171_));
 sg13g2_o21ai_1 _17268_ (.B1(_05149_),
    .Y(_08173_),
    .A1(_08154_),
    .A2(_08172_));
 sg13g2_nor2b_1 _17269_ (.A(_08173_),
    .B_N(_06303_),
    .Y(_08174_));
 sg13g2_inv_1 _17270_ (.Y(_08175_),
    .A(_07938_));
 sg13g2_nor2_2 _17271_ (.A(_08175_),
    .B(_08111_),
    .Y(_08176_));
 sg13g2_nand3_1 _17272_ (.B(_05830_),
    .C(_08116_),
    .A(_08176_),
    .Y(_08177_));
 sg13g2_inv_1 _17273_ (.Y(_08178_),
    .A(_08177_));
 sg13g2_o21ai_1 _17274_ (.B1(_07923_),
    .Y(_08179_),
    .A1(_03512_),
    .A2(_08045_));
 sg13g2_nor3_1 _17275_ (.A(_07912_),
    .B(_08034_),
    .C(_08179_),
    .Y(_08180_));
 sg13g2_a21oi_1 _17276_ (.A1(_08178_),
    .A2(_08180_),
    .Y(_08181_),
    .B1(_05155_));
 sg13g2_nand3_1 _17277_ (.B(_04595_),
    .C(_04738_),
    .A(_04731_),
    .Y(_08182_));
 sg13g2_nand2_1 _17278_ (.Y(_08183_),
    .A(_05977_),
    .B(_04606_));
 sg13g2_nand2_1 _17279_ (.Y(_08184_),
    .A(_08182_),
    .B(_08183_));
 sg13g2_nand2_1 _17280_ (.Y(_08185_),
    .A(_08184_),
    .B(_06093_));
 sg13g2_nand2_1 _17281_ (.Y(_08186_),
    .A(_08185_),
    .B(_06099_));
 sg13g2_nand2_1 _17282_ (.Y(_08187_),
    .A(_06073_),
    .B(_08186_));
 sg13g2_inv_1 _17283_ (.Y(_08188_),
    .A(net74));
 sg13g2_a21oi_2 _17284_ (.B1(_06408_),
    .Y(_08189_),
    .A2(_05961_),
    .A1(_08078_));
 sg13g2_o21ai_1 _17285_ (.B1(_05687_),
    .Y(_08190_),
    .A1(_08188_),
    .A2(_08189_));
 sg13g2_inv_1 _17286_ (.Y(_08191_),
    .A(_08190_));
 sg13g2_o21ai_1 _17287_ (.B1(_05149_),
    .Y(_08192_),
    .A1(_08187_),
    .A2(_08191_));
 sg13g2_a21oi_1 _17288_ (.A1(_08192_),
    .A2(_08173_),
    .Y(_08193_),
    .B1(_06081_));
 sg13g2_inv_1 _17289_ (.Y(_08194_),
    .A(_08193_));
 sg13g2_o21ai_1 _17290_ (.B1(_08194_),
    .Y(_08195_),
    .A1(_06083_),
    .A2(_08192_));
 sg13g2_nor3_1 _17291_ (.A(_08174_),
    .B(_08181_),
    .C(_08195_),
    .Y(_08196_));
 sg13g2_nand2b_1 _17292_ (.Y(_08197_),
    .B(net143),
    .A_N(_08196_));
 sg13g2_nor2_1 _17293_ (.A(_05150_),
    .B(_06078_),
    .Y(_08198_));
 sg13g2_nand2_1 _17294_ (.Y(_08199_),
    .A(_06084_),
    .B(net161));
 sg13g2_a21oi_2 _17295_ (.B1(_05963_),
    .Y(_08200_),
    .A2(_05961_),
    .A1(_08080_));
 sg13g2_inv_1 _17296_ (.Y(_08201_),
    .A(_05723_));
 sg13g2_o21ai_1 _17297_ (.B1(_08201_),
    .Y(_08202_),
    .A1(_08188_),
    .A2(_08200_));
 sg13g2_nand2_1 _17298_ (.Y(_08203_),
    .A(_08191_),
    .B(_08202_));
 sg13g2_a21oi_1 _17299_ (.A1(_06999_),
    .A2(net36),
    .Y(_08204_),
    .B1(_06808_));
 sg13g2_inv_1 _17300_ (.Y(_08205_),
    .A(_08204_));
 sg13g2_a21oi_1 _17301_ (.A1(_08205_),
    .A2(_04959_),
    .Y(_08206_),
    .B1(_04962_));
 sg13g2_inv_1 _17302_ (.Y(_08207_),
    .A(_08206_));
 sg13g2_a21oi_1 _17303_ (.A1(_08207_),
    .A2(net53),
    .Y(_08208_),
    .B1(_05718_));
 sg13g2_nand2b_1 _17304_ (.Y(_08209_),
    .B(_08172_),
    .A_N(_08208_));
 sg13g2_nand3_1 _17305_ (.B(_05939_),
    .C(_05512_),
    .A(_08103_),
    .Y(_08210_));
 sg13g2_inv_1 _17306_ (.Y(_08211_),
    .A(_06047_));
 sg13g2_a21oi_1 _17307_ (.A1(_08211_),
    .A2(_06066_),
    .Y(_08212_),
    .B1(_06053_));
 sg13g2_buf_1 _17308_ (.A(_08212_),
    .X(_08213_));
 sg13g2_nor2_1 _17309_ (.A(_08213_),
    .B(_06112_),
    .Y(_08214_));
 sg13g2_nor3_1 _17310_ (.A(_08094_),
    .B(_08210_),
    .C(_08214_),
    .Y(_08215_));
 sg13g2_a21oi_1 _17311_ (.A1(_06444_),
    .A2(_04650_),
    .Y(_08216_),
    .B1(_04654_));
 sg13g2_inv_1 _17312_ (.Y(_08217_),
    .A(_08216_));
 sg13g2_a21oi_1 _17313_ (.A1(_08217_),
    .A2(_05568_),
    .Y(_08218_),
    .B1(_05571_));
 sg13g2_nor2b_1 _17314_ (.A(_08218_),
    .B_N(_08154_),
    .Y(_08219_));
 sg13g2_inv_1 _17315_ (.Y(_08220_),
    .A(_00061_));
 sg13g2_nor2_1 _17316_ (.A(_08220_),
    .B(_04606_),
    .Y(_08221_));
 sg13g2_a21oi_2 _17317_ (.B1(_08221_),
    .Y(_08222_),
    .A2(_04606_),
    .A1(_05431_));
 sg13g2_a21oi_1 _17318_ (.A1(_08222_),
    .A2(_06093_),
    .Y(_08223_),
    .B1(_05501_));
 sg13g2_nor2b_1 _17319_ (.A(_08186_),
    .B_N(_08223_),
    .Y(_08224_));
 sg13g2_nor2_1 _17320_ (.A(_06112_),
    .B(_06073_),
    .Y(_08225_));
 sg13g2_nor4_1 _17321_ (.A(_08219_),
    .B(_08224_),
    .C(_08177_),
    .D(_08225_),
    .Y(_08226_));
 sg13g2_nand4_1 _17322_ (.B(_08209_),
    .C(_08215_),
    .A(_08203_),
    .Y(_08227_),
    .D(_08226_));
 sg13g2_nand2b_1 _17323_ (.Y(_08228_),
    .B(_08191_),
    .A_N(_08202_));
 sg13g2_or2_1 _17324_ (.X(_08229_),
    .B(_08223_),
    .A(_08186_));
 sg13g2_nand2b_1 _17325_ (.Y(_08230_),
    .B(_06112_),
    .A_N(_08213_));
 sg13g2_nand2_1 _17326_ (.Y(_08231_),
    .A(_08218_),
    .B(_06121_));
 sg13g2_nand3_1 _17327_ (.B(_06125_),
    .C(_08231_),
    .A(_08230_),
    .Y(_08232_));
 sg13g2_nor3_1 _17328_ (.A(_08061_),
    .B(_08072_),
    .C(_08232_),
    .Y(_08233_));
 sg13g2_nand2_1 _17329_ (.Y(_08234_),
    .A(_08218_),
    .B(_08154_));
 sg13g2_nand2_1 _17330_ (.Y(_08235_),
    .A(_08234_),
    .B(_08180_));
 sg13g2_a221oi_1 _17331_ (.B2(_08172_),
    .C1(_08235_),
    .B1(_08208_),
    .A1(_06112_),
    .Y(_08236_),
    .A2(_06072_));
 sg13g2_nand4_1 _17332_ (.B(_08229_),
    .C(_08233_),
    .A(_08228_),
    .Y(_08237_),
    .D(_08236_));
 sg13g2_or2_1 _17333_ (.X(_08238_),
    .B(_08237_),
    .A(_08227_));
 sg13g2_inv_2 _17334_ (.Y(_08239_),
    .A(_08238_));
 sg13g2_nand4_1 _17335_ (.B(_08227_),
    .C(net191),
    .A(_08237_),
    .Y(_08240_),
    .D(_06084_));
 sg13g2_buf_1 _17336_ (.A(_08240_),
    .X(_08241_));
 sg13g2_o21ai_1 _17337_ (.B1(_08241_),
    .Y(_08242_),
    .A1(_08199_),
    .A2(_08239_));
 sg13g2_o21ai_1 _17338_ (.B1(_08242_),
    .Y(_08243_),
    .A1(_06080_),
    .A2(_08198_));
 sg13g2_inv_1 _17339_ (.Y(_08244_),
    .A(\b.gen_square[32].sq.mask ));
 sg13g2_a21oi_1 _17340_ (.A1(_08197_),
    .A2(_08243_),
    .Y(_08245_),
    .B1(_08244_));
 sg13g2_nor3_1 _17341_ (.A(_06013_),
    .B(_06015_),
    .C(_06023_),
    .Y(_08246_));
 sg13g2_nand2_1 _17342_ (.Y(_08247_),
    .A(_06021_),
    .B(_08246_));
 sg13g2_inv_1 _17343_ (.Y(_08248_),
    .A(_08247_));
 sg13g2_a21oi_1 _17344_ (.A1(net133),
    .A2(_08248_),
    .Y(_08249_),
    .B1(_06028_));
 sg13g2_nor2_1 _17345_ (.A(_06106_),
    .B(_08249_),
    .Y(_08250_));
 sg13g2_nor2_1 _17346_ (.A(_08250_),
    .B(_07758_),
    .Y(_08251_));
 sg13g2_inv_1 _17347_ (.Y(_08252_),
    .A(_05837_));
 sg13g2_a21oi_1 _17348_ (.A1(net78),
    .A2(_08252_),
    .Y(_08253_),
    .B1(_04604_));
 sg13g2_nor2_1 _17349_ (.A(_08220_),
    .B(_08253_),
    .Y(_08254_));
 sg13g2_inv_1 _17350_ (.Y(_08255_),
    .A(_06488_));
 sg13g2_a21oi_2 _17351_ (.B1(_04648_),
    .Y(_08256_),
    .A2(_08255_),
    .A1(net78));
 sg13g2_nor2_1 _17352_ (.A(_04652_),
    .B(_08256_),
    .Y(_08257_));
 sg13g2_nor2_1 _17353_ (.A(_08254_),
    .B(_08257_),
    .Y(_08258_));
 sg13g2_nand2_1 _17354_ (.Y(_08259_),
    .A(_08251_),
    .B(_08258_));
 sg13g2_nor3_1 _17355_ (.A(_04798_),
    .B(_04800_),
    .C(_04807_),
    .Y(_08260_));
 sg13g2_nand2_1 _17356_ (.Y(_08261_),
    .A(_04806_),
    .B(_08260_));
 sg13g2_inv_1 _17357_ (.Y(_08262_),
    .A(_08261_));
 sg13g2_a21oi_1 _17358_ (.A1(_04263_),
    .A2(_08262_),
    .Y(_08263_),
    .B1(_04813_));
 sg13g2_nor2_1 _17359_ (.A(_04960_),
    .B(_08263_),
    .Y(_08264_));
 sg13g2_buf_2 _17360_ (.A(_08264_),
    .X(_08265_));
 sg13g2_nor2_1 _17361_ (.A(_08265_),
    .B(_05183_),
    .Y(_08266_));
 sg13g2_inv_1 _17362_ (.Y(_08267_),
    .A(_08266_));
 sg13g2_nor2_2 _17363_ (.A(_03875_),
    .B(_08256_),
    .Y(_08268_));
 sg13g2_nor2_2 _17364_ (.A(_03535_),
    .B(_08263_),
    .Y(_08269_));
 sg13g2_nor2_1 _17365_ (.A(_08268_),
    .B(_08269_),
    .Y(_08270_));
 sg13g2_inv_1 _17366_ (.Y(_08271_),
    .A(_08270_));
 sg13g2_nor2_1 _17367_ (.A(_03847_),
    .B(_08253_),
    .Y(_08272_));
 sg13g2_nor2_2 _17368_ (.A(_03362_),
    .B(_08249_),
    .Y(_08273_));
 sg13g2_nor2_1 _17369_ (.A(_08273_),
    .B(_07835_),
    .Y(_08274_));
 sg13g2_nand3b_1 _17370_ (.B(_08274_),
    .C(_07832_),
    .Y(_08275_),
    .A_N(_08272_));
 sg13g2_nor4_1 _17371_ (.A(_08259_),
    .B(_08267_),
    .C(_08271_),
    .D(_08275_),
    .Y(_08276_));
 sg13g2_inv_2 _17372_ (.Y(_08277_),
    .A(_06391_));
 sg13g2_nor2_1 _17373_ (.A(_07074_),
    .B(_07086_),
    .Y(_08278_));
 sg13g2_a21oi_1 _17374_ (.A1(_07073_),
    .A2(_08278_),
    .Y(_08279_),
    .B1(_07079_));
 sg13g2_o21ai_1 _17375_ (.B1(_07090_),
    .Y(_08280_),
    .A1(_07084_),
    .A2(_08279_));
 sg13g2_inv_1 _17376_ (.Y(_08281_),
    .A(_08280_));
 sg13g2_and3_1 _17377_ (.X(_08282_),
    .A(_06938_),
    .B(_06946_),
    .C(_06939_));
 sg13g2_nand2b_1 _17378_ (.Y(_08283_),
    .B(_06960_),
    .A_N(_08282_));
 sg13g2_nand2_1 _17379_ (.Y(_08284_),
    .A(_08283_),
    .B(_06957_));
 sg13g2_nand3_1 _17380_ (.B(_06943_),
    .C(_08284_),
    .A(_06951_),
    .Y(_08285_));
 sg13g2_inv_1 _17381_ (.Y(_08286_),
    .A(_08285_));
 sg13g2_a21oi_1 _17382_ (.A1(_08281_),
    .A2(net49),
    .Y(_08287_),
    .B1(_08286_));
 sg13g2_inv_1 _17383_ (.Y(_08288_),
    .A(_08287_));
 sg13g2_a21oi_2 _17384_ (.B1(_07590_),
    .Y(_08289_),
    .A2(net26),
    .A1(_08288_));
 sg13g2_o21ai_1 _17385_ (.B1(_07202_),
    .Y(_08290_),
    .A1(_08277_),
    .A2(_08289_));
 sg13g2_buf_1 _17386_ (.A(_08290_),
    .X(_08291_));
 sg13g2_a21oi_2 _17387_ (.B1(_07694_),
    .Y(_08292_),
    .A2(net44),
    .A1(_06766_));
 sg13g2_o21ai_1 _17388_ (.B1(_05416_),
    .Y(_08293_),
    .A1(_05757_),
    .A2(_08292_));
 sg13g2_buf_1 _17389_ (.A(_08293_),
    .X(_08294_));
 sg13g2_nand4_1 _17390_ (.B(_05252_),
    .C(_06750_),
    .A(_08291_),
    .Y(_08295_),
    .D(_08294_));
 sg13g2_nand3_1 _17391_ (.B(_05668_),
    .C(_06751_),
    .A(_08295_),
    .Y(_08296_));
 sg13g2_o21ai_1 _17392_ (.B1(_08296_),
    .Y(_08297_),
    .A1(_05812_),
    .A2(_08276_));
 sg13g2_inv_1 _17393_ (.Y(_08298_),
    .A(_08200_));
 sg13g2_nor2_1 _17394_ (.A(_05659_),
    .B(_05719_),
    .Y(_08299_));
 sg13g2_a21oi_1 _17395_ (.A1(_08298_),
    .A2(_08189_),
    .Y(_08300_),
    .B1(_08299_));
 sg13g2_inv_1 _17396_ (.Y(_08301_),
    .A(_08300_));
 sg13g2_nand2_1 _17397_ (.Y(_08302_),
    .A(_08189_),
    .B(_08200_));
 sg13g2_a22oi_1 _17398_ (.Y(_08303_),
    .B1(_05658_),
    .B2(_05719_),
    .A2(_06089_),
    .A1(_06114_));
 sg13g2_nor2_1 _17399_ (.A(_05147_),
    .B(_06088_),
    .Y(_08304_));
 sg13g2_nand2_1 _17400_ (.Y(_08305_),
    .A(_04625_),
    .B(_05478_));
 sg13g2_nand2_1 _17401_ (.Y(_08306_),
    .A(_08305_),
    .B(_04753_));
 sg13g2_nand2_1 _17402_ (.Y(_08307_),
    .A(_08306_),
    .B(_05568_));
 sg13g2_nand2_1 _17403_ (.Y(_08308_),
    .A(_08307_),
    .B(_05697_));
 sg13g2_inv_1 _17404_ (.Y(_08309_),
    .A(_08308_));
 sg13g2_nor2_1 _17405_ (.A(_08304_),
    .B(_08309_),
    .Y(_08310_));
 sg13g2_nand3_1 _17406_ (.B(_08303_),
    .C(_08310_),
    .A(_08302_),
    .Y(_08311_));
 sg13g2_o21ai_1 _17407_ (.B1(_05668_),
    .Y(_08312_),
    .A1(_08301_),
    .A2(_08311_));
 sg13g2_nand2_1 _17408_ (.Y(_08313_),
    .A(_08295_),
    .B(_05668_));
 sg13g2_a21o_1 _17409_ (.A2(_08313_),
    .A1(_08312_),
    .B1(_05683_),
    .X(_08314_));
 sg13g2_nand2b_1 _17410_ (.Y(_08315_),
    .B(_05681_),
    .A_N(_08312_));
 sg13g2_nand2_1 _17411_ (.Y(_08316_),
    .A(_08314_),
    .B(_08315_));
 sg13g2_o21ai_1 _17412_ (.B1(net143),
    .Y(_08317_),
    .A1(_08297_),
    .A2(_08316_));
 sg13g2_nand2_1 _17413_ (.Y(_08318_),
    .A(_05440_),
    .B(_08103_));
 sg13g2_a21oi_1 _17414_ (.A1(_04997_),
    .A2(net44),
    .Y(_08319_),
    .B1(_04678_));
 sg13g2_inv_1 _17415_ (.Y(_08320_),
    .A(_08319_));
 sg13g2_a21oi_2 _17416_ (.B1(_05436_),
    .Y(_08321_),
    .A2(_05407_),
    .A1(_08320_));
 sg13g2_a21oi_2 _17417_ (.B1(_05161_),
    .Y(_08322_),
    .A2(_06085_),
    .A1(_05158_));
 sg13g2_nor2_2 _17418_ (.A(_08322_),
    .B(_06114_),
    .Y(_08323_));
 sg13g2_nor2_1 _17419_ (.A(_08213_),
    .B(_06742_),
    .Y(_08324_));
 sg13g2_or4_1 _17420_ (.A(_08323_),
    .B(_08304_),
    .C(_08324_),
    .D(_08267_),
    .X(_08325_));
 sg13g2_nor3_1 _17421_ (.A(_05502_),
    .B(_08259_),
    .C(_08325_),
    .Y(_08326_));
 sg13g2_o21ai_1 _17422_ (.B1(_08326_),
    .Y(_08327_),
    .A1(_08321_),
    .A2(_08294_));
 sg13g2_a21oi_1 _17423_ (.A1(_07137_),
    .A2(net65),
    .Y(_08328_),
    .B1(_07002_));
 sg13g2_inv_1 _17424_ (.Y(_08329_),
    .A(_08328_));
 sg13g2_a21oi_2 _17425_ (.B1(_06812_),
    .Y(_08330_),
    .A2(net26),
    .A1(_08329_));
 sg13g2_inv_1 _17426_ (.Y(_08331_),
    .A(_08330_));
 sg13g2_a21oi_1 _17427_ (.A1(_08331_),
    .A2(net51),
    .Y(_08332_),
    .B1(_06433_));
 sg13g2_nor2_1 _17428_ (.A(_06750_),
    .B(_06742_),
    .Y(_08333_));
 sg13g2_nand2_1 _17429_ (.Y(_08334_),
    .A(_05943_),
    .B(_05568_));
 sg13g2_inv_1 _17430_ (.Y(_08335_),
    .A(_05571_));
 sg13g2_nand2_1 _17431_ (.Y(_08336_),
    .A(_08334_),
    .B(_08335_));
 sg13g2_inv_1 _17432_ (.Y(_08337_),
    .A(_08336_));
 sg13g2_nor2_1 _17433_ (.A(_08308_),
    .B(_08337_),
    .Y(_08338_));
 sg13g2_nor3_1 _17434_ (.A(_05511_),
    .B(_08333_),
    .C(_08338_),
    .Y(_08339_));
 sg13g2_o21ai_1 _17435_ (.B1(_08339_),
    .Y(_08340_),
    .A1(_08291_),
    .A2(_08332_));
 sg13g2_nor4_1 _17436_ (.A(_08096_),
    .B(_08318_),
    .C(_08327_),
    .D(_08340_),
    .Y(_08341_));
 sg13g2_a21oi_2 _17437_ (.B1(_05143_),
    .Y(_08342_),
    .A2(_05138_),
    .A1(_05919_));
 sg13g2_a21oi_2 _17438_ (.B1(_05963_),
    .Y(_08343_),
    .A2(net28),
    .A1(_08097_));
 sg13g2_nor2_1 _17439_ (.A(_08342_),
    .B(_08343_),
    .Y(_08344_));
 sg13g2_buf_2 _17440_ (.A(_08344_),
    .X(_08345_));
 sg13g2_nor2_2 _17441_ (.A(_05573_),
    .B(_08345_),
    .Y(_08346_));
 sg13g2_nand3_1 _17442_ (.B(_08346_),
    .C(_08300_),
    .A(_08341_),
    .Y(_08347_));
 sg13g2_a22oi_1 _17443_ (.Y(_08348_),
    .B1(_08200_),
    .B2(_08189_),
    .A2(_08309_),
    .A1(_08337_));
 sg13g2_nor2_1 _17444_ (.A(_05780_),
    .B(_08275_),
    .Y(_08349_));
 sg13g2_nand2b_1 _17445_ (.Y(_08350_),
    .B(_06742_),
    .A_N(_06750_));
 sg13g2_nor2_1 _17446_ (.A(_08213_),
    .B(_06743_),
    .Y(_08351_));
 sg13g2_nor2_1 _17447_ (.A(_08322_),
    .B(_06300_),
    .Y(_08352_));
 sg13g2_nor2_1 _17448_ (.A(_08351_),
    .B(_08352_),
    .Y(_08353_));
 sg13g2_nand4_1 _17449_ (.B(_08350_),
    .C(_08270_),
    .A(_08349_),
    .Y(_08354_),
    .D(_08353_));
 sg13g2_inv_1 _17450_ (.Y(_08355_),
    .A(_08332_));
 sg13g2_nand2b_1 _17451_ (.Y(_08356_),
    .B(_08321_),
    .A_N(_08294_));
 sg13g2_o21ai_1 _17452_ (.B1(_08356_),
    .Y(_08357_),
    .A1(_08291_),
    .A2(_08355_));
 sg13g2_nor4_1 _17453_ (.A(_05779_),
    .B(_08065_),
    .C(_08354_),
    .D(_08357_),
    .Y(_08358_));
 sg13g2_nor2_1 _17454_ (.A(_08342_),
    .B(_06893_),
    .Y(_08359_));
 sg13g2_buf_2 _17455_ (.A(_08359_),
    .X(_08360_));
 sg13g2_nor4_1 _17456_ (.A(_05771_),
    .B(_08072_),
    .C(_05763_),
    .D(_08360_),
    .Y(_08361_));
 sg13g2_nand4_1 _17457_ (.B(_08358_),
    .C(_08303_),
    .A(_08348_),
    .Y(_08362_),
    .D(_08361_));
 sg13g2_nor2_1 _17458_ (.A(_08347_),
    .B(_08362_),
    .Y(_08363_));
 sg13g2_inv_1 _17459_ (.Y(_08364_),
    .A(_08363_));
 sg13g2_nand3_1 _17460_ (.B(net144),
    .C(_05679_),
    .A(_08364_),
    .Y(_08365_));
 sg13g2_nand4_1 _17461_ (.B(net191),
    .C(_08347_),
    .A(_08362_),
    .Y(_08366_),
    .D(_05679_));
 sg13g2_buf_1 _17462_ (.A(_08366_),
    .X(_08367_));
 sg13g2_nand2_1 _17463_ (.Y(_08368_),
    .A(_08365_),
    .B(_08367_));
 sg13g2_xnor2_1 _17464_ (.Y(_08369_),
    .A(_05660_),
    .B(_05682_));
 sg13g2_nand2_1 _17465_ (.Y(_08370_),
    .A(_08368_),
    .B(_08369_));
 sg13g2_nand2_1 _17466_ (.Y(_08371_),
    .A(_08317_),
    .B(_08370_));
 sg13g2_buf_1 _17467_ (.A(\b.gen_square[33].sq.mask ),
    .X(_08372_));
 sg13g2_nand2_1 _17468_ (.Y(_08373_),
    .A(_08371_),
    .B(_08372_));
 sg13g2_nor2b_1 _17469_ (.A(_08245_),
    .B_N(_08373_),
    .Y(_08374_));
 sg13g2_nand2_1 _17470_ (.Y(_08375_),
    .A(_08151_),
    .B(_08374_));
 sg13g2_nor2_1 _17471_ (.A(_02078_),
    .B(_05370_),
    .Y(_08376_));
 sg13g2_nand2b_1 _17472_ (.Y(_08377_),
    .B(_04750_),
    .A_N(_05420_));
 sg13g2_nand2_1 _17473_ (.Y(_08378_),
    .A(_08377_),
    .B(_04746_));
 sg13g2_nand3_1 _17474_ (.B(_04745_),
    .C(_04615_),
    .A(_08378_),
    .Y(_08379_));
 sg13g2_inv_1 _17475_ (.Y(_08380_),
    .A(_08379_));
 sg13g2_a21oi_1 _17476_ (.A1(_04625_),
    .A2(_05270_),
    .Y(_08381_),
    .B1(_08380_));
 sg13g2_inv_1 _17477_ (.Y(_08382_),
    .A(_08381_));
 sg13g2_a21oi_1 _17478_ (.A1(_08382_),
    .A2(_05408_),
    .Y(_08383_),
    .B1(_05417_));
 sg13g2_inv_1 _17479_ (.Y(_08384_),
    .A(_08383_));
 sg13g2_nor2_1 _17480_ (.A(_08384_),
    .B(_07973_),
    .Y(_08385_));
 sg13g2_a21oi_1 _17481_ (.A1(_07288_),
    .A2(_07277_),
    .Y(_08386_),
    .B1(_04790_));
 sg13g2_nor2_1 _17482_ (.A(_08386_),
    .B(_04721_),
    .Y(_08387_));
 sg13g2_nand2_1 _17483_ (.Y(_08388_),
    .A(_08387_),
    .B(_04711_));
 sg13g2_nand2_1 _17484_ (.Y(_08389_),
    .A(_04723_),
    .B(_07216_));
 sg13g2_nand2_1 _17485_ (.Y(_08390_),
    .A(_08388_),
    .B(_08389_));
 sg13g2_nand2_1 _17486_ (.Y(_08391_),
    .A(_08390_),
    .B(_06734_));
 sg13g2_nand2_1 _17487_ (.Y(_08392_),
    .A(_08391_),
    .B(_06718_));
 sg13g2_nand2_1 _17488_ (.Y(_08393_),
    .A(_04466_),
    .B(_04723_));
 sg13g2_nand2_1 _17489_ (.Y(_08394_),
    .A(_04726_),
    .B(\b.gen_square[53].sq.color ));
 sg13g2_nand3_1 _17490_ (.B(_08394_),
    .C(_06734_),
    .A(_08393_),
    .Y(_08395_));
 sg13g2_nand2_1 _17491_ (.Y(_08396_),
    .A(_06662_),
    .B(_03812_));
 sg13g2_nand2_1 _17492_ (.Y(_08397_),
    .A(_08395_),
    .B(_08396_));
 sg13g2_nor2_1 _17493_ (.A(_08392_),
    .B(_08397_),
    .Y(_08398_));
 sg13g2_nor2_1 _17494_ (.A(_07205_),
    .B(_07184_),
    .Y(_08399_));
 sg13g2_nor3_1 _17495_ (.A(_08385_),
    .B(_08398_),
    .C(_08399_),
    .Y(_08400_));
 sg13g2_nor2b_1 _17496_ (.A(_05358_),
    .B_N(_08400_),
    .Y(_08401_));
 sg13g2_nor2_1 _17497_ (.A(_05437_),
    .B(_08384_),
    .Y(_08402_));
 sg13g2_a21oi_1 _17498_ (.A1(_07014_),
    .A2(_07013_),
    .Y(_08403_),
    .B1(_08392_));
 sg13g2_nor2_1 _17499_ (.A(_07205_),
    .B(_07183_),
    .Y(_08404_));
 sg13g2_nor3_1 _17500_ (.A(_08402_),
    .B(_08403_),
    .C(_08404_),
    .Y(_08405_));
 sg13g2_a21oi_1 _17501_ (.A1(_08401_),
    .A2(_08405_),
    .Y(_08406_),
    .B1(_05379_));
 sg13g2_nand2b_1 _17502_ (.Y(_08407_),
    .B(_08406_),
    .A_N(_05381_));
 sg13g2_nor2_1 _17503_ (.A(_06625_),
    .B(_07735_),
    .Y(_08408_));
 sg13g2_nor2_1 _17504_ (.A(_08265_),
    .B(_07752_),
    .Y(_08409_));
 sg13g2_nand4_1 _17505_ (.B(_06181_),
    .C(_06171_),
    .A(_06177_),
    .Y(_08410_),
    .D(_06173_));
 sg13g2_inv_1 _17506_ (.Y(_08411_),
    .A(_08410_));
 sg13g2_a21oi_1 _17507_ (.A1(net88),
    .A2(_08411_),
    .Y(_08412_),
    .B1(_07701_));
 sg13g2_nor2_2 _17508_ (.A(_06187_),
    .B(_08412_),
    .Y(_08413_));
 sg13g2_nor3_1 _17509_ (.A(_05629_),
    .B(_05631_),
    .C(_05638_),
    .Y(_08414_));
 sg13g2_nand2_1 _17510_ (.Y(_08415_),
    .A(_05637_),
    .B(_08414_));
 sg13g2_inv_1 _17511_ (.Y(_08416_),
    .A(_08415_));
 sg13g2_a21oi_1 _17512_ (.A1(net133),
    .A2(_08416_),
    .Y(_08417_),
    .B1(_05644_));
 sg13g2_nor2_2 _17513_ (.A(_05716_),
    .B(_08417_),
    .Y(_08418_));
 sg13g2_nor2_1 _17514_ (.A(_08413_),
    .B(_08418_),
    .Y(_08419_));
 sg13g2_nor2_1 _17515_ (.A(_08257_),
    .B(_06620_),
    .Y(_08420_));
 sg13g2_nand4_1 _17516_ (.B(_08409_),
    .C(_08419_),
    .A(_08408_),
    .Y(_08421_),
    .D(_08420_));
 sg13g2_nor2_2 _17517_ (.A(_03658_),
    .B(_08412_),
    .Y(_08422_));
 sg13g2_nor2_2 _17518_ (.A(_03621_),
    .B(_08417_),
    .Y(_08423_));
 sg13g2_nor2_1 _17519_ (.A(_08423_),
    .B(_07830_),
    .Y(_08424_));
 sg13g2_nand2_1 _17520_ (.Y(_08425_),
    .A(_08424_),
    .B(_06652_));
 sg13g2_nor4_1 _17521_ (.A(_08422_),
    .B(_08271_),
    .C(_07838_),
    .D(_08425_),
    .Y(_08426_));
 sg13g2_inv_1 _17522_ (.Y(_08427_),
    .A(_08426_));
 sg13g2_o21ai_1 _17523_ (.B1(_06293_),
    .Y(_08428_),
    .A1(_08421_),
    .A2(_08427_));
 sg13g2_nand2_1 _17524_ (.Y(_08429_),
    .A(_08407_),
    .B(_08428_));
 sg13g2_xnor2_1 _17525_ (.Y(_08430_),
    .A(_05360_),
    .B(_05382_));
 sg13g2_inv_1 _17526_ (.Y(_08431_),
    .A(_08405_));
 sg13g2_a21oi_2 _17527_ (.B1(_04678_),
    .Y(_08432_),
    .A2(net44),
    .A1(_06444_));
 sg13g2_inv_2 _17528_ (.Y(_08433_),
    .A(_08432_));
 sg13g2_a21oi_2 _17529_ (.B1(_06201_),
    .Y(_08434_),
    .A2(_06198_),
    .A1(_08433_));
 sg13g2_a21oi_1 _17530_ (.A1(_06510_),
    .A2(net44),
    .Y(_08435_),
    .B1(_04776_));
 sg13g2_inv_2 _17531_ (.Y(_08436_),
    .A(_08435_));
 sg13g2_a21oi_1 _17532_ (.A1(_08436_),
    .A2(_06198_),
    .Y(_08437_),
    .B1(_06611_));
 sg13g2_inv_1 _17533_ (.Y(_08438_),
    .A(_08437_));
 sg13g2_nand2_1 _17534_ (.Y(_08439_),
    .A(_07784_),
    .B(_07775_));
 sg13g2_o21ai_1 _17535_ (.B1(_08439_),
    .Y(_08440_),
    .A1(_08434_),
    .A2(_08438_));
 sg13g2_a21oi_1 _17536_ (.A1(_06835_),
    .A2(_08397_),
    .Y(_08441_),
    .B1(_06313_));
 sg13g2_inv_1 _17537_ (.Y(_08442_),
    .A(_08096_));
 sg13g2_and3_1 _17538_ (.X(_08443_),
    .A(_08441_),
    .B(_05440_),
    .C(_08442_));
 sg13g2_o21ai_1 _17539_ (.B1(_08443_),
    .Y(_08444_),
    .A1(_05533_),
    .A2(_05359_));
 sg13g2_nor4_1 _17540_ (.A(_08431_),
    .B(_08440_),
    .C(_08421_),
    .D(_08444_),
    .Y(_08445_));
 sg13g2_nor2_1 _17541_ (.A(_07715_),
    .B(_07707_),
    .Y(_08446_));
 sg13g2_inv_1 _17542_ (.Y(_08447_),
    .A(_08345_));
 sg13g2_nand2_1 _17543_ (.Y(_08448_),
    .A(_08126_),
    .B(_08447_));
 sg13g2_inv_1 _17544_ (.Y(_08449_),
    .A(_08076_));
 sg13g2_nand2_1 _17545_ (.Y(_08450_),
    .A(_06816_),
    .B(_06597_));
 sg13g2_o21ai_1 _17546_ (.B1(_08450_),
    .Y(_08451_),
    .A1(_08079_),
    .A2(_08449_));
 sg13g2_nor2_1 _17547_ (.A(_08448_),
    .B(_08451_),
    .Y(_08452_));
 sg13g2_nand3_1 _17548_ (.B(_08446_),
    .C(_08452_),
    .A(_08445_),
    .Y(_08453_));
 sg13g2_inv_1 _17549_ (.Y(_08454_),
    .A(_08453_));
 sg13g2_o21ai_1 _17550_ (.B1(_08400_),
    .Y(_08455_),
    .A1(_05534_),
    .A2(_05359_));
 sg13g2_a22oi_1 _17551_ (.Y(_08456_),
    .B1(_06597_),
    .B2(_06815_),
    .A2(_07775_),
    .A1(_07783_));
 sg13g2_a22oi_1 _17552_ (.Y(_08457_),
    .B1(_08079_),
    .B2(_08076_),
    .A2(_08437_),
    .A1(_08434_));
 sg13g2_nand2_1 _17553_ (.Y(_08458_),
    .A(_08456_),
    .B(_08457_));
 sg13g2_inv_1 _17554_ (.Y(_08459_),
    .A(_08065_));
 sg13g2_inv_1 _17555_ (.Y(_08460_),
    .A(_07017_));
 sg13g2_nand3_1 _17556_ (.B(_08067_),
    .C(_08460_),
    .A(_08459_),
    .Y(_08461_));
 sg13g2_nor3_1 _17557_ (.A(_08360_),
    .B(_05763_),
    .C(_08461_),
    .Y(_08462_));
 sg13g2_inv_2 _17558_ (.Y(_08463_),
    .A(_07807_));
 sg13g2_nand4_1 _17559_ (.B(_08068_),
    .C(_08462_),
    .A(_07810_),
    .Y(_08464_),
    .D(_08463_));
 sg13g2_nor4_1 _17560_ (.A(_08455_),
    .B(_08458_),
    .C(_08427_),
    .D(_08464_),
    .Y(_08465_));
 sg13g2_nor3_1 _17561_ (.A(_05368_),
    .B(_08454_),
    .C(_08465_),
    .Y(_08466_));
 sg13g2_nand2_1 _17562_ (.Y(_08467_),
    .A(_08466_),
    .B(_05075_));
 sg13g2_nand2_1 _17563_ (.Y(_08468_),
    .A(_08465_),
    .B(_08454_));
 sg13g2_nand3_1 _17564_ (.B(net113),
    .C(_05379_),
    .A(_08468_),
    .Y(_08469_));
 sg13g2_nand2_1 _17565_ (.Y(_08470_),
    .A(_08467_),
    .B(_08469_));
 sg13g2_a22oi_1 _17566_ (.Y(_08471_),
    .B1(_08430_),
    .B2(_08470_),
    .A2(_08429_),
    .A1(_08376_));
 sg13g2_nor3_1 _17567_ (.A(_08440_),
    .B(_08451_),
    .C(_08458_),
    .Y(_08472_));
 sg13g2_nand2b_1 _17568_ (.Y(_08473_),
    .B(_05368_),
    .A_N(_08472_));
 sg13g2_inv_1 _17569_ (.Y(_08474_),
    .A(_08406_));
 sg13g2_a21o_1 _17570_ (.A2(_08474_),
    .A1(_08473_),
    .B1(_05383_),
    .X(_08475_));
 sg13g2_o21ai_1 _17571_ (.B1(_08475_),
    .Y(_08476_),
    .A1(_06599_),
    .A2(_08473_));
 sg13g2_nand2_1 _17572_ (.Y(_08477_),
    .A(_08476_),
    .B(net95));
 sg13g2_nand2_1 _17573_ (.Y(_08478_),
    .A(_08471_),
    .B(_08477_));
 sg13g2_buf_1 _17574_ (.A(\b.gen_square[35].sq.mask ),
    .X(_08479_));
 sg13g2_nand2_1 _17575_ (.Y(_08480_),
    .A(_08478_),
    .B(_08479_));
 sg13g2_nor2b_1 _17576_ (.A(_08375_),
    .B_N(_08480_),
    .Y(_08481_));
 sg13g2_inv_1 _17577_ (.Y(_08482_),
    .A(_08481_));
 sg13g2_nor2_1 _17578_ (.A(_08013_),
    .B(_08482_),
    .Y(_08483_));
 sg13g2_inv_1 _17579_ (.Y(_08484_),
    .A(_08483_));
 sg13g2_nor2_1 _17580_ (.A(net72),
    .B(_07959_),
    .Y(_08485_));
 sg13g2_nand2b_1 _17581_ (.Y(_08486_),
    .B(_06700_),
    .A_N(_07855_));
 sg13g2_a21o_1 _17582_ (.A2(_07841_),
    .A1(_07761_),
    .B1(_04538_),
    .X(_08487_));
 sg13g2_nand2_1 _17583_ (.Y(_08488_),
    .A(_08486_),
    .B(_08487_));
 sg13g2_xnor2_1 _17584_ (.Y(_08489_),
    .A(_04533_),
    .B(_06701_));
 sg13g2_a22oi_1 _17585_ (.Y(_08490_),
    .B1(_08489_),
    .B2(_07848_),
    .A2(_08488_),
    .A1(_08485_));
 sg13g2_nand2_1 _17586_ (.Y(_08491_),
    .A(_08490_),
    .B(_07858_));
 sg13g2_nand2_1 _17587_ (.Y(_08492_),
    .A(_08491_),
    .B(_07859_));
 sg13g2_nand2b_1 _17588_ (.Y(_08493_),
    .B(_05664_),
    .A_N(_05682_));
 sg13g2_nand2_1 _17589_ (.Y(_08494_),
    .A(_08367_),
    .B(_05665_));
 sg13g2_nand3_1 _17590_ (.B(_08493_),
    .C(_08494_),
    .A(_08368_),
    .Y(_08495_));
 sg13g2_nand2_1 _17591_ (.Y(_08496_),
    .A(_08316_),
    .B(net143));
 sg13g2_nand2_1 _17592_ (.Y(_08497_),
    .A(_08495_),
    .B(_08496_));
 sg13g2_nand2_1 _17593_ (.Y(_08498_),
    .A(_08497_),
    .B(_08372_));
 sg13g2_a21oi_1 _17594_ (.A1(_05679_),
    .A2(_05669_),
    .Y(_08499_),
    .B1(_05665_));
 sg13g2_nor3_1 _17595_ (.A(net158),
    .B(_08499_),
    .C(_08363_),
    .Y(_08500_));
 sg13g2_nand3_1 _17596_ (.B(_05671_),
    .C(_08296_),
    .A(_08314_),
    .Y(_08501_));
 sg13g2_nand2_1 _17597_ (.Y(_08502_),
    .A(_08322_),
    .B(_05510_));
 sg13g2_nand3_1 _17598_ (.B(_05670_),
    .C(_08213_),
    .A(_08062_),
    .Y(_08503_));
 sg13g2_nor4_1 _17599_ (.A(_08502_),
    .B(_08102_),
    .C(_08503_),
    .D(_05439_),
    .Y(_08504_));
 sg13g2_nand3_1 _17600_ (.B(_08346_),
    .C(_08504_),
    .A(_08361_),
    .Y(_08505_));
 sg13g2_nor2_1 _17601_ (.A(net120),
    .B(_05672_),
    .Y(_08506_));
 sg13g2_nand3_1 _17602_ (.B(_08505_),
    .C(_08506_),
    .A(_08501_),
    .Y(_08507_));
 sg13g2_o21ai_1 _17603_ (.B1(_08507_),
    .Y(_08508_),
    .A1(_05663_),
    .A2(_08367_));
 sg13g2_o21ai_1 _17604_ (.B1(_08372_),
    .Y(_08509_),
    .A1(_08500_),
    .A2(_08508_));
 sg13g2_nor2_1 _17605_ (.A(_05152_),
    .B(_08241_),
    .Y(_08510_));
 sg13g2_nand3_1 _17606_ (.B(_05158_),
    .C(_08215_),
    .A(_08233_),
    .Y(_08511_));
 sg13g2_nand2_1 _17607_ (.Y(_08512_),
    .A(_08511_),
    .B(net143));
 sg13g2_nor3_1 _17608_ (.A(_05158_),
    .B(_08174_),
    .C(_08193_),
    .Y(_08513_));
 sg13g2_nor3_1 _17609_ (.A(_05159_),
    .B(_08512_),
    .C(_08513_),
    .Y(_08514_));
 sg13g2_nor2_1 _17610_ (.A(_06075_),
    .B(_06084_),
    .Y(_08515_));
 sg13g2_nor2_1 _17611_ (.A(_05153_),
    .B(_06075_),
    .Y(_08516_));
 sg13g2_nor4_1 _17612_ (.A(net158),
    .B(_08515_),
    .C(_08516_),
    .D(_08239_),
    .Y(_08517_));
 sg13g2_nor3_1 _17613_ (.A(_08510_),
    .B(_08514_),
    .C(_08517_),
    .Y(_08518_));
 sg13g2_nor2_1 _17614_ (.A(_08244_),
    .B(_08518_),
    .Y(_08519_));
 sg13g2_nand2_1 _17615_ (.Y(_08520_),
    .A(_08241_),
    .B(_06075_));
 sg13g2_nand2_1 _17616_ (.Y(_08521_),
    .A(_06079_),
    .B(_06074_));
 sg13g2_nand3_1 _17617_ (.B(_08520_),
    .C(_08521_),
    .A(_08242_),
    .Y(_08522_));
 sg13g2_nand2_1 _17618_ (.Y(_08523_),
    .A(_08195_),
    .B(_05109_));
 sg13g2_nand2_1 _17619_ (.Y(_08524_),
    .A(_08522_),
    .B(_08523_));
 sg13g2_nand2_1 _17620_ (.Y(_08525_),
    .A(_08524_),
    .B(\b.gen_square[32].sq.mask ));
 sg13g2_inv_1 _17621_ (.Y(_08526_),
    .A(_08525_));
 sg13g2_nor2_1 _17622_ (.A(_08498_),
    .B(_08526_),
    .Y(_08527_));
 sg13g2_a21oi_1 _17623_ (.A1(_08509_),
    .A2(_08519_),
    .Y(_08528_),
    .B1(_08527_));
 sg13g2_nor2_1 _17624_ (.A(_08373_),
    .B(_08245_),
    .Y(_08529_));
 sg13g2_nand2_1 _17625_ (.Y(_08530_),
    .A(_08245_),
    .B(_08373_));
 sg13g2_nor2b_1 _17626_ (.A(_08529_),
    .B_N(_08530_),
    .Y(_08531_));
 sg13g2_nand2_1 _17627_ (.Y(_08532_),
    .A(_08526_),
    .B(_08498_));
 sg13g2_nor2_1 _17628_ (.A(_08519_),
    .B(_08509_),
    .Y(_08533_));
 sg13g2_nand4_1 _17629_ (.B(_08531_),
    .C(_08532_),
    .A(_08528_),
    .Y(_08534_),
    .D(_08533_));
 sg13g2_a21oi_1 _17630_ (.A1(_08527_),
    .A2(_08530_),
    .Y(_08535_),
    .B1(_08529_));
 sg13g2_nand2_2 _17631_ (.Y(_08536_),
    .A(_08534_),
    .B(_08535_));
 sg13g2_nor2_1 _17632_ (.A(_08526_),
    .B(_08536_),
    .Y(_08537_));
 sg13g2_a21oi_1 _17633_ (.A1(_08498_),
    .A2(_08536_),
    .Y(_08538_),
    .B1(_08537_));
 sg13g2_nand2_1 _17634_ (.Y(_08539_),
    .A(_08130_),
    .B(_05841_));
 sg13g2_nand2_1 _17635_ (.Y(_08540_),
    .A(_05915_),
    .B(_05840_));
 sg13g2_nand3_1 _17636_ (.B(_08539_),
    .C(_08540_),
    .A(_08133_),
    .Y(_08541_));
 sg13g2_nand2_1 _17637_ (.Y(_08542_),
    .A(_08541_),
    .B(_08148_));
 sg13g2_nand2_1 _17638_ (.Y(_08543_),
    .A(_08542_),
    .B(_08150_));
 sg13g2_nand2_1 _17639_ (.Y(_08544_),
    .A(_08536_),
    .B(_08509_));
 sg13g2_o21ai_1 _17640_ (.B1(_08544_),
    .Y(_08545_),
    .A1(_08519_),
    .A2(_08536_));
 sg13g2_nand3_1 _17641_ (.B(net177),
    .C(_05133_),
    .A(_08129_),
    .Y(_08546_));
 sg13g2_nand3_1 _17642_ (.B(_05139_),
    .C(_08138_),
    .A(_08146_),
    .Y(_08547_));
 sg13g2_nor2_1 _17643_ (.A(_05439_),
    .B(_07975_),
    .Y(_08548_));
 sg13g2_inv_1 _17644_ (.Y(_08549_),
    .A(_08094_));
 sg13g2_nand3_1 _17645_ (.B(_08549_),
    .C(_08442_),
    .A(_08548_),
    .Y(_08550_));
 sg13g2_nor4_1 _17646_ (.A(_08104_),
    .B(_07969_),
    .C(_08550_),
    .D(_08074_),
    .Y(_08551_));
 sg13g2_o21ai_1 _17647_ (.B1(_05138_),
    .Y(_08552_),
    .A1(_05918_),
    .A2(_08551_));
 sg13g2_nand3_1 _17648_ (.B(net128),
    .C(_08552_),
    .A(_08547_),
    .Y(_08553_));
 sg13g2_o21ai_1 _17649_ (.B1(_05842_),
    .Y(_08554_),
    .A1(_05132_),
    .A2(_05129_));
 sg13g2_nand3_1 _17650_ (.B(net129),
    .C(_08554_),
    .A(_08131_),
    .Y(_08555_));
 sg13g2_nand3_1 _17651_ (.B(_08553_),
    .C(_08555_),
    .A(_08546_),
    .Y(_08556_));
 sg13g2_nand2_1 _17652_ (.Y(_08557_),
    .A(_08556_),
    .B(_08150_));
 sg13g2_inv_1 _17653_ (.Y(_08558_),
    .A(_08557_));
 sg13g2_nand2_1 _17654_ (.Y(_08559_),
    .A(_08545_),
    .B(_08558_));
 sg13g2_o21ai_1 _17655_ (.B1(_08559_),
    .Y(_08560_),
    .A1(_08543_),
    .A2(_08538_));
 sg13g2_nand2_1 _17656_ (.Y(_08561_),
    .A(_08538_),
    .B(_08543_));
 sg13g2_nor2b_1 _17657_ (.A(_08151_),
    .B_N(_08374_),
    .Y(_08562_));
 sg13g2_a21oi_1 _17658_ (.A1(_08560_),
    .A2(_08561_),
    .Y(_08563_),
    .B1(_08562_));
 sg13g2_nand2b_1 _17659_ (.Y(_08564_),
    .B(_08151_),
    .A_N(_08374_));
 sg13g2_nand2b_1 _17660_ (.Y(_08565_),
    .B(_08564_),
    .A_N(_08563_));
 sg13g2_buf_2 _17661_ (.A(_08565_),
    .X(_08566_));
 sg13g2_nor2_1 _17662_ (.A(_08543_),
    .B(_08566_),
    .Y(_08567_));
 sg13g2_a21o_1 _17663_ (.A2(_08566_),
    .A1(_08538_),
    .B1(_08567_),
    .X(_08568_));
 sg13g2_nand2_1 _17664_ (.Y(_08569_),
    .A(_08467_),
    .B(_05365_));
 sg13g2_nand2b_1 _17665_ (.Y(_08570_),
    .B(_05364_),
    .A_N(_05382_));
 sg13g2_nand3_1 _17666_ (.B(_08569_),
    .C(_08570_),
    .A(_08470_),
    .Y(_08571_));
 sg13g2_nand2_1 _17667_ (.Y(_08572_),
    .A(_08571_),
    .B(_08477_));
 sg13g2_nand2_1 _17668_ (.Y(_08573_),
    .A(_08572_),
    .B(_08479_));
 sg13g2_inv_1 _17669_ (.Y(_08574_),
    .A(_08573_));
 sg13g2_inv_1 _17670_ (.Y(_08575_),
    .A(_08568_));
 sg13g2_nand3_1 _17671_ (.B(net145),
    .C(_05369_),
    .A(_08466_),
    .Y(_08576_));
 sg13g2_nand3_1 _17672_ (.B(_05371_),
    .C(_08407_),
    .A(_08475_),
    .Y(_08577_));
 sg13g2_nor2_1 _17673_ (.A(_08448_),
    .B(_08464_),
    .Y(_08578_));
 sg13g2_nand4_1 _17674_ (.B(_05370_),
    .C(_08443_),
    .A(_08578_),
    .Y(_08579_),
    .D(_08446_));
 sg13g2_nor2_1 _17675_ (.A(net93),
    .B(_05372_),
    .Y(_08580_));
 sg13g2_nand3_1 _17676_ (.B(_08579_),
    .C(_08580_),
    .A(_08577_),
    .Y(_08581_));
 sg13g2_o21ai_1 _17677_ (.B1(_05366_),
    .Y(_08582_),
    .A1(_05363_),
    .A2(_05368_));
 sg13g2_nand3_1 _17678_ (.B(net96),
    .C(_08582_),
    .A(_08468_),
    .Y(_08583_));
 sg13g2_nand3_1 _17679_ (.B(_08581_),
    .C(_08583_),
    .A(_08576_),
    .Y(_08584_));
 sg13g2_nand2_1 _17680_ (.Y(_08585_),
    .A(_08584_),
    .B(_08479_));
 sg13g2_nor2_1 _17681_ (.A(_08558_),
    .B(_08566_),
    .Y(_08586_));
 sg13g2_a21oi_1 _17682_ (.A1(_08545_),
    .A2(_08566_),
    .Y(_08587_),
    .B1(_08586_));
 sg13g2_nor2_1 _17683_ (.A(_08585_),
    .B(_08587_),
    .Y(_08588_));
 sg13g2_o21ai_1 _17684_ (.B1(_08588_),
    .Y(_08589_),
    .A1(_08574_),
    .A2(_08575_));
 sg13g2_nand2_1 _17685_ (.Y(_08590_),
    .A(_08575_),
    .B(_08574_));
 sg13g2_xor2_1 _17686_ (.B(_08375_),
    .A(_08480_),
    .X(_08591_));
 sg13g2_nand3_1 _17687_ (.B(_08590_),
    .C(_08591_),
    .A(_08589_),
    .Y(_08592_));
 sg13g2_nand2_1 _17688_ (.Y(_08593_),
    .A(_08375_),
    .B(_08480_));
 sg13g2_nand2_2 _17689_ (.Y(_08594_),
    .A(_08592_),
    .B(_08593_));
 sg13g2_nor2_1 _17690_ (.A(_08573_),
    .B(_08594_),
    .Y(_08595_));
 sg13g2_a21oi_1 _17691_ (.A1(_08568_),
    .A2(_08594_),
    .Y(_08596_),
    .B1(_08595_));
 sg13g2_inv_2 _17692_ (.Y(_08597_),
    .A(_08596_));
 sg13g2_nand2_1 _17693_ (.Y(_08598_),
    .A(_08004_),
    .B(_08002_));
 sg13g2_nand2_1 _17694_ (.Y(_08599_),
    .A(_08004_),
    .B(_04915_));
 sg13g2_nand2b_1 _17695_ (.Y(_08600_),
    .B(_04914_),
    .A_N(_04932_));
 sg13g2_nand3_1 _17696_ (.B(_08599_),
    .C(_08600_),
    .A(_08598_),
    .Y(_08601_));
 sg13g2_a21o_1 _17697_ (.A2(_08011_),
    .A1(_08601_),
    .B1(_08012_),
    .X(_08602_));
 sg13g2_buf_1 _17698_ (.A(_08602_),
    .X(_08603_));
 sg13g2_nand2_1 _17699_ (.Y(_08604_),
    .A(_08597_),
    .B(_08603_));
 sg13g2_nand2_1 _17700_ (.Y(_08605_),
    .A(_08594_),
    .B(_08587_));
 sg13g2_o21ai_1 _17701_ (.B1(_08605_),
    .Y(_08606_),
    .A1(_08585_),
    .A2(_08594_));
 sg13g2_nand3_1 _17702_ (.B(_04921_),
    .C(_07892_),
    .A(_08009_),
    .Y(_08607_));
 sg13g2_inv_1 _17703_ (.Y(_08608_),
    .A(_07976_));
 sg13g2_nor4_1 _17704_ (.A(_04921_),
    .B(_07995_),
    .C(_08608_),
    .D(_07971_),
    .Y(_08609_));
 sg13g2_nor3_1 _17705_ (.A(_02089_),
    .B(_04922_),
    .C(_08609_),
    .Y(_08610_));
 sg13g2_o21ai_1 _17706_ (.B1(_04916_),
    .Y(_08611_),
    .A1(_04913_),
    .A2(net146));
 sg13g2_nand3_1 _17707_ (.B(_05088_),
    .C(_08611_),
    .A(_08001_),
    .Y(_08612_));
 sg13g2_o21ai_1 _17708_ (.B1(_08612_),
    .Y(_08613_),
    .A1(_04913_),
    .A2(_08004_));
 sg13g2_a21oi_1 _17709_ (.A1(_08607_),
    .A2(_08610_),
    .Y(_08614_),
    .B1(_08613_));
 sg13g2_nor2_1 _17710_ (.A(_08012_),
    .B(_08614_),
    .Y(_08615_));
 sg13g2_nor2b_1 _17711_ (.A(_08606_),
    .B_N(_08615_),
    .Y(_08616_));
 sg13g2_nand2_1 _17712_ (.Y(_08617_),
    .A(_08604_),
    .B(_08616_));
 sg13g2_nand2_1 _17713_ (.Y(_08618_),
    .A(_08481_),
    .B(_08013_));
 sg13g2_nand2b_1 _17714_ (.Y(_08619_),
    .B(_08596_),
    .A_N(_08603_));
 sg13g2_nand3_1 _17715_ (.B(_08618_),
    .C(_08619_),
    .A(_08617_),
    .Y(_08620_));
 sg13g2_nand2b_1 _17716_ (.Y(_08621_),
    .B(_08482_),
    .A_N(_08013_));
 sg13g2_nand2_2 _17717_ (.Y(_08622_),
    .A(_08620_),
    .B(_08621_));
 sg13g2_nor2_1 _17718_ (.A(_08603_),
    .B(_08622_),
    .Y(_08623_));
 sg13g2_a21oi_1 _17719_ (.A1(_08597_),
    .A2(_08622_),
    .Y(_08624_),
    .B1(_08623_));
 sg13g2_inv_2 _17720_ (.Y(_08625_),
    .A(_08624_));
 sg13g2_a22oi_1 _17721_ (.Y(_08626_),
    .B1(_07862_),
    .B2(_08625_),
    .A2(_08492_),
    .A1(_08484_));
 sg13g2_inv_2 _17722_ (.Y(_08627_),
    .A(_08622_));
 sg13g2_nand2_1 _17723_ (.Y(_08628_),
    .A(_08627_),
    .B(_08615_));
 sg13g2_nand3_1 _17724_ (.B(_05078_),
    .C(_04536_),
    .A(_07844_),
    .Y(_08629_));
 sg13g2_nor2b_1 _17725_ (.A(_07731_),
    .B_N(_07818_),
    .Y(_08630_));
 sg13g2_o21ai_1 _17726_ (.B1(_07959_),
    .Y(_08631_),
    .A1(_06698_),
    .A2(_08630_));
 sg13g2_nand3_1 _17727_ (.B(_04542_),
    .C(_08486_),
    .A(_07856_),
    .Y(_08632_));
 sg13g2_nand3_1 _17728_ (.B(net75),
    .C(_08632_),
    .A(_08631_),
    .Y(_08633_));
 sg13g2_o21ai_1 _17729_ (.B1(_06694_),
    .Y(_08634_),
    .A1(_04535_),
    .A2(net164));
 sg13g2_nand3_1 _17730_ (.B(net68),
    .C(_08634_),
    .A(_07846_),
    .Y(_08635_));
 sg13g2_nand3_1 _17731_ (.B(_08633_),
    .C(_08635_),
    .A(_08629_),
    .Y(_08636_));
 sg13g2_nor2b_1 _17732_ (.A(_07860_),
    .B_N(_08636_),
    .Y(_08637_));
 sg13g2_nand2_1 _17733_ (.Y(_08638_),
    .A(_08622_),
    .B(_08606_));
 sg13g2_nand3_1 _17734_ (.B(_08637_),
    .C(_08638_),
    .A(_08628_),
    .Y(_08639_));
 sg13g2_o21ai_1 _17735_ (.B1(_08639_),
    .Y(_08640_),
    .A1(_07862_),
    .A2(_08625_));
 sg13g2_nand2_1 _17736_ (.Y(_08641_),
    .A(_08626_),
    .B(_08640_));
 sg13g2_inv_1 _17737_ (.Y(_08642_),
    .A(_08492_));
 sg13g2_nand2_1 _17738_ (.Y(_08643_),
    .A(_08483_),
    .B(_08642_));
 sg13g2_nand2_2 _17739_ (.Y(_08644_),
    .A(_08641_),
    .B(_08643_));
 sg13g2_nor2_1 _17740_ (.A(_08625_),
    .B(_08644_),
    .Y(_08645_));
 sg13g2_a21oi_1 _17741_ (.A1(_07862_),
    .A2(_08644_),
    .Y(_08646_),
    .B1(_08645_));
 sg13g2_nor2_1 _17742_ (.A(net72),
    .B(_07717_),
    .Y(_08647_));
 sg13g2_a21oi_1 _17743_ (.A1(_06274_),
    .A2(_04699_),
    .Y(_08648_),
    .B1(_08020_));
 sg13g2_o21ai_1 _17744_ (.B1(_04948_),
    .Y(_08649_),
    .A1(_04127_),
    .A2(_08648_));
 sg13g2_nand3_1 _17745_ (.B(_06863_),
    .C(_05003_),
    .A(_08649_),
    .Y(_08650_));
 sg13g2_inv_1 _17746_ (.Y(_08651_),
    .A(_06352_));
 sg13g2_nor2b_1 _17747_ (.A(_06339_),
    .B_N(_06336_),
    .Y(_08652_));
 sg13g2_a21oi_1 _17748_ (.A1(_06338_),
    .A2(_08652_),
    .Y(_08653_),
    .B1(_06348_));
 sg13g2_o21ai_1 _17749_ (.B1(_06345_),
    .Y(_08654_),
    .A1(_08651_),
    .A2(_08653_));
 sg13g2_inv_1 _17750_ (.Y(_08655_),
    .A(_08654_));
 sg13g2_a21oi_2 _17751_ (.B1(_08166_),
    .Y(_08656_),
    .A2(net36),
    .A1(_08655_));
 sg13g2_o21ai_1 _17752_ (.B1(_05910_),
    .Y(_08657_),
    .A1(_05864_),
    .A2(_08656_));
 sg13g2_buf_1 _17753_ (.A(_08657_),
    .X(_08658_));
 sg13g2_a21oi_2 _17754_ (.B1(_06229_),
    .Y(_08659_),
    .A2(net27),
    .A1(_08658_));
 sg13g2_o21ai_1 _17755_ (.B1(_04110_),
    .Y(_08660_),
    .A1(_08650_),
    .A2(_08659_));
 sg13g2_nand2b_1 _17756_ (.Y(_08661_),
    .B(_06864_),
    .A_N(_08660_));
 sg13g2_inv_1 _17757_ (.Y(_08662_),
    .A(_07673_));
 sg13g2_a21oi_1 _17758_ (.A1(net60),
    .A2(_08662_),
    .Y(_08663_),
    .B1(_04346_));
 sg13g2_nor2_1 _17759_ (.A(_03916_),
    .B(_08663_),
    .Y(_08664_));
 sg13g2_nor3_1 _17760_ (.A(_06665_),
    .B(_06668_),
    .C(_06670_),
    .Y(_08665_));
 sg13g2_nand2_1 _17761_ (.Y(_08666_),
    .A(_06664_),
    .B(_08665_));
 sg13g2_inv_1 _17762_ (.Y(_08667_),
    .A(_08666_));
 sg13g2_a21oi_1 _17763_ (.A1(net69),
    .A2(_08667_),
    .Y(_08668_),
    .B1(_06681_));
 sg13g2_nor2_1 _17764_ (.A(_03601_),
    .B(_08668_),
    .Y(_08669_));
 sg13g2_nor4_1 _17765_ (.A(_08664_),
    .B(_07905_),
    .C(_08669_),
    .D(_05015_),
    .Y(_08670_));
 sg13g2_nor2_1 _17766_ (.A(_08040_),
    .B(_07902_),
    .Y(_08671_));
 sg13g2_nand2_1 _17767_ (.Y(_08672_),
    .A(_08670_),
    .B(_08671_));
 sg13g2_nor2_1 _17768_ (.A(_05057_),
    .B(_08663_),
    .Y(_08673_));
 sg13g2_or2_1 _17769_ (.X(_08674_),
    .B(_07936_),
    .A(_08106_));
 sg13g2_nor3_1 _17770_ (.A(_07930_),
    .B(_08673_),
    .C(_08674_),
    .Y(_08675_));
 sg13g2_nor2_2 _17771_ (.A(_06725_),
    .B(_08668_),
    .Y(_08676_));
 sg13g2_nor2_1 _17772_ (.A(_08676_),
    .B(_04528_),
    .Y(_08677_));
 sg13g2_nand2_1 _17773_ (.Y(_08678_),
    .A(_08675_),
    .B(_08677_));
 sg13g2_o21ai_1 _17774_ (.B1(_07158_),
    .Y(_08679_),
    .A1(_08672_),
    .A2(_08678_));
 sg13g2_nand2_1 _17775_ (.Y(_08680_),
    .A(_08661_),
    .B(_08679_));
 sg13g2_xnor2_1 _17776_ (.Y(_08681_),
    .A(_04099_),
    .B(_04317_));
 sg13g2_inv_1 _17777_ (.Y(_08682_),
    .A(_04226_));
 sg13g2_a21oi_1 _17778_ (.A1(_07780_),
    .A2(net50),
    .Y(_08683_),
    .B1(_07122_));
 sg13g2_a21oi_1 _17779_ (.A1(_07827_),
    .A2(net50),
    .Y(_08684_),
    .B1(_06731_));
 sg13g2_a22oi_1 _17780_ (.Y(_08685_),
    .B1(_08683_),
    .B2(_08684_),
    .A2(_04310_),
    .A1(_08682_));
 sg13g2_nor4_1 _17781_ (.A(_05062_),
    .B(_05006_),
    .C(_07801_),
    .D(_07993_),
    .Y(_08686_));
 sg13g2_inv_1 _17782_ (.Y(_08687_),
    .A(_08659_));
 sg13g2_a21oi_1 _17783_ (.A1(_06423_),
    .A2(net36),
    .Y(_08688_),
    .B1(_06808_));
 sg13g2_inv_1 _17784_ (.Y(_08689_),
    .A(_08688_));
 sg13g2_a21oi_1 _17785_ (.A1(_08689_),
    .A2(net22),
    .Y(_08690_),
    .B1(_05956_));
 sg13g2_inv_1 _17786_ (.Y(_08691_),
    .A(_08690_));
 sg13g2_a21oi_1 _17787_ (.A1(_08691_),
    .A2(_06186_),
    .Y(_08692_),
    .B1(_06189_));
 sg13g2_inv_1 _17788_ (.Y(_08693_),
    .A(_08692_));
 sg13g2_a21oi_1 _17789_ (.A1(_08687_),
    .A2(_07702_),
    .Y(_08694_),
    .B1(_08693_));
 sg13g2_inv_1 _17790_ (.Y(_08695_),
    .A(_04580_));
 sg13g2_nor2_1 _17791_ (.A(_07535_),
    .B(net32),
    .Y(_08696_));
 sg13g2_a21oi_1 _17792_ (.A1(_08695_),
    .A2(_08696_),
    .Y(_08697_),
    .B1(_04583_));
 sg13g2_buf_2 _17793_ (.A(_08697_),
    .X(_08698_));
 sg13g2_nor2_1 _17794_ (.A(_04985_),
    .B(_08698_),
    .Y(_08699_));
 sg13g2_inv_1 _17795_ (.Y(_08700_),
    .A(_04075_));
 sg13g2_a21oi_1 _17796_ (.A1(_08700_),
    .A2(_07527_),
    .Y(_08701_),
    .B1(_07526_));
 sg13g2_buf_2 _17797_ (.A(_08701_),
    .X(_08702_));
 sg13g2_nor2_1 _17798_ (.A(_04098_),
    .B(_08702_),
    .Y(_08703_));
 sg13g2_inv_1 _17799_ (.Y(_08704_),
    .A(_08703_));
 sg13g2_inv_1 _17800_ (.Y(_08705_),
    .A(_04098_));
 sg13g2_nand2_1 _17801_ (.Y(_08706_),
    .A(_08705_),
    .B(_06862_));
 sg13g2_nand2_1 _17802_ (.Y(_08707_),
    .A(_08704_),
    .B(_08706_));
 sg13g2_nor4_1 _17803_ (.A(_08699_),
    .B(_05004_),
    .C(_08707_),
    .D(_08672_),
    .Y(_08708_));
 sg13g2_inv_1 _17804_ (.Y(_08709_),
    .A(_07239_));
 sg13g2_a21oi_1 _17805_ (.A1(_08709_),
    .A2(_04248_),
    .Y(_08710_),
    .B1(_04251_));
 sg13g2_a21oi_1 _17806_ (.A1(_04496_),
    .A2(net98),
    .Y(_08711_),
    .B1(_05744_));
 sg13g2_inv_1 _17807_ (.Y(_08712_),
    .A(_08711_));
 sg13g2_a21oi_2 _17808_ (.B1(_04333_),
    .Y(_08713_),
    .A2(_04247_),
    .A1(_08712_));
 sg13g2_a22oi_1 _17809_ (.Y(_08714_),
    .B1(_08710_),
    .B2(_08713_),
    .A2(_07540_),
    .A1(_03760_));
 sg13g2_a21oi_1 _17810_ (.A1(_06444_),
    .A2(_04698_),
    .Y(_08715_),
    .B1(_04702_));
 sg13g2_inv_1 _17811_ (.Y(_08716_),
    .A(_08715_));
 sg13g2_a21oi_1 _17812_ (.A1(_08716_),
    .A2(net71),
    .Y(_08717_),
    .B1(_04131_));
 sg13g2_inv_1 _17813_ (.Y(_08718_),
    .A(_08649_));
 sg13g2_nand2_1 _17814_ (.Y(_08719_),
    .A(_08717_),
    .B(_08718_));
 sg13g2_nand4_1 _17815_ (.B(_05055_),
    .C(_08714_),
    .A(_08708_),
    .Y(_08720_),
    .D(_08719_));
 sg13g2_nor2_1 _17816_ (.A(_08694_),
    .B(_08720_),
    .Y(_08721_));
 sg13g2_nand3_1 _17817_ (.B(_08686_),
    .C(_08721_),
    .A(_08685_),
    .Y(_08722_));
 sg13g2_inv_1 _17818_ (.Y(_08723_),
    .A(_08717_));
 sg13g2_a22oi_1 _17819_ (.Y(_08724_),
    .B1(_08659_),
    .B2(_08693_),
    .A2(_08718_),
    .A1(_08723_));
 sg13g2_inv_1 _17820_ (.Y(_08725_),
    .A(_08710_));
 sg13g2_a22oi_1 _17821_ (.Y(_08726_),
    .B1(_08713_),
    .B2(_08725_),
    .A2(_07540_),
    .A1(_04985_));
 sg13g2_o21ai_1 _17822_ (.B1(_08726_),
    .Y(_08727_),
    .A1(_04311_),
    .A2(_08682_));
 sg13g2_inv_1 _17823_ (.Y(_08728_),
    .A(_08727_));
 sg13g2_nand2_1 _17824_ (.Y(_08729_),
    .A(_08724_),
    .B(_08728_));
 sg13g2_inv_1 _17825_ (.Y(_08730_),
    .A(_08684_));
 sg13g2_nand2_1 _17826_ (.Y(_08731_),
    .A(_08730_),
    .B(_08683_));
 sg13g2_inv_1 _17827_ (.Y(_08732_),
    .A(_07704_));
 sg13g2_inv_1 _17828_ (.Y(_08733_),
    .A(_04985_));
 sg13g2_nor2_1 _17829_ (.A(_08698_),
    .B(_08733_),
    .Y(_08734_));
 sg13g2_nand3b_1 _17830_ (.B(_04488_),
    .C(_08677_),
    .Y(_08735_),
    .A_N(_08734_));
 sg13g2_nand2_1 _17831_ (.Y(_08736_),
    .A(_06862_),
    .B(_04098_));
 sg13g2_nor2_2 _17832_ (.A(_08702_),
    .B(_08705_),
    .Y(_08737_));
 sg13g2_inv_1 _17833_ (.Y(_08738_),
    .A(_08737_));
 sg13g2_nand3_1 _17834_ (.B(_08736_),
    .C(_08738_),
    .A(_08675_),
    .Y(_08739_));
 sg13g2_nor3_1 _17835_ (.A(_04988_),
    .B(_08735_),
    .C(_08739_),
    .Y(_08740_));
 sg13g2_nor2_1 _17836_ (.A(_07724_),
    .B(_04134_),
    .Y(_08741_));
 sg13g2_nand4_1 _17837_ (.B(_08732_),
    .C(_08740_),
    .A(_08731_),
    .Y(_08742_),
    .D(_08741_));
 sg13g2_nor4_1 _17838_ (.A(net14),
    .B(_04408_),
    .C(_08729_),
    .D(_08742_),
    .Y(_08743_));
 sg13g2_nor2b_1 _17839_ (.A(_08722_),
    .B_N(_08743_),
    .Y(_08744_));
 sg13g2_nand2_1 _17840_ (.Y(_08745_),
    .A(_04312_),
    .B(net68));
 sg13g2_nor2_1 _17841_ (.A(_04110_),
    .B(_08743_),
    .Y(_08746_));
 sg13g2_nand3_1 _17842_ (.B(net114),
    .C(_08722_),
    .A(_08746_),
    .Y(_08747_));
 sg13g2_buf_1 _17843_ (.A(_08747_),
    .X(_08748_));
 sg13g2_o21ai_1 _17844_ (.B1(_08748_),
    .Y(_08749_),
    .A1(_08744_),
    .A2(_08745_));
 sg13g2_a22oi_1 _17845_ (.Y(_08750_),
    .B1(_08681_),
    .B2(_08749_),
    .A2(_08680_),
    .A1(_08647_));
 sg13g2_nand4_1 _17846_ (.B(_08731_),
    .C(_08714_),
    .A(_08685_),
    .Y(_08751_),
    .D(_08728_));
 sg13g2_nand2_1 _17847_ (.Y(_08752_),
    .A(_08751_),
    .B(_04110_));
 sg13g2_a21o_1 _17848_ (.A2(_08660_),
    .A1(_08752_),
    .B1(_04318_),
    .X(_08753_));
 sg13g2_o21ai_1 _17849_ (.B1(_08753_),
    .Y(_08754_),
    .A1(_04316_),
    .A2(_08752_));
 sg13g2_nand2_1 _17850_ (.Y(_08755_),
    .A(_08754_),
    .B(net67));
 sg13g2_nand2_1 _17851_ (.Y(_08756_),
    .A(_08750_),
    .B(_08755_));
 sg13g2_buf_1 _17852_ (.A(\b.gen_square[38].sq.mask ),
    .X(_08757_));
 sg13g2_nand2_1 _17853_ (.Y(_08758_),
    .A(_08756_),
    .B(_08757_));
 sg13g2_nor2_1 _17854_ (.A(_08642_),
    .B(_08484_),
    .Y(_08759_));
 sg13g2_inv_1 _17855_ (.Y(_08760_),
    .A(_08759_));
 sg13g2_nor2_1 _17856_ (.A(_08758_),
    .B(_08760_),
    .Y(_08761_));
 sg13g2_inv_1 _17857_ (.Y(_08762_),
    .A(_08761_));
 sg13g2_nand2_1 _17858_ (.Y(_08763_),
    .A(_08760_),
    .B(_08758_));
 sg13g2_nand2_1 _17859_ (.Y(_08764_),
    .A(_08762_),
    .B(_08763_));
 sg13g2_a21oi_1 _17860_ (.A1(_08628_),
    .A2(_08638_),
    .Y(_08765_),
    .B1(_08644_));
 sg13g2_a21o_1 _17861_ (.A2(_08644_),
    .A1(_08637_),
    .B1(_08765_),
    .X(_08766_));
 sg13g2_inv_1 _17862_ (.Y(_08767_),
    .A(_04102_));
 sg13g2_a21oi_1 _17863_ (.A1(_04312_),
    .A2(_08767_),
    .Y(_08768_),
    .B1(_04104_));
 sg13g2_nor3_1 _17864_ (.A(net142),
    .B(_08768_),
    .C(_08744_),
    .Y(_08769_));
 sg13g2_nand3_1 _17865_ (.B(_04108_),
    .C(_08661_),
    .A(_08753_),
    .Y(_08770_));
 sg13g2_nor2_1 _17866_ (.A(_04408_),
    .B(net14),
    .Y(_08771_));
 sg13g2_nand4_1 _17867_ (.B(_08698_),
    .C(_08702_),
    .A(_07702_),
    .Y(_08772_),
    .D(_07717_));
 sg13g2_nor3_1 _17868_ (.A(_04988_),
    .B(_08772_),
    .C(_05054_),
    .Y(_08773_));
 sg13g2_nand4_1 _17869_ (.B(_08741_),
    .C(_08771_),
    .A(_08686_),
    .Y(_08774_),
    .D(_08773_));
 sg13g2_nor2_1 _17870_ (.A(net63),
    .B(_04111_),
    .Y(_08775_));
 sg13g2_nand3_1 _17871_ (.B(_08774_),
    .C(_08775_),
    .A(_08770_),
    .Y(_08776_));
 sg13g2_o21ai_1 _17872_ (.B1(_08776_),
    .Y(_08777_),
    .A1(_04102_),
    .A2(_08748_));
 sg13g2_o21ai_1 _17873_ (.B1(_08757_),
    .Y(_08778_),
    .A1(_08769_),
    .A2(_08777_));
 sg13g2_inv_1 _17874_ (.Y(_08779_),
    .A(_04317_));
 sg13g2_a22oi_1 _17875_ (.Y(_08780_),
    .B1(_04104_),
    .B2(_08748_),
    .A2(_04103_),
    .A1(_08779_));
 sg13g2_a22oi_1 _17876_ (.Y(_08781_),
    .B1(_08749_),
    .B2(_08780_),
    .A2(_08754_),
    .A1(_05115_));
 sg13g2_nand2b_1 _17877_ (.Y(_08782_),
    .B(_08757_),
    .A_N(_08781_));
 sg13g2_xnor2_1 _17878_ (.Y(_08783_),
    .A(_08782_),
    .B(_08646_));
 sg13g2_or4_1 _17879_ (.A(_08764_),
    .B(_08766_),
    .C(_08778_),
    .D(_08783_),
    .X(_08784_));
 sg13g2_nor2_1 _17880_ (.A(_08782_),
    .B(_08646_),
    .Y(_08785_));
 sg13g2_a21oi_1 _17881_ (.A1(_08785_),
    .A2(_08763_),
    .Y(_08786_),
    .B1(_08761_));
 sg13g2_nand2_2 _17882_ (.Y(_08787_),
    .A(_08784_),
    .B(_08786_));
 sg13g2_inv_4 _17883_ (.A(_08787_),
    .Y(_08788_));
 sg13g2_nand2b_1 _17884_ (.Y(_08789_),
    .B(_08788_),
    .A_N(_08646_));
 sg13g2_nand2_1 _17885_ (.Y(_08790_),
    .A(_08787_),
    .B(_08782_));
 sg13g2_nand2_1 _17886_ (.Y(_08791_),
    .A(_08789_),
    .B(_08790_));
 sg13g2_inv_1 _17887_ (.Y(_08792_),
    .A(_08791_));
 sg13g2_nor3_1 _17888_ (.A(_06531_),
    .B(_06533_),
    .C(_06544_),
    .Y(_08793_));
 sg13g2_o21ai_1 _17889_ (.B1(net115),
    .Y(_08794_),
    .A1(_08793_),
    .A2(_06536_));
 sg13g2_o21ai_1 _17890_ (.B1(_06549_),
    .Y(_08795_),
    .A1(_06541_),
    .A2(_08794_));
 sg13g2_inv_1 _17891_ (.Y(_08796_),
    .A(_08795_));
 sg13g2_a21oi_1 _17892_ (.A1(_08796_),
    .A2(net49),
    .Y(_08797_),
    .B1(_08286_));
 sg13g2_inv_1 _17893_ (.Y(_08798_),
    .A(_08797_));
 sg13g2_inv_1 _17894_ (.Y(_08799_),
    .A(_05327_));
 sg13g2_a21oi_1 _17895_ (.A1(_08798_),
    .A2(_07100_),
    .Y(_08800_),
    .B1(_08799_));
 sg13g2_inv_1 _17896_ (.Y(_08801_),
    .A(_08800_));
 sg13g2_a21oi_1 _17897_ (.A1(_08801_),
    .A2(net33),
    .Y(_08802_),
    .B1(_06688_));
 sg13g2_inv_1 _17898_ (.Y(_08803_),
    .A(_08802_));
 sg13g2_a21oi_1 _17899_ (.A1(_06805_),
    .A2(net65),
    .Y(_08804_),
    .B1(_07002_));
 sg13g2_inv_1 _17900_ (.Y(_08805_),
    .A(_08804_));
 sg13g2_a21oi_1 _17901_ (.A1(_08805_),
    .A2(net25),
    .Y(_08806_),
    .B1(_05527_));
 sg13g2_inv_1 _17902_ (.Y(_08807_),
    .A(_08806_));
 sg13g2_a21oi_1 _17903_ (.A1(_08807_),
    .A2(_04154_),
    .Y(_08808_),
    .B1(_04224_));
 sg13g2_nor2b_1 _17904_ (.A(_08803_),
    .B_N(_08808_),
    .Y(_08809_));
 sg13g2_nand2b_1 _17905_ (.Y(_08810_),
    .B(_07497_),
    .A_N(_08702_));
 sg13g2_nor2_1 _17906_ (.A(_05062_),
    .B(_07612_),
    .Y(_08811_));
 sg13g2_inv_1 _17907_ (.Y(_08812_),
    .A(_07812_));
 sg13g2_inv_1 _17908_ (.Y(_08813_),
    .A(_07801_));
 sg13g2_nand4_1 _17909_ (.B(_08811_),
    .C(_08812_),
    .A(_08810_),
    .Y(_08814_),
    .D(_08813_));
 sg13g2_inv_1 _17910_ (.Y(_08815_),
    .A(_08388_));
 sg13g2_a21oi_1 _17911_ (.A1(_06766_),
    .A2(net77),
    .Y(_08816_),
    .B1(_08815_));
 sg13g2_inv_1 _17912_ (.Y(_08817_),
    .A(_08816_));
 sg13g2_a21oi_1 _17913_ (.A1(_08817_),
    .A2(_04248_),
    .Y(_08818_),
    .B1(_07231_));
 sg13g2_inv_1 _17914_ (.Y(_08819_),
    .A(_08818_));
 sg13g2_o21ai_1 _17915_ (.B1(_04250_),
    .Y(_08820_),
    .A1(_04249_),
    .A2(_04998_));
 sg13g2_nor2_1 _17916_ (.A(_07837_),
    .B(_06650_),
    .Y(_08821_));
 sg13g2_inv_1 _17917_ (.Y(_08822_),
    .A(_08821_));
 sg13g2_nor3_1 _17918_ (.A(_07831_),
    .B(_08422_),
    .C(_08822_),
    .Y(_08823_));
 sg13g2_o21ai_1 _17919_ (.B1(_08823_),
    .Y(_08824_),
    .A1(_08819_),
    .A2(_08820_));
 sg13g2_a21oi_1 _17920_ (.A1(_08730_),
    .A2(net34),
    .Y(_08825_),
    .B1(_04120_));
 sg13g2_inv_1 _17921_ (.Y(_08826_),
    .A(_08683_));
 sg13g2_a21oi_1 _17922_ (.A1(_08826_),
    .A2(net34),
    .Y(_08827_),
    .B1(_04321_));
 sg13g2_inv_1 _17923_ (.Y(_08828_),
    .A(_04438_));
 sg13g2_nor2_1 _17924_ (.A(_04436_),
    .B(_04357_),
    .Y(_08829_));
 sg13g2_a21oi_1 _17925_ (.A1(_07557_),
    .A2(_08828_),
    .Y(_08830_),
    .B1(_08829_));
 sg13g2_inv_1 _17926_ (.Y(_08831_),
    .A(_08830_));
 sg13g2_a21oi_1 _17927_ (.A1(_08831_),
    .A2(_04406_),
    .Y(_08832_),
    .B1(_07549_));
 sg13g2_inv_1 _17928_ (.Y(_08833_),
    .A(_08832_));
 sg13g2_nand2_1 _17929_ (.Y(_08834_),
    .A(_07534_),
    .B(_07497_));
 sg13g2_o21ai_1 _17930_ (.B1(_08834_),
    .Y(_08835_),
    .A1(_07611_),
    .A2(_08833_));
 sg13g2_a21oi_1 _17931_ (.A1(_08825_),
    .A2(_08827_),
    .Y(_08836_),
    .B1(_08835_));
 sg13g2_inv_1 _17932_ (.Y(_08837_),
    .A(_08836_));
 sg13g2_nor4_1 _17933_ (.A(_08809_),
    .B(_08814_),
    .C(_08824_),
    .D(_08837_),
    .Y(_08838_));
 sg13g2_nor2_1 _17934_ (.A(_08803_),
    .B(_08808_),
    .Y(_08839_));
 sg13g2_nor2_1 _17935_ (.A(_08702_),
    .B(_07497_),
    .Y(_08840_));
 sg13g2_nor2_1 _17936_ (.A(_07571_),
    .B(_08840_),
    .Y(_08841_));
 sg13g2_inv_1 _17937_ (.Y(_08842_),
    .A(_07724_));
 sg13g2_nand3_1 _17938_ (.B(_07721_),
    .C(_08842_),
    .A(_08841_),
    .Y(_08843_));
 sg13g2_nor2_1 _17939_ (.A(_07570_),
    .B(_08833_),
    .Y(_08844_));
 sg13g2_o21ai_1 _17940_ (.B1(_08820_),
    .Y(_08845_),
    .A1(_07653_),
    .A2(_08818_));
 sg13g2_nor4_2 _17941_ (.A(_07737_),
    .B(_07747_),
    .C(_06625_),
    .Y(_08846_),
    .D(_08413_));
 sg13g2_nand3b_1 _17942_ (.B(_08845_),
    .C(_08846_),
    .Y(_08847_),
    .A_N(_08844_));
 sg13g2_inv_1 _17943_ (.Y(_08848_),
    .A(_07534_));
 sg13g2_nand2b_1 _17944_ (.Y(_08849_),
    .B(_08827_),
    .A_N(_08825_));
 sg13g2_o21ai_1 _17945_ (.B1(_08849_),
    .Y(_08850_),
    .A1(_07497_),
    .A2(_08848_));
 sg13g2_nor4_1 _17946_ (.A(_08839_),
    .B(_08843_),
    .C(_08847_),
    .D(_08850_),
    .Y(_08851_));
 sg13g2_nor3_1 _17947_ (.A(_04570_),
    .B(_08838_),
    .C(_08851_),
    .Y(_08852_));
 sg13g2_nand2_1 _17948_ (.Y(_08853_),
    .A(_08852_),
    .B(net114));
 sg13g2_nand2_1 _17949_ (.Y(_08854_),
    .A(_08851_),
    .B(_08838_));
 sg13g2_nand3_1 _17950_ (.B(net57),
    .C(_07535_),
    .A(_08854_),
    .Y(_08855_));
 sg13g2_nand2_1 _17951_ (.Y(_08856_),
    .A(_08853_),
    .B(_08855_));
 sg13g2_nand2_1 _17952_ (.Y(_08857_),
    .A(_08853_),
    .B(_04982_));
 sg13g2_nand2_1 _17953_ (.Y(_08858_),
    .A(_07219_),
    .B(_04981_));
 sg13g2_nand3_1 _17954_ (.B(_08857_),
    .C(_08858_),
    .A(_08856_),
    .Y(_08859_));
 sg13g2_a21oi_1 _17955_ (.A1(_08803_),
    .A2(_08819_),
    .Y(_08860_),
    .B1(_07535_));
 sg13g2_nor3_1 _17956_ (.A(_08844_),
    .B(_08837_),
    .C(_08850_),
    .Y(_08861_));
 sg13g2_nor2_1 _17957_ (.A(_07535_),
    .B(_08861_),
    .Y(_08862_));
 sg13g2_o21ai_1 _17958_ (.B1(_07220_),
    .Y(_08863_),
    .A1(_08860_),
    .A2(_08862_));
 sg13g2_nand3_1 _17959_ (.B(_04980_),
    .C(_07536_),
    .A(_08862_),
    .Y(_08864_));
 sg13g2_nand2_1 _17960_ (.Y(_08865_),
    .A(_08863_),
    .B(_08864_));
 sg13g2_nand2_1 _17961_ (.Y(_08866_),
    .A(_08865_),
    .B(_05115_));
 sg13g2_nand2_1 _17962_ (.Y(_08867_),
    .A(_08859_),
    .B(_08866_));
 sg13g2_buf_1 _17963_ (.A(\b.gen_square[39].sq.mask ),
    .X(_08868_));
 sg13g2_nand2_1 _17964_ (.Y(_08869_),
    .A(_08867_),
    .B(_08868_));
 sg13g2_inv_1 _17965_ (.Y(_08870_),
    .A(_08869_));
 sg13g2_nand2b_1 _17966_ (.Y(_08871_),
    .B(_08788_),
    .A_N(_08766_));
 sg13g2_nand2_1 _17967_ (.Y(_08872_),
    .A(_08787_),
    .B(_08778_));
 sg13g2_nor2b_1 _17968_ (.A(_07222_),
    .B_N(_08860_),
    .Y(_08873_));
 sg13g2_nand3b_1 _17969_ (.B(_08863_),
    .C(_04580_),
    .Y(_08874_),
    .A_N(_08873_));
 sg13g2_nor3_1 _17970_ (.A(_04988_),
    .B(_08843_),
    .C(_08814_),
    .Y(_08875_));
 sg13g2_o21ai_1 _17971_ (.B1(_08695_),
    .Y(_08876_),
    .A1(_07535_),
    .A2(_08875_));
 sg13g2_nand3_1 _17972_ (.B(_05116_),
    .C(_08876_),
    .A(_08874_),
    .Y(_08877_));
 sg13g2_inv_1 _17973_ (.Y(_08878_),
    .A(_04982_));
 sg13g2_nand2_1 _17974_ (.Y(_08879_),
    .A(_08878_),
    .B(_04570_));
 sg13g2_nand3_1 _17975_ (.B(_05091_),
    .C(_08879_),
    .A(_08854_),
    .Y(_08880_));
 sg13g2_a21o_1 _17976_ (.A2(_08878_),
    .A1(_04573_),
    .B1(_08880_),
    .X(_08881_));
 sg13g2_nand3_1 _17977_ (.B(_05079_),
    .C(_04574_),
    .A(_08852_),
    .Y(_08882_));
 sg13g2_nand3_1 _17978_ (.B(_08881_),
    .C(_08882_),
    .A(_08877_),
    .Y(_08883_));
 sg13g2_nand2_1 _17979_ (.Y(_08884_),
    .A(_08883_),
    .B(_08868_));
 sg13g2_a21oi_1 _17980_ (.A1(_08871_),
    .A2(_08872_),
    .Y(_08885_),
    .B1(_08884_));
 sg13g2_o21ai_1 _17981_ (.B1(_08885_),
    .Y(_08886_),
    .A1(_08791_),
    .A2(_08870_));
 sg13g2_a21oi_1 _17982_ (.A1(_08823_),
    .A2(_08846_),
    .Y(_08887_),
    .B1(_04576_));
 sg13g2_nor3_1 _17983_ (.A(_08873_),
    .B(_08887_),
    .C(_08865_),
    .Y(_08888_));
 sg13g2_nor2_1 _17984_ (.A(_04571_),
    .B(_07218_),
    .Y(_08889_));
 sg13g2_o21ai_1 _17985_ (.B1(_08856_),
    .Y(_08890_),
    .A1(_07220_),
    .A2(_08889_));
 sg13g2_o21ai_1 _17986_ (.B1(_08890_),
    .Y(_08891_),
    .A1(net48),
    .A2(_08888_));
 sg13g2_nand2_1 _17987_ (.Y(_08892_),
    .A(_08891_),
    .B(_08868_));
 sg13g2_nand2_1 _17988_ (.Y(_08893_),
    .A(_08759_),
    .B(_08758_));
 sg13g2_nor2_1 _17989_ (.A(_08892_),
    .B(_08893_),
    .Y(_08894_));
 sg13g2_a21oi_1 _17990_ (.A1(_08791_),
    .A2(_08870_),
    .Y(_08895_),
    .B1(_08894_));
 sg13g2_nand2_1 _17991_ (.Y(_08896_),
    .A(_08886_),
    .B(_08895_));
 sg13g2_nand2_1 _17992_ (.Y(_08897_),
    .A(_08893_),
    .B(_08892_));
 sg13g2_nand2_2 _17993_ (.Y(_08898_),
    .A(_08896_),
    .B(_08897_));
 sg13g2_nor2_1 _17994_ (.A(_08869_),
    .B(_08898_),
    .Y(_08899_));
 sg13g2_a21oi_2 _17995_ (.B1(_08899_),
    .Y(_08900_),
    .A2(_08898_),
    .A1(_08792_));
 sg13g2_inv_1 _17996_ (.Y(_08901_),
    .A(_06333_));
 sg13g2_a21oi_2 _17997_ (.B1(_05616_),
    .Y(_08902_),
    .A2(_04835_),
    .A1(_06008_));
 sg13g2_o21ai_1 _17998_ (.B1(_06362_),
    .Y(_08903_),
    .A1(_08901_),
    .A2(_08902_));
 sg13g2_a21oi_1 _17999_ (.A1(_08903_),
    .A2(net36),
    .Y(_08904_),
    .B1(_06560_));
 sg13g2_inv_1 _18000_ (.Y(_08905_),
    .A(_08904_));
 sg13g2_a21oi_1 _18001_ (.A1(_08905_),
    .A2(net49),
    .Y(_08906_),
    .B1(_06964_));
 sg13g2_inv_1 _18002_ (.Y(_08907_),
    .A(_08906_));
 sg13g2_a21oi_1 _18003_ (.A1(_08907_),
    .A2(net64),
    .Y(_08908_),
    .B1(_07097_));
 sg13g2_inv_2 _18004_ (.Y(_08909_),
    .A(_06529_));
 sg13g2_a21oi_1 _18005_ (.A1(_07180_),
    .A2(_04835_),
    .Y(_08910_),
    .B1(_04956_));
 sg13g2_inv_1 _18006_ (.Y(_08911_),
    .A(_08910_));
 sg13g2_a21oi_1 _18007_ (.A1(_08911_),
    .A2(net37),
    .Y(_08912_),
    .B1(_06426_));
 sg13g2_inv_1 _18008_ (.Y(_08913_),
    .A(_06808_));
 sg13g2_o21ai_1 _18009_ (.B1(_08913_),
    .Y(_08914_),
    .A1(_08909_),
    .A2(_08912_));
 sg13g2_a21oi_1 _18010_ (.A1(_08914_),
    .A2(net49),
    .Y(_08915_),
    .B1(_07002_));
 sg13g2_inv_1 _18011_ (.Y(_08916_),
    .A(_08915_));
 sg13g2_a21oi_1 _18012_ (.A1(_08916_),
    .A2(net64),
    .Y(_08917_),
    .B1(_05950_));
 sg13g2_a22oi_1 _18013_ (.Y(_08918_),
    .B1(_08908_),
    .B2(_08917_),
    .A2(_04269_),
    .A1(_04001_));
 sg13g2_inv_1 _18014_ (.Y(_08919_),
    .A(_08713_));
 sg13g2_a21oi_1 _18015_ (.A1(_08919_),
    .A2(_04116_),
    .Y(_08920_),
    .B1(_04321_));
 sg13g2_inv_1 _18016_ (.Y(_08921_),
    .A(_08920_));
 sg13g2_a21oi_1 _18017_ (.A1(_08921_),
    .A2(_04153_),
    .Y(_08922_),
    .B1(_04309_));
 sg13g2_inv_1 _18018_ (.Y(_08923_),
    .A(_08922_));
 sg13g2_a21oi_1 _18019_ (.A1(_08923_),
    .A2(net62),
    .Y(_08924_),
    .B1(_04295_));
 sg13g2_a21oi_2 _18020_ (.B1(_04120_),
    .Y(_08925_),
    .A2(_04116_),
    .A1(_08725_));
 sg13g2_inv_1 _18021_ (.Y(_08926_),
    .A(_08925_));
 sg13g2_a21oi_1 _18022_ (.A1(_08926_),
    .A2(net33),
    .Y(_08927_),
    .B1(_04224_));
 sg13g2_inv_1 _18023_ (.Y(_08928_),
    .A(_08927_));
 sg13g2_a21oi_1 _18024_ (.A1(_08928_),
    .A2(net47),
    .Y(_08929_),
    .B1(_04220_));
 sg13g2_a22oi_1 _18025_ (.Y(_08930_),
    .B1(_08924_),
    .B2(_08929_),
    .A2(_07514_),
    .A1(_03221_));
 sg13g2_nand2_1 _18026_ (.Y(_08931_),
    .A(_08918_),
    .B(_08930_));
 sg13g2_inv_1 _18027_ (.Y(_08932_),
    .A(_05882_));
 sg13g2_a21oi_2 _18028_ (.B1(_05888_),
    .Y(_08933_),
    .A2(_05892_),
    .A1(_08932_));
 sg13g2_nor2_2 _18029_ (.A(_08933_),
    .B(_05952_),
    .Y(_08934_));
 sg13g2_inv_1 _18030_ (.Y(_08935_),
    .A(_08934_));
 sg13g2_inv_1 _18031_ (.Y(_08936_),
    .A(_04209_));
 sg13g2_a21oi_1 _18032_ (.A1(_08936_),
    .A2(_04288_),
    .Y(_08937_),
    .B1(_04214_));
 sg13g2_buf_2 _18033_ (.A(_08937_),
    .X(_08938_));
 sg13g2_nor2_1 _18034_ (.A(_08938_),
    .B(_06169_),
    .Y(_08939_));
 sg13g2_buf_1 _18035_ (.A(_08939_),
    .X(_08940_));
 sg13g2_inv_1 _18036_ (.Y(_08941_),
    .A(_08940_));
 sg13g2_inv_1 _18037_ (.Y(_08942_),
    .A(_06677_));
 sg13g2_a21oi_1 _18038_ (.A1(_08942_),
    .A2(_07520_),
    .Y(_08943_),
    .B1(_06681_));
 sg13g2_buf_2 _18039_ (.A(_08943_),
    .X(_08944_));
 sg13g2_nor2_1 _18040_ (.A(_08944_),
    .B(_06727_),
    .Y(_08945_));
 sg13g2_inv_1 _18041_ (.Y(_08946_),
    .A(_06156_));
 sg13g2_a21oi_1 _18042_ (.A1(_08946_),
    .A2(_06210_),
    .Y(_08947_),
    .B1(_06211_));
 sg13g2_buf_1 _18043_ (.A(_08947_),
    .X(_08948_));
 sg13g2_nor3_1 _18044_ (.A(_03231_),
    .B(_07505_),
    .C(_08948_),
    .Y(_08949_));
 sg13g2_nor2_1 _18045_ (.A(_08945_),
    .B(_08949_),
    .Y(_08950_));
 sg13g2_nand3_1 _18046_ (.B(_08941_),
    .C(_08950_),
    .A(_08935_),
    .Y(_08951_));
 sg13g2_a21oi_1 _18047_ (.A1(_08384_),
    .A2(net54),
    .Y(_08952_),
    .B1(_05387_));
 sg13g2_inv_1 _18048_ (.Y(_08953_),
    .A(_08952_));
 sg13g2_a21oi_1 _18049_ (.A1(_08953_),
    .A2(net40),
    .Y(_08954_),
    .B1(_05357_));
 sg13g2_inv_1 _18050_ (.Y(_08955_),
    .A(_08954_));
 sg13g2_a21oi_1 _18051_ (.A1(_08955_),
    .A2(_07100_),
    .Y(_08956_),
    .B1(_08799_));
 sg13g2_inv_1 _18052_ (.Y(_08957_),
    .A(_08956_));
 sg13g2_a21oi_2 _18053_ (.B1(_05287_),
    .Y(_08958_),
    .A2(_05320_),
    .A1(_05282_));
 sg13g2_nand2_1 _18054_ (.Y(_08959_),
    .A(_08957_),
    .B(_08958_));
 sg13g2_inv_1 _18055_ (.Y(_08960_),
    .A(_07974_));
 sg13g2_a21oi_1 _18056_ (.A1(_08960_),
    .A2(_05347_),
    .Y(_08961_),
    .B1(_05532_));
 sg13g2_inv_1 _18057_ (.Y(_08962_),
    .A(_08961_));
 sg13g2_a21oi_1 _18058_ (.A1(_08962_),
    .A2(net25),
    .Y(_08963_),
    .B1(_05527_));
 sg13g2_nand2_1 _18059_ (.Y(_08964_),
    .A(_08959_),
    .B(_08963_));
 sg13g2_nand2_1 _18060_ (.Y(_08965_),
    .A(_05520_),
    .B(_04009_));
 sg13g2_inv_1 _18061_ (.Y(_08966_),
    .A(_08965_));
 sg13g2_nor2_1 _18062_ (.A(_06683_),
    .B(_06727_),
    .Y(_08967_));
 sg13g2_a21oi_1 _18063_ (.A1(_05311_),
    .A2(_08966_),
    .Y(_08968_),
    .B1(_08967_));
 sg13g2_nor4_1 _18064_ (.A(_06918_),
    .B(_06917_),
    .C(_06921_),
    .D(_06932_),
    .Y(_08969_));
 sg13g2_a21o_1 _18065_ (.A2(_08969_),
    .A1(net115),
    .B1(_06994_),
    .X(_08970_));
 sg13g2_buf_1 _18066_ (.A(_08970_),
    .X(_08971_));
 sg13g2_a21oi_1 _18067_ (.A1(_08971_),
    .A2(_03870_),
    .Y(_08972_),
    .B1(_07838_));
 sg13g2_nor2_1 _18068_ (.A(_07834_),
    .B(_08422_),
    .Y(_08973_));
 sg13g2_nand2_1 _18069_ (.Y(_08974_),
    .A(_08972_),
    .B(_08973_));
 sg13g2_inv_1 _18070_ (.Y(_08975_),
    .A(_08974_));
 sg13g2_o21ai_1 _18071_ (.B1(_05310_),
    .Y(_08976_),
    .A1(_05305_),
    .A2(_05303_));
 sg13g2_inv_1 _18072_ (.Y(_08977_),
    .A(_08976_));
 sg13g2_nor2_1 _18073_ (.A(_08965_),
    .B(_08977_),
    .Y(_08978_));
 sg13g2_o21ai_1 _18074_ (.B1(_04258_),
    .Y(_08979_),
    .A1(_04165_),
    .A2(_05867_));
 sg13g2_buf_1 _18075_ (.A(_08979_),
    .X(_08980_));
 sg13g2_inv_1 _18076_ (.Y(_08981_),
    .A(_08980_));
 sg13g2_nor2_1 _18077_ (.A(_04176_),
    .B(_08981_),
    .Y(_08982_));
 sg13g2_inv_1 _18078_ (.Y(_08983_),
    .A(_07088_));
 sg13g2_a21oi_1 _18079_ (.A1(_08983_),
    .A2(_07083_),
    .Y(_08984_),
    .B1(_07091_));
 sg13g2_buf_2 _18080_ (.A(_08984_),
    .X(_08985_));
 sg13g2_a21oi_1 _18081_ (.A1(_08281_),
    .A2(_08985_),
    .Y(_08986_),
    .B1(_07137_));
 sg13g2_nor3_1 _18082_ (.A(_08978_),
    .B(_08982_),
    .C(_08986_),
    .Y(_08987_));
 sg13g2_nand4_1 _18083_ (.B(_08968_),
    .C(_08975_),
    .A(_08964_),
    .Y(_08988_),
    .D(_08987_));
 sg13g2_nor3_1 _18084_ (.A(_08931_),
    .B(_08951_),
    .C(_08988_),
    .Y(_08989_));
 sg13g2_nor2_1 _18085_ (.A(_04001_),
    .B(_04270_),
    .Y(_08990_));
 sg13g2_nor2_1 _18086_ (.A(_03221_),
    .B(_07513_),
    .Y(_08991_));
 sg13g2_inv_1 _18087_ (.Y(_08992_),
    .A(_08924_));
 sg13g2_nor2_1 _18088_ (.A(_08929_),
    .B(_08992_),
    .Y(_08993_));
 sg13g2_inv_1 _18089_ (.Y(_08994_),
    .A(_08908_));
 sg13g2_nor2_1 _18090_ (.A(_08994_),
    .B(_08917_),
    .Y(_08995_));
 sg13g2_nor4_1 _18091_ (.A(_08990_),
    .B(_08991_),
    .C(_08993_),
    .D(_08995_),
    .Y(_08996_));
 sg13g2_a21oi_1 _18092_ (.A1(_03221_),
    .A2(_06165_),
    .Y(_08997_),
    .B1(_08948_));
 sg13g2_nor2_1 _18093_ (.A(_08944_),
    .B(_07492_),
    .Y(_08998_));
 sg13g2_nor2_1 _18094_ (.A(_08997_),
    .B(_08998_),
    .Y(_08999_));
 sg13g2_inv_1 _18095_ (.Y(_09000_),
    .A(_08999_));
 sg13g2_nor2_2 _18096_ (.A(_08938_),
    .B(_06168_),
    .Y(_09001_));
 sg13g2_nor2_1 _18097_ (.A(_08933_),
    .B(_05951_),
    .Y(_09002_));
 sg13g2_buf_2 _18098_ (.A(_09002_),
    .X(_09003_));
 sg13g2_nor3_1 _18099_ (.A(_09000_),
    .B(_09001_),
    .C(_09003_),
    .Y(_09004_));
 sg13g2_inv_1 _18100_ (.Y(_09005_),
    .A(_08963_));
 sg13g2_inv_1 _18101_ (.Y(_09006_),
    .A(_08413_));
 sg13g2_nand2b_1 _18102_ (.Y(_09007_),
    .B(_09006_),
    .A_N(_07743_));
 sg13g2_nand2_1 _18103_ (.Y(_09008_),
    .A(_08971_),
    .B(_00055_));
 sg13g2_inv_1 _18104_ (.Y(_09009_),
    .A(_07752_));
 sg13g2_nand2_1 _18105_ (.Y(_09010_),
    .A(_09008_),
    .B(_09009_));
 sg13g2_nor2_1 _18106_ (.A(_09007_),
    .B(_09010_),
    .Y(_09011_));
 sg13g2_inv_1 _18107_ (.Y(_09012_),
    .A(_06683_));
 sg13g2_a22oi_1 _18108_ (.Y(_09013_),
    .B1(_06727_),
    .B2(_09012_),
    .A2(_08965_),
    .A1(_05311_));
 sg13g2_inv_1 _18109_ (.Y(_09014_),
    .A(_07137_));
 sg13g2_nor2_1 _18110_ (.A(_08985_),
    .B(_09014_),
    .Y(_09015_));
 sg13g2_nor2_1 _18111_ (.A(_08281_),
    .B(_09014_),
    .Y(_09016_));
 sg13g2_nor2_1 _18112_ (.A(_09015_),
    .B(_09016_),
    .Y(_09017_));
 sg13g2_nor2_1 _18113_ (.A(_08966_),
    .B(_08977_),
    .Y(_09018_));
 sg13g2_inv_1 _18114_ (.Y(_09019_),
    .A(_04176_));
 sg13g2_nor2_1 _18115_ (.A(_08981_),
    .B(_09019_),
    .Y(_09020_));
 sg13g2_nor2_1 _18116_ (.A(_09018_),
    .B(_09020_),
    .Y(_09021_));
 sg13g2_nand4_1 _18117_ (.B(_09013_),
    .C(_09017_),
    .A(_09011_),
    .Y(_09022_),
    .D(_09021_));
 sg13g2_a21oi_1 _18118_ (.A1(_08959_),
    .A2(_09005_),
    .Y(_09023_),
    .B1(_09022_));
 sg13g2_and3_1 _18119_ (.X(_09024_),
    .A(_08996_),
    .B(_09004_),
    .C(_09023_));
 sg13g2_nor3_1 _18120_ (.A(_04189_),
    .B(_08989_),
    .C(_09024_),
    .Y(_09025_));
 sg13g2_nand2_1 _18121_ (.Y(_09026_),
    .A(_09025_),
    .B(net162));
 sg13g2_nand2_1 _18122_ (.Y(_09027_),
    .A(_09024_),
    .B(_08989_));
 sg13g2_o21ai_1 _18123_ (.B1(_04183_),
    .Y(_09028_),
    .A1(_04180_),
    .A2(_04189_));
 sg13g2_nand3_1 _18124_ (.B(net113),
    .C(_09028_),
    .A(_09027_),
    .Y(_09029_));
 sg13g2_o21ai_1 _18125_ (.B1(_09029_),
    .Y(_09030_),
    .A1(_04180_),
    .A2(_09026_));
 sg13g2_nand3_1 _18126_ (.B(_09013_),
    .C(_08281_),
    .A(_08968_),
    .Y(_09031_));
 sg13g2_o21ai_1 _18127_ (.B1(_04189_),
    .Y(_09032_),
    .A1(_09031_),
    .A2(_08956_));
 sg13g2_nor2b_1 _18128_ (.A(_09032_),
    .B_N(_05313_),
    .Y(_09033_));
 sg13g2_inv_1 _18129_ (.Y(_09034_),
    .A(_08996_));
 sg13g2_o21ai_1 _18130_ (.B1(_04189_),
    .Y(_09035_),
    .A1(_08931_),
    .A2(_09034_));
 sg13g2_a21o_1 _18131_ (.A2(_09032_),
    .A1(_09035_),
    .B1(_04276_),
    .X(_09036_));
 sg13g2_nand3b_1 _18132_ (.B(_09036_),
    .C(_04187_),
    .Y(_09037_),
    .A_N(_09033_));
 sg13g2_inv_1 _18133_ (.Y(_09038_),
    .A(_08951_));
 sg13g2_nor2_1 _18134_ (.A(_08980_),
    .B(_08976_),
    .Y(_09039_));
 sg13g2_inv_1 _18135_ (.Y(_09040_),
    .A(_08985_));
 sg13g2_inv_1 _18136_ (.Y(_09041_),
    .A(_08958_));
 sg13g2_nor3_1 _18137_ (.A(_04187_),
    .B(_09040_),
    .C(_09041_),
    .Y(_09042_));
 sg13g2_nand4_1 _18138_ (.B(_09004_),
    .C(_09039_),
    .A(_09038_),
    .Y(_09043_),
    .D(_09042_));
 sg13g2_nor2_1 _18139_ (.A(net103),
    .B(_04190_),
    .Y(_09044_));
 sg13g2_and3_1 _18140_ (.X(_09045_),
    .A(_09037_),
    .B(_09043_),
    .C(_09044_));
 sg13g2_buf_1 _18141_ (.A(\b.gen_square[14].sq.mask ),
    .X(_09046_));
 sg13g2_o21ai_1 _18142_ (.B1(_09046_),
    .Y(_09047_),
    .A1(_09030_),
    .A2(_09045_));
 sg13g2_a21oi_1 _18143_ (.A1(_07823_),
    .A2(_06696_),
    .Y(_09048_),
    .B1(_06731_));
 sg13g2_inv_1 _18144_ (.Y(_09049_),
    .A(_09048_));
 sg13g2_a21oi_1 _18145_ (.A1(_09049_),
    .A2(_06185_),
    .Y(_09050_),
    .B1(_06189_));
 sg13g2_inv_1 _18146_ (.Y(_09051_),
    .A(_09050_));
 sg13g2_a21oi_1 _18147_ (.A1(_09051_),
    .A2(net25),
    .Y(_09052_),
    .B1(_05527_));
 sg13g2_a21oi_1 _18148_ (.A1(_07792_),
    .A2(net50),
    .Y(_09053_),
    .B1(_07122_));
 sg13g2_inv_1 _18149_ (.Y(_09054_),
    .A(_09053_));
 sg13g2_a21oi_1 _18150_ (.A1(_09054_),
    .A2(_06185_),
    .Y(_09055_),
    .B1(_07114_));
 sg13g2_inv_1 _18151_ (.Y(_09056_),
    .A(_09055_));
 sg13g2_a21oi_1 _18152_ (.A1(_09056_),
    .A2(net25),
    .Y(_09057_),
    .B1(_07106_));
 sg13g2_nand3_1 _18153_ (.B(_06165_),
    .C(_03221_),
    .A(net90),
    .Y(_09058_));
 sg13g2_nand2_1 _18154_ (.Y(_09059_),
    .A(_04195_),
    .B(\b.gen_square[14].sq.color ));
 sg13g2_nand2_1 _18155_ (.Y(_09060_),
    .A(_09058_),
    .B(_09059_));
 sg13g2_nand2_1 _18156_ (.Y(_09061_),
    .A(_07513_),
    .B(_04194_));
 sg13g2_nand2_1 _18157_ (.Y(_09062_),
    .A(_04279_),
    .B(_09061_));
 sg13g2_inv_1 _18158_ (.Y(_09063_),
    .A(_09062_));
 sg13g2_inv_1 _18159_ (.Y(_09064_),
    .A(_07092_));
 sg13g2_a22oi_1 _18160_ (.Y(_09065_),
    .B1(_09014_),
    .B2(_09064_),
    .A2(_09063_),
    .A1(_09060_));
 sg13g2_o21ai_1 _18161_ (.B1(_09065_),
    .Y(_09066_),
    .A1(_08907_),
    .A2(_08916_));
 sg13g2_a21o_1 _18162_ (.A2(_09057_),
    .A1(_09052_),
    .B1(_09066_),
    .X(_09067_));
 sg13g2_inv_1 _18163_ (.Y(_09068_),
    .A(_09067_));
 sg13g2_inv_1 _18164_ (.Y(_09069_),
    .A(_09052_));
 sg13g2_nand2_1 _18165_ (.Y(_09070_),
    .A(_06167_),
    .B(net90));
 sg13g2_nand2_1 _18166_ (.Y(_09071_),
    .A(_09070_),
    .B(_04196_));
 sg13g2_a22oi_1 _18167_ (.Y(_09072_),
    .B1(_09063_),
    .B2(_09071_),
    .A2(_09064_),
    .A1(_00048_));
 sg13g2_o21ai_1 _18168_ (.B1(_09072_),
    .Y(_09073_),
    .A1(_08907_),
    .A2(_08915_));
 sg13g2_a21oi_1 _18169_ (.A1(_09069_),
    .A2(_09057_),
    .Y(_09074_),
    .B1(_09073_));
 sg13g2_a21oi_1 _18170_ (.A1(_09068_),
    .A2(_09074_),
    .Y(_09075_),
    .B1(_05891_));
 sg13g2_inv_1 _18171_ (.Y(_09076_),
    .A(_09075_));
 sg13g2_o21ai_1 _18172_ (.B1(_05922_),
    .Y(_09077_),
    .A1(_05845_),
    .A2(_08029_));
 sg13g2_a21oi_1 _18173_ (.A1(_09077_),
    .A2(net42),
    .Y(_09078_),
    .B1(_04907_));
 sg13g2_inv_1 _18174_ (.Y(_09079_),
    .A(_09078_));
 sg13g2_inv_1 _18175_ (.Y(_09080_),
    .A(_05910_));
 sg13g2_a21oi_1 _18176_ (.A1(_09079_),
    .A2(net22),
    .Y(_09081_),
    .B1(_09080_));
 sg13g2_inv_1 _18177_ (.Y(_09082_),
    .A(_09081_));
 sg13g2_nor2_1 _18178_ (.A(_08160_),
    .B(_06999_),
    .Y(_09083_));
 sg13g2_a21oi_1 _18179_ (.A1(_06863_),
    .A2(net62),
    .Y(_09084_),
    .B1(_06217_));
 sg13g2_a21oi_1 _18180_ (.A1(_04098_),
    .A2(net62),
    .Y(_09085_),
    .B1(_04220_));
 sg13g2_nor2_1 _18181_ (.A(_04176_),
    .B(_05872_),
    .Y(_09086_));
 sg13g2_a21oi_1 _18182_ (.A1(_09084_),
    .A2(_09085_),
    .Y(_09087_),
    .B1(_09086_));
 sg13g2_inv_1 _18183_ (.Y(_09088_),
    .A(_09087_));
 sg13g2_inv_1 _18184_ (.Y(_09089_),
    .A(_09084_));
 sg13g2_nor2_1 _18185_ (.A(_05872_),
    .B(_09019_),
    .Y(_09090_));
 sg13g2_nor2_1 _18186_ (.A(_08160_),
    .B(_06998_),
    .Y(_09091_));
 sg13g2_nor2_1 _18187_ (.A(_09090_),
    .B(_09091_),
    .Y(_09092_));
 sg13g2_o21ai_1 _18188_ (.B1(_09092_),
    .Y(_09093_),
    .A1(_09085_),
    .A2(_09089_));
 sg13g2_nor3_1 _18189_ (.A(_09083_),
    .B(_09088_),
    .C(_09093_),
    .Y(_09094_));
 sg13g2_a21o_1 _18190_ (.A2(_09094_),
    .A1(_09082_),
    .B1(_05891_),
    .X(_09095_));
 sg13g2_a21o_1 _18191_ (.A2(_09095_),
    .A1(_09076_),
    .B1(_05895_),
    .X(_09096_));
 sg13g2_nand2b_1 _18192_ (.Y(_09097_),
    .B(_05893_),
    .A_N(_09095_));
 sg13g2_nand3_1 _18193_ (.B(_05882_),
    .C(_09097_),
    .A(_09096_),
    .Y(_09098_));
 sg13g2_a21oi_2 _18194_ (.B1(_06952_),
    .Y(_09099_),
    .A2(_06957_),
    .A1(_06947_));
 sg13g2_nor2_1 _18195_ (.A(_09099_),
    .B(_08804_),
    .Y(_09100_));
 sg13g2_buf_1 _18196_ (.A(_09100_),
    .X(_09101_));
 sg13g2_nor2_1 _18197_ (.A(_08958_),
    .B(_05528_),
    .Y(_09102_));
 sg13g2_buf_2 _18198_ (.A(_09102_),
    .X(_09103_));
 sg13g2_a21oi_2 _18199_ (.B1(_05861_),
    .Y(_09104_),
    .A2(_05906_),
    .A1(_05856_));
 sg13g2_nor2_1 _18200_ (.A(_09104_),
    .B(_05957_),
    .Y(_09105_));
 sg13g2_buf_2 _18201_ (.A(_09105_),
    .X(_09106_));
 sg13g2_inv_1 _18202_ (.Y(_09107_),
    .A(_04187_));
 sg13g2_a21oi_1 _18203_ (.A1(_09107_),
    .A2(_04273_),
    .Y(_09108_),
    .B1(_04192_));
 sg13g2_buf_2 _18204_ (.A(_09108_),
    .X(_09109_));
 sg13g2_nor2_1 _18205_ (.A(_09020_),
    .B(_09001_),
    .Y(_09110_));
 sg13g2_o21ai_1 _18206_ (.B1(_09110_),
    .Y(_09111_),
    .A1(_09109_),
    .A2(_09060_));
 sg13g2_nor4_1 _18207_ (.A(_09101_),
    .B(_09103_),
    .C(_09106_),
    .D(_09111_),
    .Y(_09112_));
 sg13g2_nor2_2 _18208_ (.A(_09099_),
    .B(_08805_),
    .Y(_09113_));
 sg13g2_nor2_2 _18209_ (.A(_09109_),
    .B(_09071_),
    .Y(_09114_));
 sg13g2_nor2_2 _18210_ (.A(_08958_),
    .B(_05529_),
    .Y(_09115_));
 sg13g2_nor4_1 _18211_ (.A(_08940_),
    .B(_09113_),
    .C(_09114_),
    .D(_09115_),
    .Y(_09116_));
 sg13g2_nor2_1 _18212_ (.A(_09104_),
    .B(_05958_),
    .Y(_09117_));
 sg13g2_buf_2 _18213_ (.A(_09117_),
    .X(_09118_));
 sg13g2_nor2_1 _18214_ (.A(_08982_),
    .B(_09118_),
    .Y(_09119_));
 sg13g2_a21oi_1 _18215_ (.A1(_06922_),
    .A2(_06933_),
    .Y(_09120_),
    .B1(_06994_));
 sg13g2_inv_1 _18216_ (.Y(_09121_),
    .A(_09120_));
 sg13g2_nor3_1 _18217_ (.A(_05882_),
    .B(_09040_),
    .C(_09121_),
    .Y(_09122_));
 sg13g2_nand4_1 _18218_ (.B(_09116_),
    .C(_09119_),
    .A(_09112_),
    .Y(_09123_),
    .D(_09122_));
 sg13g2_nor2_1 _18219_ (.A(net120),
    .B(_05885_),
    .Y(_09124_));
 sg13g2_nand3_1 _18220_ (.B(_09123_),
    .C(_09124_),
    .A(_09098_),
    .Y(_09125_));
 sg13g2_nand4_1 _18221_ (.B(_06532_),
    .C(_06544_),
    .A(_06540_),
    .Y(_09126_),
    .D(_06533_));
 sg13g2_o21ai_1 _18222_ (.B1(_06549_),
    .Y(_09127_),
    .A1(net79),
    .A2(_09126_));
 sg13g2_nand2_1 _18223_ (.Y(_09128_),
    .A(_09127_),
    .B(_00012_));
 sg13g2_inv_1 _18224_ (.Y(_09129_),
    .A(_09128_));
 sg13g2_or4_1 _18225_ (.A(_07934_),
    .B(_08676_),
    .C(_09129_),
    .D(_08106_),
    .X(_09130_));
 sg13g2_nor2_1 _18226_ (.A(_09120_),
    .B(_06998_),
    .Y(_09131_));
 sg13g2_inv_1 _18227_ (.Y(_09132_),
    .A(_09131_));
 sg13g2_inv_1 _18228_ (.Y(_09133_),
    .A(_05292_));
 sg13g2_nor3_1 _18229_ (.A(_05291_),
    .B(_05293_),
    .C(_09133_),
    .Y(_09134_));
 sg13g2_nand2_1 _18230_ (.Y(_09135_),
    .A(_05302_),
    .B(_09134_));
 sg13g2_inv_1 _18231_ (.Y(_09136_),
    .A(_09135_));
 sg13g2_a21oi_1 _18232_ (.A1(_04530_),
    .A2(_09136_),
    .Y(_09137_),
    .B1(_05309_));
 sg13g2_nor2_1 _18233_ (.A(_05521_),
    .B(_09137_),
    .Y(_09138_));
 sg13g2_nor2_1 _18234_ (.A(_09138_),
    .B(_08109_),
    .Y(_09139_));
 sg13g2_nand3b_1 _18235_ (.B(_09132_),
    .C(_09139_),
    .Y(_09140_),
    .A_N(_09015_));
 sg13g2_inv_1 _18236_ (.Y(_09141_),
    .A(_08343_));
 sg13g2_a21oi_1 _18237_ (.A1(_09141_),
    .A2(net42),
    .Y(_09142_),
    .B1(_04967_));
 sg13g2_inv_1 _18238_ (.Y(_09143_),
    .A(_09142_));
 sg13g2_a21oi_1 _18239_ (.A1(_09143_),
    .A2(net22),
    .Y(_09144_),
    .B1(_05956_));
 sg13g2_nor2_1 _18240_ (.A(_09082_),
    .B(_09144_),
    .Y(_09145_));
 sg13g2_nor4_1 _18241_ (.A(_09130_),
    .B(_09093_),
    .C(_09140_),
    .D(_09145_),
    .Y(_09146_));
 sg13g2_nand3_1 _18242_ (.B(_09112_),
    .C(_09146_),
    .A(_09074_),
    .Y(_09147_));
 sg13g2_nor2_1 _18243_ (.A(_04010_),
    .B(_09137_),
    .Y(_09148_));
 sg13g2_nor2b_1 _18244_ (.A(_06798_),
    .B_N(_09127_),
    .Y(_09149_));
 sg13g2_nor2_1 _18245_ (.A(_08669_),
    .B(_09149_),
    .Y(_09150_));
 sg13g2_nor2_1 _18246_ (.A(_07896_),
    .B(_08040_),
    .Y(_09151_));
 sg13g2_nand2_1 _18247_ (.Y(_09152_),
    .A(_09150_),
    .B(_09151_));
 sg13g2_nor4_1 _18248_ (.A(_07919_),
    .B(_09148_),
    .C(_09083_),
    .D(_09152_),
    .Y(_09153_));
 sg13g2_nor2_1 _18249_ (.A(_08985_),
    .B(_07137_),
    .Y(_09154_));
 sg13g2_inv_1 _18250_ (.Y(_09155_),
    .A(_09154_));
 sg13g2_nor2_1 _18251_ (.A(_09120_),
    .B(_06999_),
    .Y(_09156_));
 sg13g2_inv_1 _18252_ (.Y(_09157_),
    .A(_09156_));
 sg13g2_nand4_1 _18253_ (.B(_09155_),
    .C(_09157_),
    .A(_09153_),
    .Y(_09158_),
    .D(_09087_));
 sg13g2_a21oi_1 _18254_ (.A1(_09144_),
    .A2(_09081_),
    .Y(_09159_),
    .B1(_09158_));
 sg13g2_nand4_1 _18255_ (.B(_09116_),
    .C(_09119_),
    .A(_09068_),
    .Y(_09160_),
    .D(_09159_));
 sg13g2_nor2_1 _18256_ (.A(_09147_),
    .B(_09160_),
    .Y(_09161_));
 sg13g2_inv_1 _18257_ (.Y(_09162_),
    .A(_09161_));
 sg13g2_o21ai_1 _18258_ (.B1(_05879_),
    .Y(_09163_),
    .A1(_05876_),
    .A2(_05884_));
 sg13g2_nand3_1 _18259_ (.B(net129),
    .C(_09163_),
    .A(_09162_),
    .Y(_09164_));
 sg13g2_nand4_1 _18260_ (.B(net177),
    .C(_05891_),
    .A(_09160_),
    .Y(_09165_),
    .D(_09147_));
 sg13g2_buf_1 _18261_ (.A(_09165_),
    .X(_09166_));
 sg13g2_or2_1 _18262_ (.X(_09167_),
    .B(_09166_),
    .A(_05876_));
 sg13g2_nand3_1 _18263_ (.B(_09164_),
    .C(_09167_),
    .A(_09125_),
    .Y(_09168_));
 sg13g2_buf_1 _18264_ (.A(\b.gen_square[13].sq.mask ),
    .X(_09169_));
 sg13g2_nand2_1 _18265_ (.Y(_09170_),
    .A(_09168_),
    .B(_09169_));
 sg13g2_nand2_1 _18266_ (.Y(_09171_),
    .A(_08222_),
    .B(_06093_));
 sg13g2_nand3_1 _18267_ (.B(_05500_),
    .C(_06077_),
    .A(_09171_),
    .Y(_09172_));
 sg13g2_o21ai_1 _18268_ (.B1(_00058_),
    .Y(_09173_),
    .A1(_06076_),
    .A2(_05161_));
 sg13g2_nand2_1 _18269_ (.Y(_09174_),
    .A(_09172_),
    .B(_09173_));
 sg13g2_nand2_1 _18270_ (.Y(_09175_),
    .A(_09174_),
    .B(_06058_));
 sg13g2_inv_1 _18271_ (.Y(_09176_),
    .A(_06111_));
 sg13g2_nand2_1 _18272_ (.Y(_09177_),
    .A(_09175_),
    .B(_09176_));
 sg13g2_nand2_1 _18273_ (.Y(_09178_),
    .A(_09177_),
    .B(_06030_));
 sg13g2_inv_1 _18274_ (.Y(_09179_),
    .A(_06107_));
 sg13g2_nand2_1 _18275_ (.Y(_09180_),
    .A(_09178_),
    .B(_09179_));
 sg13g2_nand2_1 _18276_ (.Y(_09181_),
    .A(_08186_),
    .B(_06077_));
 sg13g2_nand2b_1 _18277_ (.Y(_09182_),
    .B(_09181_),
    .A_N(_06090_));
 sg13g2_buf_1 _18278_ (.A(_09182_),
    .X(_09183_));
 sg13g2_nand2_1 _18279_ (.Y(_09184_),
    .A(_09183_),
    .B(_06058_));
 sg13g2_inv_1 _18280_ (.Y(_09185_),
    .A(_06071_));
 sg13g2_nand2_2 _18281_ (.Y(_09186_),
    .A(_09184_),
    .B(_09185_));
 sg13g2_a21oi_1 _18282_ (.A1(_09186_),
    .A2(_06030_),
    .Y(_09187_),
    .B1(_06039_));
 sg13g2_nand2_1 _18283_ (.Y(_09188_),
    .A(_09180_),
    .B(_09187_));
 sg13g2_nand3_1 _18284_ (.B(_05377_),
    .C(_08396_),
    .A(_08395_),
    .Y(_09189_));
 sg13g2_nand2_1 _18285_ (.Y(_09190_),
    .A(_06512_),
    .B(\b.gen_square[35].sq.color ));
 sg13g2_nand3_1 _18286_ (.B(_06391_),
    .C(_09190_),
    .A(_09189_),
    .Y(_09191_));
 sg13g2_nand2_1 _18287_ (.Y(_09192_),
    .A(_08277_),
    .B(_03632_));
 sg13g2_nand3_1 _18288_ (.B(net38),
    .C(_09192_),
    .A(_09191_),
    .Y(_09193_));
 sg13g2_inv_1 _18289_ (.Y(_09194_),
    .A(_05582_));
 sg13g2_a21oi_1 _18290_ (.A1(_09194_),
    .A2(_05623_),
    .Y(_09195_),
    .B1(_08044_));
 sg13g2_inv_1 _18291_ (.Y(_09196_),
    .A(_09195_));
 sg13g2_nor2_1 _18292_ (.A(_03512_),
    .B(_05709_),
    .Y(_09197_));
 sg13g2_inv_1 _18293_ (.Y(_09198_),
    .A(_09197_));
 sg13g2_nand3_1 _18294_ (.B(_09196_),
    .C(_09198_),
    .A(_09193_),
    .Y(_09199_));
 sg13g2_buf_1 _18295_ (.A(_09199_),
    .X(_09200_));
 sg13g2_nand2_1 _18296_ (.Y(_09201_),
    .A(_09188_),
    .B(_09200_));
 sg13g2_nand2_1 _18297_ (.Y(_09202_),
    .A(_07981_),
    .B(_06391_));
 sg13g2_inv_1 _18298_ (.Y(_09203_),
    .A(_06433_));
 sg13g2_nand2_1 _18299_ (.Y(_09204_),
    .A(_09202_),
    .B(_09203_));
 sg13g2_nand2_1 _18300_ (.Y(_09205_),
    .A(_09204_),
    .B(net38));
 sg13g2_nand2_1 _18301_ (.Y(_09206_),
    .A(_09205_),
    .B(_05712_));
 sg13g2_nand2_1 _18302_ (.Y(_09207_),
    .A(_08392_),
    .B(_05377_));
 sg13g2_nand2_1 _18303_ (.Y(_09208_),
    .A(_09207_),
    .B(_05386_));
 sg13g2_nand2_1 _18304_ (.Y(_09209_),
    .A(_09208_),
    .B(_06391_));
 sg13g2_nand2_1 _18305_ (.Y(_09210_),
    .A(_09209_),
    .B(_07202_));
 sg13g2_a21oi_1 _18306_ (.A1(_09210_),
    .A2(net38),
    .Y(_09211_),
    .B1(_07196_));
 sg13g2_nand2_1 _18307_ (.Y(_09212_),
    .A(_09206_),
    .B(_09211_));
 sg13g2_nor4_1 _18308_ (.A(_06337_),
    .B(_06336_),
    .C(_06340_),
    .D(_06351_),
    .Y(_09213_));
 sg13g2_a21o_1 _18309_ (.A2(_09213_),
    .A1(net133),
    .B1(_06419_),
    .X(_09214_));
 sg13g2_nand2_1 _18310_ (.Y(_09215_),
    .A(_09214_),
    .B(_00013_));
 sg13g2_inv_1 _18311_ (.Y(_09216_),
    .A(_09215_));
 sg13g2_nor3_1 _18312_ (.A(_08418_),
    .B(_08265_),
    .C(_09216_),
    .Y(_09217_));
 sg13g2_inv_2 _18313_ (.Y(_09218_),
    .A(_04853_));
 sg13g2_nand3_1 _18314_ (.B(net131),
    .C(_09218_),
    .A(net133),
    .Y(_09219_));
 sg13g2_nand2_1 _18315_ (.Y(_09220_),
    .A(_04856_),
    .B(_09219_));
 sg13g2_inv_1 _18316_ (.Y(_09221_),
    .A(_09220_));
 sg13g2_inv_4 _18317_ (.A(_04953_),
    .Y(_09222_));
 sg13g2_nor2_1 _18318_ (.A(_09221_),
    .B(_09222_),
    .Y(_09223_));
 sg13g2_a21oi_1 _18319_ (.A1(_05608_),
    .A2(_05604_),
    .Y(_09224_),
    .B1(_05611_));
 sg13g2_nor2_1 _18320_ (.A(_09224_),
    .B(_05705_),
    .Y(_09225_));
 sg13g2_nor2_1 _18321_ (.A(_09223_),
    .B(_09225_),
    .Y(_09226_));
 sg13g2_nor2_1 _18322_ (.A(_06000_),
    .B(_09222_),
    .Y(_09227_));
 sg13g2_nor2_1 _18323_ (.A(_07578_),
    .B(_05705_),
    .Y(_09228_));
 sg13g2_nor2_1 _18324_ (.A(_09227_),
    .B(_09228_),
    .Y(_09229_));
 sg13g2_and3_1 _18325_ (.X(_09230_),
    .A(_09217_),
    .B(_09226_),
    .C(_09229_));
 sg13g2_nand2_1 _18326_ (.Y(_09231_),
    .A(_09212_),
    .B(_09230_));
 sg13g2_nor2_1 _18327_ (.A(_09201_),
    .B(_09231_),
    .Y(_09232_));
 sg13g2_nand2_1 _18328_ (.Y(_09233_),
    .A(_09071_),
    .B(net73));
 sg13g2_nand2b_1 _18329_ (.Y(_09234_),
    .B(_09233_),
    .A_N(_05950_));
 sg13g2_nand2_1 _18330_ (.Y(_09235_),
    .A(_09234_),
    .B(net65));
 sg13g2_nand2b_1 _18331_ (.Y(_09236_),
    .B(_09235_),
    .A_N(_07002_));
 sg13g2_nand2_1 _18332_ (.Y(_09237_),
    .A(_09236_),
    .B(_06529_));
 sg13g2_nand2_1 _18333_ (.Y(_09238_),
    .A(_09237_),
    .B(_08913_));
 sg13g2_nand2_1 _18334_ (.Y(_09239_),
    .A(_09238_),
    .B(_06333_));
 sg13g2_inv_1 _18335_ (.Y(_09240_),
    .A(_06426_));
 sg13g2_nand2_1 _18336_ (.Y(_09241_),
    .A(_09239_),
    .B(_09240_));
 sg13g2_nand2_1 _18337_ (.Y(_09242_),
    .A(_09241_),
    .B(net59));
 sg13g2_inv_1 _18338_ (.Y(_09243_),
    .A(_04956_));
 sg13g2_nand2_1 _18339_ (.Y(_09244_),
    .A(_09242_),
    .B(_09243_));
 sg13g2_nand2_1 _18340_ (.Y(_09245_),
    .A(_09062_),
    .B(net73));
 sg13g2_nand2_1 _18341_ (.Y(_09246_),
    .A(_09245_),
    .B(_07096_));
 sg13g2_nand2_1 _18342_ (.Y(_09247_),
    .A(_09246_),
    .B(_06954_));
 sg13g2_nand2_1 _18343_ (.Y(_09248_),
    .A(_09247_),
    .B(_06963_));
 sg13g2_nand2_1 _18344_ (.Y(_09249_),
    .A(_09248_),
    .B(_06529_));
 sg13g2_nand2_1 _18345_ (.Y(_09250_),
    .A(_09249_),
    .B(_06559_));
 sg13g2_a21oi_1 _18346_ (.A1(_09250_),
    .A2(_06333_),
    .Y(_09251_),
    .B1(_06363_));
 sg13g2_nor2b_1 _18347_ (.A(_09251_),
    .B_N(net59),
    .Y(_09252_));
 sg13g2_nor2_1 _18348_ (.A(_05616_),
    .B(_09252_),
    .Y(_09253_));
 sg13g2_nand2_1 _18349_ (.Y(_09254_),
    .A(_09244_),
    .B(_09253_));
 sg13g2_nand2_1 _18350_ (.Y(_09255_),
    .A(_09232_),
    .B(_09254_));
 sg13g2_a21oi_2 _18351_ (.B1(_04832_),
    .Y(_09256_),
    .A2(_04864_),
    .A1(_04827_));
 sg13g2_nor2_1 _18352_ (.A(_04026_),
    .B(net59),
    .Y(_09257_));
 sg13g2_a21oi_1 _18353_ (.A1(_06888_),
    .A2(net59),
    .Y(_09258_),
    .B1(_09257_));
 sg13g2_inv_1 _18354_ (.Y(_09259_),
    .A(_09258_));
 sg13g2_nor2_1 _18355_ (.A(_09256_),
    .B(_09259_),
    .Y(_09260_));
 sg13g2_inv_1 _18356_ (.Y(_09261_),
    .A(_06024_));
 sg13g2_nor3_1 _18357_ (.A(_06022_),
    .B(_09261_),
    .C(_04313_),
    .Y(_09262_));
 sg13g2_nor2_1 _18358_ (.A(_09262_),
    .B(_06028_),
    .Y(_09263_));
 sg13g2_buf_2 _18359_ (.A(_09263_),
    .X(_09264_));
 sg13g2_nor2_1 _18360_ (.A(_09264_),
    .B(_06108_),
    .Y(_09265_));
 sg13g2_nor2_1 _18361_ (.A(_09260_),
    .B(_09265_),
    .Y(_09266_));
 sg13g2_nor2b_1 _18362_ (.A(_09255_),
    .B_N(_09266_),
    .Y(_09267_));
 sg13g2_nand2_1 _18363_ (.Y(_09268_),
    .A(_09193_),
    .B(_09198_));
 sg13g2_nand2_1 _18364_ (.Y(_09269_),
    .A(_09211_),
    .B(_09268_));
 sg13g2_a21oi_1 _18365_ (.A1(_09177_),
    .A2(_06030_),
    .Y(_09270_),
    .B1(_06107_));
 sg13g2_nand2_1 _18366_ (.Y(_09271_),
    .A(_09270_),
    .B(_09187_));
 sg13g2_nand2_1 _18367_ (.Y(_09272_),
    .A(_09269_),
    .B(_09271_));
 sg13g2_o21ai_1 _18368_ (.B1(_05712_),
    .Y(_09273_),
    .A1(_05590_),
    .A2(_06742_));
 sg13g2_nor2_1 _18369_ (.A(_09195_),
    .B(_09273_),
    .Y(_09274_));
 sg13g2_buf_2 _18370_ (.A(_09274_),
    .X(_09275_));
 sg13g2_nor2_1 _18371_ (.A(_09221_),
    .B(_04953_),
    .Y(_09276_));
 sg13g2_nor2_1 _18372_ (.A(_04953_),
    .B(_06000_),
    .Y(_09277_));
 sg13g2_nor2_1 _18373_ (.A(_07578_),
    .B(_05706_),
    .Y(_09278_));
 sg13g2_nor2_1 _18374_ (.A(_09224_),
    .B(_05706_),
    .Y(_09279_));
 sg13g2_nor4_1 _18375_ (.A(_09276_),
    .B(_09277_),
    .C(_09278_),
    .D(_09279_),
    .Y(_09280_));
 sg13g2_nand2_1 _18376_ (.Y(_09281_),
    .A(_09214_),
    .B(_03668_));
 sg13g2_inv_1 _18377_ (.Y(_09282_),
    .A(_08269_));
 sg13g2_nand2_1 _18378_ (.Y(_09283_),
    .A(_09281_),
    .B(_09282_));
 sg13g2_nor2_1 _18379_ (.A(_08423_),
    .B(_09283_),
    .Y(_09284_));
 sg13g2_nand2_1 _18380_ (.Y(_09285_),
    .A(_09280_),
    .B(_09284_));
 sg13g2_nor2_1 _18381_ (.A(_09275_),
    .B(_09285_),
    .Y(_09286_));
 sg13g2_nor2b_1 _18382_ (.A(_09272_),
    .B_N(_09286_),
    .Y(_09287_));
 sg13g2_inv_1 _18383_ (.Y(_09288_),
    .A(\b.gen_square[12].sq.color ));
 sg13g2_nor2_1 _18384_ (.A(_09288_),
    .B(net65),
    .Y(_09289_));
 sg13g2_nand3_1 _18385_ (.B(_09059_),
    .C(net73),
    .A(_09058_),
    .Y(_09290_));
 sg13g2_inv_1 _18386_ (.Y(_09291_),
    .A(net73));
 sg13g2_nand2_1 _18387_ (.Y(_09292_),
    .A(_09291_),
    .B(_02939_));
 sg13g2_nand3_1 _18388_ (.B(_06954_),
    .C(_09292_),
    .A(_09290_),
    .Y(_09293_));
 sg13g2_nand2b_1 _18389_ (.Y(_09294_),
    .B(_09293_),
    .A_N(_09289_));
 sg13g2_nand2_1 _18390_ (.Y(_09295_),
    .A(_09294_),
    .B(_06529_));
 sg13g2_nand2_1 _18391_ (.Y(_09296_),
    .A(_08909_),
    .B(\b.gen_square[11].sq.color ));
 sg13g2_nand2_1 _18392_ (.Y(_09297_),
    .A(_09295_),
    .B(_09296_));
 sg13g2_nand2_1 _18393_ (.Y(_09298_),
    .A(_09297_),
    .B(_06333_));
 sg13g2_nor2_1 _18394_ (.A(_02393_),
    .B(_06333_),
    .Y(_09299_));
 sg13g2_inv_1 _18395_ (.Y(_09300_),
    .A(_09299_));
 sg13g2_nand2_1 _18396_ (.Y(_09301_),
    .A(_09298_),
    .B(_09300_));
 sg13g2_nand2_1 _18397_ (.Y(_09302_),
    .A(_09301_),
    .B(_04834_));
 sg13g2_nand2b_1 _18398_ (.Y(_09303_),
    .B(_09302_),
    .A_N(_09257_));
 sg13g2_nand2_1 _18399_ (.Y(_09304_),
    .A(_09303_),
    .B(_09253_));
 sg13g2_nand2_1 _18400_ (.Y(_09305_),
    .A(_09287_),
    .B(_09304_));
 sg13g2_nor2_1 _18401_ (.A(_09256_),
    .B(_04958_),
    .Y(_09306_));
 sg13g2_buf_2 _18402_ (.A(_09306_),
    .X(_09307_));
 sg13g2_nor2_1 _18403_ (.A(_09264_),
    .B(_06109_),
    .Y(_09308_));
 sg13g2_nor2_1 _18404_ (.A(_09307_),
    .B(_09308_),
    .Y(_09309_));
 sg13g2_nor2b_1 _18405_ (.A(_09305_),
    .B_N(_09309_),
    .Y(_09310_));
 sg13g2_nand2_1 _18406_ (.Y(_09311_),
    .A(_09267_),
    .B(_09310_));
 sg13g2_nor2_1 _18407_ (.A(_04261_),
    .B(_05990_),
    .Y(_09312_));
 sg13g2_nand2_1 _18408_ (.Y(_09313_),
    .A(_09311_),
    .B(_09312_));
 sg13g2_nand3_1 _18409_ (.B(_09254_),
    .C(_09266_),
    .A(_09232_),
    .Y(_09314_));
 sg13g2_nand3_1 _18410_ (.B(_09304_),
    .C(_09309_),
    .A(_09287_),
    .Y(_09315_));
 sg13g2_nor2_1 _18411_ (.A(net192),
    .B(_05990_),
    .Y(_09316_));
 sg13g2_nand3_1 _18412_ (.B(_09315_),
    .C(_09316_),
    .A(_09314_),
    .Y(_09317_));
 sg13g2_buf_1 _18413_ (.A(_09317_),
    .X(_09318_));
 sg13g2_nand2_1 _18414_ (.Y(_09319_),
    .A(_09313_),
    .B(_09318_));
 sg13g2_nand2_1 _18415_ (.Y(_09320_),
    .A(_09318_),
    .B(_05984_));
 sg13g2_nand2_1 _18416_ (.Y(_09321_),
    .A(_06004_),
    .B(_05983_));
 sg13g2_nand3_1 _18417_ (.B(_09320_),
    .C(_09321_),
    .A(_09319_),
    .Y(_09322_));
 sg13g2_nor2b_1 _18418_ (.A(_09187_),
    .B_N(_06000_),
    .Y(_09323_));
 sg13g2_nand3_1 _18419_ (.B(_09304_),
    .C(_09323_),
    .A(_09254_),
    .Y(_09324_));
 sg13g2_nand2_1 _18420_ (.Y(_09325_),
    .A(_09324_),
    .B(_05990_));
 sg13g2_nand3_1 _18421_ (.B(_09269_),
    .C(_07578_),
    .A(_09212_),
    .Y(_09326_));
 sg13g2_nand2_1 _18422_ (.Y(_09327_),
    .A(_09326_),
    .B(_05990_));
 sg13g2_nand2_1 _18423_ (.Y(_09328_),
    .A(_09325_),
    .B(_09327_));
 sg13g2_nand2_1 _18424_ (.Y(_09329_),
    .A(_09328_),
    .B(_06005_));
 sg13g2_nand3_1 _18425_ (.B(_05990_),
    .C(_06002_),
    .A(_09324_),
    .Y(_09330_));
 sg13g2_nand2_1 _18426_ (.Y(_09331_),
    .A(_09329_),
    .B(_09330_));
 sg13g2_nand2_1 _18427_ (.Y(_09332_),
    .A(_09331_),
    .B(net183));
 sg13g2_inv_1 _18428_ (.Y(_09333_),
    .A(\b.gen_square[8].sq.mask ));
 sg13g2_a21oi_1 _18429_ (.A1(_09322_),
    .A2(_09332_),
    .Y(_09334_),
    .B1(_09333_));
 sg13g2_nand2_1 _18430_ (.Y(_09335_),
    .A(_09241_),
    .B(_09251_));
 sg13g2_nand2_1 _18431_ (.Y(_09336_),
    .A(_08336_),
    .B(_05677_));
 sg13g2_nand2_1 _18432_ (.Y(_09337_),
    .A(_09336_),
    .B(_08201_));
 sg13g2_nand2_1 _18433_ (.Y(_09338_),
    .A(_09337_),
    .B(_05646_));
 sg13g2_inv_1 _18434_ (.Y(_09339_),
    .A(_05718_));
 sg13g2_nand2_1 _18435_ (.Y(_09340_),
    .A(_09338_),
    .B(_09339_));
 sg13g2_nand2_1 _18436_ (.Y(_09341_),
    .A(_09340_),
    .B(_05709_));
 sg13g2_nand2_1 _18437_ (.Y(_09342_),
    .A(_09341_),
    .B(_05712_));
 sg13g2_nand2_1 _18438_ (.Y(_09343_),
    .A(_08308_),
    .B(_05677_));
 sg13g2_nand2_1 _18439_ (.Y(_09344_),
    .A(_09343_),
    .B(_05687_));
 sg13g2_nand2_1 _18440_ (.Y(_09345_),
    .A(_09344_),
    .B(_05646_));
 sg13g2_nand2_1 _18441_ (.Y(_09346_),
    .A(_09345_),
    .B(_05656_));
 sg13g2_nand2_1 _18442_ (.Y(_09347_),
    .A(_09346_),
    .B(_05709_));
 sg13g2_nand2_1 _18443_ (.Y(_09348_),
    .A(_09347_),
    .B(_05627_));
 sg13g2_inv_2 _18444_ (.Y(_09349_),
    .A(_09348_));
 sg13g2_nand2_1 _18445_ (.Y(_09350_),
    .A(_09342_),
    .B(_09349_));
 sg13g2_inv_1 _18446_ (.Y(_09351_),
    .A(_05612_));
 sg13g2_a22oi_1 _18447_ (.Y(_09352_),
    .B1(_03558_),
    .B2(_09351_),
    .A2(_04018_),
    .A1(_06009_));
 sg13g2_nand3_1 _18448_ (.B(_09350_),
    .C(_09352_),
    .A(_09335_),
    .Y(_09353_));
 sg13g2_nand2_1 _18449_ (.Y(_09354_),
    .A(_07989_),
    .B(_04815_));
 sg13g2_inv_1 _18450_ (.Y(_09355_),
    .A(_04962_));
 sg13g2_nand2_1 _18451_ (.Y(_09356_),
    .A(_09354_),
    .B(_09355_));
 sg13g2_nand2_1 _18452_ (.Y(_09357_),
    .A(_07878_),
    .B(_04927_));
 sg13g2_nand2_1 _18453_ (.Y(_09358_),
    .A(_09357_),
    .B(_04937_));
 sg13g2_nand2_1 _18454_ (.Y(_09359_),
    .A(_09358_),
    .B(_04897_));
 sg13g2_nand2_1 _18455_ (.Y(_09360_),
    .A(_09359_),
    .B(_04906_));
 sg13g2_nand2_1 _18456_ (.Y(_09361_),
    .A(_09360_),
    .B(_04815_));
 sg13g2_nand2_1 _18457_ (.Y(_09362_),
    .A(_09361_),
    .B(_04877_));
 sg13g2_inv_1 _18458_ (.Y(_09363_),
    .A(_09362_));
 sg13g2_nand2_1 _18459_ (.Y(_09364_),
    .A(_09356_),
    .B(_09363_));
 sg13g2_nand3_1 _18460_ (.B(net58),
    .C(_07882_),
    .A(_07881_),
    .Y(_09365_));
 sg13g2_nand2_1 _18461_ (.Y(_09366_),
    .A(_06203_),
    .B(\b.gen_square[36].sq.color ));
 sg13g2_nand3_1 _18462_ (.B(_04897_),
    .C(_09366_),
    .A(_09365_),
    .Y(_09367_));
 sg13g2_inv_1 _18463_ (.Y(_09368_),
    .A(_04897_));
 sg13g2_nand2_1 _18464_ (.Y(_09369_),
    .A(_09368_),
    .B(_03639_));
 sg13g2_nand3_1 _18465_ (.B(_04815_),
    .C(_09369_),
    .A(_09367_),
    .Y(_09370_));
 sg13g2_a21oi_2 _18466_ (.B1(_04813_),
    .Y(_09371_),
    .A2(_04808_),
    .A1(_04873_));
 sg13g2_inv_1 _18467_ (.Y(_09372_),
    .A(_09371_));
 sg13g2_nor2_1 _18468_ (.A(_03535_),
    .B(_04815_),
    .Y(_09373_));
 sg13g2_inv_1 _18469_ (.Y(_09374_),
    .A(_09373_));
 sg13g2_nand3_1 _18470_ (.B(_09372_),
    .C(_09374_),
    .A(_09370_),
    .Y(_09375_));
 sg13g2_a21oi_2 _18471_ (.B1(_05713_),
    .Y(_09376_),
    .A2(_05709_),
    .A1(_06889_));
 sg13g2_nor2_1 _18472_ (.A(_09195_),
    .B(_09376_),
    .Y(_09377_));
 sg13g2_a21oi_2 _18473_ (.B1(_06331_),
    .Y(_09378_),
    .A2(_06326_),
    .A1(_06357_));
 sg13g2_o21ai_1 _18474_ (.B1(_09300_),
    .Y(_09379_),
    .A1(_08901_),
    .A2(_09273_));
 sg13g2_buf_1 _18475_ (.A(_09379_),
    .X(_09380_));
 sg13g2_nor2_1 _18476_ (.A(_09378_),
    .B(_09380_),
    .Y(_09381_));
 sg13g2_nor2_1 _18477_ (.A(_09377_),
    .B(_09381_),
    .Y(_09382_));
 sg13g2_a21oi_2 _18478_ (.B1(_06419_),
    .Y(_09383_),
    .A2(_06352_),
    .A1(_06341_));
 sg13g2_nor2_1 _18479_ (.A(_09383_),
    .B(_06422_),
    .Y(_09384_));
 sg13g2_nor2_1 _18480_ (.A(_08655_),
    .B(_06422_),
    .Y(_09385_));
 sg13g2_inv_1 _18481_ (.Y(_09386_),
    .A(_04858_));
 sg13g2_nor2_1 _18482_ (.A(_06888_),
    .B(_06876_),
    .Y(_09387_));
 sg13g2_a21o_1 _18483_ (.A2(_09386_),
    .A1(_04953_),
    .B1(_09387_),
    .X(_09388_));
 sg13g2_nand2_1 _18484_ (.Y(_09389_),
    .A(_08107_),
    .B(_07938_));
 sg13g2_nor3_1 _18485_ (.A(_08109_),
    .B(_09129_),
    .C(_09389_),
    .Y(_09390_));
 sg13g2_nor2_1 _18486_ (.A(_09264_),
    .B(_06888_),
    .Y(_09391_));
 sg13g2_inv_1 _18487_ (.Y(_09392_),
    .A(_05988_));
 sg13g2_nor2_1 _18488_ (.A(_06001_),
    .B(_04313_),
    .Y(_09393_));
 sg13g2_a21oi_1 _18489_ (.A1(_09392_),
    .A2(_09393_),
    .Y(_09394_),
    .B1(_05993_));
 sg13g2_buf_1 _18490_ (.A(_09394_),
    .X(_09395_));
 sg13g2_nor2_1 _18491_ (.A(_09395_),
    .B(_07179_),
    .Y(_09396_));
 sg13g2_nor2_1 _18492_ (.A(_09391_),
    .B(_09396_),
    .Y(_09397_));
 sg13g2_nand3_1 _18493_ (.B(_09397_),
    .C(_09226_),
    .A(_09390_),
    .Y(_09398_));
 sg13g2_nor4_1 _18494_ (.A(_09384_),
    .B(_09385_),
    .C(_09388_),
    .D(_09398_),
    .Y(_09399_));
 sg13g2_nand4_1 _18495_ (.B(_09375_),
    .C(_09382_),
    .A(_09364_),
    .Y(_09400_),
    .D(_09399_));
 sg13g2_nor2_1 _18496_ (.A(_09353_),
    .B(_09400_),
    .Y(_09401_));
 sg13g2_nand2_1 _18497_ (.Y(_09402_),
    .A(_04863_),
    .B(_01968_));
 sg13g2_nand2_1 _18498_ (.Y(_09403_),
    .A(_09301_),
    .B(_09251_));
 sg13g2_inv_4 _18499_ (.A(_09376_),
    .Y(_09404_));
 sg13g2_a21oi_2 _18500_ (.B1(_04962_),
    .Y(_09405_),
    .A2(_04815_),
    .A1(_09404_));
 sg13g2_inv_2 _18501_ (.Y(_09406_),
    .A(_09405_));
 sg13g2_nor2_1 _18502_ (.A(_09371_),
    .B(_09406_),
    .Y(_09407_));
 sg13g2_nor2_1 _18503_ (.A(_06008_),
    .B(_07180_),
    .Y(_09408_));
 sg13g2_nor2_1 _18504_ (.A(_09383_),
    .B(_06423_),
    .Y(_09409_));
 sg13g2_nor2_1 _18505_ (.A(_09409_),
    .B(_09279_),
    .Y(_09410_));
 sg13g2_inv_2 _18506_ (.Y(_09411_),
    .A(_09410_));
 sg13g2_nor3_1 _18507_ (.A(_09276_),
    .B(_09408_),
    .C(_09411_),
    .Y(_09412_));
 sg13g2_nor2_1 _18508_ (.A(_06889_),
    .B(_06876_),
    .Y(_09413_));
 sg13g2_nor2_1 _18509_ (.A(_08655_),
    .B(_06423_),
    .Y(_09414_));
 sg13g2_nor2_1 _18510_ (.A(_09413_),
    .B(_09414_),
    .Y(_09415_));
 sg13g2_nand2_1 _18511_ (.Y(_09416_),
    .A(_09386_),
    .B(_09222_));
 sg13g2_nor2_1 _18512_ (.A(_09264_),
    .B(_06889_),
    .Y(_09417_));
 sg13g2_nand2b_1 _18513_ (.Y(_09418_),
    .B(_07179_),
    .A_N(_09395_));
 sg13g2_nand2b_1 _18514_ (.Y(_09419_),
    .B(_09418_),
    .A_N(_09417_));
 sg13g2_nor2_1 _18515_ (.A(_08052_),
    .B(_09149_),
    .Y(_09420_));
 sg13g2_nand2_1 _18516_ (.Y(_09421_),
    .A(_09420_),
    .B(_07924_));
 sg13g2_nor2_1 _18517_ (.A(_09419_),
    .B(_09421_),
    .Y(_09422_));
 sg13g2_nand4_1 _18518_ (.B(_09415_),
    .C(_09416_),
    .A(_09412_),
    .Y(_09423_),
    .D(_09422_));
 sg13g2_nor2_1 _18519_ (.A(_09407_),
    .B(_09423_),
    .Y(_09424_));
 sg13g2_nand2_1 _18520_ (.Y(_09425_),
    .A(_09351_),
    .B(_03557_));
 sg13g2_nand3_1 _18521_ (.B(_09424_),
    .C(_09425_),
    .A(_09403_),
    .Y(_09426_));
 sg13g2_nand3_1 _18522_ (.B(_05712_),
    .C(_09341_),
    .A(_09349_),
    .Y(_09427_));
 sg13g2_a21oi_2 _18523_ (.B1(_06426_),
    .Y(_09428_),
    .A2(_06333_),
    .A1(_06805_));
 sg13g2_inv_2 _18524_ (.Y(_09429_),
    .A(_09428_));
 sg13g2_nor2_1 _18525_ (.A(_09378_),
    .B(_09429_),
    .Y(_09430_));
 sg13g2_buf_1 _18526_ (.A(_09430_),
    .X(_09431_));
 sg13g2_nor2_1 _18527_ (.A(_09275_),
    .B(_09431_),
    .Y(_09432_));
 sg13g2_nand2_1 _18528_ (.Y(_09433_),
    .A(_09370_),
    .B(_09374_));
 sg13g2_nand2_1 _18529_ (.Y(_09434_),
    .A(_09433_),
    .B(_09363_));
 sg13g2_nand3_1 _18530_ (.B(_09432_),
    .C(_09434_),
    .A(_09427_),
    .Y(_09435_));
 sg13g2_nor2_1 _18531_ (.A(_09426_),
    .B(_09435_),
    .Y(_09436_));
 sg13g2_nor2_1 _18532_ (.A(_09402_),
    .B(_09436_),
    .Y(_09437_));
 sg13g2_nand2b_1 _18533_ (.Y(_09438_),
    .B(_09437_),
    .A_N(_09401_));
 sg13g2_nor2b_1 _18534_ (.A(_04859_),
    .B_N(_04821_),
    .Y(_09439_));
 sg13g2_a21oi_1 _18535_ (.A1(_09438_),
    .A2(_04822_),
    .Y(_09440_),
    .B1(_09439_));
 sg13g2_nand2_1 _18536_ (.Y(_09441_),
    .A(_09401_),
    .B(_09436_));
 sg13g2_nor2_1 _18537_ (.A(_04261_),
    .B(net132),
    .Y(_09442_));
 sg13g2_nand2_1 _18538_ (.Y(_09443_),
    .A(_09441_),
    .B(_09442_));
 sg13g2_nand2_1 _18539_ (.Y(_09444_),
    .A(_09443_),
    .B(_09438_));
 sg13g2_nand2_1 _18540_ (.Y(_09445_),
    .A(_09440_),
    .B(_09444_));
 sg13g2_o21ai_1 _18541_ (.B1(_09425_),
    .Y(_09446_),
    .A1(_06008_),
    .A2(_07180_));
 sg13g2_nand2_1 _18542_ (.Y(_09447_),
    .A(_09427_),
    .B(_09403_));
 sg13g2_nor2_1 _18543_ (.A(_09446_),
    .B(_09447_),
    .Y(_09448_));
 sg13g2_nand2b_1 _18544_ (.Y(_09449_),
    .B(_09448_),
    .A_N(_09353_));
 sg13g2_nand2_1 _18545_ (.Y(_09450_),
    .A(_09449_),
    .B(net132));
 sg13g2_nor3_1 _18546_ (.A(_06875_),
    .B(_08654_),
    .C(_09386_),
    .Y(_09451_));
 sg13g2_nand3_1 _18547_ (.B(_09364_),
    .C(_09451_),
    .A(_09434_),
    .Y(_09452_));
 sg13g2_nand2_1 _18548_ (.Y(_09453_),
    .A(_09452_),
    .B(net132));
 sg13g2_nand2_1 _18549_ (.Y(_09454_),
    .A(_09450_),
    .B(_09453_));
 sg13g2_nand2_1 _18550_ (.Y(_09455_),
    .A(_09454_),
    .B(_04861_));
 sg13g2_nand3_1 _18551_ (.B(net132),
    .C(_05613_),
    .A(_09449_),
    .Y(_09456_));
 sg13g2_nand2_1 _18552_ (.Y(_09457_),
    .A(_09455_),
    .B(_09456_));
 sg13g2_nor2_1 _18553_ (.A(_02023_),
    .B(_04827_),
    .Y(_09458_));
 sg13g2_nand2_1 _18554_ (.Y(_09459_),
    .A(_09457_),
    .B(_09458_));
 sg13g2_nand2_1 _18555_ (.Y(_09460_),
    .A(_09445_),
    .B(_09459_));
 sg13g2_buf_2 _18556_ (.A(\b.gen_square[9].sq.mask ),
    .X(_09461_));
 sg13g2_nand2_1 _18557_ (.Y(_09462_),
    .A(_09460_),
    .B(_09461_));
 sg13g2_nand2_1 _18558_ (.Y(_09463_),
    .A(_09334_),
    .B(_09462_));
 sg13g2_nand2_1 _18559_ (.Y(_09464_),
    .A(_09322_),
    .B(_09332_));
 sg13g2_nand2_1 _18560_ (.Y(_09465_),
    .A(_09464_),
    .B(\b.gen_square[8].sq.mask ));
 sg13g2_inv_1 _18561_ (.Y(_09466_),
    .A(_09461_));
 sg13g2_a21oi_1 _18562_ (.A1(_09445_),
    .A2(_09459_),
    .Y(_09467_),
    .B1(_09466_));
 sg13g2_nand2_1 _18563_ (.Y(_09468_),
    .A(_09465_),
    .B(_09467_));
 sg13g2_nor2b_1 _18564_ (.A(_09327_),
    .B_N(_07188_),
    .Y(_09469_));
 sg13g2_nor2_1 _18565_ (.A(_09392_),
    .B(_09469_),
    .Y(_09470_));
 sg13g2_nand2_1 _18566_ (.Y(_09471_),
    .A(_09329_),
    .B(_09470_));
 sg13g2_inv_1 _18567_ (.Y(_09472_),
    .A(_09224_));
 sg13g2_nor4_1 _18568_ (.A(_05988_),
    .B(_09472_),
    .C(_09220_),
    .D(_09275_),
    .Y(_09473_));
 sg13g2_and4_1 _18569_ (.A(_09200_),
    .B(_09309_),
    .C(_09266_),
    .D(_09473_),
    .X(_09474_));
 sg13g2_nor3_1 _18570_ (.A(net154),
    .B(_05991_),
    .C(_09474_),
    .Y(_09475_));
 sg13g2_nand2_1 _18571_ (.Y(_09476_),
    .A(_09471_),
    .B(_09475_));
 sg13g2_inv_1 _18572_ (.Y(_09477_),
    .A(_05982_));
 sg13g2_nand2_1 _18573_ (.Y(_09478_),
    .A(_09312_),
    .B(_09477_));
 sg13g2_o21ai_1 _18574_ (.B1(_09478_),
    .Y(_09479_),
    .A1(_04261_),
    .A2(_05985_));
 sg13g2_nor2_1 _18575_ (.A(_05982_),
    .B(_09318_),
    .Y(_09480_));
 sg13g2_a21oi_1 _18576_ (.A1(_09311_),
    .A2(_09479_),
    .Y(_09481_),
    .B1(_09480_));
 sg13g2_a21oi_2 _18577_ (.B1(_09333_),
    .Y(_09482_),
    .A2(_09481_),
    .A1(_09476_));
 sg13g2_nor2b_1 _18578_ (.A(_09453_),
    .B_N(_04862_),
    .Y(_09483_));
 sg13g2_nor2_1 _18579_ (.A(_04827_),
    .B(_09483_),
    .Y(_09484_));
 sg13g2_nand2_1 _18580_ (.Y(_09485_),
    .A(_09455_),
    .B(_09484_));
 sg13g2_inv_1 _18581_ (.Y(_09486_),
    .A(_09407_));
 sg13g2_nor2_1 _18582_ (.A(_09384_),
    .B(_09225_),
    .Y(_09487_));
 sg13g2_nand4_1 _18583_ (.B(_09264_),
    .C(_09395_),
    .A(_09487_),
    .Y(_09488_),
    .D(_09221_));
 sg13g2_nor2_1 _18584_ (.A(_09411_),
    .B(_09488_),
    .Y(_09489_));
 sg13g2_nand4_1 _18585_ (.B(_09486_),
    .C(_09382_),
    .A(_09375_),
    .Y(_09490_),
    .D(_09489_));
 sg13g2_nor4_1 _18586_ (.A(_04828_),
    .B(_09275_),
    .C(_09431_),
    .D(_09490_),
    .Y(_09491_));
 sg13g2_nor3_1 _18587_ (.A(net154),
    .B(_04829_),
    .C(_09491_),
    .Y(_09492_));
 sg13g2_nand2_1 _18588_ (.Y(_09493_),
    .A(_09485_),
    .B(_09492_));
 sg13g2_nand2_1 _18589_ (.Y(_09494_),
    .A(_04863_),
    .B(_04826_));
 sg13g2_a21oi_1 _18590_ (.A1(_09494_),
    .A2(_04823_),
    .Y(_09495_),
    .B1(_04261_));
 sg13g2_nor2_1 _18591_ (.A(_04820_),
    .B(_09438_),
    .Y(_09496_));
 sg13g2_a21oi_1 _18592_ (.A1(_09441_),
    .A2(_09495_),
    .Y(_09497_),
    .B1(_09496_));
 sg13g2_nand2_1 _18593_ (.Y(_09498_),
    .A(_09493_),
    .B(_09497_));
 sg13g2_nand2_1 _18594_ (.Y(_09499_),
    .A(_09498_),
    .B(_09461_));
 sg13g2_nand2_1 _18595_ (.Y(_09500_),
    .A(_09482_),
    .B(_09499_));
 sg13g2_nand3_1 _18596_ (.B(_09468_),
    .C(_09500_),
    .A(_09463_),
    .Y(_09501_));
 sg13g2_xnor2_1 _18597_ (.Y(_09502_),
    .A(_05979_),
    .B(_06003_));
 sg13g2_nor4_1 _18598_ (.A(_05979_),
    .B(_05981_),
    .C(_09477_),
    .D(_06001_),
    .Y(_09503_));
 sg13g2_nand2_1 _18599_ (.Y(_09504_),
    .A(_09217_),
    .B(_09284_));
 sg13g2_a21oi_1 _18600_ (.A1(_09503_),
    .A2(_09504_),
    .Y(_09505_),
    .B1(_09469_));
 sg13g2_nor3_1 _18601_ (.A(_02023_),
    .B(_09392_),
    .C(_09505_),
    .Y(_09506_));
 sg13g2_a21oi_1 _18602_ (.A1(_09319_),
    .A2(_09502_),
    .Y(_09507_),
    .B1(_09506_));
 sg13g2_a21oi_1 _18603_ (.A1(_09507_),
    .A2(_09332_),
    .Y(_09508_),
    .B1(_09333_));
 sg13g2_nor3_1 _18604_ (.A(_04817_),
    .B(_04819_),
    .C(_04826_),
    .Y(_09509_));
 sg13g2_nand2_1 _18605_ (.Y(_09510_),
    .A(_04825_),
    .B(_09509_));
 sg13g2_inv_1 _18606_ (.Y(_09511_),
    .A(_09510_));
 sg13g2_nand2b_1 _18607_ (.Y(_09512_),
    .B(_09390_),
    .A_N(_09421_));
 sg13g2_a21o_1 _18608_ (.A2(_09512_),
    .A1(_09511_),
    .B1(_09483_),
    .X(_09513_));
 sg13g2_xnor2_1 _18609_ (.Y(_09514_),
    .A(_04817_),
    .B(_04859_));
 sg13g2_a22oi_1 _18610_ (.Y(_09515_),
    .B1(_09514_),
    .B2(_09444_),
    .A2(_09458_),
    .A1(_09513_));
 sg13g2_nand2_1 _18611_ (.Y(_09516_),
    .A(_09515_),
    .B(_09459_));
 sg13g2_nand2_1 _18612_ (.Y(_09517_),
    .A(_09516_),
    .B(_09461_));
 sg13g2_nor2_1 _18613_ (.A(_09508_),
    .B(_09517_),
    .Y(_09518_));
 sg13g2_nor2b_1 _18614_ (.A(_09518_),
    .B_N(_09468_),
    .Y(_09519_));
 sg13g2_inv_1 _18615_ (.Y(_09520_),
    .A(_09508_));
 sg13g2_nor2b_1 _18616_ (.A(_09520_),
    .B_N(_09517_),
    .Y(_09521_));
 sg13g2_a21oi_1 _18617_ (.A1(_09501_),
    .A2(_09519_),
    .Y(_09522_),
    .B1(_09521_));
 sg13g2_xnor2_1 _18618_ (.Y(_09523_),
    .A(_09499_),
    .B(_09482_));
 sg13g2_nand2_1 _18619_ (.Y(_09524_),
    .A(_09463_),
    .B(_09468_));
 sg13g2_nor2_1 _18620_ (.A(_09523_),
    .B(_09524_),
    .Y(_09525_));
 sg13g2_nor2_1 _18621_ (.A(_09518_),
    .B(_09521_),
    .Y(_09526_));
 sg13g2_nand2_1 _18622_ (.Y(_09527_),
    .A(_09525_),
    .B(_09526_));
 sg13g2_nand2_1 _18623_ (.Y(_09528_),
    .A(_09522_),
    .B(_09527_));
 sg13g2_nand2_1 _18624_ (.Y(_09529_),
    .A(_09528_),
    .B(_09334_));
 sg13g2_nand3_1 _18625_ (.B(_09467_),
    .C(_09527_),
    .A(_09522_),
    .Y(_09530_));
 sg13g2_nand2_1 _18626_ (.Y(_09531_),
    .A(_09529_),
    .B(_09530_));
 sg13g2_nor2_1 _18627_ (.A(_09256_),
    .B(_04957_),
    .Y(_09532_));
 sg13g2_buf_2 _18628_ (.A(_09532_),
    .X(_09533_));
 sg13g2_inv_1 _18629_ (.Y(_09534_),
    .A(_09377_));
 sg13g2_inv_1 _18630_ (.Y(_09535_),
    .A(_06546_));
 sg13g2_a21oi_2 _18631_ (.B1(_06801_),
    .Y(_09536_),
    .A2(_06542_),
    .A1(_09535_));
 sg13g2_nor2_1 _18632_ (.A(_09536_),
    .B(_06804_),
    .Y(_09537_));
 sg13g2_inv_1 _18633_ (.Y(_09538_),
    .A(_09537_));
 sg13g2_nand3_1 _18634_ (.B(_09538_),
    .C(_09487_),
    .A(_09534_),
    .Y(_09539_));
 sg13g2_a21oi_1 _18635_ (.A1(_06523_),
    .A2(_06557_),
    .Y(_09540_),
    .B1(_06527_));
 sg13g2_buf_2 _18636_ (.A(_09540_),
    .X(_09541_));
 sg13g2_nor2_1 _18637_ (.A(_09541_),
    .B(_09297_),
    .Y(_09542_));
 sg13g2_nor3_1 _18638_ (.A(_09533_),
    .B(_09539_),
    .C(_09542_),
    .Y(_09543_));
 sg13g2_nor2_2 _18639_ (.A(_09371_),
    .B(_09405_),
    .Y(_09544_));
 sg13g2_inv_1 _18640_ (.Y(_09545_),
    .A(_09544_));
 sg13g2_inv_1 _18641_ (.Y(_09546_),
    .A(_06571_));
 sg13g2_a21oi_2 _18642_ (.B1(_06577_),
    .Y(_09547_),
    .A2(_06582_),
    .A1(_09546_));
 sg13g2_nor2_1 _18643_ (.A(_03548_),
    .B(net35),
    .Y(_09548_));
 sg13g2_nand2_1 _18644_ (.Y(_09549_),
    .A(_07728_),
    .B(_06696_));
 sg13g2_nand2_1 _18645_ (.Y(_09550_),
    .A(_07952_),
    .B(\b.gen_square[37].sq.color ));
 sg13g2_nand3_1 _18646_ (.B(net55),
    .C(_09550_),
    .A(_09549_),
    .Y(_09551_));
 sg13g2_buf_1 _18647_ (.A(_09551_),
    .X(_09552_));
 sg13g2_nand2_1 _18648_ (.Y(_09553_),
    .A(_07574_),
    .B(_03650_));
 sg13g2_nand3_1 _18649_ (.B(net35),
    .C(_09553_),
    .A(_09552_),
    .Y(_09554_));
 sg13g2_nand2b_1 _18650_ (.Y(_09555_),
    .B(_09554_),
    .A_N(_09548_));
 sg13g2_inv_1 _18651_ (.Y(_09556_),
    .A(_09555_));
 sg13g2_nand2b_1 _18652_ (.Y(_09557_),
    .B(_09556_),
    .A_N(_09547_));
 sg13g2_nand3_1 _18653_ (.B(_09545_),
    .C(_09557_),
    .A(_09543_),
    .Y(_09558_));
 sg13g2_inv_1 _18654_ (.Y(_09559_),
    .A(_09558_));
 sg13g2_nor2_1 _18655_ (.A(_08796_),
    .B(_06804_),
    .Y(_09560_));
 sg13g2_inv_1 _18656_ (.Y(_09561_),
    .A(_09273_));
 sg13g2_a21oi_1 _18657_ (.A1(_06750_),
    .A2(net38),
    .Y(_09562_),
    .B1(_07196_));
 sg13g2_nor2b_1 _18658_ (.A(_09561_),
    .B_N(_09562_),
    .Y(_09563_));
 sg13g2_nand2_1 _18659_ (.Y(_09564_),
    .A(_07767_),
    .B(_06696_));
 sg13g2_nand2_1 _18660_ (.Y(_09565_),
    .A(_09564_),
    .B(_06706_));
 sg13g2_nand2_1 _18661_ (.Y(_09566_),
    .A(_09565_),
    .B(_05346_));
 sg13g2_nand2_1 _18662_ (.Y(_09567_),
    .A(_09566_),
    .B(_05356_));
 sg13g2_nand2_1 _18663_ (.Y(_09568_),
    .A(_09567_),
    .B(_06579_));
 sg13g2_nand2_1 _18664_ (.Y(_09569_),
    .A(_09568_),
    .B(_07589_));
 sg13g2_nand2_1 _18665_ (.Y(_09570_),
    .A(_07806_),
    .B(_06579_));
 sg13g2_nand2b_1 _18666_ (.Y(_09571_),
    .B(_09570_),
    .A_N(_06812_));
 sg13g2_nor2b_1 _18667_ (.A(_09569_),
    .B_N(_09571_),
    .Y(_09572_));
 sg13g2_nor4_1 _18668_ (.A(_09560_),
    .B(_09563_),
    .C(_09228_),
    .D(_09572_),
    .Y(_09573_));
 sg13g2_nand4_1 _18669_ (.B(_04837_),
    .C(_04851_),
    .A(_04843_),
    .Y(_09574_),
    .D(_04839_));
 sg13g2_o21ai_1 _18670_ (.B1(_04856_),
    .Y(_09575_),
    .A1(net61),
    .A2(_09574_));
 sg13g2_nand2_1 _18671_ (.Y(_09576_),
    .A(_09575_),
    .B(_01770_));
 sg13g2_inv_1 _18672_ (.Y(_09577_),
    .A(_09576_));
 sg13g2_inv_1 _18673_ (.Y(_09578_),
    .A(_08251_));
 sg13g2_nor4_2 _18674_ (.A(_08418_),
    .B(_09577_),
    .C(_09578_),
    .Y(_09579_),
    .D(_09010_));
 sg13g2_nand3_1 _18675_ (.B(_09573_),
    .C(_09579_),
    .A(_09559_),
    .Y(_09580_));
 sg13g2_a21oi_1 _18676_ (.A1(_05761_),
    .A2(_05844_),
    .Y(_09581_),
    .B1(_05963_));
 sg13g2_o21ai_1 _18677_ (.B1(_09203_),
    .Y(_09582_),
    .A1(_08277_),
    .A2(_09581_));
 sg13g2_buf_1 _18678_ (.A(_09582_),
    .X(_09583_));
 sg13g2_a21oi_1 _18679_ (.A1(_09583_),
    .A2(net29),
    .Y(_09584_),
    .B1(_04962_));
 sg13g2_o21ai_1 _18680_ (.B1(_06407_),
    .Y(_09585_),
    .A1(_05845_),
    .A2(_08088_));
 sg13g2_a21oi_1 _18681_ (.A1(_09585_),
    .A2(_06391_),
    .Y(_09586_),
    .B1(_06402_));
 sg13g2_o21ai_1 _18682_ (.B1(_06369_),
    .Y(_09587_),
    .A1(_04816_),
    .A2(_09586_));
 sg13g2_inv_2 _18683_ (.Y(_09588_),
    .A(_09587_));
 sg13g2_nand2b_1 _18684_ (.Y(_09589_),
    .B(_09588_),
    .A_N(_09584_));
 sg13g2_a22oi_1 _18685_ (.Y(_09590_),
    .B1(_08902_),
    .B2(_08911_),
    .A2(_06354_),
    .A1(_03669_));
 sg13g2_inv_1 _18686_ (.Y(_09591_),
    .A(_09250_));
 sg13g2_nand2_1 _18687_ (.Y(_09592_),
    .A(_09238_),
    .B(_09591_));
 sg13g2_nand3_1 _18688_ (.B(_09590_),
    .C(_09592_),
    .A(_09589_),
    .Y(_09593_));
 sg13g2_nor2_1 _18689_ (.A(_09580_),
    .B(_09593_),
    .Y(_09594_));
 sg13g2_inv_1 _18690_ (.Y(_09595_),
    .A(_09594_));
 sg13g2_nand2_1 _18691_ (.Y(_09596_),
    .A(_09588_),
    .B(_09584_));
 sg13g2_a22oi_1 _18692_ (.Y(_09597_),
    .B1(_08902_),
    .B2(_08910_),
    .A2(_06422_),
    .A1(_06354_));
 sg13g2_nand2_1 _18693_ (.Y(_09598_),
    .A(_09591_),
    .B(_09297_));
 sg13g2_nand3_1 _18694_ (.B(_09597_),
    .C(_09598_),
    .A(_09596_),
    .Y(_09599_));
 sg13g2_inv_2 _18695_ (.Y(_09600_),
    .A(_09599_));
 sg13g2_nor2_1 _18696_ (.A(_08796_),
    .B(_06805_),
    .Y(_09601_));
 sg13g2_a21oi_1 _18697_ (.A1(_09561_),
    .A2(_09562_),
    .Y(_09602_),
    .B1(_09278_));
 sg13g2_o21ai_1 _18698_ (.B1(_09602_),
    .Y(_09603_),
    .A1(_09569_),
    .A2(_09556_));
 sg13g2_nor2_1 _18699_ (.A(_09601_),
    .B(_09603_),
    .Y(_09604_));
 sg13g2_inv_1 _18700_ (.Y(_09605_),
    .A(_08972_));
 sg13g2_a21o_1 _18701_ (.A2(_09575_),
    .A1(_01759_),
    .B1(_07835_),
    .X(_09606_));
 sg13g2_nor4_1 _18702_ (.A(_08423_),
    .B(_08273_),
    .C(_09605_),
    .D(_09606_),
    .Y(_09607_));
 sg13g2_nor2_2 _18703_ (.A(_09541_),
    .B(_06810_),
    .Y(_09608_));
 sg13g2_nor2_1 _18704_ (.A(_09536_),
    .B(_06805_),
    .Y(_09609_));
 sg13g2_nor4_1 _18705_ (.A(_09609_),
    .B(_09275_),
    .C(_09411_),
    .D(_09307_),
    .Y(_09610_));
 sg13g2_nor2_2 _18706_ (.A(_09547_),
    .B(_06814_),
    .Y(_09611_));
 sg13g2_inv_4 _18707_ (.A(_09611_),
    .Y(_09612_));
 sg13g2_nand2_1 _18708_ (.Y(_09613_),
    .A(_09610_),
    .B(_09612_));
 sg13g2_nor3_1 _18709_ (.A(_09407_),
    .B(_09608_),
    .C(_09613_),
    .Y(_09614_));
 sg13g2_nand4_1 _18710_ (.B(_09604_),
    .C(_09607_),
    .A(_09600_),
    .Y(_09615_),
    .D(_09614_));
 sg13g2_nor2_1 _18711_ (.A(_09595_),
    .B(_09615_),
    .Y(_09616_));
 sg13g2_inv_2 _18712_ (.Y(_09617_),
    .A(_09616_));
 sg13g2_nand3_1 _18713_ (.B(_04044_),
    .C(_06356_),
    .A(_09617_),
    .Y(_09618_));
 sg13g2_nand4_1 _18714_ (.B(net215),
    .C(_06356_),
    .A(_09615_),
    .Y(_09619_),
    .D(_09595_));
 sg13g2_buf_1 _18715_ (.A(_09619_),
    .X(_09620_));
 sg13g2_nand2_1 _18716_ (.Y(_09621_),
    .A(_09618_),
    .B(_09620_));
 sg13g2_nand2_1 _18717_ (.Y(_09622_),
    .A(_09620_),
    .B(_06321_));
 sg13g2_nand2b_1 _18718_ (.Y(_09623_),
    .B(_06320_),
    .A_N(_06358_));
 sg13g2_nand3_1 _18719_ (.B(_09622_),
    .C(_09623_),
    .A(_09621_),
    .Y(_09624_));
 sg13g2_o21ai_1 _18720_ (.B1(_06324_),
    .Y(_09625_),
    .A1(_09599_),
    .A2(_09593_));
 sg13g2_nor3_1 _18721_ (.A(_06316_),
    .B(_06320_),
    .C(_09625_),
    .Y(_09626_));
 sg13g2_a21o_1 _18722_ (.A2(_09604_),
    .A1(_09573_),
    .B1(_06356_),
    .X(_09627_));
 sg13g2_a21o_1 _18723_ (.A2(_09627_),
    .A1(_09625_),
    .B1(_06359_),
    .X(_09628_));
 sg13g2_nand2b_1 _18724_ (.Y(_09629_),
    .B(_09628_),
    .A_N(_09626_));
 sg13g2_nand2_1 _18725_ (.Y(_09630_),
    .A(_09629_),
    .B(net183));
 sg13g2_nand2_1 _18726_ (.Y(_09631_),
    .A(_09624_),
    .B(_09630_));
 sg13g2_buf_2 _18727_ (.A(\b.gen_square[10].sq.mask ),
    .X(_09632_));
 sg13g2_nand2_1 _18728_ (.Y(_09633_),
    .A(_09631_),
    .B(_09632_));
 sg13g2_nor2_1 _18729_ (.A(net154),
    .B(_06326_),
    .Y(_09634_));
 sg13g2_nor3_1 _18730_ (.A(_06316_),
    .B(_06318_),
    .C(_06325_),
    .Y(_09635_));
 sg13g2_nand2_1 _18731_ (.Y(_09636_),
    .A(_06324_),
    .B(_09635_));
 sg13g2_a21oi_1 _18732_ (.A1(_09607_),
    .A2(_09579_),
    .Y(_09637_),
    .B1(_09636_));
 sg13g2_or2_1 _18733_ (.X(_09638_),
    .B(_09627_),
    .A(_07579_));
 sg13g2_nand2b_1 _18734_ (.Y(_09639_),
    .B(_09638_),
    .A_N(_09637_));
 sg13g2_xnor2_1 _18735_ (.Y(_09640_),
    .A(_06316_),
    .B(_06358_));
 sg13g2_a22oi_1 _18736_ (.Y(_09641_),
    .B1(_09640_),
    .B2(_09621_),
    .A2(_09639_),
    .A1(_09634_));
 sg13g2_nand2_1 _18737_ (.Y(_09642_),
    .A(_09641_),
    .B(_09630_));
 sg13g2_nand2_1 _18738_ (.Y(_09643_),
    .A(_09520_),
    .B(_09517_));
 sg13g2_inv_2 _18739_ (.Y(_09644_),
    .A(_09643_));
 sg13g2_a21oi_1 _18740_ (.A1(_09642_),
    .A2(_09632_),
    .Y(_09645_),
    .B1(_09644_));
 sg13g2_a21oi_1 _18741_ (.A1(_09531_),
    .A2(_09633_),
    .Y(_09646_),
    .B1(_09645_));
 sg13g2_nand3b_1 _18742_ (.B(_09522_),
    .C(_09527_),
    .Y(_09647_),
    .A_N(_09499_));
 sg13g2_nand2_1 _18743_ (.Y(_09648_),
    .A(_09528_),
    .B(_09482_));
 sg13g2_a21oi_1 _18744_ (.A1(_09559_),
    .A2(_09614_),
    .Y(_09649_),
    .B1(_06356_));
 sg13g2_nand3_1 _18745_ (.B(_06327_),
    .C(_09638_),
    .A(_09628_),
    .Y(_09650_));
 sg13g2_o21ai_1 _18746_ (.B1(_09650_),
    .Y(_09651_),
    .A1(_06327_),
    .A2(_09649_));
 sg13g2_a21oi_1 _18747_ (.A1(_06356_),
    .A2(_06325_),
    .Y(_09652_),
    .B1(_06321_));
 sg13g2_nor3_1 _18748_ (.A(net158),
    .B(_09652_),
    .C(_09616_),
    .Y(_09653_));
 sg13g2_nor2_1 _18749_ (.A(_06319_),
    .B(_09620_),
    .Y(_09654_));
 sg13g2_nor2_1 _18750_ (.A(_09653_),
    .B(_09654_),
    .Y(_09655_));
 sg13g2_o21ai_1 _18751_ (.B1(_09655_),
    .Y(_09656_),
    .A1(net154),
    .A2(_09651_));
 sg13g2_nand2_1 _18752_ (.Y(_09657_),
    .A(_09656_),
    .B(_09632_));
 sg13g2_inv_1 _18753_ (.Y(_09658_),
    .A(_09657_));
 sg13g2_nand3_1 _18754_ (.B(_09648_),
    .C(_09658_),
    .A(_09647_),
    .Y(_09659_));
 sg13g2_inv_2 _18755_ (.Y(_09660_),
    .A(_09633_));
 sg13g2_nand3_1 _18756_ (.B(_09530_),
    .C(_09660_),
    .A(_09529_),
    .Y(_09661_));
 sg13g2_nand2_1 _18757_ (.Y(_09662_),
    .A(_09659_),
    .B(_09661_));
 sg13g2_nand2_1 _18758_ (.Y(_09663_),
    .A(_09646_),
    .B(_09662_));
 sg13g2_nand3_1 _18759_ (.B(_09632_),
    .C(_09644_),
    .A(_09642_),
    .Y(_09664_));
 sg13g2_buf_1 _18760_ (.A(_09664_),
    .X(_09665_));
 sg13g2_nand2_1 _18761_ (.Y(_09666_),
    .A(_09663_),
    .B(_09665_));
 sg13g2_nand2_1 _18762_ (.Y(_09667_),
    .A(_09666_),
    .B(_09657_));
 sg13g2_nand2_1 _18763_ (.Y(_09668_),
    .A(_09647_),
    .B(_09648_));
 sg13g2_inv_1 _18764_ (.Y(_09669_),
    .A(_09668_));
 sg13g2_nand3_1 _18765_ (.B(_09665_),
    .C(_09669_),
    .A(_09663_),
    .Y(_09670_));
 sg13g2_buf_1 _18766_ (.A(_09670_),
    .X(_09671_));
 sg13g2_a21oi_2 _18767_ (.B1(_05718_),
    .Y(_09672_),
    .A2(net53),
    .A1(_06300_));
 sg13g2_o21ai_1 _18768_ (.B1(_09355_),
    .Y(_09673_),
    .A1(_04816_),
    .A2(_09672_));
 sg13g2_a21oi_1 _18769_ (.A1(_06306_),
    .A2(net53),
    .Y(_09674_),
    .B1(_06880_));
 sg13g2_inv_1 _18770_ (.Y(_09675_),
    .A(_09674_));
 sg13g2_a21oi_1 _18771_ (.A1(_09675_),
    .A2(net29),
    .Y(_09676_),
    .B1(_08169_));
 sg13g2_a21oi_1 _18772_ (.A1(_04480_),
    .A2(_04116_),
    .Y(_09677_),
    .B1(_04120_));
 sg13g2_inv_1 _18773_ (.Y(_09678_),
    .A(_09677_));
 sg13g2_a21oi_1 _18774_ (.A1(_09678_),
    .A2(_06185_),
    .Y(_09679_),
    .B1(_06189_));
 sg13g2_inv_1 _18775_ (.Y(_09680_),
    .A(_05956_));
 sg13g2_o21ai_1 _18776_ (.B1(_09680_),
    .Y(_09681_),
    .A1(_05864_),
    .A2(_09679_));
 sg13g2_a21oi_2 _18777_ (.B1(_06868_),
    .Y(_09682_),
    .A2(_04116_),
    .A1(_05003_));
 sg13g2_inv_1 _18778_ (.Y(_09683_),
    .A(_09682_));
 sg13g2_a21oi_1 _18779_ (.A1(_09683_),
    .A2(_06185_),
    .Y(_09684_),
    .B1(_06229_));
 sg13g2_inv_1 _18780_ (.Y(_09685_),
    .A(_09684_));
 sg13g2_a21oi_1 _18781_ (.A1(_09685_),
    .A2(_05863_),
    .Y(_09686_),
    .B1(_09080_));
 sg13g2_or2_1 _18782_ (.X(_09687_),
    .B(_09091_),
    .A(_09385_));
 sg13g2_a221oi_1 _18783_ (.B2(_09686_),
    .C1(_09687_),
    .B1(_09681_),
    .A1(_09673_),
    .Y(_09688_),
    .A2(_09676_));
 sg13g2_nor2b_1 _18784_ (.A(_09673_),
    .B_N(_09676_),
    .Y(_09689_));
 sg13g2_nor2b_1 _18785_ (.A(_09681_),
    .B_N(_09686_),
    .Y(_09690_));
 sg13g2_nor4_1 _18786_ (.A(_09689_),
    .B(_09414_),
    .C(_09083_),
    .D(_09690_),
    .Y(_09691_));
 sg13g2_a21oi_1 _18787_ (.A1(_09688_),
    .A2(_09691_),
    .Y(_09692_),
    .B1(_06556_));
 sg13g2_inv_1 _18788_ (.Y(_09693_),
    .A(_08903_));
 sg13g2_nor2_1 _18789_ (.A(_06551_),
    .B(_06805_),
    .Y(_09694_));
 sg13g2_a21oi_2 _18790_ (.B1(_07777_),
    .Y(_09695_),
    .A2(_05378_),
    .A1(_08438_));
 sg13g2_o21ai_1 _18791_ (.B1(_06595_),
    .Y(_09696_),
    .A1(_09368_),
    .A2(_09695_));
 sg13g2_buf_1 _18792_ (.A(_09696_),
    .X(_09697_));
 sg13g2_a21oi_1 _18793_ (.A1(_09697_),
    .A2(net26),
    .Y(_09698_),
    .B1(_06589_));
 sg13g2_inv_1 _18794_ (.Y(_09699_),
    .A(_09698_));
 sg13g2_inv_2 _18795_ (.Y(_09700_),
    .A(_08434_));
 sg13g2_a21oi_1 _18796_ (.A1(_09700_),
    .A2(_05377_),
    .Y(_09701_),
    .B1(_05537_));
 sg13g2_inv_1 _18797_ (.Y(_09702_),
    .A(_09701_));
 sg13g2_a21oi_1 _18798_ (.A1(_09702_),
    .A2(_04897_),
    .Y(_09703_),
    .B1(_04967_));
 sg13g2_inv_2 _18799_ (.Y(_09704_),
    .A(_09703_));
 sg13g2_a21oi_1 _18800_ (.A1(_09704_),
    .A2(net35),
    .Y(_09705_),
    .B1(_06812_));
 sg13g2_inv_2 _18801_ (.Y(_09706_),
    .A(_09705_));
 sg13g2_inv_1 _18802_ (.Y(_09707_),
    .A(_09248_));
 sg13g2_nand2_1 _18803_ (.Y(_09708_),
    .A(_09707_),
    .B(_09294_));
 sg13g2_o21ai_1 _18804_ (.B1(_09708_),
    .Y(_09709_),
    .A1(_09699_),
    .A2(_09706_));
 sg13g2_nor3_1 _18805_ (.A(_09693_),
    .B(_09694_),
    .C(_09709_),
    .Y(_09710_));
 sg13g2_a22oi_1 _18806_ (.Y(_09711_),
    .B1(_09707_),
    .B2(_09236_),
    .A2(_06550_),
    .A1(_06805_));
 sg13g2_o21ai_1 _18807_ (.B1(_09711_),
    .Y(_09712_),
    .A1(_09699_),
    .A2(_09705_));
 sg13g2_inv_1 _18808_ (.Y(_09713_),
    .A(_09712_));
 sg13g2_a21oi_1 _18809_ (.A1(_09710_),
    .A2(_09713_),
    .Y(_09714_),
    .B1(_06556_));
 sg13g2_o21ai_1 _18810_ (.B1(_06554_),
    .Y(_09715_),
    .A1(_09692_),
    .A2(_09714_));
 sg13g2_a21oi_1 _18811_ (.A1(_09692_),
    .A2(_08162_),
    .Y(_09716_),
    .B1(_06523_));
 sg13g2_nand2_1 _18812_ (.Y(_09717_),
    .A(_09715_),
    .B(_09716_));
 sg13g2_nor4_1 _18813_ (.A(_09113_),
    .B(_09431_),
    .C(_09118_),
    .D(_09611_),
    .Y(_09718_));
 sg13g2_nor2_1 _18814_ (.A(_09378_),
    .B(_09428_),
    .Y(_09719_));
 sg13g2_nor2_1 _18815_ (.A(_09547_),
    .B(_06813_),
    .Y(_09720_));
 sg13g2_buf_2 _18816_ (.A(_09720_),
    .X(_09721_));
 sg13g2_nor3_1 _18817_ (.A(_09106_),
    .B(_09719_),
    .C(_09721_),
    .Y(_09722_));
 sg13g2_nand4_1 _18818_ (.B(_09132_),
    .C(_09383_),
    .A(_09157_),
    .Y(_09723_),
    .D(_09536_));
 sg13g2_nor2_1 _18819_ (.A(_09099_),
    .B(_09294_),
    .Y(_09724_));
 sg13g2_nor3_1 _18820_ (.A(_09372_),
    .B(_09723_),
    .C(_09724_),
    .Y(_09725_));
 sg13g2_nand4_1 _18821_ (.B(_06523_),
    .C(_09722_),
    .A(_09718_),
    .Y(_09726_),
    .D(_09725_));
 sg13g2_nor2_1 _18822_ (.A(net137),
    .B(_06524_),
    .Y(_09727_));
 sg13g2_nand3_1 _18823_ (.B(_09726_),
    .C(_09727_),
    .A(_09717_),
    .Y(_09728_));
 sg13g2_nor2_1 _18824_ (.A(_08903_),
    .B(_08912_),
    .Y(_09729_));
 sg13g2_nor4_1 _18825_ (.A(_05591_),
    .B(_05592_),
    .C(_05607_),
    .D(_05603_),
    .Y(_09730_));
 sg13g2_a21o_1 _18826_ (.A2(_09730_),
    .A1(net115),
    .B1(_05611_),
    .X(_09731_));
 sg13g2_nand2_1 _18827_ (.Y(_09732_),
    .A(_09731_),
    .B(_00014_));
 sg13g2_inv_1 _18828_ (.Y(_09733_),
    .A(_09732_));
 sg13g2_nand4_1 _18829_ (.B(_07073_),
    .C(_07086_),
    .A(_07081_),
    .Y(_09734_),
    .D(_07074_));
 sg13g2_inv_1 _18830_ (.Y(_09735_),
    .A(_09734_));
 sg13g2_a21oi_2 _18831_ (.B1(_07091_),
    .Y(_09736_),
    .A2(_09735_),
    .A1(net88));
 sg13g2_nor2_2 _18832_ (.A(_07135_),
    .B(_09736_),
    .Y(_09737_));
 sg13g2_nor3_1 _18833_ (.A(_09733_),
    .B(_09737_),
    .C(_08674_),
    .Y(_09738_));
 sg13g2_inv_1 _18834_ (.Y(_09739_),
    .A(_09384_));
 sg13g2_nor2_1 _18835_ (.A(_09537_),
    .B(_09131_),
    .Y(_09740_));
 sg13g2_nand4_1 _18836_ (.B(_08176_),
    .C(_09739_),
    .A(_09738_),
    .Y(_09741_),
    .D(_09740_));
 sg13g2_nor4_1 _18837_ (.A(_09544_),
    .B(_09724_),
    .C(_09729_),
    .D(_09741_),
    .Y(_09742_));
 sg13g2_and4_1 _18838_ (.A(_09713_),
    .B(_09688_),
    .C(_09722_),
    .D(_09742_),
    .X(_09743_));
 sg13g2_nand2_1 _18839_ (.Y(_09744_),
    .A(_08912_),
    .B(_09693_));
 sg13g2_nor2_2 _18840_ (.A(_03959_),
    .B(_09736_),
    .Y(_09745_));
 sg13g2_nand2_1 _18841_ (.Y(_09746_),
    .A(_09731_),
    .B(_03557_));
 sg13g2_inv_1 _18842_ (.Y(_09747_),
    .A(_09746_));
 sg13g2_nor2_1 _18843_ (.A(_09745_),
    .B(_09747_),
    .Y(_09748_));
 sg13g2_inv_1 _18844_ (.Y(_09749_),
    .A(_09748_));
 sg13g2_nor3_1 _18845_ (.A(_08040_),
    .B(_07902_),
    .C(_08179_),
    .Y(_09750_));
 sg13g2_nor2_1 _18846_ (.A(_09609_),
    .B(_09156_),
    .Y(_09751_));
 sg13g2_nand2_1 _18847_ (.Y(_09752_),
    .A(_09750_),
    .B(_09751_));
 sg13g2_nor4_1 _18848_ (.A(_09694_),
    .B(_09749_),
    .C(_09409_),
    .D(_09752_),
    .Y(_09753_));
 sg13g2_nand4_1 _18849_ (.B(_09486_),
    .C(_09744_),
    .A(_09691_),
    .Y(_09754_),
    .D(_09753_));
 sg13g2_nand2b_1 _18850_ (.Y(_09755_),
    .B(_09718_),
    .A_N(_09709_));
 sg13g2_nor2_1 _18851_ (.A(_09754_),
    .B(_09755_),
    .Y(_09756_));
 sg13g2_nand2_1 _18852_ (.Y(_09757_),
    .A(_09743_),
    .B(_09756_));
 sg13g2_o21ai_1 _18853_ (.B1(_06519_),
    .Y(_09758_),
    .A1(_06516_),
    .A2(_06521_));
 sg13g2_nand3_1 _18854_ (.B(net161),
    .C(_09758_),
    .A(_09757_),
    .Y(_09759_));
 sg13g2_nor3_1 _18855_ (.A(_06521_),
    .B(_09756_),
    .C(_09743_),
    .Y(_09760_));
 sg13g2_nand3_1 _18856_ (.B(net191),
    .C(_06522_),
    .A(_09760_),
    .Y(_09761_));
 sg13g2_nand3_1 _18857_ (.B(_09759_),
    .C(_09761_),
    .A(_09728_),
    .Y(_09762_));
 sg13g2_buf_2 _18858_ (.A(\b.gen_square[11].sq.mask ),
    .X(_09763_));
 sg13g2_nand2_1 _18859_ (.Y(_09764_),
    .A(_09762_),
    .B(_09763_));
 sg13g2_nand3_1 _18860_ (.B(_09671_),
    .C(_09764_),
    .A(_09667_),
    .Y(_09765_));
 sg13g2_nand2_1 _18861_ (.Y(_09766_),
    .A(_09642_),
    .B(_09632_));
 sg13g2_nand2_1 _18862_ (.Y(_09767_),
    .A(_09766_),
    .B(_09644_));
 sg13g2_nor3_1 _18863_ (.A(_06513_),
    .B(_06515_),
    .C(_06522_),
    .Y(_09768_));
 sg13g2_nand2_1 _18864_ (.Y(_09769_),
    .A(_06521_),
    .B(_09768_));
 sg13g2_inv_1 _18865_ (.Y(_09770_),
    .A(_09769_));
 sg13g2_nand4_1 _18866_ (.B(_09750_),
    .C(_08176_),
    .A(_09738_),
    .Y(_09771_),
    .D(_09748_));
 sg13g2_nand2_1 _18867_ (.Y(_09772_),
    .A(_09714_),
    .B(_06555_));
 sg13g2_nand2_1 _18868_ (.Y(_09773_),
    .A(_09715_),
    .B(_09772_));
 sg13g2_a221oi_1 _18869_ (.B2(_09771_),
    .C1(_09773_),
    .B1(_09770_),
    .A1(_08162_),
    .Y(_09774_),
    .A2(_09692_));
 sg13g2_nor2_1 _18870_ (.A(_06513_),
    .B(_06552_),
    .Y(_09775_));
 sg13g2_nand2_1 _18871_ (.Y(_09776_),
    .A(_09760_),
    .B(net215));
 sg13g2_nand3_1 _18872_ (.B(net176),
    .C(_06556_),
    .A(_09757_),
    .Y(_09777_));
 sg13g2_nand2_1 _18873_ (.Y(_09778_),
    .A(_09776_),
    .B(_09777_));
 sg13g2_o21ai_1 _18874_ (.B1(_09778_),
    .Y(_09779_),
    .A1(_06554_),
    .A2(_09775_));
 sg13g2_o21ai_1 _18875_ (.B1(_09779_),
    .Y(_09780_),
    .A1(net154),
    .A2(_09774_));
 sg13g2_nand2_1 _18876_ (.Y(_09781_),
    .A(_09780_),
    .B(_09763_));
 sg13g2_nor2_1 _18877_ (.A(_09767_),
    .B(_09781_),
    .Y(_09782_));
 sg13g2_nand2_1 _18878_ (.Y(_09783_),
    .A(_09781_),
    .B(_09767_));
 sg13g2_nor2b_1 _18879_ (.A(_09782_),
    .B_N(_09783_),
    .Y(_09784_));
 sg13g2_nand2_1 _18880_ (.Y(_09785_),
    .A(_09765_),
    .B(_09784_));
 sg13g2_nand2_1 _18881_ (.Y(_09786_),
    .A(_09666_),
    .B(_09660_));
 sg13g2_nand3_1 _18882_ (.B(_09531_),
    .C(_09665_),
    .A(_09663_),
    .Y(_09787_));
 sg13g2_nand2_1 _18883_ (.Y(_09788_),
    .A(_09786_),
    .B(_09787_));
 sg13g2_a22oi_1 _18884_ (.Y(_09789_),
    .B1(_06518_),
    .B2(_09776_),
    .A2(_06553_),
    .A1(_06517_));
 sg13g2_a21oi_1 _18885_ (.A1(_09715_),
    .A2(_09772_),
    .Y(_09790_),
    .B1(net154));
 sg13g2_a21o_1 _18886_ (.A2(_09778_),
    .A1(_09789_),
    .B1(_09790_),
    .X(_09791_));
 sg13g2_nand2_1 _18887_ (.Y(_09792_),
    .A(_09791_),
    .B(_09763_));
 sg13g2_nand2_1 _18888_ (.Y(_09793_),
    .A(_09788_),
    .B(_09792_));
 sg13g2_inv_1 _18889_ (.Y(_09794_),
    .A(_09792_));
 sg13g2_nand3_1 _18890_ (.B(_09787_),
    .C(_09794_),
    .A(_09786_),
    .Y(_09795_));
 sg13g2_nand2_1 _18891_ (.Y(_09796_),
    .A(_09793_),
    .B(_09795_));
 sg13g2_nor2_1 _18892_ (.A(_09785_),
    .B(_09796_),
    .Y(_09797_));
 sg13g2_a21oi_1 _18893_ (.A1(_09667_),
    .A2(_09671_),
    .Y(_09798_),
    .B1(_09764_));
 sg13g2_nand2_1 _18894_ (.Y(_09799_),
    .A(_09797_),
    .B(_09798_));
 sg13g2_nand2_1 _18895_ (.Y(_09800_),
    .A(_09667_),
    .B(_09671_));
 sg13g2_inv_2 _18896_ (.Y(_09801_),
    .A(_09795_));
 sg13g2_a21oi_2 _18897_ (.B1(_09782_),
    .Y(_09802_),
    .A2(_09784_),
    .A1(_09801_));
 sg13g2_nand3_1 _18898_ (.B(_09800_),
    .C(_09802_),
    .A(_09799_),
    .Y(_09803_));
 sg13g2_nand2b_1 _18899_ (.Y(_09804_),
    .B(_09764_),
    .A_N(_09802_));
 sg13g2_nand2_1 _18900_ (.Y(_09805_),
    .A(_09803_),
    .B(_09804_));
 sg13g2_nand2_1 _18901_ (.Y(_09806_),
    .A(_09799_),
    .B(_09802_));
 sg13g2_nand2_1 _18902_ (.Y(_09807_),
    .A(_09806_),
    .B(_09792_));
 sg13g2_inv_1 _18903_ (.Y(_09808_),
    .A(_09788_));
 sg13g2_nand3_1 _18904_ (.B(_09808_),
    .C(_09802_),
    .A(_09799_),
    .Y(_09809_));
 sg13g2_nand2_1 _18905_ (.Y(_09810_),
    .A(_09807_),
    .B(_09809_));
 sg13g2_a21oi_1 _18906_ (.A1(_07948_),
    .A2(_04928_),
    .Y(_09811_),
    .B1(_04972_));
 sg13g2_inv_1 _18907_ (.Y(_09812_),
    .A(_09811_));
 sg13g2_a21oi_1 _18908_ (.A1(_09812_),
    .A2(net55),
    .Y(_09813_),
    .B1(_05532_));
 sg13g2_inv_1 _18909_ (.Y(_09814_),
    .A(_09813_));
 sg13g2_a21oi_1 _18910_ (.A1(_09814_),
    .A2(net22),
    .Y(_09815_),
    .B1(_05956_));
 sg13g2_o21ai_1 _18911_ (.B1(_06984_),
    .Y(_09816_),
    .A1(_06203_),
    .A2(_07951_));
 sg13g2_a21oi_1 _18912_ (.A1(_09816_),
    .A2(net40),
    .Y(_09817_),
    .B1(_06979_));
 sg13g2_inv_1 _18913_ (.Y(_09818_),
    .A(_09817_));
 sg13g2_a21oi_1 _18914_ (.A1(_09818_),
    .A2(net22),
    .Y(_09819_),
    .B1(_06971_));
 sg13g2_inv_1 _18915_ (.Y(_09820_),
    .A(_09246_));
 sg13g2_nand2_1 _18916_ (.Y(_09821_),
    .A(_09290_),
    .B(_09292_));
 sg13g2_inv_1 _18917_ (.Y(_09822_),
    .A(_09821_));
 sg13g2_a22oi_1 _18918_ (.Y(_09823_),
    .B1(_09820_),
    .B2(_09822_),
    .A2(_06935_),
    .A1(_06998_));
 sg13g2_o21ai_1 _18919_ (.B1(_09823_),
    .Y(_09824_),
    .A1(_08905_),
    .A2(_08914_));
 sg13g2_a21oi_1 _18920_ (.A1(_09815_),
    .A2(_09819_),
    .Y(_09825_),
    .B1(_09824_));
 sg13g2_nor4_1 _18921_ (.A(_08934_),
    .B(_09608_),
    .C(_09115_),
    .D(_09118_),
    .Y(_09826_));
 sg13g2_a21oi_1 _18922_ (.A1(_05252_),
    .A2(_05678_),
    .Y(_09827_),
    .B1(_06755_));
 sg13g2_o21ai_1 _18923_ (.B1(_07202_),
    .Y(_09828_),
    .A1(_08277_),
    .A2(_09827_));
 sg13g2_a21oi_1 _18924_ (.A1(_09828_),
    .A2(net26),
    .Y(_09829_),
    .B1(_07590_));
 sg13g2_inv_1 _18925_ (.Y(_09830_),
    .A(_09829_));
 sg13g2_a21oi_1 _18926_ (.A1(_08064_),
    .A2(net26),
    .Y(_09831_),
    .B1(_06812_));
 sg13g2_nor2b_1 _18927_ (.A(_09830_),
    .B_N(_09831_),
    .Y(_09832_));
 sg13g2_nand2_1 _18928_ (.Y(_09833_),
    .A(_09612_),
    .B(_09155_));
 sg13g2_a21oi_1 _18929_ (.A1(_04985_),
    .A2(_04153_),
    .Y(_09834_),
    .B1(_04224_));
 sg13g2_inv_1 _18930_ (.Y(_09835_),
    .A(_09834_));
 sg13g2_a21oi_1 _18931_ (.A1(_09835_),
    .A2(_05289_),
    .Y(_09836_),
    .B1(_05527_));
 sg13g2_a21oi_1 _18932_ (.A1(_07225_),
    .A2(_04153_),
    .Y(_09837_),
    .B1(_06688_));
 sg13g2_inv_1 _18933_ (.Y(_09838_),
    .A(_09837_));
 sg13g2_a21oi_1 _18934_ (.A1(_09838_),
    .A2(_05289_),
    .Y(_09839_),
    .B1(_08799_));
 sg13g2_a221oi_1 _18935_ (.B2(_09839_),
    .C1(_09601_),
    .B1(_09836_),
    .A1(_09014_),
    .Y(_09840_),
    .A2(_08280_));
 sg13g2_inv_1 _18936_ (.Y(_09841_),
    .A(_04159_));
 sg13g2_nor3_1 _18937_ (.A(_04156_),
    .B(_04158_),
    .C(_09841_),
    .Y(_09842_));
 sg13g2_nand2_1 _18938_ (.Y(_09843_),
    .A(_04167_),
    .B(_09842_));
 sg13g2_inv_1 _18939_ (.Y(_09844_),
    .A(_09843_));
 sg13g2_a21oi_1 _18940_ (.A1(net88),
    .A2(_09844_),
    .Y(_09845_),
    .B1(_04171_));
 sg13g2_nor2_1 _18941_ (.A(_04002_),
    .B(_09845_),
    .Y(_09846_));
 sg13g2_nor2_1 _18942_ (.A(_09846_),
    .B(_08422_),
    .Y(_09847_));
 sg13g2_inv_1 _18943_ (.Y(_09848_),
    .A(_09847_));
 sg13g2_nor4_1 _18944_ (.A(_07835_),
    .B(_07837_),
    .C(_09848_),
    .D(_09283_),
    .Y(_09849_));
 sg13g2_nand3_1 _18945_ (.B(_09849_),
    .C(_09751_),
    .A(_09840_),
    .Y(_09850_));
 sg13g2_nor3_1 _18946_ (.A(_09832_),
    .B(_09833_),
    .C(_09850_),
    .Y(_09851_));
 sg13g2_nand3_1 _18947_ (.B(_09826_),
    .C(_09851_),
    .A(_09825_),
    .Y(_09852_));
 sg13g2_inv_1 _18948_ (.Y(_09853_),
    .A(_09815_));
 sg13g2_nand2_1 _18949_ (.Y(_09854_),
    .A(_08914_),
    .B(_08904_));
 sg13g2_o21ai_1 _18950_ (.B1(_09854_),
    .Y(_09855_),
    .A1(_06998_),
    .A2(_06936_));
 sg13g2_a221oi_1 _18951_ (.B2(_09819_),
    .C1(_09855_),
    .B1(_09853_),
    .A1(_09234_),
    .Y(_09856_),
    .A2(_09820_));
 sg13g2_inv_1 _18952_ (.Y(_09857_),
    .A(_08933_));
 sg13g2_a21oi_1 _18953_ (.A1(_09857_),
    .A2(_09821_),
    .Y(_09858_),
    .B1(_09106_));
 sg13g2_nor2_2 _18954_ (.A(_09541_),
    .B(_06809_),
    .Y(_09859_));
 sg13g2_nor4_1 _18955_ (.A(_09859_),
    .B(_09015_),
    .C(_09103_),
    .D(_09721_),
    .Y(_09860_));
 sg13g2_inv_1 _18956_ (.Y(_09861_),
    .A(_09839_));
 sg13g2_nor2_1 _18957_ (.A(_09560_),
    .B(_09016_),
    .Y(_09862_));
 sg13g2_o21ai_1 _18958_ (.B1(_09862_),
    .Y(_09863_),
    .A1(_09836_),
    .A2(_09861_));
 sg13g2_nor2_1 _18959_ (.A(_07747_),
    .B(_08265_),
    .Y(_09864_));
 sg13g2_nor2b_1 _18960_ (.A(_09845_),
    .B_N(_00077_),
    .Y(_09865_));
 sg13g2_nor2_1 _18961_ (.A(_09865_),
    .B(_08413_),
    .Y(_09866_));
 sg13g2_nand4_1 _18962_ (.B(_09864_),
    .C(_09866_),
    .A(_07759_),
    .Y(_09867_),
    .D(_09215_));
 sg13g2_inv_1 _18963_ (.Y(_09868_),
    .A(_09867_));
 sg13g2_nand2_1 _18964_ (.Y(_09869_),
    .A(_09868_),
    .B(_09740_));
 sg13g2_nor2_1 _18965_ (.A(_09830_),
    .B(_09831_),
    .Y(_09870_));
 sg13g2_nor3_1 _18966_ (.A(_09863_),
    .B(_09869_),
    .C(_09870_),
    .Y(_09871_));
 sg13g2_nand4_1 _18967_ (.B(_09858_),
    .C(_09860_),
    .A(_09856_),
    .Y(_09872_),
    .D(_09871_));
 sg13g2_nor2_1 _18968_ (.A(_09852_),
    .B(_09872_),
    .Y(_09873_));
 sg13g2_inv_1 _18969_ (.Y(_09874_),
    .A(_09873_));
 sg13g2_nand3_1 _18970_ (.B(net161),
    .C(_06956_),
    .A(_09874_),
    .Y(_09875_));
 sg13g2_nand4_1 _18971_ (.B(net191),
    .C(_06956_),
    .A(_09872_),
    .Y(_09876_),
    .D(_09852_));
 sg13g2_buf_1 _18972_ (.A(_09876_),
    .X(_09877_));
 sg13g2_nand2_1 _18973_ (.Y(_09878_),
    .A(_09875_),
    .B(_09877_));
 sg13g2_nand2_1 _18974_ (.Y(_09879_),
    .A(_09877_),
    .B(_06942_));
 sg13g2_nand2b_1 _18975_ (.Y(_09880_),
    .B(_06941_),
    .A_N(_06959_));
 sg13g2_nand3_1 _18976_ (.B(_09879_),
    .C(_09880_),
    .A(_09878_),
    .Y(_09881_));
 sg13g2_a21o_1 _18977_ (.A2(_09825_),
    .A1(_09856_),
    .B1(_06956_),
    .X(_09882_));
 sg13g2_nand3b_1 _18978_ (.B(_09840_),
    .C(_09830_),
    .Y(_09883_),
    .A_N(_09863_));
 sg13g2_nand2_1 _18979_ (.Y(_09884_),
    .A(_09883_),
    .B(_06945_));
 sg13g2_a21o_1 _18980_ (.A2(_09884_),
    .A1(_09882_),
    .B1(_06960_),
    .X(_09885_));
 sg13g2_nand2b_1 _18981_ (.Y(_09886_),
    .B(_06958_),
    .A_N(_09882_));
 sg13g2_nand2_1 _18982_ (.Y(_09887_),
    .A(_09885_),
    .B(_09886_));
 sg13g2_nand2_1 _18983_ (.Y(_09888_),
    .A(_09887_),
    .B(net160));
 sg13g2_nand2_1 _18984_ (.Y(_09889_),
    .A(_09881_),
    .B(_09888_));
 sg13g2_buf_1 _18985_ (.A(\b.gen_square[12].sq.mask ),
    .X(_09890_));
 sg13g2_nand2_1 _18986_ (.Y(_09891_),
    .A(_09889_),
    .B(_09890_));
 sg13g2_inv_1 _18987_ (.Y(_09892_),
    .A(_09891_));
 sg13g2_nor2_1 _18988_ (.A(_02045_),
    .B(_06947_),
    .Y(_09893_));
 sg13g2_nand3_1 _18989_ (.B(_06945_),
    .C(_08282_),
    .A(_09883_),
    .Y(_09894_));
 sg13g2_nor3_1 _18990_ (.A(_06937_),
    .B(_06939_),
    .C(_06946_),
    .Y(_09895_));
 sg13g2_nand2_1 _18991_ (.Y(_09896_),
    .A(_06945_),
    .B(_09895_));
 sg13g2_a21o_1 _18992_ (.A2(_09868_),
    .A1(_09849_),
    .B1(_09896_),
    .X(_09897_));
 sg13g2_nand2_1 _18993_ (.Y(_09898_),
    .A(_09894_),
    .B(_09897_));
 sg13g2_xnor2_1 _18994_ (.Y(_09899_),
    .A(_06937_),
    .B(_06959_));
 sg13g2_a22oi_1 _18995_ (.Y(_09900_),
    .B1(_09899_),
    .B2(_09878_),
    .A2(_09898_),
    .A1(_09893_));
 sg13g2_nand2_1 _18996_ (.Y(_09901_),
    .A(_09900_),
    .B(_09888_));
 sg13g2_nand2_1 _18997_ (.Y(_09902_),
    .A(_09901_),
    .B(_09890_));
 sg13g2_a21oi_1 _18998_ (.A1(_09780_),
    .A2(_09763_),
    .Y(_09903_),
    .B1(_09767_));
 sg13g2_inv_1 _18999_ (.Y(_09904_),
    .A(_09903_));
 sg13g2_nor2_1 _19000_ (.A(_09902_),
    .B(_09904_),
    .Y(_09905_));
 sg13g2_a21oi_1 _19001_ (.A1(_09810_),
    .A2(_09892_),
    .Y(_09906_),
    .B1(_09905_));
 sg13g2_nand3_1 _19002_ (.B(_06948_),
    .C(_09894_),
    .A(_09885_),
    .Y(_09907_));
 sg13g2_inv_1 _19003_ (.Y(_09908_),
    .A(_09536_));
 sg13g2_nor4_1 _19004_ (.A(_06948_),
    .B(_09121_),
    .C(_09908_),
    .D(_09833_),
    .Y(_09909_));
 sg13g2_nand4_1 _19005_ (.B(_09858_),
    .C(_09860_),
    .A(_09909_),
    .Y(_09910_),
    .D(_09826_));
 sg13g2_nor2_1 _19006_ (.A(net120),
    .B(_06949_),
    .Y(_09911_));
 sg13g2_nand3_1 _19007_ (.B(_09910_),
    .C(_09911_),
    .A(_09907_),
    .Y(_09912_));
 sg13g2_o21ai_1 _19008_ (.B1(_06943_),
    .Y(_09913_),
    .A1(_06940_),
    .A2(_06945_));
 sg13g2_nand3_1 _19009_ (.B(net144),
    .C(_09913_),
    .A(_09874_),
    .Y(_09914_));
 sg13g2_nand2b_1 _19010_ (.Y(_09915_),
    .B(_06946_),
    .A_N(_09877_));
 sg13g2_nand3_1 _19011_ (.B(_09914_),
    .C(_09915_),
    .A(_09912_),
    .Y(_09916_));
 sg13g2_nand2_1 _19012_ (.Y(_09917_),
    .A(_09916_),
    .B(_09890_));
 sg13g2_a21oi_1 _19013_ (.A1(_09803_),
    .A2(_09804_),
    .Y(_09918_),
    .B1(_09917_));
 sg13g2_nand3_1 _19014_ (.B(_09809_),
    .C(_09891_),
    .A(_09807_),
    .Y(_09919_));
 sg13g2_nand2_1 _19015_ (.Y(_09920_),
    .A(_09918_),
    .B(_09919_));
 sg13g2_nand2_1 _19016_ (.Y(_09921_),
    .A(_09906_),
    .B(_09920_));
 sg13g2_nand2_1 _19017_ (.Y(_09922_),
    .A(_09904_),
    .B(_09902_));
 sg13g2_nand2_1 _19018_ (.Y(_09923_),
    .A(_09921_),
    .B(_09922_));
 sg13g2_nand2b_1 _19019_ (.Y(_09924_),
    .B(_09923_),
    .A_N(_09805_));
 sg13g2_nand3b_1 _19020_ (.B(_09921_),
    .C(_09922_),
    .Y(_09925_),
    .A_N(_09917_));
 sg13g2_nand2_1 _19021_ (.Y(_09926_),
    .A(_09924_),
    .B(_09925_));
 sg13g2_nor2_1 _19022_ (.A(_09170_),
    .B(_09926_),
    .Y(_09927_));
 sg13g2_nand2_1 _19023_ (.Y(_09928_),
    .A(_09923_),
    .B(_09810_));
 sg13g2_nand3_1 _19024_ (.B(_09922_),
    .C(_09891_),
    .A(_09921_),
    .Y(_09929_));
 sg13g2_nand3_1 _19025_ (.B(net129),
    .C(_05891_),
    .A(_09162_),
    .Y(_09930_));
 sg13g2_nand2_1 _19026_ (.Y(_09931_),
    .A(_09930_),
    .B(_09166_));
 sg13g2_nand2_1 _19027_ (.Y(_09932_),
    .A(_09166_),
    .B(_05878_));
 sg13g2_nand2b_1 _19028_ (.Y(_09933_),
    .B(_05877_),
    .A_N(_05894_));
 sg13g2_nand3_1 _19029_ (.B(_09932_),
    .C(_09933_),
    .A(_09931_),
    .Y(_09934_));
 sg13g2_nor3_1 _19030_ (.A(_05873_),
    .B(_05877_),
    .C(_09076_),
    .Y(_09935_));
 sg13g2_nand2b_1 _19031_ (.Y(_09936_),
    .B(_09096_),
    .A_N(_09935_));
 sg13g2_nand3_1 _19032_ (.B(net128),
    .C(_05882_),
    .A(_09936_),
    .Y(_09937_));
 sg13g2_nand2_1 _19033_ (.Y(_09938_),
    .A(_09934_),
    .B(_09937_));
 sg13g2_nand2_1 _19034_ (.Y(_09939_),
    .A(_09938_),
    .B(_09169_));
 sg13g2_nand3_1 _19035_ (.B(_09929_),
    .C(_09939_),
    .A(_09928_),
    .Y(_09940_));
 sg13g2_nand2_1 _19036_ (.Y(_09941_),
    .A(_09927_),
    .B(_09940_));
 sg13g2_nand2_1 _19037_ (.Y(_09942_),
    .A(_09928_),
    .B(_09929_));
 sg13g2_inv_1 _19038_ (.Y(_09943_),
    .A(_09939_));
 sg13g2_xnor2_1 _19039_ (.Y(_09944_),
    .A(_05873_),
    .B(_05894_));
 sg13g2_nand2_1 _19040_ (.Y(_09945_),
    .A(_09931_),
    .B(_09944_));
 sg13g2_inv_1 _19041_ (.Y(_09946_),
    .A(_09152_));
 sg13g2_nor2_1 _19042_ (.A(_09148_),
    .B(_07919_),
    .Y(_09947_));
 sg13g2_nand3_1 _19043_ (.B(_09947_),
    .C(_09139_),
    .A(_09946_),
    .Y(_09948_));
 sg13g2_nand4_1 _19044_ (.B(_05874_),
    .C(_05880_),
    .A(_05884_),
    .Y(_09949_),
    .D(_05876_));
 sg13g2_inv_1 _19045_ (.Y(_09950_),
    .A(_09949_));
 sg13g2_o21ai_1 _19046_ (.B1(_09950_),
    .Y(_09951_),
    .A1(_09130_),
    .A2(_09948_));
 sg13g2_nand2_1 _19047_ (.Y(_09952_),
    .A(_09097_),
    .B(_09951_));
 sg13g2_nand3_1 _19048_ (.B(net128),
    .C(_05882_),
    .A(_09952_),
    .Y(_09953_));
 sg13g2_nand3_1 _19049_ (.B(_09945_),
    .C(_09953_),
    .A(_09937_),
    .Y(_09954_));
 sg13g2_nand2_1 _19050_ (.Y(_09955_),
    .A(_09954_),
    .B(_09169_));
 sg13g2_nand2_1 _19051_ (.Y(_09956_),
    .A(_09903_),
    .B(_09902_));
 sg13g2_nor2_1 _19052_ (.A(_09955_),
    .B(_09956_),
    .Y(_09957_));
 sg13g2_a21oi_1 _19053_ (.A1(_09942_),
    .A2(_09943_),
    .Y(_09958_),
    .B1(_09957_));
 sg13g2_nand2_1 _19054_ (.Y(_09959_),
    .A(_09941_),
    .B(_09958_));
 sg13g2_nand2_1 _19055_ (.Y(_09960_),
    .A(_09956_),
    .B(_09955_));
 sg13g2_nand3b_1 _19056_ (.B(_09959_),
    .C(_09960_),
    .Y(_09961_),
    .A_N(_09170_));
 sg13g2_nand2_1 _19057_ (.Y(_09962_),
    .A(_09959_),
    .B(_09960_));
 sg13g2_nand2_1 _19058_ (.Y(_09963_),
    .A(_09962_),
    .B(_09926_));
 sg13g2_nand2_1 _19059_ (.Y(_09964_),
    .A(_09961_),
    .B(_09963_));
 sg13g2_nor2_1 _19060_ (.A(_09047_),
    .B(_09964_),
    .Y(_09965_));
 sg13g2_nand2_1 _19061_ (.Y(_09966_),
    .A(_09962_),
    .B(_09942_));
 sg13g2_nand3_1 _19062_ (.B(_09939_),
    .C(_09960_),
    .A(_09959_),
    .Y(_09967_));
 sg13g2_nand3_1 _19063_ (.B(net113),
    .C(_04272_),
    .A(_09027_),
    .Y(_09968_));
 sg13g2_nand2_1 _19064_ (.Y(_09969_),
    .A(_09026_),
    .B(_09968_));
 sg13g2_nand2_1 _19065_ (.Y(_09970_),
    .A(_09026_),
    .B(_04182_));
 sg13g2_nand2b_1 _19066_ (.Y(_09971_),
    .B(_04181_),
    .A_N(_04275_));
 sg13g2_nand3_1 _19067_ (.B(_09970_),
    .C(_09971_),
    .A(_09969_),
    .Y(_09972_));
 sg13g2_nand2b_1 _19068_ (.Y(_09973_),
    .B(_04274_),
    .A_N(_09035_));
 sg13g2_a21o_1 _19069_ (.A2(_09973_),
    .A1(_09036_),
    .B1(net103),
    .X(_09974_));
 sg13g2_nand2_1 _19070_ (.Y(_09975_),
    .A(_09972_),
    .B(_09974_));
 sg13g2_nand2_1 _19071_ (.Y(_09976_),
    .A(_09975_),
    .B(_09046_));
 sg13g2_nand3_1 _19072_ (.B(_09967_),
    .C(_09976_),
    .A(_09966_),
    .Y(_09977_));
 sg13g2_nand2_1 _19073_ (.Y(_09978_),
    .A(_09965_),
    .B(_09977_));
 sg13g2_nand2_1 _19074_ (.Y(_09979_),
    .A(_09966_),
    .B(_09967_));
 sg13g2_inv_1 _19075_ (.Y(_09980_),
    .A(_09976_));
 sg13g2_nand3_1 _19076_ (.B(_04185_),
    .C(_04180_),
    .A(_04178_),
    .Y(_09981_));
 sg13g2_nor2_1 _19077_ (.A(_09981_),
    .B(_04272_),
    .Y(_09982_));
 sg13g2_inv_1 _19078_ (.Y(_09983_),
    .A(_09982_));
 sg13g2_a21oi_1 _19079_ (.A1(_08975_),
    .A2(_09011_),
    .Y(_09984_),
    .B1(_09983_));
 sg13g2_nor2_1 _19080_ (.A(net103),
    .B(_09107_),
    .Y(_09985_));
 sg13g2_o21ai_1 _19081_ (.B1(_09985_),
    .Y(_09986_),
    .A1(_09984_),
    .A2(_09033_));
 sg13g2_xnor2_1 _19082_ (.Y(_09987_),
    .A(_04177_),
    .B(_04275_));
 sg13g2_nand2_1 _19083_ (.Y(_09988_),
    .A(_09969_),
    .B(_09987_));
 sg13g2_nand3_1 _19084_ (.B(_09986_),
    .C(_09988_),
    .A(_09974_),
    .Y(_09989_));
 sg13g2_nand2_1 _19085_ (.Y(_09990_),
    .A(_09989_),
    .B(_09046_));
 sg13g2_inv_1 _19086_ (.Y(_09991_),
    .A(_09990_));
 sg13g2_nor2b_1 _19087_ (.A(_09956_),
    .B_N(_09955_),
    .Y(_09992_));
 sg13g2_xnor2_1 _19088_ (.Y(_09993_),
    .A(_09991_),
    .B(_09992_));
 sg13g2_a21oi_1 _19089_ (.A1(_09979_),
    .A2(_09980_),
    .Y(_09994_),
    .B1(_09993_));
 sg13g2_nand2_1 _19090_ (.Y(_09995_),
    .A(_09978_),
    .B(_09994_));
 sg13g2_inv_1 _19091_ (.Y(_09996_),
    .A(_09992_));
 sg13g2_nand2_1 _19092_ (.Y(_09997_),
    .A(_09996_),
    .B(_09990_));
 sg13g2_nand3b_1 _19093_ (.B(_09995_),
    .C(_09997_),
    .Y(_09998_),
    .A_N(_09047_));
 sg13g2_nand2_2 _19094_ (.Y(_09999_),
    .A(_09995_),
    .B(_09997_));
 sg13g2_nand2_1 _19095_ (.Y(_10000_),
    .A(_09999_),
    .B(_09964_));
 sg13g2_nand2_1 _19096_ (.Y(_10001_),
    .A(_09998_),
    .B(_10000_));
 sg13g2_nor3_1 _19097_ (.A(_07896_),
    .B(_09745_),
    .C(_07902_),
    .Y(_10002_));
 sg13g2_nor3_1 _19098_ (.A(_08978_),
    .B(_09086_),
    .C(_08982_),
    .Y(_10003_));
 sg13g2_nand2_1 _19099_ (.Y(_10004_),
    .A(_10002_),
    .B(_10003_));
 sg13g2_a21oi_1 _19100_ (.A1(_08833_),
    .A2(_07499_),
    .Y(_10005_),
    .B1(_07541_));
 sg13g2_inv_1 _19101_ (.Y(_10006_),
    .A(_10005_));
 sg13g2_a21oi_1 _19102_ (.A1(_10006_),
    .A2(_07494_),
    .Y(_10007_),
    .B1(_07533_));
 sg13g2_inv_1 _19103_ (.Y(_10008_),
    .A(_10007_));
 sg13g2_a21oi_1 _19104_ (.A1(_10008_),
    .A2(_07491_),
    .Y(_10009_),
    .B1(_07523_));
 sg13g2_inv_1 _19105_ (.Y(_10010_),
    .A(_10009_));
 sg13g2_a21oi_2 _19106_ (.B1(_07500_),
    .Y(_10011_),
    .A2(_07499_),
    .A1(_07611_));
 sg13g2_inv_1 _19107_ (.Y(_10012_),
    .A(_10011_));
 sg13g2_a21oi_1 _19108_ (.A1(_10012_),
    .A2(_07494_),
    .Y(_10013_),
    .B1(_07496_));
 sg13g2_a21oi_1 _19109_ (.A1(_10013_),
    .A2(_07491_),
    .Y(_10014_),
    .B1(_07492_));
 sg13g2_a21oi_1 _19110_ (.A1(_10010_),
    .A2(_08944_),
    .Y(_10015_),
    .B1(_10014_));
 sg13g2_o21ai_1 _19111_ (.B1(_04937_),
    .Y(_10016_),
    .A1(_06203_),
    .A2(_07870_));
 sg13g2_buf_1 _19112_ (.A(_10016_),
    .X(_10017_));
 sg13g2_a21oi_1 _19113_ (.A1(_10017_),
    .A2(_06186_),
    .Y(_10018_),
    .B1(_06229_));
 sg13g2_inv_1 _19114_ (.Y(_10019_),
    .A(_10018_));
 sg13g2_a21oi_1 _19115_ (.A1(_10019_),
    .A2(net47),
    .Y(_10020_),
    .B1(_06217_));
 sg13g2_inv_1 _19116_ (.Y(_10021_),
    .A(_10020_));
 sg13g2_nand2_1 _19117_ (.Y(_10022_),
    .A(_10021_),
    .B(_08938_));
 sg13g2_a21oi_1 _19118_ (.A1(_06468_),
    .A2(net58),
    .Y(_10023_),
    .B1(_04972_));
 sg13g2_inv_1 _19119_ (.Y(_10024_),
    .A(_10023_));
 sg13g2_a21oi_1 _19120_ (.A1(_10024_),
    .A2(net27),
    .Y(_10025_),
    .B1(_06189_));
 sg13g2_inv_1 _19121_ (.Y(_10026_),
    .A(_10025_));
 sg13g2_a21oi_1 _19122_ (.A1(_10026_),
    .A2(net47),
    .Y(_10027_),
    .B1(_04220_));
 sg13g2_and2_1 _19123_ (.A(_10022_),
    .B(_10027_),
    .X(_10028_));
 sg13g2_nor4_1 _19124_ (.A(_09114_),
    .B(_10004_),
    .C(_10015_),
    .D(_10028_),
    .Y(_10029_));
 sg13g2_inv_1 _19125_ (.Y(_10030_),
    .A(_08917_));
 sg13g2_a21oi_1 _19126_ (.A1(_10030_),
    .A2(net81),
    .Y(_10031_),
    .B1(_04197_));
 sg13g2_a21oi_1 _19127_ (.A1(_08994_),
    .A2(net81),
    .Y(_10032_),
    .B1(_04280_));
 sg13g2_nor2_1 _19128_ (.A(_07509_),
    .B(_08965_),
    .Y(_10033_));
 sg13g2_a21oi_1 _19129_ (.A1(_10031_),
    .A2(_10032_),
    .Y(_10034_),
    .B1(_10033_));
 sg13g2_and2_1 _19130_ (.A(_10029_),
    .B(_10034_),
    .X(_10035_));
 sg13g2_nor2_2 _19131_ (.A(_09109_),
    .B(_04198_),
    .Y(_10036_));
 sg13g2_a21oi_1 _19132_ (.A1(_10021_),
    .A2(_08938_),
    .Y(_10037_),
    .B1(_10027_));
 sg13g2_inv_1 _19133_ (.Y(_10038_),
    .A(_08944_));
 sg13g2_o21ai_1 _19134_ (.B1(_10014_),
    .Y(_10039_),
    .A1(_10038_),
    .A2(_10009_));
 sg13g2_inv_1 _19135_ (.Y(_10040_),
    .A(_09090_));
 sg13g2_nor3_1 _19136_ (.A(_07934_),
    .B(_09737_),
    .C(_07936_),
    .Y(_10041_));
 sg13g2_nand4_1 _19137_ (.B(_10040_),
    .C(_09021_),
    .A(_10039_),
    .Y(_10042_),
    .D(_10041_));
 sg13g2_nor2_1 _19138_ (.A(_07509_),
    .B(_08966_),
    .Y(_10043_));
 sg13g2_nor2b_1 _19139_ (.A(_10031_),
    .B_N(_10032_),
    .Y(_10044_));
 sg13g2_nor2_1 _19140_ (.A(_10043_),
    .B(_10044_),
    .Y(_10045_));
 sg13g2_inv_1 _19141_ (.Y(_10046_),
    .A(_10045_));
 sg13g2_nor4_1 _19142_ (.A(_10036_),
    .B(_10037_),
    .C(_10042_),
    .D(_10046_),
    .Y(_10047_));
 sg13g2_nor3_1 _19143_ (.A(net159),
    .B(_10035_),
    .C(_10047_),
    .Y(_10048_));
 sg13g2_nand2_1 _19144_ (.Y(_10049_),
    .A(_10048_),
    .B(net145));
 sg13g2_nand2_1 _19145_ (.Y(_10050_),
    .A(_10047_),
    .B(_10035_));
 sg13g2_inv_1 _19146_ (.Y(_10051_),
    .A(_06163_));
 sg13g2_o21ai_1 _19147_ (.B1(_10051_),
    .Y(_10052_),
    .A1(_06154_),
    .A2(net159));
 sg13g2_nand3_1 _19148_ (.B(net86),
    .C(_10052_),
    .A(_10050_),
    .Y(_10053_));
 sg13g2_o21ai_1 _19149_ (.B1(_10053_),
    .Y(_10054_),
    .A1(_06154_),
    .A2(_10049_));
 sg13g2_nand3_1 _19150_ (.B(_10034_),
    .C(_10010_),
    .A(_10045_),
    .Y(_10055_));
 sg13g2_inv_1 _19151_ (.Y(_10056_),
    .A(net159));
 sg13g2_a21oi_1 _19152_ (.A1(_10021_),
    .A2(_05872_),
    .Y(_10057_),
    .B1(_10056_));
 sg13g2_a21oi_1 _19153_ (.A1(_10055_),
    .A2(_06158_),
    .Y(_10058_),
    .B1(_10057_));
 sg13g2_or2_1 _19154_ (.X(_10059_),
    .B(_10058_),
    .A(_06207_));
 sg13g2_nand2b_1 _19155_ (.Y(_10060_),
    .B(_10057_),
    .A_N(_06205_));
 sg13g2_nand3_1 _19156_ (.B(_06156_),
    .C(_10060_),
    .A(_10059_),
    .Y(_10061_));
 sg13g2_inv_1 _19157_ (.Y(_10062_),
    .A(_09109_));
 sg13g2_nor3_1 _19158_ (.A(_06156_),
    .B(_10062_),
    .C(_10038_),
    .Y(_10063_));
 sg13g2_nand3_1 _19159_ (.B(_08938_),
    .C(_09039_),
    .A(_10063_),
    .Y(_10064_));
 sg13g2_nor2_1 _19160_ (.A(net93),
    .B(_06159_),
    .Y(_10065_));
 sg13g2_and3_1 _19161_ (.X(_10066_),
    .A(_10061_),
    .B(_10064_),
    .C(_10065_));
 sg13g2_buf_1 _19162_ (.A(\b.gen_square[15].sq.mask ),
    .X(_10067_));
 sg13g2_o21ai_1 _19163_ (.B1(_10067_),
    .Y(_10068_),
    .A1(_10054_),
    .A2(_10066_));
 sg13g2_nor2_1 _19164_ (.A(_10068_),
    .B(_10001_),
    .Y(_10069_));
 sg13g2_nand2_1 _19165_ (.Y(_10070_),
    .A(_09999_),
    .B(_09979_));
 sg13g2_nand3_1 _19166_ (.B(_09997_),
    .C(_09976_),
    .A(_09995_),
    .Y(_10071_));
 sg13g2_nand3_1 _19167_ (.B(net96),
    .C(_10056_),
    .A(_10050_),
    .Y(_10072_));
 sg13g2_nand2_1 _19168_ (.Y(_10073_),
    .A(_10049_),
    .B(_10072_));
 sg13g2_nand2_1 _19169_ (.Y(_10074_),
    .A(_10049_),
    .B(_06163_));
 sg13g2_nand2b_1 _19170_ (.Y(_10075_),
    .B(_06162_),
    .A_N(_06206_));
 sg13g2_nand3_1 _19171_ (.B(_10074_),
    .C(_10075_),
    .A(_10073_),
    .Y(_10076_));
 sg13g2_nand3_1 _19172_ (.B(_06158_),
    .C(_07510_),
    .A(_10055_),
    .Y(_10077_));
 sg13g2_nand2_1 _19173_ (.Y(_10078_),
    .A(_10059_),
    .B(_10077_));
 sg13g2_nor2_1 _19174_ (.A(net93),
    .B(_08946_),
    .Y(_10079_));
 sg13g2_nand2_1 _19175_ (.Y(_10080_),
    .A(_10078_),
    .B(_10079_));
 sg13g2_nand2_1 _19176_ (.Y(_10081_),
    .A(_10076_),
    .B(_10080_));
 sg13g2_nand2_1 _19177_ (.Y(_10082_),
    .A(_10081_),
    .B(_10067_));
 sg13g2_nand3_1 _19178_ (.B(_10071_),
    .C(_10082_),
    .A(_10070_),
    .Y(_10083_));
 sg13g2_nand2_1 _19179_ (.Y(_10084_),
    .A(_10069_),
    .B(_10083_));
 sg13g2_nand2_1 _19180_ (.Y(_10085_),
    .A(_10070_),
    .B(_10071_));
 sg13g2_inv_1 _19181_ (.Y(_10086_),
    .A(_10082_));
 sg13g2_nor3_1 _19182_ (.A(_06153_),
    .B(_06151_),
    .C(_06204_),
    .Y(_10087_));
 sg13g2_nand2_1 _19183_ (.Y(_10088_),
    .A(net159),
    .B(_10087_));
 sg13g2_a21oi_1 _19184_ (.A1(_10041_),
    .A2(_10002_),
    .Y(_10089_),
    .B1(_10088_));
 sg13g2_nand2b_1 _19185_ (.Y(_10090_),
    .B(_10060_),
    .A_N(_10089_));
 sg13g2_xnor2_1 _19186_ (.Y(_10091_),
    .A(_06153_),
    .B(_06206_));
 sg13g2_a22oi_1 _19187_ (.Y(_10092_),
    .B1(_10091_),
    .B2(_10073_),
    .A2(_10079_),
    .A1(_10090_));
 sg13g2_nand2_1 _19188_ (.Y(_10093_),
    .A(_10092_),
    .B(_10080_));
 sg13g2_nand2_1 _19189_ (.Y(_10094_),
    .A(_10093_),
    .B(_10067_));
 sg13g2_nor2_1 _19190_ (.A(_09991_),
    .B(_09996_),
    .Y(_10095_));
 sg13g2_inv_1 _19191_ (.Y(_10096_),
    .A(_10095_));
 sg13g2_nor2_1 _19192_ (.A(_10094_),
    .B(_10096_),
    .Y(_10097_));
 sg13g2_a21oi_1 _19193_ (.A1(_10085_),
    .A2(_10086_),
    .Y(_10098_),
    .B1(_10097_));
 sg13g2_nand2_1 _19194_ (.Y(_10099_),
    .A(_10084_),
    .B(_10098_));
 sg13g2_nand2_1 _19195_ (.Y(_10100_),
    .A(_10096_),
    .B(_10094_));
 sg13g2_nand2_1 _19196_ (.Y(_10101_),
    .A(_10099_),
    .B(_10100_));
 sg13g2_buf_2 _19197_ (.A(_10101_),
    .X(_10102_));
 sg13g2_nand2b_1 _19198_ (.Y(_10103_),
    .B(_10102_),
    .A_N(_10001_));
 sg13g2_nand3_1 _19199_ (.B(_10100_),
    .C(_10068_),
    .A(_10099_),
    .Y(_10104_));
 sg13g2_nand2_1 _19200_ (.Y(_10105_),
    .A(_10103_),
    .B(_10104_));
 sg13g2_nor2_1 _19201_ (.A(_07130_),
    .B(_07082_),
    .Y(_10106_));
 sg13g2_a21o_1 _19202_ (.A2(_07074_),
    .A1(_07131_),
    .B1(net158),
    .X(_10107_));
 sg13g2_a21oi_1 _19203_ (.A1(_09830_),
    .A2(net49),
    .Y(_10108_),
    .B1(_08286_));
 sg13g2_inv_1 _19204_ (.Y(_10109_),
    .A(_10108_));
 sg13g2_a21oi_1 _19205_ (.A1(_09831_),
    .A2(_06955_),
    .Y(_10110_),
    .B1(_09289_));
 sg13g2_inv_1 _19206_ (.Y(_10111_),
    .A(_10110_));
 sg13g2_nor2_1 _19207_ (.A(_10109_),
    .B(_10111_),
    .Y(_10112_));
 sg13g2_nor4_1 _19208_ (.A(_09003_),
    .B(_10036_),
    .C(_09020_),
    .D(_09724_),
    .Y(_10113_));
 sg13g2_a21oi_1 _19209_ (.A1(_06727_),
    .A2(net90),
    .Y(_10114_),
    .B1(_04197_));
 sg13g2_a21oi_1 _19210_ (.A1(_06683_),
    .A2(net90),
    .Y(_10115_),
    .B1(_05317_));
 sg13g2_inv_1 _19211_ (.Y(_10116_),
    .A(_10115_));
 sg13g2_nor2_1 _19212_ (.A(_10114_),
    .B(_10116_),
    .Y(_10117_));
 sg13g2_inv_1 _19213_ (.Y(_10118_),
    .A(_10088_));
 sg13g2_a21oi_1 _19214_ (.A1(_04530_),
    .A2(_10118_),
    .Y(_10119_),
    .B1(_06211_));
 sg13g2_nor2_1 _19215_ (.A(_06166_),
    .B(_10119_),
    .Y(_10120_));
 sg13g2_a21oi_1 _19216_ (.A1(net133),
    .A2(_09770_),
    .Y(_10121_),
    .B1(_06527_));
 sg13g2_nor2_2 _19217_ (.A(_06806_),
    .B(_10121_),
    .Y(_10122_));
 sg13g2_nor2_1 _19218_ (.A(_07747_),
    .B(_10122_),
    .Y(_10123_));
 sg13g2_nand3b_1 _19219_ (.B(_10123_),
    .C(_09009_),
    .Y(_10124_),
    .A_N(_10120_));
 sg13g2_nor3_1 _19220_ (.A(_10117_),
    .B(_09131_),
    .C(_10124_),
    .Y(_10125_));
 sg13g2_nand3b_1 _19221_ (.B(_10113_),
    .C(_10125_),
    .Y(_10126_),
    .A_N(_10112_));
 sg13g2_nor2_1 _19222_ (.A(_05701_),
    .B(_09351_),
    .Y(_10127_));
 sg13g2_a21oi_1 _19223_ (.A1(_06000_),
    .A2(_05704_),
    .Y(_10128_),
    .B1(_10127_));
 sg13g2_inv_1 _19224_ (.Y(_10129_),
    .A(_10128_));
 sg13g2_nor2_1 _19225_ (.A(_06417_),
    .B(_06354_),
    .Y(_10130_));
 sg13g2_a21oi_1 _19226_ (.A1(_10129_),
    .A2(_06421_),
    .Y(_10131_),
    .B1(_10130_));
 sg13g2_inv_1 _19227_ (.Y(_10132_),
    .A(_10131_));
 sg13g2_nor2_1 _19228_ (.A(_06799_),
    .B(_06550_),
    .Y(_10133_));
 sg13g2_a21oi_1 _19229_ (.A1(_10132_),
    .A2(_06803_),
    .Y(_10134_),
    .B1(_10133_));
 sg13g2_inv_1 _19230_ (.Y(_10135_),
    .A(_10134_));
 sg13g2_nor2_1 _19231_ (.A(_06992_),
    .B(_06935_),
    .Y(_10136_));
 sg13g2_a21oi_1 _19232_ (.A1(_10135_),
    .A2(_06996_),
    .Y(_10137_),
    .B1(_10136_));
 sg13g2_inv_4 _19233_ (.A(_05704_),
    .Y(_10138_));
 sg13g2_nand2_1 _19234_ (.Y(_10139_),
    .A(_10138_),
    .B(_00014_));
 sg13g2_o21ai_1 _19235_ (.B1(_10139_),
    .Y(_10140_),
    .A1(_10138_),
    .A2(_09222_));
 sg13g2_buf_1 _19236_ (.A(_10140_),
    .X(_10141_));
 sg13g2_nor2b_1 _19237_ (.A(_06421_),
    .B_N(_00013_),
    .Y(_10142_));
 sg13g2_a21o_1 _19238_ (.A2(_06421_),
    .A1(_10141_),
    .B1(_10142_),
    .X(_10143_));
 sg13g2_buf_2 _19239_ (.A(_10143_),
    .X(_10144_));
 sg13g2_nor2b_1 _19240_ (.A(_06803_),
    .B_N(_00012_),
    .Y(_10145_));
 sg13g2_a21oi_2 _19241_ (.B1(_10145_),
    .Y(_10146_),
    .A2(_06803_),
    .A1(_10144_));
 sg13g2_a21oi_1 _19242_ (.A1(_10146_),
    .A2(_06996_),
    .Y(_10147_),
    .B1(_06998_));
 sg13g2_o21ai_1 _19243_ (.B1(_07096_),
    .Y(_10148_),
    .A1(_09291_),
    .A2(_09057_));
 sg13g2_a21oi_1 _19244_ (.A1(_09069_),
    .A2(net64),
    .Y(_10149_),
    .B1(_05950_));
 sg13g2_nand2_1 _19245_ (.Y(_10150_),
    .A(_07509_),
    .B(_04173_));
 sg13g2_nand3_1 _19246_ (.B(_04162_),
    .C(_04268_),
    .A(_04258_),
    .Y(_10151_));
 sg13g2_nand2_1 _19247_ (.Y(_10152_),
    .A(_10150_),
    .B(_10151_));
 sg13g2_nand2_1 _19248_ (.Y(_10153_),
    .A(_05522_),
    .B(_04173_));
 sg13g2_nand2_1 _19249_ (.Y(_10154_),
    .A(_04174_),
    .B(_00077_));
 sg13g2_nand2_1 _19250_ (.Y(_10155_),
    .A(_10153_),
    .B(_10154_));
 sg13g2_nand2b_1 _19251_ (.Y(_10156_),
    .B(_10155_),
    .A_N(_10152_));
 sg13g2_o21ai_1 _19252_ (.B1(_10156_),
    .Y(_10157_),
    .A1(_10148_),
    .A2(_10149_));
 sg13g2_a21oi_1 _19253_ (.A1(_10137_),
    .A2(_10147_),
    .Y(_10158_),
    .B1(_10157_));
 sg13g2_nor2b_1 _19254_ (.A(_10126_),
    .B_N(_10158_),
    .Y(_10159_));
 sg13g2_inv_1 _19255_ (.Y(_10160_),
    .A(_10159_));
 sg13g2_inv_1 _19256_ (.Y(_10161_),
    .A(_10147_));
 sg13g2_inv_1 _19257_ (.Y(_10162_),
    .A(_10148_));
 sg13g2_nand3_1 _19258_ (.B(_05520_),
    .C(_04009_),
    .A(_04173_),
    .Y(_10163_));
 sg13g2_a21oi_1 _19259_ (.A1(_10163_),
    .A2(_04176_),
    .Y(_10164_),
    .B1(_10152_));
 sg13g2_a221oi_1 _19260_ (.B2(_10162_),
    .C1(_10164_),
    .B1(_10149_),
    .A1(_10137_),
    .Y(_10165_),
    .A2(_10161_));
 sg13g2_nor2_1 _19261_ (.A(_08981_),
    .B(_10155_),
    .Y(_10166_));
 sg13g2_nor4_1 _19262_ (.A(_10166_),
    .B(_09114_),
    .C(_09156_),
    .D(_08934_),
    .Y(_10167_));
 sg13g2_o21ai_1 _19263_ (.B1(_10167_),
    .Y(_10168_),
    .A1(_09099_),
    .A2(_10110_));
 sg13g2_inv_1 _19264_ (.Y(_10169_),
    .A(_10168_));
 sg13g2_nor2_1 _19265_ (.A(_03231_),
    .B(_10119_),
    .Y(_10170_));
 sg13g2_nor2_2 _19266_ (.A(_02598_),
    .B(_10121_),
    .Y(_10171_));
 sg13g2_nor2_1 _19267_ (.A(_10170_),
    .B(_10171_),
    .Y(_10172_));
 sg13g2_nand2_1 _19268_ (.Y(_10173_),
    .A(_07839_),
    .B(_10172_));
 sg13g2_a221oi_1 _19269_ (.B2(_10108_),
    .C1(_10173_),
    .B1(_10111_),
    .A1(_10114_),
    .Y(_10174_),
    .A2(_10115_));
 sg13g2_nand3_1 _19270_ (.B(_10169_),
    .C(_10174_),
    .A(_10165_),
    .Y(_10175_));
 sg13g2_nor2_1 _19271_ (.A(_10160_),
    .B(_10175_),
    .Y(_10176_));
 sg13g2_nor3_1 _19272_ (.A(_10106_),
    .B(_10107_),
    .C(_10176_),
    .Y(_10177_));
 sg13g2_nand4_1 _19273_ (.B(_10160_),
    .C(net177),
    .A(_10175_),
    .Y(_10178_),
    .D(_07082_));
 sg13g2_buf_1 _19274_ (.A(_10178_),
    .X(_10179_));
 sg13g2_nor2_1 _19275_ (.A(_07074_),
    .B(_10179_),
    .Y(_10180_));
 sg13g2_a21oi_1 _19276_ (.A1(_10109_),
    .A2(_10116_),
    .Y(_10181_),
    .B1(_07082_));
 sg13g2_a21oi_1 _19277_ (.A1(_10165_),
    .A2(_10158_),
    .Y(_10182_),
    .B1(_07082_));
 sg13g2_o21ai_1 _19278_ (.B1(_07079_),
    .Y(_10183_),
    .A1(_10181_),
    .A2(_10182_));
 sg13g2_nand3_1 _19279_ (.B(_07073_),
    .C(_08278_),
    .A(_10181_),
    .Y(_10184_));
 sg13g2_nand3_1 _19280_ (.B(_07088_),
    .C(_10184_),
    .A(_10183_),
    .Y(_10185_));
 sg13g2_nand4_1 _19281_ (.B(_08983_),
    .C(_10113_),
    .A(_10169_),
    .Y(_10186_),
    .D(_09132_));
 sg13g2_nor2_1 _19282_ (.A(net120),
    .B(_07089_),
    .Y(_10187_));
 sg13g2_nand3_1 _19283_ (.B(_10186_),
    .C(_10187_),
    .A(_10185_),
    .Y(_10188_));
 sg13g2_nand2b_1 _19284_ (.Y(_10189_),
    .B(_10188_),
    .A_N(_10180_));
 sg13g2_buf_1 _19285_ (.A(\b.gen_square[5].sq.mask ),
    .X(_10190_));
 sg13g2_o21ai_1 _19286_ (.B1(_10190_),
    .Y(_10191_),
    .A1(_10177_),
    .A2(_10189_));
 sg13g2_nor2_1 _19287_ (.A(_06992_),
    .B(_06932_),
    .Y(_10192_));
 sg13g2_o21ai_1 _19288_ (.B1(net161),
    .Y(_10193_),
    .A1(_06921_),
    .A2(_06992_));
 sg13g2_a21oi_1 _19289_ (.A1(_09853_),
    .A2(_06955_),
    .Y(_10194_),
    .B1(_07002_));
 sg13g2_inv_1 _19290_ (.Y(_10195_),
    .A(_10194_));
 sg13g2_inv_1 _19291_ (.Y(_10196_),
    .A(_09819_));
 sg13g2_a21oi_1 _19292_ (.A1(_10196_),
    .A2(net49),
    .Y(_10197_),
    .B1(_06964_));
 sg13g2_nand2_1 _19293_ (.Y(_10198_),
    .A(_10152_),
    .B(_07133_));
 sg13g2_nand2_1 _19294_ (.Y(_10199_),
    .A(_07092_),
    .B(_07131_));
 sg13g2_nand2_1 _19295_ (.Y(_10200_),
    .A(_10198_),
    .B(_10199_));
 sg13g2_nand3_1 _19296_ (.B(_07133_),
    .C(_10154_),
    .A(_10153_),
    .Y(_10201_));
 sg13g2_nand2_1 _19297_ (.Y(_10202_),
    .A(_10201_),
    .B(_07137_));
 sg13g2_nor2_1 _19298_ (.A(_10200_),
    .B(_10202_),
    .Y(_10203_));
 sg13g2_a21oi_1 _19299_ (.A1(_10195_),
    .A2(_10197_),
    .Y(_10204_),
    .B1(_10203_));
 sg13g2_inv_1 _19300_ (.Y(_10205_),
    .A(_10146_));
 sg13g2_a21oi_1 _19301_ (.A1(_10205_),
    .A2(_09908_),
    .Y(_10206_),
    .B1(_09542_));
 sg13g2_inv_1 _19302_ (.Y(_10207_),
    .A(_09085_));
 sg13g2_a21oi_1 _19303_ (.A1(_10207_),
    .A2(net64),
    .Y(_10208_),
    .B1(_05950_));
 sg13g2_a21oi_1 _19304_ (.A1(_09089_),
    .A2(_05890_),
    .Y(_10209_),
    .B1(_05899_));
 sg13g2_nor2_1 _19305_ (.A(_09857_),
    .B(_10209_),
    .Y(_10210_));
 sg13g2_a21oi_1 _19306_ (.A1(net88),
    .A2(_09982_),
    .Y(_10211_),
    .B1(_04192_));
 sg13g2_inv_1 _19307_ (.Y(_10212_),
    .A(_10211_));
 sg13g2_nand2_1 _19308_ (.Y(_10213_),
    .A(_10212_),
    .B(_00038_));
 sg13g2_inv_1 _19309_ (.Y(_10214_),
    .A(_10213_));
 sg13g2_inv_1 _19310_ (.Y(_10215_),
    .A(_09636_));
 sg13g2_a21oi_2 _19311_ (.B1(_06331_),
    .Y(_10216_),
    .A2(_10215_),
    .A1(net115));
 sg13g2_o21ai_1 _19312_ (.B1(_07939_),
    .Y(_10217_),
    .A1(_06424_),
    .A2(_10216_));
 sg13g2_nor3_1 _19313_ (.A(_07936_),
    .B(_10214_),
    .C(_10217_),
    .Y(_10218_));
 sg13g2_o21ai_1 _19314_ (.B1(_10218_),
    .Y(_10219_),
    .A1(_10208_),
    .A2(_10210_));
 sg13g2_o21ai_1 _19315_ (.B1(_08165_),
    .Y(_10220_),
    .A1(_08909_),
    .A2(_09676_));
 sg13g2_o21ai_1 _19316_ (.B1(_09296_),
    .Y(_10221_),
    .A1(_08909_),
    .A2(_09673_));
 sg13g2_nor2_1 _19317_ (.A(_10220_),
    .B(_10221_),
    .Y(_10222_));
 sg13g2_nor2_1 _19318_ (.A(_10146_),
    .B(_10135_),
    .Y(_10223_));
 sg13g2_nor3_1 _19319_ (.A(_10219_),
    .B(_10222_),
    .C(_10223_),
    .Y(_10224_));
 sg13g2_nand3_1 _19320_ (.B(_07133_),
    .C(_04176_),
    .A(_10163_),
    .Y(_10225_));
 sg13g2_nand2_1 _19321_ (.Y(_10226_),
    .A(_07134_),
    .B(_03959_));
 sg13g2_nand2_1 _19322_ (.Y(_10227_),
    .A(_10225_),
    .B(_10226_));
 sg13g2_a21oi_1 _19323_ (.A1(_10227_),
    .A2(_09040_),
    .Y(_10228_),
    .B1(_09101_));
 sg13g2_nand4_1 _19324_ (.B(_10206_),
    .C(_10224_),
    .A(_10204_),
    .Y(_10229_),
    .D(_10228_));
 sg13g2_inv_1 _19325_ (.Y(_10230_),
    .A(_09541_));
 sg13g2_nand2_1 _19326_ (.Y(_10231_),
    .A(_10146_),
    .B(_09908_));
 sg13g2_inv_1 _19327_ (.Y(_10232_),
    .A(_09113_));
 sg13g2_nand4_1 _19328_ (.B(_10232_),
    .C(_08935_),
    .A(_10231_),
    .Y(_10233_),
    .D(_09155_));
 sg13g2_a21oi_1 _19329_ (.A1(_10230_),
    .A2(_10221_),
    .Y(_10234_),
    .B1(_10233_));
 sg13g2_inv_1 _19330_ (.Y(_10235_),
    .A(_10234_));
 sg13g2_nand2b_1 _19331_ (.Y(_10236_),
    .B(_10221_),
    .A_N(_10220_));
 sg13g2_nand2_1 _19332_ (.Y(_10237_),
    .A(_10209_),
    .B(_10208_));
 sg13g2_nor2_1 _19333_ (.A(_02393_),
    .B(_10216_),
    .Y(_10238_));
 sg13g2_nor2_1 _19334_ (.A(_07919_),
    .B(_10238_),
    .Y(_10239_));
 sg13g2_inv_1 _19335_ (.Y(_10240_),
    .A(_10239_));
 sg13g2_nor2_1 _19336_ (.A(_03080_),
    .B(_10211_),
    .Y(_10241_));
 sg13g2_nor2_1 _19337_ (.A(_10241_),
    .B(_07902_),
    .Y(_10242_));
 sg13g2_inv_1 _19338_ (.Y(_10243_),
    .A(_10242_));
 sg13g2_nor2_1 _19339_ (.A(_10240_),
    .B(_10243_),
    .Y(_10244_));
 sg13g2_nand3_1 _19340_ (.B(_10237_),
    .C(_10244_),
    .A(_10236_),
    .Y(_10245_));
 sg13g2_a22oi_1 _19341_ (.Y(_10246_),
    .B1(_10197_),
    .B2(_10194_),
    .A2(_10146_),
    .A1(_10134_));
 sg13g2_o21ai_1 _19342_ (.B1(_10246_),
    .Y(_10247_),
    .A1(_10200_),
    .A2(_10227_));
 sg13g2_nor3_1 _19343_ (.A(_10235_),
    .B(_10245_),
    .C(_10247_),
    .Y(_10248_));
 sg13g2_inv_1 _19344_ (.Y(_10249_),
    .A(_10248_));
 sg13g2_nor2_1 _19345_ (.A(_10229_),
    .B(_10249_),
    .Y(_10250_));
 sg13g2_nor3_1 _19346_ (.A(_10192_),
    .B(_10193_),
    .C(_10250_),
    .Y(_10251_));
 sg13g2_inv_1 _19347_ (.Y(_10252_),
    .A(_10209_));
 sg13g2_a21oi_1 _19348_ (.A1(_10220_),
    .A2(_10252_),
    .Y(_10253_),
    .B1(_06932_));
 sg13g2_nor2_1 _19349_ (.A(_10223_),
    .B(_10247_),
    .Y(_10254_));
 sg13g2_a21oi_1 _19350_ (.A1(_10254_),
    .A2(_10204_),
    .Y(_10255_),
    .B1(_06932_));
 sg13g2_o21ai_1 _19351_ (.B1(_06929_),
    .Y(_10256_),
    .A1(_10253_),
    .A2(_10255_));
 sg13g2_nand3_1 _19352_ (.B(_06919_),
    .C(_08157_),
    .A(_10253_),
    .Y(_10257_));
 sg13g2_nand3_1 _19353_ (.B(_06923_),
    .C(_10257_),
    .A(_10256_),
    .Y(_10258_));
 sg13g2_nor2_1 _19354_ (.A(_06923_),
    .B(_09003_),
    .Y(_10259_));
 sg13g2_nand4_1 _19355_ (.B(_10206_),
    .C(_10228_),
    .A(_10234_),
    .Y(_10260_),
    .D(_10259_));
 sg13g2_nor2_1 _19356_ (.A(net137),
    .B(_06924_),
    .Y(_10261_));
 sg13g2_nand3_1 _19357_ (.B(_10260_),
    .C(_10261_),
    .A(_10258_),
    .Y(_10262_));
 sg13g2_nand4_1 _19358_ (.B(net191),
    .C(_10229_),
    .A(_10249_),
    .Y(_10263_),
    .D(_06932_));
 sg13g2_buf_1 _19359_ (.A(_10263_),
    .X(_10264_));
 sg13g2_nand2b_1 _19360_ (.Y(_10265_),
    .B(_06921_),
    .A_N(_10264_));
 sg13g2_nand3b_1 _19361_ (.B(_10262_),
    .C(_10265_),
    .Y(_10266_),
    .A_N(_10251_));
 sg13g2_buf_1 _19362_ (.A(\b.gen_square[4].sq.mask ),
    .X(_10267_));
 sg13g2_nand2_1 _19363_ (.Y(_10268_),
    .A(_10266_),
    .B(_10267_));
 sg13g2_inv_1 _19364_ (.Y(_10269_),
    .A(_09719_));
 sg13g2_nand2_1 _19365_ (.Y(_10270_),
    .A(_10269_),
    .B(_09538_));
 sg13g2_o21ai_1 _19366_ (.B1(_08165_),
    .Y(_10271_),
    .A1(_08909_),
    .A2(_09686_));
 sg13g2_a21oi_1 _19367_ (.A1(_09681_),
    .A2(_06530_),
    .Y(_10272_),
    .B1(_06808_));
 sg13g2_a21oi_1 _19368_ (.A1(_10271_),
    .A2(_09541_),
    .Y(_10273_),
    .B1(_10272_));
 sg13g2_a21oi_1 _19369_ (.A1(_10141_),
    .A2(_09472_),
    .Y(_10274_),
    .B1(_09260_));
 sg13g2_inv_1 _19370_ (.Y(_10275_),
    .A(_09896_));
 sg13g2_a21oi_1 _19371_ (.A1(_04508_),
    .A2(_10275_),
    .Y(_10276_),
    .B1(_06952_));
 sg13g2_nor2_2 _19372_ (.A(_07000_),
    .B(_10276_),
    .Y(_10277_));
 sg13g2_a21o_1 _19373_ (.A2(_09503_),
    .A1(_04508_),
    .B1(_05993_),
    .X(_10278_));
 sg13g2_nand2_1 _19374_ (.Y(_10279_),
    .A(_10278_),
    .B(_00066_));
 sg13g2_inv_1 _19375_ (.Y(_10280_),
    .A(_10279_));
 sg13g2_nor3_1 _19376_ (.A(_10277_),
    .B(_10280_),
    .C(_08113_),
    .Y(_10281_));
 sg13g2_inv_1 _19377_ (.Y(_10282_),
    .A(_10141_));
 sg13g2_nor2_1 _19378_ (.A(_10129_),
    .B(_10282_),
    .Y(_10283_));
 sg13g2_inv_1 _19379_ (.Y(_10284_),
    .A(_10283_));
 sg13g2_a21oi_1 _19380_ (.A1(_06876_),
    .A2(net43),
    .Y(_10285_),
    .B1(_04867_));
 sg13g2_nand2_1 _19381_ (.Y(_10286_),
    .A(_09258_),
    .B(_10285_));
 sg13g2_nand4_1 _19382_ (.B(_10281_),
    .C(_10284_),
    .A(_10274_),
    .Y(_10287_),
    .D(_10286_));
 sg13g2_o21ai_1 _19383_ (.B1(_09240_),
    .Y(_10288_),
    .A1(_08901_),
    .A2(_09584_));
 sg13g2_a21oi_1 _19384_ (.A1(_09587_),
    .A2(net37),
    .Y(_10289_),
    .B1(_06363_));
 sg13g2_nand2_1 _19385_ (.Y(_10290_),
    .A(_10288_),
    .B(_10289_));
 sg13g2_nand2_1 _19386_ (.Y(_10291_),
    .A(_10200_),
    .B(_06996_));
 sg13g2_inv_1 _19387_ (.Y(_10292_),
    .A(_10136_));
 sg13g2_nand2_1 _19388_ (.Y(_10293_),
    .A(_10291_),
    .B(_10292_));
 sg13g2_nand2_1 _19389_ (.Y(_10294_),
    .A(_10293_),
    .B(_06803_));
 sg13g2_inv_1 _19390_ (.Y(_10295_),
    .A(_10133_));
 sg13g2_nand2_1 _19391_ (.Y(_10296_),
    .A(_10294_),
    .B(_10295_));
 sg13g2_inv_1 _19392_ (.Y(_10297_),
    .A(_10296_));
 sg13g2_nand3_1 _19393_ (.B(_06996_),
    .C(_07137_),
    .A(_10201_),
    .Y(_10298_));
 sg13g2_inv_1 _19394_ (.Y(_10299_),
    .A(_06996_));
 sg13g2_nand2_1 _19395_ (.Y(_10300_),
    .A(_10299_),
    .B(_00055_));
 sg13g2_nand2_1 _19396_ (.Y(_10301_),
    .A(_10298_),
    .B(_10300_));
 sg13g2_nand2_1 _19397_ (.Y(_10302_),
    .A(_10301_),
    .B(_06803_));
 sg13g2_inv_1 _19398_ (.Y(_10303_),
    .A(_10145_));
 sg13g2_nand2_1 _19399_ (.Y(_10304_),
    .A(_10302_),
    .B(_10303_));
 sg13g2_nand2_1 _19400_ (.Y(_10305_),
    .A(_10297_),
    .B(_10304_));
 sg13g2_nand2_1 _19401_ (.Y(_10306_),
    .A(_10290_),
    .B(_10305_));
 sg13g2_nor3_1 _19402_ (.A(_10273_),
    .B(_10287_),
    .C(_10306_),
    .Y(_10307_));
 sg13g2_nand2b_1 _19403_ (.Y(_10308_),
    .B(_10307_),
    .A_N(_10270_));
 sg13g2_nand3_1 _19404_ (.B(_06996_),
    .C(_10226_),
    .A(_10225_),
    .Y(_10309_));
 sg13g2_nand2_1 _19405_ (.Y(_10310_),
    .A(_10299_),
    .B(_03870_));
 sg13g2_nand2_1 _19406_ (.Y(_10311_),
    .A(_10309_),
    .B(_10310_));
 sg13g2_nand2_1 _19407_ (.Y(_10312_),
    .A(_10311_),
    .B(_06803_));
 sg13g2_nand2_1 _19408_ (.Y(_10313_),
    .A(_10312_),
    .B(_06805_));
 sg13g2_nor2b_1 _19409_ (.A(_10288_),
    .B_N(_10289_),
    .Y(_10314_));
 sg13g2_a21oi_1 _19410_ (.A1(_10297_),
    .A2(_10313_),
    .Y(_10315_),
    .B1(_10314_));
 sg13g2_inv_1 _19411_ (.Y(_10316_),
    .A(_09256_));
 sg13g2_inv_1 _19412_ (.Y(_10317_),
    .A(_09431_));
 sg13g2_inv_1 _19413_ (.Y(_10318_),
    .A(_09608_));
 sg13g2_nand2_1 _19414_ (.Y(_10319_),
    .A(_10282_),
    .B(_09472_));
 sg13g2_nand4_1 _19415_ (.B(_10317_),
    .C(_10318_),
    .A(_10231_),
    .Y(_10320_),
    .D(_10319_));
 sg13g2_a21oi_1 _19416_ (.A1(_10316_),
    .A2(_09259_),
    .Y(_10321_),
    .B1(_10320_));
 sg13g2_nand2b_1 _19417_ (.Y(_10322_),
    .B(_10272_),
    .A_N(_10271_));
 sg13g2_nand2_1 _19418_ (.Y(_10323_),
    .A(_09259_),
    .B(_10285_));
 sg13g2_nor2_1 _19419_ (.A(_09288_),
    .B(_10276_),
    .Y(_10324_));
 sg13g2_inv_1 _19420_ (.Y(_10325_),
    .A(_10324_));
 sg13g2_nand2_1 _19421_ (.Y(_10326_),
    .A(_10278_),
    .B(\b.gen_square[8].sq.color ));
 sg13g2_and3_1 _19422_ (.X(_10327_),
    .A(_08047_),
    .B(_10325_),
    .C(_10326_));
 sg13g2_nand3_1 _19423_ (.B(_10323_),
    .C(_10327_),
    .A(_10322_),
    .Y(_10328_));
 sg13g2_a21oi_1 _19424_ (.A1(_10128_),
    .A2(_10282_),
    .Y(_10329_),
    .B1(_10328_));
 sg13g2_nand3_1 _19425_ (.B(_10321_),
    .C(_10329_),
    .A(_10315_),
    .Y(_10330_));
 sg13g2_nand4_1 _19426_ (.B(_10330_),
    .C(_05072_),
    .A(_10308_),
    .Y(_10331_),
    .D(_06351_));
 sg13g2_buf_1 _19427_ (.A(_10331_),
    .X(_10332_));
 sg13g2_a22oi_1 _19428_ (.Y(_10333_),
    .B1(_06417_),
    .B2(_10332_),
    .A2(_06349_),
    .A1(_06347_));
 sg13g2_nor2_1 _19429_ (.A(_10330_),
    .B(_10308_),
    .Y(_10334_));
 sg13g2_inv_2 _19430_ (.Y(_10335_),
    .A(_10334_));
 sg13g2_nand3_1 _19431_ (.B(_04044_),
    .C(_06351_),
    .A(_10335_),
    .Y(_10336_));
 sg13g2_nand2_1 _19432_ (.Y(_10337_),
    .A(_10336_),
    .B(_10332_));
 sg13g2_inv_1 _19433_ (.Y(_10338_),
    .A(_10285_));
 sg13g2_a21oi_1 _19434_ (.A1(_10271_),
    .A2(_10338_),
    .Y(_10339_),
    .B1(_06351_));
 sg13g2_nor2_1 _19435_ (.A(_10128_),
    .B(_10306_),
    .Y(_10340_));
 sg13g2_a21oi_1 _19436_ (.A1(_10315_),
    .A2(_10340_),
    .Y(_10341_),
    .B1(_06351_));
 sg13g2_o21ai_1 _19437_ (.B1(_06348_),
    .Y(_10342_),
    .A1(_10339_),
    .A2(_10341_));
 sg13g2_nand2_1 _19438_ (.Y(_10343_),
    .A(_10341_),
    .B(_06350_));
 sg13g2_a21oi_1 _19439_ (.A1(_10342_),
    .A2(_10343_),
    .Y(_10344_),
    .B1(net154));
 sg13g2_a21o_1 _19440_ (.A2(_10337_),
    .A1(_10333_),
    .B1(_10344_),
    .X(_10345_));
 sg13g2_nand2_1 _19441_ (.Y(_10346_),
    .A(_10345_),
    .B(\b.gen_square[2].sq.mask ));
 sg13g2_nor2_1 _19442_ (.A(_06424_),
    .B(_10216_),
    .Y(_10347_));
 sg13g2_nor2_1 _19443_ (.A(_10347_),
    .B(_08111_),
    .Y(_10348_));
 sg13g2_inv_1 _19444_ (.Y(_10349_),
    .A(_10348_));
 sg13g2_nor2_1 _19445_ (.A(_09395_),
    .B(_06104_),
    .Y(_10350_));
 sg13g2_nor2_1 _19446_ (.A(_09225_),
    .B(_10350_),
    .Y(_10351_));
 sg13g2_inv_1 _19447_ (.Y(_10352_),
    .A(_10351_));
 sg13g2_nor2_1 _19448_ (.A(_10349_),
    .B(_10352_),
    .Y(_10353_));
 sg13g2_inv_1 _19449_ (.Y(_10354_),
    .A(_10353_));
 sg13g2_nand2_1 _19450_ (.Y(_10355_),
    .A(_09180_),
    .B(_05995_));
 sg13g2_inv_1 _19451_ (.Y(_10356_),
    .A(_06103_));
 sg13g2_nand2_1 _19452_ (.Y(_10357_),
    .A(_10355_),
    .B(_10356_));
 sg13g2_nand2_1 _19453_ (.Y(_10358_),
    .A(_09186_),
    .B(_06030_));
 sg13g2_nand2b_1 _19454_ (.Y(_10359_),
    .B(_10358_),
    .A_N(_06039_));
 sg13g2_a21oi_2 _19455_ (.B1(_06010_),
    .Y(_10360_),
    .A2(_05995_),
    .A1(_10359_));
 sg13g2_nand2_1 _19456_ (.Y(_10361_),
    .A(_10357_),
    .B(_10360_));
 sg13g2_inv_1 _19457_ (.Y(_10362_),
    .A(_09533_));
 sg13g2_nand2_1 _19458_ (.Y(_10363_),
    .A(_10361_),
    .B(_10362_));
 sg13g2_nand2_1 _19459_ (.Y(_10364_),
    .A(_09356_),
    .B(net59));
 sg13g2_nand2_1 _19460_ (.Y(_10365_),
    .A(_10364_),
    .B(_09243_));
 sg13g2_nand2_1 _19461_ (.Y(_10366_),
    .A(_09362_),
    .B(net59));
 sg13g2_nand2_1 _19462_ (.Y(_10367_),
    .A(_10366_),
    .B(_04866_));
 sg13g2_inv_2 _19463_ (.Y(_10368_),
    .A(_10367_));
 sg13g2_nand2_1 _19464_ (.Y(_10369_),
    .A(_10365_),
    .B(_10368_));
 sg13g2_nand2_1 _19465_ (.Y(_10370_),
    .A(_10304_),
    .B(_06421_));
 sg13g2_inv_1 _19466_ (.Y(_10371_),
    .A(_10142_));
 sg13g2_nand2_1 _19467_ (.Y(_10372_),
    .A(_10370_),
    .B(_10371_));
 sg13g2_nand2_1 _19468_ (.Y(_10373_),
    .A(_10372_),
    .B(_05704_));
 sg13g2_nand2_1 _19469_ (.Y(_10374_),
    .A(_10373_),
    .B(_10139_));
 sg13g2_nand2_1 _19470_ (.Y(_10375_),
    .A(_10296_),
    .B(_06421_));
 sg13g2_inv_1 _19471_ (.Y(_10376_),
    .A(_10130_));
 sg13g2_nand2_1 _19472_ (.Y(_10377_),
    .A(_10375_),
    .B(_10376_));
 sg13g2_a21oi_1 _19473_ (.A1(_10377_),
    .A2(_05704_),
    .Y(_10378_),
    .B1(_10127_));
 sg13g2_nand2_1 _19474_ (.Y(_10379_),
    .A(_10374_),
    .B(_10378_));
 sg13g2_nand2_1 _19475_ (.Y(_10380_),
    .A(_10369_),
    .B(_10379_));
 sg13g2_nor3_1 _19476_ (.A(_10354_),
    .B(_10363_),
    .C(_10380_),
    .Y(_10381_));
 sg13g2_a21oi_1 _19477_ (.A1(_09180_),
    .A2(_05995_),
    .Y(_10382_),
    .B1(_06103_));
 sg13g2_nand2_1 _19478_ (.Y(_10383_),
    .A(_10382_),
    .B(_10360_));
 sg13g2_nand2_1 _19479_ (.Y(_10384_),
    .A(_10313_),
    .B(_06421_));
 sg13g2_nand2_1 _19480_ (.Y(_10385_),
    .A(_10384_),
    .B(_06423_));
 sg13g2_nand2_1 _19481_ (.Y(_10386_),
    .A(_10385_),
    .B(_05704_));
 sg13g2_nand2_1 _19482_ (.Y(_10387_),
    .A(_10386_),
    .B(_05706_));
 sg13g2_nand2_1 _19483_ (.Y(_10388_),
    .A(_10387_),
    .B(_10378_));
 sg13g2_nand2_1 _19484_ (.Y(_10389_),
    .A(_10383_),
    .B(_10388_));
 sg13g2_a21oi_1 _19485_ (.A1(_09356_),
    .A2(net43),
    .Y(_10390_),
    .B1(_04956_));
 sg13g2_nand2_1 _19486_ (.Y(_10391_),
    .A(_10390_),
    .B(_10368_));
 sg13g2_nor2_2 _19487_ (.A(_08046_),
    .B(_10238_),
    .Y(_10392_));
 sg13g2_nor2_1 _19488_ (.A(_09395_),
    .B(_06105_),
    .Y(_10393_));
 sg13g2_nand2b_1 _19489_ (.Y(_10394_),
    .B(_10319_),
    .A_N(_10393_));
 sg13g2_nor2_1 _19490_ (.A(_09307_),
    .B(_10394_),
    .Y(_10395_));
 sg13g2_nand3_1 _19491_ (.B(_10392_),
    .C(_10395_),
    .A(_10391_),
    .Y(_10396_));
 sg13g2_nor2_1 _19492_ (.A(_10389_),
    .B(_10396_),
    .Y(_10397_));
 sg13g2_nand2_1 _19493_ (.Y(_10398_),
    .A(_10381_),
    .B(_10397_));
 sg13g2_nor2_1 _19494_ (.A(_04261_),
    .B(net131),
    .Y(_10399_));
 sg13g2_nand2_1 _19495_ (.Y(_10400_),
    .A(_10398_),
    .B(_10399_));
 sg13g2_inv_1 _19496_ (.Y(_10401_),
    .A(_10379_));
 sg13g2_nor2_1 _19497_ (.A(_10367_),
    .B(_10390_),
    .Y(_10402_));
 sg13g2_nor2_1 _19498_ (.A(_10401_),
    .B(_10402_),
    .Y(_10403_));
 sg13g2_a21oi_1 _19499_ (.A1(_10357_),
    .A2(_10360_),
    .Y(_10404_),
    .B1(_09533_));
 sg13g2_nand3_1 _19500_ (.B(_10404_),
    .C(_10353_),
    .A(_10403_),
    .Y(_10405_));
 sg13g2_a21oi_1 _19501_ (.A1(_10367_),
    .A2(_09256_),
    .Y(_10406_),
    .B1(_10365_));
 sg13g2_nor2b_1 _19502_ (.A(_10406_),
    .B_N(_10383_),
    .Y(_10407_));
 sg13g2_nand2_1 _19503_ (.Y(_10408_),
    .A(_10388_),
    .B(_10392_));
 sg13g2_nor2_1 _19504_ (.A(_10394_),
    .B(_10408_),
    .Y(_10409_));
 sg13g2_nand2_1 _19505_ (.Y(_10410_),
    .A(_10407_),
    .B(_10409_));
 sg13g2_nor2_1 _19506_ (.A(net192),
    .B(net131),
    .Y(_10411_));
 sg13g2_nand3_1 _19507_ (.B(_10410_),
    .C(_10411_),
    .A(_10405_),
    .Y(_10412_));
 sg13g2_buf_1 _19508_ (.A(_10412_),
    .X(_10413_));
 sg13g2_nand2_1 _19509_ (.Y(_10414_),
    .A(_10400_),
    .B(_10413_));
 sg13g2_nand2_1 _19510_ (.Y(_10415_),
    .A(_10413_),
    .B(_04841_));
 sg13g2_nand2_1 _19511_ (.Y(_10416_),
    .A(_04847_),
    .B(_04840_));
 sg13g2_nand3_1 _19512_ (.B(_10415_),
    .C(_10416_),
    .A(_10414_),
    .Y(_10417_));
 sg13g2_inv_1 _19513_ (.Y(_10418_),
    .A(_10360_));
 sg13g2_nand3_1 _19514_ (.B(_10379_),
    .C(_10418_),
    .A(_10388_),
    .Y(_10419_));
 sg13g2_nand2_1 _19515_ (.Y(_10420_),
    .A(_10419_),
    .B(net131));
 sg13g2_nand2_1 _19516_ (.Y(_10421_),
    .A(_10368_),
    .B(net131));
 sg13g2_nand2_1 _19517_ (.Y(_10422_),
    .A(_10420_),
    .B(_10421_));
 sg13g2_nand2_1 _19518_ (.Y(_10423_),
    .A(_10422_),
    .B(_05997_));
 sg13g2_nand3_1 _19519_ (.B(_04843_),
    .C(_05996_),
    .A(_10419_),
    .Y(_10424_));
 sg13g2_nand2_1 _19520_ (.Y(_10425_),
    .A(_10423_),
    .B(_10424_));
 sg13g2_nor2_1 _19521_ (.A(_02023_),
    .B(_09218_),
    .Y(_10426_));
 sg13g2_nand2_1 _19522_ (.Y(_10427_),
    .A(_10425_),
    .B(_10426_));
 sg13g2_buf_1 _19523_ (.A(\b.gen_square[0].sq.mask ),
    .X(_10428_));
 sg13g2_inv_1 _19524_ (.Y(_10429_),
    .A(_10428_));
 sg13g2_a21oi_1 _19525_ (.A1(_10417_),
    .A2(_10427_),
    .Y(_10430_),
    .B1(_10429_));
 sg13g2_a21oi_1 _19526_ (.A1(_10296_),
    .A2(_06421_),
    .Y(_10431_),
    .B1(_10130_));
 sg13g2_a21o_1 _19527_ (.A2(_10431_),
    .A1(_10385_),
    .B1(_09277_),
    .X(_10432_));
 sg13g2_nand2_1 _19528_ (.Y(_10433_),
    .A(_09342_),
    .B(net59));
 sg13g2_nand2_1 _19529_ (.Y(_10434_),
    .A(_10433_),
    .B(_09243_));
 sg13g2_a21oi_1 _19530_ (.A1(_09348_),
    .A2(net59),
    .Y(_10435_),
    .B1(_05616_));
 sg13g2_nor2b_1 _19531_ (.A(_10434_),
    .B_N(_10435_),
    .Y(_10436_));
 sg13g2_nor2_1 _19532_ (.A(_10432_),
    .B(_10436_),
    .Y(_10437_));
 sg13g2_nand2_1 _19533_ (.Y(_10438_),
    .A(_10372_),
    .B(_10431_));
 sg13g2_nand2b_1 _19534_ (.Y(_10439_),
    .B(_10438_),
    .A_N(_09227_));
 sg13g2_a21oi_1 _19535_ (.A1(_10434_),
    .A2(_10435_),
    .Y(_10440_),
    .B1(_10439_));
 sg13g2_nand2_1 _19536_ (.Y(_10441_),
    .A(_10437_),
    .B(_10440_));
 sg13g2_nand2_1 _19537_ (.Y(_10442_),
    .A(_10441_),
    .B(_05602_));
 sg13g2_nand2_1 _19538_ (.Y(_10443_),
    .A(_09555_),
    .B(net37));
 sg13g2_nand2_1 _19539_ (.Y(_10444_),
    .A(_10443_),
    .B(_09300_));
 sg13g2_a21oi_1 _19540_ (.A1(_09569_),
    .A2(net37),
    .Y(_10445_),
    .B1(_07583_));
 sg13g2_nand2_1 _19541_ (.Y(_10446_),
    .A(_10444_),
    .B(_10445_));
 sg13g2_nand2_1 _19542_ (.Y(_10447_),
    .A(_09571_),
    .B(_06334_));
 sg13g2_nand2_1 _19543_ (.Y(_10448_),
    .A(_10447_),
    .B(_09240_));
 sg13g2_nand2_1 _19544_ (.Y(_10449_),
    .A(_10448_),
    .B(_10445_));
 sg13g2_nand3_1 _19545_ (.B(_10449_),
    .C(_07191_),
    .A(_10446_),
    .Y(_10450_));
 sg13g2_nand2_1 _19546_ (.Y(_10451_),
    .A(_10450_),
    .B(_05602_));
 sg13g2_nand2_1 _19547_ (.Y(_10452_),
    .A(_10442_),
    .B(_10451_));
 sg13g2_nand2_1 _19548_ (.Y(_10453_),
    .A(_10452_),
    .B(_05599_));
 sg13g2_nand3_1 _19549_ (.B(_05602_),
    .C(_05595_),
    .A(_10441_),
    .Y(_10454_));
 sg13g2_nand2_1 _19550_ (.Y(_10455_),
    .A(_10453_),
    .B(_10454_));
 sg13g2_nor2_1 _19551_ (.A(_02023_),
    .B(_05608_),
    .Y(_10456_));
 sg13g2_nand2_1 _19552_ (.Y(_10457_),
    .A(_10455_),
    .B(_10456_));
 sg13g2_nor2_1 _19553_ (.A(_09383_),
    .B(_10144_),
    .Y(_10458_));
 sg13g2_nor4_1 _19554_ (.A(_09307_),
    .B(_09431_),
    .C(_09276_),
    .D(_10458_),
    .Y(_10459_));
 sg13g2_nor3_1 _19555_ (.A(_08273_),
    .B(_08269_),
    .C(_10171_),
    .Y(_10460_));
 sg13g2_nand2_1 _19556_ (.Y(_10461_),
    .A(_07179_),
    .B(_07190_));
 sg13g2_and3_1 _19557_ (.X(_10462_),
    .A(_10460_),
    .B(_10461_),
    .C(_09418_));
 sg13g2_nand3_1 _19558_ (.B(_10459_),
    .C(_10462_),
    .A(_10446_),
    .Y(_10463_));
 sg13g2_nor3_1 _19559_ (.A(_10432_),
    .B(_10463_),
    .C(_10436_),
    .Y(_10464_));
 sg13g2_nor4_1 _19560_ (.A(_09533_),
    .B(_09223_),
    .C(_09384_),
    .D(_09381_),
    .Y(_10465_));
 sg13g2_nor2_1 _19561_ (.A(_07191_),
    .B(_07179_),
    .Y(_10466_));
 sg13g2_nor2_1 _19562_ (.A(_08250_),
    .B(_10122_),
    .Y(_10467_));
 sg13g2_nand2b_1 _19563_ (.Y(_10468_),
    .B(_10467_),
    .A_N(_08265_));
 sg13g2_nor3_1 _19564_ (.A(_10466_),
    .B(_09396_),
    .C(_10468_),
    .Y(_10469_));
 sg13g2_nand3_1 _19565_ (.B(_10465_),
    .C(_10469_),
    .A(_10449_),
    .Y(_10470_));
 sg13g2_a21oi_1 _19566_ (.A1(_09342_),
    .A2(net43),
    .Y(_10471_),
    .B1(_04956_));
 sg13g2_nor2b_1 _19567_ (.A(_10471_),
    .B_N(_10435_),
    .Y(_10472_));
 sg13g2_nor3_1 _19568_ (.A(_10439_),
    .B(_10470_),
    .C(_10472_),
    .Y(_10473_));
 sg13g2_nand2_1 _19569_ (.Y(_10474_),
    .A(_10464_),
    .B(_10473_));
 sg13g2_nor2_1 _19570_ (.A(_04261_),
    .B(_05602_),
    .Y(_10475_));
 sg13g2_nand2_1 _19571_ (.Y(_10476_),
    .A(_10474_),
    .B(_10475_));
 sg13g2_nand2b_1 _19572_ (.Y(_10477_),
    .B(_10437_),
    .A_N(_10463_));
 sg13g2_nand2b_1 _19573_ (.Y(_10478_),
    .B(_10440_),
    .A_N(_10470_));
 sg13g2_nor2_1 _19574_ (.A(net192),
    .B(_05602_),
    .Y(_10479_));
 sg13g2_nand3_1 _19575_ (.B(_10478_),
    .C(_10479_),
    .A(_10477_),
    .Y(_10480_));
 sg13g2_buf_1 _19576_ (.A(_10480_),
    .X(_10481_));
 sg13g2_nand2_1 _19577_ (.Y(_10482_),
    .A(_10476_),
    .B(_10481_));
 sg13g2_nand2_1 _19578_ (.Y(_10483_),
    .A(_10481_),
    .B(_05701_));
 sg13g2_nand2_1 _19579_ (.Y(_10484_),
    .A(_05598_),
    .B(_05594_));
 sg13g2_nand3_1 _19580_ (.B(_10483_),
    .C(_10484_),
    .A(_10482_),
    .Y(_10485_));
 sg13g2_nand2_1 _19581_ (.Y(_10486_),
    .A(_10457_),
    .B(_10485_));
 sg13g2_buf_2 _19582_ (.A(\b.gen_square[1].sq.mask ),
    .X(_10487_));
 sg13g2_nand2_2 _19583_ (.Y(_10488_),
    .A(_10486_),
    .B(_10487_));
 sg13g2_nand2_1 _19584_ (.Y(_10489_),
    .A(_10430_),
    .B(_10488_));
 sg13g2_nand3_1 _19585_ (.B(_05602_),
    .C(_07575_),
    .A(_10450_),
    .Y(_10490_));
 sg13g2_nor2b_1 _19586_ (.A(_05608_),
    .B_N(_10490_),
    .Y(_10491_));
 sg13g2_nand2_1 _19587_ (.Y(_10492_),
    .A(_10453_),
    .B(_10491_));
 sg13g2_and4_1 _19588_ (.A(_05608_),
    .B(_10459_),
    .C(_09395_),
    .D(_10465_),
    .X(_10493_));
 sg13g2_nor3_1 _19589_ (.A(_02023_),
    .B(_05609_),
    .C(_10493_),
    .Y(_10494_));
 sg13g2_nand2_1 _19590_ (.Y(_10495_),
    .A(_10492_),
    .B(_10494_));
 sg13g2_nor2_1 _19591_ (.A(_05701_),
    .B(_05603_),
    .Y(_10496_));
 sg13g2_o21ai_1 _19592_ (.B1(_04044_),
    .Y(_10497_),
    .A1(_05607_),
    .A2(_05701_));
 sg13g2_nor2_1 _19593_ (.A(_10496_),
    .B(_10497_),
    .Y(_10498_));
 sg13g2_nor2_1 _19594_ (.A(_05593_),
    .B(_10481_),
    .Y(_10499_));
 sg13g2_a21oi_1 _19595_ (.A1(_10474_),
    .A2(_10498_),
    .Y(_10500_),
    .B1(_10499_));
 sg13g2_nand2_1 _19596_ (.Y(_10501_),
    .A(_10495_),
    .B(_10500_));
 sg13g2_nand2_1 _19597_ (.Y(_10502_),
    .A(_10501_),
    .B(_10487_));
 sg13g2_a22oi_1 _19598_ (.Y(_10503_),
    .B1(_04848_),
    .B2(_10399_),
    .A2(_04841_),
    .A1(_04044_));
 sg13g2_a21oi_1 _19599_ (.A1(_10381_),
    .A2(_10397_),
    .Y(_10504_),
    .B1(_10503_));
 sg13g2_nor2_1 _19600_ (.A(_04839_),
    .B(_10413_),
    .Y(_10505_));
 sg13g2_nor2_1 _19601_ (.A(_10504_),
    .B(_10505_),
    .Y(_10506_));
 sg13g2_nor2_1 _19602_ (.A(_04849_),
    .B(_10421_),
    .Y(_10507_));
 sg13g2_nor2_1 _19603_ (.A(_09218_),
    .B(_10507_),
    .Y(_10508_));
 sg13g2_nand2_1 _19604_ (.Y(_10509_),
    .A(_10423_),
    .B(_10508_));
 sg13g2_nor4_1 _19605_ (.A(_04853_),
    .B(_10316_),
    .C(_10352_),
    .D(_10394_),
    .Y(_10510_));
 sg13g2_nor3_1 _19606_ (.A(_02023_),
    .B(_04854_),
    .C(_10510_),
    .Y(_10511_));
 sg13g2_nand2_1 _19607_ (.Y(_10512_),
    .A(_10509_),
    .B(_10511_));
 sg13g2_nand2_1 _19608_ (.Y(_10513_),
    .A(_10506_),
    .B(_10512_));
 sg13g2_nand2_1 _19609_ (.Y(_10514_),
    .A(_10513_),
    .B(_10428_));
 sg13g2_inv_1 _19610_ (.Y(_10515_),
    .A(_10514_));
 sg13g2_nor2_1 _19611_ (.A(_10502_),
    .B(_10515_),
    .Y(_10516_));
 sg13g2_nand2_1 _19612_ (.Y(_10517_),
    .A(_10489_),
    .B(_10516_));
 sg13g2_inv_1 _19613_ (.Y(_10518_),
    .A(_10430_));
 sg13g2_nand2b_1 _19614_ (.Y(_10519_),
    .B(_10518_),
    .A_N(_10488_));
 sg13g2_nand2_1 _19615_ (.Y(_10520_),
    .A(_10517_),
    .B(_10519_));
 sg13g2_a21oi_1 _19616_ (.A1(_10348_),
    .A2(_10392_),
    .Y(_10521_),
    .B1(_09574_));
 sg13g2_nor2_1 _19617_ (.A(_10521_),
    .B(_10507_),
    .Y(_10522_));
 sg13g2_nor2b_1 _19618_ (.A(_10522_),
    .B_N(_10426_),
    .Y(_10523_));
 sg13g2_a21oi_1 _19619_ (.A1(_10425_),
    .A2(_10426_),
    .Y(_10524_),
    .B1(_10523_));
 sg13g2_xnor2_1 _19620_ (.Y(_10525_),
    .A(_04836_),
    .B(_04846_));
 sg13g2_nand2_1 _19621_ (.Y(_10526_),
    .A(_10414_),
    .B(_10525_));
 sg13g2_a21oi_1 _19622_ (.A1(_10524_),
    .A2(_10526_),
    .Y(_10527_),
    .B1(_10429_));
 sg13g2_xnor2_1 _19623_ (.Y(_10528_),
    .A(_05591_),
    .B(_05597_));
 sg13g2_inv_1 _19624_ (.Y(_10529_),
    .A(_10460_));
 sg13g2_o21ai_1 _19625_ (.B1(_09730_),
    .Y(_10530_),
    .A1(_10468_),
    .A2(_10529_));
 sg13g2_inv_1 _19626_ (.Y(_10531_),
    .A(_10456_));
 sg13g2_a21oi_1 _19627_ (.A1(_10490_),
    .A2(_10530_),
    .Y(_10532_),
    .B1(_10531_));
 sg13g2_a21oi_1 _19628_ (.A1(_10482_),
    .A2(_10528_),
    .Y(_10533_),
    .B1(_10532_));
 sg13g2_nand2_1 _19629_ (.Y(_10534_),
    .A(_10533_),
    .B(_10457_));
 sg13g2_nand2_1 _19630_ (.Y(_10535_),
    .A(_10534_),
    .B(_10487_));
 sg13g2_nand2_1 _19631_ (.Y(_10536_),
    .A(_10527_),
    .B(_10535_));
 sg13g2_nand2_1 _19632_ (.Y(_10537_),
    .A(_10520_),
    .B(_10536_));
 sg13g2_nand2_1 _19633_ (.Y(_10538_),
    .A(_10524_),
    .B(_10526_));
 sg13g2_nand2_1 _19634_ (.Y(_10539_),
    .A(_10538_),
    .B(_10428_));
 sg13g2_inv_1 _19635_ (.Y(_10540_),
    .A(_10487_));
 sg13g2_a21oi_1 _19636_ (.A1(_10533_),
    .A2(_10457_),
    .Y(_10541_),
    .B1(_10540_));
 sg13g2_nand2_2 _19637_ (.Y(_10542_),
    .A(_10539_),
    .B(_10541_));
 sg13g2_nand3_1 _19638_ (.B(_10518_),
    .C(_10542_),
    .A(_10537_),
    .Y(_10543_));
 sg13g2_nand2_1 _19639_ (.Y(_10544_),
    .A(_10536_),
    .B(_10542_));
 sg13g2_inv_1 _19640_ (.Y(_10545_),
    .A(_10516_));
 sg13g2_nor2b_1 _19641_ (.A(_10544_),
    .B_N(_10545_),
    .Y(_10546_));
 sg13g2_xor2_1 _19642_ (.B(_10430_),
    .A(_10488_),
    .X(_10547_));
 sg13g2_nand2_1 _19643_ (.Y(_10548_),
    .A(_10546_),
    .B(_10547_));
 sg13g2_nor2b_1 _19644_ (.A(_10489_),
    .B_N(_10542_),
    .Y(_10549_));
 sg13g2_nor2b_1 _19645_ (.A(_10549_),
    .B_N(_10536_),
    .Y(_10550_));
 sg13g2_nand3_1 _19646_ (.B(_10488_),
    .C(_10550_),
    .A(_10548_),
    .Y(_10551_));
 sg13g2_nand2_1 _19647_ (.Y(_10552_),
    .A(_10543_),
    .B(_10551_));
 sg13g2_xnor2_1 _19648_ (.Y(_10553_),
    .A(_10346_),
    .B(_10552_));
 sg13g2_nand3_1 _19649_ (.B(_10542_),
    .C(_10515_),
    .A(_10537_),
    .Y(_10554_));
 sg13g2_inv_1 _19650_ (.Y(_10555_),
    .A(_10502_));
 sg13g2_nand3_1 _19651_ (.B(_10555_),
    .C(_10550_),
    .A(_10548_),
    .Y(_10556_));
 sg13g2_nand2_1 _19652_ (.Y(_10557_),
    .A(_10554_),
    .B(_10556_));
 sg13g2_nand3_1 _19653_ (.B(_06338_),
    .C(_08652_),
    .A(_10339_),
    .Y(_10558_));
 sg13g2_nand3_1 _19654_ (.B(_06342_),
    .C(_10558_),
    .A(_10342_),
    .Y(_10559_));
 sg13g2_inv_1 _19655_ (.Y(_10560_),
    .A(_09859_));
 sg13g2_nor2_1 _19656_ (.A(_06342_),
    .B(_10270_),
    .Y(_10561_));
 sg13g2_nand4_1 _19657_ (.B(_10560_),
    .C(_10274_),
    .A(_10321_),
    .Y(_10562_),
    .D(_10561_));
 sg13g2_nor2_1 _19658_ (.A(net154),
    .B(_06343_),
    .Y(_10563_));
 sg13g2_nand3_1 _19659_ (.B(_10562_),
    .C(_10563_),
    .A(_10559_),
    .Y(_10564_));
 sg13g2_nor2_1 _19660_ (.A(_06339_),
    .B(_10332_),
    .Y(_10565_));
 sg13g2_nand2_1 _19661_ (.Y(_10566_),
    .A(_06418_),
    .B(_06335_));
 sg13g2_nand3_1 _19662_ (.B(_05082_),
    .C(_10566_),
    .A(_10335_),
    .Y(_10567_));
 sg13g2_a21oi_1 _19663_ (.A1(_06339_),
    .A2(_06418_),
    .Y(_10568_),
    .B1(_10567_));
 sg13g2_nor2_1 _19664_ (.A(_10565_),
    .B(_10568_),
    .Y(_10569_));
 sg13g2_inv_1 _19665_ (.Y(_10570_),
    .A(\b.gen_square[2].sq.mask ));
 sg13g2_a21o_1 _19666_ (.A2(_10569_),
    .A1(_10564_),
    .B1(_10570_),
    .X(_10571_));
 sg13g2_buf_1 _19667_ (.A(_10571_),
    .X(_10572_));
 sg13g2_nor2_1 _19668_ (.A(_10541_),
    .B(_10527_),
    .Y(_10573_));
 sg13g2_nand2_1 _19669_ (.Y(_10574_),
    .A(_10281_),
    .B(_10327_));
 sg13g2_nand2_1 _19670_ (.Y(_10575_),
    .A(_10574_),
    .B(_09213_));
 sg13g2_nand3_1 _19671_ (.B(_10558_),
    .C(_10575_),
    .A(_10343_),
    .Y(_10576_));
 sg13g2_nor2b_1 _19672_ (.A(_10576_),
    .B_N(_10342_),
    .Y(_10577_));
 sg13g2_nand2b_1 _19673_ (.Y(_10578_),
    .B(_02012_),
    .A_N(_10577_));
 sg13g2_xnor2_1 _19674_ (.Y(_10579_),
    .A(_06337_),
    .B(_06346_));
 sg13g2_nand2_1 _19675_ (.Y(_10580_),
    .A(_10337_),
    .B(_10579_));
 sg13g2_a21oi_1 _19676_ (.A1(_10578_),
    .A2(_10580_),
    .Y(_10581_),
    .B1(_10570_));
 sg13g2_xnor2_1 _19677_ (.Y(_10582_),
    .A(_10573_),
    .B(_10581_));
 sg13g2_a21oi_1 _19678_ (.A1(_10557_),
    .A2(_10572_),
    .Y(_10583_),
    .B1(_10582_));
 sg13g2_nor2_1 _19679_ (.A(_10572_),
    .B(_10557_),
    .Y(_10584_));
 sg13g2_nand3_1 _19680_ (.B(_10583_),
    .C(_10584_),
    .A(_10553_),
    .Y(_10585_));
 sg13g2_buf_1 _19681_ (.A(_10585_),
    .X(_10586_));
 sg13g2_inv_2 _19682_ (.Y(_10587_),
    .A(_10552_));
 sg13g2_nor2_1 _19683_ (.A(_10346_),
    .B(_10587_),
    .Y(_10588_));
 sg13g2_inv_2 _19684_ (.Y(_10589_),
    .A(_10582_));
 sg13g2_nand2_1 _19685_ (.Y(_10590_),
    .A(_10581_),
    .B(_10573_));
 sg13g2_inv_2 _19686_ (.Y(_10591_),
    .A(_10590_));
 sg13g2_a21oi_2 _19687_ (.B1(_10591_),
    .Y(_10592_),
    .A2(_10589_),
    .A1(_10588_));
 sg13g2_nand2_1 _19688_ (.Y(_10593_),
    .A(_10586_),
    .B(_10592_));
 sg13g2_inv_1 _19689_ (.Y(_10594_),
    .A(_10346_));
 sg13g2_nand2_1 _19690_ (.Y(_10595_),
    .A(_10593_),
    .B(_10594_));
 sg13g2_nand3_1 _19691_ (.B(_10587_),
    .C(_10592_),
    .A(_10586_),
    .Y(_10596_));
 sg13g2_nand2_1 _19692_ (.Y(_10597_),
    .A(_10595_),
    .B(_10596_));
 sg13g2_inv_1 _19693_ (.Y(_10598_),
    .A(_09836_));
 sg13g2_a21oi_1 _19694_ (.A1(_10598_),
    .A2(net65),
    .Y(_10599_),
    .B1(_07002_));
 sg13g2_a21oi_1 _19695_ (.A1(_09861_),
    .A2(net65),
    .Y(_10600_),
    .B1(_08286_));
 sg13g2_inv_1 _19696_ (.Y(_10601_),
    .A(_10600_));
 sg13g2_nor2_1 _19697_ (.A(_10599_),
    .B(_10601_),
    .Y(_10602_));
 sg13g2_inv_1 _19698_ (.Y(_10603_),
    .A(_09383_));
 sg13g2_a21oi_1 _19699_ (.A1(_10144_),
    .A2(_10603_),
    .Y(_10604_),
    .B1(_09101_));
 sg13g2_inv_1 _19700_ (.Y(_10605_),
    .A(_09381_));
 sg13g2_inv_1 _19701_ (.Y(_10606_),
    .A(_10311_));
 sg13g2_a21oi_1 _19702_ (.A1(_10606_),
    .A2(_09121_),
    .Y(_10607_),
    .B1(_09859_));
 sg13g2_and3_1 _19703_ (.X(_10608_),
    .A(_10604_),
    .B(_10605_),
    .C(_10607_));
 sg13g2_inv_1 _19704_ (.Y(_10609_),
    .A(_10608_));
 sg13g2_o21ai_1 _19705_ (.B1(_07582_),
    .Y(_10610_),
    .A1(_08901_),
    .A2(_09562_));
 sg13g2_inv_1 _19706_ (.Y(_10611_),
    .A(_10144_));
 sg13g2_nor2_1 _19707_ (.A(_10132_),
    .B(_10611_),
    .Y(_10612_));
 sg13g2_a21oi_1 _19708_ (.A1(_04510_),
    .A2(_09950_),
    .Y(_10613_),
    .B1(_05888_));
 sg13g2_nor2_2 _19709_ (.A(_05948_),
    .B(_10613_),
    .Y(_10614_));
 sg13g2_a21oi_1 _19710_ (.A1(_04510_),
    .A2(_09511_),
    .Y(_10615_),
    .B1(_04832_));
 sg13g2_nor2_1 _19711_ (.A(_04954_),
    .B(_10615_),
    .Y(_10616_));
 sg13g2_nor2_1 _19712_ (.A(_10614_),
    .B(_10616_),
    .Y(_10617_));
 sg13g2_and2_1 _19713_ (.A(_08409_),
    .B(_10617_),
    .X(_10618_));
 sg13g2_nor2b_1 _19714_ (.A(_10612_),
    .B_N(_10618_),
    .Y(_10619_));
 sg13g2_o21ai_1 _19715_ (.B1(_10619_),
    .Y(_10620_),
    .A1(_10610_),
    .A2(_09380_));
 sg13g2_a21oi_1 _19716_ (.A1(_09699_),
    .A2(_06530_),
    .Y(_10621_),
    .B1(_06560_));
 sg13g2_inv_1 _19717_ (.Y(_10622_),
    .A(_10621_));
 sg13g2_a21oi_1 _19718_ (.A1(_09706_),
    .A2(net36),
    .Y(_10623_),
    .B1(_06808_));
 sg13g2_nand2b_1 _19719_ (.Y(_10624_),
    .B(_10301_),
    .A_N(_10293_));
 sg13g2_o21ai_1 _19720_ (.B1(_10624_),
    .Y(_10625_),
    .A1(_10622_),
    .A2(_10623_));
 sg13g2_nor4_1 _19721_ (.A(_10602_),
    .B(_10609_),
    .C(_10620_),
    .D(_10625_),
    .Y(_10626_));
 sg13g2_nor2b_1 _19722_ (.A(_09378_),
    .B_N(_09380_),
    .Y(_10627_));
 sg13g2_nor2_1 _19723_ (.A(_09113_),
    .B(_10458_),
    .Y(_10628_));
 sg13g2_nand3_1 _19724_ (.B(_10318_),
    .C(_09157_),
    .A(_10628_),
    .Y(_10629_));
 sg13g2_inv_1 _19725_ (.Y(_10630_),
    .A(_10610_));
 sg13g2_a22oi_1 _19726_ (.Y(_10631_),
    .B1(_10599_),
    .B2(_10600_),
    .A2(_09380_),
    .A1(_10630_));
 sg13g2_nor2_2 _19727_ (.A(_04026_),
    .B(_10615_),
    .Y(_10632_));
 sg13g2_nor2_2 _19728_ (.A(_02939_),
    .B(_10613_),
    .Y(_10633_));
 sg13g2_nor2_1 _19729_ (.A(_10633_),
    .B(_07838_),
    .Y(_10634_));
 sg13g2_inv_1 _19730_ (.Y(_10635_),
    .A(_10634_));
 sg13g2_nor3_1 _19731_ (.A(_08269_),
    .B(_10632_),
    .C(_10635_),
    .Y(_10636_));
 sg13g2_nand2_1 _19732_ (.Y(_10637_),
    .A(_10631_),
    .B(_10636_));
 sg13g2_a22oi_1 _19733_ (.Y(_10638_),
    .B1(_10621_),
    .B2(_10623_),
    .A2(_10611_),
    .A1(_10131_));
 sg13g2_o21ai_1 _19734_ (.B1(_10638_),
    .Y(_10639_),
    .A1(_10293_),
    .A2(_10606_));
 sg13g2_nor4_1 _19735_ (.A(_10627_),
    .B(_10629_),
    .C(_10637_),
    .D(_10639_),
    .Y(_10640_));
 sg13g2_nor3_1 _19736_ (.A(_06540_),
    .B(_10626_),
    .C(_10640_),
    .Y(_10641_));
 sg13g2_nand2_1 _19737_ (.Y(_10642_),
    .A(_10641_),
    .B(_05072_));
 sg13g2_nand2_1 _19738_ (.Y(_10643_),
    .A(_10640_),
    .B(_10626_));
 sg13g2_nand3_1 _19739_ (.B(_05082_),
    .C(_06541_),
    .A(_10643_),
    .Y(_10644_));
 sg13g2_nand2_1 _19740_ (.Y(_10645_),
    .A(_10642_),
    .B(_10644_));
 sg13g2_nand2_1 _19741_ (.Y(_10646_),
    .A(_10642_),
    .B(_06799_));
 sg13g2_nand2_1 _19742_ (.Y(_10647_),
    .A(_06535_),
    .B(_06537_));
 sg13g2_nand3_1 _19743_ (.B(_10646_),
    .C(_10647_),
    .A(_10645_),
    .Y(_10648_));
 sg13g2_a21oi_1 _19744_ (.A1(_10601_),
    .A2(_10610_),
    .Y(_10649_),
    .B1(_06541_));
 sg13g2_nor3_1 _19745_ (.A(_10625_),
    .B(_10612_),
    .C(_10639_),
    .Y(_10650_));
 sg13g2_nor2_1 _19746_ (.A(_06541_),
    .B(_10650_),
    .Y(_10651_));
 sg13g2_o21ai_1 _19747_ (.B1(_06536_),
    .Y(_10652_),
    .A1(_10649_),
    .A2(_10651_));
 sg13g2_nand2_1 _19748_ (.Y(_10653_),
    .A(_10651_),
    .B(_06538_));
 sg13g2_nand2_1 _19749_ (.Y(_10654_),
    .A(_06546_),
    .B(net160));
 sg13g2_a21o_1 _19750_ (.A2(_10653_),
    .A1(_10652_),
    .B1(_10654_),
    .X(_10655_));
 sg13g2_nand2_1 _19751_ (.Y(_10656_),
    .A(_10648_),
    .B(_10655_));
 sg13g2_buf_1 _19752_ (.A(\b.gen_square[3].sq.mask ),
    .X(_10657_));
 sg13g2_nand2_1 _19753_ (.Y(_10658_),
    .A(_10656_),
    .B(_10657_));
 sg13g2_nor2b_1 _19754_ (.A(_10581_),
    .B_N(_10573_),
    .Y(_10659_));
 sg13g2_xnor2_1 _19755_ (.Y(_10660_),
    .A(_06531_),
    .B(_06534_));
 sg13g2_nand2_1 _19756_ (.Y(_10661_),
    .A(_10649_),
    .B(_08793_));
 sg13g2_a21o_1 _19757_ (.A2(_10618_),
    .A1(_10636_),
    .B1(_09126_),
    .X(_10662_));
 sg13g2_a21oi_1 _19758_ (.A1(_10661_),
    .A2(_10662_),
    .Y(_10663_),
    .B1(_10654_));
 sg13g2_a21oi_1 _19759_ (.A1(_10645_),
    .A2(_10660_),
    .Y(_10664_),
    .B1(_10663_));
 sg13g2_inv_1 _19760_ (.Y(_10665_),
    .A(_10657_));
 sg13g2_a21o_1 _19761_ (.A2(_10655_),
    .A1(_10664_),
    .B1(_10665_),
    .X(_10666_));
 sg13g2_buf_1 _19762_ (.A(_10666_),
    .X(_10667_));
 sg13g2_nor2b_1 _19763_ (.A(_10659_),
    .B_N(_10667_),
    .Y(_10668_));
 sg13g2_a21oi_1 _19764_ (.A1(_10597_),
    .A2(_10658_),
    .Y(_10669_),
    .B1(_10668_));
 sg13g2_inv_1 _19765_ (.Y(_10670_),
    .A(_10658_));
 sg13g2_nand3_1 _19766_ (.B(_10596_),
    .C(_10670_),
    .A(_10595_),
    .Y(_10671_));
 sg13g2_inv_1 _19767_ (.Y(_10672_),
    .A(_10557_));
 sg13g2_nand3_1 _19768_ (.B(_10672_),
    .C(_10592_),
    .A(_10586_),
    .Y(_10673_));
 sg13g2_nand2b_1 _19769_ (.Y(_10674_),
    .B(_10572_),
    .A_N(_10592_));
 sg13g2_nand2_1 _19770_ (.Y(_10675_),
    .A(_10673_),
    .B(_10674_));
 sg13g2_nor2_1 _19771_ (.A(_10627_),
    .B(_10629_),
    .Y(_10676_));
 sg13g2_a21oi_1 _19772_ (.A1(_10676_),
    .A2(_10608_),
    .Y(_10677_),
    .B1(_06541_));
 sg13g2_nand3_1 _19773_ (.B(_06546_),
    .C(_10661_),
    .A(_10652_),
    .Y(_10678_));
 sg13g2_o21ai_1 _19774_ (.B1(_10678_),
    .Y(_10679_),
    .A1(_06546_),
    .A2(_10677_));
 sg13g2_nor2_1 _19775_ (.A(_06533_),
    .B(_10642_),
    .Y(_10680_));
 sg13g2_nand2_1 _19776_ (.Y(_10681_),
    .A(_06800_),
    .B(_06540_));
 sg13g2_nand3_1 _19777_ (.B(_05083_),
    .C(_10681_),
    .A(_10643_),
    .Y(_10682_));
 sg13g2_a21oi_1 _19778_ (.A1(_06533_),
    .A2(_06800_),
    .Y(_10683_),
    .B1(_10682_));
 sg13g2_nor2_1 _19779_ (.A(_10680_),
    .B(_10683_),
    .Y(_10684_));
 sg13g2_o21ai_1 _19780_ (.B1(_10684_),
    .Y(_10685_),
    .A1(_02045_),
    .A2(_10679_));
 sg13g2_nand2_1 _19781_ (.Y(_10686_),
    .A(_10685_),
    .B(_10657_));
 sg13g2_inv_1 _19782_ (.Y(_10687_),
    .A(_10686_));
 sg13g2_nand2_1 _19783_ (.Y(_10688_),
    .A(_10675_),
    .B(_10687_));
 sg13g2_nand2_1 _19784_ (.Y(_10689_),
    .A(_10671_),
    .B(_10688_));
 sg13g2_nand2_1 _19785_ (.Y(_10690_),
    .A(_10669_),
    .B(_10689_));
 sg13g2_nand2b_1 _19786_ (.Y(_10691_),
    .B(_10659_),
    .A_N(_10667_));
 sg13g2_buf_8 _19787_ (.A(_10691_),
    .X(_10692_));
 sg13g2_nand2_1 _19788_ (.Y(_10693_),
    .A(_10690_),
    .B(_10692_));
 sg13g2_nand2_1 _19789_ (.Y(_10694_),
    .A(_10693_),
    .B(_10687_));
 sg13g2_inv_1 _19790_ (.Y(_10695_),
    .A(_10675_));
 sg13g2_nand3_1 _19791_ (.B(_10692_),
    .C(_10695_),
    .A(_10690_),
    .Y(_10696_));
 sg13g2_nand2_1 _19792_ (.Y(_10697_),
    .A(_10694_),
    .B(_10696_));
 sg13g2_nor2_1 _19793_ (.A(_10268_),
    .B(_10697_),
    .Y(_10698_));
 sg13g2_nand2_1 _19794_ (.Y(_10699_),
    .A(_10693_),
    .B(_10658_));
 sg13g2_inv_1 _19795_ (.Y(_10700_),
    .A(_10597_));
 sg13g2_nand3_1 _19796_ (.B(_10692_),
    .C(_10700_),
    .A(_10690_),
    .Y(_10701_));
 sg13g2_inv_1 _19797_ (.Y(_10702_),
    .A(_10250_));
 sg13g2_nand3_1 _19798_ (.B(_05083_),
    .C(_06932_),
    .A(_10702_),
    .Y(_10703_));
 sg13g2_nand2_1 _19799_ (.Y(_10704_),
    .A(_10703_),
    .B(_10264_));
 sg13g2_nand2_1 _19800_ (.Y(_10705_),
    .A(_10264_),
    .B(_06992_));
 sg13g2_nand2_1 _19801_ (.Y(_10706_),
    .A(_06928_),
    .B(_06930_));
 sg13g2_nand3_1 _19802_ (.B(_10705_),
    .C(_10706_),
    .A(_10704_),
    .Y(_10707_));
 sg13g2_nand2_1 _19803_ (.Y(_10708_),
    .A(_10255_),
    .B(_06931_));
 sg13g2_nand2_1 _19804_ (.Y(_10709_),
    .A(_10256_),
    .B(_10708_));
 sg13g2_nand3_1 _19805_ (.B(net160),
    .C(_06923_),
    .A(_10709_),
    .Y(_10710_));
 sg13g2_nand2_1 _19806_ (.Y(_10711_),
    .A(_10707_),
    .B(_10710_));
 sg13g2_nand2_1 _19807_ (.Y(_10712_),
    .A(_10711_),
    .B(_10267_));
 sg13g2_nand3_1 _19808_ (.B(_10701_),
    .C(_10712_),
    .A(_10699_),
    .Y(_10713_));
 sg13g2_nand2_1 _19809_ (.Y(_10714_),
    .A(_10698_),
    .B(_10713_));
 sg13g2_nand2_1 _19810_ (.Y(_10715_),
    .A(_10699_),
    .B(_10701_));
 sg13g2_inv_1 _19811_ (.Y(_10716_),
    .A(_10712_));
 sg13g2_nand2_1 _19812_ (.Y(_10717_),
    .A(_10218_),
    .B(_10244_));
 sg13g2_nand2_1 _19813_ (.Y(_10718_),
    .A(_10717_),
    .B(_08969_));
 sg13g2_nand2_1 _19814_ (.Y(_10719_),
    .A(_10257_),
    .B(_10718_));
 sg13g2_o21ai_1 _19815_ (.B1(_05108_),
    .Y(_10720_),
    .A1(_10719_),
    .A2(_10709_));
 sg13g2_nor2_1 _19816_ (.A(_06918_),
    .B(_06927_),
    .Y(_10721_));
 sg13g2_o21ai_1 _19817_ (.B1(_10704_),
    .Y(_10722_),
    .A1(_06929_),
    .A2(_10721_));
 sg13g2_inv_1 _19818_ (.Y(_10723_),
    .A(_10267_));
 sg13g2_a21o_1 _19819_ (.A2(_10722_),
    .A1(_10720_),
    .B1(_10723_),
    .X(_10724_));
 sg13g2_buf_1 _19820_ (.A(_10724_),
    .X(_10725_));
 sg13g2_nand2_1 _19821_ (.Y(_10726_),
    .A(_10667_),
    .B(_10659_));
 sg13g2_nor2_1 _19822_ (.A(_10725_),
    .B(_10726_),
    .Y(_10727_));
 sg13g2_a21oi_1 _19823_ (.A1(_10715_),
    .A2(_10716_),
    .Y(_10728_),
    .B1(_10727_));
 sg13g2_nand2_1 _19824_ (.Y(_10729_),
    .A(_10714_),
    .B(_10728_));
 sg13g2_nand2_1 _19825_ (.Y(_10730_),
    .A(_10726_),
    .B(_10725_));
 sg13g2_nand2_1 _19826_ (.Y(_10731_),
    .A(_10729_),
    .B(_10730_));
 sg13g2_nand2_1 _19827_ (.Y(_10732_),
    .A(_10731_),
    .B(_10697_));
 sg13g2_inv_1 _19828_ (.Y(_10733_),
    .A(_10268_));
 sg13g2_nand3_1 _19829_ (.B(_10730_),
    .C(_10733_),
    .A(_10729_),
    .Y(_10734_));
 sg13g2_nand2_1 _19830_ (.Y(_10735_),
    .A(_10732_),
    .B(_10734_));
 sg13g2_nor2_1 _19831_ (.A(_10191_),
    .B(_10735_),
    .Y(_10736_));
 sg13g2_nand2_1 _19832_ (.Y(_10737_),
    .A(_10731_),
    .B(_10715_));
 sg13g2_nand3_1 _19833_ (.B(_10712_),
    .C(_10730_),
    .A(_10729_),
    .Y(_10738_));
 sg13g2_inv_1 _19834_ (.Y(_10739_),
    .A(_10176_));
 sg13g2_nand3_1 _19835_ (.B(net144),
    .C(_07082_),
    .A(_10739_),
    .Y(_10740_));
 sg13g2_nand2_1 _19836_ (.Y(_10741_),
    .A(_10740_),
    .B(_10179_));
 sg13g2_nand2_1 _19837_ (.Y(_10742_),
    .A(_10179_),
    .B(_07130_));
 sg13g2_nand2_1 _19838_ (.Y(_10743_),
    .A(_07078_),
    .B(_07075_));
 sg13g2_nand3_1 _19839_ (.B(_10742_),
    .C(_10743_),
    .A(_10741_),
    .Y(_10744_));
 sg13g2_nand3_1 _19840_ (.B(_07073_),
    .C(_07076_),
    .A(_10182_),
    .Y(_10745_));
 sg13g2_nand2_1 _19841_ (.Y(_10746_),
    .A(_10183_),
    .B(_10745_));
 sg13g2_nand2_1 _19842_ (.Y(_10747_),
    .A(_10746_),
    .B(net128));
 sg13g2_nand2_1 _19843_ (.Y(_10748_),
    .A(_10744_),
    .B(_10747_));
 sg13g2_nand2_1 _19844_ (.Y(_10749_),
    .A(_10748_),
    .B(_10190_));
 sg13g2_nand3_1 _19845_ (.B(_10738_),
    .C(_10749_),
    .A(_10737_),
    .Y(_10750_));
 sg13g2_nand2_1 _19846_ (.Y(_10751_),
    .A(_10736_),
    .B(_10750_));
 sg13g2_nand2_1 _19847_ (.Y(_10752_),
    .A(_10737_),
    .B(_10738_));
 sg13g2_inv_1 _19848_ (.Y(_10753_),
    .A(_10749_));
 sg13g2_nor2_1 _19849_ (.A(_07072_),
    .B(_07077_),
    .Y(_10754_));
 sg13g2_o21ai_1 _19850_ (.B1(_10741_),
    .Y(_10755_),
    .A1(_07079_),
    .A2(_10754_));
 sg13g2_o21ai_1 _19851_ (.B1(_09735_),
    .Y(_10756_),
    .A1(_10173_),
    .A2(_10124_));
 sg13g2_nand2_1 _19852_ (.Y(_10757_),
    .A(_10184_),
    .B(_10756_));
 sg13g2_o21ai_1 _19853_ (.B1(net128),
    .Y(_10758_),
    .A1(_10757_),
    .A2(_10746_));
 sg13g2_inv_1 _19854_ (.Y(_10759_),
    .A(_10190_));
 sg13g2_a21o_1 _19855_ (.A2(_10758_),
    .A1(_10755_),
    .B1(_10759_),
    .X(_10760_));
 sg13g2_buf_1 _19856_ (.A(_10760_),
    .X(_10761_));
 sg13g2_nor2b_1 _19857_ (.A(_10726_),
    .B_N(_10725_),
    .Y(_10762_));
 sg13g2_inv_1 _19858_ (.Y(_10763_),
    .A(_10762_));
 sg13g2_nor2_1 _19859_ (.A(_10761_),
    .B(_10763_),
    .Y(_10764_));
 sg13g2_a21oi_1 _19860_ (.A1(_10752_),
    .A2(_10753_),
    .Y(_10765_),
    .B1(_10764_));
 sg13g2_nand2_1 _19861_ (.Y(_10766_),
    .A(_10751_),
    .B(_10765_));
 sg13g2_nand2_2 _19862_ (.Y(_10767_),
    .A(_10763_),
    .B(_10761_));
 sg13g2_nand2_2 _19863_ (.Y(_10768_),
    .A(_10766_),
    .B(_10767_));
 sg13g2_inv_1 _19864_ (.Y(_10769_),
    .A(_10735_));
 sg13g2_nand2_1 _19865_ (.Y(_10770_),
    .A(_10768_),
    .B(_10769_));
 sg13g2_nand3_1 _19866_ (.B(_10767_),
    .C(_10191_),
    .A(_10766_),
    .Y(_10771_));
 sg13g2_buf_1 _19867_ (.A(_10771_),
    .X(_10772_));
 sg13g2_inv_1 _19868_ (.Y(_10773_),
    .A(_08929_));
 sg13g2_a21oi_1 _19869_ (.A1(_10773_),
    .A2(_04253_),
    .Y(_10774_),
    .B1(_04197_));
 sg13g2_inv_1 _19870_ (.Y(_10775_),
    .A(_10774_));
 sg13g2_a21oi_1 _19871_ (.A1(_08992_),
    .A2(_04253_),
    .Y(_10776_),
    .B1(_04280_));
 sg13g2_nor2_1 _19872_ (.A(_10062_),
    .B(_10776_),
    .Y(_10777_));
 sg13g2_nand2b_1 _19873_ (.Y(_10778_),
    .B(_10325_),
    .A_N(_08669_));
 sg13g2_nor2_1 _19874_ (.A(_07902_),
    .B(_10778_),
    .Y(_10779_));
 sg13g2_nand2b_1 _19875_ (.Y(_10780_),
    .B(_03221_),
    .A_N(_06212_));
 sg13g2_nor2_1 _19876_ (.A(_10033_),
    .B(_08949_),
    .Y(_10781_));
 sg13g2_inv_1 _19877_ (.Y(_10782_),
    .A(_08978_));
 sg13g2_nand4_1 _19878_ (.B(_10780_),
    .C(_10781_),
    .A(_10779_),
    .Y(_10783_),
    .D(_10782_));
 sg13g2_a21oi_1 _19879_ (.A1(_09082_),
    .A2(_07071_),
    .Y(_10784_),
    .B1(_05899_));
 sg13g2_nor2_1 _19880_ (.A(_09857_),
    .B(_10784_),
    .Y(_10785_));
 sg13g2_inv_1 _19881_ (.Y(_10786_),
    .A(_09144_));
 sg13g2_a21oi_1 _19882_ (.A1(_10786_),
    .A2(_07071_),
    .Y(_10787_),
    .B1(_05950_));
 sg13g2_nor2b_1 _19883_ (.A(_10785_),
    .B_N(_10787_),
    .Y(_10788_));
 sg13g2_o21ai_1 _19884_ (.B1(_10199_),
    .Y(_10789_),
    .A1(_07134_),
    .A2(_10137_));
 sg13g2_buf_1 _19885_ (.A(_10789_),
    .X(_10790_));
 sg13g2_a21oi_1 _19886_ (.A1(_10161_),
    .A2(_07133_),
    .Y(_10791_),
    .B1(_09014_));
 sg13g2_a21oi_1 _19887_ (.A1(_10790_),
    .A2(_08985_),
    .Y(_10792_),
    .B1(_10791_));
 sg13g2_nor3_1 _19888_ (.A(_10783_),
    .B(_10788_),
    .C(_10792_),
    .Y(_10793_));
 sg13g2_o21ai_1 _19889_ (.B1(_10793_),
    .Y(_10794_),
    .A1(_10775_),
    .A2(_10777_));
 sg13g2_nand2_1 _19890_ (.Y(_10795_),
    .A(_10790_),
    .B(_08985_));
 sg13g2_inv_1 _19891_ (.Y(_10796_),
    .A(_10777_));
 sg13g2_nor2_1 _19892_ (.A(_03221_),
    .B(_06212_),
    .Y(_10797_));
 sg13g2_nor3_1 _19893_ (.A(_08676_),
    .B(_10277_),
    .C(_07936_),
    .Y(_10798_));
 sg13g2_nand2b_1 _19894_ (.Y(_10799_),
    .B(_10798_),
    .A_N(_10043_));
 sg13g2_nor4_1 _19895_ (.A(_10797_),
    .B(_08997_),
    .C(_09018_),
    .D(_10799_),
    .Y(_10800_));
 sg13g2_o21ai_1 _19896_ (.B1(_10800_),
    .Y(_10801_),
    .A1(_10787_),
    .A2(_10785_));
 sg13g2_a221oi_1 _19897_ (.B2(_10775_),
    .C1(_10801_),
    .B1(_10796_),
    .A1(_10791_),
    .Y(_10802_),
    .A2(_10795_));
 sg13g2_nand2b_1 _19898_ (.Y(_10803_),
    .B(_10802_),
    .A_N(_10794_));
 sg13g2_nand2_1 _19899_ (.Y(_10804_),
    .A(_04162_),
    .B(_04167_));
 sg13g2_a21oi_1 _19900_ (.A1(_04162_),
    .A2(_04159_),
    .Y(_10805_),
    .B1(net158));
 sg13g2_nand3_1 _19901_ (.B(_10804_),
    .C(_10805_),
    .A(_10803_),
    .Y(_10806_));
 sg13g2_nand2_1 _19902_ (.Y(_10807_),
    .A(_10790_),
    .B(_07509_));
 sg13g2_o21ai_1 _19903_ (.B1(_04167_),
    .Y(_10808_),
    .A1(_10807_),
    .A2(_10776_));
 sg13g2_inv_1 _19904_ (.Y(_10809_),
    .A(_10784_));
 sg13g2_a21oi_1 _19905_ (.A1(_10809_),
    .A2(_06212_),
    .Y(_10810_),
    .B1(_05865_));
 sg13g2_inv_1 _19906_ (.Y(_10811_),
    .A(_10810_));
 sg13g2_a21o_1 _19907_ (.A2(_10811_),
    .A1(_10808_),
    .B1(_04266_),
    .X(_10812_));
 sg13g2_nand3_1 _19908_ (.B(_04157_),
    .C(_05868_),
    .A(_10810_),
    .Y(_10813_));
 sg13g2_nand3_1 _19909_ (.B(_04165_),
    .C(_10813_),
    .A(_10812_),
    .Y(_10814_));
 sg13g2_nand4_1 _19910_ (.B(_08977_),
    .C(_09109_),
    .A(_08985_),
    .Y(_10815_),
    .D(_08948_));
 sg13g2_nor3_1 _19911_ (.A(_04165_),
    .B(_09857_),
    .C(_10815_),
    .Y(_10816_));
 sg13g2_nor3_1 _19912_ (.A(net103),
    .B(_04168_),
    .C(_10816_),
    .Y(_10817_));
 sg13g2_nand2_1 _19913_ (.Y(_10818_),
    .A(_10814_),
    .B(_10817_));
 sg13g2_nand2_1 _19914_ (.Y(_10819_),
    .A(_10806_),
    .B(_10818_));
 sg13g2_nor2_1 _19915_ (.A(_04167_),
    .B(_10802_),
    .Y(_10820_));
 sg13g2_nand3_1 _19916_ (.B(_05074_),
    .C(_10794_),
    .A(_10820_),
    .Y(_10821_));
 sg13g2_buf_1 _19917_ (.A(_10821_),
    .X(_10822_));
 sg13g2_nor2_1 _19918_ (.A(_04159_),
    .B(_10822_),
    .Y(_10823_));
 sg13g2_buf_1 _19919_ (.A(\b.gen_square[6].sq.mask ),
    .X(_10824_));
 sg13g2_o21ai_1 _19920_ (.B1(_10824_),
    .Y(_10825_),
    .A1(_10819_),
    .A2(_10823_));
 sg13g2_nand3_1 _19921_ (.B(_10772_),
    .C(_10825_),
    .A(_10770_),
    .Y(_10826_));
 sg13g2_nor2_1 _19922_ (.A(_04156_),
    .B(_04265_),
    .Y(_10827_));
 sg13g2_nand3_1 _19923_ (.B(net113),
    .C(_05865_),
    .A(_10803_),
    .Y(_10828_));
 sg13g2_nand2_1 _19924_ (.Y(_10829_),
    .A(_10822_),
    .B(_10828_));
 sg13g2_o21ai_1 _19925_ (.B1(_10829_),
    .Y(_10830_),
    .A1(_05869_),
    .A2(_10827_));
 sg13g2_a21o_1 _19926_ (.A2(_10798_),
    .A1(_10779_),
    .B1(_09843_),
    .X(_10831_));
 sg13g2_nand2_1 _19927_ (.Y(_10832_),
    .A(_10813_),
    .B(_10831_));
 sg13g2_nand3_1 _19928_ (.B(_05111_),
    .C(_04165_),
    .A(_10832_),
    .Y(_10833_));
 sg13g2_o21ai_1 _19929_ (.B1(_10812_),
    .Y(_10834_),
    .A1(_04264_),
    .A2(_10808_));
 sg13g2_nand2_1 _19930_ (.Y(_10835_),
    .A(_10834_),
    .B(_05111_));
 sg13g2_nand3_1 _19931_ (.B(_10833_),
    .C(_10835_),
    .A(_10830_),
    .Y(_10836_));
 sg13g2_nand2_1 _19932_ (.Y(_10837_),
    .A(_10836_),
    .B(_10824_));
 sg13g2_inv_1 _19933_ (.Y(_10838_),
    .A(_10837_));
 sg13g2_nand2_1 _19934_ (.Y(_10839_),
    .A(_10762_),
    .B(_10761_));
 sg13g2_xnor2_1 _19935_ (.Y(_10840_),
    .A(_10838_),
    .B(_10839_));
 sg13g2_nand2_1 _19936_ (.Y(_10841_),
    .A(_10826_),
    .B(_10840_));
 sg13g2_nand2b_1 _19937_ (.Y(_10842_),
    .B(_10768_),
    .A_N(_10752_));
 sg13g2_nand3_1 _19938_ (.B(_10767_),
    .C(_10753_),
    .A(_10766_),
    .Y(_10843_));
 sg13g2_nand2_1 _19939_ (.Y(_10844_),
    .A(_10822_),
    .B(_04161_));
 sg13g2_nand2b_1 _19940_ (.Y(_10845_),
    .B(_04160_),
    .A_N(_04265_));
 sg13g2_nand3_1 _19941_ (.B(_10844_),
    .C(_10845_),
    .A(_10829_),
    .Y(_10846_));
 sg13g2_nand2_1 _19942_ (.Y(_10847_),
    .A(_10846_),
    .B(_10835_));
 sg13g2_nand2_1 _19943_ (.Y(_10848_),
    .A(_10847_),
    .B(_10824_));
 sg13g2_inv_1 _19944_ (.Y(_10849_),
    .A(_10848_));
 sg13g2_nand3_1 _19945_ (.B(_10843_),
    .C(_10849_),
    .A(_10842_),
    .Y(_10850_));
 sg13g2_nand2_1 _19946_ (.Y(_10851_),
    .A(_10768_),
    .B(_10752_));
 sg13g2_nand3_1 _19947_ (.B(_10767_),
    .C(_10749_),
    .A(_10766_),
    .Y(_10852_));
 sg13g2_nand3_1 _19948_ (.B(_10852_),
    .C(_10848_),
    .A(_10851_),
    .Y(_10853_));
 sg13g2_nand2_1 _19949_ (.Y(_10854_),
    .A(_10850_),
    .B(_10853_));
 sg13g2_nor2_1 _19950_ (.A(_10841_),
    .B(_10854_),
    .Y(_10855_));
 sg13g2_a21oi_1 _19951_ (.A1(_10770_),
    .A2(_10772_),
    .Y(_10856_),
    .B1(_10825_));
 sg13g2_nand2_1 _19952_ (.Y(_10857_),
    .A(_10855_),
    .B(_10856_));
 sg13g2_nand2_1 _19953_ (.Y(_10858_),
    .A(_10770_),
    .B(_10772_));
 sg13g2_nor2_1 _19954_ (.A(_10837_),
    .B(_10839_),
    .Y(_10859_));
 sg13g2_nor2b_1 _19955_ (.A(_10850_),
    .B_N(_10840_),
    .Y(_10860_));
 sg13g2_nor2_1 _19956_ (.A(_10859_),
    .B(_10860_),
    .Y(_10861_));
 sg13g2_nand3_1 _19957_ (.B(_10858_),
    .C(_10861_),
    .A(_10857_),
    .Y(_10862_));
 sg13g2_o21ai_1 _19958_ (.B1(_10825_),
    .Y(_10863_),
    .A1(_10859_),
    .A2(_10860_));
 sg13g2_nand2_1 _19959_ (.Y(_10864_),
    .A(_10862_),
    .B(_10863_));
 sg13g2_nand2_1 _19960_ (.Y(_10865_),
    .A(_10857_),
    .B(_10861_));
 sg13g2_nand2_1 _19961_ (.Y(_10866_),
    .A(_10865_),
    .B(_10848_));
 sg13g2_nand2_1 _19962_ (.Y(_10867_),
    .A(_10842_),
    .B(_10843_));
 sg13g2_inv_1 _19963_ (.Y(_10868_),
    .A(_10867_));
 sg13g2_nand3_1 _19964_ (.B(_10868_),
    .C(_10861_),
    .A(_10857_),
    .Y(_10869_));
 sg13g2_nand2_1 _19965_ (.Y(_10870_),
    .A(_10866_),
    .B(_10869_));
 sg13g2_o21ai_1 _19966_ (.B1(_06167_),
    .Y(_10871_),
    .A1(_06165_),
    .A2(_10014_));
 sg13g2_inv_1 _19967_ (.Y(_10872_),
    .A(_10871_));
 sg13g2_a21oi_1 _19968_ (.A1(_10010_),
    .A2(_07505_),
    .Y(_10873_),
    .B1(_07515_));
 sg13g2_inv_1 _19969_ (.Y(_10874_),
    .A(_10151_));
 sg13g2_a21oi_1 _19970_ (.A1(_10790_),
    .A2(_04173_),
    .Y(_10875_),
    .B1(_10874_));
 sg13g2_inv_1 _19971_ (.Y(_10876_),
    .A(_10154_));
 sg13g2_a21oi_1 _19972_ (.A1(_10791_),
    .A2(_04173_),
    .Y(_10877_),
    .B1(_10876_));
 sg13g2_inv_1 _19973_ (.Y(_10878_),
    .A(_10877_));
 sg13g2_a22oi_1 _19974_ (.Y(_10879_),
    .B1(_10875_),
    .B2(_10878_),
    .A2(_10873_),
    .A1(_10872_));
 sg13g2_a22oi_1 _19975_ (.Y(_10880_),
    .B1(_10877_),
    .B2(_10875_),
    .A2(_10871_),
    .A1(_10873_));
 sg13g2_inv_2 _19976_ (.Y(_10881_),
    .A(_05302_));
 sg13g2_a21oi_1 _19977_ (.A1(_10879_),
    .A2(_10880_),
    .Y(_10882_),
    .B1(_10881_));
 sg13g2_a21oi_1 _19978_ (.A1(_08957_),
    .A2(net81),
    .Y(_10883_),
    .B1(_05317_));
 sg13g2_nand2_1 _19979_ (.Y(_10884_),
    .A(_10883_),
    .B(_05302_));
 sg13g2_nand2b_1 _19980_ (.Y(_10885_),
    .B(_10884_),
    .A_N(_10882_));
 sg13g2_nand2_1 _19981_ (.Y(_10886_),
    .A(_10885_),
    .B(_05299_));
 sg13g2_nand3_1 _19982_ (.B(_05296_),
    .C(_07506_),
    .A(_10882_),
    .Y(_10887_));
 sg13g2_a21oi_1 _19983_ (.A1(_10886_),
    .A2(_10887_),
    .Y(_10888_),
    .B1(net93));
 sg13g2_a21oi_1 _19984_ (.A1(_09005_),
    .A2(net81),
    .Y(_10889_),
    .B1(_04197_));
 sg13g2_nand2_1 _19985_ (.Y(_10890_),
    .A(_10889_),
    .B(_10883_));
 sg13g2_nor2_1 _19986_ (.A(_07837_),
    .B(_10633_),
    .Y(_10891_));
 sg13g2_inv_1 _19987_ (.Y(_10892_),
    .A(_09114_));
 sg13g2_nand2b_1 _19988_ (.Y(_10893_),
    .B(_07490_),
    .A_N(_08948_));
 sg13g2_nand2_1 _19989_ (.Y(_10894_),
    .A(_10892_),
    .B(_10893_));
 sg13g2_nor2_1 _19990_ (.A(_10166_),
    .B(_10894_),
    .Y(_10895_));
 sg13g2_nand4_1 _19991_ (.B(_10890_),
    .C(_10891_),
    .A(_10880_),
    .Y(_10896_),
    .D(_10895_));
 sg13g2_nor2_1 _19992_ (.A(_08948_),
    .B(_07490_),
    .Y(_10897_));
 sg13g2_a221oi_1 _19993_ (.B2(_08980_),
    .C1(_10897_),
    .B1(_10878_),
    .A1(_05524_),
    .Y(_10898_),
    .A2(_10062_));
 sg13g2_nor2b_1 _19994_ (.A(_10889_),
    .B_N(_10883_),
    .Y(_10899_));
 sg13g2_nor2_1 _19995_ (.A(_07747_),
    .B(_10614_),
    .Y(_10900_));
 sg13g2_nor2b_1 _19996_ (.A(_10899_),
    .B_N(_10900_),
    .Y(_10901_));
 sg13g2_and3_1 _19997_ (.X(_10902_),
    .A(_10898_),
    .B(_10879_),
    .C(_10901_));
 sg13g2_nor2b_1 _19998_ (.A(_10896_),
    .B_N(_10902_),
    .Y(_10903_));
 sg13g2_inv_1 _19999_ (.Y(_10904_),
    .A(_10903_));
 sg13g2_nor2_1 _20000_ (.A(_07381_),
    .B(_05302_),
    .Y(_10905_));
 sg13g2_nand3b_1 _20001_ (.B(_10881_),
    .C(_10896_),
    .Y(_10906_),
    .A_N(_10902_));
 sg13g2_nor2_1 _20002_ (.A(_04046_),
    .B(_10906_),
    .Y(_10907_));
 sg13g2_a21o_1 _20003_ (.A2(_10905_),
    .A1(_10904_),
    .B1(_10907_),
    .X(_10908_));
 sg13g2_o21ai_1 _20004_ (.B1(_05518_),
    .Y(_10909_),
    .A1(_04046_),
    .A2(_10906_));
 sg13g2_nand2_1 _20005_ (.Y(_10910_),
    .A(_05298_),
    .B(_05517_));
 sg13g2_nand3_1 _20006_ (.B(_10909_),
    .C(_10910_),
    .A(_10908_),
    .Y(_10911_));
 sg13g2_nand2b_1 _20007_ (.Y(_10912_),
    .B(_10911_),
    .A_N(_10888_));
 sg13g2_buf_1 _20008_ (.A(\b.gen_square[7].sq.mask ),
    .X(_10913_));
 sg13g2_nand2_1 _20009_ (.Y(_10914_),
    .A(_10912_),
    .B(_10913_));
 sg13g2_inv_1 _20010_ (.Y(_10915_),
    .A(_10914_));
 sg13g2_nor2b_1 _20011_ (.A(_10884_),
    .B_N(_05295_),
    .Y(_10916_));
 sg13g2_a21oi_1 _20012_ (.A1(_10885_),
    .A2(_05299_),
    .Y(_10917_),
    .B1(_10916_));
 sg13g2_a21o_1 _20013_ (.A2(_10900_),
    .A1(_10891_),
    .B1(_09135_),
    .X(_10918_));
 sg13g2_and3_1 _20014_ (.X(_10919_),
    .A(_10917_),
    .B(_10918_),
    .C(_10887_));
 sg13g2_nor2_1 _20015_ (.A(_05291_),
    .B(_05297_),
    .Y(_10920_));
 sg13g2_o21ai_1 _20016_ (.B1(_10908_),
    .Y(_10921_),
    .A1(_05299_),
    .A2(_10920_));
 sg13g2_o21ai_1 _20017_ (.B1(_10921_),
    .Y(_10922_),
    .A1(net83),
    .A2(_10919_));
 sg13g2_nand2_1 _20018_ (.Y(_10923_),
    .A(_10922_),
    .B(_10913_));
 sg13g2_nor2_1 _20019_ (.A(_10838_),
    .B(_10839_),
    .Y(_10924_));
 sg13g2_inv_1 _20020_ (.Y(_10925_),
    .A(_10924_));
 sg13g2_nor2_1 _20021_ (.A(_10923_),
    .B(_10925_),
    .Y(_10926_));
 sg13g2_a21oi_1 _20022_ (.A1(_10870_),
    .A2(_10915_),
    .Y(_10927_),
    .B1(_10926_));
 sg13g2_inv_1 _20023_ (.Y(_10928_),
    .A(_10913_));
 sg13g2_nand2_1 _20024_ (.Y(_10929_),
    .A(_10898_),
    .B(_10895_));
 sg13g2_a21oi_1 _20025_ (.A1(_10929_),
    .A2(_05302_),
    .Y(_10930_),
    .B1(_05305_));
 sg13g2_a21oi_1 _20026_ (.A1(_10917_),
    .A2(_05305_),
    .Y(_10931_),
    .B1(_10930_));
 sg13g2_a22oi_1 _20027_ (.Y(_10932_),
    .B1(_09133_),
    .B2(_10905_),
    .A2(_05518_),
    .A1(net96));
 sg13g2_nor2_1 _20028_ (.A(_10932_),
    .B(_10903_),
    .Y(_10933_));
 sg13g2_a221oi_1 _20029_ (.B2(_09133_),
    .C1(_10933_),
    .B1(_10907_),
    .A1(_10931_),
    .Y(_10934_),
    .A2(_05113_));
 sg13g2_nor2_1 _20030_ (.A(_10928_),
    .B(_10934_),
    .Y(_10935_));
 sg13g2_inv_1 _20031_ (.Y(_10936_),
    .A(_10935_));
 sg13g2_a21oi_1 _20032_ (.A1(_10862_),
    .A2(_10863_),
    .Y(_10937_),
    .B1(_10936_));
 sg13g2_nand3_1 _20033_ (.B(_10869_),
    .C(_10914_),
    .A(_10866_),
    .Y(_10938_));
 sg13g2_nand2_1 _20034_ (.Y(_10939_),
    .A(_10937_),
    .B(_10938_));
 sg13g2_nand2_1 _20035_ (.Y(_10940_),
    .A(_10927_),
    .B(_10939_));
 sg13g2_nand2_1 _20036_ (.Y(_10941_),
    .A(_10925_),
    .B(_10923_));
 sg13g2_nand2_1 _20037_ (.Y(_10942_),
    .A(_10940_),
    .B(_10941_));
 sg13g2_buf_8 _20038_ (.A(_10942_),
    .X(_10943_));
 sg13g2_nand2b_1 _20039_ (.Y(_10944_),
    .B(_10943_),
    .A_N(_10864_));
 sg13g2_nand3_1 _20040_ (.B(_10941_),
    .C(_10935_),
    .A(_10940_),
    .Y(_10945_));
 sg13g2_nand2_1 _20041_ (.Y(_10946_),
    .A(_10944_),
    .B(_10945_));
 sg13g2_nor2_1 _20042_ (.A(_10105_),
    .B(_10946_),
    .Y(_10947_));
 sg13g2_nand2b_1 _20043_ (.Y(_10948_),
    .B(_10943_),
    .A_N(_10870_));
 sg13g2_nand3_1 _20044_ (.B(_10941_),
    .C(_10915_),
    .A(_10940_),
    .Y(_10949_));
 sg13g2_nand2_1 _20045_ (.Y(_10950_),
    .A(_10948_),
    .B(_10949_));
 sg13g2_nand2_1 _20046_ (.Y(_10951_),
    .A(_10102_),
    .B(_10085_));
 sg13g2_nand3_1 _20047_ (.B(_10100_),
    .C(_10082_),
    .A(_10099_),
    .Y(_10952_));
 sg13g2_nand2_1 _20048_ (.Y(_10953_),
    .A(_10951_),
    .B(_10952_));
 sg13g2_nand2_1 _20049_ (.Y(_10954_),
    .A(_10950_),
    .B(_10953_));
 sg13g2_nand2_1 _20050_ (.Y(_10955_),
    .A(_10947_),
    .B(_10954_));
 sg13g2_nand2_1 _20051_ (.Y(_10956_),
    .A(_10943_),
    .B(_10870_));
 sg13g2_nand3_1 _20052_ (.B(_10941_),
    .C(_10914_),
    .A(_10940_),
    .Y(_10957_));
 sg13g2_nand2_1 _20053_ (.Y(_10958_),
    .A(_10956_),
    .B(_10957_));
 sg13g2_nand2b_1 _20054_ (.Y(_10959_),
    .B(_10102_),
    .A_N(_10085_));
 sg13g2_nand3_1 _20055_ (.B(_10100_),
    .C(_10086_),
    .A(_10099_),
    .Y(_10960_));
 sg13g2_nand2_1 _20056_ (.Y(_10961_),
    .A(_10959_),
    .B(_10960_));
 sg13g2_nand2_1 _20057_ (.Y(_10962_),
    .A(_10095_),
    .B(_10094_));
 sg13g2_inv_1 _20058_ (.Y(_10963_),
    .A(_10962_));
 sg13g2_nand2_1 _20059_ (.Y(_10964_),
    .A(_10924_),
    .B(_10923_));
 sg13g2_nor2_1 _20060_ (.A(_10963_),
    .B(_10964_),
    .Y(_10965_));
 sg13g2_a21oi_1 _20061_ (.A1(_10958_),
    .A2(_10961_),
    .Y(_10966_),
    .B1(_10965_));
 sg13g2_nand2_2 _20062_ (.Y(_10967_),
    .A(_10955_),
    .B(_10966_));
 sg13g2_nand2_2 _20063_ (.Y(_10968_),
    .A(_10964_),
    .B(_10963_));
 sg13g2_nand2_1 _20064_ (.Y(_10969_),
    .A(_10967_),
    .B(_10968_));
 sg13g2_buf_8 _20065_ (.A(_10969_),
    .X(_10970_));
 sg13g2_inv_1 _20066_ (.Y(_10971_),
    .A(_10946_));
 sg13g2_nand2_1 _20067_ (.Y(_10972_),
    .A(_10970_),
    .B(_10971_));
 sg13g2_nand3_1 _20068_ (.B(_10968_),
    .C(_10105_),
    .A(_10967_),
    .Y(_10973_));
 sg13g2_buf_8 _20069_ (.A(_10973_),
    .X(_10974_));
 sg13g2_a21oi_1 _20070_ (.A1(_09406_),
    .A2(_06580_),
    .Y(_10975_),
    .B1(_06812_));
 sg13g2_inv_1 _20071_ (.Y(_10976_),
    .A(_10975_));
 sg13g2_a21oi_1 _20072_ (.A1(_10976_),
    .A2(net22),
    .Y(_10977_),
    .B1(_05956_));
 sg13g2_inv_1 _20073_ (.Y(_10978_),
    .A(_10977_));
 sg13g2_a21oi_1 _20074_ (.A1(_10978_),
    .A2(net25),
    .Y(_10979_),
    .B1(_05527_));
 sg13g2_inv_1 _20075_ (.Y(_10980_),
    .A(_10979_));
 sg13g2_inv_1 _20076_ (.Y(_10981_),
    .A(_05627_));
 sg13g2_a21oi_1 _20077_ (.A1(_06037_),
    .A2(net38),
    .Y(_10982_),
    .B1(_10981_));
 sg13g2_inv_1 _20078_ (.Y(_10983_),
    .A(_10982_));
 sg13g2_a21oi_1 _20079_ (.A1(_10983_),
    .A2(net29),
    .Y(_10984_),
    .B1(_06370_));
 sg13g2_inv_1 _20080_ (.Y(_10985_),
    .A(_10984_));
 sg13g2_a21oi_1 _20081_ (.A1(_10985_),
    .A2(_06580_),
    .Y(_10986_),
    .B1(_06589_));
 sg13g2_inv_1 _20082_ (.Y(_10987_),
    .A(_10986_));
 sg13g2_a21oi_1 _20083_ (.A1(_10987_),
    .A2(net22),
    .Y(_10988_),
    .B1(_06971_));
 sg13g2_inv_1 _20084_ (.Y(_10989_),
    .A(_10988_));
 sg13g2_a21oi_1 _20085_ (.A1(_10989_),
    .A2(net25),
    .Y(_10990_),
    .B1(_07106_));
 sg13g2_a22oi_1 _20086_ (.Y(_10991_),
    .B1(_04281_),
    .B2(_04199_),
    .A2(_07522_),
    .A1(_06727_));
 sg13g2_o21ai_1 _20087_ (.B1(_10991_),
    .Y(_10992_),
    .A1(_08927_),
    .A2(_08923_));
 sg13g2_a21oi_1 _20088_ (.A1(_10980_),
    .A2(_10990_),
    .Y(_10993_),
    .B1(_10992_));
 sg13g2_inv_1 _20089_ (.Y(_10994_),
    .A(_10993_));
 sg13g2_a22oi_1 _20090_ (.Y(_10995_),
    .B1(_10990_),
    .B2(_10979_),
    .A2(_04281_),
    .A1(_04198_));
 sg13g2_a22oi_1 _20091_ (.Y(_10996_),
    .B1(_08922_),
    .B2(_08927_),
    .A2(_07522_),
    .A1(_07492_));
 sg13g2_nand2_1 _20092_ (.Y(_10997_),
    .A(_10995_),
    .B(_10996_));
 sg13g2_o21ai_1 _20093_ (.B1(net116),
    .Y(_10998_),
    .A1(_10994_),
    .A2(_10997_));
 sg13g2_nand2b_1 _20094_ (.Y(_10999_),
    .B(_08736_),
    .A_N(_10797_));
 sg13g2_a21oi_1 _20095_ (.A1(_06999_),
    .A2(net64),
    .Y(_11000_),
    .B1(_05950_));
 sg13g2_a21oi_1 _20096_ (.A1(_08160_),
    .A2(net64),
    .Y(_11001_),
    .B1(_05899_));
 sg13g2_nand2_1 _20097_ (.Y(_11002_),
    .A(_08706_),
    .B(_10780_));
 sg13g2_a221oi_1 _20098_ (.B2(_10018_),
    .C1(_11002_),
    .B1(_10025_),
    .A1(_11000_),
    .Y(_11003_),
    .A2(_11001_));
 sg13g2_inv_1 _20099_ (.Y(_11004_),
    .A(_11000_));
 sg13g2_a22oi_1 _20100_ (.Y(_11005_),
    .B1(_10018_),
    .B2(_10026_),
    .A2(_11001_),
    .A1(_11004_));
 sg13g2_nand3b_1 _20101_ (.B(_11003_),
    .C(_11005_),
    .Y(_11006_),
    .A_N(_10999_));
 sg13g2_nand2_1 _20102_ (.Y(_11007_),
    .A(_11006_),
    .B(net116));
 sg13g2_a21o_1 _20103_ (.A2(_11007_),
    .A1(_10998_),
    .B1(_04291_),
    .X(_11008_));
 sg13g2_nand3_1 _20104_ (.B(net116),
    .C(_06213_),
    .A(_11006_),
    .Y(_11009_));
 sg13g2_nand3_1 _20105_ (.B(_04209_),
    .C(_11009_),
    .A(_11008_),
    .Y(_11010_));
 sg13g2_nor4_1 _20106_ (.A(_07801_),
    .B(_08703_),
    .C(_09114_),
    .D(_09115_),
    .Y(_11011_));
 sg13g2_nor2_1 _20107_ (.A(_08934_),
    .B(_07815_),
    .Y(_11012_));
 sg13g2_nor2_1 _20108_ (.A(_10036_),
    .B(_09003_),
    .Y(_11013_));
 sg13g2_nand4_1 _20109_ (.B(_08936_),
    .C(_08944_),
    .A(_11013_),
    .Y(_11014_),
    .D(_08948_));
 sg13g2_nor2_1 _20110_ (.A(_07724_),
    .B(_07704_),
    .Y(_11015_));
 sg13g2_nor2b_1 _20111_ (.A(_11014_),
    .B_N(_11015_),
    .Y(_11016_));
 sg13g2_nor2_1 _20112_ (.A(_08737_),
    .B(_09103_),
    .Y(_11017_));
 sg13g2_nand4_1 _20113_ (.B(_11012_),
    .C(_11016_),
    .A(_11011_),
    .Y(_11018_),
    .D(_11017_));
 sg13g2_nor2_1 _20114_ (.A(net93),
    .B(_04212_),
    .Y(_11019_));
 sg13g2_nand3_1 _20115_ (.B(_11018_),
    .C(_11019_),
    .A(_11010_),
    .Y(_11020_));
 sg13g2_inv_1 _20116_ (.Y(_11021_),
    .A(_11011_));
 sg13g2_nor2_1 _20117_ (.A(_08040_),
    .B(_10324_),
    .Y(_11022_));
 sg13g2_inv_1 _20118_ (.Y(_11023_),
    .A(_11022_));
 sg13g2_nor4_1 _20119_ (.A(_09745_),
    .B(_09148_),
    .C(_11023_),
    .D(_05020_),
    .Y(_11024_));
 sg13g2_nand4_1 _20120_ (.B(_11012_),
    .C(_11024_),
    .A(_11003_),
    .Y(_11025_),
    .D(_08950_));
 sg13g2_nor3_1 _20121_ (.A(_10997_),
    .B(_11021_),
    .C(_11025_),
    .Y(_11026_));
 sg13g2_nor2_1 _20122_ (.A(_04548_),
    .B(_10277_),
    .Y(_11027_));
 sg13g2_nor2_1 _20123_ (.A(_09737_),
    .B(_08106_),
    .Y(_11028_));
 sg13g2_nor2_1 _20124_ (.A(_09138_),
    .B(_04585_),
    .Y(_11029_));
 sg13g2_and3_1 _20125_ (.X(_11030_),
    .A(_11027_),
    .B(_11028_),
    .C(_11029_));
 sg13g2_inv_1 _20126_ (.Y(_11031_),
    .A(_11030_));
 sg13g2_nor3_1 _20127_ (.A(_10999_),
    .B(_09000_),
    .C(_11031_),
    .Y(_11032_));
 sg13g2_nand4_1 _20128_ (.B(_11015_),
    .C(_11032_),
    .A(_11005_),
    .Y(_11033_),
    .D(_11013_));
 sg13g2_nor4_1 _20129_ (.A(_08737_),
    .B(_09103_),
    .C(_11033_),
    .D(_10994_),
    .Y(_11034_));
 sg13g2_nand2_1 _20130_ (.Y(_11035_),
    .A(_11026_),
    .B(_11034_));
 sg13g2_o21ai_1 _20131_ (.B1(_04206_),
    .Y(_11036_),
    .A1(_04203_),
    .A2(_04211_));
 sg13g2_nand3_1 _20132_ (.B(net86),
    .C(_11036_),
    .A(_11035_),
    .Y(_11037_));
 sg13g2_nor3_1 _20133_ (.A(net116),
    .B(_11034_),
    .C(_11026_),
    .Y(_11038_));
 sg13g2_nand2_1 _20134_ (.Y(_11039_),
    .A(_11038_),
    .B(_05076_));
 sg13g2_or2_1 _20135_ (.X(_11040_),
    .B(_11039_),
    .A(_04203_));
 sg13g2_nand3_1 _20136_ (.B(_11037_),
    .C(_11040_),
    .A(_11020_),
    .Y(_11041_));
 sg13g2_buf_1 _20137_ (.A(\b.gen_square[22].sq.mask ),
    .X(_11042_));
 sg13g2_nand2_1 _20138_ (.Y(_11043_),
    .A(_11041_),
    .B(_11042_));
 sg13g2_nor2_1 _20139_ (.A(\b.gen_square[22].sq.color ),
    .B(net62),
    .Y(_11044_));
 sg13g2_nand2_1 _20140_ (.Y(_11045_),
    .A(_06727_),
    .B(_04216_));
 sg13g2_nand2b_1 _20141_ (.Y(_11046_),
    .B(_11045_),
    .A_N(_11044_));
 sg13g2_nor2_1 _20142_ (.A(\b.gen_square[21].sq.color ),
    .B(_05289_),
    .Y(_11047_));
 sg13g2_a21oi_2 _20143_ (.B1(_11047_),
    .Y(_11048_),
    .A2(_05289_),
    .A1(_11046_));
 sg13g2_nor2_1 _20144_ (.A(_05864_),
    .B(_11048_),
    .Y(_11049_));
 sg13g2_a21oi_2 _20145_ (.B1(_11049_),
    .Y(_11050_),
    .A2(_05864_),
    .A1(_03567_));
 sg13g2_a21oi_2 _20146_ (.B1(_09548_),
    .Y(_11051_),
    .A2(net35),
    .A1(_11050_));
 sg13g2_inv_4 _20147_ (.A(_11051_),
    .Y(_11052_));
 sg13g2_inv_1 _20148_ (.Y(_11053_),
    .A(net35));
 sg13g2_a21oi_1 _20149_ (.A1(net62),
    .A2(_07521_),
    .Y(_11054_),
    .B1(_04295_));
 sg13g2_o21ai_1 _20150_ (.B1(_07105_),
    .Y(_11055_),
    .A1(_05290_),
    .A2(_11054_));
 sg13g2_buf_1 _20151_ (.A(_11055_),
    .X(_11056_));
 sg13g2_a21oi_1 _20152_ (.A1(_11056_),
    .A2(_05863_),
    .Y(_11057_),
    .B1(_06971_));
 sg13g2_o21ai_1 _20153_ (.B1(_06588_),
    .Y(_11058_),
    .A1(_11053_),
    .A2(_11057_));
 sg13g2_inv_1 _20154_ (.Y(_11059_),
    .A(_11058_));
 sg13g2_inv_1 _20155_ (.Y(_11060_),
    .A(_09586_));
 sg13g2_nand2_1 _20156_ (.Y(_11061_),
    .A(_06427_),
    .B(_06364_));
 sg13g2_o21ai_1 _20157_ (.B1(_11061_),
    .Y(_11062_),
    .A1(_09583_),
    .A2(_11060_));
 sg13g2_a221oi_1 _20158_ (.B2(_11059_),
    .C1(_11062_),
    .B1(_11052_),
    .A1(_09376_),
    .Y(_11063_),
    .A2(_10982_));
 sg13g2_nand2_1 _20159_ (.Y(_11064_),
    .A(_09404_),
    .B(_10982_));
 sg13g2_o21ai_1 _20160_ (.B1(_11064_),
    .Y(_11065_),
    .A1(_06365_),
    .A2(_06427_));
 sg13g2_a221oi_1 _20161_ (.B2(_11051_),
    .C1(_11065_),
    .B1(_11059_),
    .A1(_09583_),
    .Y(_11066_),
    .A2(_09586_));
 sg13g2_a21o_1 _20162_ (.A2(_11066_),
    .A1(_11063_),
    .B1(_04872_),
    .X(_11067_));
 sg13g2_and2_1 _20163_ (.A(_09367_),
    .B(_09369_),
    .X(_11068_));
 sg13g2_inv_1 _20164_ (.Y(_11069_),
    .A(_09360_));
 sg13g2_nor2_1 _20165_ (.A(_08168_),
    .B(_08205_),
    .Y(_11070_));
 sg13g2_a21o_1 _20166_ (.A2(_04957_),
    .A1(_04868_),
    .B1(_11070_),
    .X(_11071_));
 sg13g2_a221oi_1 _20167_ (.B2(_11069_),
    .C1(_11071_),
    .B1(_11068_),
    .A1(_09672_),
    .Y(_11072_),
    .A2(_09674_));
 sg13g2_nand2_1 _20168_ (.Y(_11073_),
    .A(_04958_),
    .B(_04868_));
 sg13g2_o21ai_1 _20169_ (.B1(_11073_),
    .Y(_11074_),
    .A1(_09675_),
    .A2(_09672_));
 sg13g2_a221oi_1 _20170_ (.B2(_11069_),
    .C1(_11074_),
    .B1(_07989_),
    .A1(_08205_),
    .Y(_11075_),
    .A2(_08167_));
 sg13g2_a21o_1 _20171_ (.A2(_11075_),
    .A1(_11072_),
    .B1(_04872_),
    .X(_11076_));
 sg13g2_a21o_1 _20172_ (.A2(_11076_),
    .A1(_11067_),
    .B1(_04870_),
    .X(_11077_));
 sg13g2_or2_1 _20173_ (.X(_11078_),
    .B(_11076_),
    .A(_04871_));
 sg13g2_nand3_1 _20174_ (.B(_04809_),
    .C(_11078_),
    .A(_11077_),
    .Y(_11079_));
 sg13g2_inv_1 _20175_ (.Y(_11080_),
    .A(_04810_));
 sg13g2_inv_1 _20176_ (.Y(_11081_),
    .A(_08072_));
 sg13g2_inv_1 _20177_ (.Y(_11082_),
    .A(_09307_));
 sg13g2_nand4_1 _20178_ (.B(_11081_),
    .C(_11082_),
    .A(_09432_),
    .Y(_11083_),
    .D(_10318_));
 sg13g2_o21ai_1 _20179_ (.B1(_08068_),
    .Y(_11084_),
    .A1(_09547_),
    .A2(_11051_));
 sg13g2_nor3_1 _20180_ (.A(_08065_),
    .B(_11083_),
    .C(_11084_),
    .Y(_11085_));
 sg13g2_nand3_1 _20181_ (.B(_08103_),
    .C(_10362_),
    .A(_10560_),
    .Y(_11086_));
 sg13g2_o21ai_1 _20182_ (.B1(_09557_),
    .Y(_11087_),
    .A1(_07965_),
    .A2(_11068_));
 sg13g2_nor3_1 _20183_ (.A(_08096_),
    .B(_11086_),
    .C(_11087_),
    .Y(_11088_));
 sg13g2_nand2_1 _20184_ (.Y(_11089_),
    .A(_10269_),
    .B(_09534_));
 sg13g2_nor2_1 _20185_ (.A(_04809_),
    .B(_11089_),
    .Y(_11090_));
 sg13g2_nand3_1 _20186_ (.B(_11088_),
    .C(_11090_),
    .A(_11085_),
    .Y(_11091_));
 sg13g2_nand4_1 _20187_ (.B(net160),
    .C(_11080_),
    .A(_11079_),
    .Y(_11092_),
    .D(_11091_));
 sg13g2_nand2_1 _20188_ (.Y(_11093_),
    .A(_10279_),
    .B(_06297_));
 sg13g2_nor2_1 _20189_ (.A(_05828_),
    .B(_08106_),
    .Y(_11094_));
 sg13g2_nand3_1 _20190_ (.B(_09732_),
    .C(_09128_),
    .A(_11094_),
    .Y(_11095_));
 sg13g2_nor4_1 _20191_ (.A(_08108_),
    .B(_10277_),
    .C(_11093_),
    .D(_11095_),
    .Y(_11096_));
 sg13g2_nor2b_1 _20192_ (.A(_11089_),
    .B_N(_11096_),
    .Y(_11097_));
 sg13g2_nand4_1 _20193_ (.B(_11075_),
    .C(_11088_),
    .A(_11066_),
    .Y(_11098_),
    .D(_11097_));
 sg13g2_inv_1 _20194_ (.Y(_11099_),
    .A(_06461_));
 sg13g2_nand2_1 _20195_ (.Y(_11100_),
    .A(_10326_),
    .B(_11099_));
 sg13g2_inv_1 _20196_ (.Y(_11101_),
    .A(_09420_));
 sg13g2_nor2_1 _20197_ (.A(_05815_),
    .B(_09747_),
    .Y(_11102_));
 sg13g2_inv_1 _20198_ (.Y(_11103_),
    .A(_11102_));
 sg13g2_nor4_1 _20199_ (.A(_11100_),
    .B(_11101_),
    .C(_11023_),
    .D(_11103_),
    .Y(_11104_));
 sg13g2_nand4_1 _20200_ (.B(_11072_),
    .C(_11104_),
    .A(_11063_),
    .Y(_11105_),
    .D(_11085_));
 sg13g2_nor2_1 _20201_ (.A(_11098_),
    .B(_11105_),
    .Y(_11106_));
 sg13g2_inv_1 _20202_ (.Y(_11107_),
    .A(_11106_));
 sg13g2_o21ai_1 _20203_ (.B1(_04804_),
    .Y(_11108_),
    .A1(_04801_),
    .A2(_04806_));
 sg13g2_nand3_1 _20204_ (.B(net161),
    .C(_11108_),
    .A(_11107_),
    .Y(_11109_));
 sg13g2_nand4_1 _20205_ (.B(net191),
    .C(_04872_),
    .A(_11105_),
    .Y(_11110_),
    .D(_11098_));
 sg13g2_buf_1 _20206_ (.A(_11110_),
    .X(_11111_));
 sg13g2_nand2b_1 _20207_ (.Y(_11112_),
    .B(_04807_),
    .A_N(_11111_));
 sg13g2_nand3_1 _20208_ (.B(_11109_),
    .C(_11112_),
    .A(_11092_),
    .Y(_11113_));
 sg13g2_buf_1 _20209_ (.A(\b.gen_square[18].sq.mask ),
    .X(_11114_));
 sg13g2_nand2_1 _20210_ (.Y(_11115_),
    .A(_11113_),
    .B(_11114_));
 sg13g2_a21oi_1 _20211_ (.A1(_11058_),
    .A2(net29),
    .Y(_11116_),
    .B1(_06370_));
 sg13g2_o21ai_1 _20212_ (.B1(_05627_),
    .Y(_11117_),
    .A1(_05590_),
    .A2(_11116_));
 sg13g2_a21oi_1 _20213_ (.A1(_11052_),
    .A2(net29),
    .Y(_11118_),
    .B1(_09373_));
 sg13g2_o21ai_1 _20214_ (.B1(_09198_),
    .Y(_11119_),
    .A1(_05590_),
    .A2(_11118_));
 sg13g2_nand2b_1 _20215_ (.Y(_11120_),
    .B(_11119_),
    .A_N(_11117_));
 sg13g2_o21ai_1 _20216_ (.B1(_11120_),
    .Y(_11121_),
    .A1(_09177_),
    .A2(_09186_));
 sg13g2_inv_1 _20217_ (.Y(_11122_),
    .A(_08016_));
 sg13g2_a21oi_1 _20218_ (.A1(_11122_),
    .A2(net28),
    .Y(_11123_),
    .B1(_05963_));
 sg13g2_inv_1 _20219_ (.Y(_11124_),
    .A(_11123_));
 sg13g2_a21oi_1 _20220_ (.A1(_11124_),
    .A2(_05647_),
    .Y(_11125_),
    .B1(_05718_));
 sg13g2_a21oi_1 _20221_ (.A1(_08120_),
    .A2(_05844_),
    .Y(_11126_),
    .B1(_06883_));
 sg13g2_inv_1 _20222_ (.Y(_11127_),
    .A(_11126_));
 sg13g2_a21oi_1 _20223_ (.A1(_11127_),
    .A2(_05647_),
    .Y(_11128_),
    .B1(_06880_));
 sg13g2_o21ai_1 _20224_ (.B1(_07923_),
    .Y(_11129_),
    .A1(_02393_),
    .A2(_10216_));
 sg13g2_nor2_1 _20225_ (.A(_11129_),
    .B(_11103_),
    .Y(_11130_));
 sg13g2_a21oi_1 _20226_ (.A1(_06423_),
    .A2(net43),
    .Y(_11131_),
    .B1(_04956_));
 sg13g2_a21oi_1 _20227_ (.A1(_08655_),
    .A2(net43),
    .Y(_11132_),
    .B1(_04867_));
 sg13g2_nand2_1 _20228_ (.Y(_11133_),
    .A(_11131_),
    .B(_11132_));
 sg13g2_nand2_1 _20229_ (.Y(_11134_),
    .A(_11130_),
    .B(_11133_));
 sg13g2_a21oi_1 _20230_ (.A1(_11125_),
    .A2(_11128_),
    .Y(_11135_),
    .B1(_11134_));
 sg13g2_o21ai_1 _20231_ (.B1(_11135_),
    .Y(_11136_),
    .A1(_06105_),
    .A2(_06012_));
 sg13g2_nand2_1 _20232_ (.Y(_11137_),
    .A(_11119_),
    .B(_09196_));
 sg13g2_nor2_1 _20233_ (.A(_10393_),
    .B(_09307_),
    .Y(_11138_));
 sg13g2_nand4_1 _20234_ (.B(_11081_),
    .C(_08230_),
    .A(_11137_),
    .Y(_11139_),
    .D(_11138_));
 sg13g2_nor3_1 _20235_ (.A(_11121_),
    .B(_11136_),
    .C(_11139_),
    .Y(_11140_));
 sg13g2_nand2b_1 _20236_ (.Y(_11141_),
    .B(_09200_),
    .A_N(_08214_));
 sg13g2_nor2_1 _20237_ (.A(_08175_),
    .B(_10347_),
    .Y(_11142_));
 sg13g2_inv_1 _20238_ (.Y(_11143_),
    .A(_11142_));
 sg13g2_nor3_1 _20239_ (.A(_05828_),
    .B(_09733_),
    .C(_11143_),
    .Y(_11144_));
 sg13g2_nand2b_1 _20240_ (.Y(_11145_),
    .B(_11132_),
    .A_N(_11131_));
 sg13g2_nand2_1 _20241_ (.Y(_11146_),
    .A(_06105_),
    .B(_06011_));
 sg13g2_nand3_1 _20242_ (.B(_11145_),
    .C(_11146_),
    .A(_11144_),
    .Y(_11147_));
 sg13g2_inv_1 _20243_ (.Y(_11148_),
    .A(_11128_));
 sg13g2_nor3_1 _20244_ (.A(_10350_),
    .B(_08102_),
    .C(_09533_),
    .Y(_11149_));
 sg13g2_o21ai_1 _20245_ (.B1(_11149_),
    .Y(_11150_),
    .A1(_11148_),
    .A2(_11125_));
 sg13g2_nand2b_1 _20246_ (.Y(_11151_),
    .B(_09177_),
    .A_N(_09186_));
 sg13g2_o21ai_1 _20247_ (.B1(_11151_),
    .Y(_11152_),
    .A1(_11117_),
    .A2(_11119_));
 sg13g2_nor4_1 _20248_ (.A(_11141_),
    .B(_11147_),
    .C(_11150_),
    .D(_11152_),
    .Y(_11153_));
 sg13g2_nand2_1 _20249_ (.Y(_11154_),
    .A(_11140_),
    .B(_11153_));
 sg13g2_nand2_1 _20250_ (.Y(_11155_),
    .A(_06019_),
    .B(_06021_));
 sg13g2_nand3_1 _20251_ (.B(net176),
    .C(_11155_),
    .A(_11154_),
    .Y(_11156_));
 sg13g2_a21oi_1 _20252_ (.A1(_06016_),
    .A2(_06019_),
    .Y(_11157_),
    .B1(_11156_));
 sg13g2_o21ai_1 _20253_ (.B1(_06021_),
    .Y(_11158_),
    .A1(_11132_),
    .A2(_11128_));
 sg13g2_nor2b_1 _20254_ (.A(_11158_),
    .B_N(_06872_),
    .Y(_11159_));
 sg13g2_nand3_1 _20255_ (.B(_06012_),
    .C(_09186_),
    .A(_11117_),
    .Y(_11160_));
 sg13g2_nand2_1 _20256_ (.Y(_11161_),
    .A(_11160_),
    .B(_06021_));
 sg13g2_nand2_1 _20257_ (.Y(_11162_),
    .A(_11161_),
    .B(_11158_));
 sg13g2_nand2_1 _20258_ (.Y(_11163_),
    .A(_11162_),
    .B(_06034_));
 sg13g2_nand3b_1 _20259_ (.B(_11163_),
    .C(_09261_),
    .Y(_11164_),
    .A_N(_11159_));
 sg13g2_nor2_1 _20260_ (.A(_11141_),
    .B(_11139_),
    .Y(_11165_));
 sg13g2_nand3_1 _20261_ (.B(_06024_),
    .C(_11149_),
    .A(_11165_),
    .Y(_11166_));
 sg13g2_nand4_1 _20262_ (.B(_11166_),
    .C(net183),
    .A(_11164_),
    .Y(_11167_),
    .D(_06025_));
 sg13g2_nor3_1 _20263_ (.A(_06021_),
    .B(_11153_),
    .C(_11140_),
    .Y(_11168_));
 sg13g2_nand3_1 _20264_ (.B(net215),
    .C(_06023_),
    .A(_11168_),
    .Y(_11169_));
 sg13g2_nand2_1 _20265_ (.Y(_11170_),
    .A(_11167_),
    .B(_11169_));
 sg13g2_buf_1 _20266_ (.A(\b.gen_square[16].sq.mask ),
    .X(_11171_));
 sg13g2_o21ai_1 _20267_ (.B1(_11171_),
    .Y(_11172_),
    .A1(_11157_),
    .A2(_11170_));
 sg13g2_nand2_1 _20268_ (.Y(_11173_),
    .A(_11168_),
    .B(net215));
 sg13g2_nand3_1 _20269_ (.B(net176),
    .C(_06022_),
    .A(_11154_),
    .Y(_11174_));
 sg13g2_nand2_1 _20270_ (.Y(_11175_),
    .A(_11173_),
    .B(_11174_));
 sg13g2_nand2_1 _20271_ (.Y(_11176_),
    .A(_11173_),
    .B(_06018_));
 sg13g2_nand2_1 _20272_ (.Y(_11177_),
    .A(_06033_),
    .B(_06017_));
 sg13g2_nand3_1 _20273_ (.B(_11176_),
    .C(_11177_),
    .A(_11175_),
    .Y(_11178_));
 sg13g2_inv_1 _20274_ (.Y(_11179_),
    .A(_06031_));
 sg13g2_o21ai_1 _20275_ (.B1(_11163_),
    .Y(_11180_),
    .A1(_11179_),
    .A2(_11161_));
 sg13g2_nand3_1 _20276_ (.B(net183),
    .C(_09261_),
    .A(_11180_),
    .Y(_11181_));
 sg13g2_nand2_1 _20277_ (.Y(_11182_),
    .A(_11178_),
    .B(_11181_));
 sg13g2_nand2_1 _20278_ (.Y(_11183_),
    .A(_11182_),
    .B(_11171_));
 sg13g2_inv_1 _20279_ (.Y(_11184_),
    .A(_11183_));
 sg13g2_a21oi_1 _20280_ (.A1(_09338_),
    .A2(_09339_),
    .Y(_11185_),
    .B1(_09346_));
 sg13g2_a221oi_1 _20281_ (.B2(_11116_),
    .C1(_11185_),
    .B1(_11118_),
    .A1(_05708_),
    .Y(_11186_),
    .A2(_05617_));
 sg13g2_nor2_1 _20282_ (.A(_08333_),
    .B(_10466_),
    .Y(_11187_));
 sg13g2_o21ai_1 _20283_ (.B1(_11187_),
    .Y(_11188_),
    .A1(_06037_),
    .A2(_06888_));
 sg13g2_nor2_1 _20284_ (.A(_09577_),
    .B(_10122_),
    .Y(_11189_));
 sg13g2_nand4_1 _20285_ (.B(_05164_),
    .C(_07759_),
    .A(_11189_),
    .Y(_11190_),
    .D(_09215_));
 sg13g2_nor4_1 _20286_ (.A(_08324_),
    .B(_09391_),
    .C(_09396_),
    .D(_09533_),
    .Y(_11191_));
 sg13g2_nand2b_1 _20287_ (.Y(_11192_),
    .B(_11191_),
    .A_N(_11190_));
 sg13g2_nand2_1 _20288_ (.Y(_11193_),
    .A(_09191_),
    .B(_09192_));
 sg13g2_nand2b_1 _20289_ (.Y(_11194_),
    .B(_11193_),
    .A_N(_08062_));
 sg13g2_nand2_1 _20290_ (.Y(_11195_),
    .A(_11194_),
    .B(_10269_));
 sg13g2_a21oi_1 _20291_ (.A1(net37),
    .A2(_08796_),
    .Y(_11196_),
    .B1(_07583_));
 sg13g2_inv_1 _20292_ (.Y(_11197_),
    .A(_11196_));
 sg13g2_nand2b_1 _20293_ (.Y(_11198_),
    .B(_09204_),
    .A_N(_09210_));
 sg13g2_o21ai_1 _20294_ (.B1(_11198_),
    .Y(_11199_),
    .A1(_09428_),
    .A2(_11197_));
 sg13g2_nor4_1 _20295_ (.A(_11188_),
    .B(_11192_),
    .C(_11195_),
    .D(_11199_),
    .Y(_11200_));
 sg13g2_nor2b_1 _20296_ (.A(_08102_),
    .B_N(_09375_),
    .Y(_11201_));
 sg13g2_nand3_1 _20297_ (.B(_11200_),
    .C(_11201_),
    .A(_11186_),
    .Y(_11202_));
 sg13g2_inv_1 _20298_ (.Y(_11203_),
    .A(_11118_));
 sg13g2_nor4_1 _20299_ (.A(_08351_),
    .B(_09419_),
    .C(_09307_),
    .D(_09431_),
    .Y(_11204_));
 sg13g2_nand3_1 _20300_ (.B(_08459_),
    .C(_11081_),
    .A(_11204_),
    .Y(_11205_));
 sg13g2_a21oi_1 _20301_ (.A1(_11203_),
    .A2(_09372_),
    .Y(_11206_),
    .B1(_11205_));
 sg13g2_nand2_1 _20302_ (.Y(_11207_),
    .A(_05707_),
    .B(_05617_));
 sg13g2_o21ai_1 _20303_ (.B1(_11207_),
    .Y(_11208_),
    .A1(_09346_),
    .A2(_09340_));
 sg13g2_a21oi_1 _20304_ (.A1(_11203_),
    .A2(_11116_),
    .Y(_11209_),
    .B1(_11208_));
 sg13g2_nand2_1 _20305_ (.Y(_11210_),
    .A(_10461_),
    .B(_08350_));
 sg13g2_nor2_1 _20306_ (.A(_11197_),
    .B(_09429_),
    .Y(_11211_));
 sg13g2_nor2_1 _20307_ (.A(_11193_),
    .B(_09210_),
    .Y(_11212_));
 sg13g2_nor3_1 _20308_ (.A(_11210_),
    .B(_11211_),
    .C(_11212_),
    .Y(_11213_));
 sg13g2_nand2_1 _20309_ (.Y(_11214_),
    .A(_06038_),
    .B(\b.gen_square[16].sq.color ));
 sg13g2_nand2b_1 _20310_ (.Y(_11215_),
    .B(_09281_),
    .A_N(_10171_));
 sg13g2_nor3_1 _20311_ (.A(_05207_),
    .B(_11215_),
    .C(_09606_),
    .Y(_11216_));
 sg13g2_and3_1 _20312_ (.X(_11217_),
    .A(_11213_),
    .B(_11214_),
    .C(_11216_));
 sg13g2_nand3_1 _20313_ (.B(_11209_),
    .C(_11217_),
    .A(_11206_),
    .Y(_11218_));
 sg13g2_nand4_1 _20314_ (.B(net215),
    .C(_05622_),
    .A(_11202_),
    .Y(_11219_),
    .D(_11218_));
 sg13g2_buf_1 _20315_ (.A(_11219_),
    .X(_11220_));
 sg13g2_a22oi_1 _20316_ (.Y(_11221_),
    .B1(_05588_),
    .B2(_11220_),
    .A2(_05619_),
    .A1(_05587_));
 sg13g2_nor2_1 _20317_ (.A(_11218_),
    .B(_11202_),
    .Y(_11222_));
 sg13g2_inv_2 _20318_ (.Y(_11223_),
    .A(_11222_));
 sg13g2_nand3_1 _20319_ (.B(net176),
    .C(_05622_),
    .A(_11223_),
    .Y(_11224_));
 sg13g2_nand2_1 _20320_ (.Y(_11225_),
    .A(_11224_),
    .B(_11220_));
 sg13g2_nand2_1 _20321_ (.Y(_11226_),
    .A(_11221_),
    .B(_11225_));
 sg13g2_nor2b_1 _20322_ (.A(_11199_),
    .B_N(_11187_),
    .Y(_11227_));
 sg13g2_a21oi_1 _20323_ (.A1(_11227_),
    .A2(_11213_),
    .Y(_11228_),
    .B1(_05622_));
 sg13g2_nor2b_1 _20324_ (.A(_06038_),
    .B_N(_11209_),
    .Y(_11229_));
 sg13g2_a21oi_1 _20325_ (.A1(_11186_),
    .A2(_11229_),
    .Y(_11230_),
    .B1(_05622_));
 sg13g2_o21ai_1 _20326_ (.B1(_05620_),
    .Y(_11231_),
    .A1(_11228_),
    .A2(_11230_));
 sg13g2_nand2_1 _20327_ (.Y(_11232_),
    .A(_11230_),
    .B(_05621_));
 sg13g2_nand2_1 _20328_ (.Y(_11233_),
    .A(_05582_),
    .B(net183));
 sg13g2_a21o_1 _20329_ (.A2(_11232_),
    .A1(_11231_),
    .B1(_11233_),
    .X(_11234_));
 sg13g2_nand2_1 _20330_ (.Y(_11235_),
    .A(_11226_),
    .B(_11234_));
 sg13g2_buf_2 _20331_ (.A(\b.gen_square[17].sq.mask ),
    .X(_11236_));
 sg13g2_nand2_1 _20332_ (.Y(_11237_),
    .A(_11235_),
    .B(_11236_));
 sg13g2_nand2_1 _20333_ (.Y(_11238_),
    .A(_11184_),
    .B(_11237_));
 sg13g2_o21ai_1 _20334_ (.B1(_05625_),
    .Y(_11239_),
    .A1(_05580_),
    .A2(_05577_));
 sg13g2_nand3_1 _20335_ (.B(net176),
    .C(_11239_),
    .A(_11223_),
    .Y(_11240_));
 sg13g2_o21ai_1 _20336_ (.B1(_11240_),
    .Y(_11241_),
    .A1(_05580_),
    .A2(_11220_));
 sg13g2_nand2_1 _20337_ (.Y(_11242_),
    .A(_11228_),
    .B(_07193_));
 sg13g2_nand3_1 _20338_ (.B(_05582_),
    .C(_11242_),
    .A(_11231_),
    .Y(_11243_));
 sg13g2_inv_1 _20339_ (.Y(_11244_),
    .A(_11191_));
 sg13g2_nor3_1 _20340_ (.A(_05582_),
    .B(_11244_),
    .C(_11195_),
    .Y(_11245_));
 sg13g2_nand3_1 _20341_ (.B(_11201_),
    .C(_11245_),
    .A(_11206_),
    .Y(_11246_));
 sg13g2_nor2_1 _20342_ (.A(_02034_),
    .B(_05583_),
    .Y(_11247_));
 sg13g2_and3_1 _20343_ (.X(_11248_),
    .A(_11243_),
    .B(_11246_),
    .C(_11247_));
 sg13g2_o21ai_1 _20344_ (.B1(_11236_),
    .Y(_11249_),
    .A1(_11241_),
    .A2(_11248_));
 sg13g2_inv_1 _20345_ (.Y(_11250_),
    .A(_11249_));
 sg13g2_nand3_1 _20346_ (.B(_11250_),
    .C(_11172_),
    .A(_11238_),
    .Y(_11251_));
 sg13g2_inv_1 _20347_ (.Y(_11252_),
    .A(_11237_));
 sg13g2_xnor2_1 _20348_ (.Y(_11253_),
    .A(_05579_),
    .B(_05618_));
 sg13g2_nand2b_1 _20349_ (.Y(_11254_),
    .B(_11216_),
    .A_N(_11190_));
 sg13g2_nand2_1 _20350_ (.Y(_11255_),
    .A(_11254_),
    .B(_08043_));
 sg13g2_a21oi_1 _20351_ (.A1(_11242_),
    .A2(_11255_),
    .Y(_11256_),
    .B1(_11233_));
 sg13g2_a21oi_1 _20352_ (.A1(_11225_),
    .A2(_11253_),
    .Y(_11257_),
    .B1(_11256_));
 sg13g2_nand2_1 _20353_ (.Y(_11258_),
    .A(_11257_),
    .B(_11234_));
 sg13g2_nand2_1 _20354_ (.Y(_11259_),
    .A(_11258_),
    .B(_11236_));
 sg13g2_nor2_1 _20355_ (.A(_06013_),
    .B(_06032_),
    .Y(_11260_));
 sg13g2_o21ai_1 _20356_ (.B1(_11175_),
    .Y(_11261_),
    .A1(_06034_),
    .A2(_11260_));
 sg13g2_a21oi_1 _20357_ (.A1(_11130_),
    .A2(_11144_),
    .Y(_11262_),
    .B1(_08247_));
 sg13g2_nor3_1 _20358_ (.A(_11159_),
    .B(_11262_),
    .C(_11180_),
    .Y(_11263_));
 sg13g2_nand3b_1 _20359_ (.B(net183),
    .C(_09261_),
    .Y(_11264_),
    .A_N(_11263_));
 sg13g2_inv_1 _20360_ (.Y(_11265_),
    .A(_11171_));
 sg13g2_a21oi_1 _20361_ (.A1(_11261_),
    .A2(_11264_),
    .Y(_11266_),
    .B1(_11265_));
 sg13g2_nor2_1 _20362_ (.A(_11259_),
    .B(_11266_),
    .Y(_11267_));
 sg13g2_a21oi_1 _20363_ (.A1(_11183_),
    .A2(_11252_),
    .Y(_11268_),
    .B1(_11267_));
 sg13g2_nand2_1 _20364_ (.Y(_11269_),
    .A(_11251_),
    .B(_11268_));
 sg13g2_nand2_1 _20365_ (.Y(_11270_),
    .A(_11266_),
    .B(_11259_));
 sg13g2_nand2_1 _20366_ (.Y(_11271_),
    .A(_11269_),
    .B(_11270_));
 sg13g2_nand2b_1 _20367_ (.Y(_11272_),
    .B(_11271_),
    .A_N(_11172_));
 sg13g2_nand3_1 _20368_ (.B(_11250_),
    .C(_11270_),
    .A(_11269_),
    .Y(_11273_));
 sg13g2_nand2_1 _20369_ (.Y(_11274_),
    .A(_11272_),
    .B(_11273_));
 sg13g2_nor2_1 _20370_ (.A(_11115_),
    .B(_11274_),
    .Y(_11275_));
 sg13g2_nand2_1 _20371_ (.Y(_11276_),
    .A(_11271_),
    .B(_11183_));
 sg13g2_nand3_1 _20372_ (.B(_11237_),
    .C(_11270_),
    .A(_11269_),
    .Y(_11277_));
 sg13g2_nand3_1 _20373_ (.B(net161),
    .C(_04872_),
    .A(_11107_),
    .Y(_11278_));
 sg13g2_nand2_1 _20374_ (.Y(_11279_),
    .A(_11278_),
    .B(_11111_));
 sg13g2_nand2_1 _20375_ (.Y(_11280_),
    .A(_11111_),
    .B(_04803_));
 sg13g2_nand2b_1 _20376_ (.Y(_11281_),
    .B(_04802_),
    .A_N(_04869_));
 sg13g2_nand3_1 _20377_ (.B(_11280_),
    .C(_11281_),
    .A(_11279_),
    .Y(_11282_));
 sg13g2_o21ai_1 _20378_ (.B1(_11077_),
    .Y(_11283_),
    .A1(_06367_),
    .A2(_11067_));
 sg13g2_nand2_1 _20379_ (.Y(_11284_),
    .A(_11283_),
    .B(net160));
 sg13g2_nand2_1 _20380_ (.Y(_11285_),
    .A(_11282_),
    .B(_11284_));
 sg13g2_nand2_1 _20381_ (.Y(_11286_),
    .A(_11285_),
    .B(_11114_));
 sg13g2_nand3_1 _20382_ (.B(_11277_),
    .C(_11286_),
    .A(_11276_),
    .Y(_11287_));
 sg13g2_nand2_1 _20383_ (.Y(_11288_),
    .A(_11275_),
    .B(_11287_));
 sg13g2_nand2_1 _20384_ (.Y(_11289_),
    .A(_11276_),
    .B(_11277_));
 sg13g2_inv_1 _20385_ (.Y(_11290_),
    .A(_11286_));
 sg13g2_nor2_1 _20386_ (.A(net137),
    .B(_04808_),
    .Y(_11291_));
 sg13g2_a21o_1 _20387_ (.A2(_11104_),
    .A1(_11096_),
    .B1(_08261_),
    .X(_11292_));
 sg13g2_nand2_1 _20388_ (.Y(_11293_),
    .A(_11078_),
    .B(_11292_));
 sg13g2_xnor2_1 _20389_ (.Y(_11294_),
    .A(_04798_),
    .B(_04869_));
 sg13g2_a22oi_1 _20390_ (.Y(_11295_),
    .B1(_11294_),
    .B2(_11279_),
    .A2(_11293_),
    .A1(_11291_));
 sg13g2_inv_1 _20391_ (.Y(_11296_),
    .A(_11114_));
 sg13g2_a21o_1 _20392_ (.A2(_11284_),
    .A1(_11295_),
    .B1(_11296_),
    .X(_11297_));
 sg13g2_buf_1 _20393_ (.A(_11297_),
    .X(_11298_));
 sg13g2_nor2b_1 _20394_ (.A(_11266_),
    .B_N(_11259_),
    .Y(_11299_));
 sg13g2_inv_1 _20395_ (.Y(_11300_),
    .A(_11299_));
 sg13g2_nor2_1 _20396_ (.A(_11298_),
    .B(_11300_),
    .Y(_11301_));
 sg13g2_a21oi_1 _20397_ (.A1(_11289_),
    .A2(_11290_),
    .Y(_11302_),
    .B1(_11301_));
 sg13g2_nand2_1 _20398_ (.Y(_11303_),
    .A(_11288_),
    .B(_11302_));
 sg13g2_nand2_1 _20399_ (.Y(_11304_),
    .A(_11300_),
    .B(_11298_));
 sg13g2_nand3b_1 _20400_ (.B(_11303_),
    .C(_11304_),
    .Y(_11305_),
    .A_N(_11115_));
 sg13g2_nand2_1 _20401_ (.Y(_11306_),
    .A(_11303_),
    .B(_11304_));
 sg13g2_nand2_1 _20402_ (.Y(_11307_),
    .A(_11306_),
    .B(_11274_));
 sg13g2_nand2_1 _20403_ (.Y(_11308_),
    .A(_11305_),
    .B(_11307_));
 sg13g2_nor2_1 _20404_ (.A(_09405_),
    .B(_10985_),
    .Y(_11309_));
 sg13g2_nor2b_1 _20405_ (.A(_11309_),
    .B_N(_09697_),
    .Y(_11310_));
 sg13g2_inv_1 _20406_ (.Y(_11311_),
    .A(_11050_));
 sg13g2_a22oi_1 _20407_ (.Y(_11312_),
    .B1(_11057_),
    .B2(_11311_),
    .A2(_06561_),
    .A1(_06810_));
 sg13g2_a22oi_1 _20408_ (.Y(_11313_),
    .B1(_10984_),
    .B2(_09405_),
    .A2(_06561_),
    .A1(_06809_));
 sg13g2_nand2_1 _20409_ (.Y(_11314_),
    .A(_11050_),
    .B(_11057_));
 sg13g2_nand4_1 _20410_ (.B(_11312_),
    .C(_11313_),
    .A(_11310_),
    .Y(_11315_),
    .D(_11314_));
 sg13g2_nand2_1 _20411_ (.Y(_11316_),
    .A(_11315_),
    .B(net126));
 sg13g2_inv_1 _20412_ (.Y(_11317_),
    .A(_09828_));
 sg13g2_a22oi_1 _20413_ (.Y(_11318_),
    .B1(_08063_),
    .B2(_11317_),
    .A2(_07584_),
    .A1(_07598_));
 sg13g2_nand4_1 _20414_ (.B(_09566_),
    .C(_05356_),
    .A(_09552_),
    .Y(_11319_),
    .D(_09553_));
 sg13g2_nand2_1 _20415_ (.Y(_11320_),
    .A(_08328_),
    .B(_08287_));
 sg13g2_nand3_1 _20416_ (.B(_11319_),
    .C(_11320_),
    .A(_11318_),
    .Y(_11321_));
 sg13g2_nor2_1 _20417_ (.A(_08288_),
    .B(_08328_),
    .Y(_11322_));
 sg13g2_a22oi_1 _20418_ (.Y(_11323_),
    .B1(_11317_),
    .B2(_08064_),
    .A2(_07584_),
    .A1(_07599_));
 sg13g2_nand2b_1 _20419_ (.Y(_11324_),
    .B(_07806_),
    .A_N(_09567_));
 sg13g2_nand3b_1 _20420_ (.B(_11323_),
    .C(_11324_),
    .Y(_11325_),
    .A_N(_11322_));
 sg13g2_o21ai_1 _20421_ (.B1(net126),
    .Y(_11326_),
    .A1(_11321_),
    .A2(_11325_));
 sg13g2_a21o_1 _20422_ (.A2(_11326_),
    .A1(_11316_),
    .B1(_06585_),
    .X(_11327_));
 sg13g2_nand2b_1 _20423_ (.Y(_11328_),
    .B(_07586_),
    .A_N(_11326_));
 sg13g2_nand3_1 _20424_ (.B(_06571_),
    .C(_11328_),
    .A(_11327_),
    .Y(_11329_));
 sg13g2_nand4_1 _20425_ (.B(_08463_),
    .C(_10232_),
    .A(_08459_),
    .Y(_11330_),
    .D(_10317_));
 sg13g2_o21ai_1 _20426_ (.B1(_08068_),
    .Y(_11331_),
    .A1(_09104_),
    .A2(_11311_));
 sg13g2_nor4_1 _20427_ (.A(_09407_),
    .B(_09608_),
    .C(_11330_),
    .D(_11331_),
    .Y(_11332_));
 sg13g2_a21oi_1 _20428_ (.A1(_09552_),
    .A2(_09553_),
    .Y(_11333_),
    .B1(_07708_));
 sg13g2_nor2_1 _20429_ (.A(_09104_),
    .B(_11050_),
    .Y(_11334_));
 sg13g2_nor4_1 _20430_ (.A(_09101_),
    .B(_11333_),
    .C(_11334_),
    .D(_07967_),
    .Y(_11335_));
 sg13g2_nor4_1 _20431_ (.A(_09719_),
    .B(_09859_),
    .C(_08096_),
    .D(_09544_),
    .Y(_11336_));
 sg13g2_nand4_1 _20432_ (.B(_09546_),
    .C(_11335_),
    .A(_11332_),
    .Y(_11337_),
    .D(_11336_));
 sg13g2_nor2_1 _20433_ (.A(_02056_),
    .B(_06574_),
    .Y(_11338_));
 sg13g2_nand3_1 _20434_ (.B(_11337_),
    .C(_11338_),
    .A(_11329_),
    .Y(_11339_));
 sg13g2_inv_1 _20435_ (.Y(_11340_),
    .A(_11313_));
 sg13g2_o21ai_1 _20436_ (.B1(_11314_),
    .Y(_11341_),
    .A1(_09697_),
    .A2(_09704_));
 sg13g2_nand2_1 _20437_ (.Y(_11342_),
    .A(_08971_),
    .B(_03870_));
 sg13g2_nand2b_1 _20438_ (.Y(_11343_),
    .B(_11342_),
    .A_N(_10633_));
 sg13g2_nand2b_1 _20439_ (.Y(_11344_),
    .B(_09281_),
    .A_N(_08423_));
 sg13g2_nor2_1 _20440_ (.A(_08422_),
    .B(_05205_),
    .Y(_11345_));
 sg13g2_nand2b_1 _20441_ (.Y(_11346_),
    .B(_11345_),
    .A_N(_11344_));
 sg13g2_nor4_1 _20442_ (.A(_06646_),
    .B(_10632_),
    .C(_11343_),
    .D(_11346_),
    .Y(_11347_));
 sg13g2_nand2_1 _20443_ (.Y(_11348_),
    .A(_11332_),
    .B(_11347_));
 sg13g2_nor4_1 _20444_ (.A(_11321_),
    .B(_11340_),
    .C(_11341_),
    .D(_11348_),
    .Y(_11349_));
 sg13g2_nor2_1 _20445_ (.A(_09697_),
    .B(_09703_),
    .Y(_11350_));
 sg13g2_inv_1 _20446_ (.Y(_11351_),
    .A(_11335_));
 sg13g2_inv_1 _20447_ (.Y(_11352_),
    .A(_11325_));
 sg13g2_inv_1 _20448_ (.Y(_11353_),
    .A(_09008_));
 sg13g2_nor2_1 _20449_ (.A(_09216_),
    .B(_11353_),
    .Y(_11354_));
 sg13g2_nand4_1 _20450_ (.B(_08419_),
    .C(_06642_),
    .A(_11354_),
    .Y(_11355_),
    .D(_10617_));
 sg13g2_nor2_1 _20451_ (.A(_11309_),
    .B(_11355_),
    .Y(_11356_));
 sg13g2_nand4_1 _20452_ (.B(_11312_),
    .C(_11336_),
    .A(_11352_),
    .Y(_11357_),
    .D(_11356_));
 sg13g2_nor3_1 _20453_ (.A(_11350_),
    .B(_11351_),
    .C(_11357_),
    .Y(_11358_));
 sg13g2_nand2_1 _20454_ (.Y(_11359_),
    .A(_11349_),
    .B(_11358_));
 sg13g2_o21ai_1 _20455_ (.B1(_06568_),
    .Y(_11360_),
    .A1(_06564_),
    .A2(net126));
 sg13g2_nand3_1 _20456_ (.B(_05084_),
    .C(_11360_),
    .A(_11359_),
    .Y(_11361_));
 sg13g2_nor3_1 _20457_ (.A(net126),
    .B(_11358_),
    .C(_11349_),
    .Y(_11362_));
 sg13g2_nand3_1 _20458_ (.B(_05073_),
    .C(_07914_),
    .A(_11362_),
    .Y(_11363_));
 sg13g2_nand3_1 _20459_ (.B(_11361_),
    .C(_11363_),
    .A(_11339_),
    .Y(_11364_));
 sg13g2_buf_1 _20460_ (.A(\b.gen_square[19].sq.mask ),
    .X(_11365_));
 sg13g2_nand2_1 _20461_ (.Y(_11366_),
    .A(_11364_),
    .B(_11365_));
 sg13g2_nor2_1 _20462_ (.A(_11366_),
    .B(_11308_),
    .Y(_11367_));
 sg13g2_nand2_1 _20463_ (.Y(_11368_),
    .A(_11306_),
    .B(_11289_));
 sg13g2_nand3_1 _20464_ (.B(_11304_),
    .C(_11286_),
    .A(_11303_),
    .Y(_11369_));
 sg13g2_nand2_1 _20465_ (.Y(_11370_),
    .A(_11362_),
    .B(_05073_));
 sg13g2_nand3_1 _20466_ (.B(net144),
    .C(_06581_),
    .A(_11359_),
    .Y(_11371_));
 sg13g2_nand2_1 _20467_ (.Y(_11372_),
    .A(_11370_),
    .B(_11371_));
 sg13g2_nand2_1 _20468_ (.Y(_11373_),
    .A(_11370_),
    .B(_06567_));
 sg13g2_nand2b_1 _20469_ (.Y(_11374_),
    .B(_06565_),
    .A_N(_06584_));
 sg13g2_nand3_1 _20470_ (.B(_11373_),
    .C(_11374_),
    .A(_11372_),
    .Y(_11375_));
 sg13g2_nand3_1 _20471_ (.B(net126),
    .C(_06583_),
    .A(_11315_),
    .Y(_11376_));
 sg13g2_nand2_1 _20472_ (.Y(_11377_),
    .A(_06571_),
    .B(_05108_));
 sg13g2_a21o_1 _20473_ (.A2(_11376_),
    .A1(_11327_),
    .B1(_11377_),
    .X(_11378_));
 sg13g2_nand2_1 _20474_ (.Y(_11379_),
    .A(_11375_),
    .B(_11378_));
 sg13g2_nand2_1 _20475_ (.Y(_11380_),
    .A(_11379_),
    .B(_11365_));
 sg13g2_nand3_1 _20476_ (.B(_11369_),
    .C(_11380_),
    .A(_11368_),
    .Y(_11381_));
 sg13g2_nand2_1 _20477_ (.Y(_11382_),
    .A(_11367_),
    .B(_11381_));
 sg13g2_nand2_1 _20478_ (.Y(_11383_),
    .A(_11368_),
    .B(_11369_));
 sg13g2_inv_1 _20479_ (.Y(_11384_),
    .A(_11380_));
 sg13g2_xnor2_1 _20480_ (.Y(_11385_),
    .A(_06566_),
    .B(_06584_));
 sg13g2_nand2b_1 _20481_ (.Y(_11386_),
    .B(_11347_),
    .A_N(_11355_));
 sg13g2_nand2b_1 _20482_ (.Y(_11387_),
    .B(_11386_),
    .A_N(_07916_));
 sg13g2_a21oi_1 _20483_ (.A1(_11328_),
    .A2(_11387_),
    .Y(_11388_),
    .B1(_11377_));
 sg13g2_a21oi_1 _20484_ (.A1(_11372_),
    .A2(_11385_),
    .Y(_11389_),
    .B1(_11388_));
 sg13g2_nand2_1 _20485_ (.Y(_11390_),
    .A(_11389_),
    .B(_11378_));
 sg13g2_nand2_1 _20486_ (.Y(_11391_),
    .A(_11390_),
    .B(_11365_));
 sg13g2_nand2_1 _20487_ (.Y(_11392_),
    .A(_11299_),
    .B(_11298_));
 sg13g2_nor2_1 _20488_ (.A(_11391_),
    .B(_11392_),
    .Y(_11393_));
 sg13g2_a21oi_1 _20489_ (.A1(_11383_),
    .A2(_11384_),
    .Y(_11394_),
    .B1(_11393_));
 sg13g2_nand2_1 _20490_ (.Y(_11395_),
    .A(_11382_),
    .B(_11394_));
 sg13g2_nand2_1 _20491_ (.Y(_11396_),
    .A(_11392_),
    .B(_11391_));
 sg13g2_nand2_1 _20492_ (.Y(_11397_),
    .A(_11395_),
    .B(_11396_));
 sg13g2_nand2b_1 _20493_ (.Y(_11398_),
    .B(_11397_),
    .A_N(_11308_));
 sg13g2_nand3_1 _20494_ (.B(_11396_),
    .C(_11366_),
    .A(_11395_),
    .Y(_11399_));
 sg13g2_buf_1 _20495_ (.A(_11399_),
    .X(_11400_));
 sg13g2_nor2_1 _20496_ (.A(_08958_),
    .B(_11048_),
    .Y(_11401_));
 sg13g2_nor4_1 _20497_ (.A(_09721_),
    .B(_09101_),
    .C(_11401_),
    .D(_07715_),
    .Y(_11402_));
 sg13g2_nor4_1 _20498_ (.A(_07704_),
    .B(_09003_),
    .C(_09859_),
    .D(_07967_),
    .Y(_11403_));
 sg13g2_nand2_1 _20499_ (.Y(_11404_),
    .A(_11402_),
    .B(_11403_));
 sg13g2_nor2_1 _20500_ (.A(_10975_),
    .B(_10987_),
    .Y(_11405_));
 sg13g2_nor2_1 _20501_ (.A(_06966_),
    .B(_07003_),
    .Y(_11406_));
 sg13g2_nor2_1 _20502_ (.A(_11048_),
    .B(_11056_),
    .Y(_11407_));
 sg13g2_nor2_1 _20503_ (.A(_09818_),
    .B(_09813_),
    .Y(_11408_));
 sg13g2_nor4_1 _20504_ (.A(_11405_),
    .B(_11406_),
    .C(_11407_),
    .D(_11408_),
    .Y(_11409_));
 sg13g2_a22oi_1 _20505_ (.Y(_11410_),
    .B1(_08656_),
    .B2(_08689_),
    .A2(_05900_),
    .A1(_05952_));
 sg13g2_o21ai_1 _20506_ (.B1(_11410_),
    .Y(_11411_),
    .A1(_09685_),
    .A2(_09679_));
 sg13g2_a21oi_1 _20507_ (.A1(_09143_),
    .A2(_09078_),
    .Y(_11412_),
    .B1(_11411_));
 sg13g2_nor2_1 _20508_ (.A(_10214_),
    .B(_04548_),
    .Y(_11413_));
 sg13g2_inv_1 _20509_ (.Y(_11414_),
    .A(_11413_));
 sg13g2_nor3_1 _20510_ (.A(_09129_),
    .B(_09737_),
    .C(_11143_),
    .Y(_11415_));
 sg13g2_inv_1 _20511_ (.Y(_11416_),
    .A(_11415_));
 sg13g2_nor4_1 _20512_ (.A(_07934_),
    .B(_06296_),
    .C(_11414_),
    .D(_11416_),
    .Y(_11417_));
 sg13g2_nand3_1 _20513_ (.B(_11412_),
    .C(_11417_),
    .A(_11409_),
    .Y(_11418_));
 sg13g2_nor2_1 _20514_ (.A(_11404_),
    .B(_11418_),
    .Y(_11419_));
 sg13g2_nor2_1 _20515_ (.A(_05854_),
    .B(_11419_),
    .Y(_11420_));
 sg13g2_nor2_1 _20516_ (.A(_10987_),
    .B(_10976_),
    .Y(_11421_));
 sg13g2_nor2_1 _20517_ (.A(_06966_),
    .B(_07004_),
    .Y(_11422_));
 sg13g2_nor2b_1 _20518_ (.A(_11056_),
    .B_N(_11048_),
    .Y(_11423_));
 sg13g2_nor2_1 _20519_ (.A(_09818_),
    .B(_09814_),
    .Y(_11424_));
 sg13g2_nor4_1 _20520_ (.A(_11421_),
    .B(_11422_),
    .C(_11423_),
    .D(_11424_),
    .Y(_11425_));
 sg13g2_nand2_1 _20521_ (.Y(_11426_),
    .A(_08688_),
    .B(_08656_));
 sg13g2_o21ai_1 _20522_ (.B1(_11426_),
    .Y(_11427_),
    .A1(_09079_),
    .A2(_09143_));
 sg13g2_a221oi_1 _20523_ (.B2(_09684_),
    .C1(_11427_),
    .B1(_09679_),
    .A1(_05951_),
    .Y(_11428_),
    .A2(_05900_));
 sg13g2_nor2_1 _20524_ (.A(_10241_),
    .B(_06461_),
    .Y(_11429_));
 sg13g2_nor2_1 _20525_ (.A(_07896_),
    .B(_05019_),
    .Y(_11430_));
 sg13g2_nand2_1 _20526_ (.Y(_11431_),
    .A(_11429_),
    .B(_11430_));
 sg13g2_nor4_1 _20527_ (.A(_09149_),
    .B(_09745_),
    .C(_11129_),
    .D(_11431_),
    .Y(_11432_));
 sg13g2_nor2_1 _20528_ (.A(_08934_),
    .B(_09113_),
    .Y(_11433_));
 sg13g2_nand2_1 _20529_ (.Y(_11434_),
    .A(_11048_),
    .B(_09041_));
 sg13g2_nand4_1 _20530_ (.B(_08463_),
    .C(_11433_),
    .A(_09612_),
    .Y(_11435_),
    .D(_11434_));
 sg13g2_nor4_1 _20531_ (.A(_07815_),
    .B(_07990_),
    .C(_09608_),
    .D(_11435_),
    .Y(_11436_));
 sg13g2_nand4_1 _20532_ (.B(_11428_),
    .C(_11432_),
    .A(_11425_),
    .Y(_11437_),
    .D(_11436_));
 sg13g2_nand3_1 _20533_ (.B(_05074_),
    .C(_11437_),
    .A(_11420_),
    .Y(_11438_));
 sg13g2_buf_1 _20534_ (.A(_11438_),
    .X(_11439_));
 sg13g2_nand2b_1 _20535_ (.Y(_11440_),
    .B(_11419_),
    .A_N(_11437_));
 sg13g2_o21ai_1 _20536_ (.B1(_05852_),
    .Y(_11441_),
    .A1(_05849_),
    .A2(_05854_));
 sg13g2_nand3_1 _20537_ (.B(_05085_),
    .C(_11441_),
    .A(_11440_),
    .Y(_11442_));
 sg13g2_o21ai_1 _20538_ (.B1(_11442_),
    .Y(_11443_),
    .A1(_05849_),
    .A2(_11439_));
 sg13g2_a21o_1 _20539_ (.A2(_11412_),
    .A1(_11428_),
    .B1(_05905_),
    .X(_11444_));
 sg13g2_nor2_1 _20540_ (.A(_05904_),
    .B(_11444_),
    .Y(_11445_));
 sg13g2_a21o_1 _20541_ (.A2(_11409_),
    .A1(_11425_),
    .B1(_05905_),
    .X(_11446_));
 sg13g2_a21o_1 _20542_ (.A2(_11444_),
    .A1(_11446_),
    .B1(_05902_),
    .X(_11447_));
 sg13g2_nand3b_1 _20543_ (.B(_11447_),
    .C(_05857_),
    .Y(_11448_),
    .A_N(_11445_));
 sg13g2_nor2b_1 _20544_ (.A(_11404_),
    .B_N(_11436_),
    .Y(_11449_));
 sg13g2_o21ai_1 _20545_ (.B1(_05856_),
    .Y(_11450_),
    .A1(_05905_),
    .A2(_11449_));
 sg13g2_and3_1 _20546_ (.X(_11451_),
    .A(_11448_),
    .B(_05110_),
    .C(_11450_));
 sg13g2_buf_1 _20547_ (.A(\b.gen_square[20].sq.mask ),
    .X(_11452_));
 sg13g2_o21ai_1 _20548_ (.B1(_11452_),
    .Y(_11453_),
    .A1(_11443_),
    .A2(_11451_));
 sg13g2_nand3_1 _20549_ (.B(_11400_),
    .C(_11453_),
    .A(_11398_),
    .Y(_11454_));
 sg13g2_o21ai_1 _20550_ (.B1(_11447_),
    .Y(_11455_),
    .A1(_06968_),
    .A2(_11446_));
 sg13g2_nand2_1 _20551_ (.Y(_11456_),
    .A(_11455_),
    .B(_05110_));
 sg13g2_a21oi_1 _20552_ (.A1(_11417_),
    .A2(_11432_),
    .Y(_11457_),
    .B1(_07749_));
 sg13g2_nor2_1 _20553_ (.A(_02056_),
    .B(_05856_),
    .Y(_11458_));
 sg13g2_o21ai_1 _20554_ (.B1(_11458_),
    .Y(_11459_),
    .A1(_11457_),
    .A2(_11445_));
 sg13g2_nand3_1 _20555_ (.B(_05085_),
    .C(_05905_),
    .A(_11440_),
    .Y(_11460_));
 sg13g2_nand2_1 _20556_ (.Y(_11461_),
    .A(_11460_),
    .B(_11439_));
 sg13g2_xnor2_1 _20557_ (.Y(_11462_),
    .A(_05846_),
    .B(_05901_));
 sg13g2_nand2_1 _20558_ (.Y(_11463_),
    .A(_11461_),
    .B(_11462_));
 sg13g2_nand3_1 _20559_ (.B(_11459_),
    .C(_11463_),
    .A(_11456_),
    .Y(_11464_));
 sg13g2_nand2_1 _20560_ (.Y(_11465_),
    .A(_11464_),
    .B(_11452_));
 sg13g2_nor2b_1 _20561_ (.A(_11392_),
    .B_N(_11391_),
    .Y(_11466_));
 sg13g2_xnor2_1 _20562_ (.Y(_11467_),
    .A(_11465_),
    .B(_11466_));
 sg13g2_nand2_1 _20563_ (.Y(_11468_),
    .A(_11454_),
    .B(_11467_));
 sg13g2_nand2b_1 _20564_ (.Y(_11469_),
    .B(_05850_),
    .A_N(_05901_));
 sg13g2_nand2_1 _20565_ (.Y(_11470_),
    .A(_11439_),
    .B(_05851_));
 sg13g2_nand3_1 _20566_ (.B(_11469_),
    .C(_11470_),
    .A(_11461_),
    .Y(_11471_));
 sg13g2_nand2_1 _20567_ (.Y(_11472_),
    .A(_11471_),
    .B(_11456_));
 sg13g2_nand2_1 _20568_ (.Y(_11473_),
    .A(_11472_),
    .B(_11452_));
 sg13g2_nand2b_1 _20569_ (.Y(_11474_),
    .B(_11397_),
    .A_N(_11383_));
 sg13g2_nand3_1 _20570_ (.B(_11384_),
    .C(_11396_),
    .A(_11395_),
    .Y(_11475_));
 sg13g2_nand3b_1 _20571_ (.B(_11474_),
    .C(_11475_),
    .Y(_11476_),
    .A_N(_11473_));
 sg13g2_nand2_1 _20572_ (.Y(_11477_),
    .A(_11474_),
    .B(_11475_));
 sg13g2_nand2_1 _20573_ (.Y(_11478_),
    .A(_11477_),
    .B(_11473_));
 sg13g2_nand2_1 _20574_ (.Y(_11479_),
    .A(_11476_),
    .B(_11478_));
 sg13g2_nor2_1 _20575_ (.A(_11468_),
    .B(_11479_),
    .Y(_11480_));
 sg13g2_a21oi_1 _20576_ (.A1(_11398_),
    .A2(_11400_),
    .Y(_11481_),
    .B1(_11453_));
 sg13g2_nand2_1 _20577_ (.Y(_11482_),
    .A(_11480_),
    .B(_11481_));
 sg13g2_nor2b_1 _20578_ (.A(_11465_),
    .B_N(_11466_),
    .Y(_11483_));
 sg13g2_nor2b_1 _20579_ (.A(_11476_),
    .B_N(_11467_),
    .Y(_11484_));
 sg13g2_nor2_1 _20580_ (.A(_11483_),
    .B(_11484_),
    .Y(_11485_));
 sg13g2_nand2_1 _20581_ (.Y(_11486_),
    .A(_11398_),
    .B(_11400_));
 sg13g2_nand3_1 _20582_ (.B(_11485_),
    .C(_11486_),
    .A(_11482_),
    .Y(_11487_));
 sg13g2_o21ai_1 _20583_ (.B1(_11453_),
    .Y(_11488_),
    .A1(_11483_),
    .A2(_11484_));
 sg13g2_nand2_1 _20584_ (.Y(_11489_),
    .A(_11487_),
    .B(_11488_));
 sg13g2_nand2_1 _20585_ (.Y(_11490_),
    .A(_11482_),
    .B(_11485_));
 sg13g2_nand2_1 _20586_ (.Y(_11491_),
    .A(_11490_),
    .B(_11473_));
 sg13g2_inv_1 _20587_ (.Y(_11492_),
    .A(_11477_));
 sg13g2_nand3_1 _20588_ (.B(_11485_),
    .C(_11492_),
    .A(_11482_),
    .Y(_11493_));
 sg13g2_nand2_1 _20589_ (.Y(_11494_),
    .A(_11491_),
    .B(_11493_));
 sg13g2_nor2_1 _20590_ (.A(_07099_),
    .B(_07138_),
    .Y(_11495_));
 sg13g2_inv_1 _20591_ (.Y(_11496_),
    .A(_11046_));
 sg13g2_inv_1 _20592_ (.Y(_11497_),
    .A(_11054_));
 sg13g2_nor2_1 _20593_ (.A(_11496_),
    .B(_11497_),
    .Y(_11498_));
 sg13g2_nor2_1 _20594_ (.A(_10977_),
    .B(_10989_),
    .Y(_11499_));
 sg13g2_nor2_1 _20595_ (.A(_09056_),
    .B(_09050_),
    .Y(_11500_));
 sg13g2_nor4_1 _20596_ (.A(_11495_),
    .B(_11498_),
    .C(_11499_),
    .D(_11500_),
    .Y(_11501_));
 sg13g2_o21ai_1 _20597_ (.B1(_08732_),
    .Y(_11502_),
    .A1(_08938_),
    .A2(_11496_));
 sg13g2_or4_1 _20598_ (.A(_07724_),
    .B(_10036_),
    .C(_09101_),
    .D(_07715_),
    .X(_11503_));
 sg13g2_nor4_1 _20599_ (.A(_09106_),
    .B(_09003_),
    .C(_11502_),
    .D(_11503_),
    .Y(_11504_));
 sg13g2_nand2_1 _20600_ (.Y(_11505_),
    .A(_08805_),
    .B(_08797_));
 sg13g2_o21ai_1 _20601_ (.B1(_11505_),
    .Y(_11506_),
    .A1(_08961_),
    .A2(_08955_));
 sg13g2_a22oi_1 _20602_ (.Y(_11507_),
    .B1(_09835_),
    .B2(_09837_),
    .A2(_05318_),
    .A1(_05524_));
 sg13g2_nor2b_1 _20603_ (.A(_11506_),
    .B_N(_11507_),
    .Y(_11508_));
 sg13g2_nor4_1 _20604_ (.A(_09865_),
    .B(_07246_),
    .C(_10122_),
    .D(_07758_),
    .Y(_11509_));
 sg13g2_nor2_1 _20605_ (.A(_10120_),
    .B(_06641_),
    .Y(_11510_));
 sg13g2_nor2_1 _20606_ (.A(_07743_),
    .B(_11353_),
    .Y(_11511_));
 sg13g2_and3_1 _20607_ (.X(_11512_),
    .A(_11509_),
    .B(_11510_),
    .C(_11511_));
 sg13g2_nand4_1 _20608_ (.B(_11504_),
    .C(_11508_),
    .A(_11501_),
    .Y(_11513_),
    .D(_11512_));
 sg13g2_nor2_1 _20609_ (.A(_07099_),
    .B(_07139_),
    .Y(_11514_));
 sg13g2_nor2_1 _20610_ (.A(_11046_),
    .B(_11497_),
    .Y(_11515_));
 sg13g2_nor2_1 _20611_ (.A(_10989_),
    .B(_10978_),
    .Y(_11516_));
 sg13g2_nor2_1 _20612_ (.A(_09056_),
    .B(_09051_),
    .Y(_11517_));
 sg13g2_nor4_1 _20613_ (.A(_11514_),
    .B(_11515_),
    .C(_11516_),
    .D(_11517_),
    .Y(_11518_));
 sg13g2_nor2_1 _20614_ (.A(_08798_),
    .B(_08805_),
    .Y(_11519_));
 sg13g2_nand2_1 _20615_ (.Y(_11520_),
    .A(_05523_),
    .B(_05318_));
 sg13g2_o21ai_1 _20616_ (.B1(_11520_),
    .Y(_11521_),
    .A1(_09835_),
    .A2(_09838_));
 sg13g2_nor2_1 _20617_ (.A(_08955_),
    .B(_08962_),
    .Y(_11522_));
 sg13g2_nor3_1 _20618_ (.A(_11519_),
    .B(_11521_),
    .C(_11522_),
    .Y(_11523_));
 sg13g2_nand2b_1 _20619_ (.Y(_11524_),
    .B(_11342_),
    .A_N(_09846_));
 sg13g2_nand2_1 _20620_ (.Y(_11525_),
    .A(_07836_),
    .B(_07161_));
 sg13g2_nor4_1 _20621_ (.A(_10170_),
    .B(_10171_),
    .C(_11524_),
    .D(_11525_),
    .Y(_11526_));
 sg13g2_nand2b_1 _20622_ (.Y(_11527_),
    .B(_11496_),
    .A_N(_08938_));
 sg13g2_nand4_1 _20623_ (.B(_08813_),
    .C(_10892_),
    .A(_11433_),
    .Y(_11528_),
    .D(_11527_));
 sg13g2_nor4_1 _20624_ (.A(_07815_),
    .B(_07807_),
    .C(_09118_),
    .D(_11528_),
    .Y(_11529_));
 sg13g2_nand4_1 _20625_ (.B(_11523_),
    .C(_11526_),
    .A(_11518_),
    .Y(_11530_),
    .D(_11529_));
 sg13g2_nor2_1 _20626_ (.A(_11513_),
    .B(_11530_),
    .Y(_11531_));
 sg13g2_inv_1 _20627_ (.Y(_11532_),
    .A(_11531_));
 sg13g2_nand3_1 _20628_ (.B(net113),
    .C(_05319_),
    .A(_11532_),
    .Y(_11533_));
 sg13g2_nand4_1 _20629_ (.B(_11513_),
    .C(net162),
    .A(_11530_),
    .Y(_11534_),
    .D(_05319_));
 sg13g2_buf_1 _20630_ (.A(_11534_),
    .X(_11535_));
 sg13g2_nand2_1 _20631_ (.Y(_11536_),
    .A(_11533_),
    .B(_11535_));
 sg13g2_nand2_1 _20632_ (.Y(_11537_),
    .A(_11535_),
    .B(_05277_));
 sg13g2_nand2b_1 _20633_ (.Y(_11538_),
    .B(_05276_),
    .A_N(_05323_));
 sg13g2_nand3_1 _20634_ (.B(_11537_),
    .C(_11538_),
    .A(_11536_),
    .Y(_11539_));
 sg13g2_a21oi_1 _20635_ (.A1(_11518_),
    .A2(_11501_),
    .Y(_11540_),
    .B1(_05319_));
 sg13g2_inv_1 _20636_ (.Y(_11541_),
    .A(_11540_));
 sg13g2_a21o_1 _20637_ (.A2(_11523_),
    .A1(_11508_),
    .B1(_05319_),
    .X(_11542_));
 sg13g2_a21o_1 _20638_ (.A2(_11542_),
    .A1(_11541_),
    .B1(_05324_),
    .X(_11543_));
 sg13g2_o21ai_1 _20639_ (.B1(_11543_),
    .Y(_11544_),
    .A1(_07102_),
    .A2(_11541_));
 sg13g2_nand2_1 _20640_ (.Y(_11545_),
    .A(_11544_),
    .B(net112));
 sg13g2_nand2_1 _20641_ (.Y(_11546_),
    .A(_11539_),
    .B(_11545_));
 sg13g2_buf_1 _20642_ (.A(\b.gen_square[21].sq.mask ),
    .X(_11547_));
 sg13g2_nand2_1 _20643_ (.Y(_11548_),
    .A(_11546_),
    .B(_11547_));
 sg13g2_inv_1 _20644_ (.Y(_11549_),
    .A(_11548_));
 sg13g2_xnor2_1 _20645_ (.Y(_11550_),
    .A(_05272_),
    .B(_05323_));
 sg13g2_nand2_1 _20646_ (.Y(_11551_),
    .A(_11536_),
    .B(_11550_));
 sg13g2_a21oi_1 _20647_ (.A1(_11512_),
    .A2(_11526_),
    .Y(_11552_),
    .B1(_07898_));
 sg13g2_nor2_1 _20648_ (.A(_05322_),
    .B(_11542_),
    .Y(_11553_));
 sg13g2_nor2_1 _20649_ (.A(_02067_),
    .B(_05282_),
    .Y(_11554_));
 sg13g2_o21ai_1 _20650_ (.B1(_11554_),
    .Y(_11555_),
    .A1(_11552_),
    .A2(_11553_));
 sg13g2_nand3_1 _20651_ (.B(_11551_),
    .C(_11555_),
    .A(_11545_),
    .Y(_11556_));
 sg13g2_nand2_1 _20652_ (.Y(_11557_),
    .A(_11556_),
    .B(_11547_));
 sg13g2_nand2_1 _20653_ (.Y(_11558_),
    .A(_11466_),
    .B(_11465_));
 sg13g2_nor2_1 _20654_ (.A(_11557_),
    .B(_11558_),
    .Y(_11559_));
 sg13g2_a21oi_1 _20655_ (.A1(_11494_),
    .A2(_11549_),
    .Y(_11560_),
    .B1(_11559_));
 sg13g2_o21ai_1 _20656_ (.B1(_05278_),
    .Y(_11561_),
    .A1(_05275_),
    .A2(_05280_));
 sg13g2_nand3_1 _20657_ (.B(net96),
    .C(_11561_),
    .A(_11532_),
    .Y(_11562_));
 sg13g2_o21ai_1 _20658_ (.B1(_11562_),
    .Y(_11563_),
    .A1(_05275_),
    .A2(_11535_));
 sg13g2_nand3b_1 _20659_ (.B(_11543_),
    .C(_05283_),
    .Y(_11564_),
    .A_N(_11553_));
 sg13g2_inv_1 _20660_ (.Y(_11565_),
    .A(_05284_));
 sg13g2_nand3_1 _20661_ (.B(_05282_),
    .C(_11529_),
    .A(_11504_),
    .Y(_11566_));
 sg13g2_and4_1 _20662_ (.A(_05112_),
    .B(_11564_),
    .C(_11565_),
    .D(_11566_),
    .X(_11567_));
 sg13g2_o21ai_1 _20663_ (.B1(_11547_),
    .Y(_11568_),
    .A1(_11563_),
    .A2(_11567_));
 sg13g2_a21oi_1 _20664_ (.A1(_11487_),
    .A2(_11488_),
    .Y(_11569_),
    .B1(_11568_));
 sg13g2_nand3_1 _20665_ (.B(_11493_),
    .C(_11548_),
    .A(_11491_),
    .Y(_11570_));
 sg13g2_nand2_1 _20666_ (.Y(_11571_),
    .A(_11569_),
    .B(_11570_));
 sg13g2_nand2_1 _20667_ (.Y(_11572_),
    .A(_11560_),
    .B(_11571_));
 sg13g2_nand2_1 _20668_ (.Y(_11573_),
    .A(_11558_),
    .B(_11557_));
 sg13g2_nand2_1 _20669_ (.Y(_11574_),
    .A(_11572_),
    .B(_11573_));
 sg13g2_nand2b_1 _20670_ (.Y(_11575_),
    .B(_11574_),
    .A_N(_11489_));
 sg13g2_nand3b_1 _20671_ (.B(_11572_),
    .C(_11573_),
    .Y(_11576_),
    .A_N(_11568_));
 sg13g2_nand2_1 _20672_ (.Y(_11577_),
    .A(_11575_),
    .B(_11576_));
 sg13g2_nor2_1 _20673_ (.A(_11043_),
    .B(_11577_),
    .Y(_11578_));
 sg13g2_nand2_1 _20674_ (.Y(_11579_),
    .A(_11574_),
    .B(_11494_));
 sg13g2_nand3_1 _20675_ (.B(_11573_),
    .C(_11548_),
    .A(_11572_),
    .Y(_11580_));
 sg13g2_nand3_1 _20676_ (.B(net96),
    .C(_04284_),
    .A(_11035_),
    .Y(_11581_));
 sg13g2_nand2_1 _20677_ (.Y(_11582_),
    .A(_11039_),
    .B(_11581_));
 sg13g2_nand2_1 _20678_ (.Y(_11583_),
    .A(_11039_),
    .B(_04205_));
 sg13g2_nand2b_1 _20679_ (.Y(_11584_),
    .B(_04204_),
    .A_N(_04290_));
 sg13g2_nand3_1 _20680_ (.B(_11583_),
    .C(_11584_),
    .A(_11582_),
    .Y(_11585_));
 sg13g2_nand2b_1 _20681_ (.Y(_11586_),
    .B(_04289_),
    .A_N(_10998_));
 sg13g2_nand2_1 _20682_ (.Y(_11587_),
    .A(_11008_),
    .B(_11586_));
 sg13g2_nand2_1 _20683_ (.Y(_11588_),
    .A(_11587_),
    .B(net95));
 sg13g2_nand2_1 _20684_ (.Y(_11589_),
    .A(_11585_),
    .B(_11588_));
 sg13g2_nand2_1 _20685_ (.Y(_11590_),
    .A(_11589_),
    .B(_11042_));
 sg13g2_nand3_1 _20686_ (.B(_11580_),
    .C(_11590_),
    .A(_11579_),
    .Y(_11591_));
 sg13g2_nand2_1 _20687_ (.Y(_11592_),
    .A(_11578_),
    .B(_11591_));
 sg13g2_nand2_1 _20688_ (.Y(_11593_),
    .A(_11579_),
    .B(_11580_));
 sg13g2_inv_1 _20689_ (.Y(_11594_),
    .A(_11590_));
 sg13g2_nor2_1 _20690_ (.A(_02078_),
    .B(_08936_),
    .Y(_11595_));
 sg13g2_nand2_1 _20691_ (.Y(_11596_),
    .A(_11024_),
    .B(_11030_));
 sg13g2_nand2_1 _20692_ (.Y(_11597_),
    .A(_11596_),
    .B(_07745_));
 sg13g2_nand2_1 _20693_ (.Y(_11598_),
    .A(_11009_),
    .B(_11597_));
 sg13g2_xnor2_1 _20694_ (.Y(_11599_),
    .A(_04200_),
    .B(_04290_));
 sg13g2_a22oi_1 _20695_ (.Y(_11600_),
    .B1(_11599_),
    .B2(_11582_),
    .A2(_11598_),
    .A1(_11595_));
 sg13g2_nand2_1 _20696_ (.Y(_11601_),
    .A(_11600_),
    .B(_11588_));
 sg13g2_nand2_1 _20697_ (.Y(_11602_),
    .A(_11601_),
    .B(_11042_));
 sg13g2_inv_1 _20698_ (.Y(_11603_),
    .A(_11602_));
 sg13g2_nor2b_1 _20699_ (.A(_11558_),
    .B_N(_11557_),
    .Y(_11604_));
 sg13g2_xnor2_1 _20700_ (.Y(_11605_),
    .A(_11603_),
    .B(_11604_));
 sg13g2_a21oi_1 _20701_ (.A1(_11593_),
    .A2(_11594_),
    .Y(_11606_),
    .B1(_11605_));
 sg13g2_nand2_1 _20702_ (.Y(_11607_),
    .A(_11592_),
    .B(_11606_));
 sg13g2_inv_1 _20703_ (.Y(_11608_),
    .A(_11604_));
 sg13g2_nand2_1 _20704_ (.Y(_11609_),
    .A(_11608_),
    .B(_11602_));
 sg13g2_nand3b_1 _20705_ (.B(_11607_),
    .C(_11609_),
    .Y(_11610_),
    .A_N(_11043_));
 sg13g2_nand2_1 _20706_ (.Y(_11611_),
    .A(_11607_),
    .B(_11609_));
 sg13g2_nand2_1 _20707_ (.Y(_11612_),
    .A(_11611_),
    .B(_11577_));
 sg13g2_nand2_1 _20708_ (.Y(_11613_),
    .A(_11610_),
    .B(_11612_));
 sg13g2_nor2_1 _20709_ (.A(_06722_),
    .B(_07519_),
    .Y(_11614_));
 sg13g2_nor2_1 _20710_ (.A(_06670_),
    .B(_06722_),
    .Y(_11615_));
 sg13g2_a21oi_1 _20711_ (.A1(_08281_),
    .A2(net81),
    .Y(_11616_),
    .B1(_05317_));
 sg13g2_inv_1 _20712_ (.Y(_11617_),
    .A(_11616_));
 sg13g2_a21oi_1 _20713_ (.A1(_07137_),
    .A2(net81),
    .Y(_11618_),
    .B1(_04197_));
 sg13g2_nor2_1 _20714_ (.A(_11617_),
    .B(_11618_),
    .Y(_11619_));
 sg13g2_o21ai_1 _20715_ (.B1(_06706_),
    .Y(_11620_),
    .A1(_07952_),
    .A2(_07697_));
 sg13g2_a21oi_1 _20716_ (.A1(_11620_),
    .A2(net33),
    .Y(_11621_),
    .B1(_06688_));
 sg13g2_inv_1 _20717_ (.Y(_11622_),
    .A(_11621_));
 sg13g2_a21oi_1 _20718_ (.A1(_07690_),
    .A2(_06697_),
    .Y(_11623_),
    .B1(_06731_));
 sg13g2_inv_1 _20719_ (.Y(_11624_),
    .A(_11623_));
 sg13g2_a21oi_1 _20720_ (.A1(_11624_),
    .A2(_04154_),
    .Y(_11625_),
    .B1(_04224_));
 sg13g2_nor2_1 _20721_ (.A(_11622_),
    .B(_11625_),
    .Y(_11626_));
 sg13g2_nor2_1 _20722_ (.A(_10013_),
    .B(_10008_),
    .Y(_11627_));
 sg13g2_inv_1 _20723_ (.Y(_11628_),
    .A(_11627_));
 sg13g2_nor2_1 _20724_ (.A(_10614_),
    .B(_07246_),
    .Y(_11629_));
 sg13g2_nand2_1 _20725_ (.Y(_11630_),
    .A(_11629_),
    .B(_09866_));
 sg13g2_inv_1 _20726_ (.Y(_11631_),
    .A(_11630_));
 sg13g2_nand3_1 _20727_ (.B(_08842_),
    .C(_11631_),
    .A(_11628_),
    .Y(_11632_));
 sg13g2_a21oi_1 _20728_ (.A1(_10980_),
    .A2(_04217_),
    .Y(_11633_),
    .B1(_04220_));
 sg13g2_inv_1 _20729_ (.Y(_11634_),
    .A(_10990_));
 sg13g2_a21oi_1 _20730_ (.A1(_11634_),
    .A2(net47),
    .Y(_11635_),
    .B1(_04295_));
 sg13g2_nand2b_1 _20731_ (.Y(_11636_),
    .B(_11635_),
    .A_N(_11633_));
 sg13g2_nand2b_1 _20732_ (.Y(_11637_),
    .B(_07516_),
    .A_N(_07490_));
 sg13g2_nor4_1 _20733_ (.A(_09001_),
    .B(_10036_),
    .C(_10897_),
    .D(_08840_),
    .Y(_11638_));
 sg13g2_nand3_1 _20734_ (.B(_11637_),
    .C(_11638_),
    .A(_11636_),
    .Y(_11639_));
 sg13g2_nor4_1 _20735_ (.A(_11619_),
    .B(_11626_),
    .C(_11632_),
    .D(_11639_),
    .Y(_11640_));
 sg13g2_inv_1 _20736_ (.Y(_11641_),
    .A(_11640_));
 sg13g2_nor2b_1 _20737_ (.A(_10008_),
    .B_N(_10013_),
    .Y(_11642_));
 sg13g2_a221oi_1 _20738_ (.B2(_11635_),
    .C1(_11642_),
    .B1(_11633_),
    .A1(_07490_),
    .Y(_11643_),
    .A2(_07516_));
 sg13g2_a22oi_1 _20739_ (.Y(_11644_),
    .B1(_11621_),
    .B2(_11625_),
    .A2(_11616_),
    .A1(_11618_));
 sg13g2_nor2_1 _20740_ (.A(_10633_),
    .B(_07160_),
    .Y(_11645_));
 sg13g2_inv_1 _20741_ (.Y(_11646_),
    .A(_11645_));
 sg13g2_nor2_1 _20742_ (.A(_09848_),
    .B(_11646_),
    .Y(_11647_));
 sg13g2_nand3_1 _20743_ (.B(_10892_),
    .C(_10893_),
    .A(_08810_),
    .Y(_11648_));
 sg13g2_nor3_1 _20744_ (.A(_07801_),
    .B(_08940_),
    .C(_11648_),
    .Y(_11649_));
 sg13g2_nand4_1 _20745_ (.B(_11644_),
    .C(_11647_),
    .A(_11643_),
    .Y(_11650_),
    .D(_11649_));
 sg13g2_nor2_1 _20746_ (.A(_11641_),
    .B(_11650_),
    .Y(_11651_));
 sg13g2_nor4_1 _20747_ (.A(_07412_),
    .B(_11614_),
    .C(_11615_),
    .D(_11651_),
    .Y(_11652_));
 sg13g2_nand4_1 _20748_ (.B(_11641_),
    .C(_05077_),
    .A(_11650_),
    .Y(_11653_),
    .D(_07519_));
 sg13g2_buf_1 _20749_ (.A(_11653_),
    .X(_11654_));
 sg13g2_a21oi_1 _20750_ (.A1(_11622_),
    .A2(_11617_),
    .Y(_11655_),
    .B1(_07519_));
 sg13g2_inv_1 _20751_ (.Y(_11656_),
    .A(_11655_));
 sg13g2_nor2_1 _20752_ (.A(_06672_),
    .B(_11656_),
    .Y(_11657_));
 sg13g2_nand4_1 _20753_ (.B(_11636_),
    .C(_11628_),
    .A(_11643_),
    .Y(_11658_),
    .D(_11637_));
 sg13g2_nand2_1 _20754_ (.Y(_11659_),
    .A(_11658_),
    .B(_06664_));
 sg13g2_a21o_1 _20755_ (.A2(_11656_),
    .A1(_11659_),
    .B1(_06669_),
    .X(_11660_));
 sg13g2_nand3b_1 _20756_ (.B(_11660_),
    .C(_06677_),
    .Y(_11661_),
    .A_N(_11657_));
 sg13g2_nand4_1 _20757_ (.B(_08942_),
    .C(_08842_),
    .A(_11649_),
    .Y(_11662_),
    .D(_11638_));
 sg13g2_nor2_1 _20758_ (.A(net72),
    .B(_06678_),
    .Y(_11663_));
 sg13g2_nand3_1 _20759_ (.B(_11662_),
    .C(_11663_),
    .A(_11661_),
    .Y(_11664_));
 sg13g2_o21ai_1 _20760_ (.B1(_11664_),
    .Y(_11665_),
    .A1(_06666_),
    .A2(_11654_));
 sg13g2_buf_1 _20761_ (.A(\b.gen_square[23].sq.mask ),
    .X(_11666_));
 sg13g2_o21ai_1 _20762_ (.B1(_11666_),
    .Y(_11667_),
    .A1(_11652_),
    .A2(_11665_));
 sg13g2_nor2_1 _20763_ (.A(_11667_),
    .B(_11613_),
    .Y(_11668_));
 sg13g2_nand2_1 _20764_ (.Y(_11669_),
    .A(_11611_),
    .B(_11593_));
 sg13g2_nand3_1 _20765_ (.B(_11609_),
    .C(_11590_),
    .A(_11607_),
    .Y(_11670_));
 sg13g2_inv_1 _20766_ (.Y(_11671_),
    .A(_11651_));
 sg13g2_nand3_1 _20767_ (.B(net76),
    .C(_07519_),
    .A(_11671_),
    .Y(_11672_));
 sg13g2_nand2_1 _20768_ (.Y(_11673_),
    .A(_11672_),
    .B(_11654_));
 sg13g2_nand2_1 _20769_ (.Y(_11674_),
    .A(_11654_),
    .B(_06722_));
 sg13g2_nand2b_1 _20770_ (.Y(_11675_),
    .B(_06721_),
    .A_N(_06667_));
 sg13g2_nand3_1 _20771_ (.B(_11674_),
    .C(_11675_),
    .A(_11673_),
    .Y(_11676_));
 sg13g2_nand3_1 _20772_ (.B(_06664_),
    .C(_07517_),
    .A(_11658_),
    .Y(_11677_));
 sg13g2_nand2_1 _20773_ (.Y(_11678_),
    .A(_11660_),
    .B(_11677_));
 sg13g2_nor2_1 _20774_ (.A(net83),
    .B(_08942_),
    .Y(_11679_));
 sg13g2_nand2_1 _20775_ (.Y(_11680_),
    .A(_11678_),
    .B(_11679_));
 sg13g2_nand2_1 _20776_ (.Y(_11681_),
    .A(_11676_),
    .B(_11680_));
 sg13g2_nand2_1 _20777_ (.Y(_11682_),
    .A(_11681_),
    .B(_11666_));
 sg13g2_nand3_1 _20778_ (.B(_11670_),
    .C(_11682_),
    .A(_11669_),
    .Y(_11683_));
 sg13g2_nand2_1 _20779_ (.Y(_11684_),
    .A(_11668_),
    .B(_11683_));
 sg13g2_nand2_1 _20780_ (.Y(_11685_),
    .A(_11669_),
    .B(_11670_));
 sg13g2_inv_1 _20781_ (.Y(_11686_),
    .A(_11682_));
 sg13g2_xnor2_1 _20782_ (.Y(_11687_),
    .A(_06668_),
    .B(_06667_));
 sg13g2_nand2_1 _20783_ (.Y(_11688_),
    .A(_11673_),
    .B(_11687_));
 sg13g2_a21oi_1 _20784_ (.A1(_11647_),
    .A2(_11631_),
    .Y(_11689_),
    .B1(_08666_));
 sg13g2_o21ai_1 _20785_ (.B1(_11679_),
    .Y(_11690_),
    .A1(_11689_),
    .A2(_11657_));
 sg13g2_nand3_1 _20786_ (.B(_11688_),
    .C(_11690_),
    .A(_11680_),
    .Y(_11691_));
 sg13g2_nand2_2 _20787_ (.Y(_11692_),
    .A(_11691_),
    .B(_11666_));
 sg13g2_nor2_1 _20788_ (.A(_11603_),
    .B(_11608_),
    .Y(_11693_));
 sg13g2_inv_1 _20789_ (.Y(_11694_),
    .A(_11693_));
 sg13g2_nor2_1 _20790_ (.A(_11692_),
    .B(_11694_),
    .Y(_11695_));
 sg13g2_a21oi_1 _20791_ (.A1(_11685_),
    .A2(_11686_),
    .Y(_11696_),
    .B1(_11695_));
 sg13g2_nand2_1 _20792_ (.Y(_11697_),
    .A(_11684_),
    .B(_11696_));
 sg13g2_nand2_2 _20793_ (.Y(_11698_),
    .A(_11694_),
    .B(_11692_));
 sg13g2_nand2_2 _20794_ (.Y(_11699_),
    .A(_11697_),
    .B(_11698_));
 sg13g2_nand2b_1 _20795_ (.Y(_11700_),
    .B(_11699_),
    .A_N(_11613_));
 sg13g2_nand3_1 _20796_ (.B(_11698_),
    .C(_11667_),
    .A(_11697_),
    .Y(_11701_));
 sg13g2_nand2_1 _20797_ (.Y(_11702_),
    .A(_11700_),
    .B(_11701_));
 sg13g2_nand3_1 _20798_ (.B(_10974_),
    .C(_11702_),
    .A(_10972_),
    .Y(_11703_));
 sg13g2_nand2_2 _20799_ (.Y(_11704_),
    .A(_11693_),
    .B(_11692_));
 sg13g2_nor2_1 _20800_ (.A(_10962_),
    .B(_10964_),
    .Y(_11705_));
 sg13g2_xor2_1 _20801_ (.B(_11705_),
    .A(_11704_),
    .X(_11706_));
 sg13g2_nand2_1 _20802_ (.Y(_11707_),
    .A(_11703_),
    .B(_11706_));
 sg13g2_nand2_1 _20803_ (.Y(_11708_),
    .A(_10970_),
    .B(_10950_));
 sg13g2_nand3_1 _20804_ (.B(_10961_),
    .C(_10968_),
    .A(_10967_),
    .Y(_11709_));
 sg13g2_nand2b_1 _20805_ (.Y(_11710_),
    .B(_11699_),
    .A_N(_11685_));
 sg13g2_nand3_1 _20806_ (.B(_11686_),
    .C(_11698_),
    .A(_11697_),
    .Y(_11711_));
 sg13g2_nand2_1 _20807_ (.Y(_11712_),
    .A(_11710_),
    .B(_11711_));
 sg13g2_nand3_1 _20808_ (.B(_11709_),
    .C(_11712_),
    .A(_11708_),
    .Y(_11713_));
 sg13g2_nand2_1 _20809_ (.Y(_11714_),
    .A(_10970_),
    .B(_10958_));
 sg13g2_nand3_1 _20810_ (.B(_10953_),
    .C(_10968_),
    .A(_10967_),
    .Y(_11715_));
 sg13g2_nand2_1 _20811_ (.Y(_11716_),
    .A(_11699_),
    .B(_11685_));
 sg13g2_nand3_1 _20812_ (.B(_11682_),
    .C(_11698_),
    .A(_11697_),
    .Y(_11717_));
 sg13g2_nand2_1 _20813_ (.Y(_11718_),
    .A(_11716_),
    .B(_11717_));
 sg13g2_nand3_1 _20814_ (.B(_11715_),
    .C(_11718_),
    .A(_11714_),
    .Y(_11719_));
 sg13g2_nand2_1 _20815_ (.Y(_11720_),
    .A(_11713_),
    .B(_11719_));
 sg13g2_nor2_1 _20816_ (.A(_11707_),
    .B(_11720_),
    .Y(_11721_));
 sg13g2_a21oi_1 _20817_ (.A1(_10972_),
    .A2(_10974_),
    .Y(_11722_),
    .B1(_11702_));
 sg13g2_nand2_1 _20818_ (.Y(_11723_),
    .A(_11721_),
    .B(_11722_));
 sg13g2_nor2b_1 _20819_ (.A(_11713_),
    .B_N(_11706_),
    .Y(_11724_));
 sg13g2_a21oi_1 _20820_ (.A1(_11704_),
    .A2(_11705_),
    .Y(_11725_),
    .B1(_11724_));
 sg13g2_nand2_1 _20821_ (.Y(_11726_),
    .A(_11723_),
    .B(_11725_));
 sg13g2_buf_8 _20822_ (.A(_11726_),
    .X(_11727_));
 sg13g2_nand2_1 _20823_ (.Y(_11728_),
    .A(_11727_),
    .B(_11702_));
 sg13g2_nand2_1 _20824_ (.Y(_11729_),
    .A(_10972_),
    .B(_10974_));
 sg13g2_nand3_1 _20825_ (.B(_11729_),
    .C(_11725_),
    .A(_11723_),
    .Y(_11730_));
 sg13g2_buf_1 _20826_ (.A(_11730_),
    .X(_11731_));
 sg13g2_nor2_1 _20827_ (.A(_05015_),
    .B(_07912_),
    .Y(_11732_));
 sg13g2_nor2_1 _20828_ (.A(_10324_),
    .B(_07902_),
    .Y(_11733_));
 sg13g2_nor2_1 _20829_ (.A(_05019_),
    .B(_05815_),
    .Y(_11734_));
 sg13g2_nand4_1 _20830_ (.B(_10392_),
    .C(_11733_),
    .A(_11732_),
    .Y(_11735_),
    .D(_11734_));
 sg13g2_inv_1 _20831_ (.Y(_11736_),
    .A(_04878_));
 sg13g2_inv_1 _20832_ (.Y(_11737_),
    .A(_09358_));
 sg13g2_nand2_1 _20833_ (.Y(_11738_),
    .A(_09365_),
    .B(_09366_));
 sg13g2_inv_1 _20834_ (.Y(_11739_),
    .A(_09077_));
 sg13g2_nand2_1 _20835_ (.Y(_11740_),
    .A(_08343_),
    .B(_11739_));
 sg13g2_o21ai_1 _20836_ (.B1(_11740_),
    .Y(_11741_),
    .A1(_05958_),
    .A2(_05912_));
 sg13g2_a221oi_1 _20837_ (.B2(_11738_),
    .C1(_11741_),
    .B1(_11737_),
    .A1(_11736_),
    .Y(_11742_),
    .A2(_04963_));
 sg13g2_a22oi_1 _20838_ (.Y(_11743_),
    .B1(_09695_),
    .B2(_09701_),
    .A2(_06590_),
    .A1(_06813_));
 sg13g2_a21oi_1 _20839_ (.A1(_08071_),
    .A2(net51),
    .Y(_11744_),
    .B1(_06433_));
 sg13g2_a21oi_1 _20840_ (.A1(_06069_),
    .A2(net53),
    .Y(_11745_),
    .B1(_05657_));
 sg13g2_inv_1 _20841_ (.Y(_11746_),
    .A(_11745_));
 sg13g2_a21oi_1 _20842_ (.A1(_11746_),
    .A2(net51),
    .Y(_11747_),
    .B1(_06402_));
 sg13g2_a21oi_1 _20843_ (.A1(_04153_),
    .A2(_07531_),
    .Y(_11748_),
    .B1(_04309_));
 sg13g2_o21ai_1 _20844_ (.B1(_07113_),
    .Y(_11749_),
    .A1(_06184_),
    .A2(_11748_));
 sg13g2_buf_1 _20845_ (.A(_11749_),
    .X(_11750_));
 sg13g2_a21oi_2 _20846_ (.B1(_06979_),
    .Y(_11751_),
    .A2(net55),
    .A1(_11750_));
 sg13g2_a22oi_1 _20847_ (.Y(_11752_),
    .B1(_11751_),
    .B2(_07713_),
    .A2(_11747_),
    .A1(_11744_));
 sg13g2_nand3_1 _20848_ (.B(_11743_),
    .C(_11752_),
    .A(_11742_),
    .Y(_11753_));
 sg13g2_inv_1 _20849_ (.Y(_11754_),
    .A(_07983_));
 sg13g2_nand3_1 _20850_ (.B(_08459_),
    .C(_09486_),
    .A(_09612_),
    .Y(_11755_));
 sg13g2_nor3_1 _20851_ (.A(_08360_),
    .B(_09118_),
    .C(_11755_),
    .Y(_11756_));
 sg13g2_nand4_1 _20852_ (.B(_11754_),
    .C(_08463_),
    .A(_07810_),
    .Y(_11757_),
    .D(_11756_));
 sg13g2_nor3_1 _20853_ (.A(_11735_),
    .B(_11753_),
    .C(_11757_),
    .Y(_11758_));
 sg13g2_nand2_1 _20854_ (.Y(_11759_),
    .A(_07986_),
    .B(_11737_));
 sg13g2_o21ai_1 _20855_ (.B1(_11759_),
    .Y(_11760_),
    .A1(_05957_),
    .A2(_05912_));
 sg13g2_a22oi_1 _20856_ (.Y(_11761_),
    .B1(_11736_),
    .B2(_04964_),
    .A2(_11739_),
    .A1(_09141_));
 sg13g2_nor2b_1 _20857_ (.A(_11760_),
    .B_N(_11761_),
    .Y(_11762_));
 sg13g2_inv_1 _20858_ (.Y(_11763_),
    .A(_11762_));
 sg13g2_inv_1 _20859_ (.Y(_11764_),
    .A(_07713_));
 sg13g2_a22oi_1 _20860_ (.Y(_11765_),
    .B1(_09695_),
    .B2(_09702_),
    .A2(_11751_),
    .A1(_11764_));
 sg13g2_inv_1 _20861_ (.Y(_11766_),
    .A(_11744_));
 sg13g2_a22oi_1 _20862_ (.Y(_11767_),
    .B1(_06814_),
    .B2(_06590_),
    .A2(_11747_),
    .A1(_11766_));
 sg13g2_nand2_1 _20863_ (.Y(_11768_),
    .A(_11765_),
    .B(_11767_));
 sg13g2_nor3_1 _20864_ (.A(_05828_),
    .B(_07936_),
    .C(_10349_),
    .Y(_11769_));
 sg13g2_nor2_1 _20865_ (.A(_04528_),
    .B(_05829_),
    .Y(_11770_));
 sg13g2_nand3_1 _20866_ (.B(_11770_),
    .C(_11027_),
    .A(_11769_),
    .Y(_11771_));
 sg13g2_nor4_1 _20867_ (.A(_08345_),
    .B(_09106_),
    .C(_09544_),
    .D(_08608_),
    .Y(_11772_));
 sg13g2_inv_1 _20868_ (.Y(_11773_),
    .A(_09721_));
 sg13g2_or2_1 _20869_ (.X(_11774_),
    .B(_11738_),
    .A(_07705_));
 sg13g2_nand4_1 _20870_ (.B(_08442_),
    .C(_11773_),
    .A(_11772_),
    .Y(_11775_),
    .D(_11774_));
 sg13g2_nor4_1 _20871_ (.A(_11763_),
    .B(_11768_),
    .C(_11771_),
    .D(_11775_),
    .Y(_11776_));
 sg13g2_nor3_1 _20872_ (.A(_04887_),
    .B(_11758_),
    .C(_11776_),
    .Y(_11777_));
 sg13g2_nand2_1 _20873_ (.Y(_11778_),
    .A(_11777_),
    .B(net162));
 sg13g2_nand2_1 _20874_ (.Y(_11779_),
    .A(_11776_),
    .B(_11758_));
 sg13g2_nand3_1 _20875_ (.B(net129),
    .C(_04903_),
    .A(_11779_),
    .Y(_11780_));
 sg13g2_nand2_1 _20876_ (.Y(_11781_),
    .A(_11778_),
    .B(_11780_));
 sg13g2_nand2_1 _20877_ (.Y(_11782_),
    .A(_11778_),
    .B(_04884_));
 sg13g2_nand2b_1 _20878_ (.Y(_11783_),
    .B(_04883_),
    .A_N(_04900_));
 sg13g2_nand3_1 _20879_ (.B(_11782_),
    .C(_11783_),
    .A(_11781_),
    .Y(_11784_));
 sg13g2_nand2_1 _20880_ (.Y(_11785_),
    .A(_11743_),
    .B(_11752_));
 sg13g2_o21ai_1 _20881_ (.B1(_04887_),
    .Y(_11786_),
    .A1(_11785_),
    .A2(_11768_));
 sg13g2_nor3_1 _20882_ (.A(_04879_),
    .B(_04883_),
    .C(_11786_),
    .Y(_11787_));
 sg13g2_a21o_1 _20883_ (.A2(_11762_),
    .A1(_11742_),
    .B1(_04903_),
    .X(_11788_));
 sg13g2_a21o_1 _20884_ (.A2(_11788_),
    .A1(_11786_),
    .B1(_04901_),
    .X(_11789_));
 sg13g2_buf_1 _20885_ (.A(_11789_),
    .X(_11790_));
 sg13g2_nand2b_1 _20886_ (.Y(_11791_),
    .B(_11790_),
    .A_N(_11787_));
 sg13g2_nand2_1 _20887_ (.Y(_11792_),
    .A(_11791_),
    .B(net112));
 sg13g2_nand2_1 _20888_ (.Y(_11793_),
    .A(_11784_),
    .B(_11792_));
 sg13g2_buf_1 _20889_ (.A(\b.gen_square[27].sq.mask ),
    .X(_11794_));
 sg13g2_nand2_1 _20890_ (.Y(_11795_),
    .A(_11793_),
    .B(_11794_));
 sg13g2_inv_1 _20891_ (.Y(_11796_),
    .A(_11795_));
 sg13g2_nand2_1 _20892_ (.Y(_11797_),
    .A(_07182_),
    .B(_09196_));
 sg13g2_nand2_1 _20893_ (.Y(_11798_),
    .A(_11797_),
    .B(_08549_));
 sg13g2_nor3_1 _20894_ (.A(_08102_),
    .B(_11798_),
    .C(_09721_),
    .Y(_11799_));
 sg13g2_nand2_1 _20895_ (.Y(_11800_),
    .A(_09189_),
    .B(_09190_));
 sg13g2_nor2_1 _20896_ (.A(_07972_),
    .B(_11800_),
    .Y(_11801_));
 sg13g2_inv_1 _20897_ (.Y(_11802_),
    .A(_11801_));
 sg13g2_nand4_1 _20898_ (.B(_08447_),
    .C(_11802_),
    .A(_11799_),
    .Y(_11803_),
    .D(_09545_));
 sg13g2_a22oi_1 _20899_ (.Y(_11804_),
    .B1(_07197_),
    .B2(_07182_),
    .A2(_09827_),
    .A1(_08059_));
 sg13g2_inv_1 _20900_ (.Y(_11805_),
    .A(_11804_));
 sg13g2_inv_1 _20901_ (.Y(_11806_),
    .A(_08289_));
 sg13g2_inv_1 _20902_ (.Y(_11807_),
    .A(_09208_));
 sg13g2_nand2_1 _20903_ (.Y(_11808_),
    .A(_11807_),
    .B(_07981_));
 sg13g2_o21ai_1 _20904_ (.B1(_11808_),
    .Y(_11809_),
    .A1(_08330_),
    .A2(_11806_));
 sg13g2_nor2_1 _20905_ (.A(_11805_),
    .B(_11809_),
    .Y(_11810_));
 sg13g2_or2_1 _20906_ (.X(_11811_),
    .B(_05183_),
    .A(_06620_));
 sg13g2_nand3b_1 _20907_ (.B(_10467_),
    .C(_09009_),
    .Y(_11812_),
    .A_N(_10616_));
 sg13g2_nor4_1 _20908_ (.A(_11811_),
    .B(_06641_),
    .C(_05163_),
    .D(_11812_),
    .Y(_11813_));
 sg13g2_nand2_1 _20909_ (.Y(_11814_),
    .A(_11810_),
    .B(_11813_));
 sg13g2_nor2_1 _20910_ (.A(_09581_),
    .B(_09585_),
    .Y(_11815_));
 sg13g2_a22oi_1 _20911_ (.Y(_11816_),
    .B1(_06371_),
    .B2(_06430_),
    .A2(_11745_),
    .A1(_08071_));
 sg13g2_inv_1 _20912_ (.Y(_11817_),
    .A(_11816_));
 sg13g2_o21ai_1 _20913_ (.B1(_06595_),
    .Y(_11818_),
    .A1(_09368_),
    .A2(_11751_));
 sg13g2_buf_1 _20914_ (.A(_11818_),
    .X(_11819_));
 sg13g2_o21ai_1 _20915_ (.B1(_07988_),
    .Y(_11820_),
    .A1(_09368_),
    .A2(_07713_));
 sg13g2_inv_1 _20916_ (.Y(_11821_),
    .A(_11820_));
 sg13g2_nor2_1 _20917_ (.A(_11819_),
    .B(_11821_),
    .Y(_11822_));
 sg13g2_nor3_1 _20918_ (.A(_11815_),
    .B(_11817_),
    .C(_11822_),
    .Y(_11823_));
 sg13g2_inv_1 _20919_ (.Y(_11824_),
    .A(_11823_));
 sg13g2_nor4_1 _20920_ (.A(_07967_),
    .B(_11803_),
    .C(_11814_),
    .D(_11824_),
    .Y(_11825_));
 sg13g2_a22oi_1 _20921_ (.Y(_11826_),
    .B1(_08330_),
    .B2(_08289_),
    .A2(_11800_),
    .A1(_11807_));
 sg13g2_a22oi_1 _20922_ (.Y(_11827_),
    .B1(_07197_),
    .B2(_07181_),
    .A2(_09827_),
    .A1(_08058_));
 sg13g2_nand2_1 _20923_ (.Y(_11828_),
    .A(_11826_),
    .B(_11827_));
 sg13g2_nand2b_1 _20924_ (.Y(_11829_),
    .B(_11821_),
    .A_N(_11819_));
 sg13g2_a22oi_1 _20925_ (.Y(_11830_),
    .B1(_06371_),
    .B2(_06429_),
    .A2(_11745_),
    .A1(_08070_));
 sg13g2_nand2b_1 _20926_ (.Y(_11831_),
    .B(_09581_),
    .A_N(_09585_));
 sg13g2_nand3_1 _20927_ (.B(_11830_),
    .C(_11831_),
    .A(_11829_),
    .Y(_11832_));
 sg13g2_nor2_1 _20928_ (.A(_11828_),
    .B(_11832_),
    .Y(_11833_));
 sg13g2_nor2_1 _20929_ (.A(_05204_),
    .B(_06646_),
    .Y(_11834_));
 sg13g2_inv_1 _20930_ (.Y(_11835_),
    .A(_11834_));
 sg13g2_nor2_1 _20931_ (.A(_05208_),
    .B(_10171_),
    .Y(_11836_));
 sg13g2_inv_1 _20932_ (.Y(_11837_),
    .A(_11836_));
 sg13g2_nor2_1 _20933_ (.A(_08273_),
    .B(_07838_),
    .Y(_11838_));
 sg13g2_nor2_1 _20934_ (.A(_06651_),
    .B(_10632_),
    .Y(_11839_));
 sg13g2_nand2_1 _20935_ (.Y(_11840_),
    .A(_11838_),
    .B(_11839_));
 sg13g2_nor3_1 _20936_ (.A(_11835_),
    .B(_11837_),
    .C(_11840_),
    .Y(_11841_));
 sg13g2_nor3_1 _20937_ (.A(_09275_),
    .B(_08061_),
    .C(_08072_),
    .Y(_11842_));
 sg13g2_nand3_1 _20938_ (.B(_09612_),
    .C(_11842_),
    .A(_09486_),
    .Y(_11843_));
 sg13g2_nor4_1 _20939_ (.A(_07983_),
    .B(_08360_),
    .C(_07990_),
    .D(_11843_),
    .Y(_11844_));
 sg13g2_and3_1 _20940_ (.X(_11845_),
    .A(_11833_),
    .B(_11841_),
    .C(_11844_));
 sg13g2_nor3_1 _20941_ (.A(net127),
    .B(_11825_),
    .C(_11845_),
    .Y(_11846_));
 sg13g2_nand2_1 _20942_ (.Y(_11847_),
    .A(_11846_),
    .B(net191));
 sg13g2_nand2_1 _20943_ (.Y(_11848_),
    .A(_11845_),
    .B(_11825_));
 sg13g2_nand3_1 _20944_ (.B(net144),
    .C(_06397_),
    .A(_11848_),
    .Y(_11849_));
 sg13g2_nand2_1 _20945_ (.Y(_11850_),
    .A(_11847_),
    .B(_11849_));
 sg13g2_nand2_1 _20946_ (.Y(_11851_),
    .A(_11847_),
    .B(_06378_));
 sg13g2_nand2b_1 _20947_ (.Y(_11852_),
    .B(_06377_),
    .A_N(_06393_));
 sg13g2_nand3_1 _20948_ (.B(_11851_),
    .C(_11852_),
    .A(_11850_),
    .Y(_11853_));
 sg13g2_o21ai_1 _20949_ (.B1(net127),
    .Y(_11854_),
    .A1(_11832_),
    .A2(_11824_));
 sg13g2_inv_1 _20950_ (.Y(_11855_),
    .A(_11810_));
 sg13g2_o21ai_1 _20951_ (.B1(net127),
    .Y(_11856_),
    .A1(_11828_),
    .A2(_11855_));
 sg13g2_a21o_1 _20952_ (.A2(_11856_),
    .A1(_11854_),
    .B1(_06394_),
    .X(_11857_));
 sg13g2_o21ai_1 _20953_ (.B1(_11857_),
    .Y(_11858_),
    .A1(_06396_),
    .A2(_11854_));
 sg13g2_nand2_1 _20954_ (.Y(_11859_),
    .A(_11858_),
    .B(_05109_));
 sg13g2_nand2_1 _20955_ (.Y(_11860_),
    .A(_11853_),
    .B(_11859_));
 sg13g2_buf_1 _20956_ (.A(\b.gen_square[26].sq.mask ),
    .X(_11861_));
 sg13g2_nand2_1 _20957_ (.Y(_11862_),
    .A(_11860_),
    .B(_11861_));
 sg13g2_inv_1 _20958_ (.Y(_11863_),
    .A(_11862_));
 sg13g2_o21ai_1 _20959_ (.B1(_06379_),
    .Y(_11864_),
    .A1(_06376_),
    .A2(_06381_));
 sg13g2_nand3_1 _20960_ (.B(net144),
    .C(_11864_),
    .A(_11848_),
    .Y(_11865_));
 sg13g2_o21ai_1 _20961_ (.B1(_11865_),
    .Y(_11866_),
    .A1(_06376_),
    .A2(_11847_));
 sg13g2_nor3_1 _20962_ (.A(_06384_),
    .B(_07967_),
    .C(_11803_),
    .Y(_11867_));
 sg13g2_a21oi_1 _20963_ (.A1(_11867_),
    .A2(_11844_),
    .Y(_11868_),
    .B1(net120));
 sg13g2_nand2b_1 _20964_ (.Y(_11869_),
    .B(_11868_),
    .A_N(_06385_));
 sg13g2_or2_1 _20965_ (.X(_11870_),
    .B(_11856_),
    .A(_07199_));
 sg13g2_nand3_1 _20966_ (.B(_06384_),
    .C(_11870_),
    .A(_11857_),
    .Y(_11871_));
 sg13g2_nor2b_1 _20967_ (.A(_11869_),
    .B_N(_11871_),
    .Y(_11872_));
 sg13g2_o21ai_1 _20968_ (.B1(_11861_),
    .Y(_11873_),
    .A1(_11866_),
    .A2(_11872_));
 sg13g2_inv_1 _20969_ (.Y(_11874_),
    .A(_11873_));
 sg13g2_buf_1 _20970_ (.A(\b.gen_square[24].sq.mask ),
    .X(_11875_));
 sg13g2_inv_1 _20971_ (.Y(_11876_),
    .A(_11875_));
 sg13g2_nor2_1 _20972_ (.A(_09183_),
    .B(_09174_),
    .Y(_11877_));
 sg13g2_a21oi_1 _20973_ (.A1(_11819_),
    .A2(net51),
    .Y(_11878_),
    .B1(_06402_));
 sg13g2_o21ai_1 _20974_ (.B1(_05656_),
    .Y(_11879_),
    .A1(_08155_),
    .A2(_11878_));
 sg13g2_a21oi_1 _20975_ (.A1(_11820_),
    .A2(net51),
    .Y(_11880_),
    .B1(_06433_));
 sg13g2_o21ai_1 _20976_ (.B1(_09339_),
    .Y(_11881_),
    .A1(_08155_),
    .A2(_11880_));
 sg13g2_nor2_1 _20977_ (.A(_11879_),
    .B(_11881_),
    .Y(_11882_));
 sg13g2_nor2_1 _20978_ (.A(_11877_),
    .B(_11882_),
    .Y(_11883_));
 sg13g2_nand2_1 _20979_ (.Y(_11884_),
    .A(_06040_),
    .B(_06108_));
 sg13g2_nor2_1 _20980_ (.A(_08061_),
    .B(_09308_),
    .Y(_11885_));
 sg13g2_inv_1 _20981_ (.Y(_11886_),
    .A(_08352_));
 sg13g2_nand3_1 _20982_ (.B(_11886_),
    .C(_11081_),
    .A(_11885_),
    .Y(_11887_));
 sg13g2_nor2_1 _20983_ (.A(_09275_),
    .B(_11887_),
    .Y(_11888_));
 sg13g2_a21oi_1 _20984_ (.A1(_09429_),
    .A2(_05710_),
    .Y(_11889_),
    .B1(_05713_));
 sg13g2_a21oi_1 _20985_ (.A1(_11197_),
    .A2(net38),
    .Y(_11890_),
    .B1(_07196_));
 sg13g2_inv_1 _20986_ (.Y(_11891_),
    .A(_08321_));
 sg13g2_a21oi_1 _20987_ (.A1(_11891_),
    .A2(_05677_),
    .Y(_11892_),
    .B1(_05723_));
 sg13g2_a21oi_1 _20988_ (.A1(_08294_),
    .A2(_05677_),
    .Y(_11893_),
    .B1(_06755_));
 sg13g2_nand3_1 _20989_ (.B(_05206_),
    .C(_09282_),
    .A(_11839_),
    .Y(_11894_));
 sg13g2_a221oi_1 _20990_ (.B2(_11893_),
    .C1(_11894_),
    .B1(_11892_),
    .A1(_11889_),
    .Y(_11895_),
    .A2(_11890_));
 sg13g2_nand4_1 _20991_ (.B(_11884_),
    .C(_11888_),
    .A(_11883_),
    .Y(_11896_),
    .D(_11895_));
 sg13g2_nand2b_1 _20992_ (.Y(_11897_),
    .B(_11893_),
    .A_N(_11892_));
 sg13g2_nor4_1 _20993_ (.A(_06620_),
    .B(_05146_),
    .C(_08265_),
    .D(_10616_),
    .Y(_11898_));
 sg13g2_inv_1 _20994_ (.Y(_11899_),
    .A(_11898_));
 sg13g2_nor2b_1 _20995_ (.A(_11889_),
    .B_N(_11890_),
    .Y(_11900_));
 sg13g2_a21oi_1 _20996_ (.A1(_06041_),
    .A2(_09264_),
    .Y(_11901_),
    .B1(_06108_));
 sg13g2_nor3_1 _20997_ (.A(_11899_),
    .B(_11900_),
    .C(_11901_),
    .Y(_11902_));
 sg13g2_inv_1 _20998_ (.Y(_11903_),
    .A(_11798_));
 sg13g2_nor2_1 _20999_ (.A(_08323_),
    .B(_08102_),
    .Y(_11904_));
 sg13g2_nand4_1 _21000_ (.B(_11902_),
    .C(_11903_),
    .A(_11897_),
    .Y(_11905_),
    .D(_11904_));
 sg13g2_nand2b_1 _21001_ (.Y(_11906_),
    .B(_11881_),
    .A_N(_11879_));
 sg13g2_nand2b_1 _21002_ (.Y(_11907_),
    .B(_09174_),
    .A_N(_09183_));
 sg13g2_nand3b_1 _21003_ (.B(_11906_),
    .C(_11907_),
    .Y(_11908_),
    .A_N(_11905_));
 sg13g2_nand4_1 _21004_ (.B(net215),
    .C(_06065_),
    .A(_11896_),
    .Y(_11909_),
    .D(_11908_));
 sg13g2_buf_1 _21005_ (.A(_11909_),
    .X(_11910_));
 sg13g2_nor2_1 _21006_ (.A(_06045_),
    .B(_11910_),
    .Y(_11911_));
 sg13g2_nor3_1 _21007_ (.A(_06047_),
    .B(_11798_),
    .C(_09265_),
    .Y(_11912_));
 sg13g2_and3_1 _21008_ (.X(_11913_),
    .A(_11888_),
    .B(_11904_),
    .C(_11912_));
 sg13g2_o21ai_1 _21009_ (.B1(_06049_),
    .Y(_11914_),
    .A1(_11890_),
    .A2(_11893_));
 sg13g2_nor2_1 _21010_ (.A(_06748_),
    .B(_11914_),
    .Y(_11915_));
 sg13g2_nand3_1 _21011_ (.B(_06041_),
    .C(_09183_),
    .A(_11879_),
    .Y(_11916_));
 sg13g2_nand2_1 _21012_ (.Y(_11917_),
    .A(_11916_),
    .B(_06049_));
 sg13g2_a21oi_1 _21013_ (.A1(_11917_),
    .A2(_11914_),
    .Y(_11918_),
    .B1(_06062_));
 sg13g2_nor3_1 _21014_ (.A(_08211_),
    .B(_11915_),
    .C(_11918_),
    .Y(_11919_));
 sg13g2_nor4_1 _21015_ (.A(net137),
    .B(_06050_),
    .C(_11913_),
    .D(_11919_),
    .Y(_11920_));
 sg13g2_nor2_1 _21016_ (.A(_06056_),
    .B(_06065_),
    .Y(_11921_));
 sg13g2_nor2b_1 _21017_ (.A(_06056_),
    .B_N(_06045_),
    .Y(_11922_));
 sg13g2_or2_1 _21018_ (.X(_11923_),
    .B(_11896_),
    .A(_11908_));
 sg13g2_buf_1 _21019_ (.A(_11923_),
    .X(_11924_));
 sg13g2_inv_1 _21020_ (.Y(_11925_),
    .A(_11924_));
 sg13g2_nor4_1 _21021_ (.A(_07381_),
    .B(_11921_),
    .C(_11922_),
    .D(_11925_),
    .Y(_11926_));
 sg13g2_nor3_1 _21022_ (.A(_11911_),
    .B(_11920_),
    .C(_11926_),
    .Y(_11927_));
 sg13g2_nor2_1 _21023_ (.A(_11876_),
    .B(_11927_),
    .Y(_11928_));
 sg13g2_nand2_1 _21024_ (.Y(_11929_),
    .A(_08206_),
    .B(_08170_));
 sg13g2_o21ai_1 _21025_ (.B1(_11929_),
    .Y(_11930_),
    .A1(_11127_),
    .A2(_11124_));
 sg13g2_nor2_1 _21026_ (.A(_06306_),
    .B(_06300_),
    .Y(_11931_));
 sg13g2_nor2_1 _21027_ (.A(_09413_),
    .B(_11931_),
    .Y(_11932_));
 sg13g2_nor2b_1 _21028_ (.A(_11930_),
    .B_N(_11932_),
    .Y(_11933_));
 sg13g2_nand2_1 _21029_ (.Y(_11934_),
    .A(_08207_),
    .B(_08170_));
 sg13g2_nor2_1 _21030_ (.A(_06306_),
    .B(_06114_),
    .Y(_11935_));
 sg13g2_nor2_1 _21031_ (.A(_09387_),
    .B(_11935_),
    .Y(_11936_));
 sg13g2_nand2_1 _21032_ (.Y(_11937_),
    .A(_11934_),
    .B(_11936_));
 sg13g2_a21oi_1 _21033_ (.A1(_11124_),
    .A2(_11126_),
    .Y(_11938_),
    .B1(_11937_));
 sg13g2_a21oi_1 _21034_ (.A1(_11933_),
    .A2(_11938_),
    .Y(_11939_),
    .B1(_05652_));
 sg13g2_inv_1 _21035_ (.Y(_11940_),
    .A(_09344_));
 sg13g2_inv_1 _21036_ (.Y(_11941_),
    .A(_11880_));
 sg13g2_nand2_1 _21037_ (.Y(_11942_),
    .A(_06070_),
    .B(_03611_));
 sg13g2_o21ai_1 _21038_ (.B1(_11942_),
    .Y(_11943_),
    .A1(_05628_),
    .A2(_05714_));
 sg13g2_a221oi_1 _21039_ (.B2(_11878_),
    .C1(_11943_),
    .B1(_11941_),
    .A1(_09337_),
    .Y(_11944_),
    .A2(_11940_));
 sg13g2_inv_1 _21040_ (.Y(_11945_),
    .A(_09337_));
 sg13g2_a22oi_1 _21041_ (.Y(_11946_),
    .B1(_11878_),
    .B2(_11880_),
    .A2(_11940_),
    .A1(_11945_));
 sg13g2_inv_1 _21042_ (.Y(_11947_),
    .A(_05628_));
 sg13g2_a22oi_1 _21043_ (.Y(_11948_),
    .B1(_11947_),
    .B2(_05714_),
    .A2(_06742_),
    .A1(_06070_));
 sg13g2_and2_1 _21044_ (.A(_11946_),
    .B(_11948_),
    .X(_11949_));
 sg13g2_a21oi_1 _21045_ (.A1(_11944_),
    .A2(_11949_),
    .Y(_11950_),
    .B1(_05652_));
 sg13g2_o21ai_1 _21046_ (.B1(_05650_),
    .Y(_11951_),
    .A1(_11939_),
    .A2(_11950_));
 sg13g2_nand2_1 _21047_ (.Y(_11952_),
    .A(_11950_),
    .B(_05651_));
 sg13g2_a21oi_1 _21048_ (.A1(_11951_),
    .A2(_11952_),
    .Y(_11953_),
    .B1(net137));
 sg13g2_nand2_1 _21049_ (.Y(_11954_),
    .A(_05652_),
    .B(net176));
 sg13g2_nor4_1 _21050_ (.A(_08061_),
    .B(_09275_),
    .C(_08360_),
    .D(_08065_),
    .Y(_11955_));
 sg13g2_nand2_1 _21051_ (.Y(_11956_),
    .A(_09486_),
    .B(_11886_));
 sg13g2_nor2_1 _21052_ (.A(_06464_),
    .B(_07912_),
    .Y(_11957_));
 sg13g2_inv_1 _21053_ (.Y(_11958_),
    .A(_11957_));
 sg13g2_nor3_1 _21054_ (.A(_11100_),
    .B(_11958_),
    .C(_10240_),
    .Y(_11959_));
 sg13g2_nor2_1 _21055_ (.A(_09417_),
    .B(_08351_),
    .Y(_11960_));
 sg13g2_nand3_1 _21056_ (.B(_11959_),
    .C(_11960_),
    .A(_11948_),
    .Y(_11961_));
 sg13g2_nor2_1 _21057_ (.A(_11956_),
    .B(_11961_),
    .Y(_11962_));
 sg13g2_nand4_1 _21058_ (.B(_11933_),
    .C(_11955_),
    .A(_11946_),
    .Y(_11963_),
    .D(_11962_));
 sg13g2_nor4_1 _21059_ (.A(_06289_),
    .B(_05829_),
    .C(_10217_),
    .D(_11093_),
    .Y(_11964_));
 sg13g2_nor2_1 _21060_ (.A(_08323_),
    .B(_09544_),
    .Y(_11965_));
 sg13g2_nor2_1 _21061_ (.A(_09391_),
    .B(_08324_),
    .Y(_11966_));
 sg13g2_nand4_1 _21062_ (.B(_11964_),
    .C(_11965_),
    .A(_11938_),
    .Y(_11967_),
    .D(_11966_));
 sg13g2_nor3_1 _21063_ (.A(_11798_),
    .B(_08345_),
    .C(_08096_),
    .Y(_11968_));
 sg13g2_nand3b_1 _21064_ (.B(_11944_),
    .C(_11968_),
    .Y(_11969_),
    .A_N(_11967_));
 sg13g2_or2_1 _21065_ (.X(_11970_),
    .B(_11969_),
    .A(_11963_));
 sg13g2_buf_1 _21066_ (.A(_11970_),
    .X(_11971_));
 sg13g2_inv_1 _21067_ (.Y(_11972_),
    .A(_11971_));
 sg13g2_nand4_1 _21068_ (.B(net215),
    .C(_05652_),
    .A(_11969_),
    .Y(_11973_),
    .D(_11963_));
 sg13g2_buf_1 _21069_ (.A(_11973_),
    .X(_11974_));
 sg13g2_o21ai_1 _21070_ (.B1(_11974_),
    .Y(_11975_),
    .A1(_11954_),
    .A2(_11972_));
 sg13g2_nand2_1 _21071_ (.Y(_11976_),
    .A(_11974_),
    .B(_05634_));
 sg13g2_nand2_1 _21072_ (.Y(_11977_),
    .A(_05649_),
    .B(_05633_));
 sg13g2_nand3_1 _21073_ (.B(_11976_),
    .C(_11977_),
    .A(_11975_),
    .Y(_11978_));
 sg13g2_nand2b_1 _21074_ (.Y(_11979_),
    .B(_11978_),
    .A_N(_11953_));
 sg13g2_buf_1 _21075_ (.A(\b.gen_square[25].sq.mask ),
    .X(_11980_));
 sg13g2_nand2_1 _21076_ (.Y(_11981_),
    .A(_11979_),
    .B(_11980_));
 sg13g2_a22oi_1 _21077_ (.Y(_11982_),
    .B1(_06056_),
    .B2(_11910_),
    .A2(_06055_),
    .A1(_06060_));
 sg13g2_nand3_1 _21078_ (.B(net176),
    .C(_06065_),
    .A(_11924_),
    .Y(_11983_));
 sg13g2_nand2_1 _21079_ (.Y(_11984_),
    .A(_11983_),
    .B(_11910_));
 sg13g2_inv_1 _21080_ (.Y(_11985_),
    .A(_11918_));
 sg13g2_o21ai_1 _21081_ (.B1(_11985_),
    .Y(_11986_),
    .A1(_06064_),
    .A2(_11917_));
 sg13g2_nor2b_1 _21082_ (.A(net137),
    .B_N(_11986_),
    .Y(_11987_));
 sg13g2_a21o_1 _21083_ (.A2(_11984_),
    .A1(_11982_),
    .B1(_11987_),
    .X(_11988_));
 sg13g2_nand2_1 _21084_ (.Y(_11989_),
    .A(_11988_),
    .B(_11875_));
 sg13g2_xnor2_1 _21085_ (.Y(_11990_),
    .A(_11981_),
    .B(_11989_));
 sg13g2_nor2_1 _21086_ (.A(_05629_),
    .B(_05648_),
    .Y(_11991_));
 sg13g2_o21ai_1 _21087_ (.B1(_11975_),
    .Y(_11992_),
    .A1(_05650_),
    .A2(_11991_));
 sg13g2_nand2_1 _21088_ (.Y(_11993_),
    .A(_11939_),
    .B(_06877_));
 sg13g2_a21o_1 _21089_ (.A2(_11959_),
    .A1(_11964_),
    .B1(_08415_),
    .X(_11994_));
 sg13g2_nand4_1 _21090_ (.B(_11952_),
    .C(_11993_),
    .A(_11951_),
    .Y(_11995_),
    .D(_11994_));
 sg13g2_nand2_1 _21091_ (.Y(_11996_),
    .A(_11995_),
    .B(net160));
 sg13g2_nand2_1 _21092_ (.Y(_11997_),
    .A(_11992_),
    .B(_11996_));
 sg13g2_nand2_1 _21093_ (.Y(_11998_),
    .A(_11997_),
    .B(_11980_));
 sg13g2_nor2_1 _21094_ (.A(_06044_),
    .B(_06059_),
    .Y(_11999_));
 sg13g2_o21ai_1 _21095_ (.B1(_11984_),
    .Y(_12000_),
    .A1(_06061_),
    .A2(_11999_));
 sg13g2_o21ai_1 _21096_ (.B1(_08050_),
    .Y(_12001_),
    .A1(_11894_),
    .A2(_11899_));
 sg13g2_o21ai_1 _21097_ (.B1(_12001_),
    .Y(_12002_),
    .A1(_06748_),
    .A2(_11914_));
 sg13g2_o21ai_1 _21098_ (.B1(net160),
    .Y(_12003_),
    .A1(_12002_),
    .A2(_11986_));
 sg13g2_a21oi_1 _21099_ (.A1(_12000_),
    .A2(_12003_),
    .Y(_12004_),
    .B1(_11876_));
 sg13g2_nor2_1 _21100_ (.A(_11998_),
    .B(_12004_),
    .Y(_12005_));
 sg13g2_nand2_1 _21101_ (.Y(_12006_),
    .A(_12004_),
    .B(_11998_));
 sg13g2_nor2b_1 _21102_ (.A(_12005_),
    .B_N(_12006_),
    .Y(_12007_));
 sg13g2_nand3_1 _21103_ (.B(_05640_),
    .C(_11993_),
    .A(_11951_),
    .Y(_12008_));
 sg13g2_nand4_1 _21104_ (.B(_05639_),
    .C(_08213_),
    .A(_11965_),
    .Y(_12009_),
    .D(_09264_));
 sg13g2_nor2_1 _21105_ (.A(_11956_),
    .B(_12009_),
    .Y(_12010_));
 sg13g2_nand3_1 _21106_ (.B(_11955_),
    .C(_11968_),
    .A(_12010_),
    .Y(_12011_));
 sg13g2_nor2_1 _21107_ (.A(net137),
    .B(_05641_),
    .Y(_12012_));
 sg13g2_nand3_1 _21108_ (.B(_12011_),
    .C(_12012_),
    .A(_12008_),
    .Y(_12013_));
 sg13g2_o21ai_1 _21109_ (.B1(_05635_),
    .Y(_12014_),
    .A1(_05632_),
    .A2(_05637_));
 sg13g2_nand3_1 _21110_ (.B(net161),
    .C(_12014_),
    .A(_11971_),
    .Y(_12015_));
 sg13g2_nand2b_1 _21111_ (.Y(_12016_),
    .B(_05638_),
    .A_N(_11974_));
 sg13g2_nand3_1 _21112_ (.B(_12015_),
    .C(_12016_),
    .A(_12013_),
    .Y(_12017_));
 sg13g2_nand2_1 _21113_ (.Y(_12018_),
    .A(_12017_),
    .B(_11980_));
 sg13g2_nand2_1 _21114_ (.Y(_12019_),
    .A(_12018_),
    .B(_11928_));
 sg13g2_nand3_1 _21115_ (.B(_12007_),
    .C(_12019_),
    .A(_11990_),
    .Y(_12020_));
 sg13g2_nor2_1 _21116_ (.A(_11928_),
    .B(_12018_),
    .Y(_12021_));
 sg13g2_a21oi_1 _21117_ (.A1(_11988_),
    .A2(_11875_),
    .Y(_12022_),
    .B1(_11981_));
 sg13g2_a21oi_1 _21118_ (.A1(_12022_),
    .A2(_12006_),
    .Y(_12023_),
    .B1(_12005_));
 sg13g2_nand2_1 _21119_ (.Y(_00632_),
    .A(_12020_),
    .B(_12023_));
 sg13g2_o21ai_1 _21120_ (.B1(_00632_),
    .Y(_00633_),
    .A1(_12020_),
    .A2(_12021_));
 sg13g2_buf_1 _21121_ (.A(_00633_),
    .X(_00634_));
 sg13g2_nor2_1 _21122_ (.A(_12018_),
    .B(_00634_),
    .Y(_00635_));
 sg13g2_a21oi_1 _21123_ (.A1(_11928_),
    .A2(_00634_),
    .Y(_00636_),
    .B1(_00635_));
 sg13g2_nor2b_1 _21124_ (.A(_00634_),
    .B_N(_11981_),
    .Y(_00637_));
 sg13g2_a21o_1 _21125_ (.A2(_00634_),
    .A1(_11989_),
    .B1(_00637_),
    .X(_00638_));
 sg13g2_buf_1 _21126_ (.A(_00638_),
    .X(_00639_));
 sg13g2_a22oi_1 _21127_ (.Y(_00640_),
    .B1(_11863_),
    .B2(_00639_),
    .A2(_00636_),
    .A1(_11874_));
 sg13g2_nor2_1 _21128_ (.A(net120),
    .B(_06383_),
    .Y(_00641_));
 sg13g2_a21o_1 _21129_ (.A2(_11841_),
    .A1(_11813_),
    .B1(_07921_),
    .X(_00642_));
 sg13g2_nand2_1 _21130_ (.Y(_00643_),
    .A(_11870_),
    .B(_00642_));
 sg13g2_xnor2_1 _21131_ (.Y(_00644_),
    .A(_06373_),
    .B(_06393_));
 sg13g2_a22oi_1 _21132_ (.Y(_00645_),
    .B1(_00644_),
    .B2(_11850_),
    .A2(_00643_),
    .A1(_00641_));
 sg13g2_nand2_1 _21133_ (.Y(_00646_),
    .A(_00645_),
    .B(_11859_));
 sg13g2_nand2_1 _21134_ (.Y(_00647_),
    .A(_00646_),
    .B(_11861_));
 sg13g2_nand2b_1 _21135_ (.Y(_00648_),
    .B(_11998_),
    .A_N(_12004_));
 sg13g2_inv_1 _21136_ (.Y(_00649_),
    .A(_00639_));
 sg13g2_a22oi_1 _21137_ (.Y(_00650_),
    .B1(_11862_),
    .B2(_00649_),
    .A2(_00648_),
    .A1(_00647_));
 sg13g2_nand2b_1 _21138_ (.Y(_00651_),
    .B(_00650_),
    .A_N(_00640_));
 sg13g2_inv_1 _21139_ (.Y(_00652_),
    .A(_00647_));
 sg13g2_nand2b_1 _21140_ (.Y(_00653_),
    .B(_00652_),
    .A_N(_00648_));
 sg13g2_nand2_1 _21141_ (.Y(_00654_),
    .A(_00651_),
    .B(_00653_));
 sg13g2_buf_2 _21142_ (.A(_00654_),
    .X(_00655_));
 sg13g2_nor2_1 _21143_ (.A(_00639_),
    .B(_00655_),
    .Y(_00656_));
 sg13g2_a21oi_1 _21144_ (.A1(_11863_),
    .A2(_00655_),
    .Y(_00657_),
    .B1(_00656_));
 sg13g2_nand3_1 _21145_ (.B(net162),
    .C(_04888_),
    .A(_11777_),
    .Y(_00658_));
 sg13g2_nand2b_1 _21146_ (.Y(_00659_),
    .B(_04899_),
    .A_N(_11788_));
 sg13g2_nand3_1 _21147_ (.B(_04890_),
    .C(_00659_),
    .A(_11790_),
    .Y(_00660_));
 sg13g2_inv_1 _21148_ (.Y(_00661_),
    .A(_04891_));
 sg13g2_nor2_1 _21149_ (.A(_11775_),
    .B(_11757_),
    .Y(_00662_));
 sg13g2_a21oi_1 _21150_ (.A1(_00662_),
    .A2(_04889_),
    .Y(_00663_),
    .B1(_02067_));
 sg13g2_nand3_1 _21151_ (.B(_00661_),
    .C(_00663_),
    .A(_00660_),
    .Y(_00664_));
 sg13g2_o21ai_1 _21152_ (.B1(_04885_),
    .Y(_00665_),
    .A1(_04882_),
    .A2(_04887_));
 sg13g2_nand3_1 _21153_ (.B(_05086_),
    .C(_00665_),
    .A(_11779_),
    .Y(_00666_));
 sg13g2_nand3_1 _21154_ (.B(_00664_),
    .C(_00666_),
    .A(_00658_),
    .Y(_00667_));
 sg13g2_nand2_1 _21155_ (.Y(_00668_),
    .A(_00667_),
    .B(_11794_));
 sg13g2_nand2_1 _21156_ (.Y(_00669_),
    .A(_00655_),
    .B(_11874_));
 sg13g2_o21ai_1 _21157_ (.B1(_00669_),
    .Y(_00670_),
    .A1(_00636_),
    .A2(_00655_));
 sg13g2_nor2_1 _21158_ (.A(_00668_),
    .B(_00670_),
    .Y(_00671_));
 sg13g2_o21ai_1 _21159_ (.B1(_00671_),
    .Y(_00672_),
    .A1(_11796_),
    .A2(_00657_));
 sg13g2_nor2_1 _21160_ (.A(_00652_),
    .B(_00648_),
    .Y(_00673_));
 sg13g2_inv_1 _21161_ (.Y(_00674_),
    .A(_11794_));
 sg13g2_nor2b_1 _21162_ (.A(_11787_),
    .B_N(_00659_),
    .Y(_00675_));
 sg13g2_o21ai_1 _21163_ (.B1(_07756_),
    .Y(_00676_),
    .A1(_11735_),
    .A2(_11771_));
 sg13g2_nand3_1 _21164_ (.B(_11790_),
    .C(_00676_),
    .A(_00675_),
    .Y(_00677_));
 sg13g2_o21ai_1 _21165_ (.B1(_04880_),
    .Y(_00678_),
    .A1(_04881_),
    .A2(_04882_));
 sg13g2_a22oi_1 _21166_ (.Y(_00679_),
    .B1(_11780_),
    .B2(_11778_),
    .A2(_00678_),
    .A1(_04901_));
 sg13g2_a21oi_1 _21167_ (.A1(net112),
    .A2(_00677_),
    .Y(_00680_),
    .B1(_00679_));
 sg13g2_nor2_1 _21168_ (.A(_00674_),
    .B(_00680_),
    .Y(_00681_));
 sg13g2_a22oi_1 _21169_ (.Y(_00682_),
    .B1(_11796_),
    .B2(_00657_),
    .A2(_00681_),
    .A1(_00673_));
 sg13g2_nand2_1 _21170_ (.Y(_00683_),
    .A(_00672_),
    .B(_00682_));
 sg13g2_inv_1 _21171_ (.Y(_00684_),
    .A(_00673_));
 sg13g2_nand2b_1 _21172_ (.Y(_00685_),
    .B(_00684_),
    .A_N(_00681_));
 sg13g2_nand4_1 _21173_ (.B(_11794_),
    .C(_00685_),
    .A(_00683_),
    .Y(_00686_),
    .D(_00667_));
 sg13g2_nand2_1 _21174_ (.Y(_00687_),
    .A(_00683_),
    .B(_00685_));
 sg13g2_nand2_1 _21175_ (.Y(_00688_),
    .A(_00687_),
    .B(_00670_));
 sg13g2_nor2_1 _21176_ (.A(_08953_),
    .B(_08960_),
    .Y(_00689_));
 sg13g2_inv_1 _21177_ (.Y(_00690_),
    .A(_09565_));
 sg13g2_nand2_1 _21178_ (.Y(_00691_),
    .A(_09549_),
    .B(_09550_));
 sg13g2_nor2_1 _21179_ (.A(_05328_),
    .B(_05529_),
    .Y(_00692_));
 sg13g2_a221oi_1 _21180_ (.B2(_07591_),
    .C1(_00692_),
    .B1(_07600_),
    .A1(_00690_),
    .Y(_00693_),
    .A2(_00691_));
 sg13g2_nor2b_1 _21181_ (.A(_00689_),
    .B_N(_00693_),
    .Y(_00694_));
 sg13g2_inv_1 _21182_ (.Y(_00695_),
    .A(_00694_));
 sg13g2_nor2_1 _21183_ (.A(_11750_),
    .B(_07712_),
    .Y(_00696_));
 sg13g2_inv_1 _21184_ (.Y(_00697_),
    .A(_11747_));
 sg13g2_a21oi_1 _21185_ (.A1(_00697_),
    .A2(net42),
    .Y(_00698_),
    .B1(_06596_));
 sg13g2_a21oi_1 _21186_ (.A1(_11766_),
    .A2(_04898_),
    .Y(_00699_),
    .B1(_04967_));
 sg13g2_a22oi_1 _21187_ (.Y(_00700_),
    .B1(_00698_),
    .B2(_00699_),
    .A2(_06972_),
    .A1(_07005_));
 sg13g2_nand2b_1 _21188_ (.Y(_00701_),
    .B(_09811_),
    .A_N(_09816_));
 sg13g2_nand3b_1 _21189_ (.B(_00700_),
    .C(_00701_),
    .Y(_00702_),
    .A_N(_00696_));
 sg13g2_nor4_1 _21190_ (.A(_07815_),
    .B(_07990_),
    .C(_09118_),
    .D(_07809_),
    .Y(_00703_));
 sg13g2_nor2_1 _21191_ (.A(_07993_),
    .B(_09115_),
    .Y(_00704_));
 sg13g2_nand4_1 _21192_ (.B(_11754_),
    .C(_00704_),
    .A(_00703_),
    .Y(_00705_),
    .D(_09612_));
 sg13g2_nor3_1 _21193_ (.A(_00695_),
    .B(_00702_),
    .C(_00705_),
    .Y(_00706_));
 sg13g2_nand2_1 _21194_ (.Y(_00707_),
    .A(_05206_),
    .B(_09282_));
 sg13g2_nor4_1 _21195_ (.A(_08822_),
    .B(_11646_),
    .C(_00707_),
    .D(_11837_),
    .Y(_00708_));
 sg13g2_nand2_1 _21196_ (.Y(_00709_),
    .A(_00706_),
    .B(_00708_));
 sg13g2_nand2_1 _21197_ (.Y(_00710_),
    .A(_00690_),
    .B(_07804_));
 sg13g2_o21ai_1 _21198_ (.B1(_00710_),
    .Y(_00711_),
    .A1(_05328_),
    .A2(_05528_));
 sg13g2_nor3_1 _21199_ (.A(_06625_),
    .B(_05146_),
    .C(_08267_),
    .Y(_00712_));
 sg13g2_nand3_1 _21200_ (.B(_10123_),
    .C(_11629_),
    .A(_00712_),
    .Y(_00713_));
 sg13g2_nand2b_1 _21201_ (.Y(_00714_),
    .B(_07712_),
    .A_N(_11750_));
 sg13g2_o21ai_1 _21202_ (.B1(_00714_),
    .Y(_00715_),
    .A1(_06973_),
    .A2(_07005_));
 sg13g2_nand2_1 _21203_ (.Y(_00716_),
    .A(_07601_),
    .B(_07591_));
 sg13g2_o21ai_1 _21204_ (.B1(_00716_),
    .Y(_00717_),
    .A1(_07974_),
    .A2(_08953_));
 sg13g2_nor4_1 _21205_ (.A(_00711_),
    .B(_00713_),
    .C(_00715_),
    .D(_00717_),
    .Y(_00718_));
 sg13g2_nor4_1 _21206_ (.A(_09106_),
    .B(_09721_),
    .C(_07975_),
    .D(_07967_),
    .Y(_00719_));
 sg13g2_inv_1 _21207_ (.Y(_00720_),
    .A(_00698_));
 sg13g2_nor2_1 _21208_ (.A(_00699_),
    .B(_00720_),
    .Y(_00721_));
 sg13g2_inv_1 _21209_ (.Y(_00722_),
    .A(_07707_));
 sg13g2_nor2_1 _21210_ (.A(_07960_),
    .B(_00691_),
    .Y(_00723_));
 sg13g2_nor3_1 _21211_ (.A(_00723_),
    .B(_07704_),
    .C(_09103_),
    .Y(_00724_));
 sg13g2_nand2_1 _21212_ (.Y(_00725_),
    .A(_00722_),
    .B(_00724_));
 sg13g2_nor2_1 _21213_ (.A(_09816_),
    .B(_09811_),
    .Y(_00726_));
 sg13g2_nor3_1 _21214_ (.A(_00721_),
    .B(_00725_),
    .C(_00726_),
    .Y(_00727_));
 sg13g2_nand3_1 _21215_ (.B(_00719_),
    .C(_00727_),
    .A(_00718_),
    .Y(_00728_));
 sg13g2_nand4_1 _21216_ (.B(net162),
    .C(_05352_),
    .A(_00709_),
    .Y(_00729_),
    .D(_00728_));
 sg13g2_buf_1 _21217_ (.A(_00729_),
    .X(_00730_));
 sg13g2_nand2b_1 _21218_ (.Y(_00731_),
    .B(_05338_),
    .A_N(_00730_));
 sg13g2_nor2_1 _21219_ (.A(_05340_),
    .B(_00725_),
    .Y(_00732_));
 sg13g2_nand3b_1 _21220_ (.B(_00719_),
    .C(_00732_),
    .Y(_00733_),
    .A_N(_00705_));
 sg13g2_nand2b_1 _21221_ (.Y(_00734_),
    .B(_00694_),
    .A_N(_00711_));
 sg13g2_o21ai_1 _21222_ (.B1(_05337_),
    .Y(_00735_),
    .A1(_00717_),
    .A2(_00734_));
 sg13g2_or3_1 _21223_ (.A(_00715_),
    .B(_00721_),
    .C(_00726_),
    .X(_00736_));
 sg13g2_o21ai_1 _21224_ (.B1(_05337_),
    .Y(_00737_),
    .A1(_00736_),
    .A2(_00702_));
 sg13g2_a21o_1 _21225_ (.A2(_00737_),
    .A1(_00735_),
    .B1(_05350_),
    .X(_00738_));
 sg13g2_nor2b_1 _21226_ (.A(_00735_),
    .B_N(_05348_),
    .Y(_00739_));
 sg13g2_inv_1 _21227_ (.Y(_00740_),
    .A(_00739_));
 sg13g2_nand3_1 _21228_ (.B(_05340_),
    .C(_00740_),
    .A(_00738_),
    .Y(_00741_));
 sg13g2_inv_1 _21229_ (.Y(_00742_),
    .A(_05341_));
 sg13g2_nand4_1 _21230_ (.B(_00741_),
    .C(net112),
    .A(_00733_),
    .Y(_00743_),
    .D(_00742_));
 sg13g2_or2_1 _21231_ (.X(_00744_),
    .B(_00709_),
    .A(_00728_));
 sg13g2_buf_1 _21232_ (.A(_00744_),
    .X(_00745_));
 sg13g2_o21ai_1 _21233_ (.B1(_05335_),
    .Y(_00746_),
    .A1(_05332_),
    .A2(_05337_));
 sg13g2_nand3_1 _21234_ (.B(_05087_),
    .C(_00746_),
    .A(_00745_),
    .Y(_00747_));
 sg13g2_nand3_1 _21235_ (.B(_00743_),
    .C(_00747_),
    .A(_00731_),
    .Y(_00748_));
 sg13g2_buf_1 _21236_ (.A(\b.gen_square[28].sq.mask ),
    .X(_00749_));
 sg13g2_nand2_1 _21237_ (.Y(_00750_),
    .A(_00748_),
    .B(_00749_));
 sg13g2_inv_1 _21238_ (.Y(_00751_),
    .A(_00750_));
 sg13g2_nand3_1 _21239_ (.B(_00688_),
    .C(_00751_),
    .A(_00686_),
    .Y(_00752_));
 sg13g2_nand2b_1 _21240_ (.Y(_00753_),
    .B(_00687_),
    .A_N(_00657_));
 sg13g2_nand3_1 _21241_ (.B(_11796_),
    .C(_00685_),
    .A(_00683_),
    .Y(_00754_));
 sg13g2_nand3_1 _21242_ (.B(_05086_),
    .C(_05352_),
    .A(_00745_),
    .Y(_00755_));
 sg13g2_nand2_1 _21243_ (.Y(_00756_),
    .A(_00755_),
    .B(_00730_));
 sg13g2_nand2_1 _21244_ (.Y(_00757_),
    .A(_00730_),
    .B(_05334_));
 sg13g2_nand2b_1 _21245_ (.Y(_00758_),
    .B(_05333_),
    .A_N(_05349_));
 sg13g2_nand3_1 _21246_ (.B(_00757_),
    .C(_00758_),
    .A(_00756_),
    .Y(_00759_));
 sg13g2_o21ai_1 _21247_ (.B1(_00738_),
    .Y(_00760_),
    .A1(_06975_),
    .A2(_00737_));
 sg13g2_nand2_1 _21248_ (.Y(_00761_),
    .A(_00760_),
    .B(net112));
 sg13g2_nand2_1 _21249_ (.Y(_00762_),
    .A(_00759_),
    .B(_00761_));
 sg13g2_nand2_1 _21250_ (.Y(_00763_),
    .A(_00762_),
    .B(_00749_));
 sg13g2_inv_1 _21251_ (.Y(_00764_),
    .A(_00763_));
 sg13g2_nand3_1 _21252_ (.B(_00754_),
    .C(_00764_),
    .A(_00753_),
    .Y(_00765_));
 sg13g2_nand2_1 _21253_ (.Y(_00766_),
    .A(_00752_),
    .B(_00765_));
 sg13g2_nor2_1 _21254_ (.A(_00681_),
    .B(_00684_),
    .Y(_00767_));
 sg13g2_inv_1 _21255_ (.Y(_00768_),
    .A(_00767_));
 sg13g2_inv_1 _21256_ (.Y(_00769_),
    .A(_00708_));
 sg13g2_o21ai_1 _21257_ (.B1(_08037_),
    .Y(_00770_),
    .A1(_00713_),
    .A2(_00769_));
 sg13g2_nand2_1 _21258_ (.Y(_00771_),
    .A(_05340_),
    .B(net112));
 sg13g2_a21oi_1 _21259_ (.A1(_00740_),
    .A2(_00770_),
    .Y(_00773_),
    .B1(_00771_));
 sg13g2_nand2b_1 _21260_ (.Y(_00774_),
    .B(_00761_),
    .A_N(_00773_));
 sg13g2_o21ai_1 _21261_ (.B1(_05330_),
    .Y(_00775_),
    .A1(_05331_),
    .A2(_05332_));
 sg13g2_a22oi_1 _21262_ (.Y(_00776_),
    .B1(_00730_),
    .B2(_00755_),
    .A2(_00775_),
    .A1(_05350_));
 sg13g2_o21ai_1 _21263_ (.B1(_00749_),
    .Y(_00777_),
    .A1(_00774_),
    .A2(_00776_));
 sg13g2_buf_1 _21264_ (.A(_00777_),
    .X(_00778_));
 sg13g2_nand2_1 _21265_ (.Y(_00779_),
    .A(_00753_),
    .B(_00754_));
 sg13g2_a22oi_1 _21266_ (.Y(_00780_),
    .B1(_00763_),
    .B2(_00779_),
    .A2(_00778_),
    .A1(_00768_));
 sg13g2_nand2_1 _21267_ (.Y(_00781_),
    .A(_00766_),
    .B(_00780_));
 sg13g2_nand2b_1 _21268_ (.Y(_00782_),
    .B(_00767_),
    .A_N(_00778_));
 sg13g2_nand2_1 _21269_ (.Y(_00784_),
    .A(_00781_),
    .B(_00782_));
 sg13g2_nand2_1 _21270_ (.Y(_00785_),
    .A(_00784_),
    .B(_00750_));
 sg13g2_nand2_1 _21271_ (.Y(_00786_),
    .A(_00686_),
    .B(_00688_));
 sg13g2_inv_1 _21272_ (.Y(_00787_),
    .A(_00786_));
 sg13g2_nand3_1 _21273_ (.B(_00782_),
    .C(_00787_),
    .A(_00781_),
    .Y(_00788_));
 sg13g2_buf_1 _21274_ (.A(_00788_),
    .X(_00789_));
 sg13g2_inv_1 _21275_ (.Y(_00790_),
    .A(_00699_));
 sg13g2_a21oi_1 _21276_ (.A1(_00790_),
    .A2(net40),
    .Y(_00791_),
    .B1(_05532_));
 sg13g2_a21oi_1 _21277_ (.A1(_00720_),
    .A2(net40),
    .Y(_00792_),
    .B1(_06979_));
 sg13g2_nor2_1 _21278_ (.A(_07108_),
    .B(_07141_),
    .Y(_00793_));
 sg13g2_nor2_1 _21279_ (.A(_09054_),
    .B(_09049_),
    .Y(_00795_));
 sg13g2_or2_1 _21280_ (.X(_00796_),
    .B(_00795_),
    .A(_00793_));
 sg13g2_a221oi_1 _21281_ (.B2(_00792_),
    .C1(_00796_),
    .B1(_00791_),
    .A1(_07709_),
    .Y(_00797_),
    .A2(_11748_));
 sg13g2_inv_1 _21282_ (.Y(_00798_),
    .A(_00791_));
 sg13g2_inv_1 _21283_ (.Y(_00799_),
    .A(_07709_));
 sg13g2_nand2_1 _21284_ (.Y(_00800_),
    .A(_00799_),
    .B(_11748_));
 sg13g2_o21ai_1 _21285_ (.B1(_00800_),
    .Y(_00801_),
    .A1(_07108_),
    .A2(_07140_));
 sg13g2_a221oi_1 _21286_ (.B2(_00792_),
    .C1(_00801_),
    .B1(_00798_),
    .A1(_09049_),
    .Y(_00802_),
    .A2(_09053_));
 sg13g2_a21o_1 _21287_ (.A2(_00802_),
    .A1(_00797_),
    .B1(_06221_),
    .X(_00803_));
 sg13g2_a22oi_1 _21288_ (.Y(_00804_),
    .B1(_09682_),
    .B2(_09677_),
    .A2(_06218_),
    .A1(_06168_));
 sg13g2_o21ai_1 _21289_ (.B1(_00804_),
    .Y(_00806_),
    .A1(_08658_),
    .A2(_08691_));
 sg13g2_nor2_1 _21290_ (.A(_10017_),
    .B(_10024_),
    .Y(_00807_));
 sg13g2_nor2_1 _21291_ (.A(_00806_),
    .B(_00807_),
    .Y(_00808_));
 sg13g2_inv_1 _21292_ (.Y(_00809_),
    .A(_00808_));
 sg13g2_inv_1 _21293_ (.Y(_00810_),
    .A(_08658_));
 sg13g2_a22oi_1 _21294_ (.Y(_00811_),
    .B1(_09682_),
    .B2(_09678_),
    .A2(_06218_),
    .A1(_06169_));
 sg13g2_inv_1 _21295_ (.Y(_00812_),
    .A(_00811_));
 sg13g2_a21oi_1 _21296_ (.A1(_08691_),
    .A2(_00810_),
    .Y(_00813_),
    .B1(_00812_));
 sg13g2_o21ai_1 _21297_ (.B1(_00813_),
    .Y(_00814_),
    .A1(_10023_),
    .A2(_10017_));
 sg13g2_o21ai_1 _21298_ (.B1(_06177_),
    .Y(_00815_),
    .A1(_00809_),
    .A2(_00814_));
 sg13g2_a21o_1 _21299_ (.A2(_00815_),
    .A1(_00803_),
    .B1(_06225_),
    .X(_00817_));
 sg13g2_nand2b_1 _21300_ (.Y(_00818_),
    .B(_06223_),
    .A_N(_00815_));
 sg13g2_nand3_1 _21301_ (.B(_06175_),
    .C(_00818_),
    .A(_00817_),
    .Y(_00819_));
 sg13g2_nor3_1 _21302_ (.A(_08940_),
    .B(_09118_),
    .C(_07809_),
    .Y(_00820_));
 sg13g2_nor4_1 _21303_ (.A(_07812_),
    .B(_07993_),
    .C(_07801_),
    .D(_09115_),
    .Y(_00821_));
 sg13g2_nand3_1 _21304_ (.B(_08463_),
    .C(_00821_),
    .A(_00820_),
    .Y(_00822_));
 sg13g2_inv_1 _21305_ (.Y(_00823_),
    .A(_00822_));
 sg13g2_nor2_1 _21306_ (.A(_09103_),
    .B(_07715_),
    .Y(_00824_));
 sg13g2_nand2b_1 _21307_ (.Y(_00825_),
    .B(_08842_),
    .A_N(_09001_));
 sg13g2_nor3_1 _21308_ (.A(_07720_),
    .B(_00825_),
    .C(_09106_),
    .Y(_00826_));
 sg13g2_nand2_1 _21309_ (.Y(_00828_),
    .A(_00722_),
    .B(_00826_));
 sg13g2_nor3_1 _21310_ (.A(_06175_),
    .B(net14),
    .C(_00828_),
    .Y(_00829_));
 sg13g2_nand3_1 _21311_ (.B(_00824_),
    .C(_00829_),
    .A(_00823_),
    .Y(_00830_));
 sg13g2_nor2_1 _21312_ (.A(net83),
    .B(_06178_),
    .Y(_00831_));
 sg13g2_nand3_1 _21313_ (.B(_00830_),
    .C(_00831_),
    .A(_00819_),
    .Y(_00832_));
 sg13g2_nor2_1 _21314_ (.A(_06904_),
    .B(_05015_),
    .Y(_00833_));
 sg13g2_nand2_1 _21315_ (.Y(_00834_),
    .A(_11429_),
    .B(_00833_));
 sg13g2_nor4_1 _21316_ (.A(_05017_),
    .B(_07919_),
    .C(_10778_),
    .D(_00834_),
    .Y(_00835_));
 sg13g2_nand4_1 _21317_ (.B(_00797_),
    .C(_00808_),
    .A(_00823_),
    .Y(_00836_),
    .D(_00835_));
 sg13g2_nor4_1 _21318_ (.A(_07029_),
    .B(_04585_),
    .C(_04528_),
    .D(_06296_),
    .Y(_00837_));
 sg13g2_nor2_1 _21319_ (.A(_08676_),
    .B(_10277_),
    .Y(_00839_));
 sg13g2_nand4_1 _21320_ (.B(_07939_),
    .C(_10213_),
    .A(_00837_),
    .Y(_00840_),
    .D(_00839_));
 sg13g2_nor4_1 _21321_ (.A(net14),
    .B(_00840_),
    .C(_00828_),
    .D(_00814_),
    .Y(_00841_));
 sg13g2_and3_1 _21322_ (.X(_00842_),
    .A(_00802_),
    .B(_00824_),
    .C(_00841_));
 sg13g2_nand2b_1 _21323_ (.Y(_00843_),
    .B(_00842_),
    .A_N(_00836_));
 sg13g2_o21ai_1 _21324_ (.B1(_06220_),
    .Y(_00844_),
    .A1(_06173_),
    .A2(_06177_));
 sg13g2_nand3_1 _21325_ (.B(net86),
    .C(_00844_),
    .A(_00843_),
    .Y(_00845_));
 sg13g2_nor2_1 _21326_ (.A(_06177_),
    .B(_00842_),
    .Y(_00846_));
 sg13g2_nand3_1 _21327_ (.B(net145),
    .C(_00846_),
    .A(_00836_),
    .Y(_00847_));
 sg13g2_or2_1 _21328_ (.X(_00848_),
    .B(_00847_),
    .A(_06173_));
 sg13g2_nand3_1 _21329_ (.B(_00845_),
    .C(_00848_),
    .A(_00832_),
    .Y(_00850_));
 sg13g2_buf_1 _21330_ (.A(\b.gen_square[29].sq.mask ),
    .X(_00851_));
 sg13g2_nand2_1 _21331_ (.Y(_00852_),
    .A(_00850_),
    .B(_00851_));
 sg13g2_nand3_1 _21332_ (.B(_00789_),
    .C(_00852_),
    .A(_00785_),
    .Y(_00853_));
 sg13g2_nor2_1 _21333_ (.A(net93),
    .B(_07700_),
    .Y(_00854_));
 sg13g2_inv_1 _21334_ (.Y(_00855_),
    .A(_00835_));
 sg13g2_o21ai_1 _21335_ (.B1(_08411_),
    .Y(_00856_),
    .A1(_00855_),
    .A2(_00840_));
 sg13g2_nand2_1 _21336_ (.Y(_00857_),
    .A(_00818_),
    .B(_00856_));
 sg13g2_xnor2_1 _21337_ (.Y(_00858_),
    .A(_06172_),
    .B(_06224_));
 sg13g2_nand3_1 _21338_ (.B(_05087_),
    .C(_06221_),
    .A(_00843_),
    .Y(_00859_));
 sg13g2_nand2_1 _21339_ (.Y(_00861_),
    .A(_00859_),
    .B(_00847_));
 sg13g2_a22oi_1 _21340_ (.Y(_00862_),
    .B1(_00858_),
    .B2(_00861_),
    .A2(_00857_),
    .A1(_00854_));
 sg13g2_o21ai_1 _21341_ (.B1(_00817_),
    .Y(_00863_),
    .A1(_07110_),
    .A2(_00803_));
 sg13g2_nand2_1 _21342_ (.Y(_00864_),
    .A(_00863_),
    .B(net85));
 sg13g2_nand2_1 _21343_ (.Y(_00865_),
    .A(_00862_),
    .B(_00864_));
 sg13g2_nand2_1 _21344_ (.Y(_00866_),
    .A(_00865_),
    .B(_00851_));
 sg13g2_inv_1 _21345_ (.Y(_00867_),
    .A(_00866_));
 sg13g2_nand2_1 _21346_ (.Y(_00868_),
    .A(_00767_),
    .B(_00778_));
 sg13g2_xnor2_1 _21347_ (.Y(_00869_),
    .A(_00867_),
    .B(_00868_));
 sg13g2_nand2_1 _21348_ (.Y(_00870_),
    .A(_00853_),
    .B(_00869_));
 sg13g2_nand2_1 _21349_ (.Y(_00872_),
    .A(_00784_),
    .B(_00764_));
 sg13g2_nand3_1 _21350_ (.B(_00779_),
    .C(_00782_),
    .A(_00781_),
    .Y(_00873_));
 sg13g2_nand2_1 _21351_ (.Y(_00874_),
    .A(_00872_),
    .B(_00873_));
 sg13g2_nand2_1 _21352_ (.Y(_00875_),
    .A(_00847_),
    .B(_06183_));
 sg13g2_nand2b_1 _21353_ (.Y(_00876_),
    .B(_06182_),
    .A_N(_06224_));
 sg13g2_nand3_1 _21354_ (.B(_00875_),
    .C(_00876_),
    .A(_00861_),
    .Y(_00877_));
 sg13g2_nand2_1 _21355_ (.Y(_00878_),
    .A(_00877_),
    .B(_00864_));
 sg13g2_nand2_1 _21356_ (.Y(_00879_),
    .A(_00878_),
    .B(_00851_));
 sg13g2_nand2_1 _21357_ (.Y(_00880_),
    .A(_00874_),
    .B(_00879_));
 sg13g2_inv_1 _21358_ (.Y(_00881_),
    .A(_00879_));
 sg13g2_nand3_1 _21359_ (.B(_00873_),
    .C(_00881_),
    .A(_00872_),
    .Y(_00883_));
 sg13g2_nand2_1 _21360_ (.Y(_00884_),
    .A(_00880_),
    .B(_00883_));
 sg13g2_nor2_1 _21361_ (.A(_00870_),
    .B(_00884_),
    .Y(_00885_));
 sg13g2_a21oi_1 _21362_ (.A1(_00785_),
    .A2(_00789_),
    .Y(_00886_),
    .B1(_00852_));
 sg13g2_nand2_1 _21363_ (.Y(_00887_),
    .A(_00885_),
    .B(_00886_));
 sg13g2_inv_1 _21364_ (.Y(_00888_),
    .A(_00868_));
 sg13g2_nor2b_1 _21365_ (.A(_00883_),
    .B_N(_00869_),
    .Y(_00889_));
 sg13g2_a21oi_2 _21366_ (.B1(_00889_),
    .Y(_00890_),
    .A2(_00888_),
    .A1(_00867_));
 sg13g2_nand2_1 _21367_ (.Y(_00891_),
    .A(_00785_),
    .B(_00789_));
 sg13g2_nand3_1 _21368_ (.B(_00890_),
    .C(_00891_),
    .A(_00887_),
    .Y(_00892_));
 sg13g2_nand2b_1 _21369_ (.Y(_00894_),
    .B(_00852_),
    .A_N(_00890_));
 sg13g2_nand2_1 _21370_ (.Y(_00895_),
    .A(_00892_),
    .B(_00894_));
 sg13g2_nand2_1 _21371_ (.Y(_00896_),
    .A(_00887_),
    .B(_00890_));
 sg13g2_nand2_1 _21372_ (.Y(_00897_),
    .A(_00896_),
    .B(_00879_));
 sg13g2_inv_1 _21373_ (.Y(_00898_),
    .A(_00874_));
 sg13g2_nand3_1 _21374_ (.B(_00890_),
    .C(_00898_),
    .A(_00887_),
    .Y(_00899_));
 sg13g2_nand2_1 _21375_ (.Y(_00900_),
    .A(_00897_),
    .B(_00899_));
 sg13g2_inv_1 _21376_ (.Y(_00901_),
    .A(_11620_));
 sg13g2_a21oi_1 _21377_ (.A1(_06683_),
    .A2(_08944_),
    .Y(_00902_),
    .B1(_07492_));
 sg13g2_nor2_1 _21378_ (.A(_06625_),
    .B(_07250_),
    .Y(_00903_));
 sg13g2_inv_1 _21379_ (.Y(_00905_),
    .A(_00903_));
 sg13g2_nor3_1 _21380_ (.A(_07752_),
    .B(_10614_),
    .C(_00905_),
    .Y(_00906_));
 sg13g2_nor2b_1 _21381_ (.A(_00902_),
    .B_N(_00906_),
    .Y(_00907_));
 sg13g2_nand2_1 _21382_ (.Y(_00908_),
    .A(_08807_),
    .B(_08800_));
 sg13g2_nor2_1 _21383_ (.A(_07225_),
    .B(_08733_),
    .Y(_00909_));
 sg13g2_nor4_1 _21384_ (.A(_10120_),
    .B(_00909_),
    .C(_08737_),
    .D(_06641_),
    .Y(_00910_));
 sg13g2_nand4_1 _21385_ (.B(_00908_),
    .C(_07721_),
    .A(_00907_),
    .Y(_00911_),
    .D(_00910_));
 sg13g2_a21oi_1 _21386_ (.A1(_11624_),
    .A2(_00901_),
    .Y(_00912_),
    .B1(_00911_));
 sg13g2_inv_1 _21387_ (.Y(_00913_),
    .A(_04221_));
 sg13g2_a22oi_1 _21388_ (.Y(_00914_),
    .B1(_04296_),
    .B2(_00913_),
    .A2(_07532_),
    .A1(_04098_));
 sg13g2_o21ai_1 _21389_ (.B1(_00914_),
    .Y(_00916_),
    .A1(_08925_),
    .A2(_08921_));
 sg13g2_inv_1 _21390_ (.Y(_00917_),
    .A(_00916_));
 sg13g2_nor3_1 _21391_ (.A(_09001_),
    .B(_07962_),
    .C(_09103_),
    .Y(_00918_));
 sg13g2_nand3_1 _21392_ (.B(_00917_),
    .C(_00918_),
    .A(_00912_),
    .Y(_00919_));
 sg13g2_a21oi_1 _21393_ (.A1(_00798_),
    .A2(net27),
    .Y(_00920_),
    .B1(_06189_));
 sg13g2_inv_1 _21394_ (.Y(_00921_),
    .A(_00792_));
 sg13g2_a21oi_1 _21395_ (.A1(_00921_),
    .A2(net27),
    .Y(_00922_),
    .B1(_07114_));
 sg13g2_inv_1 _21396_ (.Y(_00923_),
    .A(_00922_));
 sg13g2_nor2_1 _21397_ (.A(_00920_),
    .B(_00923_),
    .Y(_00924_));
 sg13g2_nor4_1 _21398_ (.A(_08734_),
    .B(_07704_),
    .C(_00919_),
    .D(_00924_),
    .Y(_00925_));
 sg13g2_inv_1 _21399_ (.Y(_00927_),
    .A(_00925_));
 sg13g2_nor2b_1 _21400_ (.A(_00923_),
    .B_N(_00920_),
    .Y(_00928_));
 sg13g2_inv_1 _21401_ (.Y(_00929_),
    .A(_00928_));
 sg13g2_nand2_1 _21402_ (.Y(_00930_),
    .A(_04221_),
    .B(_04296_));
 sg13g2_nor4_1 _21403_ (.A(_07812_),
    .B(_08699_),
    .C(_08940_),
    .D(_07815_),
    .Y(_00931_));
 sg13g2_nor2_1 _21404_ (.A(_04985_),
    .B(_07225_),
    .Y(_00932_));
 sg13g2_inv_1 _21405_ (.Y(_00933_),
    .A(_00704_));
 sg13g2_nand2_1 _21406_ (.Y(_00934_),
    .A(_08806_),
    .B(_08800_));
 sg13g2_nor4_1 _21407_ (.A(_08967_),
    .B(_08703_),
    .C(_08945_),
    .D(_10635_),
    .Y(_00935_));
 sg13g2_nor2_1 _21408_ (.A(_06650_),
    .B(_07170_),
    .Y(_00936_));
 sg13g2_inv_1 _21409_ (.Y(_00938_),
    .A(_00936_));
 sg13g2_nor3_1 _21410_ (.A(_06646_),
    .B(_10170_),
    .C(_00938_),
    .Y(_00939_));
 sg13g2_nand3_1 _21411_ (.B(_00935_),
    .C(_00939_),
    .A(_00934_),
    .Y(_00940_));
 sg13g2_a22oi_1 _21412_ (.Y(_00941_),
    .B1(_08925_),
    .B2(_08920_),
    .A2(_07532_),
    .A1(_08705_));
 sg13g2_o21ai_1 _21413_ (.B1(_00941_),
    .Y(_00942_),
    .A1(_11624_),
    .A2(_11620_));
 sg13g2_nor4_1 _21414_ (.A(_00932_),
    .B(_00933_),
    .C(_00940_),
    .D(_00942_),
    .Y(_00943_));
 sg13g2_nand4_1 _21415_ (.B(_00930_),
    .C(_00931_),
    .A(_00929_),
    .Y(_00944_),
    .D(_00943_));
 sg13g2_nor2_1 _21416_ (.A(_00927_),
    .B(_00944_),
    .Y(_00945_));
 sg13g2_inv_1 _21417_ (.Y(_00946_),
    .A(_00945_));
 sg13g2_nand3_1 _21418_ (.B(net76),
    .C(_04299_),
    .A(_00946_),
    .Y(_00947_));
 sg13g2_nand4_1 _21419_ (.B(_00927_),
    .C(net130),
    .A(_00944_),
    .Y(_00948_),
    .D(_04299_));
 sg13g2_buf_1 _21420_ (.A(_00948_),
    .X(_00949_));
 sg13g2_o21ai_1 _21421_ (.B1(_00949_),
    .Y(_00950_),
    .A1(_04139_),
    .A2(_00947_));
 sg13g2_o21ai_1 _21422_ (.B1(_00950_),
    .Y(_00951_),
    .A1(_04304_),
    .A2(_04302_));
 sg13g2_nand3b_1 _21423_ (.B(_00941_),
    .C(_00930_),
    .Y(_00952_),
    .A_N(_00916_));
 sg13g2_o21ai_1 _21424_ (.B1(_04148_),
    .Y(_00953_),
    .A1(_00952_),
    .A2(_00922_));
 sg13g2_nand3_1 _21425_ (.B(_06683_),
    .C(_07225_),
    .A(_08801_),
    .Y(_00954_));
 sg13g2_o21ai_1 _21426_ (.B1(_04148_),
    .Y(_00955_),
    .A1(_00954_),
    .A2(_00901_));
 sg13g2_a21o_1 _21427_ (.A2(_00955_),
    .A1(_00953_),
    .B1(_04305_),
    .X(_00956_));
 sg13g2_o21ai_1 _21428_ (.B1(_00956_),
    .Y(_00957_),
    .A1(_04303_),
    .A2(_00953_));
 sg13g2_nand2_1 _21429_ (.Y(_00959_),
    .A(_00957_),
    .B(net75));
 sg13g2_nand2_1 _21430_ (.Y(_00960_),
    .A(_00951_),
    .B(_00959_));
 sg13g2_buf_1 _21431_ (.A(\b.gen_square[30].sq.mask ),
    .X(_00961_));
 sg13g2_nand2_1 _21432_ (.Y(_00962_),
    .A(_00960_),
    .B(_00961_));
 sg13g2_inv_1 _21433_ (.Y(_00963_),
    .A(_00962_));
 sg13g2_nor2_1 _21434_ (.A(_02100_),
    .B(_07722_),
    .Y(_00964_));
 sg13g2_nand2b_1 _21435_ (.Y(_00965_),
    .B(_06684_),
    .A_N(_00955_));
 sg13g2_nand4_1 _21436_ (.B(_00906_),
    .C(_10634_),
    .A(_00939_),
    .Y(_00966_),
    .D(_11510_));
 sg13g2_nand2_1 _21437_ (.Y(_00967_),
    .A(_00966_),
    .B(_07894_));
 sg13g2_nand2_1 _21438_ (.Y(_00968_),
    .A(_00965_),
    .B(_00967_));
 sg13g2_xnor2_1 _21439_ (.Y(_00970_),
    .A(_04135_),
    .B(_04304_));
 sg13g2_nand2_1 _21440_ (.Y(_00971_),
    .A(_00947_),
    .B(_00949_));
 sg13g2_a22oi_1 _21441_ (.Y(_00972_),
    .B1(_00970_),
    .B2(_00971_),
    .A2(_00968_),
    .A1(_00964_));
 sg13g2_nand2_1 _21442_ (.Y(_00973_),
    .A(_00972_),
    .B(_00959_));
 sg13g2_nand2_1 _21443_ (.Y(_00974_),
    .A(_00973_),
    .B(_00961_));
 sg13g2_nor2_1 _21444_ (.A(_00867_),
    .B(_00868_),
    .Y(_00975_));
 sg13g2_inv_1 _21445_ (.Y(_00976_),
    .A(_00975_));
 sg13g2_nor2_1 _21446_ (.A(_00974_),
    .B(_00976_),
    .Y(_00977_));
 sg13g2_a21oi_1 _21447_ (.A1(_00900_),
    .A2(_00963_),
    .Y(_00978_),
    .B1(_00977_));
 sg13g2_nand3_1 _21448_ (.B(_04146_),
    .C(_00965_),
    .A(_00956_),
    .Y(_00979_));
 sg13g2_inv_1 _21449_ (.Y(_00981_),
    .A(_04149_));
 sg13g2_nand3_1 _21450_ (.B(_07722_),
    .C(_08944_),
    .A(_08702_),
    .Y(_00982_));
 sg13g2_inv_1 _21451_ (.Y(_00983_),
    .A(_00918_));
 sg13g2_nor3_1 _21452_ (.A(_07720_),
    .B(_00982_),
    .C(_00983_),
    .Y(_00984_));
 sg13g2_nor2_1 _21453_ (.A(_08734_),
    .B(_07704_),
    .Y(_00985_));
 sg13g2_nand4_1 _21454_ (.B(_00931_),
    .C(_00704_),
    .A(_00984_),
    .Y(_00986_),
    .D(_00985_));
 sg13g2_nand4_1 _21455_ (.B(_05114_),
    .C(_00981_),
    .A(_00979_),
    .Y(_00987_),
    .D(_00986_));
 sg13g2_or2_1 _21456_ (.X(_00988_),
    .B(_00949_),
    .A(_04137_));
 sg13g2_o21ai_1 _21457_ (.B1(_04140_),
    .Y(_00989_),
    .A1(_04137_),
    .A2(_04148_));
 sg13g2_nand3_1 _21458_ (.B(_05090_),
    .C(_00989_),
    .A(_00946_),
    .Y(_00990_));
 sg13g2_nand3_1 _21459_ (.B(_00988_),
    .C(_00990_),
    .A(_00987_),
    .Y(_00992_));
 sg13g2_nand2_1 _21460_ (.Y(_00993_),
    .A(_00992_),
    .B(_00961_));
 sg13g2_a21oi_1 _21461_ (.A1(_00892_),
    .A2(_00894_),
    .Y(_00994_),
    .B1(_00993_));
 sg13g2_nand3_1 _21462_ (.B(_00899_),
    .C(_00962_),
    .A(_00897_),
    .Y(_00995_));
 sg13g2_nand2_1 _21463_ (.Y(_00996_),
    .A(_00994_),
    .B(_00995_));
 sg13g2_nand2_1 _21464_ (.Y(_00997_),
    .A(_00978_),
    .B(_00996_));
 sg13g2_nand2_1 _21465_ (.Y(_00998_),
    .A(_00976_),
    .B(_00974_));
 sg13g2_nand2_1 _21466_ (.Y(_00999_),
    .A(_00997_),
    .B(_00998_));
 sg13g2_nand2b_1 _21467_ (.Y(_01000_),
    .B(_00999_),
    .A_N(_00895_));
 sg13g2_nand3b_1 _21468_ (.B(_00997_),
    .C(_00998_),
    .Y(_01001_),
    .A_N(_00993_));
 sg13g2_nand2_1 _21469_ (.Y(_01003_),
    .A(_01000_),
    .B(_01001_));
 sg13g2_a21oi_1 _21470_ (.A1(_08649_),
    .A2(net34),
    .Y(_01004_),
    .B1(_06868_));
 sg13g2_inv_1 _21471_ (.Y(_01005_),
    .A(_01004_));
 sg13g2_inv_1 _21472_ (.Y(_01006_),
    .A(_11001_));
 sg13g2_a21oi_1 _21473_ (.A1(_01006_),
    .A2(net47),
    .Y(_01007_),
    .B1(_06217_));
 sg13g2_inv_1 _21474_ (.Y(_01008_),
    .A(_01007_));
 sg13g2_a21oi_1 _21475_ (.A1(_01005_),
    .A2(_01008_),
    .Y(_01009_),
    .B1(_06855_));
 sg13g2_inv_1 _21476_ (.Y(_01010_),
    .A(_01009_));
 sg13g2_nor2_1 _21477_ (.A(_06859_),
    .B(_01010_),
    .Y(_01011_));
 sg13g2_nor2_1 _21478_ (.A(_10011_),
    .B(_10006_),
    .Y(_01012_));
 sg13g2_inv_1 _21479_ (.Y(_01014_),
    .A(_07493_));
 sg13g2_inv_1 _21480_ (.Y(_01015_),
    .A(_07525_));
 sg13g2_o21ai_1 _21481_ (.B1(_04225_),
    .Y(_01016_),
    .A1(_04155_),
    .A2(_00920_));
 sg13g2_a21oi_1 _21482_ (.A1(_00923_),
    .A2(net33),
    .Y(_01017_),
    .B1(_04309_));
 sg13g2_nor2b_1 _21483_ (.A(_01016_),
    .B_N(_01017_),
    .Y(_01018_));
 sg13g2_a221oi_1 _21484_ (.B2(_10005_),
    .C1(_01018_),
    .B1(_10011_),
    .A1(_01014_),
    .Y(_01019_),
    .A2(_01015_));
 sg13g2_a22oi_1 _21485_ (.Y(_01020_),
    .B1(_01017_),
    .B2(_01016_),
    .A2(_01015_),
    .A1(_07493_));
 sg13g2_nand2_1 _21486_ (.Y(_01021_),
    .A(_01019_),
    .B(_01020_));
 sg13g2_o21ai_1 _21487_ (.B1(_04081_),
    .Y(_01022_),
    .A1(_01012_),
    .A2(_01021_));
 sg13g2_a21o_1 _21488_ (.A2(_01010_),
    .A1(_01022_),
    .B1(_06857_),
    .X(_01023_));
 sg13g2_nand3b_1 _21489_ (.B(_01023_),
    .C(_04075_),
    .Y(_01025_),
    .A_N(_01011_));
 sg13g2_nor2_1 _21490_ (.A(_08945_),
    .B(_08940_),
    .Y(_01026_));
 sg13g2_o21ai_1 _21491_ (.B1(_01026_),
    .Y(_01027_),
    .A1(_08698_),
    .A2(_10012_));
 sg13g2_nor3_1 _21492_ (.A(_07812_),
    .B(_07801_),
    .C(_01027_),
    .Y(_01028_));
 sg13g2_nor2_1 _21493_ (.A(_08698_),
    .B(_10011_),
    .Y(_01029_));
 sg13g2_nor3_1 _21494_ (.A(_08998_),
    .B(_00825_),
    .C(_01029_),
    .Y(_01030_));
 sg13g2_nand4_1 _21495_ (.B(_08700_),
    .C(_07721_),
    .A(_01028_),
    .Y(_01031_),
    .D(_01030_));
 sg13g2_nor2_1 _21496_ (.A(_02100_),
    .B(_04082_),
    .Y(_01032_));
 sg13g2_nand3_1 _21497_ (.B(_01031_),
    .C(_01032_),
    .A(_01025_),
    .Y(_01033_));
 sg13g2_a21oi_1 _21498_ (.A1(_08723_),
    .A2(_04117_),
    .Y(_01034_),
    .B1(_04120_));
 sg13g2_a21oi_1 _21499_ (.A1(_11004_),
    .A2(net47),
    .Y(_01036_),
    .B1(_04220_));
 sg13g2_inv_1 _21500_ (.Y(_01037_),
    .A(_01036_));
 sg13g2_nor2_1 _21501_ (.A(_06906_),
    .B(_10243_),
    .Y(_01038_));
 sg13g2_o21ai_1 _21502_ (.B1(_01038_),
    .Y(_01039_),
    .A1(_01008_),
    .A2(_01037_));
 sg13g2_a21oi_1 _21503_ (.A1(_01034_),
    .A2(_01004_),
    .Y(_01040_),
    .B1(_01039_));
 sg13g2_nand3_1 _21504_ (.B(_01040_),
    .C(_01028_),
    .A(_01019_),
    .Y(_01041_));
 sg13g2_nor3_1 _21505_ (.A(_07029_),
    .B(_07936_),
    .C(_11414_),
    .Y(_01042_));
 sg13g2_inv_1 _21506_ (.Y(_01043_),
    .A(_01042_));
 sg13g2_nand2_1 _21507_ (.Y(_01044_),
    .A(_01037_),
    .B(_01007_));
 sg13g2_o21ai_1 _21508_ (.B1(_01044_),
    .Y(_01045_),
    .A1(_01005_),
    .A2(_01034_));
 sg13g2_nor4_1 _21509_ (.A(_07720_),
    .B(_01012_),
    .C(_01043_),
    .D(_01045_),
    .Y(_01047_));
 sg13g2_nand3_1 _21510_ (.B(_01030_),
    .C(_01047_),
    .A(_01020_),
    .Y(_01048_));
 sg13g2_and3_1 _21511_ (.X(_01049_),
    .A(_01041_),
    .B(_06855_),
    .C(_01048_));
 sg13g2_nand2_1 _21512_ (.Y(_01050_),
    .A(_01049_),
    .B(_05078_));
 sg13g2_inv_1 _21513_ (.Y(_01051_),
    .A(_01050_));
 sg13g2_nor2_1 _21514_ (.A(_04095_),
    .B(_06855_),
    .Y(_01052_));
 sg13g2_nor2_1 _21515_ (.A(_07738_),
    .B(_04095_),
    .Y(_01053_));
 sg13g2_nor2_1 _21516_ (.A(_01048_),
    .B(_01041_),
    .Y(_01054_));
 sg13g2_nor4_1 _21517_ (.A(_07412_),
    .B(_01052_),
    .C(_01053_),
    .D(_01054_),
    .Y(_01055_));
 sg13g2_a21oi_1 _21518_ (.A1(_01051_),
    .A2(_07738_),
    .Y(_01056_),
    .B1(_01055_));
 sg13g2_buf_1 _21519_ (.A(\b.gen_square[31].sq.mask ),
    .X(_01058_));
 sg13g2_inv_1 _21520_ (.Y(_01059_),
    .A(_01058_));
 sg13g2_a21o_1 _21521_ (.A2(_01056_),
    .A1(_01033_),
    .B1(_01059_),
    .X(_01060_));
 sg13g2_nor2_1 _21522_ (.A(_01060_),
    .B(_01003_),
    .Y(_01061_));
 sg13g2_nand2_1 _21523_ (.Y(_01062_),
    .A(_00999_),
    .B(_00900_));
 sg13g2_nand3_1 _21524_ (.B(_00998_),
    .C(_00962_),
    .A(_00997_),
    .Y(_01063_));
 sg13g2_inv_1 _21525_ (.Y(_01064_),
    .A(_04095_));
 sg13g2_inv_1 _21526_ (.Y(_01065_),
    .A(_06856_));
 sg13g2_inv_1 _21527_ (.Y(_01066_),
    .A(_01054_));
 sg13g2_nand3_1 _21528_ (.B(_05090_),
    .C(_06855_),
    .A(_01066_),
    .Y(_01067_));
 sg13g2_a22oi_1 _21529_ (.Y(_01068_),
    .B1(_01067_),
    .B2(_01050_),
    .A2(_04094_),
    .A1(_01065_));
 sg13g2_o21ai_1 _21530_ (.B1(_01068_),
    .Y(_01069_),
    .A1(_01064_),
    .A2(_01051_));
 sg13g2_o21ai_1 _21531_ (.B1(_01023_),
    .Y(_01070_),
    .A1(_07528_),
    .A2(_01022_));
 sg13g2_nand2_1 _21532_ (.Y(_01071_),
    .A(_01070_),
    .B(_05114_));
 sg13g2_nand2_1 _21533_ (.Y(_01072_),
    .A(_01069_),
    .B(_01071_));
 sg13g2_nand2_1 _21534_ (.Y(_01073_),
    .A(_01072_),
    .B(_01058_));
 sg13g2_nand3_1 _21535_ (.B(_01063_),
    .C(_01073_),
    .A(_01062_),
    .Y(_01074_));
 sg13g2_nand2_1 _21536_ (.Y(_01075_),
    .A(_01061_),
    .B(_01074_));
 sg13g2_nand2_1 _21537_ (.Y(_01076_),
    .A(_01062_),
    .B(_01063_));
 sg13g2_inv_1 _21538_ (.Y(_01077_),
    .A(_01073_));
 sg13g2_nand2_1 _21539_ (.Y(_01079_),
    .A(_01076_),
    .B(_01077_));
 sg13g2_nand2_1 _21540_ (.Y(_01080_),
    .A(_01065_),
    .B(_04093_));
 sg13g2_a22oi_1 _21541_ (.Y(_01081_),
    .B1(_01067_),
    .B2(_01050_),
    .A2(_01080_),
    .A1(_06857_));
 sg13g2_a21oi_1 _21542_ (.A1(_01042_),
    .A2(_01038_),
    .Y(_01082_),
    .B1(_07740_));
 sg13g2_nor3_1 _21543_ (.A(_01011_),
    .B(_01082_),
    .C(_01070_),
    .Y(_01083_));
 sg13g2_nor2_1 _21544_ (.A(_02111_),
    .B(_01083_),
    .Y(_01084_));
 sg13g2_o21ai_1 _21545_ (.B1(_01058_),
    .Y(_01085_),
    .A1(_01081_),
    .A2(_01084_));
 sg13g2_buf_1 _21546_ (.A(_01085_),
    .X(_01086_));
 sg13g2_nand2_1 _21547_ (.Y(_01087_),
    .A(_00975_),
    .B(_00974_));
 sg13g2_xor2_1 _21548_ (.B(_01087_),
    .A(_01086_),
    .X(_01088_));
 sg13g2_nand3_1 _21549_ (.B(_01079_),
    .C(_01088_),
    .A(_01075_),
    .Y(_01090_));
 sg13g2_buf_1 _21550_ (.A(_01090_),
    .X(_01091_));
 sg13g2_nand2_1 _21551_ (.Y(_01092_),
    .A(_01087_),
    .B(_01086_));
 sg13g2_nand2_1 _21552_ (.Y(_01093_),
    .A(_01091_),
    .B(_01092_));
 sg13g2_nand2b_1 _21553_ (.Y(_01094_),
    .B(_01093_),
    .A_N(_01003_));
 sg13g2_nand3_1 _21554_ (.B(_01092_),
    .C(_01060_),
    .A(_01091_),
    .Y(_01095_));
 sg13g2_nand2_1 _21555_ (.Y(_01096_),
    .A(_01094_),
    .B(_01095_));
 sg13g2_nand3_1 _21556_ (.B(_11731_),
    .C(_01096_),
    .A(_11728_),
    .Y(_01097_));
 sg13g2_nor2b_2 _21557_ (.A(_01087_),
    .B_N(_01086_),
    .Y(_01098_));
 sg13g2_inv_1 _21558_ (.Y(_01099_),
    .A(_11705_));
 sg13g2_nor2_1 _21559_ (.A(_11704_),
    .B(_01099_),
    .Y(_01101_));
 sg13g2_xnor2_1 _21560_ (.Y(_01102_),
    .A(_01098_),
    .B(_01101_));
 sg13g2_nand2_1 _21561_ (.Y(_01103_),
    .A(_01097_),
    .B(_01102_));
 sg13g2_nand2_1 _21562_ (.Y(_01104_),
    .A(_11727_),
    .B(_11712_));
 sg13g2_nand2_1 _21563_ (.Y(_01105_),
    .A(_11708_),
    .B(_11709_));
 sg13g2_nand3_1 _21564_ (.B(_01105_),
    .C(_11725_),
    .A(_11723_),
    .Y(_01106_));
 sg13g2_nand2_1 _21565_ (.Y(_01107_),
    .A(_01104_),
    .B(_01106_));
 sg13g2_nand2b_1 _21566_ (.Y(_01108_),
    .B(_01093_),
    .A_N(_01076_));
 sg13g2_nand3_1 _21567_ (.B(_01092_),
    .C(_01077_),
    .A(_01091_),
    .Y(_01109_));
 sg13g2_nand2_1 _21568_ (.Y(_01110_),
    .A(_01108_),
    .B(_01109_));
 sg13g2_inv_1 _21569_ (.Y(_01112_),
    .A(_01110_));
 sg13g2_nand2_1 _21570_ (.Y(_01113_),
    .A(_01107_),
    .B(_01112_));
 sg13g2_nand3_1 _21571_ (.B(_01106_),
    .C(_01110_),
    .A(_01104_),
    .Y(_01114_));
 sg13g2_nand2_1 _21572_ (.Y(_01115_),
    .A(_01113_),
    .B(_01114_));
 sg13g2_nor2_1 _21573_ (.A(_01103_),
    .B(_01115_),
    .Y(_01116_));
 sg13g2_a21oi_1 _21574_ (.A1(_11728_),
    .A2(_11731_),
    .Y(_01117_),
    .B1(_01096_));
 sg13g2_nand2_1 _21575_ (.Y(_01118_),
    .A(_01116_),
    .B(_01117_));
 sg13g2_nor3_1 _21576_ (.A(_01098_),
    .B(_11704_),
    .C(_01099_),
    .Y(_01119_));
 sg13g2_nor2b_1 _21577_ (.A(_01114_),
    .B_N(_01102_),
    .Y(_01120_));
 sg13g2_nor2_1 _21578_ (.A(_01119_),
    .B(_01120_),
    .Y(_01121_));
 sg13g2_nand2_1 _21579_ (.Y(_01123_),
    .A(_01118_),
    .B(_01121_));
 sg13g2_nand2_1 _21580_ (.Y(_01124_),
    .A(_01123_),
    .B(_01112_));
 sg13g2_inv_1 _21581_ (.Y(_01125_),
    .A(_01107_));
 sg13g2_nand3_1 _21582_ (.B(_01125_),
    .C(_01121_),
    .A(_01118_),
    .Y(_01126_));
 sg13g2_nand2_2 _21583_ (.Y(_01127_),
    .A(_01124_),
    .B(_01126_));
 sg13g2_xnor2_1 _21584_ (.Y(_01128_),
    .A(_08900_),
    .B(_01127_));
 sg13g2_nor2b_1 _21585_ (.A(_08893_),
    .B_N(_08892_),
    .Y(_01129_));
 sg13g2_inv_1 _21586_ (.Y(_01130_),
    .A(_01129_));
 sg13g2_nand2_1 _21587_ (.Y(_01131_),
    .A(_01101_),
    .B(_01098_));
 sg13g2_xnor2_1 _21588_ (.Y(_01132_),
    .A(_01130_),
    .B(_01131_));
 sg13g2_inv_1 _21589_ (.Y(_01134_),
    .A(_01132_));
 sg13g2_nand2_1 _21590_ (.Y(_01135_),
    .A(_11728_),
    .B(_11731_));
 sg13g2_nand3_1 _21591_ (.B(_01135_),
    .C(_01121_),
    .A(_01118_),
    .Y(_01136_));
 sg13g2_o21ai_1 _21592_ (.B1(_01096_),
    .Y(_01137_),
    .A1(_01119_),
    .A2(_01120_));
 sg13g2_nand2_1 _21593_ (.Y(_01138_),
    .A(_01136_),
    .B(_01137_));
 sg13g2_nand2_1 _21594_ (.Y(_01139_),
    .A(_08871_),
    .B(_08872_));
 sg13g2_nand2_1 _21595_ (.Y(_01140_),
    .A(_08898_),
    .B(_01139_));
 sg13g2_nand3_1 _21596_ (.B(_08897_),
    .C(_08884_),
    .A(_08896_),
    .Y(_01141_));
 sg13g2_nand2_1 _21597_ (.Y(_01142_),
    .A(_01140_),
    .B(_01141_));
 sg13g2_nor2b_1 _21598_ (.A(_01138_),
    .B_N(_01142_),
    .Y(_01143_));
 sg13g2_nor2_1 _21599_ (.A(_01134_),
    .B(_01143_),
    .Y(_01145_));
 sg13g2_a21oi_1 _21600_ (.A1(_01136_),
    .A2(_01137_),
    .Y(_01146_),
    .B1(_01142_));
 sg13g2_nand3_1 _21601_ (.B(_01145_),
    .C(_01146_),
    .A(_01128_),
    .Y(_01147_));
 sg13g2_buf_1 _21602_ (.A(_01147_),
    .X(_01148_));
 sg13g2_nor2_1 _21603_ (.A(_01129_),
    .B(_01131_),
    .Y(_01149_));
 sg13g2_inv_2 _21604_ (.Y(_01150_),
    .A(_01127_));
 sg13g2_nor3_1 _21605_ (.A(_08900_),
    .B(_01134_),
    .C(_01150_),
    .Y(_01151_));
 sg13g2_nor2_1 _21606_ (.A(_01149_),
    .B(_01151_),
    .Y(_01152_));
 sg13g2_nand2_1 _21607_ (.Y(_01153_),
    .A(_01148_),
    .B(_01152_));
 sg13g2_buf_8 _21608_ (.A(_01153_),
    .X(_01154_));
 sg13g2_nand2_1 _21609_ (.Y(_01156_),
    .A(_01154_),
    .B(_01142_));
 sg13g2_nand3_1 _21610_ (.B(_01138_),
    .C(_01152_),
    .A(_01148_),
    .Y(_01157_));
 sg13g2_buf_8 _21611_ (.A(_01157_),
    .X(_01158_));
 sg13g2_nand3_1 _21612_ (.B(_07225_),
    .C(_07765_),
    .A(_08817_),
    .Y(_01159_));
 sg13g2_o21ai_1 _21613_ (.B1(net165),
    .Y(_01160_),
    .A1(_01159_),
    .A2(_07594_));
 sg13g2_nor2_1 _21614_ (.A(_07227_),
    .B(_01160_),
    .Y(_01161_));
 sg13g2_nand2_1 _21615_ (.Y(_01162_),
    .A(_07548_),
    .B(_03839_));
 sg13g2_o21ai_1 _21616_ (.B1(_01162_),
    .Y(_01163_),
    .A1(_07239_),
    .A2(_08712_));
 sg13g2_nor2_1 _21617_ (.A(_04227_),
    .B(_04323_),
    .Y(_01164_));
 sg13g2_nor2_1 _21618_ (.A(_01163_),
    .B(_01164_),
    .Y(_01165_));
 sg13g2_inv_1 _21619_ (.Y(_01167_),
    .A(_01165_));
 sg13g2_a21oi_1 _21620_ (.A1(_06097_),
    .A2(net52),
    .Y(_01168_),
    .B1(_05698_));
 sg13g2_inv_1 _21621_ (.Y(_01169_),
    .A(_01168_));
 sg13g2_a21oi_1 _21622_ (.A1(_01169_),
    .A2(net39),
    .Y(_01170_),
    .B1(_08087_));
 sg13g2_inv_1 _21623_ (.Y(_01171_),
    .A(_01170_));
 sg13g2_a21oi_1 _21624_ (.A1(_01171_),
    .A2(_06199_),
    .Y(_01172_),
    .B1(_06611_));
 sg13g2_inv_1 _21625_ (.Y(_01173_),
    .A(_01172_));
 sg13g2_a21oi_1 _21626_ (.A1(_01173_),
    .A2(net66),
    .Y(_01174_),
    .B1(_06990_));
 sg13g2_o21ai_1 _21627_ (.B1(_07127_),
    .Y(_01175_),
    .A1(_04127_),
    .A2(_01174_));
 sg13g2_buf_1 _21628_ (.A(_01175_),
    .X(_01176_));
 sg13g2_a22oi_1 _21629_ (.Y(_01178_),
    .B1(_07239_),
    .B2(_08711_),
    .A2(_07548_),
    .A1(_04407_));
 sg13g2_nor2_1 _21630_ (.A(_04228_),
    .B(_04323_),
    .Y(_01179_));
 sg13g2_inv_1 _21631_ (.Y(_01180_),
    .A(_01179_));
 sg13g2_nand3_1 _21632_ (.B(_01178_),
    .C(_01180_),
    .A(_01176_),
    .Y(_01181_));
 sg13g2_o21ai_1 _21633_ (.B1(net165),
    .Y(_01182_),
    .A1(_01167_),
    .A2(_01181_));
 sg13g2_a21o_1 _21634_ (.A2(_01160_),
    .A1(_01182_),
    .B1(_04329_),
    .X(_01183_));
 sg13g2_nand3b_1 _21635_ (.B(_01183_),
    .C(_04239_),
    .Y(_01184_),
    .A_N(_01161_));
 sg13g2_nor2_1 _21636_ (.A(_05067_),
    .B(_07993_),
    .Y(_01185_));
 sg13g2_inv_1 _21637_ (.Y(_01186_),
    .A(_01185_));
 sg13g2_nor2_1 _21638_ (.A(_07720_),
    .B(net14),
    .Y(_01187_));
 sg13g2_nor2_1 _21639_ (.A(_07241_),
    .B(_04999_),
    .Y(_01188_));
 sg13g2_nand4_1 _21640_ (.B(_08698_),
    .C(_01188_),
    .A(_01187_),
    .Y(_01189_),
    .D(_04401_));
 sg13g2_nor2_1 _21641_ (.A(_01186_),
    .B(_01189_),
    .Y(_01190_));
 sg13g2_nor2_1 _21642_ (.A(_04442_),
    .B(_04134_),
    .Y(_01191_));
 sg13g2_nor4_1 _21643_ (.A(_07150_),
    .B(_05005_),
    .C(_07812_),
    .D(_05054_),
    .Y(_01192_));
 sg13g2_nand4_1 _21644_ (.B(_04978_),
    .C(_01191_),
    .A(_01190_),
    .Y(_01193_),
    .D(_01192_));
 sg13g2_nor2_1 _21645_ (.A(net63),
    .B(_04242_),
    .Y(_01194_));
 sg13g2_nand3_1 _21646_ (.B(_01193_),
    .C(_01194_),
    .A(_01184_),
    .Y(_01195_));
 sg13g2_a21oi_1 _21647_ (.A1(_05770_),
    .A2(net39),
    .Y(_01196_),
    .B1(_05436_));
 sg13g2_inv_1 _21648_ (.Y(_01197_),
    .A(_01196_));
 sg13g2_a21oi_1 _21649_ (.A1(_01197_),
    .A2(net21),
    .Y(_01199_),
    .B1(_06201_));
 sg13g2_inv_1 _21650_ (.Y(_01200_),
    .A(_01199_));
 sg13g2_a21oi_1 _21651_ (.A1(_01200_),
    .A2(_06735_),
    .Y(_01201_),
    .B1(_06737_));
 sg13g2_inv_1 _21652_ (.Y(_01202_),
    .A(_01201_));
 sg13g2_a21oi_1 _21653_ (.A1(_01202_),
    .A2(_04129_),
    .Y(_01203_),
    .B1(_04131_));
 sg13g2_inv_1 _21654_ (.Y(_01204_),
    .A(_01203_));
 sg13g2_nor2_1 _21655_ (.A(_01176_),
    .B(_01204_),
    .Y(_01205_));
 sg13g2_nand2_1 _21656_ (.Y(_01206_),
    .A(_04998_),
    .B(_08816_));
 sg13g2_nor2_1 _21657_ (.A(_07765_),
    .B(_04440_),
    .Y(_01207_));
 sg13g2_nor4_1 _21658_ (.A(_01207_),
    .B(_00932_),
    .C(_08699_),
    .D(_05006_),
    .Y(_01208_));
 sg13g2_nor2_1 _21659_ (.A(_07165_),
    .B(_07830_),
    .Y(_01210_));
 sg13g2_nand3_1 _21660_ (.B(_01210_),
    .C(_08973_),
    .A(_06647_),
    .Y(_01211_));
 sg13g2_inv_1 _21661_ (.Y(_01212_),
    .A(_01211_));
 sg13g2_and4_1 _21662_ (.A(_01206_),
    .B(_01208_),
    .C(_01212_),
    .D(_01178_),
    .X(_01213_));
 sg13g2_o21ai_1 _21663_ (.B1(_01213_),
    .Y(_01214_),
    .A1(_07595_),
    .A2(_07605_));
 sg13g2_nor3_1 _21664_ (.A(_01186_),
    .B(_01179_),
    .C(_01214_),
    .Y(_01215_));
 sg13g2_nand3b_1 _21665_ (.B(_01215_),
    .C(_01192_),
    .Y(_01216_),
    .A_N(_01205_));
 sg13g2_o21ai_1 _21666_ (.B1(_07247_),
    .Y(_01217_),
    .A1(_06630_),
    .A2(_06634_));
 sg13g2_nor4_1 _21667_ (.A(_00909_),
    .B(_08734_),
    .C(_09007_),
    .D(_01217_),
    .Y(_01218_));
 sg13g2_nor2_1 _21668_ (.A(_07765_),
    .B(_04441_),
    .Y(_01219_));
 sg13g2_nor4_1 _21669_ (.A(_01219_),
    .B(_07735_),
    .C(_06641_),
    .D(_04408_),
    .Y(_01221_));
 sg13g2_nand4_1 _21670_ (.B(_01218_),
    .C(_01188_),
    .A(_01187_),
    .Y(_01222_),
    .D(_01221_));
 sg13g2_nor2_1 _21671_ (.A(_01176_),
    .B(_01203_),
    .Y(_01223_));
 sg13g2_inv_1 _21672_ (.Y(_01224_),
    .A(_04998_));
 sg13g2_a22oi_1 _21673_ (.Y(_01225_),
    .B1(_07594_),
    .B2(_07605_),
    .A2(_08816_),
    .A1(_01224_));
 sg13g2_nand3b_1 _21674_ (.B(_01225_),
    .C(_01191_),
    .Y(_01226_),
    .A_N(_01223_));
 sg13g2_nor3_1 _21675_ (.A(_01167_),
    .B(_01222_),
    .C(_01226_),
    .Y(_01227_));
 sg13g2_nand2b_1 _21676_ (.Y(_01228_),
    .B(_01227_),
    .A_N(_01216_));
 sg13g2_o21ai_1 _21677_ (.B1(_04235_),
    .Y(_01229_),
    .A1(_04232_),
    .A2(_04241_));
 sg13g2_nand3_1 _21678_ (.B(_05091_),
    .C(_01229_),
    .A(_01228_),
    .Y(_01230_));
 sg13g2_nor2_1 _21679_ (.A(net165),
    .B(_01227_),
    .Y(_01232_));
 sg13g2_nand3_1 _21680_ (.B(net114),
    .C(_01216_),
    .A(_01232_),
    .Y(_01233_));
 sg13g2_nand2b_1 _21681_ (.Y(_01234_),
    .B(_07226_),
    .A_N(_01233_));
 sg13g2_nand3_1 _21682_ (.B(_01230_),
    .C(_01234_),
    .A(_01195_),
    .Y(_01235_));
 sg13g2_buf_1 _21683_ (.A(\b.gen_square[46].sq.mask ),
    .X(_01236_));
 sg13g2_nand2_1 _21684_ (.Y(_01237_),
    .A(_01235_),
    .B(_01236_));
 sg13g2_nand2b_1 _21685_ (.Y(_01238_),
    .B(_05050_),
    .A_N(_07876_));
 sg13g2_o21ai_1 _21686_ (.B1(_01238_),
    .Y(_01239_),
    .A1(_04121_),
    .A2(_06870_));
 sg13g2_a221oi_1 _21687_ (.B2(_04939_),
    .C1(_01239_),
    .B1(_04974_),
    .A1(_08716_),
    .Y(_01240_),
    .A2(_08648_));
 sg13g2_a21oi_1 _21688_ (.A1(_07547_),
    .A2(_04247_),
    .Y(_01241_),
    .B1(_04333_));
 sg13g2_a21oi_1 _21689_ (.A1(_04480_),
    .A2(_04247_),
    .Y(_01243_),
    .B1(_04251_));
 sg13g2_inv_1 _21690_ (.Y(_01244_),
    .A(_01243_));
 sg13g2_a22oi_1 _21691_ (.Y(_01245_),
    .B1(_01241_),
    .B2(_01244_),
    .A2(_07791_),
    .A1(_07794_));
 sg13g2_a22oi_1 _21692_ (.Y(_01246_),
    .B1(_07123_),
    .B2(_07145_),
    .A2(_01174_),
    .A1(_01202_));
 sg13g2_nor4_1 _21693_ (.A(_07934_),
    .B(_04585_),
    .C(_08106_),
    .D(_06296_),
    .Y(_01247_));
 sg13g2_nor4_1 _21694_ (.A(_08673_),
    .B(_07030_),
    .C(_07926_),
    .D(_04567_),
    .Y(_01248_));
 sg13g2_and2_1 _21695_ (.A(_01247_),
    .B(_01248_),
    .X(_01249_));
 sg13g2_nand4_1 _21696_ (.B(_01245_),
    .C(_01246_),
    .A(_01240_),
    .Y(_01250_),
    .D(_01249_));
 sg13g2_inv_1 _21697_ (.Y(_01251_),
    .A(_07880_));
 sg13g2_nor2_1 _21698_ (.A(_07149_),
    .B(_01251_),
    .Y(_01252_));
 sg13g2_inv_1 _21699_ (.Y(_01254_),
    .A(_01252_));
 sg13g2_nand4_1 _21700_ (.B(_07258_),
    .C(_01254_),
    .A(_05000_),
    .Y(_01255_),
    .D(_07721_));
 sg13g2_nor4_1 _21701_ (.A(net14),
    .B(_06795_),
    .C(_07707_),
    .D(_01255_),
    .Y(_01256_));
 sg13g2_nor2b_1 _21702_ (.A(_01250_),
    .B_N(_01256_),
    .Y(_01257_));
 sg13g2_nor2_1 _21703_ (.A(_06900_),
    .B(_06461_),
    .Y(_01258_));
 sg13g2_nor2_1 _21704_ (.A(_05017_),
    .B(_05016_),
    .Y(_01259_));
 sg13g2_nor2_1 _21705_ (.A(_08664_),
    .B(_07911_),
    .Y(_01260_));
 sg13g2_nand4_1 _21706_ (.B(_01258_),
    .C(_01259_),
    .A(_09151_),
    .Y(_01261_),
    .D(_01260_));
 sg13g2_a22oi_1 _21707_ (.Y(_01262_),
    .B1(_07123_),
    .B2(_07144_),
    .A2(_01241_),
    .A1(_01243_));
 sg13g2_a22oi_1 _21708_ (.Y(_01263_),
    .B1(_01174_),
    .B2(_01201_),
    .A2(_07791_),
    .A1(_07793_));
 sg13g2_nand2_1 _21709_ (.Y(_01265_),
    .A(_01262_),
    .B(_01263_));
 sg13g2_nand2_1 _21710_ (.Y(_01266_),
    .A(_08715_),
    .B(_08648_));
 sg13g2_o21ai_1 _21711_ (.B1(_01266_),
    .Y(_01267_),
    .A1(_07880_),
    .A2(_07876_));
 sg13g2_a221oi_1 _21712_ (.B2(_04939_),
    .C1(_01267_),
    .B1(_04973_),
    .A1(_06869_),
    .Y(_01268_),
    .A2(_04121_));
 sg13g2_nand2b_1 _21713_ (.Y(_01269_),
    .B(_01268_),
    .A_N(_01265_));
 sg13g2_nor4_1 _21714_ (.A(_06830_),
    .B(_07150_),
    .C(_07812_),
    .D(_07809_),
    .Y(_01270_));
 sg13g2_inv_1 _21715_ (.Y(_01271_),
    .A(_07993_));
 sg13g2_nand4_1 _21716_ (.B(_01271_),
    .C(_08460_),
    .A(_01270_),
    .Y(_01272_),
    .D(_05068_));
 sg13g2_nor3_1 _21717_ (.A(_01261_),
    .B(_01269_),
    .C(_01272_),
    .Y(_01273_));
 sg13g2_nor3_1 _21718_ (.A(_04041_),
    .B(_01257_),
    .C(_01273_),
    .Y(_01274_));
 sg13g2_nand2_1 _21719_ (.Y(_01276_),
    .A(_01274_),
    .B(net114));
 sg13g2_nand2_1 _21720_ (.Y(_01277_),
    .A(_01273_),
    .B(_01257_));
 sg13g2_nand3_1 _21721_ (.B(net68),
    .C(_04042_),
    .A(_01277_),
    .Y(_01278_));
 sg13g2_nand2_1 _21722_ (.Y(_01279_),
    .A(_01276_),
    .B(_01278_));
 sg13g2_nand2_1 _21723_ (.Y(_01280_),
    .A(_01276_),
    .B(_04125_));
 sg13g2_nand2b_1 _21724_ (.Y(_01281_),
    .B(_04124_),
    .A_N(_04942_));
 sg13g2_nand3_1 _21725_ (.B(_01280_),
    .C(_01281_),
    .A(_01279_),
    .Y(_01282_));
 sg13g2_nand2_1 _21726_ (.Y(_01283_),
    .A(_01246_),
    .B(_01245_));
 sg13g2_o21ai_1 _21727_ (.B1(_04041_),
    .Y(_01284_),
    .A1(_01265_),
    .A2(_01283_));
 sg13g2_nor3_1 _21728_ (.A(_04055_),
    .B(_04124_),
    .C(_01284_),
    .Y(_01285_));
 sg13g2_a21o_1 _21729_ (.A2(_01268_),
    .A1(_01240_),
    .B1(_04042_),
    .X(_01287_));
 sg13g2_a21o_1 _21730_ (.A2(_01284_),
    .A1(_01287_),
    .B1(_04943_),
    .X(_01288_));
 sg13g2_nand2b_1 _21731_ (.Y(_01289_),
    .B(_01288_),
    .A_N(_01285_));
 sg13g2_nand2_1 _21732_ (.Y(_01290_),
    .A(_01289_),
    .B(net67));
 sg13g2_inv_1 _21733_ (.Y(_01291_),
    .A(\b.gen_square[45].sq.mask ));
 sg13g2_a21o_1 _21734_ (.A2(_01290_),
    .A1(_01282_),
    .B1(_01291_),
    .X(_01292_));
 sg13g2_buf_1 _21735_ (.A(_01292_),
    .X(_01293_));
 sg13g2_inv_1 _21736_ (.Y(_01294_),
    .A(\b.gen_square[41].sq.mask ));
 sg13g2_inv_1 _21737_ (.Y(_01295_),
    .A(_08306_));
 sg13g2_inv_1 _21738_ (.Y(_01296_),
    .A(_01241_));
 sg13g2_inv_1 _21739_ (.Y(_01298_),
    .A(_07127_));
 sg13g2_a21oi_1 _21740_ (.A1(_01296_),
    .A2(net71),
    .Y(_01299_),
    .B1(_01298_));
 sg13g2_o21ai_1 _21741_ (.B1(_06989_),
    .Y(_01300_),
    .A1(_06662_),
    .A2(_01299_));
 sg13g2_a21oi_1 _21742_ (.A1(_01300_),
    .A2(_06198_),
    .Y(_01301_),
    .B1(_06611_));
 sg13g2_inv_1 _21743_ (.Y(_01302_),
    .A(_01301_));
 sg13g2_a21oi_2 _21744_ (.B1(_08087_),
    .Y(_01303_),
    .A2(net39),
    .A1(_01302_));
 sg13g2_a21oi_1 _21745_ (.A1(_01244_),
    .A2(net71),
    .Y(_01304_),
    .B1(_04131_));
 sg13g2_o21ai_1 _21746_ (.B1(_07014_),
    .Y(_01305_),
    .A1(_06662_),
    .A2(_01304_));
 sg13g2_a21oi_1 _21747_ (.A1(_01305_),
    .A2(_06198_),
    .Y(_01306_),
    .B1(_06201_));
 sg13g2_o21ai_1 _21748_ (.B1(_05759_),
    .Y(_01307_),
    .A1(_05757_),
    .A2(_01306_));
 sg13g2_buf_1 _21749_ (.A(_01307_),
    .X(_01309_));
 sg13g2_inv_1 _21750_ (.Y(_01310_),
    .A(_01309_));
 sg13g2_a22oi_1 _21751_ (.Y(_01311_),
    .B1(_01303_),
    .B2(_01310_),
    .A2(_01295_),
    .A1(_05944_));
 sg13g2_a22oi_1 _21752_ (.Y(_01312_),
    .B1(_01303_),
    .B2(_01309_),
    .A2(_05689_),
    .A1(_05725_));
 sg13g2_inv_1 _21753_ (.Y(_01313_),
    .A(_06097_));
 sg13g2_a22oi_1 _21754_ (.Y(_01314_),
    .B1(_05689_),
    .B2(_05724_),
    .A2(_01313_),
    .A1(_05498_));
 sg13g2_a22oi_1 _21755_ (.Y(_01315_),
    .B1(_01295_),
    .B2(_05943_),
    .A2(_01313_),
    .A1(_05500_));
 sg13g2_nand4_1 _21756_ (.B(_01312_),
    .C(_01314_),
    .A(_01311_),
    .Y(_01316_),
    .D(_01315_));
 sg13g2_nand2_1 _21757_ (.Y(_01317_),
    .A(_01316_),
    .B(net190));
 sg13g2_nor2_1 _21758_ (.A(_08153_),
    .B(_08216_),
    .Y(_01318_));
 sg13g2_inv_1 _21759_ (.Y(_01320_),
    .A(_01318_));
 sg13g2_nand3_1 _21760_ (.B(_08028_),
    .C(_06306_),
    .A(_01320_),
    .Y(_01321_));
 sg13g2_nor2_1 _21761_ (.A(_05923_),
    .B(_05964_),
    .Y(_01322_));
 sg13g2_inv_1 _21762_ (.Y(_01323_),
    .A(_05923_));
 sg13g2_a22oi_1 _21763_ (.Y(_01324_),
    .B1(_05964_),
    .B2(_01323_),
    .A2(_08152_),
    .A1(_08216_));
 sg13g2_nand2b_1 _21764_ (.Y(_01325_),
    .B(_01324_),
    .A_N(_01322_));
 sg13g2_o21ai_1 _21765_ (.B1(net190),
    .Y(_01326_),
    .A1(_01321_),
    .A2(_01325_));
 sg13g2_a21o_1 _21766_ (.A2(_01326_),
    .A1(_01317_),
    .B1(_05694_),
    .X(_01327_));
 sg13g2_nand2b_1 _21767_ (.Y(_01328_),
    .B(_05924_),
    .A_N(_01326_));
 sg13g2_nand3_1 _21768_ (.B(_05552_),
    .C(_01328_),
    .A(_01327_),
    .Y(_01329_));
 sg13g2_nor4_1 _21769_ (.A(_05768_),
    .B(_06123_),
    .C(_08061_),
    .D(_05763_),
    .Y(_01330_));
 sg13g2_nor2_1 _21770_ (.A(_05945_),
    .B(_05439_),
    .Y(_01331_));
 sg13g2_nand3_1 _21771_ (.B(_05553_),
    .C(_05506_),
    .A(_08342_),
    .Y(_01332_));
 sg13g2_nor2_1 _21772_ (.A(_05546_),
    .B(_08094_),
    .Y(_01333_));
 sg13g2_inv_1 _21773_ (.Y(_01334_),
    .A(_01333_));
 sg13g2_nor3_1 _21774_ (.A(_08502_),
    .B(_01332_),
    .C(_01334_),
    .Y(_01335_));
 sg13g2_nand3_1 _21775_ (.B(_01331_),
    .C(_01335_),
    .A(_01330_),
    .Y(_01336_));
 sg13g2_nor2_1 _21776_ (.A(net120),
    .B(_05558_),
    .Y(_01337_));
 sg13g2_nand3_1 _21777_ (.B(_01336_),
    .C(_01337_),
    .A(_01329_),
    .Y(_01338_));
 sg13g2_nor2_1 _21778_ (.A(_08028_),
    .B(_04608_),
    .Y(_01339_));
 sg13g2_inv_1 _21779_ (.Y(_01341_),
    .A(_05776_));
 sg13g2_o21ai_1 _21780_ (.B1(_01341_),
    .Y(_01342_),
    .A1(_08342_),
    .A2(_06893_));
 sg13g2_and3_1 _21781_ (.X(_01343_),
    .A(_08053_),
    .B(_07923_),
    .C(_06462_));
 sg13g2_nand2_1 _21782_ (.Y(_01344_),
    .A(_11099_),
    .B(_05824_));
 sg13g2_nor2_1 _21783_ (.A(_11931_),
    .B(_01344_),
    .Y(_01345_));
 sg13g2_nand4_1 _21784_ (.B(_01345_),
    .C(_11886_),
    .A(_01343_),
    .Y(_01346_),
    .D(_06125_));
 sg13g2_nand2_1 _21785_ (.Y(_01347_),
    .A(_01314_),
    .B(_01324_));
 sg13g2_nor4_1 _21786_ (.A(_01339_),
    .B(_01342_),
    .C(_01346_),
    .D(_01347_),
    .Y(_01348_));
 sg13g2_and3_1 _21787_ (.X(_01349_),
    .A(_01348_),
    .B(_01311_),
    .C(_01330_));
 sg13g2_nor2_1 _21788_ (.A(_07926_),
    .B(_06296_),
    .Y(_01350_));
 sg13g2_nor2_1 _21789_ (.A(_08028_),
    .B(_04607_),
    .Y(_01352_));
 sg13g2_inv_1 _21790_ (.Y(_01353_),
    .A(_01352_));
 sg13g2_nand2_1 _21791_ (.Y(_01354_),
    .A(_01350_),
    .B(_01353_));
 sg13g2_nor2_1 _21792_ (.A(_06285_),
    .B(_05831_),
    .Y(_01355_));
 sg13g2_nor2b_1 _21793_ (.A(_09389_),
    .B_N(_01355_),
    .Y(_01356_));
 sg13g2_nand2b_1 _21794_ (.Y(_01357_),
    .B(_01356_),
    .A_N(_05513_));
 sg13g2_nor4_1 _21795_ (.A(_11935_),
    .B(_08323_),
    .C(_01354_),
    .D(_01357_),
    .Y(_01358_));
 sg13g2_nand3_1 _21796_ (.B(_01315_),
    .C(_01320_),
    .A(_01358_),
    .Y(_01359_));
 sg13g2_nor3_1 _21797_ (.A(_08345_),
    .B(_01359_),
    .C(_01322_),
    .Y(_01360_));
 sg13g2_and4_1 _21798_ (.A(_01333_),
    .B(_01312_),
    .C(_01331_),
    .D(_01360_),
    .X(_01361_));
 sg13g2_nand2_1 _21799_ (.Y(_01363_),
    .A(_01349_),
    .B(_01361_));
 sg13g2_o21ai_1 _21800_ (.B1(_05566_),
    .Y(_01364_),
    .A1(_05550_),
    .A2(net190));
 sg13g2_nand3_1 _21801_ (.B(net129),
    .C(_01364_),
    .A(_01363_),
    .Y(_01365_));
 sg13g2_nor3_1 _21802_ (.A(net190),
    .B(_01361_),
    .C(_01349_),
    .Y(_01366_));
 sg13g2_nand3_1 _21803_ (.B(net177),
    .C(_06615_),
    .A(_01366_),
    .Y(_01367_));
 sg13g2_nand3_1 _21804_ (.B(_01365_),
    .C(_01367_),
    .A(_01338_),
    .Y(_01368_));
 sg13g2_nor2b_1 _21805_ (.A(_01294_),
    .B_N(_01368_),
    .Y(_01369_));
 sg13g2_inv_1 _21806_ (.Y(_01370_),
    .A(_08184_));
 sg13g2_inv_1 _21807_ (.Y(_01371_),
    .A(_01303_));
 sg13g2_a21oi_1 _21808_ (.A1(_01371_),
    .A2(net52),
    .Y(_01372_),
    .B1(_05698_));
 sg13g2_a21oi_1 _21809_ (.A1(_01309_),
    .A2(net52),
    .Y(_01374_),
    .B1(_05571_));
 sg13g2_a22oi_1 _21810_ (.Y(_01375_),
    .B1(_01372_),
    .B2(_01374_),
    .A2(_01370_),
    .A1(_08222_));
 sg13g2_inv_1 _21811_ (.Y(_01376_),
    .A(_08061_));
 sg13g2_nor2_1 _21812_ (.A(_03859_),
    .B(_04625_),
    .Y(_01377_));
 sg13g2_a21oi_1 _21813_ (.A1(_05501_),
    .A2(_04625_),
    .Y(_01378_),
    .B1(_01377_));
 sg13g2_nor2_1 _21814_ (.A(_05941_),
    .B(_01378_),
    .Y(_01379_));
 sg13g2_inv_1 _21815_ (.Y(_01380_),
    .A(_01379_));
 sg13g2_inv_1 _21816_ (.Y(_01381_),
    .A(_08222_));
 sg13g2_nor2_1 _21817_ (.A(_05506_),
    .B(_01381_),
    .Y(_01382_));
 sg13g2_nor2_1 _21818_ (.A(_08352_),
    .B(_01382_),
    .Y(_01383_));
 sg13g2_nand3_1 _21819_ (.B(_01380_),
    .C(_01383_),
    .A(_01376_),
    .Y(_01385_));
 sg13g2_a21oi_1 _21820_ (.A1(_01374_),
    .A2(_06121_),
    .Y(_01386_),
    .B1(_01385_));
 sg13g2_a21oi_1 _21821_ (.A1(_08355_),
    .A2(net74),
    .Y(_01387_),
    .B1(_05723_));
 sg13g2_a21oi_1 _21822_ (.A1(_08291_),
    .A2(net74),
    .Y(_01388_),
    .B1(_06755_));
 sg13g2_a21oi_1 _21823_ (.A1(_05491_),
    .A2(net87),
    .Y(_01389_),
    .B1(_01377_));
 sg13g2_a21o_1 _21824_ (.A2(_04626_),
    .A1(_05231_),
    .B1(_08380_),
    .X(_01390_));
 sg13g2_buf_1 _21825_ (.A(_01390_),
    .X(_01391_));
 sg13g2_inv_1 _21826_ (.Y(_01392_),
    .A(_06649_));
 sg13g2_nor3_1 _21827_ (.A(_08268_),
    .B(_08423_),
    .C(_01392_),
    .Y(_01393_));
 sg13g2_o21ai_1 _21828_ (.B1(_01393_),
    .Y(_01394_),
    .A1(_01389_),
    .A2(_01391_));
 sg13g2_a221oi_1 _21829_ (.B2(_01388_),
    .C1(_01394_),
    .B1(_01387_),
    .A1(_06091_),
    .Y(_01396_),
    .A2(_06116_));
 sg13g2_and3_1 _21830_ (.X(_01397_),
    .A(_01375_),
    .B(_01386_),
    .C(_01396_));
 sg13g2_inv_1 _21831_ (.Y(_01398_),
    .A(_01374_));
 sg13g2_a22oi_1 _21832_ (.Y(_01399_),
    .B1(_01372_),
    .B2(_01398_),
    .A2(_01370_),
    .A1(_01381_));
 sg13g2_nor2_1 _21833_ (.A(_05506_),
    .B(_08222_),
    .Y(_01400_));
 sg13g2_inv_1 _21834_ (.Y(_01401_),
    .A(_01378_));
 sg13g2_nor2_1 _21835_ (.A(_05941_),
    .B(_01401_),
    .Y(_01402_));
 sg13g2_inv_1 _21836_ (.Y(_01403_),
    .A(_01402_));
 sg13g2_nand2_1 _21837_ (.Y(_01404_),
    .A(_01403_),
    .B(_08549_));
 sg13g2_nor4_1 _21838_ (.A(_01400_),
    .B(_05573_),
    .C(_08323_),
    .D(_01404_),
    .Y(_01405_));
 sg13g2_inv_1 _21839_ (.Y(_01407_),
    .A(_01389_));
 sg13g2_nor2_1 _21840_ (.A(_01407_),
    .B(_01391_),
    .Y(_01408_));
 sg13g2_nor4_1 _21841_ (.A(_06629_),
    .B(_08257_),
    .C(_05146_),
    .D(_08418_),
    .Y(_01409_));
 sg13g2_inv_1 _21842_ (.Y(_01410_),
    .A(_01409_));
 sg13g2_nor2_1 _21843_ (.A(_06116_),
    .B(_06092_),
    .Y(_01411_));
 sg13g2_inv_1 _21844_ (.Y(_01412_),
    .A(_01388_));
 sg13g2_nor2_1 _21845_ (.A(_01412_),
    .B(_01387_),
    .Y(_01413_));
 sg13g2_nor4_1 _21846_ (.A(_01408_),
    .B(_01410_),
    .C(_01411_),
    .D(_01413_),
    .Y(_01414_));
 sg13g2_and3_1 _21847_ (.X(_01415_),
    .A(_01399_),
    .B(_01405_),
    .C(_01414_));
 sg13g2_nor3_1 _21848_ (.A(_05233_),
    .B(_01397_),
    .C(_01415_),
    .Y(_01416_));
 sg13g2_nand2_1 _21849_ (.Y(_01418_),
    .A(_01416_),
    .B(net177));
 sg13g2_nand2_1 _21850_ (.Y(_01419_),
    .A(_01415_),
    .B(_01397_));
 sg13g2_nand3_1 _21851_ (.B(net144),
    .C(_05508_),
    .A(_01419_),
    .Y(_01420_));
 sg13g2_nand2_1 _21852_ (.Y(_01421_),
    .A(_01418_),
    .B(_01420_));
 sg13g2_nand2_1 _21853_ (.Y(_01422_),
    .A(_01418_),
    .B(_05496_));
 sg13g2_nand2_1 _21854_ (.Y(_01423_),
    .A(_05239_),
    .B(_05495_));
 sg13g2_nand3_1 _21855_ (.B(_01422_),
    .C(_01423_),
    .A(_01421_),
    .Y(_01424_));
 sg13g2_a21oi_1 _21856_ (.A1(_01412_),
    .A2(_01391_),
    .Y(_01425_),
    .B1(_05508_));
 sg13g2_nor2b_1 _21857_ (.A(_06091_),
    .B_N(_01375_),
    .Y(_01426_));
 sg13g2_a21oi_1 _21858_ (.A1(_01426_),
    .A2(_01399_),
    .Y(_01427_),
    .B1(_05508_));
 sg13g2_o21ai_1 _21859_ (.B1(_05240_),
    .Y(_01429_),
    .A1(_01425_),
    .A2(_01427_));
 sg13g2_nand3_1 _21860_ (.B(_05235_),
    .C(_06094_),
    .A(_01427_),
    .Y(_01430_));
 sg13g2_nand2_1 _21861_ (.Y(_01431_),
    .A(_01429_),
    .B(_01430_));
 sg13g2_nand2_1 _21862_ (.Y(_01432_),
    .A(_01431_),
    .B(net143));
 sg13g2_buf_1 _21863_ (.A(\b.gen_square[40].sq.mask ),
    .X(_01433_));
 sg13g2_inv_1 _21864_ (.Y(_01434_),
    .A(_01433_));
 sg13g2_a21o_1 _21865_ (.A2(_01432_),
    .A1(_01424_),
    .B1(_01434_),
    .X(_01435_));
 sg13g2_buf_1 _21866_ (.A(_01435_),
    .X(_01436_));
 sg13g2_nand2_1 _21867_ (.Y(_01437_),
    .A(_01366_),
    .B(net177));
 sg13g2_nand3_1 _21868_ (.B(net144),
    .C(_05556_),
    .A(_01363_),
    .Y(_01438_));
 sg13g2_nand2_1 _21869_ (.Y(_01439_),
    .A(_01437_),
    .B(_01438_));
 sg13g2_nand2_1 _21870_ (.Y(_01440_),
    .A(_01437_),
    .B(_05565_));
 sg13g2_nand2b_1 _21871_ (.Y(_01441_),
    .B(_05564_),
    .A_N(_05693_));
 sg13g2_nand3_1 _21872_ (.B(_01440_),
    .C(_01441_),
    .A(_01439_),
    .Y(_01442_));
 sg13g2_nand3_1 _21873_ (.B(net190),
    .C(_05692_),
    .A(_01316_),
    .Y(_01443_));
 sg13g2_nand2_1 _21874_ (.Y(_01444_),
    .A(_01327_),
    .B(_01443_));
 sg13g2_nand2_1 _21875_ (.Y(_01445_),
    .A(_01444_),
    .B(net128));
 sg13g2_a21o_1 _21876_ (.A2(_01445_),
    .A1(_01442_),
    .B1(_01294_),
    .X(_01446_));
 sg13g2_inv_1 _21877_ (.Y(_01447_),
    .A(_01446_));
 sg13g2_nand2_1 _21878_ (.Y(_01448_),
    .A(_01436_),
    .B(_01447_));
 sg13g2_nor2b_1 _21879_ (.A(_01344_),
    .B_N(_01350_),
    .Y(_01450_));
 sg13g2_and3_1 _21880_ (.X(_01451_),
    .A(_01343_),
    .B(_01356_),
    .C(_01450_));
 sg13g2_o21ai_1 _21881_ (.B1(_01328_),
    .Y(_01452_),
    .A1(_06617_),
    .A2(_01451_));
 sg13g2_o21ai_1 _21882_ (.B1(net143),
    .Y(_01453_),
    .A1(_01452_),
    .A2(_01444_));
 sg13g2_xnor2_1 _21883_ (.Y(_01454_),
    .A(_05549_),
    .B(_05693_));
 sg13g2_nand2_1 _21884_ (.Y(_01455_),
    .A(_01439_),
    .B(_01454_));
 sg13g2_a21o_1 _21885_ (.A2(_01455_),
    .A1(_01453_),
    .B1(_01294_),
    .X(_01456_));
 sg13g2_buf_1 _21886_ (.A(_01456_),
    .X(_01457_));
 sg13g2_a21oi_1 _21887_ (.A1(_01409_),
    .A2(_01393_),
    .Y(_01458_),
    .B1(_06286_));
 sg13g2_nand2b_1 _21888_ (.Y(_01459_),
    .B(_01425_),
    .A_N(_05243_));
 sg13g2_nand2b_1 _21889_ (.Y(_01461_),
    .B(_01459_),
    .A_N(_01458_));
 sg13g2_o21ai_1 _21890_ (.B1(net143),
    .Y(_01462_),
    .A1(_01461_),
    .A2(_01431_));
 sg13g2_nor2_1 _21891_ (.A(_05234_),
    .B(_05238_),
    .Y(_01463_));
 sg13g2_o21ai_1 _21892_ (.B1(_01421_),
    .Y(_01464_),
    .A1(_05240_),
    .A2(_01463_));
 sg13g2_nand2_1 _21893_ (.Y(_01465_),
    .A(_01462_),
    .B(_01464_));
 sg13g2_nand2_1 _21894_ (.Y(_01466_),
    .A(_01465_),
    .B(_01433_));
 sg13g2_xor2_1 _21895_ (.B(_01466_),
    .A(_01457_),
    .X(_01467_));
 sg13g2_nand2b_1 _21896_ (.Y(_01468_),
    .B(_01466_),
    .A_N(_01457_));
 sg13g2_o21ai_1 _21897_ (.B1(_01468_),
    .Y(_01469_),
    .A1(_01448_),
    .A2(_01467_));
 sg13g2_xnor2_1 _21898_ (.Y(_01470_),
    .A(_01447_),
    .B(_01436_));
 sg13g2_nor2_1 _21899_ (.A(_01467_),
    .B(_01470_),
    .Y(_01472_));
 sg13g2_o21ai_1 _21900_ (.B1(_06098_),
    .Y(_01473_),
    .A1(_05237_),
    .A2(_05233_));
 sg13g2_nand3_1 _21901_ (.B(net129),
    .C(_01473_),
    .A(_01419_),
    .Y(_01474_));
 sg13g2_o21ai_1 _21902_ (.B1(_01474_),
    .Y(_01475_),
    .A1(_05237_),
    .A2(_01418_));
 sg13g2_a21oi_1 _21903_ (.A1(_01386_),
    .A2(_01405_),
    .Y(_01476_),
    .B1(_05508_));
 sg13g2_nand3_1 _21904_ (.B(_05247_),
    .C(_01459_),
    .A(_01429_),
    .Y(_01477_));
 sg13g2_o21ai_1 _21905_ (.B1(_01477_),
    .Y(_01478_),
    .A1(_05247_),
    .A2(_01476_));
 sg13g2_nor2_1 _21906_ (.A(net103),
    .B(_01478_),
    .Y(_01479_));
 sg13g2_o21ai_1 _21907_ (.B1(_01433_),
    .Y(_01480_),
    .A1(_01475_),
    .A2(_01479_));
 sg13g2_nand3_1 _21908_ (.B(_01480_),
    .C(_01369_),
    .A(_01472_),
    .Y(_01481_));
 sg13g2_nor2b_1 _21909_ (.A(_01469_),
    .B_N(_01481_),
    .Y(_01482_));
 sg13g2_buf_1 _21910_ (.A(_01482_),
    .X(_01483_));
 sg13g2_nand2_1 _21911_ (.Y(_01484_),
    .A(_01483_),
    .B(_01480_));
 sg13g2_o21ai_1 _21912_ (.B1(_01484_),
    .Y(_01485_),
    .A1(_01369_),
    .A2(_01483_));
 sg13g2_nor2_1 _21913_ (.A(net103),
    .B(_05400_),
    .Y(_01486_));
 sg13g2_or2_1 _21914_ (.X(_01487_),
    .B(_07735_),
    .A(_08254_));
 sg13g2_inv_1 _21915_ (.Y(_01488_),
    .A(_06641_));
 sg13g2_inv_1 _21916_ (.Y(_01489_),
    .A(_05163_));
 sg13g2_nand4_1 _21917_ (.B(_01488_),
    .C(_05202_),
    .A(_07759_),
    .Y(_01490_),
    .D(_01489_));
 sg13g2_nor4_1 _21918_ (.A(_01487_),
    .B(_08418_),
    .C(_06629_),
    .D(_01490_),
    .Y(_01491_));
 sg13g2_nor2_1 _21919_ (.A(_05209_),
    .B(_07835_),
    .Y(_01493_));
 sg13g2_nand2_1 _21920_ (.Y(_01494_),
    .A(_01493_),
    .B(_08424_));
 sg13g2_nor4_1 _21921_ (.A(_08272_),
    .B(_06648_),
    .C(_11835_),
    .D(_01494_),
    .Y(_01495_));
 sg13g2_a21oi_1 _21922_ (.A1(_01491_),
    .A2(_01495_),
    .Y(_01496_),
    .B1(_05817_));
 sg13g2_nand2_1 _21923_ (.Y(_01497_),
    .A(_08319_),
    .B(_08292_));
 sg13g2_o21ai_1 _21924_ (.B1(_01497_),
    .Y(_01498_),
    .A1(_05433_),
    .A2(_08382_));
 sg13g2_a221oi_1 _21925_ (.B2(_05388_),
    .C1(_01498_),
    .B1(_05538_),
    .A1(_06756_),
    .Y(_01499_),
    .A2(_06744_));
 sg13g2_a22oi_1 _21926_ (.Y(_01500_),
    .B1(_08292_),
    .B2(_08320_),
    .A2(_08381_),
    .A1(_05433_));
 sg13g2_o21ai_1 _21927_ (.B1(_01500_),
    .Y(_01501_),
    .A1(_06757_),
    .A2(_06744_));
 sg13g2_a21oi_1 _21928_ (.A1(_05539_),
    .A2(_05388_),
    .Y(_01502_),
    .B1(_01501_));
 sg13g2_a21oi_1 _21929_ (.A1(_01499_),
    .A2(_01502_),
    .Y(_01504_),
    .B1(_05409_));
 sg13g2_nand2b_1 _21930_ (.Y(_01505_),
    .B(_01504_),
    .A_N(_05411_));
 sg13g2_nand2b_1 _21931_ (.Y(_01506_),
    .B(_01505_),
    .A_N(_01496_));
 sg13g2_xnor2_1 _21932_ (.Y(_01507_),
    .A(_05390_),
    .B(_05412_));
 sg13g2_a22oi_1 _21933_ (.Y(_01508_),
    .B1(_06409_),
    .B2(_06436_),
    .A2(_01168_),
    .A1(_05769_));
 sg13g2_inv_1 _21934_ (.Y(_01509_),
    .A(_08086_));
 sg13g2_a22oi_1 _21935_ (.Y(_01510_),
    .B1(_01301_),
    .B2(_01306_),
    .A2(_01509_),
    .A1(_05758_));
 sg13g2_nand2_1 _21936_ (.Y(_01511_),
    .A(_01508_),
    .B(_01510_));
 sg13g2_inv_1 _21937_ (.Y(_01512_),
    .A(_01511_));
 sg13g2_inv_1 _21938_ (.Y(_01513_),
    .A(_06454_));
 sg13g2_nand4_1 _21939_ (.B(_01513_),
    .C(_01376_),
    .A(_05772_),
    .Y(_01515_),
    .D(_06124_));
 sg13g2_nor4_1 _21940_ (.A(_07983_),
    .B(_06470_),
    .C(_08360_),
    .D(_01515_),
    .Y(_01516_));
 sg13g2_nand4_1 _21941_ (.B(_01499_),
    .C(_01495_),
    .A(_01512_),
    .Y(_01517_),
    .D(_01516_));
 sg13g2_inv_1 _21942_ (.Y(_01518_),
    .A(_08346_));
 sg13g2_inv_1 _21943_ (.Y(_01519_),
    .A(_07975_));
 sg13g2_nand2_1 _21944_ (.Y(_01520_),
    .A(_01519_),
    .B(_06314_));
 sg13g2_nand2_1 _21945_ (.Y(_01521_),
    .A(_06437_),
    .B(_06409_));
 sg13g2_o21ai_1 _21946_ (.B1(_01521_),
    .Y(_01522_),
    .A1(_01306_),
    .A2(_01302_));
 sg13g2_inv_1 _21947_ (.Y(_01523_),
    .A(_05758_));
 sg13g2_a22oi_1 _21948_ (.Y(_01524_),
    .B1(_05770_),
    .B2(_01168_),
    .A2(_01509_),
    .A1(_01523_));
 sg13g2_nor3_1 _21949_ (.A(_06250_),
    .B(_05945_),
    .C(_01334_),
    .Y(_01525_));
 sg13g2_nand4_1 _21950_ (.B(_01524_),
    .C(_01491_),
    .A(_01502_),
    .Y(_01526_),
    .D(_01525_));
 sg13g2_nor4_1 _21951_ (.A(_01518_),
    .B(_01520_),
    .C(_01522_),
    .D(_01526_),
    .Y(_01527_));
 sg13g2_nor2b_1 _21952_ (.A(_01517_),
    .B_N(_01527_),
    .Y(_01528_));
 sg13g2_nand2_1 _21953_ (.Y(_01529_),
    .A(_05409_),
    .B(net113));
 sg13g2_nor2_1 _21954_ (.A(_05398_),
    .B(_01527_),
    .Y(_01530_));
 sg13g2_nand3_1 _21955_ (.B(net162),
    .C(_01517_),
    .A(_01530_),
    .Y(_01531_));
 sg13g2_buf_1 _21956_ (.A(_01531_),
    .X(_01532_));
 sg13g2_o21ai_1 _21957_ (.B1(_01532_),
    .Y(_01533_),
    .A1(_01528_),
    .A2(_01529_));
 sg13g2_a22oi_1 _21958_ (.Y(_01534_),
    .B1(_01507_),
    .B2(_01533_),
    .A2(_01506_),
    .A1(_01486_));
 sg13g2_nand2b_1 _21959_ (.Y(_01536_),
    .B(_01524_),
    .A_N(_01522_));
 sg13g2_o21ai_1 _21960_ (.B1(_05398_),
    .Y(_01537_),
    .A1(_01511_),
    .A2(_01536_));
 sg13g2_inv_1 _21961_ (.Y(_01538_),
    .A(_01504_));
 sg13g2_a21o_1 _21962_ (.A2(_01538_),
    .A1(_01537_),
    .B1(_05413_),
    .X(_01539_));
 sg13g2_o21ai_1 _21963_ (.B1(_01539_),
    .Y(_01540_),
    .A1(_06411_),
    .A2(_01537_));
 sg13g2_nand2_1 _21964_ (.Y(_01541_),
    .A(_01540_),
    .B(net112));
 sg13g2_nand2_1 _21965_ (.Y(_01542_),
    .A(_01534_),
    .B(_01541_));
 sg13g2_buf_1 _21966_ (.A(\b.gen_square[42].sq.mask ),
    .X(_01543_));
 sg13g2_nand2_1 _21967_ (.Y(_01544_),
    .A(_01542_),
    .B(_01543_));
 sg13g2_nand2_1 _21968_ (.Y(_01545_),
    .A(_01466_),
    .B(_01457_));
 sg13g2_nand3_1 _21969_ (.B(_05401_),
    .C(_01505_),
    .A(_01539_),
    .Y(_01547_));
 sg13g2_inv_1 _21970_ (.Y(_01548_),
    .A(_05402_));
 sg13g2_inv_1 _21971_ (.Y(_01549_),
    .A(_01525_));
 sg13g2_nor3_1 _21972_ (.A(_05401_),
    .B(_01549_),
    .C(_01520_),
    .Y(_01550_));
 sg13g2_nand3_1 _21973_ (.B(_01516_),
    .C(_08346_),
    .A(_01550_),
    .Y(_01551_));
 sg13g2_nand4_1 _21974_ (.B(net95),
    .C(_01548_),
    .A(_01547_),
    .Y(_01552_),
    .D(_01551_));
 sg13g2_a21oi_1 _21975_ (.A1(_05409_),
    .A2(_05399_),
    .Y(_01553_),
    .B1(_05395_));
 sg13g2_nor3_1 _21976_ (.A(net158),
    .B(_01553_),
    .C(_01528_),
    .Y(_01554_));
 sg13g2_nor2_1 _21977_ (.A(_05393_),
    .B(_01532_),
    .Y(_01555_));
 sg13g2_nor2_1 _21978_ (.A(_01554_),
    .B(_01555_),
    .Y(_01556_));
 sg13g2_inv_1 _21979_ (.Y(_01558_),
    .A(_01543_));
 sg13g2_a21oi_1 _21980_ (.A1(_01552_),
    .A2(_01556_),
    .Y(_01559_),
    .B1(_01558_));
 sg13g2_nor2_1 _21981_ (.A(_05412_),
    .B(_06410_),
    .Y(_01560_));
 sg13g2_o21ai_1 _21982_ (.B1(_01560_),
    .Y(_01561_),
    .A1(_05394_),
    .A2(_01532_));
 sg13g2_nand2_1 _21983_ (.Y(_01562_),
    .A(_01561_),
    .B(_01533_));
 sg13g2_nand2_1 _21984_ (.Y(_01563_),
    .A(_01562_),
    .B(_01541_));
 sg13g2_nand2_1 _21985_ (.Y(_01564_),
    .A(_01563_),
    .B(_01543_));
 sg13g2_inv_1 _21986_ (.Y(_01565_),
    .A(_01564_));
 sg13g2_nor2_1 _21987_ (.A(_01447_),
    .B(_01483_),
    .Y(_01566_));
 sg13g2_a21o_1 _21988_ (.A2(_01483_),
    .A1(_01436_),
    .B1(_01566_),
    .X(_01567_));
 sg13g2_buf_1 _21989_ (.A(_01567_),
    .X(_01569_));
 sg13g2_a22oi_1 _21990_ (.Y(_01570_),
    .B1(_01565_),
    .B2(_01569_),
    .A2(_01485_),
    .A1(_01559_));
 sg13g2_inv_1 _21991_ (.Y(_01571_),
    .A(_01569_));
 sg13g2_a22oi_1 _21992_ (.Y(_01572_),
    .B1(_01564_),
    .B2(_01571_),
    .A2(_01545_),
    .A1(_01544_));
 sg13g2_nand2b_1 _21993_ (.Y(_01573_),
    .B(_01572_),
    .A_N(_01570_));
 sg13g2_o21ai_1 _21994_ (.B1(_01573_),
    .Y(_01574_),
    .A1(_01544_),
    .A2(_01545_));
 sg13g2_buf_2 _21995_ (.A(_01574_),
    .X(_01575_));
 sg13g2_nand2_1 _21996_ (.Y(_01576_),
    .A(_01575_),
    .B(_01559_));
 sg13g2_o21ai_1 _21997_ (.B1(_01576_),
    .Y(_01577_),
    .A1(_01485_),
    .A2(_01575_));
 sg13g2_inv_1 _21998_ (.Y(_01578_),
    .A(_06605_));
 sg13g2_a22oi_1 _21999_ (.Y(_01579_),
    .B1(_01578_),
    .B2(_06817_),
    .A2(_01170_),
    .A1(_01196_));
 sg13g2_nor2_1 _22000_ (.A(_01300_),
    .B(_01305_),
    .Y(_01580_));
 sg13g2_a21oi_1 _22001_ (.A1(_08432_),
    .A2(_08435_),
    .Y(_01581_),
    .B1(_01580_));
 sg13g2_and2_1 _22002_ (.A(_01579_),
    .B(_01581_),
    .X(_01582_));
 sg13g2_nor2b_1 _22003_ (.A(_01300_),
    .B_N(_01305_),
    .Y(_01583_));
 sg13g2_nor2_1 _22004_ (.A(_01196_),
    .B(_01171_),
    .Y(_01584_));
 sg13g2_nor2_1 _22005_ (.A(_08436_),
    .B(_08432_),
    .Y(_01585_));
 sg13g2_nor2_1 _22006_ (.A(_06605_),
    .B(_06817_),
    .Y(_01586_));
 sg13g2_nor4_1 _22007_ (.A(_01583_),
    .B(_01584_),
    .C(_01585_),
    .D(_01586_),
    .Y(_01587_));
 sg13g2_a21o_1 _22008_ (.A2(_01587_),
    .A1(_01582_),
    .B1(_06237_),
    .X(_01588_));
 sg13g2_nor2_1 _22009_ (.A(_06893_),
    .B(_06885_),
    .Y(_01590_));
 sg13g2_a221oi_1 _22010_ (.B2(_08021_),
    .C1(_01590_),
    .B1(_08014_),
    .A1(_05544_),
    .Y(_01591_),
    .A2(_07868_));
 sg13g2_nor2_1 _22011_ (.A(_08022_),
    .B(_08014_),
    .Y(_01592_));
 sg13g2_a221oi_1 _22012_ (.B2(_06884_),
    .C1(_01592_),
    .B1(_06893_),
    .A1(_05767_),
    .Y(_01593_),
    .A2(_07868_));
 sg13g2_nand3_1 _22013_ (.B(_01593_),
    .C(_06232_),
    .A(_01591_),
    .Y(_01594_));
 sg13g2_nand2_1 _22014_ (.Y(_01595_),
    .A(_01594_),
    .B(net94));
 sg13g2_a21o_1 _22015_ (.A2(_01595_),
    .A1(_01588_),
    .B1(_06235_),
    .X(_01596_));
 sg13g2_nand3_1 _22016_ (.B(net94),
    .C(_06233_),
    .A(_01594_),
    .Y(_01597_));
 sg13g2_nand3_1 _22017_ (.B(_05177_),
    .C(_01597_),
    .A(_01596_),
    .Y(_01598_));
 sg13g2_nor4_1 _22018_ (.A(_05768_),
    .B(_06830_),
    .C(_08360_),
    .D(_07809_),
    .Y(_01599_));
 sg13g2_nor4_1 _22019_ (.A(_06454_),
    .B(_07017_),
    .C(_05763_),
    .D(_07983_),
    .Y(_01600_));
 sg13g2_nand2_1 _22020_ (.Y(_01601_),
    .A(_01599_),
    .B(_01600_));
 sg13g2_inv_1 _22021_ (.Y(_01602_),
    .A(_01601_));
 sg13g2_nor3_1 _22022_ (.A(_05546_),
    .B(_06250_),
    .C(_06825_),
    .Y(_01603_));
 sg13g2_nand3_1 _22023_ (.B(_08447_),
    .C(_01603_),
    .A(_06796_),
    .Y(_01604_));
 sg13g2_nor3_1 _22024_ (.A(_05177_),
    .B(_07707_),
    .C(_01604_),
    .Y(_01605_));
 sg13g2_nand3_1 _22025_ (.B(_08548_),
    .C(_01605_),
    .A(_01602_),
    .Y(_01606_));
 sg13g2_nor2_1 _22026_ (.A(net83),
    .B(_05178_),
    .Y(_01607_));
 sg13g2_nand3_1 _22027_ (.B(_01606_),
    .C(_01607_),
    .A(_01598_),
    .Y(_01608_));
 sg13g2_nor2_1 _22028_ (.A(_06232_),
    .B(_06193_),
    .Y(_01609_));
 sg13g2_nor2b_1 _22029_ (.A(_01609_),
    .B_N(_01591_),
    .Y(_01611_));
 sg13g2_nor4_1 _22030_ (.A(_05019_),
    .B(_08040_),
    .C(_05016_),
    .D(_05815_),
    .Y(_01612_));
 sg13g2_nor2_1 _22031_ (.A(_08034_),
    .B(_07905_),
    .Y(_01613_));
 sg13g2_nand4_1 _22032_ (.B(_01613_),
    .C(_07923_),
    .A(_01612_),
    .Y(_01614_),
    .D(_05824_));
 sg13g2_inv_1 _22033_ (.Y(_01615_),
    .A(_01614_));
 sg13g2_nand4_1 _22034_ (.B(_01611_),
    .C(_01615_),
    .A(_01602_),
    .Y(_01616_),
    .D(_01582_));
 sg13g2_nand2b_1 _22035_ (.Y(_01617_),
    .B(_06193_),
    .A_N(_06232_));
 sg13g2_nor2b_1 _22036_ (.A(_07930_),
    .B_N(_08116_),
    .Y(_01618_));
 sg13g2_inv_1 _22037_ (.Y(_01619_),
    .A(_01618_));
 sg13g2_nand3_1 _22038_ (.B(_07938_),
    .C(_05832_),
    .A(_11094_),
    .Y(_01620_));
 sg13g2_nor4_1 _22039_ (.A(_01619_),
    .B(_04548_),
    .C(_04567_),
    .D(_01620_),
    .Y(_01622_));
 sg13g2_nand4_1 _22040_ (.B(_00722_),
    .C(_01617_),
    .A(_01593_),
    .Y(_01623_),
    .D(_01622_));
 sg13g2_nor2_1 _22041_ (.A(_01604_),
    .B(_01623_),
    .Y(_01624_));
 sg13g2_and3_1 _22042_ (.X(_01625_),
    .A(_01587_),
    .B(_08548_),
    .C(_01624_));
 sg13g2_nand2b_1 _22043_ (.Y(_01626_),
    .B(_01625_),
    .A_N(_01616_));
 sg13g2_o21ai_1 _22044_ (.B1(_06196_),
    .Y(_01627_),
    .A1(_05170_),
    .A2(net94));
 sg13g2_nand3_1 _22045_ (.B(_05089_),
    .C(_01627_),
    .A(_01626_),
    .Y(_01628_));
 sg13g2_nor2_1 _22046_ (.A(net94),
    .B(_01625_),
    .Y(_01629_));
 sg13g2_nand3_1 _22047_ (.B(net145),
    .C(_01629_),
    .A(_01616_),
    .Y(_01630_));
 sg13g2_nand2b_1 _22048_ (.Y(_01631_),
    .B(_05171_),
    .A_N(_01630_));
 sg13g2_nand3_1 _22049_ (.B(_01628_),
    .C(_01631_),
    .A(_01608_),
    .Y(_01632_));
 sg13g2_buf_1 _22050_ (.A(\b.gen_square[43].sq.mask ),
    .X(_01633_));
 sg13g2_nand2_1 _22051_ (.Y(_01634_),
    .A(_01632_),
    .B(_01633_));
 sg13g2_nand3_1 _22052_ (.B(net86),
    .C(_06237_),
    .A(_01626_),
    .Y(_01635_));
 sg13g2_nand2_1 _22053_ (.Y(_01636_),
    .A(_01635_),
    .B(_01630_));
 sg13g2_nand2_1 _22054_ (.Y(_01637_),
    .A(_01630_),
    .B(_06195_));
 sg13g2_nand2b_1 _22055_ (.Y(_01638_),
    .B(_06194_),
    .A_N(_06234_));
 sg13g2_nand3_1 _22056_ (.B(_01637_),
    .C(_01638_),
    .A(_01636_),
    .Y(_01639_));
 sg13g2_o21ai_1 _22057_ (.B1(_01596_),
    .Y(_01640_),
    .A1(_06607_),
    .A2(_01588_));
 sg13g2_nand2_1 _22058_ (.Y(_01641_),
    .A(_01640_),
    .B(net85));
 sg13g2_nand2_1 _22059_ (.Y(_01643_),
    .A(_01639_),
    .B(_01641_));
 sg13g2_nand2_1 _22060_ (.Y(_01644_),
    .A(_01643_),
    .B(_01633_));
 sg13g2_nor2_1 _22061_ (.A(_01569_),
    .B(_01575_),
    .Y(_01645_));
 sg13g2_a21oi_1 _22062_ (.A1(_01565_),
    .A2(_01575_),
    .Y(_01646_),
    .B1(_01645_));
 sg13g2_inv_2 _22063_ (.Y(_01647_),
    .A(_01646_));
 sg13g2_a22oi_1 _22064_ (.Y(_01648_),
    .B1(_01644_),
    .B2(_01647_),
    .A2(_01634_),
    .A1(_01577_));
 sg13g2_nor2_1 _22065_ (.A(net83),
    .B(_05176_),
    .Y(_01649_));
 sg13g2_a21o_1 _22066_ (.A2(_01622_),
    .A1(_01615_),
    .B1(_05173_),
    .X(_01650_));
 sg13g2_nand2_1 _22067_ (.Y(_01651_),
    .A(_01597_),
    .B(_01650_));
 sg13g2_xnor2_1 _22068_ (.Y(_01652_),
    .A(_05168_),
    .B(_06234_));
 sg13g2_a22oi_1 _22069_ (.Y(_01654_),
    .B1(_01652_),
    .B2(_01636_),
    .A2(_01651_),
    .A1(_01649_));
 sg13g2_nand2_1 _22070_ (.Y(_01655_),
    .A(_01654_),
    .B(_01641_));
 sg13g2_nand2_1 _22071_ (.Y(_01656_),
    .A(_01655_),
    .B(_01633_));
 sg13g2_inv_1 _22072_ (.Y(_01657_),
    .A(_01544_));
 sg13g2_nor2_1 _22073_ (.A(_01657_),
    .B(_01545_),
    .Y(_01658_));
 sg13g2_xnor2_1 _22074_ (.Y(_01659_),
    .A(_01656_),
    .B(_01658_));
 sg13g2_nor2_1 _22075_ (.A(_01644_),
    .B(_01647_),
    .Y(_01660_));
 sg13g2_inv_1 _22076_ (.Y(_01661_),
    .A(_01660_));
 sg13g2_nor2_1 _22077_ (.A(_01634_),
    .B(_01577_),
    .Y(_01662_));
 sg13g2_nand4_1 _22078_ (.B(_01659_),
    .C(_01661_),
    .A(_01648_),
    .Y(_01663_),
    .D(_01662_));
 sg13g2_nor3_1 _22079_ (.A(_01656_),
    .B(_01657_),
    .C(_01545_),
    .Y(_01665_));
 sg13g2_a21oi_1 _22080_ (.A1(_01660_),
    .A2(_01659_),
    .Y(_01666_),
    .B1(_01665_));
 sg13g2_nand2_1 _22081_ (.Y(_01667_),
    .A(_01663_),
    .B(_01666_));
 sg13g2_buf_2 _22082_ (.A(_01667_),
    .X(_01668_));
 sg13g2_nand2_1 _22083_ (.Y(_01669_),
    .A(_01668_),
    .B(_01634_));
 sg13g2_o21ai_1 _22084_ (.B1(_01669_),
    .Y(_01670_),
    .A1(_01577_),
    .A2(_01668_));
 sg13g2_inv_1 _22085_ (.Y(_01671_),
    .A(_01304_));
 sg13g2_a22oi_1 _22086_ (.Y(_01672_),
    .B1(_01172_),
    .B2(_01200_),
    .A2(_01299_),
    .A1(_01671_));
 sg13g2_o21ai_1 _22087_ (.B1(_01672_),
    .Y(_01673_),
    .A1(_06986_),
    .A2(_07009_));
 sg13g2_nor2_1 _22088_ (.A(_06313_),
    .B(_07707_),
    .Y(_01674_));
 sg13g2_inv_1 _22089_ (.Y(_01676_),
    .A(_01674_));
 sg13g2_nand2_1 _22090_ (.Y(_01677_),
    .A(_08393_),
    .B(_08394_));
 sg13g2_nor2_1 _22091_ (.A(_04990_),
    .B(_01677_),
    .Y(_01678_));
 sg13g2_nor4_1 _22092_ (.A(_06825_),
    .B(_01678_),
    .C(net14),
    .D(_04134_),
    .Y(_01679_));
 sg13g2_nand3_1 _22093_ (.B(_06251_),
    .C(_01519_),
    .A(_01679_),
    .Y(_01680_));
 sg13g2_nor2_1 _22094_ (.A(_07950_),
    .B(_06823_),
    .Y(_01681_));
 sg13g2_inv_1 _22095_ (.Y(_01682_),
    .A(_05066_));
 sg13g2_nand2_1 _22096_ (.Y(_01683_),
    .A(_06452_),
    .B(_07695_));
 sg13g2_o21ai_1 _22097_ (.B1(_01683_),
    .Y(_01684_),
    .A1(_01682_),
    .A2(_08390_));
 sg13g2_a221oi_1 _22098_ (.B2(_07206_),
    .C1(_01684_),
    .B1(_07186_),
    .A1(_06708_),
    .Y(_01685_),
    .A2(_06733_));
 sg13g2_inv_1 _22099_ (.Y(_01687_),
    .A(_07737_));
 sg13g2_o21ai_1 _22100_ (.B1(_01687_),
    .Y(_01688_),
    .A1(_04652_),
    .A2(_08256_));
 sg13g2_nor2_1 _22101_ (.A(_07246_),
    .B(_05146_),
    .Y(_01689_));
 sg13g2_nand3_1 _22102_ (.B(_07759_),
    .C(_09006_),
    .A(_01689_),
    .Y(_01690_));
 sg13g2_nor4_1 _22103_ (.A(_01688_),
    .B(_05201_),
    .C(_06635_),
    .D(_01690_),
    .Y(_01691_));
 sg13g2_nand3b_1 _22104_ (.B(_01685_),
    .C(_01691_),
    .Y(_01692_),
    .A_N(_01681_));
 sg13g2_nor4_1 _22105_ (.A(_01673_),
    .B(_01676_),
    .C(_01680_),
    .D(_01692_),
    .Y(_01693_));
 sg13g2_a22oi_1 _22106_ (.Y(_01694_),
    .B1(_07206_),
    .B2(_07185_),
    .A2(_07695_),
    .A1(_06248_));
 sg13g2_inv_1 _22107_ (.Y(_01695_),
    .A(_08390_));
 sg13g2_a22oi_1 _22108_ (.Y(_01696_),
    .B1(_06708_),
    .B2(_06732_),
    .A2(_01695_),
    .A1(_01677_));
 sg13g2_and2_1 _22109_ (.A(_01694_),
    .B(_01696_),
    .X(_01697_));
 sg13g2_inv_1 _22110_ (.Y(_01698_),
    .A(_01697_));
 sg13g2_nor2_1 _22111_ (.A(_07950_),
    .B(_06828_),
    .Y(_01699_));
 sg13g2_a221oi_1 _22112_ (.B2(_01172_),
    .C1(_01699_),
    .B1(_01199_),
    .A1(_01304_),
    .Y(_01700_),
    .A2(_01299_));
 sg13g2_o21ai_1 _22113_ (.B1(_01700_),
    .Y(_01701_),
    .A1(_06986_),
    .A2(_07010_));
 sg13g2_nor2_1 _22114_ (.A(_07831_),
    .B(_08268_),
    .Y(_01702_));
 sg13g2_nand4_1 _22115_ (.B(_07621_),
    .C(_01702_),
    .A(_01493_),
    .Y(_01703_),
    .D(_11345_));
 sg13g2_nor4_1 _22116_ (.A(_06830_),
    .B(_06470_),
    .C(_05054_),
    .D(_07809_),
    .Y(_01704_));
 sg13g2_nand4_1 _22117_ (.B(_01513_),
    .C(_11754_),
    .A(_01704_),
    .Y(_01705_),
    .D(_01185_));
 sg13g2_nor4_1 _22118_ (.A(_01698_),
    .B(_01701_),
    .C(_01703_),
    .D(_01705_),
    .Y(_01706_));
 sg13g2_nor3_1 _22119_ (.A(_04513_),
    .B(_01693_),
    .C(_01706_),
    .Y(_01707_));
 sg13g2_nand2_1 _22120_ (.Y(_01708_),
    .A(_01707_),
    .B(net130));
 sg13g2_nand2_1 _22121_ (.Y(_01709_),
    .A(_01706_),
    .B(_01693_));
 sg13g2_nand3_1 _22122_ (.B(net76),
    .C(_06713_),
    .A(_01709_),
    .Y(_01710_));
 sg13g2_nand2_1 _22123_ (.Y(_01711_),
    .A(_01708_),
    .B(_01710_));
 sg13g2_xnor2_1 _22124_ (.Y(_01712_),
    .A(_04514_),
    .B(_06709_));
 sg13g2_a21oi_1 _22125_ (.A1(_01685_),
    .A2(_01697_),
    .Y(_01713_),
    .B1(_06713_));
 sg13g2_nand2_1 _22126_ (.Y(_01714_),
    .A(_01713_),
    .B(_06712_));
 sg13g2_nand2b_1 _22127_ (.Y(_01715_),
    .B(_01691_),
    .A_N(_01703_));
 sg13g2_nand2_1 _22128_ (.Y(_01716_),
    .A(_01715_),
    .B(_04519_));
 sg13g2_nand2_1 _22129_ (.Y(_01718_),
    .A(_04521_),
    .B(net75));
 sg13g2_a21oi_1 _22130_ (.A1(_01714_),
    .A2(_01716_),
    .Y(_01719_),
    .B1(_01718_));
 sg13g2_a21oi_1 _22131_ (.A1(_01711_),
    .A2(_01712_),
    .Y(_01720_),
    .B1(_01719_));
 sg13g2_nor3_1 _22132_ (.A(_01673_),
    .B(_01681_),
    .C(_01701_),
    .Y(_01721_));
 sg13g2_nor2_1 _22133_ (.A(_06713_),
    .B(_01721_),
    .Y(_01722_));
 sg13g2_o21ai_1 _22134_ (.B1(_06711_),
    .Y(_01723_),
    .A1(_01713_),
    .A2(_01722_));
 sg13g2_nand2_1 _22135_ (.Y(_01724_),
    .A(_01722_),
    .B(_06987_));
 sg13g2_a21o_1 _22136_ (.A2(_01724_),
    .A1(_01723_),
    .B1(_01718_),
    .X(_01725_));
 sg13g2_inv_1 _22137_ (.Y(_01726_),
    .A(\b.gen_square[44].sq.mask ));
 sg13g2_a21o_1 _22138_ (.A2(_01725_),
    .A1(_01720_),
    .B1(_01726_),
    .X(_01727_));
 sg13g2_buf_1 _22139_ (.A(_01727_),
    .X(_01729_));
 sg13g2_nand2_1 _22140_ (.Y(_01730_),
    .A(_01658_),
    .B(_01656_));
 sg13g2_nand2_1 _22141_ (.Y(_01731_),
    .A(_01708_),
    .B(_06660_));
 sg13g2_nand2_1 _22142_ (.Y(_01732_),
    .A(_06710_),
    .B(_06659_));
 sg13g2_nand3_1 _22143_ (.B(_01731_),
    .C(_01732_),
    .A(_01711_),
    .Y(_01733_));
 sg13g2_a21o_1 _22144_ (.A2(_01725_),
    .A1(_01733_),
    .B1(_01726_),
    .X(_01734_));
 sg13g2_buf_1 _22145_ (.A(_01734_),
    .X(_01735_));
 sg13g2_nor2_1 _22146_ (.A(_01647_),
    .B(_01668_),
    .Y(_01736_));
 sg13g2_a21oi_1 _22147_ (.A1(_01644_),
    .A2(_01668_),
    .Y(_01737_),
    .B1(_01736_));
 sg13g2_nand3_1 _22148_ (.B(_04521_),
    .C(_01714_),
    .A(_01723_),
    .Y(_01738_));
 sg13g2_nor4_1 _22149_ (.A(_04521_),
    .B(_01676_),
    .C(_01680_),
    .D(_01705_),
    .Y(_01739_));
 sg13g2_nor3_1 _22150_ (.A(net72),
    .B(_04522_),
    .C(_01739_),
    .Y(_01740_));
 sg13g2_o21ai_1 _22151_ (.B1(_06716_),
    .Y(_01741_),
    .A1(_04517_),
    .A2(_04513_));
 sg13g2_nand3_1 _22152_ (.B(net76),
    .C(_01741_),
    .A(_01709_),
    .Y(_01742_));
 sg13g2_o21ai_1 _22153_ (.B1(_01742_),
    .Y(_01743_),
    .A1(_04517_),
    .A2(_01708_));
 sg13g2_a21oi_1 _22154_ (.A1(_01738_),
    .A2(_01740_),
    .Y(_01744_),
    .B1(_01743_));
 sg13g2_nor2_1 _22155_ (.A(_01726_),
    .B(_01744_),
    .Y(_01745_));
 sg13g2_nand2_1 _22156_ (.Y(_01746_),
    .A(_01670_),
    .B(_01745_));
 sg13g2_o21ai_1 _22157_ (.B1(_01746_),
    .Y(_01747_),
    .A1(_01735_),
    .A2(_01737_));
 sg13g2_a22oi_1 _22158_ (.Y(_01748_),
    .B1(_01735_),
    .B2(_01737_),
    .A2(_01730_),
    .A1(_01729_));
 sg13g2_nand2_1 _22159_ (.Y(_01749_),
    .A(_01747_),
    .B(_01748_));
 sg13g2_o21ai_1 _22160_ (.B1(_01749_),
    .Y(_01750_),
    .A1(_01729_),
    .A2(_01730_));
 sg13g2_buf_2 _22161_ (.A(_01750_),
    .X(_01751_));
 sg13g2_nand2_1 _22162_ (.Y(_01752_),
    .A(_01751_),
    .B(_01745_));
 sg13g2_o21ai_1 _22163_ (.B1(_01752_),
    .Y(_01753_),
    .A1(_01670_),
    .A2(_01751_));
 sg13g2_nor2_1 _22164_ (.A(_04056_),
    .B(_01276_),
    .Y(_01754_));
 sg13g2_nand2b_1 _22165_ (.Y(_01755_),
    .B(_04941_),
    .A_N(_01287_));
 sg13g2_nand3_1 _22166_ (.B(_04058_),
    .C(_01755_),
    .A(_01288_),
    .Y(_01756_));
 sg13g2_nor2b_1 _22167_ (.A(_01272_),
    .B_N(_01256_),
    .Y(_01757_));
 sg13g2_o21ai_1 _22168_ (.B1(_04059_),
    .Y(_01758_),
    .A1(_04042_),
    .A2(_01757_));
 sg13g2_nand3_1 _22169_ (.B(net67),
    .C(_01758_),
    .A(_01756_),
    .Y(_01760_));
 sg13g2_nor2b_1 _22170_ (.A(_01754_),
    .B_N(_01760_),
    .Y(_01761_));
 sg13g2_o21ai_1 _22171_ (.B1(_04946_),
    .Y(_01762_),
    .A1(_04056_),
    .A2(_04041_));
 sg13g2_nand3_1 _22172_ (.B(net57),
    .C(_01762_),
    .A(_01277_),
    .Y(_01763_));
 sg13g2_a21oi_1 _22173_ (.A1(_01761_),
    .A2(_01763_),
    .Y(_01764_),
    .B1(_01291_));
 sg13g2_nor2b_1 _22174_ (.A(_01753_),
    .B_N(_01764_),
    .Y(_01765_));
 sg13g2_nor2_1 _22175_ (.A(_01737_),
    .B(_01751_),
    .Y(_01766_));
 sg13g2_a21oi_2 _22176_ (.B1(_01766_),
    .Y(_01767_),
    .A2(_01751_),
    .A1(_01735_));
 sg13g2_nor2_1 _22177_ (.A(_01293_),
    .B(_01767_),
    .Y(_01768_));
 sg13g2_inv_1 _22178_ (.Y(_01769_),
    .A(_01730_));
 sg13g2_nand2_1 _22179_ (.Y(_01771_),
    .A(_01769_),
    .B(_01729_));
 sg13g2_nor2_1 _22180_ (.A(_02111_),
    .B(_04059_),
    .Y(_01772_));
 sg13g2_inv_1 _22181_ (.Y(_01773_),
    .A(_01249_));
 sg13g2_o21ai_1 _22182_ (.B1(_06622_),
    .Y(_01774_),
    .A1(_01261_),
    .A2(_01773_));
 sg13g2_nand2_1 _22183_ (.Y(_01775_),
    .A(_01755_),
    .B(_01774_));
 sg13g2_xnor2_1 _22184_ (.Y(_01776_),
    .A(_04055_),
    .B(_04942_));
 sg13g2_a22oi_1 _22185_ (.Y(_01777_),
    .B1(_01776_),
    .B2(_01279_),
    .A2(_01775_),
    .A1(_01772_));
 sg13g2_a21o_1 _22186_ (.A2(_01290_),
    .A1(_01777_),
    .B1(_01291_),
    .X(_01778_));
 sg13g2_buf_1 _22187_ (.A(_01778_),
    .X(_01779_));
 sg13g2_a22oi_1 _22188_ (.Y(_01780_),
    .B1(_01293_),
    .B2(_01767_),
    .A2(_01779_),
    .A1(_01771_));
 sg13g2_o21ai_1 _22189_ (.B1(_01780_),
    .Y(_01782_),
    .A1(_01765_),
    .A2(_01768_));
 sg13g2_inv_1 _22190_ (.Y(_01783_),
    .A(_01771_));
 sg13g2_nand2b_1 _22191_ (.Y(_01784_),
    .B(_01783_),
    .A_N(_01779_));
 sg13g2_nand2_1 _22192_ (.Y(_01785_),
    .A(_01782_),
    .B(_01784_));
 sg13g2_nor2_1 _22193_ (.A(_01767_),
    .B(_01785_),
    .Y(_01786_));
 sg13g2_a21oi_1 _22194_ (.A1(_01293_),
    .A2(_01785_),
    .Y(_01787_),
    .B1(_01786_));
 sg13g2_inv_2 _22195_ (.Y(_01788_),
    .A(_01787_));
 sg13g2_nand3_1 _22196_ (.B(net57),
    .C(_04325_),
    .A(_01228_),
    .Y(_01789_));
 sg13g2_nand2_1 _22197_ (.Y(_01790_),
    .A(_01789_),
    .B(_01233_));
 sg13g2_nand2_1 _22198_ (.Y(_01791_),
    .A(_01233_),
    .B(_04234_));
 sg13g2_nand2b_1 _22199_ (.Y(_01793_),
    .B(_04233_),
    .A_N(_04328_));
 sg13g2_nand3_1 _22200_ (.B(_01791_),
    .C(_01793_),
    .A(_01790_),
    .Y(_01794_));
 sg13g2_nand2b_1 _22201_ (.Y(_01795_),
    .B(_04327_),
    .A_N(_01182_));
 sg13g2_nand2_1 _22202_ (.Y(_01796_),
    .A(_01183_),
    .B(_01795_));
 sg13g2_nand2_1 _22203_ (.Y(_01797_),
    .A(_01796_),
    .B(net67));
 sg13g2_nand2_1 _22204_ (.Y(_01798_),
    .A(_01794_),
    .B(_01797_));
 sg13g2_nand2_1 _22205_ (.Y(_01799_),
    .A(_01798_),
    .B(_01236_));
 sg13g2_inv_1 _22206_ (.Y(_01800_),
    .A(_01799_));
 sg13g2_mux2_1 _22207_ (.A0(_01753_),
    .A1(_01764_),
    .S(_01785_),
    .X(_01801_));
 sg13g2_nor2_1 _22208_ (.A(_01237_),
    .B(_01801_),
    .Y(_01802_));
 sg13g2_o21ai_1 _22209_ (.B1(_01802_),
    .Y(_01804_),
    .A1(_01788_),
    .A2(_01800_));
 sg13g2_nor2_1 _22210_ (.A(_09007_),
    .B(_01217_),
    .Y(_01805_));
 sg13g2_nor2_1 _22211_ (.A(_06641_),
    .B(_07735_),
    .Y(_01806_));
 sg13g2_nand3_1 _22212_ (.B(_01805_),
    .C(_01806_),
    .A(_01212_),
    .Y(_01807_));
 sg13g2_a21oi_1 _22213_ (.A1(_06902_),
    .A2(_01807_),
    .Y(_01808_),
    .B1(_01161_));
 sg13g2_nor2b_1 _22214_ (.A(_01796_),
    .B_N(_01808_),
    .Y(_01809_));
 sg13g2_xnor2_1 _22215_ (.Y(_01810_),
    .A(_04229_),
    .B(_04328_));
 sg13g2_nand2_1 _22216_ (.Y(_01811_),
    .A(_01790_),
    .B(_01810_));
 sg13g2_o21ai_1 _22217_ (.B1(_01811_),
    .Y(_01812_),
    .A1(net63),
    .A2(_01809_));
 sg13g2_nand2_1 _22218_ (.Y(_01813_),
    .A(_01812_),
    .B(_01236_));
 sg13g2_nand2_1 _22219_ (.Y(_01815_),
    .A(_01783_),
    .B(_01779_));
 sg13g2_nor2_1 _22220_ (.A(_01813_),
    .B(_01815_),
    .Y(_01816_));
 sg13g2_a21oi_1 _22221_ (.A1(_01788_),
    .A2(_01800_),
    .Y(_01817_),
    .B1(_01816_));
 sg13g2_nand2_1 _22222_ (.Y(_01818_),
    .A(_01804_),
    .B(_01817_));
 sg13g2_nand2_1 _22223_ (.Y(_01819_),
    .A(_01815_),
    .B(_01813_));
 sg13g2_nand2_1 _22224_ (.Y(_01820_),
    .A(_01818_),
    .B(_01819_));
 sg13g2_buf_2 _22225_ (.A(_01820_),
    .X(_01821_));
 sg13g2_nand2_1 _22226_ (.Y(_01822_),
    .A(_01821_),
    .B(_01801_));
 sg13g2_o21ai_1 _22227_ (.B1(_01822_),
    .Y(_01823_),
    .A1(_01237_),
    .A2(_01821_));
 sg13g2_nor2_1 _22228_ (.A(_01800_),
    .B(_01821_),
    .Y(_01824_));
 sg13g2_a21oi_1 _22229_ (.A1(_01788_),
    .A2(_01821_),
    .Y(_01826_),
    .B1(_01824_));
 sg13g2_inv_1 _22230_ (.Y(_01827_),
    .A(_07543_));
 sg13g2_a21oi_1 _22231_ (.A1(_01176_),
    .A2(net82),
    .Y(_01828_),
    .B1(_04333_));
 sg13g2_a21oi_1 _22232_ (.A1(_01204_),
    .A2(net82),
    .Y(_01829_),
    .B1(_04251_));
 sg13g2_inv_1 _22233_ (.Y(_01830_),
    .A(_01829_));
 sg13g2_a22oi_1 _22234_ (.Y(_01831_),
    .B1(_01828_),
    .B2(_01830_),
    .A2(_01827_),
    .A1(_07502_));
 sg13g2_nor2_1 _22235_ (.A(_04435_),
    .B(_07568_),
    .Y(_01832_));
 sg13g2_nor4_1 _22236_ (.A(_04988_),
    .B(_07720_),
    .C(_01832_),
    .D(_01029_),
    .Y(_01833_));
 sg13g2_a21oi_1 _22237_ (.A1(_04382_),
    .A2(net84),
    .Y(_01834_),
    .B1(_07879_));
 sg13g2_inv_1 _22238_ (.Y(_01835_),
    .A(_07875_));
 sg13g2_a21oi_1 _22239_ (.A1(_04478_),
    .A2(net84),
    .Y(_01837_),
    .B1(_01835_));
 sg13g2_inv_1 _22240_ (.Y(_01838_),
    .A(net34));
 sg13g2_inv_1 _22241_ (.Y(_01839_),
    .A(_04120_));
 sg13g2_o21ai_1 _22242_ (.B1(_01839_),
    .Y(_01840_),
    .A1(_01838_),
    .A2(_08692_));
 sg13g2_a21oi_1 _22243_ (.A1(_08687_),
    .A2(_04117_),
    .Y(_01841_),
    .B1(_06868_));
 sg13g2_nor2_1 _22244_ (.A(_07568_),
    .B(_08831_),
    .Y(_01842_));
 sg13g2_nor3_1 _22245_ (.A(_07930_),
    .B(_07934_),
    .C(_07032_),
    .Y(_01843_));
 sg13g2_nand3b_1 _22246_ (.B(_01843_),
    .C(_01254_),
    .Y(_01844_),
    .A_N(_01842_));
 sg13g2_a221oi_1 _22247_ (.B2(_01841_),
    .C1(_01844_),
    .B1(_01840_),
    .A1(_01834_),
    .Y(_01845_),
    .A2(_01837_));
 sg13g2_and3_1 _22248_ (.X(_01846_),
    .A(_01831_),
    .B(_01833_),
    .C(_01845_));
 sg13g2_inv_1 _22249_ (.Y(_01848_),
    .A(_01841_));
 sg13g2_nor2_1 _22250_ (.A(_01848_),
    .B(_01840_),
    .Y(_01849_));
 sg13g2_nor2_1 _22251_ (.A(_07149_),
    .B(_01834_),
    .Y(_01850_));
 sg13g2_inv_1 _22252_ (.Y(_01851_),
    .A(_04435_));
 sg13g2_inv_1 _22253_ (.Y(_01852_),
    .A(_08698_));
 sg13g2_a22oi_1 _22254_ (.Y(_01853_),
    .B1(_01852_),
    .B2(_10011_),
    .A2(_07568_),
    .A1(_01851_));
 sg13g2_nand3b_1 _22255_ (.B(_01853_),
    .C(_07813_),
    .Y(_01854_),
    .A_N(_01850_));
 sg13g2_inv_1 _22256_ (.Y(_01855_),
    .A(_01837_));
 sg13g2_nor4_1 _22257_ (.A(_07905_),
    .B(_07896_),
    .C(_06900_),
    .D(_05019_),
    .Y(_01856_));
 sg13g2_o21ai_1 _22258_ (.B1(_01856_),
    .Y(_01857_),
    .A1(_01834_),
    .A2(_01855_));
 sg13g2_nand2_1 _22259_ (.Y(_01859_),
    .A(_01829_),
    .B(_01828_));
 sg13g2_a22oi_1 _22260_ (.Y(_01860_),
    .B1(_07501_),
    .B2(_01827_),
    .A2(_08830_),
    .A1(_07568_));
 sg13g2_and2_1 _22261_ (.A(_01859_),
    .B(_01860_),
    .X(_01861_));
 sg13g2_inv_1 _22262_ (.Y(_01862_),
    .A(_01861_));
 sg13g2_nor4_1 _22263_ (.A(_01849_),
    .B(_01854_),
    .C(_01857_),
    .D(_01862_),
    .Y(_01863_));
 sg13g2_nor3_1 _22264_ (.A(_04391_),
    .B(_01846_),
    .C(_01863_),
    .Y(_01864_));
 sg13g2_nand2_1 _22265_ (.Y(_01865_),
    .A(_01864_),
    .B(_05079_));
 sg13g2_nand2_1 _22266_ (.Y(_01866_),
    .A(_01863_),
    .B(_01846_));
 sg13g2_nand3_1 _22267_ (.B(net57),
    .C(_04392_),
    .A(_01866_),
    .Y(_01867_));
 sg13g2_nand2_1 _22268_ (.Y(_01868_),
    .A(_01865_),
    .B(_01867_));
 sg13g2_nand2_1 _22269_ (.Y(_01870_),
    .A(_01865_),
    .B(_04403_));
 sg13g2_nand2_1 _22270_ (.Y(_01871_),
    .A(_04482_),
    .B(_04402_));
 sg13g2_nand3_1 _22271_ (.B(_01870_),
    .C(_01871_),
    .A(_01868_),
    .Y(_01872_));
 sg13g2_inv_1 _22272_ (.Y(_01873_),
    .A(_07544_));
 sg13g2_nand2_1 _22273_ (.Y(_01874_),
    .A(_01831_),
    .B(_01861_));
 sg13g2_o21ai_1 _22274_ (.B1(_04391_),
    .Y(_01875_),
    .A1(_01842_),
    .A2(_01874_));
 sg13g2_a21oi_1 _22275_ (.A1(_01848_),
    .A2(_01855_),
    .Y(_01876_),
    .B1(_04392_));
 sg13g2_nand2b_1 _22276_ (.Y(_01877_),
    .B(_01875_),
    .A_N(_01876_));
 sg13g2_nand2_1 _22277_ (.Y(_01878_),
    .A(_01877_),
    .B(_04483_));
 sg13g2_o21ai_1 _22278_ (.B1(_01878_),
    .Y(_01879_),
    .A1(_01873_),
    .A2(_01875_));
 sg13g2_nand2_1 _22279_ (.Y(_01881_),
    .A(_01879_),
    .B(net56));
 sg13g2_inv_1 _22280_ (.Y(_01882_),
    .A(\b.gen_square[47].sq.mask ));
 sg13g2_a21o_1 _22281_ (.A2(_01881_),
    .A1(_01872_),
    .B1(_01882_),
    .X(_01883_));
 sg13g2_buf_1 _22282_ (.A(_01883_),
    .X(_01884_));
 sg13g2_o21ai_1 _22283_ (.B1(_04404_),
    .Y(_01885_),
    .A1(_04387_),
    .A2(_04391_));
 sg13g2_nand3_1 _22284_ (.B(net41),
    .C(_01885_),
    .A(_01866_),
    .Y(_01886_));
 sg13g2_o21ai_1 _22285_ (.B1(_01886_),
    .Y(_01887_),
    .A1(_04387_),
    .A2(_01865_));
 sg13g2_nand2_1 _22286_ (.Y(_01888_),
    .A(_01876_),
    .B(_04484_));
 sg13g2_nand3_1 _22287_ (.B(_04394_),
    .C(_01888_),
    .A(_01878_),
    .Y(_01889_));
 sg13g2_nor2_1 _22288_ (.A(_01252_),
    .B(_01854_),
    .Y(_01890_));
 sg13g2_nand3_1 _22289_ (.B(_04389_),
    .C(_01833_),
    .A(_01890_),
    .Y(_01892_));
 sg13g2_nor2_1 _22290_ (.A(_02122_),
    .B(_04395_),
    .Y(_01893_));
 sg13g2_and3_1 _22291_ (.X(_01894_),
    .A(_01889_),
    .B(_01892_),
    .C(_01893_));
 sg13g2_o21ai_1 _22292_ (.B1(\b.gen_square[47].sq.mask ),
    .Y(_01895_),
    .A1(_01887_),
    .A2(_01894_));
 sg13g2_a22oi_1 _22293_ (.Y(_01896_),
    .B1(_01823_),
    .B2(_01895_),
    .A2(_01884_),
    .A1(_01826_));
 sg13g2_a21oi_1 _22294_ (.A1(_01843_),
    .A2(_01856_),
    .Y(_01897_),
    .B1(_07167_));
 sg13g2_nand2b_1 _22295_ (.Y(_01898_),
    .B(_01888_),
    .A_N(_01897_));
 sg13g2_o21ai_1 _22296_ (.B1(_05116_),
    .Y(_01899_),
    .A1(_01898_),
    .A2(_01879_));
 sg13g2_nor2_1 _22297_ (.A(_04385_),
    .B(_04481_),
    .Y(_01900_));
 sg13g2_o21ai_1 _22298_ (.B1(_01868_),
    .Y(_01901_),
    .A1(_04483_),
    .A2(_01900_));
 sg13g2_a21o_1 _22299_ (.A2(_01901_),
    .A1(_01899_),
    .B1(_01882_),
    .X(_01903_));
 sg13g2_buf_1 _22300_ (.A(_01903_),
    .X(_01904_));
 sg13g2_nor2b_1 _22301_ (.A(_01815_),
    .B_N(_01813_),
    .Y(_01905_));
 sg13g2_xnor2_1 _22302_ (.Y(_01906_),
    .A(_01904_),
    .B(_01905_));
 sg13g2_nor2_1 _22303_ (.A(_01884_),
    .B(_01826_),
    .Y(_01907_));
 sg13g2_inv_1 _22304_ (.Y(_01908_),
    .A(_01907_));
 sg13g2_nor2_1 _22305_ (.A(_01895_),
    .B(_01823_),
    .Y(_01909_));
 sg13g2_nand4_1 _22306_ (.B(_01906_),
    .C(_01908_),
    .A(_01896_),
    .Y(_01910_),
    .D(_01909_));
 sg13g2_nor2b_1 _22307_ (.A(_01904_),
    .B_N(_01905_),
    .Y(_01911_));
 sg13g2_a21oi_1 _22308_ (.A1(_01907_),
    .A2(_01906_),
    .Y(_01912_),
    .B1(_01911_));
 sg13g2_nand2_2 _22309_ (.Y(_01914_),
    .A(_01910_),
    .B(_01912_));
 sg13g2_nand2_1 _22310_ (.Y(_01915_),
    .A(_01914_),
    .B(_01895_));
 sg13g2_o21ai_1 _22311_ (.B1(_01915_),
    .Y(_01916_),
    .A1(_01823_),
    .A2(_01914_));
 sg13g2_nand3_1 _22312_ (.B(_01158_),
    .C(_01916_),
    .A(_01156_),
    .Y(_01917_));
 sg13g2_nand2_1 _22313_ (.Y(_01918_),
    .A(_01905_),
    .B(_01904_));
 sg13g2_nor2_1 _22314_ (.A(_01130_),
    .B(_01131_),
    .Y(_01919_));
 sg13g2_nor2_1 _22315_ (.A(_01918_),
    .B(_01919_),
    .Y(_01920_));
 sg13g2_inv_1 _22316_ (.Y(_01921_),
    .A(_01919_));
 sg13g2_nor2b_1 _22317_ (.A(_01921_),
    .B_N(_01918_),
    .Y(_01922_));
 sg13g2_nor2_1 _22318_ (.A(_01920_),
    .B(_01922_),
    .Y(_01923_));
 sg13g2_nand2_1 _22319_ (.Y(_01925_),
    .A(_01917_),
    .B(_01923_));
 sg13g2_nand2_1 _22320_ (.Y(_01926_),
    .A(_01154_),
    .B(_08900_));
 sg13g2_nand3_1 _22321_ (.B(_01127_),
    .C(_01152_),
    .A(_01148_),
    .Y(_01927_));
 sg13g2_nor2_1 _22322_ (.A(_01826_),
    .B(_01914_),
    .Y(_01928_));
 sg13g2_a21oi_1 _22323_ (.A1(_01884_),
    .A2(_01914_),
    .Y(_01929_),
    .B1(_01928_));
 sg13g2_inv_1 _22324_ (.Y(_01930_),
    .A(_01929_));
 sg13g2_nand3_1 _22325_ (.B(_01927_),
    .C(_01930_),
    .A(_01926_),
    .Y(_01931_));
 sg13g2_inv_1 _22326_ (.Y(_01932_),
    .A(_08900_));
 sg13g2_nand2_1 _22327_ (.Y(_01933_),
    .A(_01154_),
    .B(_01932_));
 sg13g2_nand3_1 _22328_ (.B(_01150_),
    .C(_01152_),
    .A(_01148_),
    .Y(_01934_));
 sg13g2_nand3_1 _22329_ (.B(_01934_),
    .C(_01929_),
    .A(_01933_),
    .Y(_01936_));
 sg13g2_nand2_1 _22330_ (.Y(_01937_),
    .A(_01931_),
    .B(_01936_));
 sg13g2_nor2_1 _22331_ (.A(_01925_),
    .B(_01937_),
    .Y(_01938_));
 sg13g2_a21oi_1 _22332_ (.A1(_01156_),
    .A2(_01158_),
    .Y(_01939_),
    .B1(_01916_));
 sg13g2_nand2_1 _22333_ (.Y(_01940_),
    .A(_01938_),
    .B(_01939_));
 sg13g2_inv_1 _22334_ (.Y(_01941_),
    .A(_01936_));
 sg13g2_a21oi_2 _22335_ (.B1(_01922_),
    .Y(_01942_),
    .A2(_01923_),
    .A1(_01941_));
 sg13g2_nand2_1 _22336_ (.Y(_01943_),
    .A(_01940_),
    .B(_01942_));
 sg13g2_buf_1 _22337_ (.A(_01943_),
    .X(_01944_));
 sg13g2_nand2_1 _22338_ (.Y(_01945_),
    .A(net13),
    .B(_01930_));
 sg13g2_nand2_1 _22339_ (.Y(_01947_),
    .A(_01926_),
    .B(_01927_));
 sg13g2_nand3_1 _22340_ (.B(_01947_),
    .C(_01942_),
    .A(_01940_),
    .Y(_01948_));
 sg13g2_nand2_1 _22341_ (.Y(_01949_),
    .A(_01945_),
    .B(_01948_));
 sg13g2_xnor2_1 _22342_ (.Y(_01950_),
    .A(_07689_),
    .B(_01949_));
 sg13g2_nand2_1 _22343_ (.Y(_01951_),
    .A(_07686_),
    .B(_07668_));
 sg13g2_o21ai_1 _22344_ (.B1(_01951_),
    .Y(_01952_),
    .A1(_07666_),
    .A2(_07686_));
 sg13g2_nand2_1 _22345_ (.Y(_01953_),
    .A(_01156_),
    .B(_01158_));
 sg13g2_nand3_1 _22346_ (.B(_01953_),
    .C(_01942_),
    .A(_01940_),
    .Y(_01954_));
 sg13g2_nand2b_1 _22347_ (.Y(_01955_),
    .B(_01916_),
    .A_N(_01942_));
 sg13g2_nand2_1 _22348_ (.Y(_01956_),
    .A(_01954_),
    .B(_01955_));
 sg13g2_nor2_1 _22349_ (.A(_01952_),
    .B(_01956_),
    .Y(_01958_));
 sg13g2_nor2_1 _22350_ (.A(_07681_),
    .B(_07684_),
    .Y(_01959_));
 sg13g2_inv_1 _22351_ (.Y(_01960_),
    .A(_01959_));
 sg13g2_nor2_1 _22352_ (.A(_01918_),
    .B(_01921_),
    .Y(_01961_));
 sg13g2_nor2_1 _22353_ (.A(_01960_),
    .B(_01961_),
    .Y(_01962_));
 sg13g2_inv_2 _22354_ (.Y(_01963_),
    .A(_01961_));
 sg13g2_nor2_1 _22355_ (.A(_01959_),
    .B(_01963_),
    .Y(_01964_));
 sg13g2_nor2_1 _22356_ (.A(_01962_),
    .B(_01964_),
    .Y(_01965_));
 sg13g2_nor2b_1 _22357_ (.A(_01958_),
    .B_N(_01965_),
    .Y(_01966_));
 sg13g2_nand2_1 _22358_ (.Y(_01967_),
    .A(_01950_),
    .B(_01966_));
 sg13g2_nand2_1 _22359_ (.Y(_01969_),
    .A(_01949_),
    .B(_07688_));
 sg13g2_inv_1 _22360_ (.Y(_01970_),
    .A(_01964_));
 sg13g2_nand2_1 _22361_ (.Y(_01971_),
    .A(_01969_),
    .B(_01970_));
 sg13g2_nand2b_1 _22362_ (.Y(_01972_),
    .B(_01971_),
    .A_N(_01962_));
 sg13g2_nand2_1 _22363_ (.Y(_01973_),
    .A(_01967_),
    .B(_01972_));
 sg13g2_nand2_1 _22364_ (.Y(_01974_),
    .A(_01956_),
    .B(_01952_));
 sg13g2_nand3_1 _22365_ (.B(_01966_),
    .C(_01974_),
    .A(_01950_),
    .Y(_01975_));
 sg13g2_buf_1 _22366_ (.A(_01975_),
    .X(_01976_));
 sg13g2_nand2_1 _22367_ (.Y(_01977_),
    .A(_01973_),
    .B(_01976_));
 sg13g2_buf_8 _22368_ (.A(_01977_),
    .X(_01978_));
 sg13g2_inv_1 _22369_ (.Y(_01980_),
    .A(_01956_));
 sg13g2_nand2_1 _22370_ (.Y(_01981_),
    .A(_01978_),
    .B(_01980_));
 sg13g2_nand3_1 _22371_ (.B(_01976_),
    .C(_01952_),
    .A(_01973_),
    .Y(_01982_));
 sg13g2_nand2_1 _22372_ (.Y(_01983_),
    .A(_01981_),
    .B(_01982_));
 sg13g2_inv_1 _22373_ (.Y(_01984_),
    .A(_04464_));
 sg13g2_inv_1 _22374_ (.Y(_01985_),
    .A(_05064_));
 sg13g2_a21oi_2 _22375_ (.B1(_01985_),
    .Y(_01986_),
    .A2(_01984_),
    .A1(_07558_));
 sg13g2_inv_1 _22376_ (.Y(_01987_),
    .A(_01986_));
 sg13g2_a221oi_1 _22377_ (.B2(_01851_),
    .C1(_01850_),
    .B1(_04441_),
    .A1(_01987_),
    .Y(_01988_),
    .A2(_07615_));
 sg13g2_nor2_1 _22378_ (.A(_04459_),
    .B(_01987_),
    .Y(_01989_));
 sg13g2_nor3_1 _22379_ (.A(_04442_),
    .B(_01989_),
    .C(_01252_),
    .Y(_01991_));
 sg13g2_a21oi_1 _22380_ (.A1(_01988_),
    .A2(_01991_),
    .Y(_01992_),
    .B1(_04427_));
 sg13g2_a21oi_1 _22381_ (.A1(_05023_),
    .A2(net84),
    .Y(_01993_),
    .B1(_01835_));
 sg13g2_inv_1 _22382_ (.Y(_01994_),
    .A(_01993_));
 sg13g2_nor2_1 _22383_ (.A(_04427_),
    .B(_01994_),
    .Y(_01995_));
 sg13g2_a21oi_1 _22384_ (.A1(_07504_),
    .A2(_08828_),
    .Y(_01996_),
    .B1(_04441_));
 sg13g2_a21oi_1 _22385_ (.A1(_07551_),
    .A2(_08828_),
    .Y(_01997_),
    .B1(_08829_));
 sg13g2_inv_1 _22386_ (.Y(_01998_),
    .A(_05460_));
 sg13g2_nor3_1 _22387_ (.A(_05459_),
    .B(_05477_),
    .C(_05466_),
    .Y(_01999_));
 sg13g2_a21oi_1 _22388_ (.A1(_01998_),
    .A2(_05977_),
    .Y(_02000_),
    .B1(_01999_));
 sg13g2_inv_1 _22389_ (.Y(_02002_),
    .A(_02000_));
 sg13g2_inv_1 _22390_ (.Y(_02003_),
    .A(_05487_));
 sg13g2_nor2_1 _22391_ (.A(_05486_),
    .B(_06279_),
    .Y(_02004_));
 sg13g2_a21oi_1 _22392_ (.A1(_02002_),
    .A2(_02003_),
    .Y(_02005_),
    .B1(_02004_));
 sg13g2_inv_1 _22393_ (.Y(_02006_),
    .A(_02005_));
 sg13g2_nor2_1 _22394_ (.A(_06259_),
    .B(_06783_),
    .Y(_02007_));
 sg13g2_a21oi_1 _22395_ (.A1(_02006_),
    .A2(_06262_),
    .Y(_02008_),
    .B1(_02007_));
 sg13g2_inv_1 _22396_ (.Y(_02009_),
    .A(_02008_));
 sg13g2_nor2_1 _22397_ (.A(_04992_),
    .B(_06911_),
    .Y(_02010_));
 sg13g2_a21oi_1 _22398_ (.A1(_02009_),
    .A2(_04995_),
    .Y(_02011_),
    .B1(_02010_));
 sg13g2_inv_1 _22399_ (.Y(_02013_),
    .A(_02011_));
 sg13g2_nor2_1 _22400_ (.A(_04378_),
    .B(_07156_),
    .Y(_02014_));
 sg13g2_a21oi_1 _22401_ (.A1(_02013_),
    .A2(_04380_),
    .Y(_02015_),
    .B1(_02014_));
 sg13g2_inv_1 _22402_ (.Y(_02016_),
    .A(_02015_));
 sg13g2_nor2_1 _22403_ (.A(_04462_),
    .B(_04495_),
    .Y(_02017_));
 sg13g2_a21oi_1 _22404_ (.A1(_02016_),
    .A2(_01984_),
    .Y(_02018_),
    .B1(_02017_));
 sg13g2_inv_1 _22405_ (.Y(_02019_),
    .A(_02018_));
 sg13g2_a21oi_1 _22406_ (.A1(_05444_),
    .A2(_01998_),
    .Y(_02020_),
    .B1(_05464_));
 sg13g2_inv_1 _22407_ (.Y(_02021_),
    .A(_02020_));
 sg13g2_a21oi_1 _22408_ (.A1(_02021_),
    .A2(_02003_),
    .Y(_02022_),
    .B1(_05491_));
 sg13g2_nor2_1 _22409_ (.A(_05185_),
    .B(_06262_),
    .Y(_02024_));
 sg13g2_a21oi_1 _22410_ (.A1(_02022_),
    .A2(_06262_),
    .Y(_02025_),
    .B1(_02024_));
 sg13g2_inv_1 _22411_ (.Y(_02026_),
    .A(_02025_));
 sg13g2_nor2_1 _22412_ (.A(_04549_),
    .B(_04995_),
    .Y(_02027_));
 sg13g2_a21oi_1 _22413_ (.A1(_02026_),
    .A2(_04995_),
    .Y(_02028_),
    .B1(_02027_));
 sg13g2_inv_1 _22414_ (.Y(_02029_),
    .A(_02028_));
 sg13g2_nor2_1 _22415_ (.A(_06630_),
    .B(_04380_),
    .Y(_02030_));
 sg13g2_a21oi_1 _22416_ (.A1(_02029_),
    .A2(_04380_),
    .Y(_02031_),
    .B1(_02030_));
 sg13g2_inv_1 _22417_ (.Y(_02032_),
    .A(_02031_));
 sg13g2_o21ai_1 _22418_ (.B1(_05064_),
    .Y(_02033_),
    .A1(_04464_),
    .A2(_02032_));
 sg13g2_nor2_1 _22419_ (.A(_02019_),
    .B(_02033_),
    .Y(_02035_));
 sg13g2_a21oi_1 _22420_ (.A1(_01996_),
    .A2(_01997_),
    .Y(_02036_),
    .B1(_02035_));
 sg13g2_inv_1 _22421_ (.Y(_02037_),
    .A(_01996_));
 sg13g2_a22oi_1 _22422_ (.Y(_02038_),
    .B1(_02033_),
    .B2(_02018_),
    .A2(_01997_),
    .A1(_02037_));
 sg13g2_a21oi_1 _22423_ (.A1(_02036_),
    .A2(_02038_),
    .Y(_02039_),
    .B1(_04427_));
 sg13g2_o21ai_1 _22424_ (.B1(_04501_),
    .Y(_02040_),
    .A1(_01995_),
    .A2(_02039_));
 sg13g2_nand2_1 _22425_ (.Y(_02041_),
    .A(_01995_),
    .B(_04498_));
 sg13g2_nand3_1 _22426_ (.B(_04415_),
    .C(_02041_),
    .A(_02040_),
    .Y(_02042_));
 sg13g2_o21ai_1 _22427_ (.B1(_02042_),
    .Y(_02043_),
    .A1(_04415_),
    .A2(_01992_));
 sg13g2_nor2_1 _22428_ (.A(net48),
    .B(_02043_),
    .Y(_02044_));
 sg13g2_a21oi_1 _22429_ (.A1(_04975_),
    .A2(net84),
    .Y(_02046_),
    .B1(_07879_));
 sg13g2_a21oi_1 _22430_ (.A1(_02046_),
    .A2(_01993_),
    .Y(_02047_),
    .B1(_07932_));
 sg13g2_nand3_1 _22431_ (.B(_02036_),
    .C(_01991_),
    .A(_02047_),
    .Y(_02048_));
 sg13g2_inv_1 _22432_ (.Y(_02049_),
    .A(_02048_));
 sg13g2_inv_1 _22433_ (.Y(_02050_),
    .A(_02046_));
 sg13g2_a21oi_1 _22434_ (.A1(_02050_),
    .A2(_01993_),
    .Y(_02051_),
    .B1(_07907_));
 sg13g2_and3_1 _22435_ (.X(_02052_),
    .A(_02051_),
    .B(_02038_),
    .C(_01988_));
 sg13g2_nor3_1 _22436_ (.A(_04416_),
    .B(_02049_),
    .C(_02052_),
    .Y(_02053_));
 sg13g2_inv_1 _22437_ (.Y(_02054_),
    .A(_04413_));
 sg13g2_nand3_1 _22438_ (.B(net97),
    .C(_02054_),
    .A(_02053_),
    .Y(_02055_));
 sg13g2_nor2b_1 _22439_ (.A(_02044_),
    .B_N(_02055_),
    .Y(_02057_));
 sg13g2_nand2_1 _22440_ (.Y(_02058_),
    .A(_02052_),
    .B(_02049_));
 sg13g2_and3_1 _22441_ (.X(_02059_),
    .A(_02058_),
    .B(net41),
    .C(_07553_));
 sg13g2_o21ai_1 _22442_ (.B1(_02059_),
    .Y(_02060_),
    .A1(_02054_),
    .A2(_04423_));
 sg13g2_buf_1 _22443_ (.A(\b.gen_square[63].sq.mask ),
    .X(_02061_));
 sg13g2_inv_1 _22444_ (.Y(_02062_),
    .A(_02061_));
 sg13g2_a21oi_1 _22445_ (.A1(_02057_),
    .A2(_02060_),
    .Y(_02063_),
    .B1(_02062_));
 sg13g2_buf_1 _22446_ (.A(\b.gen_square[61].sq.mask ),
    .X(_02064_));
 sg13g2_inv_1 _22447_ (.Y(_02065_),
    .A(_02064_));
 sg13g2_a21oi_1 _22448_ (.A1(_07237_),
    .A2(net77),
    .Y(_02066_),
    .B1(_04728_));
 sg13g2_a21oi_1 _22449_ (.A1(_07128_),
    .A2(net77),
    .Y(_02068_),
    .B1(_04796_));
 sg13g2_nand2b_1 _22450_ (.Y(_02069_),
    .B(_02068_),
    .A_N(_02066_));
 sg13g2_inv_1 _22451_ (.Y(_02070_),
    .A(_06894_));
 sg13g2_nor2_1 _22452_ (.A(\b.gen_square[52].sq.color ),
    .B(net23),
    .Y(_02071_));
 sg13g2_a21o_1 _22453_ (.A2(net23),
    .A1(_02070_),
    .B1(_02071_),
    .X(_02072_));
 sg13g2_buf_1 _22454_ (.A(_02072_),
    .X(_02073_));
 sg13g2_inv_1 _22455_ (.Y(_02074_),
    .A(_02073_));
 sg13g2_nor2_1 _22456_ (.A(_06822_),
    .B(_02074_),
    .Y(_02075_));
 sg13g2_nor3_1 _22457_ (.A(_01989_),
    .B(_07241_),
    .C(_02075_),
    .Y(_02076_));
 sg13g2_nor2b_1 _22458_ (.A(_04999_),
    .B_N(_02076_),
    .Y(_02077_));
 sg13g2_a21oi_1 _22459_ (.A1(_01986_),
    .A2(_04380_),
    .Y(_02079_),
    .B1(_02030_));
 sg13g2_inv_1 _22460_ (.Y(_02080_),
    .A(_02079_));
 sg13g2_a21oi_1 _22461_ (.A1(_02080_),
    .A2(_04995_),
    .Y(_02081_),
    .B1(_02027_));
 sg13g2_buf_1 _22462_ (.A(_02081_),
    .X(_02082_));
 sg13g2_inv_1 _22463_ (.Y(_02083_),
    .A(_02082_));
 sg13g2_a21oi_1 _22464_ (.A1(_07039_),
    .A2(net23),
    .Y(_02084_),
    .B1(_08020_));
 sg13g2_nand2_1 _22465_ (.Y(_02085_),
    .A(_02029_),
    .B(_02011_));
 sg13g2_a21oi_1 _22466_ (.A1(_01984_),
    .A2(_07557_),
    .Y(_02086_),
    .B1(_02017_));
 sg13g2_nand2_1 _22467_ (.Y(_02087_),
    .A(_01986_),
    .B(_02086_));
 sg13g2_o21ai_1 _22468_ (.B1(_05049_),
    .Y(_02088_),
    .A1(_05048_),
    .A2(_04407_));
 sg13g2_a21oi_1 _22469_ (.A1(_05003_),
    .A2(net84),
    .Y(_02090_),
    .B1(_01835_));
 sg13g2_nor2_1 _22470_ (.A(_08673_),
    .B(_07926_),
    .Y(_02091_));
 sg13g2_nor2_1 _22471_ (.A(_07029_),
    .B(_04528_),
    .Y(_02092_));
 sg13g2_nand2_1 _22472_ (.Y(_02093_),
    .A(_02091_),
    .B(_02092_));
 sg13g2_a21oi_1 _22473_ (.A1(_02088_),
    .A2(_02090_),
    .Y(_02094_),
    .B1(_02093_));
 sg13g2_nand3_1 _22474_ (.B(_02087_),
    .C(_02094_),
    .A(_02085_),
    .Y(_02095_));
 sg13g2_a221oi_1 _22475_ (.B2(_02084_),
    .C1(_02095_),
    .B1(_02073_),
    .A1(_02083_),
    .Y(_02096_),
    .A2(_06788_));
 sg13g2_nand3_1 _22476_ (.B(_02077_),
    .C(_02096_),
    .A(_02069_),
    .Y(_02097_));
 sg13g2_nand3_1 _22477_ (.B(net97),
    .C(_04362_),
    .A(_02097_),
    .Y(_02098_));
 sg13g2_nor2_1 _22478_ (.A(_02013_),
    .B(_02029_),
    .Y(_02099_));
 sg13g2_nand2_1 _22479_ (.Y(_02101_),
    .A(_02082_),
    .B(_06788_));
 sg13g2_inv_1 _22480_ (.Y(_02102_),
    .A(_05067_));
 sg13g2_inv_1 _22481_ (.Y(_02103_),
    .A(_07150_));
 sg13g2_nand2_1 _22482_ (.Y(_02104_),
    .A(_01987_),
    .B(_07615_));
 sg13g2_and4_1 _22483_ (.A(_02101_),
    .B(_02102_),
    .C(_02103_),
    .D(_02104_),
    .X(_02105_));
 sg13g2_o21ai_1 _22484_ (.B1(_02105_),
    .Y(_02106_),
    .A1(_06822_),
    .A2(_02073_));
 sg13g2_nor2b_1 _22485_ (.A(_02088_),
    .B_N(_02090_),
    .Y(_02107_));
 sg13g2_a21oi_1 _22486_ (.A1(_02074_),
    .A2(_02084_),
    .Y(_02108_),
    .B1(_02107_));
 sg13g2_nand3_1 _22487_ (.B(_00833_),
    .C(_01260_),
    .A(_02108_),
    .Y(_02109_));
 sg13g2_inv_1 _22488_ (.Y(_02110_),
    .A(_02086_));
 sg13g2_nand2_1 _22489_ (.Y(_02112_),
    .A(_02066_),
    .B(_02068_));
 sg13g2_o21ai_1 _22490_ (.B1(_02112_),
    .Y(_02113_),
    .A1(_02110_),
    .A2(_01986_));
 sg13g2_nor4_1 _22491_ (.A(_02099_),
    .B(_02106_),
    .C(_02109_),
    .D(_02113_),
    .Y(_02114_));
 sg13g2_or2_1 _22492_ (.X(_02115_),
    .B(_02114_),
    .A(_02098_));
 sg13g2_buf_1 _22493_ (.A(_02115_),
    .X(_02116_));
 sg13g2_nor2_1 _22494_ (.A(_04366_),
    .B(_02116_),
    .Y(_02117_));
 sg13g2_o21ai_1 _22495_ (.B1(_04368_),
    .Y(_02118_),
    .A1(_06787_),
    .A2(_02082_));
 sg13g2_inv_1 _22496_ (.Y(_02119_),
    .A(_02077_));
 sg13g2_nor3_1 _22497_ (.A(_02106_),
    .B(_02118_),
    .C(_02119_),
    .Y(_02120_));
 sg13g2_o21ai_1 _22498_ (.B1(_04361_),
    .Y(_02121_),
    .A1(_02090_),
    .A2(_02084_));
 sg13g2_o21ai_1 _22499_ (.B1(_04369_),
    .Y(_02123_),
    .A1(_04471_),
    .A2(_02121_));
 sg13g2_nand2_1 _22500_ (.Y(_02124_),
    .A(_02013_),
    .B(_02110_));
 sg13g2_o21ai_1 _22501_ (.B1(_04361_),
    .Y(_02125_),
    .A1(_02124_),
    .A2(_02068_));
 sg13g2_a21oi_1 _22502_ (.A1(_02125_),
    .A2(_02121_),
    .Y(_02126_),
    .B1(_04475_));
 sg13g2_nor2_1 _22503_ (.A(_02123_),
    .B(_02126_),
    .Y(_02127_));
 sg13g2_nor4_1 _22504_ (.A(net48),
    .B(_04372_),
    .C(_02120_),
    .D(_02127_),
    .Y(_02128_));
 sg13g2_nor2_1 _22505_ (.A(_04378_),
    .B(_04362_),
    .Y(_02129_));
 sg13g2_nor2_1 _22506_ (.A(_04367_),
    .B(_04378_),
    .Y(_02130_));
 sg13g2_nor2b_1 _22507_ (.A(_02097_),
    .B_N(_02114_),
    .Y(_02131_));
 sg13g2_nor4_1 _22508_ (.A(net142),
    .B(_02129_),
    .C(_02130_),
    .D(_02131_),
    .Y(_02132_));
 sg13g2_nor3_1 _22509_ (.A(_02117_),
    .B(_02128_),
    .C(_02132_),
    .Y(_02134_));
 sg13g2_nor2_1 _22510_ (.A(_02065_),
    .B(_02134_),
    .Y(_02135_));
 sg13g2_inv_1 _22511_ (.Y(_02136_),
    .A(\b.gen_square[60].sq.mask ));
 sg13g2_inv_1 _22512_ (.Y(_02137_),
    .A(_07232_));
 sg13g2_a21oi_1 _22513_ (.A1(_02137_),
    .A2(net77),
    .Y(_02138_),
    .B1(_08815_));
 sg13g2_a21oi_1 _22514_ (.A1(_06772_),
    .A2(net31),
    .Y(_02139_),
    .B1(_07694_));
 sg13g2_nor2_1 _22515_ (.A(_02138_),
    .B(_02139_),
    .Y(_02140_));
 sg13g2_nor2_1 _22516_ (.A(_06784_),
    .B(_02140_),
    .Y(_02141_));
 sg13g2_a21oi_1 _22517_ (.A1(_02110_),
    .A2(_04380_),
    .Y(_02142_),
    .B1(_02014_));
 sg13g2_inv_1 _22518_ (.Y(_02143_),
    .A(_02142_));
 sg13g2_a21oi_1 _22519_ (.A1(_07022_),
    .A2(net23),
    .Y(_02145_),
    .B1(_04702_));
 sg13g2_inv_1 _22520_ (.Y(_02146_),
    .A(_06991_));
 sg13g2_a21oi_1 _22521_ (.A1(_02146_),
    .A2(net23),
    .Y(_02147_),
    .B1(_04787_));
 sg13g2_nand2_1 _22522_ (.Y(_02148_),
    .A(_02145_),
    .B(_02147_));
 sg13g2_o21ai_1 _22523_ (.B1(_02148_),
    .Y(_02149_),
    .A1(_02143_),
    .A2(_02080_));
 sg13g2_inv_1 _22524_ (.Y(_02150_),
    .A(_02145_));
 sg13g2_a22oi_1 _22525_ (.Y(_02151_),
    .B1(_02147_),
    .B2(_02150_),
    .A2(_02080_),
    .A1(_02142_));
 sg13g2_inv_1 _22526_ (.Y(_02152_),
    .A(_02151_));
 sg13g2_nor3_1 _22527_ (.A(_02149_),
    .B(_02008_),
    .C(_02152_),
    .Y(_02153_));
 sg13g2_nor2_1 _22528_ (.A(_06784_),
    .B(_02153_),
    .Y(_02154_));
 sg13g2_o21ai_1 _22529_ (.B1(_06762_),
    .Y(_02156_),
    .A1(_02141_),
    .A2(_02154_));
 sg13g2_nand2b_1 _22530_ (.Y(_02157_),
    .B(_02141_),
    .A_N(_06764_));
 sg13g2_nand3_1 _22531_ (.B(_04562_),
    .C(_02157_),
    .A(_02156_),
    .Y(_02158_));
 sg13g2_nor2_1 _22532_ (.A(_06257_),
    .B(_02025_),
    .Y(_02159_));
 sg13g2_inv_1 _22533_ (.Y(_02160_),
    .A(_06746_));
 sg13g2_nor2_1 _22534_ (.A(\b.gen_square[51].sq.color ),
    .B(net31),
    .Y(_02161_));
 sg13g2_a21o_1 _22535_ (.A2(net31),
    .A1(_02160_),
    .B1(_02161_),
    .X(_02162_));
 sg13g2_inv_1 _22536_ (.Y(_02163_),
    .A(_02162_));
 sg13g2_inv_1 _22537_ (.Y(_02164_),
    .A(_04999_));
 sg13g2_o21ai_1 _22538_ (.B1(_02164_),
    .Y(_02165_),
    .A1(_06247_),
    .A2(_02163_));
 sg13g2_nor3_1 _22539_ (.A(_04562_),
    .B(_02159_),
    .C(_02165_),
    .Y(_02167_));
 sg13g2_nor2_1 _22540_ (.A(_06247_),
    .B(_02162_),
    .Y(_02168_));
 sg13g2_nor2_1 _22541_ (.A(_04376_),
    .B(_02080_),
    .Y(_02169_));
 sg13g2_nor2_1 _22542_ (.A(_06257_),
    .B(_02026_),
    .Y(_02170_));
 sg13g2_nor4_1 _22543_ (.A(_06830_),
    .B(_05067_),
    .C(_02169_),
    .D(_02170_),
    .Y(_02171_));
 sg13g2_nor2b_1 _22544_ (.A(_02168_),
    .B_N(_02171_),
    .Y(_02172_));
 sg13g2_nor2_1 _22545_ (.A(_04376_),
    .B(_02079_),
    .Y(_02173_));
 sg13g2_nor2_1 _22546_ (.A(_06825_),
    .B(_02173_),
    .Y(_02174_));
 sg13g2_nand3_1 _22547_ (.B(_02172_),
    .C(_02174_),
    .A(_02167_),
    .Y(_02175_));
 sg13g2_nor2_1 _22548_ (.A(net48),
    .B(_04563_),
    .Y(_02176_));
 sg13g2_nand3_1 _22549_ (.B(_02175_),
    .C(_02176_),
    .A(_02158_),
    .Y(_02178_));
 sg13g2_nor2b_1 _22550_ (.A(_02163_),
    .B_N(_02139_),
    .Y(_02179_));
 sg13g2_nand2_1 _22551_ (.Y(_02180_),
    .A(_02026_),
    .B(_02008_));
 sg13g2_a21oi_1 _22552_ (.A1(_07259_),
    .A2(net77),
    .Y(_02181_),
    .B1(_04728_));
 sg13g2_nand2b_1 _22553_ (.Y(_02182_),
    .B(_02138_),
    .A_N(_02181_));
 sg13g2_nor3_1 _22554_ (.A(_05183_),
    .B(_06625_),
    .C(_01688_),
    .Y(_02183_));
 sg13g2_nand3_1 _22555_ (.B(_02182_),
    .C(_02183_),
    .A(_02180_),
    .Y(_02184_));
 sg13g2_nor4_1 _22556_ (.A(_02159_),
    .B(_02179_),
    .C(_02184_),
    .D(_02165_),
    .Y(_02185_));
 sg13g2_and3_1 _22557_ (.X(_02186_),
    .A(_02151_),
    .B(_02174_),
    .C(_02185_));
 sg13g2_inv_1 _22558_ (.Y(_02187_),
    .A(_02172_));
 sg13g2_nand3_1 _22559_ (.B(_07832_),
    .C(_07622_),
    .A(_01702_),
    .Y(_02189_));
 sg13g2_a221oi_1 _22560_ (.B2(_02139_),
    .C1(_02189_),
    .B1(_02163_),
    .A1(_02138_),
    .Y(_02190_),
    .A2(_02181_));
 sg13g2_o21ai_1 _22561_ (.B1(_02190_),
    .Y(_02191_),
    .A1(_02026_),
    .A2(_02009_));
 sg13g2_nor3_1 _22562_ (.A(_02187_),
    .B(_02191_),
    .C(_02149_),
    .Y(_02192_));
 sg13g2_nand2_1 _22563_ (.Y(_02193_),
    .A(_02186_),
    .B(_02192_));
 sg13g2_nand2_1 _22564_ (.Y(_02194_),
    .A(_04993_),
    .B(_04552_));
 sg13g2_nand3_1 _22565_ (.B(net57),
    .C(_02194_),
    .A(_02193_),
    .Y(_02195_));
 sg13g2_a21o_1 _22566_ (.A2(_04993_),
    .A1(_04555_),
    .B1(_02195_),
    .X(_02196_));
 sg13g2_nor3_1 _22567_ (.A(_04552_),
    .B(_02192_),
    .C(_02186_),
    .Y(_02197_));
 sg13g2_nand3_1 _22568_ (.B(net97),
    .C(_04556_),
    .A(_02197_),
    .Y(_02198_));
 sg13g2_nand3_1 _22569_ (.B(_02196_),
    .C(_02198_),
    .A(_02178_),
    .Y(_02200_));
 sg13g2_nor2b_1 _22570_ (.A(_02136_),
    .B_N(_02200_),
    .Y(_02201_));
 sg13g2_buf_1 _22571_ (.A(\b.gen_square[59].sq.mask ),
    .X(_02202_));
 sg13g2_inv_1 _22572_ (.Y(_02203_),
    .A(_02202_));
 sg13g2_nor2_1 _22573_ (.A(\b.gen_square[50].sq.color ),
    .B(net45),
    .Y(_02204_));
 sg13g2_a21o_1 _22574_ (.A2(net45),
    .A1(_06302_),
    .B1(_02204_),
    .X(_02205_));
 sg13g2_buf_1 _22575_ (.A(_02205_),
    .X(_02206_));
 sg13g2_inv_1 _22576_ (.Y(_02207_),
    .A(_05543_));
 sg13g2_a21oi_1 _22577_ (.A1(_02206_),
    .A2(_02207_),
    .Y(_02208_),
    .B1(_06825_));
 sg13g2_inv_1 _22578_ (.Y(_02209_),
    .A(_02208_));
 sg13g2_o21ai_1 _22579_ (.B1(_06251_),
    .Y(_02211_),
    .A1(_06787_),
    .A2(_02082_));
 sg13g2_nand2b_1 _22580_ (.Y(_02212_),
    .B(_05196_),
    .A_N(_02211_));
 sg13g2_nor2_1 _22581_ (.A(_05543_),
    .B(_02206_),
    .Y(_02213_));
 sg13g2_nand2_1 _22582_ (.Y(_02214_),
    .A(_02101_),
    .B(_05766_));
 sg13g2_nor4_1 _22583_ (.A(_06454_),
    .B(_06830_),
    .C(_02213_),
    .D(_02214_),
    .Y(_02215_));
 sg13g2_inv_1 _22584_ (.Y(_02216_),
    .A(_02215_));
 sg13g2_nor4_1 _22585_ (.A(_05492_),
    .B(_02209_),
    .C(_02212_),
    .D(_02216_),
    .Y(_02217_));
 sg13g2_o21ai_1 _22586_ (.B1(_07866_),
    .Y(_02218_),
    .A1(_08085_),
    .A2(_06307_));
 sg13g2_inv_1 _22587_ (.Y(_02219_),
    .A(_02218_));
 sg13g2_inv_1 _22588_ (.Y(_02220_),
    .A(_06871_));
 sg13g2_a21oi_1 _22589_ (.A1(_02220_),
    .A2(net23),
    .Y(_02221_),
    .B1(_08020_));
 sg13g2_o21ai_1 _22590_ (.B1(_05187_),
    .Y(_02222_),
    .A1(_02219_),
    .A2(_02221_));
 sg13g2_nor2_1 _22591_ (.A(_06268_),
    .B(_02222_),
    .Y(_02223_));
 sg13g2_a21o_1 _22592_ (.A2(_04995_),
    .A1(_02143_),
    .B1(_02010_),
    .X(_02224_));
 sg13g2_buf_1 _22593_ (.A(_02224_),
    .X(_02225_));
 sg13g2_nand2_1 _22594_ (.Y(_02226_),
    .A(_02225_),
    .B(_02006_));
 sg13g2_a21oi_1 _22595_ (.A1(_06838_),
    .A2(net31),
    .Y(_02227_),
    .B1(_04776_));
 sg13g2_o21ai_1 _22596_ (.B1(_05187_),
    .Y(_02228_),
    .A1(_02226_),
    .A2(_02227_));
 sg13g2_a21oi_1 _22597_ (.A1(_02228_),
    .A2(_02222_),
    .Y(_02229_),
    .B1(_06272_));
 sg13g2_nor3_1 _22598_ (.A(_05196_),
    .B(_02223_),
    .C(_02229_),
    .Y(_02230_));
 sg13g2_nor4_1 _22599_ (.A(net63),
    .B(_05197_),
    .C(_02217_),
    .D(_02230_),
    .Y(_02232_));
 sg13g2_a21oi_1 _22600_ (.A1(_07040_),
    .A2(net23),
    .Y(_02233_),
    .B1(_04702_));
 sg13g2_nand2b_1 _22601_ (.Y(_02234_),
    .B(_02221_),
    .A_N(_02233_));
 sg13g2_nand2_1 _22602_ (.Y(_02235_),
    .A(_02206_),
    .B(_02219_));
 sg13g2_nor2b_1 _22603_ (.A(_01619_),
    .B_N(_11770_),
    .Y(_02236_));
 sg13g2_o21ai_1 _22604_ (.B1(_02022_),
    .Y(_02237_),
    .A1(_07373_),
    .A2(_02005_));
 sg13g2_nand4_1 _22605_ (.B(_02235_),
    .C(_02236_),
    .A(_02234_),
    .Y(_02238_),
    .D(_02237_));
 sg13g2_a21oi_1 _22606_ (.A1(_06820_),
    .A2(net31),
    .Y(_02239_),
    .B1(_04678_));
 sg13g2_nand2b_1 _22607_ (.Y(_02240_),
    .B(_02227_),
    .A_N(_02239_));
 sg13g2_o21ai_1 _22608_ (.B1(_02240_),
    .Y(_02241_),
    .A1(_02225_),
    .A2(_02082_));
 sg13g2_nor4_1 _22609_ (.A(_02211_),
    .B(_02209_),
    .C(_02238_),
    .D(_02241_),
    .Y(_02243_));
 sg13g2_inv_1 _22610_ (.Y(_02244_),
    .A(_02243_));
 sg13g2_nor2_1 _22611_ (.A(_02006_),
    .B(_02022_),
    .Y(_02245_));
 sg13g2_nand2_1 _22612_ (.Y(_02246_),
    .A(_02221_),
    .B(_02233_));
 sg13g2_nand2b_1 _22613_ (.Y(_02247_),
    .B(_02219_),
    .A_N(_02206_));
 sg13g2_nand4_1 _22614_ (.B(_02247_),
    .C(_11732_),
    .A(_02246_),
    .Y(_02248_),
    .D(_01613_));
 sg13g2_inv_1 _22615_ (.Y(_02249_),
    .A(_02225_));
 sg13g2_a22oi_1 _22616_ (.Y(_02250_),
    .B1(_02227_),
    .B2(_02239_),
    .A2(_02082_),
    .A1(_02249_));
 sg13g2_inv_1 _22617_ (.Y(_02251_),
    .A(_02250_));
 sg13g2_nor4_1 _22618_ (.A(_02245_),
    .B(_02216_),
    .C(_02248_),
    .D(_02251_),
    .Y(_02252_));
 sg13g2_inv_1 _22619_ (.Y(_02254_),
    .A(_02252_));
 sg13g2_nand4_1 _22620_ (.B(net114),
    .C(_06254_),
    .A(_02244_),
    .Y(_02255_),
    .D(_02254_));
 sg13g2_buf_1 _22621_ (.A(_02255_),
    .X(_02256_));
 sg13g2_nor2_1 _22622_ (.A(_05190_),
    .B(_02256_),
    .Y(_02257_));
 sg13g2_nor2_1 _22623_ (.A(_06259_),
    .B(_06254_),
    .Y(_02258_));
 sg13g2_nor2_1 _22624_ (.A(_05191_),
    .B(_06259_),
    .Y(_02259_));
 sg13g2_nor2_1 _22625_ (.A(_02254_),
    .B(_02244_),
    .Y(_02260_));
 sg13g2_nor4_1 _22626_ (.A(net142),
    .B(_02258_),
    .C(_02259_),
    .D(_02260_),
    .Y(_02261_));
 sg13g2_nor3_1 _22627_ (.A(_02232_),
    .B(_02257_),
    .C(_02261_),
    .Y(_02262_));
 sg13g2_nor2_1 _22628_ (.A(_02203_),
    .B(_02262_),
    .Y(_02263_));
 sg13g2_inv_1 _22629_ (.Y(_02265_),
    .A(\b.gen_square[57].sq.mask ));
 sg13g2_a21oi_1 _22630_ (.A1(_06446_),
    .A2(_04651_),
    .Y(_02266_),
    .B1(_04654_));
 sg13g2_inv_1 _22631_ (.Y(_02267_),
    .A(_02266_));
 sg13g2_a21oi_1 _22632_ (.A1(_06243_),
    .A2(_04651_),
    .Y(_02268_),
    .B1(_07867_));
 sg13g2_a21oi_1 _22633_ (.A1(_05700_),
    .A2(net87),
    .Y(_02269_),
    .B1(_04754_));
 sg13g2_o21ai_1 _22634_ (.B1(_04628_),
    .Y(_02270_),
    .A1(_04627_),
    .A2(_05726_));
 sg13g2_a22oi_1 _22635_ (.Y(_02271_),
    .B1(_02269_),
    .B2(_02270_),
    .A2(_02268_),
    .A1(_02267_));
 sg13g2_nor2b_1 _22636_ (.A(_05445_),
    .B_N(_05978_),
    .Y(_02272_));
 sg13g2_a21oi_1 _22637_ (.A1(_02083_),
    .A2(_06262_),
    .Y(_02273_),
    .B1(_02024_));
 sg13g2_a21oi_1 _22638_ (.A1(_02273_),
    .A2(_02003_),
    .Y(_02274_),
    .B1(_05491_));
 sg13g2_inv_1 _22639_ (.Y(_02275_),
    .A(_02274_));
 sg13g2_a21oi_1 _22640_ (.A1(_02225_),
    .A2(_06262_),
    .Y(_02276_),
    .B1(_02007_));
 sg13g2_inv_1 _22641_ (.Y(_02277_),
    .A(_02276_));
 sg13g2_a21oi_1 _22642_ (.A1(_02277_),
    .A2(_02003_),
    .Y(_02278_),
    .B1(_02004_));
 sg13g2_inv_1 _22643_ (.Y(_02279_),
    .A(_02278_));
 sg13g2_nor2_1 _22644_ (.A(_02275_),
    .B(_02279_),
    .Y(_02280_));
 sg13g2_nor4_1 _22645_ (.A(_05546_),
    .B(_05945_),
    .C(_05492_),
    .D(_02280_),
    .Y(_02281_));
 sg13g2_nor4_1 _22646_ (.A(_06289_),
    .B(_01352_),
    .C(_05507_),
    .D(_07928_),
    .Y(_02282_));
 sg13g2_nand4_1 _22647_ (.B(_02272_),
    .C(_02281_),
    .A(_02271_),
    .Y(_02283_),
    .D(_02282_));
 sg13g2_inv_1 _22648_ (.Y(_02284_),
    .A(_05453_));
 sg13g2_inv_1 _22649_ (.Y(_02286_),
    .A(_05941_));
 sg13g2_nor2_1 _22650_ (.A(_02286_),
    .B(_02269_),
    .Y(_02287_));
 sg13g2_nor2_1 _22651_ (.A(_07911_),
    .B(_11958_),
    .Y(_02288_));
 sg13g2_nor2_1 _22652_ (.A(_05781_),
    .B(_01339_),
    .Y(_02289_));
 sg13g2_nand3_1 _22653_ (.B(_01341_),
    .C(_02289_),
    .A(_02288_),
    .Y(_02290_));
 sg13g2_inv_1 _22654_ (.Y(_02291_),
    .A(_02268_));
 sg13g2_a21oi_1 _22655_ (.A1(_02291_),
    .A2(_05543_),
    .Y(_02292_),
    .B1(_02267_));
 sg13g2_a21oi_1 _22656_ (.A1(_02279_),
    .A2(_05484_),
    .Y(_02293_),
    .B1(_02274_));
 sg13g2_nor4_1 _22657_ (.A(_06131_),
    .B(_02290_),
    .C(_02292_),
    .D(_02293_),
    .Y(_02294_));
 sg13g2_o21ai_1 _22658_ (.B1(_02294_),
    .Y(_02295_),
    .A1(_02270_),
    .A2(_02287_));
 sg13g2_nand3_1 _22659_ (.B(_02284_),
    .C(_02295_),
    .A(_02283_),
    .Y(_02297_));
 sg13g2_nor2_1 _22660_ (.A(net192),
    .B(_02297_),
    .Y(_02298_));
 sg13g2_nor2_1 _22661_ (.A(_05931_),
    .B(_05459_),
    .Y(_02299_));
 sg13g2_or2_1 _22662_ (.X(_02300_),
    .B(_02283_),
    .A(_02295_));
 sg13g2_buf_1 _22663_ (.A(_02300_),
    .X(_02301_));
 sg13g2_nand2b_1 _22664_ (.Y(_02302_),
    .B(_05453_),
    .A_N(_05459_));
 sg13g2_nand3_1 _22665_ (.B(net76),
    .C(_02302_),
    .A(_02301_),
    .Y(_02303_));
 sg13g2_nand2_1 _22666_ (.Y(_02304_),
    .A(_02279_),
    .B(_05977_));
 sg13g2_o21ai_1 _22667_ (.B1(_05453_),
    .Y(_02305_),
    .A1(_02304_),
    .A2(_02269_));
 sg13g2_a21oi_1 _22668_ (.A1(_02291_),
    .A2(_08028_),
    .Y(_02306_),
    .B1(_02284_));
 sg13g2_inv_1 _22669_ (.Y(_02308_),
    .A(_02306_));
 sg13g2_a21o_1 _22670_ (.A2(_02308_),
    .A1(_02305_),
    .B1(_05475_),
    .X(_02309_));
 sg13g2_nand2b_1 _22671_ (.Y(_02310_),
    .B(_02306_),
    .A_N(_05932_));
 sg13g2_nand3_1 _22672_ (.B(_05451_),
    .C(_02310_),
    .A(_02309_),
    .Y(_02311_));
 sg13g2_nor3_1 _22673_ (.A(_05451_),
    .B(_02286_),
    .C(_07373_),
    .Y(_02312_));
 sg13g2_nand3_1 _22674_ (.B(_05543_),
    .C(_07332_),
    .A(_02312_),
    .Y(_02313_));
 sg13g2_nor2_1 _22675_ (.A(net83),
    .B(_05454_),
    .Y(_02314_));
 sg13g2_nand3_1 _22676_ (.B(_02313_),
    .C(_02314_),
    .A(_02311_),
    .Y(_02315_));
 sg13g2_o21ai_1 _22677_ (.B1(_02315_),
    .Y(_02316_),
    .A1(_02299_),
    .A2(_02303_));
 sg13g2_a21oi_1 _22678_ (.A1(_05931_),
    .A2(_02298_),
    .Y(_02317_),
    .B1(_02316_));
 sg13g2_nor2_1 _22679_ (.A(_02265_),
    .B(_02317_),
    .Y(_02319_));
 sg13g2_nor3_1 _22680_ (.A(_05782_),
    .B(_01382_),
    .C(_01379_),
    .Y(_02320_));
 sg13g2_inv_1 _22681_ (.Y(_02321_),
    .A(_02320_));
 sg13g2_nor2_1 _22682_ (.A(_08268_),
    .B(_06651_),
    .Y(_02322_));
 sg13g2_inv_1 _22683_ (.Y(_02323_),
    .A(_02322_));
 sg13g2_a21oi_1 _22684_ (.A1(_05540_),
    .A2(net87),
    .Y(_02324_),
    .B1(_01377_));
 sg13g2_a21oi_1 _22685_ (.A1(_05516_),
    .A2(net87),
    .Y(_02325_),
    .B1(_08380_));
 sg13g2_nor2b_1 _22686_ (.A(_02324_),
    .B_N(_02325_),
    .Y(_02326_));
 sg13g2_inv_1 _22687_ (.Y(_02327_),
    .A(_08182_));
 sg13g2_a21oi_1 _22688_ (.A1(_06130_),
    .A2(_04606_),
    .Y(_02328_),
    .B1(_02327_));
 sg13g2_a21oi_1 _22689_ (.A1(_06117_),
    .A2(_04606_),
    .Y(_02329_),
    .B1(_08221_));
 sg13g2_a21oi_1 _22690_ (.A1(_02275_),
    .A2(_01998_),
    .Y(_02330_),
    .B1(_05464_));
 sg13g2_a21o_1 _22691_ (.A2(_01998_),
    .A1(_02279_),
    .B1(_01999_),
    .X(_02331_));
 sg13g2_nor2_1 _22692_ (.A(_02330_),
    .B(_02331_),
    .Y(_02332_));
 sg13g2_a21oi_1 _22693_ (.A1(_02328_),
    .A2(_02329_),
    .Y(_02333_),
    .B1(_02332_));
 sg13g2_inv_1 _22694_ (.Y(_02334_),
    .A(_02333_));
 sg13g2_nor4_1 _22695_ (.A(_02321_),
    .B(_02323_),
    .C(_02326_),
    .D(_02334_),
    .Y(_02335_));
 sg13g2_inv_1 _22696_ (.Y(_02336_),
    .A(_02335_));
 sg13g2_inv_1 _22697_ (.Y(_02337_),
    .A(_02329_));
 sg13g2_nor2b_1 _22698_ (.A(_02331_),
    .B_N(_02330_),
    .Y(_02338_));
 sg13g2_a21oi_1 _22699_ (.A1(_02328_),
    .A2(_02337_),
    .Y(_02340_),
    .B1(_02338_));
 sg13g2_nor3_1 _22700_ (.A(_05470_),
    .B(_01400_),
    .C(_01402_),
    .Y(_02341_));
 sg13g2_inv_1 _22701_ (.Y(_02342_),
    .A(_08420_));
 sg13g2_a21oi_1 _22702_ (.A1(_02324_),
    .A2(_02325_),
    .Y(_02343_),
    .B1(_02342_));
 sg13g2_nand3_1 _22703_ (.B(_02341_),
    .C(_02343_),
    .A(_02340_),
    .Y(_02344_));
 sg13g2_and3_1 _22704_ (.X(_02345_),
    .A(_02336_),
    .B(_05441_),
    .C(_02344_));
 sg13g2_buf_1 _22705_ (.A(_02345_),
    .X(_02346_));
 sg13g2_inv_1 _22706_ (.Y(_02347_),
    .A(_05427_));
 sg13g2_a21oi_1 _22707_ (.A1(_02346_),
    .A2(net130),
    .Y(_02348_),
    .B1(_02347_));
 sg13g2_nor2_1 _22708_ (.A(_02344_),
    .B(_02336_),
    .Y(_02349_));
 sg13g2_nor2_1 _22709_ (.A(_05263_),
    .B(_02349_),
    .Y(_02351_));
 sg13g2_a22oi_1 _22710_ (.Y(_02352_),
    .B1(net130),
    .B2(_02346_),
    .A2(net86),
    .A1(_02351_));
 sg13g2_nand2b_1 _22711_ (.Y(_02353_),
    .B(_05426_),
    .A_N(_05255_));
 sg13g2_nand2b_1 _22712_ (.Y(_02354_),
    .B(_02353_),
    .A_N(_02352_));
 sg13g2_a21o_1 _22713_ (.A2(_02340_),
    .A1(_02333_),
    .B1(_05441_),
    .X(_02355_));
 sg13g2_nand2_1 _22714_ (.Y(_02356_),
    .A(_02325_),
    .B(_05263_));
 sg13g2_a21o_1 _22715_ (.A2(_02356_),
    .A1(_02355_),
    .B1(_05257_),
    .X(_02357_));
 sg13g2_o21ai_1 _22716_ (.B1(_02357_),
    .Y(_02358_),
    .A1(_05973_),
    .A2(_02355_));
 sg13g2_nand3_1 _22717_ (.B(net85),
    .C(_05266_),
    .A(_02358_),
    .Y(_02359_));
 sg13g2_o21ai_1 _22718_ (.B1(_02359_),
    .Y(_02360_),
    .A1(_02348_),
    .A2(_02354_));
 sg13g2_buf_1 _22719_ (.A(\b.gen_square[56].sq.mask ),
    .X(_02362_));
 sg13g2_nand2_1 _22720_ (.Y(_02363_),
    .A(_02360_),
    .B(_02362_));
 sg13g2_nand3_1 _22721_ (.B(net76),
    .C(_02284_),
    .A(_02301_),
    .Y(_02364_));
 sg13g2_inv_1 _22722_ (.Y(_02365_),
    .A(_02298_));
 sg13g2_nand2_1 _22723_ (.Y(_02366_),
    .A(_02364_),
    .B(_02365_));
 sg13g2_nand2_1 _22724_ (.Y(_02367_),
    .A(_02365_),
    .B(_05459_));
 sg13g2_nand2b_1 _22725_ (.Y(_02368_),
    .B(_05458_),
    .A_N(_05474_));
 sg13g2_nand3_1 _22726_ (.B(_02367_),
    .C(_02368_),
    .A(_02366_),
    .Y(_02369_));
 sg13g2_nand2_1 _22727_ (.Y(_02370_),
    .A(_05451_),
    .B(net85));
 sg13g2_o21ai_1 _22728_ (.B1(_02309_),
    .Y(_02371_),
    .A1(_05473_),
    .A2(_02305_));
 sg13g2_nand2b_1 _22729_ (.Y(_02373_),
    .B(_02371_),
    .A_N(_02370_));
 sg13g2_a21o_1 _22730_ (.A2(_02373_),
    .A1(_02369_),
    .B1(_02265_),
    .X(_02374_));
 sg13g2_buf_1 _22731_ (.A(_02374_),
    .X(_02375_));
 sg13g2_nor2b_1 _22732_ (.A(_02363_),
    .B_N(_02375_),
    .Y(_02376_));
 sg13g2_inv_1 _22733_ (.Y(_02377_),
    .A(_02362_));
 sg13g2_inv_1 _22734_ (.Y(_02378_),
    .A(_05254_));
 sg13g2_a21oi_1 _22735_ (.A1(_02351_),
    .A2(_02378_),
    .Y(_02379_),
    .B1(_05427_));
 sg13g2_a21oi_1 _22736_ (.A1(_05427_),
    .A2(_02349_),
    .Y(_02380_),
    .B1(_02379_));
 sg13g2_nor2_1 _22737_ (.A(_05260_),
    .B(_02356_),
    .Y(_02381_));
 sg13g2_inv_1 _22738_ (.Y(_02382_),
    .A(_02381_));
 sg13g2_nand3_1 _22739_ (.B(_05266_),
    .C(_02382_),
    .A(_02357_),
    .Y(_02383_));
 sg13g2_nand2_1 _22740_ (.Y(_02384_),
    .A(_02341_),
    .B(_02320_));
 sg13g2_a21o_1 _22741_ (.A2(_05263_),
    .A1(_02384_),
    .B1(_05266_),
    .X(_02385_));
 sg13g2_nand3_1 _22742_ (.B(net85),
    .C(_02385_),
    .A(_02383_),
    .Y(_02386_));
 sg13g2_nand3_1 _22743_ (.B(net130),
    .C(_02378_),
    .A(_02346_),
    .Y(_02387_));
 sg13g2_nand2_1 _22744_ (.Y(_02388_),
    .A(_02386_),
    .B(_02387_));
 sg13g2_a21oi_1 _22745_ (.A1(net76),
    .A2(_02380_),
    .Y(_02389_),
    .B1(_02388_));
 sg13g2_o21ai_1 _22746_ (.B1(_02319_),
    .Y(_02390_),
    .A1(_02377_),
    .A2(_02389_));
 sg13g2_xnor2_1 _22747_ (.Y(_02391_),
    .A(_05425_),
    .B(_05255_));
 sg13g2_o21ai_1 _22748_ (.B1(_06283_),
    .Y(_02392_),
    .A1(_02323_),
    .A2(_02342_));
 sg13g2_nand3b_1 _22749_ (.B(_02392_),
    .C(_02382_),
    .Y(_02394_),
    .A_N(_02358_));
 sg13g2_nand3_1 _22750_ (.B(net85),
    .C(_05266_),
    .A(_02394_),
    .Y(_02395_));
 sg13g2_o21ai_1 _22751_ (.B1(_02395_),
    .Y(_02396_),
    .A1(_02391_),
    .A2(_02352_));
 sg13g2_nand2_1 _22752_ (.Y(_02397_),
    .A(_02396_),
    .B(_02362_));
 sg13g2_xnor2_1 _22753_ (.Y(_02398_),
    .A(_05448_),
    .B(_05474_));
 sg13g2_nor2_1 _22754_ (.A(_06289_),
    .B(_07928_),
    .Y(_02399_));
 sg13g2_a21o_1 _22755_ (.A2(_02399_),
    .A1(_02288_),
    .B1(_06626_),
    .X(_02400_));
 sg13g2_a21oi_1 _22756_ (.A1(_02310_),
    .A2(_02400_),
    .Y(_02401_),
    .B1(_02370_));
 sg13g2_a21oi_1 _22757_ (.A1(_02366_),
    .A2(_02398_),
    .Y(_02402_),
    .B1(_02401_));
 sg13g2_nand2_1 _22758_ (.Y(_02403_),
    .A(_02402_),
    .B(_02373_));
 sg13g2_nand2_1 _22759_ (.Y(_02405_),
    .A(_02403_),
    .B(\b.gen_square[57].sq.mask ));
 sg13g2_inv_1 _22760_ (.Y(_02406_),
    .A(_02405_));
 sg13g2_inv_1 _22761_ (.Y(_02407_),
    .A(_02363_));
 sg13g2_nor2_1 _22762_ (.A(_02375_),
    .B(_02407_),
    .Y(_02408_));
 sg13g2_a21oi_1 _22763_ (.A1(_02397_),
    .A2(_02406_),
    .Y(_02409_),
    .B1(_02408_));
 sg13g2_o21ai_1 _22764_ (.B1(_02409_),
    .Y(_02410_),
    .A1(_02376_),
    .A2(_02390_));
 sg13g2_inv_1 _22765_ (.Y(_02411_),
    .A(_02397_));
 sg13g2_nand2_1 _22766_ (.Y(_02412_),
    .A(_02411_),
    .B(_02405_));
 sg13g2_nand2_1 _22767_ (.Y(_02413_),
    .A(_02410_),
    .B(_02412_));
 sg13g2_inv_1 _22768_ (.Y(_02414_),
    .A(_02413_));
 sg13g2_nor3_1 _22769_ (.A(_02377_),
    .B(_02389_),
    .C(_02414_),
    .Y(_02416_));
 sg13g2_a21o_1 _22770_ (.A2(_02414_),
    .A1(_02319_),
    .B1(_02416_),
    .X(_02417_));
 sg13g2_buf_1 _22771_ (.A(\b.gen_square[58].sq.mask ),
    .X(_02418_));
 sg13g2_inv_1 _22772_ (.Y(_02419_),
    .A(_02418_));
 sg13g2_nor2_1 _22773_ (.A(_05546_),
    .B(_02159_),
    .Y(_02420_));
 sg13g2_inv_1 _22774_ (.Y(_02421_),
    .A(_02420_));
 sg13g2_nand3_1 _22775_ (.B(_05481_),
    .C(_06266_),
    .A(_01403_),
    .Y(_02422_));
 sg13g2_nor4_1 _22776_ (.A(_05768_),
    .B(_06454_),
    .C(_05782_),
    .D(_02170_),
    .Y(_02423_));
 sg13g2_nand2_1 _22777_ (.Y(_02424_),
    .A(_02423_),
    .B(_01380_));
 sg13g2_nor4_1 _22778_ (.A(_02421_),
    .B(_06250_),
    .C(_02422_),
    .D(_02424_),
    .Y(_02425_));
 sg13g2_a21oi_1 _22779_ (.A1(_05252_),
    .A2(net87),
    .Y(_02427_),
    .B1(_08380_));
 sg13g2_a21oi_1 _22780_ (.A1(_06719_),
    .A2(net31),
    .Y(_02428_),
    .B1(_07694_));
 sg13g2_o21ai_1 _22781_ (.B1(_05214_),
    .Y(_02429_),
    .A1(_02427_),
    .A2(_02428_));
 sg13g2_nor2_1 _22782_ (.A(_05222_),
    .B(_02429_),
    .Y(_02430_));
 sg13g2_nand2_1 _22783_ (.Y(_02431_),
    .A(_02277_),
    .B(_02002_));
 sg13g2_a21oi_1 _22784_ (.A1(_06416_),
    .A2(net45),
    .Y(_02432_),
    .B1(_04765_));
 sg13g2_o21ai_1 _22785_ (.B1(_05214_),
    .Y(_02433_),
    .A1(_02431_),
    .A2(_02432_));
 sg13g2_a21oi_1 _22786_ (.A1(_02433_),
    .A2(_02429_),
    .Y(_02434_),
    .B1(_05219_));
 sg13g2_nor3_1 _22787_ (.A(_02430_),
    .B(_05481_),
    .C(_02434_),
    .Y(_02435_));
 sg13g2_nor4_1 _22788_ (.A(net72),
    .B(_05227_),
    .C(_02425_),
    .D(_02435_),
    .Y(_02436_));
 sg13g2_nor2_1 _22789_ (.A(_02002_),
    .B(_02020_),
    .Y(_02438_));
 sg13g2_a21oi_1 _22790_ (.A1(_06770_),
    .A2(net31),
    .Y(_02439_),
    .B1(_04678_));
 sg13g2_a22oi_1 _22791_ (.Y(_02440_),
    .B1(_02428_),
    .B2(_02439_),
    .A2(_01401_),
    .A1(_02427_));
 sg13g2_nor2_1 _22792_ (.A(_06651_),
    .B(_05208_),
    .Y(_02441_));
 sg13g2_nor2_1 _22793_ (.A(_08272_),
    .B(_07830_),
    .Y(_02442_));
 sg13g2_nand3_1 _22794_ (.B(_02441_),
    .C(_02442_),
    .A(_02440_),
    .Y(_02443_));
 sg13g2_a21oi_1 _22795_ (.A1(_06439_),
    .A2(net45),
    .Y(_02444_),
    .B1(_04654_));
 sg13g2_a22oi_1 _22796_ (.Y(_02445_),
    .B1(_02432_),
    .B2(_02444_),
    .A2(_02273_),
    .A1(_02276_));
 sg13g2_inv_1 _22797_ (.Y(_02446_),
    .A(_02445_));
 sg13g2_nor4_1 _22798_ (.A(_02438_),
    .B(_02424_),
    .C(_02443_),
    .D(_02446_),
    .Y(_02447_));
 sg13g2_inv_1 _22799_ (.Y(_02449_),
    .A(_02447_));
 sg13g2_nand2b_1 _22800_ (.Y(_02450_),
    .B(_02428_),
    .A_N(_02439_));
 sg13g2_nand2b_1 _22801_ (.Y(_02451_),
    .B(_02276_),
    .A_N(_02273_));
 sg13g2_nor2b_1 _22802_ (.A(_01401_),
    .B_N(_02427_),
    .Y(_02452_));
 sg13g2_a21oi_1 _22803_ (.A1(_02002_),
    .A2(_05469_),
    .Y(_02453_),
    .B1(_02021_));
 sg13g2_nor2_1 _22804_ (.A(_11811_),
    .B(_01487_),
    .Y(_02454_));
 sg13g2_nand2_1 _22805_ (.Y(_02455_),
    .A(_02454_),
    .B(_01403_));
 sg13g2_nor4_1 _22806_ (.A(_02452_),
    .B(_06250_),
    .C(_02453_),
    .D(_02455_),
    .Y(_02456_));
 sg13g2_nand3_1 _22807_ (.B(_02451_),
    .C(_02456_),
    .A(_02450_),
    .Y(_02457_));
 sg13g2_nor2b_1 _22808_ (.A(_02444_),
    .B_N(_02432_),
    .Y(_02458_));
 sg13g2_nor3_1 _22809_ (.A(_02421_),
    .B(_02457_),
    .C(_02458_),
    .Y(_02460_));
 sg13g2_inv_1 _22810_ (.Y(_02461_),
    .A(_02460_));
 sg13g2_nand4_1 _22811_ (.B(net130),
    .C(_05482_),
    .A(_02449_),
    .Y(_02462_),
    .D(_02461_));
 sg13g2_buf_1 _22812_ (.A(_02462_),
    .X(_02463_));
 sg13g2_nor2_1 _22813_ (.A(_05216_),
    .B(_02463_),
    .Y(_02464_));
 sg13g2_nor2_1 _22814_ (.A(_05486_),
    .B(_05482_),
    .Y(_02465_));
 sg13g2_nor2_1 _22815_ (.A(_05221_),
    .B(_05486_),
    .Y(_02466_));
 sg13g2_nor2_1 _22816_ (.A(_02461_),
    .B(_02449_),
    .Y(_02467_));
 sg13g2_nor4_1 _22817_ (.A(net142),
    .B(_02465_),
    .C(_02466_),
    .D(_02467_),
    .Y(_02468_));
 sg13g2_nor3_1 _22818_ (.A(_02436_),
    .B(_02464_),
    .C(_02468_),
    .Y(_02469_));
 sg13g2_nor2_1 _22819_ (.A(_02419_),
    .B(_02469_),
    .Y(_02471_));
 sg13g2_nand2_1 _22820_ (.Y(_02472_),
    .A(_05482_),
    .B(net68));
 sg13g2_o21ai_1 _22821_ (.B1(_02463_),
    .Y(_02473_),
    .A1(_02467_),
    .A2(_02472_));
 sg13g2_nand2_1 _22822_ (.Y(_02474_),
    .A(_02463_),
    .B(_05486_));
 sg13g2_nand2b_1 _22823_ (.Y(_02475_),
    .B(_05485_),
    .A_N(_05217_));
 sg13g2_nand3_1 _22824_ (.B(_02474_),
    .C(_02475_),
    .A(_02473_),
    .Y(_02476_));
 sg13g2_nor3_1 _22825_ (.A(_05218_),
    .B(_05485_),
    .C(_02433_),
    .Y(_02477_));
 sg13g2_or2_1 _22826_ (.X(_02478_),
    .B(_02434_),
    .A(_02477_));
 sg13g2_nand3_1 _22827_ (.B(net75),
    .C(_05226_),
    .A(_02478_),
    .Y(_02479_));
 sg13g2_nand2_1 _22828_ (.Y(_02480_),
    .A(_02476_),
    .B(_02479_));
 sg13g2_nand2_1 _22829_ (.Y(_02482_),
    .A(_02480_),
    .B(_02418_));
 sg13g2_nor2_1 _22830_ (.A(_02375_),
    .B(_02413_),
    .Y(_02483_));
 sg13g2_a21oi_1 _22831_ (.A1(_02407_),
    .A2(_02413_),
    .Y(_02484_),
    .B1(_02483_));
 sg13g2_inv_1 _22832_ (.Y(_02485_),
    .A(_02484_));
 sg13g2_nor2_1 _22833_ (.A(_02482_),
    .B(_02485_),
    .Y(_02486_));
 sg13g2_nor2b_1 _22834_ (.A(_02417_),
    .B_N(_02471_),
    .Y(_02487_));
 sg13g2_nand3_1 _22835_ (.B(_02441_),
    .C(_02442_),
    .A(_02454_),
    .Y(_02488_));
 sg13g2_a21oi_1 _22836_ (.A1(_02488_),
    .A2(_05821_),
    .Y(_02489_),
    .B1(_02430_));
 sg13g2_nor2b_1 _22837_ (.A(_02478_),
    .B_N(_02489_),
    .Y(_02490_));
 sg13g2_inv_1 _22838_ (.Y(_02491_),
    .A(_05219_));
 sg13g2_nor2_1 _22839_ (.A(_05218_),
    .B(_05217_),
    .Y(_02493_));
 sg13g2_o21ai_1 _22840_ (.B1(_02473_),
    .Y(_02494_),
    .A1(_02491_),
    .A2(_02493_));
 sg13g2_o21ai_1 _22841_ (.B1(_02494_),
    .Y(_02495_),
    .A1(net72),
    .A2(_02490_));
 sg13g2_nand2_1 _22842_ (.Y(_02496_),
    .A(_02495_),
    .B(_02418_));
 sg13g2_nor2_1 _22843_ (.A(_02406_),
    .B(_02411_),
    .Y(_02497_));
 sg13g2_inv_1 _22844_ (.Y(_02498_),
    .A(_02497_));
 sg13g2_a22oi_1 _22845_ (.Y(_02499_),
    .B1(_02482_),
    .B2(_02485_),
    .A2(_02498_),
    .A1(_02496_));
 sg13g2_o21ai_1 _22846_ (.B1(_02499_),
    .Y(_02500_),
    .A1(_02486_),
    .A2(_02487_));
 sg13g2_inv_1 _22847_ (.Y(_02501_),
    .A(_02496_));
 sg13g2_nand2_1 _22848_ (.Y(_02502_),
    .A(_02497_),
    .B(_02501_));
 sg13g2_nand2_1 _22849_ (.Y(_02504_),
    .A(_02500_),
    .B(_02502_));
 sg13g2_mux2_1 _22850_ (.A0(_02417_),
    .A1(_02471_),
    .S(_02504_),
    .X(_02505_));
 sg13g2_inv_1 _22851_ (.Y(_02506_),
    .A(_02260_));
 sg13g2_nand3_1 _22852_ (.B(net68),
    .C(_06254_),
    .A(_02506_),
    .Y(_02507_));
 sg13g2_nand2_1 _22853_ (.Y(_02508_),
    .A(_02507_),
    .B(_02256_));
 sg13g2_nand2_1 _22854_ (.Y(_02509_),
    .A(_02256_),
    .B(_06259_));
 sg13g2_nand2_1 _22855_ (.Y(_02510_),
    .A(_06270_),
    .B(_06258_));
 sg13g2_nand3_1 _22856_ (.B(_02509_),
    .C(_02510_),
    .A(_02508_),
    .Y(_02511_));
 sg13g2_nand2b_1 _22857_ (.Y(_02512_),
    .B(_06506_),
    .A_N(_02228_));
 sg13g2_nand2b_1 _22858_ (.Y(_02513_),
    .B(_02512_),
    .A_N(_02229_));
 sg13g2_nand2_1 _22859_ (.Y(_02515_),
    .A(_02513_),
    .B(net67));
 sg13g2_nand2_1 _22860_ (.Y(_02516_),
    .A(_02511_),
    .B(_02515_));
 sg13g2_nand2_1 _22861_ (.Y(_02517_),
    .A(_02516_),
    .B(_02202_));
 sg13g2_inv_1 _22862_ (.Y(_02518_),
    .A(_02517_));
 sg13g2_inv_1 _22863_ (.Y(_02519_),
    .A(_02482_));
 sg13g2_nor2_1 _22864_ (.A(_02484_),
    .B(_02504_),
    .Y(_02520_));
 sg13g2_a21o_1 _22865_ (.A2(_02504_),
    .A1(_02519_),
    .B1(_02520_),
    .X(_02521_));
 sg13g2_inv_1 _22866_ (.Y(_02522_),
    .A(_02521_));
 sg13g2_nor2b_1 _22867_ (.A(_02505_),
    .B_N(_02263_),
    .Y(_02523_));
 sg13g2_o21ai_1 _22868_ (.B1(_02523_),
    .Y(_02524_),
    .A1(_02518_),
    .A2(_02522_));
 sg13g2_nand3_1 _22869_ (.B(_11732_),
    .C(_01613_),
    .A(_02236_),
    .Y(_02525_));
 sg13g2_a21oi_1 _22870_ (.A1(_02525_),
    .A2(_05194_),
    .Y(_02526_),
    .B1(_02223_));
 sg13g2_nor2b_1 _22871_ (.A(_02513_),
    .B_N(_02526_),
    .Y(_02527_));
 sg13g2_nor2_1 _22872_ (.A(_05188_),
    .B(_06269_),
    .Y(_02528_));
 sg13g2_o21ai_1 _22873_ (.B1(_02508_),
    .Y(_02529_),
    .A1(_06271_),
    .A2(_02528_));
 sg13g2_o21ai_1 _22874_ (.B1(_02529_),
    .Y(_02530_),
    .A1(net63),
    .A2(_02527_));
 sg13g2_nand2_1 _22875_ (.Y(_02531_),
    .A(_02530_),
    .B(_02202_));
 sg13g2_nor2_1 _22876_ (.A(_02501_),
    .B(_02498_),
    .Y(_02532_));
 sg13g2_nand2b_1 _22877_ (.Y(_02533_),
    .B(_02532_),
    .A_N(_02531_));
 sg13g2_nand2_1 _22878_ (.Y(_02534_),
    .A(_02522_),
    .B(_02518_));
 sg13g2_nand3_1 _22879_ (.B(_02533_),
    .C(_02534_),
    .A(_02524_),
    .Y(_02536_));
 sg13g2_o21ai_1 _22880_ (.B1(_02531_),
    .Y(_02537_),
    .A1(_02501_),
    .A2(_02498_));
 sg13g2_nand2_2 _22881_ (.Y(_02538_),
    .A(_02536_),
    .B(_02537_));
 sg13g2_mux2_1 _22882_ (.A0(_02263_),
    .A1(_02505_),
    .S(_02538_),
    .X(_02539_));
 sg13g2_nor2_1 _22883_ (.A(_02517_),
    .B(_02538_),
    .Y(_02540_));
 sg13g2_a21o_1 _22884_ (.A2(_02538_),
    .A1(_02521_),
    .B1(_02540_),
    .X(_02541_));
 sg13g2_inv_1 _22885_ (.Y(_02542_),
    .A(_02541_));
 sg13g2_nand2_1 _22886_ (.Y(_02543_),
    .A(_02197_),
    .B(net97));
 sg13g2_nand2_1 _22887_ (.Y(_02544_),
    .A(_02543_),
    .B(_04992_));
 sg13g2_nand3_1 _22888_ (.B(net57),
    .C(_06784_),
    .A(_02193_),
    .Y(_02545_));
 sg13g2_a22oi_1 _22889_ (.Y(_02546_),
    .B1(_02545_),
    .B2(_02543_),
    .A2(_06761_),
    .A1(_04991_));
 sg13g2_nand4_1 _22890_ (.B(_04560_),
    .C(_04554_),
    .A(_02154_),
    .Y(_02547_),
    .D(_04555_));
 sg13g2_a21o_1 _22891_ (.A2(_02156_),
    .A1(_02547_),
    .B1(net63),
    .X(_02548_));
 sg13g2_inv_1 _22892_ (.Y(_02549_),
    .A(_02548_));
 sg13g2_a21o_1 _22893_ (.A2(_02546_),
    .A1(_02544_),
    .B1(_02549_),
    .X(_02550_));
 sg13g2_nand2_1 _22894_ (.Y(_02551_),
    .A(_02550_),
    .B(\b.gen_square[60].sq.mask ));
 sg13g2_inv_1 _22895_ (.Y(_02552_),
    .A(_02551_));
 sg13g2_nor2b_1 _22896_ (.A(_02539_),
    .B_N(_02201_),
    .Y(_02553_));
 sg13g2_o21ai_1 _22897_ (.B1(_02553_),
    .Y(_02554_),
    .A1(_02542_),
    .A2(_02552_));
 sg13g2_nor2_1 _22898_ (.A(net48),
    .B(_04561_),
    .Y(_02555_));
 sg13g2_nor2b_1 _22899_ (.A(_02189_),
    .B_N(_02183_),
    .Y(_02557_));
 sg13g2_o21ai_1 _22900_ (.B1(_02157_),
    .Y(_02558_),
    .A1(_02557_),
    .A2(_04558_));
 sg13g2_nand2_1 _22901_ (.Y(_02559_),
    .A(_02543_),
    .B(_02545_));
 sg13g2_xnor2_1 _22902_ (.Y(_02560_),
    .A(_04553_),
    .B(_06760_));
 sg13g2_a221oi_1 _22903_ (.B2(_02560_),
    .C1(_02549_),
    .B1(_02559_),
    .A1(_02555_),
    .Y(_02561_),
    .A2(_02558_));
 sg13g2_nor2_1 _22904_ (.A(_02136_),
    .B(_02561_),
    .Y(_02562_));
 sg13g2_nand3_1 _22905_ (.B(_02531_),
    .C(_02562_),
    .A(_02532_),
    .Y(_02563_));
 sg13g2_nand2_1 _22906_ (.Y(_02564_),
    .A(_02532_),
    .B(_02531_));
 sg13g2_nand2b_1 _22907_ (.Y(_02565_),
    .B(_02564_),
    .A_N(_02562_));
 sg13g2_nand2_1 _22908_ (.Y(_02566_),
    .A(_02542_),
    .B(_02552_));
 sg13g2_nand4_1 _22909_ (.B(_02563_),
    .C(_02565_),
    .A(_02554_),
    .Y(_02567_),
    .D(_02566_));
 sg13g2_nand2_2 _22910_ (.Y(_02568_),
    .A(_02567_),
    .B(_02565_));
 sg13g2_mux2_1 _22911_ (.A0(_02201_),
    .A1(_02539_),
    .S(_02568_),
    .X(_02569_));
 sg13g2_nor2_1 _22912_ (.A(_02562_),
    .B(_02564_),
    .Y(_02570_));
 sg13g2_nor2_1 _22913_ (.A(_04364_),
    .B(_04472_),
    .Y(_02571_));
 sg13g2_nand2_1 _22914_ (.Y(_02572_),
    .A(_04362_),
    .B(net41));
 sg13g2_o21ai_1 _22915_ (.B1(_02116_),
    .Y(_02573_),
    .A1(_02572_),
    .A2(_02131_));
 sg13g2_o21ai_1 _22916_ (.B1(_02573_),
    .Y(_02574_),
    .A1(_04474_),
    .A2(_02571_));
 sg13g2_nand2_1 _22917_ (.Y(_02575_),
    .A(_01260_),
    .B(_00833_));
 sg13g2_o21ai_1 _22918_ (.B1(_06633_),
    .Y(_02576_),
    .A1(_02575_),
    .A2(_02093_));
 sg13g2_o21ai_1 _22919_ (.B1(_02576_),
    .Y(_02578_),
    .A1(_04471_),
    .A2(_02121_));
 sg13g2_nand2b_1 _22920_ (.Y(_02579_),
    .B(_07152_),
    .A_N(_02125_));
 sg13g2_nand2b_1 _22921_ (.Y(_02580_),
    .B(_02579_),
    .A_N(_02126_));
 sg13g2_o21ai_1 _22922_ (.B1(net56),
    .Y(_02581_),
    .A1(_02578_),
    .A2(_02580_));
 sg13g2_nand2_1 _22923_ (.Y(_02582_),
    .A(_02574_),
    .B(_02581_));
 sg13g2_nand2_1 _22924_ (.Y(_02583_),
    .A(_02582_),
    .B(_02064_));
 sg13g2_inv_1 _22925_ (.Y(_02584_),
    .A(_02583_));
 sg13g2_nor2b_1 _22926_ (.A(_02569_),
    .B_N(_02135_),
    .Y(_02585_));
 sg13g2_nor2_1 _22927_ (.A(_02551_),
    .B(_02568_),
    .Y(_02586_));
 sg13g2_a21o_1 _22928_ (.A2(_02568_),
    .A1(_02541_),
    .B1(_02586_),
    .X(_02587_));
 sg13g2_buf_1 _22929_ (.A(_02587_),
    .X(_02588_));
 sg13g2_nand2_1 _22930_ (.Y(_02589_),
    .A(_02116_),
    .B(_04378_));
 sg13g2_nand2_1 _22931_ (.Y(_02590_),
    .A(_04473_),
    .B(_04377_));
 sg13g2_nand3_1 _22932_ (.B(_02589_),
    .C(_02590_),
    .A(_02573_),
    .Y(_02591_));
 sg13g2_nand2_1 _22933_ (.Y(_02592_),
    .A(_02580_),
    .B(net56));
 sg13g2_nand2_1 _22934_ (.Y(_02593_),
    .A(_02591_),
    .B(_02592_));
 sg13g2_nand2_1 _22935_ (.Y(_02594_),
    .A(_02593_),
    .B(_02064_));
 sg13g2_nand2_1 _22936_ (.Y(_02595_),
    .A(_02588_),
    .B(_02594_));
 sg13g2_nand2_1 _22937_ (.Y(_02596_),
    .A(_02570_),
    .B(_02584_));
 sg13g2_o21ai_1 _22938_ (.B1(_02596_),
    .Y(_02597_),
    .A1(_02594_),
    .A2(_02588_));
 sg13g2_a21o_1 _22939_ (.A2(_02595_),
    .A1(_02585_),
    .B1(_02597_),
    .X(_02599_));
 sg13g2_o21ai_1 _22940_ (.B1(_02599_),
    .Y(_02600_),
    .A1(_02570_),
    .A2(_02584_));
 sg13g2_buf_1 _22941_ (.A(_02600_),
    .X(_02601_));
 sg13g2_mux2_1 _22942_ (.A0(_02135_),
    .A1(_02569_),
    .S(_02601_),
    .X(_02602_));
 sg13g2_inv_1 _22943_ (.Y(_02603_),
    .A(\b.gen_square[62].sq.mask ));
 sg13g2_inv_1 _22944_ (.Y(_02604_),
    .A(_04252_));
 sg13g2_a21oi_1 _22945_ (.A1(_02604_),
    .A2(_05727_),
    .Y(_02605_),
    .B1(_05728_));
 sg13g2_inv_1 _22946_ (.Y(_02606_),
    .A(_02605_));
 sg13g2_a21oi_1 _22947_ (.A1(_04335_),
    .A2(_05727_),
    .Y(_02607_),
    .B1(_05744_));
 sg13g2_a221oi_1 _22948_ (.B2(_02607_),
    .C1(_07559_),
    .B1(_02606_),
    .A1(_02032_),
    .Y(_02608_),
    .A2(_02015_));
 sg13g2_nor2_1 _22949_ (.A(_07241_),
    .B(_02173_),
    .Y(_02610_));
 sg13g2_a21oi_1 _22950_ (.A1(_07765_),
    .A2(_04435_),
    .Y(_02611_),
    .B1(_04441_));
 sg13g2_nor4_1 _22951_ (.A(_06625_),
    .B(_02611_),
    .C(_07250_),
    .D(_07735_),
    .Y(_02612_));
 sg13g2_inv_1 _22952_ (.Y(_02613_),
    .A(_08394_));
 sg13g2_a21oi_1 _22953_ (.A1(_07187_),
    .A2(_04724_),
    .Y(_02614_),
    .B1(_02613_));
 sg13g2_o21ai_1 _22954_ (.B1(_08388_),
    .Y(_02615_),
    .A1(_04726_),
    .A2(_07209_));
 sg13g2_nand2_1 _22955_ (.Y(_02616_),
    .A(_02615_),
    .B(_04990_));
 sg13g2_a22oi_1 _22956_ (.Y(_02617_),
    .B1(_02614_),
    .B2(_02616_),
    .A2(_04431_),
    .A1(_04426_));
 sg13g2_nand4_1 _22957_ (.B(_02610_),
    .C(_02612_),
    .A(_02608_),
    .Y(_02618_),
    .D(_02617_));
 sg13g2_nand2b_1 _22958_ (.Y(_02619_),
    .B(_02616_),
    .A_N(_02614_));
 sg13g2_nor2_1 _22959_ (.A(_07830_),
    .B(_00938_),
    .Y(_02621_));
 sg13g2_nand2b_1 _22960_ (.Y(_02622_),
    .B(_02621_),
    .A_N(_01207_));
 sg13g2_nor4_1 _22961_ (.A(_07619_),
    .B(_05005_),
    .C(_02169_),
    .D(_02622_),
    .Y(_02623_));
 sg13g2_nand3_1 _22962_ (.B(_02103_),
    .C(_02623_),
    .A(_02619_),
    .Y(_02624_));
 sg13g2_a22oi_1 _22963_ (.Y(_02625_),
    .B1(_02605_),
    .B2(_02607_),
    .A2(_02015_),
    .A1(_02031_));
 sg13g2_inv_1 _22964_ (.Y(_02626_),
    .A(_02625_));
 sg13g2_nor2_1 _22965_ (.A(_02624_),
    .B(_02626_),
    .Y(_02627_));
 sg13g2_nand2b_1 _22966_ (.Y(_02628_),
    .B(_02627_),
    .A_N(_02618_));
 sg13g2_nand2b_1 _22967_ (.Y(_02629_),
    .B(_04451_),
    .A_N(_04462_));
 sg13g2_and3_1 _22968_ (.X(_02630_),
    .A(_02628_),
    .B(_05092_),
    .C(_02629_));
 sg13g2_o21ai_1 _22969_ (.B1(_02630_),
    .Y(_02632_),
    .A1(_07211_),
    .A2(_04462_));
 sg13g2_a21oi_1 _22970_ (.A1(_02615_),
    .A2(_07765_),
    .Y(_02633_),
    .B1(_04452_));
 sg13g2_nor2_1 _22971_ (.A(_07617_),
    .B(_02626_),
    .Y(_02634_));
 sg13g2_a21oi_1 _22972_ (.A1(_02608_),
    .A2(_02634_),
    .Y(_02635_),
    .B1(_04452_));
 sg13g2_inv_1 _22973_ (.Y(_02636_),
    .A(_04492_));
 sg13g2_o21ai_1 _22974_ (.B1(_02636_),
    .Y(_02637_),
    .A1(_02633_),
    .A2(_02635_));
 sg13g2_nand2b_1 _22975_ (.Y(_02638_),
    .B(_02633_),
    .A_N(_07212_));
 sg13g2_nand3_1 _22976_ (.B(_04448_),
    .C(_02638_),
    .A(_02637_),
    .Y(_02639_));
 sg13g2_nor3_1 _22977_ (.A(_04989_),
    .B(_01851_),
    .C(_07654_),
    .Y(_02640_));
 sg13g2_nand4_1 _22978_ (.B(_04449_),
    .C(_04376_),
    .A(_02640_),
    .Y(_02641_),
    .D(_07149_));
 sg13g2_nor2_1 _22979_ (.A(net48),
    .B(_04455_),
    .Y(_02643_));
 sg13g2_nand3_1 _22980_ (.B(_02641_),
    .C(_02643_),
    .A(_02639_),
    .Y(_02644_));
 sg13g2_nand3b_1 _22981_ (.B(_02618_),
    .C(_04452_),
    .Y(_02645_),
    .A_N(_02627_));
 sg13g2_nor2_1 _22982_ (.A(net192),
    .B(_02645_),
    .Y(_02646_));
 sg13g2_nand2_1 _22983_ (.Y(_02647_),
    .A(_02646_),
    .B(_07211_));
 sg13g2_nand3_1 _22984_ (.B(_02644_),
    .C(_02647_),
    .A(_02632_),
    .Y(_02648_));
 sg13g2_nor2b_1 _22985_ (.A(_02603_),
    .B_N(_02648_),
    .Y(_02649_));
 sg13g2_inv_1 _22986_ (.Y(_02650_),
    .A(_02570_));
 sg13g2_nor2_1 _22987_ (.A(_02584_),
    .B(_02650_),
    .Y(_02651_));
 sg13g2_inv_1 _22988_ (.Y(_02652_),
    .A(_02651_));
 sg13g2_nand3_1 _22989_ (.B(_05092_),
    .C(_04452_),
    .A(_02628_),
    .Y(_02654_));
 sg13g2_inv_1 _22990_ (.Y(_02655_),
    .A(_02646_));
 sg13g2_nand2_1 _22991_ (.Y(_02656_),
    .A(_02654_),
    .B(_02655_));
 sg13g2_xnor2_1 _22992_ (.Y(_02657_),
    .A(_04445_),
    .B(_04491_));
 sg13g2_nor2_1 _22993_ (.A(_07735_),
    .B(_00905_),
    .Y(_02658_));
 sg13g2_a21o_1 _22994_ (.A2(_02658_),
    .A1(_02621_),
    .B1(_06897_),
    .X(_02659_));
 sg13g2_nand2_1 _22995_ (.Y(_02660_),
    .A(_04448_),
    .B(net56));
 sg13g2_a21oi_1 _22996_ (.A1(_02638_),
    .A2(_02659_),
    .Y(_02661_),
    .B1(_02660_));
 sg13g2_a21oi_1 _22997_ (.A1(_02656_),
    .A2(_02657_),
    .Y(_02662_),
    .B1(_02661_));
 sg13g2_nand4_1 _22998_ (.B(_04460_),
    .C(_04443_),
    .A(_02635_),
    .Y(_02663_),
    .D(_04446_));
 sg13g2_a21o_1 _22999_ (.A2(_02637_),
    .A1(_02663_),
    .B1(_02660_),
    .X(_02665_));
 sg13g2_a21o_1 _23000_ (.A2(_02665_),
    .A1(_02662_),
    .B1(_02603_),
    .X(_02666_));
 sg13g2_buf_1 _23001_ (.A(_02666_),
    .X(_02667_));
 sg13g2_nand2_1 _23002_ (.Y(_02668_),
    .A(_02601_),
    .B(_02588_));
 sg13g2_o21ai_1 _23003_ (.B1(_02668_),
    .Y(_02669_),
    .A1(_02594_),
    .A2(_02601_));
 sg13g2_inv_1 _23004_ (.Y(_02670_),
    .A(_02669_));
 sg13g2_nand2_1 _23005_ (.Y(_02671_),
    .A(_02655_),
    .B(_04462_));
 sg13g2_nand2b_1 _23006_ (.Y(_02672_),
    .B(_04461_),
    .A_N(_04491_));
 sg13g2_nand3_1 _23007_ (.B(_02671_),
    .C(_02672_),
    .A(_02656_),
    .Y(_02673_));
 sg13g2_a21o_1 _23008_ (.A2(_02665_),
    .A1(_02673_),
    .B1(_02603_),
    .X(_02674_));
 sg13g2_inv_1 _23009_ (.Y(_02676_),
    .A(_02674_));
 sg13g2_nor2_1 _23010_ (.A(_02667_),
    .B(_02652_),
    .Y(_02677_));
 sg13g2_a21oi_1 _23011_ (.A1(_02670_),
    .A2(_02676_),
    .Y(_02678_),
    .B1(_02677_));
 sg13g2_nor2b_1 _23012_ (.A(_02602_),
    .B_N(_02649_),
    .Y(_02679_));
 sg13g2_o21ai_1 _23013_ (.B1(_02679_),
    .Y(_02680_),
    .A1(_02670_),
    .A2(_02676_));
 sg13g2_a22oi_1 _23014_ (.Y(_02681_),
    .B1(_02678_),
    .B2(_02680_),
    .A2(_02667_),
    .A1(_02652_));
 sg13g2_buf_1 _23015_ (.A(_02681_),
    .X(_02682_));
 sg13g2_mux2_1 _23016_ (.A0(_02602_),
    .A1(_02649_),
    .S(_02682_),
    .X(_02683_));
 sg13g2_nand2_1 _23017_ (.Y(_02684_),
    .A(_02053_),
    .B(net97));
 sg13g2_a22oi_1 _23018_ (.Y(_02685_),
    .B1(_04423_),
    .B2(_02684_),
    .A2(_04422_),
    .A1(_04500_));
 sg13g2_nand3_1 _23019_ (.B(net41),
    .C(_04427_),
    .A(_02058_),
    .Y(_02686_));
 sg13g2_nand2_1 _23020_ (.Y(_02687_),
    .A(_02684_),
    .B(_02686_));
 sg13g2_nand2_1 _23021_ (.Y(_02688_),
    .A(_02685_),
    .B(_02687_));
 sg13g2_nand4_1 _23022_ (.B(_04421_),
    .C(_04410_),
    .A(_02039_),
    .Y(_02689_),
    .D(_04413_));
 sg13g2_nand2_1 _23023_ (.Y(_02690_),
    .A(_04415_),
    .B(net56));
 sg13g2_a21o_1 _23024_ (.A2(_02040_),
    .A1(_02689_),
    .B1(_02690_),
    .X(_02691_));
 sg13g2_a21o_1 _23025_ (.A2(_02691_),
    .A1(_02688_),
    .B1(_02062_),
    .X(_02692_));
 sg13g2_inv_1 _23026_ (.Y(_02693_),
    .A(_02692_));
 sg13g2_nor2_1 _23027_ (.A(_02669_),
    .B(_02682_),
    .Y(_02694_));
 sg13g2_a21oi_1 _23028_ (.A1(_02674_),
    .A2(_02682_),
    .Y(_02695_),
    .B1(_02694_));
 sg13g2_inv_1 _23029_ (.Y(_02697_),
    .A(_02695_));
 sg13g2_nor2b_1 _23030_ (.A(_02683_),
    .B_N(_02063_),
    .Y(_02698_));
 sg13g2_o21ai_1 _23031_ (.B1(_02698_),
    .Y(_02699_),
    .A1(_02693_),
    .A2(_02697_));
 sg13g2_nand2_1 _23032_ (.Y(_02700_),
    .A(_02651_),
    .B(_02667_));
 sg13g2_nor2_1 _23033_ (.A(_04412_),
    .B(_04499_),
    .Y(_02701_));
 sg13g2_o21ai_1 _23034_ (.B1(_02687_),
    .Y(_02702_),
    .A1(_04501_),
    .A2(_02701_));
 sg13g2_o21ai_1 _23035_ (.B1(_07163_),
    .Y(_02703_),
    .A1(_07907_),
    .A2(_07932_));
 sg13g2_a21o_1 _23036_ (.A2(_02703_),
    .A1(_02041_),
    .B1(_02690_),
    .X(_02704_));
 sg13g2_nand3_1 _23037_ (.B(_02691_),
    .C(_02704_),
    .A(_02702_),
    .Y(_02705_));
 sg13g2_nand2_1 _23038_ (.Y(_02706_),
    .A(_02705_),
    .B(_02061_));
 sg13g2_nand2_1 _23039_ (.Y(_02707_),
    .A(_02700_),
    .B(_02706_));
 sg13g2_nand4_1 _23040_ (.B(_02061_),
    .C(_02667_),
    .A(_02651_),
    .Y(_02708_),
    .D(_02705_));
 sg13g2_nand2_1 _23041_ (.Y(_02709_),
    .A(_02697_),
    .B(_02693_));
 sg13g2_nand4_1 _23042_ (.B(_02707_),
    .C(_02708_),
    .A(_02699_),
    .Y(_02710_),
    .D(_02709_));
 sg13g2_nand2_1 _23043_ (.Y(_02711_),
    .A(_02710_),
    .B(_02707_));
 sg13g2_mux2_1 _23044_ (.A0(_02063_),
    .A1(_02683_),
    .S(_02711_),
    .X(_02712_));
 sg13g2_nor2b_1 _23045_ (.A(_01983_),
    .B_N(_02712_),
    .Y(_02713_));
 sg13g2_nand2_1 _23046_ (.Y(_02714_),
    .A(_01978_),
    .B(_01949_));
 sg13g2_nand3_1 _23047_ (.B(_01976_),
    .C(_07689_),
    .A(_01973_),
    .Y(_02715_));
 sg13g2_nor2_1 _23048_ (.A(_02692_),
    .B(_02711_),
    .Y(_02716_));
 sg13g2_a21oi_1 _23049_ (.A1(_02695_),
    .A2(_02711_),
    .Y(_02718_),
    .B1(_02716_));
 sg13g2_nand3_1 _23050_ (.B(_02715_),
    .C(_02718_),
    .A(_02714_),
    .Y(_02719_));
 sg13g2_nand2_1 _23051_ (.Y(_02720_),
    .A(_02713_),
    .B(_02719_));
 sg13g2_nand2_1 _23052_ (.Y(_02721_),
    .A(_02714_),
    .B(_02715_));
 sg13g2_nand2b_1 _23053_ (.Y(_02722_),
    .B(_02721_),
    .A_N(_02718_));
 sg13g2_nand2_1 _23054_ (.Y(_02723_),
    .A(_02720_),
    .B(_02722_));
 sg13g2_nor2b_1 _23055_ (.A(_02700_),
    .B_N(_02706_),
    .Y(_02724_));
 sg13g2_o21ai_1 _23056_ (.B1(_02724_),
    .Y(_02725_),
    .A1(_01960_),
    .A2(_01963_));
 sg13g2_nand2_1 _23057_ (.Y(_02726_),
    .A(_02723_),
    .B(_02725_));
 sg13g2_buf_8 _23058_ (.A(_02726_),
    .X(_02727_));
 sg13g2_nor2_1 _23059_ (.A(_01960_),
    .B(_01963_),
    .Y(_02728_));
 sg13g2_nand2b_1 _23060_ (.Y(_02729_),
    .B(_02728_),
    .A_N(_02724_));
 sg13g2_buf_8 _23061_ (.A(_02729_),
    .X(_02730_));
 sg13g2_nand2_1 _23062_ (.Y(_02731_),
    .A(_02727_),
    .B(_02730_));
 sg13g2_buf_8 _23063_ (.A(_02731_),
    .X(_02732_));
 sg13g2_inv_1 _23064_ (.Y(_02733_),
    .A(_02682_));
 sg13g2_inv_1 _23065_ (.Y(_02734_),
    .A(_02568_));
 sg13g2_inv_1 _23066_ (.Y(_02735_),
    .A(_02504_));
 sg13g2_inv_1 _23067_ (.Y(_02736_),
    .A(_02538_));
 sg13g2_a21oi_1 _23068_ (.A1(_02414_),
    .A2(_02735_),
    .Y(_02737_),
    .B1(_02736_));
 sg13g2_o21ai_1 _23069_ (.B1(_02601_),
    .Y(_02739_),
    .A1(_02734_),
    .A2(_02737_));
 sg13g2_a22oi_1 _23070_ (.Y(_02740_),
    .B1(_02707_),
    .B2(_02710_),
    .A2(_02739_),
    .A1(_02733_));
 sg13g2_nand2_1 _23071_ (.Y(_02741_),
    .A(_02732_),
    .B(_02740_));
 sg13g2_inv_2 _23072_ (.Y(_02742_),
    .A(_01154_));
 sg13g2_inv_2 _23073_ (.Y(_02743_),
    .A(_01123_));
 sg13g2_inv_1 _23074_ (.Y(_02744_),
    .A(_00784_));
 sg13g2_o21ai_1 _23075_ (.B1(_00687_),
    .Y(_02745_),
    .A1(_00634_),
    .A2(_00655_));
 sg13g2_a21o_1 _23076_ (.A2(_02745_),
    .A1(_02744_),
    .B1(_00896_),
    .X(_02746_));
 sg13g2_a22oi_1 _23077_ (.Y(_02747_),
    .B1(_01092_),
    .B2(_01091_),
    .A2(_02746_),
    .A1(_00999_));
 sg13g2_nand2_1 _23078_ (.Y(_02748_),
    .A(_10537_),
    .B(_10542_));
 sg13g2_inv_1 _23079_ (.Y(_02749_),
    .A(_10593_));
 sg13g2_a21oi_1 _23080_ (.A1(_02748_),
    .A2(_02749_),
    .Y(_02750_),
    .B1(_10693_));
 sg13g2_nand2b_1 _23081_ (.Y(_02751_),
    .B(_10731_),
    .A_N(_02750_));
 sg13g2_a21oi_1 _23082_ (.A1(_10768_),
    .A2(_02751_),
    .Y(_02752_),
    .B1(_10865_));
 sg13g2_nand2b_1 _23083_ (.Y(_02753_),
    .B(_10943_),
    .A_N(_02752_));
 sg13g2_nor2_1 _23084_ (.A(_09528_),
    .B(_09666_),
    .Y(_02754_));
 sg13g2_o21ai_1 _23085_ (.B1(_09923_),
    .Y(_02755_),
    .A1(_09806_),
    .A2(_02754_));
 sg13g2_nand2_1 _23086_ (.Y(_02756_),
    .A(_09962_),
    .B(_02755_));
 sg13g2_nand2_1 _23087_ (.Y(_02757_),
    .A(_09999_),
    .B(_02756_));
 sg13g2_a21oi_1 _23088_ (.A1(_10102_),
    .A2(_02757_),
    .Y(_02758_),
    .B1(_10970_));
 sg13g2_a21oi_1 _23089_ (.A1(_10970_),
    .A2(_02753_),
    .Y(_02760_),
    .B1(_02758_));
 sg13g2_inv_1 _23090_ (.Y(_02761_),
    .A(_11611_));
 sg13g2_inv_1 _23091_ (.Y(_02762_),
    .A(_11490_));
 sg13g2_inv_1 _23092_ (.Y(_02763_),
    .A(_11306_));
 sg13g2_o21ai_1 _23093_ (.B1(_11397_),
    .Y(_02764_),
    .A1(_11271_),
    .A2(_02763_));
 sg13g2_a22oi_1 _23094_ (.Y(_02765_),
    .B1(_11573_),
    .B2(_11572_),
    .A2(_02764_),
    .A1(_02762_));
 sg13g2_o21ai_1 _23095_ (.B1(_11699_),
    .Y(_02766_),
    .A1(_02761_),
    .A2(_02765_));
 sg13g2_nand2_1 _23096_ (.Y(_02767_),
    .A(_11727_),
    .B(_02766_));
 sg13g2_o21ai_1 _23097_ (.B1(_02767_),
    .Y(_02768_),
    .A1(_11727_),
    .A2(_02760_));
 sg13g2_nand2_1 _23098_ (.Y(_02769_),
    .A(_02743_),
    .B(_02768_));
 sg13g2_o21ai_1 _23099_ (.B1(_02769_),
    .Y(_02771_),
    .A1(_02743_),
    .A2(_02747_));
 sg13g2_a22oi_1 _23100_ (.Y(_02772_),
    .B1(_08593_),
    .B2(_08592_),
    .A2(_08566_),
    .A1(_08536_));
 sg13g2_inv_1 _23101_ (.Y(_02773_),
    .A(_08644_));
 sg13g2_o21ai_1 _23102_ (.B1(_02773_),
    .Y(_02774_),
    .A1(_08627_),
    .A2(_02772_));
 sg13g2_a22oi_1 _23103_ (.Y(_02775_),
    .B1(_08897_),
    .B2(_08896_),
    .A2(_02774_),
    .A1(_08788_));
 sg13g2_nor2_1 _23104_ (.A(_02775_),
    .B(_02742_),
    .Y(_02776_));
 sg13g2_a21oi_1 _23105_ (.A1(_02742_),
    .A2(_02771_),
    .Y(_02777_),
    .B1(_02776_));
 sg13g2_nor2_1 _23106_ (.A(_01483_),
    .B(_01575_),
    .Y(_02778_));
 sg13g2_nor2_1 _23107_ (.A(_02778_),
    .B(_01668_),
    .Y(_02779_));
 sg13g2_inv_1 _23108_ (.Y(_02780_),
    .A(_01785_));
 sg13g2_o21ai_1 _23109_ (.B1(_02780_),
    .Y(_02782_),
    .A1(_01751_),
    .A2(_02779_));
 sg13g2_a21oi_1 _23110_ (.A1(_01821_),
    .A2(_02782_),
    .Y(_02783_),
    .B1(_01914_));
 sg13g2_nand2b_1 _23111_ (.Y(_02784_),
    .B(net13),
    .A_N(_02783_));
 sg13g2_o21ai_1 _23112_ (.B1(_02784_),
    .Y(_02785_),
    .A1(net13),
    .A2(_02777_));
 sg13g2_inv_1 _23113_ (.Y(_02786_),
    .A(_07445_));
 sg13g2_inv_1 _23114_ (.Y(_02787_),
    .A(_07360_));
 sg13g2_a21oi_1 _23115_ (.A1(_02787_),
    .A2(_07393_),
    .Y(_02788_),
    .B1(_07424_));
 sg13g2_o21ai_1 _23116_ (.B1(_07466_),
    .Y(_02789_),
    .A1(_02786_),
    .A2(_02788_));
 sg13g2_nand2b_1 _23117_ (.Y(_02790_),
    .B(_02789_),
    .A_N(_07486_));
 sg13g2_a21oi_1 _23118_ (.A1(_07686_),
    .A2(_02790_),
    .Y(_02791_),
    .B1(net12));
 sg13g2_a21oi_1 _23119_ (.A1(net12),
    .A2(_02785_),
    .Y(_02793_),
    .B1(_02791_));
 sg13g2_nand3_1 _23120_ (.B(_02730_),
    .C(_02793_),
    .A(_02727_),
    .Y(_02794_));
 sg13g2_nand2_1 _23121_ (.Y(_02795_),
    .A(_02741_),
    .B(_02794_));
 sg13g2_nor2_1 _23122_ (.A(\state[10] ),
    .B(\state[2] ),
    .Y(_02796_));
 sg13g2_inv_1 _23123_ (.Y(_02797_),
    .A(_02796_));
 sg13g2_buf_1 _23124_ (.A(_02797_),
    .X(_02798_));
 sg13g2_nor2_2 _23125_ (.A(_02798_),
    .B(_01198_),
    .Y(_02799_));
 sg13g2_inv_4 _23126_ (.A(_02799_),
    .Y(_02800_));
 sg13g2_nand2_1 _23127_ (.Y(_02801_),
    .A(_02795_),
    .B(_02800_));
 sg13g2_nand3_1 _23128_ (.B(_02796_),
    .C(_01535_),
    .A(_01449_),
    .Y(_02802_));
 sg13g2_buf_1 _23129_ (.A(_02802_),
    .X(_02804_));
 sg13g2_inv_2 _23130_ (.Y(_02805_),
    .A(_02804_));
 sg13g2_inv_2 _23131_ (.Y(_02806_),
    .A(_11727_));
 sg13g2_nand2_1 _23132_ (.Y(_02807_),
    .A(_02743_),
    .B(_02806_));
 sg13g2_nor2_1 _23133_ (.A(_01154_),
    .B(net13),
    .Y(_02808_));
 sg13g2_a22oi_1 _23134_ (.Y(_02809_),
    .B1(_01976_),
    .B2(_01973_),
    .A2(_02808_),
    .A1(_02807_));
 sg13g2_nand3_1 _23135_ (.B(_02730_),
    .C(_02809_),
    .A(_02727_),
    .Y(_02810_));
 sg13g2_nor2_1 _23136_ (.A(_02800_),
    .B(_02810_),
    .Y(_02811_));
 sg13g2_nor2_1 _23137_ (.A(_02805_),
    .B(_02811_),
    .Y(_02812_));
 sg13g2_nand2_1 _23138_ (.Y(_02813_),
    .A(_02801_),
    .B(_02812_));
 sg13g2_nand2_1 _23139_ (.Y(_02815_),
    .A(_02805_),
    .B(\data_out[0] ));
 sg13g2_nand2_1 _23140_ (.Y(_00598_),
    .A(_02813_),
    .B(_02815_));
 sg13g2_nand2_1 _23141_ (.Y(_02816_),
    .A(net12),
    .B(_02808_));
 sg13g2_nor3_1 _23142_ (.A(_02800_),
    .B(_02816_),
    .C(_02732_),
    .Y(_02817_));
 sg13g2_nor2_1 _23143_ (.A(_02805_),
    .B(_02817_),
    .Y(_02818_));
 sg13g2_nand2_1 _23144_ (.Y(_02819_),
    .A(_02601_),
    .B(_02568_));
 sg13g2_a21oi_1 _23145_ (.A1(_02735_),
    .A2(_02538_),
    .Y(_02820_),
    .B1(_02819_));
 sg13g2_nand2_1 _23146_ (.Y(_02821_),
    .A(_02711_),
    .B(_02733_));
 sg13g2_nor2_1 _23147_ (.A(_02820_),
    .B(_02821_),
    .Y(_02822_));
 sg13g2_nand2_1 _23148_ (.Y(_02823_),
    .A(_02732_),
    .B(_02822_));
 sg13g2_nand3_1 _23149_ (.B(_10692_),
    .C(_02749_),
    .A(_10690_),
    .Y(_02825_));
 sg13g2_nand2_1 _23150_ (.Y(_02826_),
    .A(_10768_),
    .B(_10731_));
 sg13g2_inv_1 _23151_ (.Y(_02827_),
    .A(_02826_));
 sg13g2_a21oi_1 _23152_ (.A1(_02825_),
    .A2(_02827_),
    .Y(_02828_),
    .B1(_10865_));
 sg13g2_a22oi_1 _23153_ (.Y(_02829_),
    .B1(_10968_),
    .B2(_10967_),
    .A2(_02828_),
    .A1(_10943_));
 sg13g2_a22oi_1 _23154_ (.Y(_02830_),
    .B1(_09960_),
    .B2(_09959_),
    .A2(_09921_),
    .A1(_09922_));
 sg13g2_o21ai_1 _23155_ (.B1(_02830_),
    .Y(_02831_),
    .A1(_09666_),
    .A2(_09806_));
 sg13g2_nand3_1 _23156_ (.B(_09999_),
    .C(_02831_),
    .A(_10102_),
    .Y(_02832_));
 sg13g2_nor2b_1 _23157_ (.A(_10970_),
    .B_N(_02832_),
    .Y(_02833_));
 sg13g2_o21ai_1 _23158_ (.B1(_02806_),
    .Y(_02834_),
    .A1(_02829_),
    .A2(_02833_));
 sg13g2_nand2_1 _23159_ (.Y(_02836_),
    .A(_11574_),
    .B(_02762_));
 sg13g2_a21oi_1 _23160_ (.A1(_11306_),
    .A2(_11397_),
    .Y(_02837_),
    .B1(_02836_));
 sg13g2_nand2_1 _23161_ (.Y(_02838_),
    .A(_11699_),
    .B(_11611_));
 sg13g2_o21ai_1 _23162_ (.B1(_11727_),
    .Y(_02839_),
    .A1(_02837_),
    .A2(_02838_));
 sg13g2_a21oi_1 _23163_ (.A1(_02834_),
    .A2(_02839_),
    .Y(_02840_),
    .B1(_01123_));
 sg13g2_inv_1 _23164_ (.Y(_02841_),
    .A(_00655_));
 sg13g2_nand3_1 _23165_ (.B(_02744_),
    .C(_00890_),
    .A(_00887_),
    .Y(_02842_));
 sg13g2_a21oi_1 _23166_ (.A1(_02841_),
    .A2(_00687_),
    .Y(_02843_),
    .B1(_02842_));
 sg13g2_nand2_1 _23167_ (.Y(_02844_),
    .A(_01093_),
    .B(_00999_));
 sg13g2_nor2_1 _23168_ (.A(_02843_),
    .B(_02844_),
    .Y(_02845_));
 sg13g2_nor2_1 _23169_ (.A(_02845_),
    .B(_02743_),
    .Y(_02847_));
 sg13g2_o21ai_1 _23170_ (.B1(_02742_),
    .Y(_02848_),
    .A1(_02840_),
    .A2(_02847_));
 sg13g2_nand2_1 _23171_ (.Y(_02849_),
    .A(_02773_),
    .B(_08622_));
 sg13g2_a21oi_1 _23172_ (.A1(_08566_),
    .A2(_08594_),
    .Y(_02850_),
    .B1(_02849_));
 sg13g2_nand2_1 _23173_ (.Y(_02851_),
    .A(_08898_),
    .B(_08788_));
 sg13g2_o21ai_1 _23174_ (.B1(_01154_),
    .Y(_02852_),
    .A1(_02850_),
    .A2(_02851_));
 sg13g2_a21oi_1 _23175_ (.A1(_02848_),
    .A2(_02852_),
    .Y(_02853_),
    .B1(net13));
 sg13g2_nor2_1 _23176_ (.A(_01575_),
    .B(_01668_),
    .Y(_02854_));
 sg13g2_nand2b_1 _23177_ (.Y(_02855_),
    .B(_02780_),
    .A_N(_01751_));
 sg13g2_nor2_1 _23178_ (.A(_02854_),
    .B(_02855_),
    .Y(_02856_));
 sg13g2_nand3_1 _23179_ (.B(_01821_),
    .C(_01912_),
    .A(_01910_),
    .Y(_02858_));
 sg13g2_o21ai_1 _23180_ (.B1(net13),
    .Y(_02859_),
    .A1(_02856_),
    .A2(_02858_));
 sg13g2_nand2b_1 _23181_ (.Y(_02860_),
    .B(_02859_),
    .A_N(_02853_));
 sg13g2_inv_1 _23182_ (.Y(_02861_),
    .A(_07393_));
 sg13g2_a21oi_1 _23183_ (.A1(_07465_),
    .A2(_07462_),
    .Y(_02862_),
    .B1(_02786_));
 sg13g2_o21ai_1 _23184_ (.B1(_02862_),
    .Y(_02863_),
    .A1(_02861_),
    .A2(_07424_));
 sg13g2_a21oi_1 _23185_ (.A1(_07683_),
    .A2(_07685_),
    .Y(_02864_),
    .B1(_07486_));
 sg13g2_a21oi_1 _23186_ (.A1(_02863_),
    .A2(_02864_),
    .Y(_02865_),
    .B1(net12));
 sg13g2_a21oi_1 _23187_ (.A1(net12),
    .A2(_02860_),
    .Y(_02866_),
    .B1(_02865_));
 sg13g2_nand3_1 _23188_ (.B(_02730_),
    .C(_02866_),
    .A(_02727_),
    .Y(_02867_));
 sg13g2_nand2_1 _23189_ (.Y(_02868_),
    .A(_02823_),
    .B(_02867_));
 sg13g2_nand2_1 _23190_ (.Y(_02869_),
    .A(_02868_),
    .B(_02800_));
 sg13g2_nand2_1 _23191_ (.Y(_02870_),
    .A(_02818_),
    .B(_02869_));
 sg13g2_nand2_1 _23192_ (.Y(_02871_),
    .A(_02805_),
    .B(\data_out[1] ));
 sg13g2_nand2_1 _23193_ (.Y(_00599_),
    .A(_02870_),
    .B(_02871_));
 sg13g2_nand4_1 _23194_ (.B(_02728_),
    .C(_01981_),
    .A(_02721_),
    .Y(_02872_),
    .D(_01982_));
 sg13g2_nor3_1 _23195_ (.A(_02800_),
    .B(_02872_),
    .C(_02732_),
    .Y(_02873_));
 sg13g2_nor2_1 _23196_ (.A(_02805_),
    .B(_02873_),
    .Y(_02874_));
 sg13g2_nor2_1 _23197_ (.A(_02819_),
    .B(_02821_),
    .Y(_02875_));
 sg13g2_nand2_1 _23198_ (.Y(_02876_),
    .A(_02732_),
    .B(_02875_));
 sg13g2_nand3_1 _23199_ (.B(_09999_),
    .C(_02830_),
    .A(_10102_),
    .Y(_02878_));
 sg13g2_nand4_1 _23200_ (.B(_10861_),
    .C(_10857_),
    .A(_10943_),
    .Y(_02879_),
    .D(_02827_));
 sg13g2_mux2_1 _23201_ (.A0(_02878_),
    .A1(_02879_),
    .S(_10970_),
    .X(_02880_));
 sg13g2_nand2_1 _23202_ (.Y(_02881_),
    .A(_02806_),
    .B(_02880_));
 sg13g2_o21ai_1 _23203_ (.B1(_11727_),
    .Y(_02882_),
    .A1(_02836_),
    .A2(_02838_));
 sg13g2_a21oi_1 _23204_ (.A1(_02881_),
    .A2(_02882_),
    .Y(_02883_),
    .B1(_01123_));
 sg13g2_nor2_1 _23205_ (.A(_02842_),
    .B(_02844_),
    .Y(_02884_));
 sg13g2_nor2_1 _23206_ (.A(_02884_),
    .B(_02743_),
    .Y(_02885_));
 sg13g2_o21ai_1 _23207_ (.B1(_02742_),
    .Y(_02886_),
    .A1(_02883_),
    .A2(_02885_));
 sg13g2_o21ai_1 _23208_ (.B1(_01154_),
    .Y(_02887_),
    .A1(_02849_),
    .A2(_02851_));
 sg13g2_a21oi_1 _23209_ (.A1(_02886_),
    .A2(_02887_),
    .Y(_02888_),
    .B1(net13));
 sg13g2_o21ai_1 _23210_ (.B1(net13),
    .Y(_02889_),
    .A1(_02855_),
    .A2(_02858_));
 sg13g2_nand2b_1 _23211_ (.Y(_02890_),
    .B(_02889_),
    .A_N(_02888_));
 sg13g2_a21oi_1 _23212_ (.A1(_02862_),
    .A2(_02864_),
    .Y(_02891_),
    .B1(net12));
 sg13g2_a21oi_1 _23213_ (.A1(net12),
    .A2(_02890_),
    .Y(_02892_),
    .B1(_02891_));
 sg13g2_nand3_1 _23214_ (.B(_02730_),
    .C(_02892_),
    .A(_02727_),
    .Y(_02893_));
 sg13g2_nand3_1 _23215_ (.B(_02893_),
    .C(_02800_),
    .A(_02876_),
    .Y(_02894_));
 sg13g2_nor2_1 _23216_ (.A(\data_out[2] ),
    .B(_02804_),
    .Y(_02895_));
 sg13g2_a21oi_1 _23217_ (.A1(_02874_),
    .A2(_02894_),
    .Y(_00600_),
    .B1(_02895_));
 sg13g2_inv_1 _23218_ (.Y(_02896_),
    .A(\data_out[3] ));
 sg13g2_o21ai_1 _23219_ (.B1(_02743_),
    .Y(_02898_),
    .A1(_10970_),
    .A2(_11727_));
 sg13g2_a21oi_1 _23220_ (.A1(_02742_),
    .A2(_02898_),
    .Y(_02899_),
    .B1(_01944_));
 sg13g2_nand2b_1 _23221_ (.Y(_02900_),
    .B(net12),
    .A_N(_02899_));
 sg13g2_nand3_1 _23222_ (.B(_02730_),
    .C(_02900_),
    .A(_02727_),
    .Y(_02901_));
 sg13g2_nand3_1 _23223_ (.B(\b.gen_square[62].sq.mask ),
    .C(_04455_),
    .A(_02628_),
    .Y(_02902_));
 sg13g2_nand3_1 _23224_ (.B(_10067_),
    .C(_06159_),
    .A(_10050_),
    .Y(_02903_));
 sg13g2_nand3_1 _23225_ (.B(_10824_),
    .C(_04168_),
    .A(_10803_),
    .Y(_02904_));
 sg13g2_nand3_1 _23226_ (.B(_02903_),
    .C(_02904_),
    .A(_02902_),
    .Y(_02905_));
 sg13g2_nand3_1 _23227_ (.B(\b.gen_square[57].sq.mask ),
    .C(_05454_),
    .A(_02301_),
    .Y(_02906_));
 sg13g2_nand3_1 _23228_ (.B(_11875_),
    .C(_06050_),
    .A(_11924_),
    .Y(_02907_));
 sg13g2_nand3_1 _23229_ (.B(\b.gen_square[8].sq.mask ),
    .C(_05991_),
    .A(_09311_),
    .Y(_02908_));
 sg13g2_nand3_1 _23230_ (.B(_09046_),
    .C(_04190_),
    .A(_09027_),
    .Y(_02909_));
 sg13g2_nand4_1 _23231_ (.B(_02907_),
    .C(_02908_),
    .A(_02906_),
    .Y(_02910_),
    .D(_02909_));
 sg13g2_nand3_1 _23232_ (.B(_02202_),
    .C(_05197_),
    .A(_02506_),
    .Y(_02911_));
 sg13g2_nand3_1 _23233_ (.B(\b.gen_square[32].sq.mask ),
    .C(_05159_),
    .A(_08238_),
    .Y(_02912_));
 sg13g2_nand3_1 _23234_ (.B(_05120_),
    .C(_05041_),
    .A(_05081_),
    .Y(_02913_));
 sg13g2_nand3_1 _23235_ (.B(_09461_),
    .C(_04829_),
    .A(_09441_),
    .Y(_02914_));
 sg13g2_nand4_1 _23236_ (.B(_02912_),
    .C(_02913_),
    .A(_02911_),
    .Y(_02915_),
    .D(_02914_));
 sg13g2_nand3b_1 _23237_ (.B(_02064_),
    .C(_04372_),
    .Y(_02916_),
    .A_N(_02131_));
 sg13g2_nand3b_1 _23238_ (.B(_02418_),
    .C(_05227_),
    .Y(_02917_),
    .A_N(_02467_));
 sg13g2_nand4_1 _23239_ (.B(_11171_),
    .C(_06022_),
    .A(_11154_),
    .Y(_02919_),
    .D(_06024_));
 sg13g2_nand4_1 _23240_ (.B(_05808_),
    .C(_04621_),
    .A(_05797_),
    .Y(_02920_),
    .D(_04619_));
 sg13g2_nand4_1 _23241_ (.B(_02917_),
    .C(_02919_),
    .A(_02916_),
    .Y(_02921_),
    .D(_02920_));
 sg13g2_nand3_1 _23242_ (.B(_11452_),
    .C(_05858_),
    .A(_11440_),
    .Y(_02922_));
 sg13g2_nand3_1 _23243_ (.B(_01236_),
    .C(_04242_),
    .A(_01228_),
    .Y(_02923_));
 sg13g2_nand3_1 _23244_ (.B(_11365_),
    .C(_06574_),
    .A(_11359_),
    .Y(_02924_));
 sg13g2_nand3_1 _23245_ (.B(_11861_),
    .C(_06385_),
    .A(_11848_),
    .Y(_02925_));
 sg13g2_nand4_1 _23246_ (.B(_02923_),
    .C(_02924_),
    .A(_02922_),
    .Y(_02926_),
    .D(_02925_));
 sg13g2_nand3_1 _23247_ (.B(_07859_),
    .C(_04543_),
    .A(_07846_),
    .Y(_02927_));
 sg13g2_nand3_1 _23248_ (.B(_08150_),
    .C(_05140_),
    .A(_08131_),
    .Y(_02928_));
 sg13g2_nand3_1 _23249_ (.B(\b.gen_square[44].sq.mask ),
    .C(_04522_),
    .A(_01709_),
    .Y(_02929_));
 sg13g2_nand3_1 _23250_ (.B(_00851_),
    .C(_06178_),
    .A(_00843_),
    .Y(_02930_));
 sg13g2_nand4_1 _23251_ (.B(_02928_),
    .C(_02929_),
    .A(_02927_),
    .Y(_02931_),
    .D(_02930_));
 sg13g2_nor2_1 _23252_ (.A(_00674_),
    .B(_00661_),
    .Y(_02932_));
 sg13g2_nor2b_1 _23253_ (.A(_00742_),
    .B_N(_00749_),
    .Y(_02933_));
 sg13g2_a22oi_1 _23254_ (.Y(_02934_),
    .B1(_02933_),
    .B2(_00745_),
    .A2(_02932_),
    .A1(_11779_));
 sg13g2_nand3_1 _23255_ (.B(_01633_),
    .C(_05178_),
    .A(_01626_),
    .Y(_02935_));
 sg13g2_nand3_1 _23256_ (.B(\b.gen_square[36].sq.mask ),
    .C(_04922_),
    .A(_08001_),
    .Y(_02936_));
 sg13g2_nand3_1 _23257_ (.B(_08479_),
    .C(_05372_),
    .A(_08468_),
    .Y(_02937_));
 sg13g2_nand4_1 _23258_ (.B(_02935_),
    .C(_02936_),
    .A(_02934_),
    .Y(_02938_),
    .D(_02937_));
 sg13g2_or2_1 _23259_ (.X(_02940_),
    .B(_02938_),
    .A(_02931_));
 sg13g2_nor3_1 _23260_ (.A(_11296_),
    .B(_11080_),
    .C(_11106_),
    .Y(_02941_));
 sg13g2_nor3_1 _23261_ (.A(_01558_),
    .B(_01548_),
    .C(_01528_),
    .Y(_02942_));
 sg13g2_and3_1 _23262_ (.X(_02943_),
    .A(_11532_),
    .B(_11547_),
    .C(_05284_));
 sg13g2_nor3_1 _23263_ (.A(_07067_),
    .B(_07434_),
    .C(_07045_),
    .Y(_02944_));
 sg13g2_nor4_1 _23264_ (.A(_02941_),
    .B(_02942_),
    .C(_02943_),
    .D(_02944_),
    .Y(_02945_));
 sg13g2_nand3_1 _23265_ (.B(\b.gen_square[45].sq.mask ),
    .C(_04060_),
    .A(_01277_),
    .Y(_02946_));
 sg13g2_nand3_1 _23266_ (.B(_06852_),
    .C(_04669_),
    .A(_06844_),
    .Y(_02947_));
 sg13g2_nand3_1 _23267_ (.B(_00961_),
    .C(_04149_),
    .A(_00946_),
    .Y(_02948_));
 sg13g2_and3_1 _23268_ (.X(_02949_),
    .A(_02946_),
    .B(_02947_),
    .C(_02948_));
 sg13g2_nand2_1 _23269_ (.Y(_02951_),
    .A(_02945_),
    .B(_02949_));
 sg13g2_nor4_1 _23270_ (.A(_02921_),
    .B(_02926_),
    .C(_02940_),
    .D(_02951_),
    .Y(_02952_));
 sg13g2_and3_1 _23271_ (.X(_02953_),
    .A(_02058_),
    .B(_02061_),
    .C(_04417_));
 sg13g2_nand3_1 _23272_ (.B(_09890_),
    .C(_06949_),
    .A(_09874_),
    .Y(_02954_));
 sg13g2_nand3_1 _23273_ (.B(_08372_),
    .C(_05672_),
    .A(_08364_),
    .Y(_02955_));
 sg13g2_nand3_1 _23274_ (.B(\b.gen_square[41].sq.mask ),
    .C(_05558_),
    .A(_01363_),
    .Y(_02956_));
 sg13g2_nand3_1 _23275_ (.B(_09763_),
    .C(_06524_),
    .A(_09757_),
    .Y(_02957_));
 sg13g2_nand4_1 _23276_ (.B(_02955_),
    .C(_02956_),
    .A(_02954_),
    .Y(_02958_),
    .D(_02957_));
 sg13g2_nand3_1 _23277_ (.B(\b.gen_square[50].sq.mask ),
    .C(_04645_),
    .A(_06476_),
    .Y(_02959_));
 sg13g2_nand3_1 _23278_ (.B(_11042_),
    .C(_04212_),
    .A(_11035_),
    .Y(_02960_));
 sg13g2_nand3_1 _23279_ (.B(_11236_),
    .C(_05583_),
    .A(_11223_),
    .Y(_02962_));
 sg13g2_nand3_1 _23280_ (.B(_09169_),
    .C(_05885_),
    .A(_09162_),
    .Y(_02963_));
 sg13g2_nand4_1 _23281_ (.B(_02960_),
    .C(_02962_),
    .A(_02959_),
    .Y(_02964_),
    .D(_02963_));
 sg13g2_nand3b_1 _23282_ (.B(_08757_),
    .C(_04111_),
    .Y(_02965_),
    .A_N(_08744_));
 sg13g2_nand3_1 _23283_ (.B(_09632_),
    .C(_06328_),
    .A(_09617_),
    .Y(_02966_));
 sg13g2_nand3_1 _23284_ (.B(_07292_),
    .C(_04718_),
    .A(_07267_),
    .Y(_02967_));
 sg13g2_nand3_1 _23285_ (.B(_11980_),
    .C(_05641_),
    .A(_11971_),
    .Y(_02968_));
 sg13g2_nand4_1 _23286_ (.B(_02966_),
    .C(_02967_),
    .A(_02965_),
    .Y(_02969_),
    .D(_02968_));
 sg13g2_nor4_1 _23287_ (.A(_02953_),
    .B(_02958_),
    .C(_02964_),
    .D(_02969_),
    .Y(_02970_));
 sg13g2_nand2_1 _23288_ (.Y(_02971_),
    .A(_02952_),
    .B(_02970_));
 sg13g2_nor4_1 _23289_ (.A(_02905_),
    .B(_02910_),
    .C(_02915_),
    .D(_02971_),
    .Y(_02973_));
 sg13g2_nand3_1 _23290_ (.B(_11666_),
    .C(_06678_),
    .A(_11671_),
    .Y(_02974_));
 sg13g2_nand3_1 _23291_ (.B(\b.gen_square[60].sq.mask ),
    .C(_04563_),
    .A(_02193_),
    .Y(_02975_));
 sg13g2_nand3_1 _23292_ (.B(_10487_),
    .C(_05609_),
    .A(_10474_),
    .Y(_02976_));
 sg13g2_nand3_1 _23293_ (.B(_10428_),
    .C(_04854_),
    .A(_10398_),
    .Y(_02977_));
 sg13g2_nand4_1 _23294_ (.B(_02975_),
    .C(_02976_),
    .A(_02974_),
    .Y(_02978_),
    .D(_02977_));
 sg13g2_nand3_1 _23295_ (.B(_01058_),
    .C(_04082_),
    .A(_01066_),
    .Y(_02979_));
 sg13g2_nand3_1 _23296_ (.B(_08868_),
    .C(_04581_),
    .A(_08854_),
    .Y(_02980_));
 sg13g2_nand3_1 _23297_ (.B(_06147_),
    .C(_04601_),
    .A(_06137_),
    .Y(_02981_));
 sg13g2_nand3_1 _23298_ (.B(_07646_),
    .C(_07657_),
    .A(_07627_),
    .Y(_02982_));
 sg13g2_nand4_1 _23299_ (.B(_02980_),
    .C(_02981_),
    .A(_02979_),
    .Y(_02984_),
    .D(_02982_));
 sg13g2_nand3_1 _23300_ (.B(_10657_),
    .C(_06547_),
    .A(_10643_),
    .Y(_02985_));
 sg13g2_nand3_1 _23301_ (.B(_10190_),
    .C(_07089_),
    .A(_10739_),
    .Y(_02986_));
 sg13g2_nand3_1 _23302_ (.B(_10267_),
    .C(_06924_),
    .A(_10702_),
    .Y(_02987_));
 sg13g2_nand3_1 _23303_ (.B(\b.gen_square[47].sq.mask ),
    .C(_04395_),
    .A(_01866_),
    .Y(_02988_));
 sg13g2_nand4_1 _23304_ (.B(_02986_),
    .C(_02987_),
    .A(_02985_),
    .Y(_02989_),
    .D(_02988_));
 sg13g2_nand3_1 _23305_ (.B(_10913_),
    .C(_05306_),
    .A(_10904_),
    .Y(_02990_));
 sg13g2_nand3_1 _23306_ (.B(_01433_),
    .C(_05248_),
    .A(_01419_),
    .Y(_02991_));
 sg13g2_nand3_1 _23307_ (.B(\b.gen_square[2].sq.mask ),
    .C(_06343_),
    .A(_10335_),
    .Y(_02992_));
 sg13g2_nand3b_1 _23308_ (.B(_02362_),
    .C(_05267_),
    .Y(_02993_),
    .A_N(_02349_));
 sg13g2_nand4_1 _23309_ (.B(_02991_),
    .C(_02992_),
    .A(_02990_),
    .Y(_02995_),
    .D(_02993_));
 sg13g2_nor4_1 _23310_ (.A(_02978_),
    .B(_02984_),
    .C(_02989_),
    .D(_02995_),
    .Y(_02996_));
 sg13g2_a21o_1 _23311_ (.A2(_02996_),
    .A1(_02973_),
    .B1(net142),
    .X(_02997_));
 sg13g2_a21oi_1 _23312_ (.A1(_02997_),
    .A2(_02799_),
    .Y(_02998_),
    .B1(_02805_));
 sg13g2_o21ai_1 _23313_ (.B1(_02998_),
    .Y(_02999_),
    .A1(_02799_),
    .A2(_02901_));
 sg13g2_o21ai_1 _23314_ (.B1(_02999_),
    .Y(_00601_),
    .A1(_02896_),
    .A2(_02804_));
 sg13g2_buf_2 _23315_ (.A(\state[7] ),
    .X(_03000_));
 sg13g2_inv_1 _23316_ (.Y(_03001_),
    .A(_03000_));
 sg13g2_nand3_1 _23317_ (.B(_01406_),
    .C(data_out_valid),
    .A(_03001_),
    .Y(_03002_));
 sg13g2_nand2_1 _23318_ (.Y(_00602_),
    .A(_02805_),
    .B(_03002_));
 sg13g2_a21oi_1 _23319_ (.A1(_00273_),
    .A2(_00980_),
    .Y(_03004_),
    .B1(_00011_));
 sg13g2_nor2_1 _23320_ (.A(net2),
    .B(_03004_),
    .Y(_00603_));
 sg13g2_nand2_1 _23321_ (.Y(_03005_),
    .A(_00991_),
    .B(_01013_));
 sg13g2_buf_2 _23322_ (.A(_03005_),
    .X(_03006_));
 sg13g2_nor2_1 _23323_ (.A(\spi.sdi_r[0] ),
    .B(_03006_),
    .Y(_03007_));
 sg13g2_a21oi_1 _23324_ (.A1(_01155_),
    .A2(_03006_),
    .Y(_00604_),
    .B1(_03007_));
 sg13g2_nor2_1 _23325_ (.A(\spi.sdi_r[1] ),
    .B(_03006_),
    .Y(_03008_));
 sg13g2_a21oi_1 _23326_ (.A1(_01546_),
    .A2(_03006_),
    .Y(_00605_),
    .B1(_03008_));
 sg13g2_inv_1 _23327_ (.Y(_03009_),
    .A(_00893_));
 sg13g2_nor2_1 _23328_ (.A(\spi.sdi_r[2] ),
    .B(_03006_),
    .Y(_03010_));
 sg13g2_a21oi_1 _23329_ (.A1(_03009_),
    .A2(_03006_),
    .Y(_00606_),
    .B1(_03010_));
 sg13g2_nor2_1 _23330_ (.A(\spi.sdi_r[3] ),
    .B(_03006_),
    .Y(_03012_));
 sg13g2_a21oi_1 _23331_ (.A1(_00915_),
    .A2(_03006_),
    .Y(_00607_),
    .B1(_03012_));
 sg13g2_mux2_1 _23332_ (.A0(\spi.sdi_r[0] ),
    .A1(net4),
    .S(_01013_),
    .X(_00608_));
 sg13g2_mux2_1 _23333_ (.A0(\spi.sdi_r[1] ),
    .A1(net5),
    .S(_01013_),
    .X(_00609_));
 sg13g2_mux2_1 _23334_ (.A0(\spi.sdi_r[2] ),
    .A1(net6),
    .S(_01013_),
    .X(_00610_));
 sg13g2_mux2_1 _23335_ (.A0(\spi.sdi_r[3] ),
    .A1(net7),
    .S(_01013_),
    .X(_00611_));
 sg13g2_nand3_1 _23336_ (.B(_02794_),
    .C(net189),
    .A(_02741_),
    .Y(_03013_));
 sg13g2_nor2_1 _23337_ (.A(_03000_),
    .B(net189),
    .Y(_03014_));
 sg13g2_buf_1 _23338_ (.A(_03014_),
    .X(_03015_));
 sg13g2_inv_1 _23339_ (.Y(_03017_),
    .A(_03015_));
 sg13g2_o21ai_1 _23340_ (.B1(_01728_),
    .Y(_03018_),
    .A1(_01351_),
    .A2(_03017_));
 sg13g2_a21oi_2 _23341_ (.B1(_03018_),
    .Y(_03019_),
    .A2(net189),
    .A1(_01035_));
 sg13g2_inv_1 _23342_ (.Y(_03020_),
    .A(_03019_));
 sg13g2_a221oi_1 _23343_ (.B2(_03015_),
    .C1(_03020_),
    .B1(_00805_),
    .A1(_03000_),
    .Y(_03021_),
    .A2(\ss2[0] ));
 sg13g2_nor2_1 _23344_ (.A(_01891_),
    .B(_03019_),
    .Y(_03022_));
 sg13g2_a21oi_1 _23345_ (.A1(_03013_),
    .A2(_03021_),
    .Y(_00612_),
    .B1(_03022_));
 sg13g2_nand3_1 _23346_ (.B(_02867_),
    .C(net189),
    .A(_02823_),
    .Y(_03023_));
 sg13g2_a221oi_1 _23347_ (.B2(_03015_),
    .C1(_03020_),
    .B1(_00816_),
    .A1(_03000_),
    .Y(_03024_),
    .A2(\ss2[1] ));
 sg13g2_nor2_1 _23348_ (.A(_01902_),
    .B(_03019_),
    .Y(_03025_));
 sg13g2_a21oi_1 _23349_ (.A1(_03023_),
    .A2(_03024_),
    .Y(_00613_),
    .B1(_03025_));
 sg13g2_nand3_1 _23350_ (.B(_02893_),
    .C(net189),
    .A(_02876_),
    .Y(_03026_));
 sg13g2_a221oi_1 _23351_ (.B2(_03015_),
    .C1(_03020_),
    .B1(_00893_),
    .A1(_03000_),
    .Y(_03027_),
    .A2(\ss2[2] ));
 sg13g2_nor2_1 _23352_ (.A(_01858_),
    .B(_03019_),
    .Y(_03028_));
 sg13g2_a21oi_1 _23353_ (.A1(_03026_),
    .A2(_03027_),
    .Y(_00614_),
    .B1(_03028_));
 sg13g2_a221oi_1 _23354_ (.B2(_03015_),
    .C1(_03020_),
    .B1(_00904_),
    .A1(_03000_),
    .Y(_03029_),
    .A2(\ss2[3] ));
 sg13g2_nand2_1 _23355_ (.Y(_03030_),
    .A(_02901_),
    .B(net189));
 sg13g2_a22oi_1 _23356_ (.Y(_00615_),
    .B1(_03029_),
    .B2(_03030_),
    .A2(_03020_),
    .A1(_03568_));
 sg13g2_o21ai_1 _23357_ (.B1(_01514_),
    .Y(_03031_),
    .A1(\state[3] ),
    .A2(_03017_));
 sg13g2_a21o_1 _23358_ (.A2(net189),
    .A1(_01035_),
    .B1(_03031_),
    .X(_03032_));
 sg13g2_buf_1 _23359_ (.A(_03032_),
    .X(_03034_));
 sg13g2_a221oi_1 _23360_ (.B2(_03015_),
    .C1(_03034_),
    .B1(_00805_),
    .A1(_03000_),
    .Y(_03035_),
    .A2(\ss2[4] ));
 sg13g2_nand2_1 _23361_ (.Y(_03036_),
    .A(_02810_),
    .B(_02798_));
 sg13g2_a22oi_1 _23362_ (.Y(_00616_),
    .B1(_03035_),
    .B2(_03036_),
    .A2(_03034_),
    .A1(_03371_));
 sg13g2_a221oi_1 _23363_ (.B2(_03015_),
    .C1(_03034_),
    .B1(_00816_),
    .A1(_03000_),
    .Y(_03037_),
    .A2(\ss2[5] ));
 sg13g2_o21ai_1 _23364_ (.B1(net189),
    .Y(_03038_),
    .A1(_02816_),
    .A2(_02732_));
 sg13g2_a22oi_1 _23365_ (.Y(_00617_),
    .B1(_03037_),
    .B2(_03038_),
    .A2(_03034_),
    .A1(_03694_));
 sg13g2_nor2_1 _23366_ (.A(\ss2[0] ),
    .B(net121),
    .Y(_03039_));
 sg13g2_a21oi_1 _23367_ (.A1(_02426_),
    .A2(net121),
    .Y(_00618_),
    .B1(_03039_));
 sg13g2_nor2_1 _23368_ (.A(\ss2[1] ),
    .B(net121),
    .Y(_03040_));
 sg13g2_a21oi_1 _23369_ (.A1(_02950_),
    .A2(net121),
    .Y(_00619_),
    .B1(_03040_));
 sg13g2_nor2_1 _23370_ (.A(\ss2[2] ),
    .B(_01057_),
    .Y(_03041_));
 sg13g2_a21oi_1 _23371_ (.A1(_02404_),
    .A2(net121),
    .Y(_00620_),
    .B1(_03041_));
 sg13g2_nor2_1 _23372_ (.A(\ss2[3] ),
    .B(_01057_),
    .Y(_03042_));
 sg13g2_a21oi_1 _23373_ (.A1(_03568_),
    .A2(net121),
    .Y(_00621_),
    .B1(_03042_));
 sg13g2_nor2_1 _23374_ (.A(\ss2[4] ),
    .B(_01057_),
    .Y(_03043_));
 sg13g2_a21oi_1 _23375_ (.A1(_03371_),
    .A2(_00000_),
    .Y(_00622_),
    .B1(_03043_));
 sg13g2_nor2_1 _23376_ (.A(\ss2[5] ),
    .B(_01057_),
    .Y(_03044_));
 sg13g2_a21oi_1 _23377_ (.A1(_03694_),
    .A2(net121),
    .Y(_00623_),
    .B1(_03044_));
 sg13g2_a21oi_2 _23378_ (.B1(net184),
    .Y(_03045_),
    .A2(_00772_),
    .A1(_01373_));
 sg13g2_nand2_1 _23379_ (.Y(_03047_),
    .A(_03045_),
    .B(net97));
 sg13g2_o21ai_1 _23380_ (.B1(_03047_),
    .Y(_00624_),
    .A1(_01373_),
    .A2(_01621_));
 sg13g2_a21oi_1 _23381_ (.A1(_01557_),
    .A2(_01362_),
    .Y(_03048_),
    .B1(_00783_));
 sg13g2_nand2_1 _23382_ (.Y(_03049_),
    .A(_03045_),
    .B(_01979_));
 sg13g2_o21ai_1 _23383_ (.B1(_03049_),
    .Y(_00625_),
    .A1(_03045_),
    .A2(_03048_));
 sg13g2_nand2_1 _23384_ (.Y(_03050_),
    .A(_03045_),
    .B(_00274_));
 sg13g2_nor2_1 _23385_ (.A(_01286_),
    .B(_01308_),
    .Y(_03051_));
 sg13g2_nand3_1 _23386_ (.B(net184),
    .C(_01362_),
    .A(_03051_),
    .Y(_03052_));
 sg13g2_nand2_1 _23387_ (.Y(_00626_),
    .A(_03050_),
    .B(_03052_));
 sg13g2_nand2_1 _23388_ (.Y(_03053_),
    .A(_00772_),
    .B(_00783_));
 sg13g2_buf_2 _23389_ (.A(_03053_),
    .X(_03054_));
 sg13g2_nand2_1 _23390_ (.Y(_03055_),
    .A(_03054_),
    .B(\b.gen_square[0].sq.write_bus[0] ));
 sg13g2_o21ai_1 _23391_ (.B1(_03055_),
    .Y(_00627_),
    .A1(_01155_),
    .A2(_03054_));
 sg13g2_nand2_1 _23392_ (.Y(_03056_),
    .A(_03054_),
    .B(\b.gen_square[0].sq.write_bus[1] ));
 sg13g2_o21ai_1 _23393_ (.B1(_03056_),
    .Y(_00628_),
    .A1(_01546_),
    .A2(_03054_));
 sg13g2_nand2_1 _23394_ (.Y(_03057_),
    .A(_03054_),
    .B(\b.gen_square[0].sq.write_bus[2] ));
 sg13g2_o21ai_1 _23395_ (.B1(_03057_),
    .Y(_00629_),
    .A1(_03009_),
    .A2(_03054_));
 sg13g2_nor2_1 _23396_ (.A(_00904_),
    .B(_03054_),
    .Y(_03058_));
 sg13g2_a21oi_1 _23397_ (.A1(_02759_),
    .A2(_03054_),
    .Y(_00630_),
    .B1(_03058_));
 sg13g2_nor3_1 _23398_ (.A(_00904_),
    .B(_00069_),
    .C(_03009_),
    .Y(_03059_));
 sg13g2_nand3_1 _23399_ (.B(_00772_),
    .C(_01546_),
    .A(_03059_),
    .Y(_03061_));
 sg13g2_mux2_1 _23400_ (.A0(_00805_),
    .A1(net136),
    .S(_03061_),
    .X(_00631_));
 sg13g2_nor3_1 _23401_ (.A(_01979_),
    .B(net192),
    .C(_01957_),
    .Y(_03062_));
 sg13g2_inv_1 _23402_ (.Y(_03063_),
    .A(_03062_));
 sg13g2_buf_1 _23403_ (.A(_03063_),
    .X(_03064_));
 sg13g2_buf_1 _23404_ (.A(net141),
    .X(_03065_));
 sg13g2_nor2b_1 _23405_ (.A(net125),
    .B_N(net131),
    .Y(_03066_));
 sg13g2_inv_1 _23406_ (.Y(_03067_),
    .A(_01935_));
 sg13g2_a21oi_1 _23407_ (.A1(_03066_),
    .A2(_03067_),
    .Y(_03068_),
    .B1(_10429_));
 sg13g2_nor2_1 _23408_ (.A(\mask_mode[2] ),
    .B(_01642_),
    .Y(_03069_));
 sg13g2_inv_1 _23409_ (.Y(_03070_),
    .A(_03069_));
 sg13g2_buf_2 _23410_ (.A(_03070_),
    .X(_03071_));
 sg13g2_nor2_1 _23411_ (.A(_01264_),
    .B(net175),
    .Y(_03072_));
 sg13g2_inv_1 _23412_ (.Y(_03073_),
    .A(_03072_));
 sg13g2_buf_1 _23413_ (.A(_03073_),
    .X(_03074_));
 sg13g2_buf_1 _23414_ (.A(net124),
    .X(_03075_));
 sg13g2_inv_1 _23415_ (.Y(_03076_),
    .A(_03068_));
 sg13g2_o21ai_1 _23416_ (.B1(_03076_),
    .Y(_03077_),
    .A1(net209),
    .A2(_04844_));
 sg13g2_buf_1 _23417_ (.A(net175),
    .X(_03078_));
 sg13g2_nand3_1 _23418_ (.B(_03067_),
    .C(net157),
    .A(_03077_),
    .Y(_03079_));
 sg13g2_nor2_1 _23419_ (.A(_01220_),
    .B(_03072_),
    .Y(_03081_));
 sg13g2_buf_1 _23420_ (.A(_03081_),
    .X(_03082_));
 sg13g2_buf_1 _23421_ (.A(net123),
    .X(_03083_));
 sg13g2_nand2_1 _23422_ (.Y(_03084_),
    .A(_03079_),
    .B(net110));
 sg13g2_o21ai_1 _23423_ (.B1(_03084_),
    .Y(_00275_),
    .A1(_03068_),
    .A2(net111));
 sg13g2_buf_1 _23424_ (.A(_03062_),
    .X(_03085_));
 sg13g2_buf_1 _23425_ (.A(net156),
    .X(_03086_));
 sg13g2_nand2_1 _23426_ (.Y(_03087_),
    .A(net140),
    .B(_06324_));
 sg13g2_o21ai_1 _23427_ (.B1(_09632_),
    .Y(_03088_),
    .A1(_03087_),
    .A2(_02481_));
 sg13g2_buf_1 _23428_ (.A(_03069_),
    .X(_03089_));
 sg13g2_buf_1 _23429_ (.A(_03089_),
    .X(_03091_));
 sg13g2_buf_1 _23430_ (.A(_01642_),
    .X(_03092_));
 sg13g2_nand3_1 _23431_ (.B(_06324_),
    .C(net214),
    .A(_06322_),
    .Y(_03093_));
 sg13g2_o21ai_1 _23432_ (.B1(_03093_),
    .Y(_03094_),
    .A1(net174),
    .A2(_03088_));
 sg13g2_a21oi_1 _23433_ (.A1(_03094_),
    .A2(_02470_),
    .Y(_03095_),
    .B1(net229));
 sg13g2_buf_2 _23434_ (.A(net124),
    .X(_03096_));
 sg13g2_mux2_1 _23435_ (.A0(_03088_),
    .A1(_03095_),
    .S(net109),
    .X(_00276_));
 sg13g2_nand2_1 _23436_ (.Y(_03097_),
    .A(net140),
    .B(_06521_));
 sg13g2_o21ai_1 _23437_ (.B1(_09763_),
    .Y(_03098_),
    .A1(_03097_),
    .A2(_02642_));
 sg13g2_nand3_1 _23438_ (.B(_06521_),
    .C(net214),
    .A(_06519_),
    .Y(_03099_));
 sg13g2_o21ai_1 _23439_ (.B1(_03099_),
    .Y(_03101_),
    .A1(net174),
    .A2(_03098_));
 sg13g2_inv_1 _23440_ (.Y(_03102_),
    .A(_02642_));
 sg13g2_a21oi_1 _23441_ (.A1(_03101_),
    .A2(_03102_),
    .Y(_03103_),
    .B1(net229));
 sg13g2_mux2_1 _23442_ (.A0(_03098_),
    .A1(_03103_),
    .S(net109),
    .X(_00277_));
 sg13g2_buf_1 _23443_ (.A(net156),
    .X(_03104_));
 sg13g2_nand2_1 _23444_ (.Y(_03105_),
    .A(net139),
    .B(_06945_));
 sg13g2_o21ai_1 _23445_ (.B1(_09890_),
    .Y(_03106_),
    .A1(_02814_),
    .A2(_03105_));
 sg13g2_nand3_1 _23446_ (.B(_06945_),
    .C(net214),
    .A(_06943_),
    .Y(_03107_));
 sg13g2_o21ai_1 _23447_ (.B1(_03107_),
    .Y(_03108_),
    .A1(net174),
    .A2(_03106_));
 sg13g2_a21oi_1 _23448_ (.A1(_03108_),
    .A2(_02824_),
    .Y(_03109_),
    .B1(net229));
 sg13g2_mux2_1 _23449_ (.A0(_03106_),
    .A1(_03109_),
    .S(net109),
    .X(_00278_));
 sg13g2_nand2_1 _23450_ (.Y(_03111_),
    .A(net140),
    .B(_05884_));
 sg13g2_o21ai_1 _23451_ (.B1(_09169_),
    .Y(_03112_),
    .A1(_03111_),
    .A2(_02994_));
 sg13g2_nand3_1 _23452_ (.B(_05884_),
    .C(net214),
    .A(_05879_),
    .Y(_03113_));
 sg13g2_o21ai_1 _23453_ (.B1(_03113_),
    .Y(_03114_),
    .A1(net174),
    .A2(_03112_));
 sg13g2_inv_1 _23454_ (.Y(_03115_),
    .A(_02994_));
 sg13g2_a21oi_1 _23455_ (.A1(_03114_),
    .A2(_03115_),
    .Y(_03116_),
    .B1(net229));
 sg13g2_buf_1 _23456_ (.A(net124),
    .X(_03117_));
 sg13g2_mux2_1 _23457_ (.A0(_03112_),
    .A1(_03116_),
    .S(net108),
    .X(_00279_));
 sg13g2_nand2_1 _23458_ (.Y(_03118_),
    .A(net140),
    .B(_04189_));
 sg13g2_o21ai_1 _23459_ (.B1(_09046_),
    .Y(_03120_),
    .A1(_03118_),
    .A2(_03119_));
 sg13g2_nand3_1 _23460_ (.B(_04189_),
    .C(net214),
    .A(_04183_),
    .Y(_03121_));
 sg13g2_o21ai_1 _23461_ (.B1(_03121_),
    .Y(_03122_),
    .A1(_03091_),
    .A2(_03120_));
 sg13g2_inv_1 _23462_ (.Y(_03123_),
    .A(_03119_));
 sg13g2_a21oi_1 _23463_ (.A1(_03122_),
    .A2(_03123_),
    .Y(_03124_),
    .B1(net229));
 sg13g2_mux2_1 _23464_ (.A0(_03120_),
    .A1(_03124_),
    .S(net108),
    .X(_00280_));
 sg13g2_nand2_1 _23465_ (.Y(_03125_),
    .A(_03086_),
    .B(net159));
 sg13g2_o21ai_1 _23466_ (.B1(_10067_),
    .Y(_03126_),
    .A1(_03125_),
    .A2(_03260_));
 sg13g2_nand3_1 _23467_ (.B(net159),
    .C(_03092_),
    .A(_10051_),
    .Y(_03127_));
 sg13g2_o21ai_1 _23468_ (.B1(_03127_),
    .Y(_03128_),
    .A1(net174),
    .A2(_03126_));
 sg13g2_inv_1 _23469_ (.Y(_03130_),
    .A(_03260_));
 sg13g2_a21oi_1 _23470_ (.A1(_03128_),
    .A2(_03130_),
    .Y(_03131_),
    .B1(net229));
 sg13g2_mux2_1 _23471_ (.A0(_03126_),
    .A1(_03131_),
    .S(net108),
    .X(_00281_));
 sg13g2_nor2_1 _23472_ (.A(_06022_),
    .B(net125),
    .Y(_03132_));
 sg13g2_inv_1 _23473_ (.Y(_03133_),
    .A(_03409_));
 sg13g2_a21oi_1 _23474_ (.A1(_03132_),
    .A2(_03133_),
    .Y(_03134_),
    .B1(_11265_));
 sg13g2_inv_1 _23475_ (.Y(_03135_),
    .A(_03134_));
 sg13g2_o21ai_1 _23476_ (.B1(_03135_),
    .Y(_03136_),
    .A1(net209),
    .A2(_11155_));
 sg13g2_nand3_1 _23477_ (.B(_03133_),
    .C(net157),
    .A(_03136_),
    .Y(_03137_));
 sg13g2_nand2_1 _23478_ (.Y(_03138_),
    .A(_03137_),
    .B(net110));
 sg13g2_o21ai_1 _23479_ (.B1(_03138_),
    .Y(_00282_),
    .A1(net111),
    .A2(_03134_));
 sg13g2_nand2_1 _23480_ (.Y(_03140_),
    .A(net139),
    .B(_05577_));
 sg13g2_o21ai_1 _23481_ (.B1(_11236_),
    .Y(_03141_),
    .A1(_03528_),
    .A2(_03140_));
 sg13g2_nand3_1 _23482_ (.B(_05577_),
    .C(net214),
    .A(_05625_),
    .Y(_03142_));
 sg13g2_o21ai_1 _23483_ (.B1(_03142_),
    .Y(_03143_),
    .A1(net174),
    .A2(_03141_));
 sg13g2_inv_1 _23484_ (.Y(_03144_),
    .A(_03528_));
 sg13g2_a21oi_1 _23485_ (.A1(_03143_),
    .A2(_03144_),
    .Y(_03145_),
    .B1(_01231_));
 sg13g2_mux2_1 _23486_ (.A0(_03141_),
    .A1(_03145_),
    .S(net108),
    .X(_00283_));
 sg13g2_nand2_1 _23487_ (.Y(_03146_),
    .A(net139),
    .B(_04806_));
 sg13g2_o21ai_1 _23488_ (.B1(_11114_),
    .Y(_03147_),
    .A1(_03537_),
    .A2(_03146_));
 sg13g2_nand3_1 _23489_ (.B(_04806_),
    .C(net214),
    .A(_04804_),
    .Y(_03149_));
 sg13g2_o21ai_1 _23490_ (.B1(_03149_),
    .Y(_03150_),
    .A1(net174),
    .A2(_03147_));
 sg13g2_inv_1 _23491_ (.Y(_03151_),
    .A(_03537_));
 sg13g2_a21oi_1 _23492_ (.A1(_03150_),
    .A2(_03151_),
    .Y(_03152_),
    .B1(net229));
 sg13g2_mux2_1 _23493_ (.A0(_03147_),
    .A1(_03152_),
    .S(net108),
    .X(_00284_));
 sg13g2_nand2_1 _23494_ (.Y(_03153_),
    .A(_03104_),
    .B(_06573_));
 sg13g2_o21ai_1 _23495_ (.B1(_11365_),
    .Y(_03154_),
    .A1(_03550_),
    .A2(_03153_));
 sg13g2_nand3_1 _23496_ (.B(_06573_),
    .C(net214),
    .A(_06568_),
    .Y(_03155_));
 sg13g2_o21ai_1 _23497_ (.B1(_03155_),
    .Y(_03156_),
    .A1(net174),
    .A2(_03154_));
 sg13g2_inv_1 _23498_ (.Y(_03157_),
    .A(_03550_));
 sg13g2_a21oi_1 _23499_ (.A1(_03156_),
    .A2(_03157_),
    .Y(_03158_),
    .B1(net229));
 sg13g2_mux2_1 _23500_ (.A0(_03154_),
    .A1(_03158_),
    .S(net108),
    .X(_00285_));
 sg13g2_buf_1 _23501_ (.A(net125),
    .X(_03159_));
 sg13g2_nor2_1 _23502_ (.A(_05603_),
    .B(net107),
    .Y(_03160_));
 sg13g2_inv_1 _23503_ (.Y(_03161_),
    .A(_03559_));
 sg13g2_a21oi_1 _23504_ (.A1(_03160_),
    .A2(_03161_),
    .Y(_03162_),
    .B1(_10540_));
 sg13g2_buf_1 _23505_ (.A(net175),
    .X(_03163_));
 sg13g2_nand2_1 _23506_ (.Y(_03164_),
    .A(_03161_),
    .B(net155));
 sg13g2_buf_1 _23507_ (.A(_01642_),
    .X(_03165_));
 sg13g2_buf_1 _23508_ (.A(net213),
    .X(_03166_));
 sg13g2_a21oi_1 _23509_ (.A1(net187),
    .A2(_10496_),
    .Y(_03168_),
    .B1(_03162_));
 sg13g2_buf_1 _23510_ (.A(net123),
    .X(_03169_));
 sg13g2_o21ai_1 _23511_ (.B1(net106),
    .Y(_03170_),
    .A1(_03164_),
    .A2(_03168_));
 sg13g2_o21ai_1 _23512_ (.B1(_03170_),
    .Y(_00286_),
    .A1(net111),
    .A2(_03162_));
 sg13g2_nand2_1 _23513_ (.Y(_03171_),
    .A(_03086_),
    .B(_05854_));
 sg13g2_o21ai_1 _23514_ (.B1(_11452_),
    .Y(_03172_),
    .A1(_03171_),
    .A2(_03572_));
 sg13g2_buf_1 _23515_ (.A(_01642_),
    .X(_03173_));
 sg13g2_nand3_1 _23516_ (.B(_05854_),
    .C(_03173_),
    .A(_05852_),
    .Y(_03174_));
 sg13g2_o21ai_1 _23517_ (.B1(_03174_),
    .Y(_03175_),
    .A1(_03091_),
    .A2(_03172_));
 sg13g2_inv_1 _23518_ (.Y(_03176_),
    .A(_03572_));
 sg13g2_buf_1 _23519_ (.A(_01220_),
    .X(_03177_));
 sg13g2_buf_1 _23520_ (.A(net211),
    .X(_03178_));
 sg13g2_a21oi_1 _23521_ (.A1(_03175_),
    .A2(_03176_),
    .Y(_03179_),
    .B1(_03178_));
 sg13g2_mux2_1 _23522_ (.A0(_03172_),
    .A1(_03179_),
    .S(net108),
    .X(_00287_));
 sg13g2_buf_1 _23523_ (.A(_03085_),
    .X(_03180_));
 sg13g2_nand2_1 _23524_ (.Y(_03181_),
    .A(_03180_),
    .B(_05280_));
 sg13g2_o21ai_1 _23525_ (.B1(_11547_),
    .Y(_03182_),
    .A1(_03181_),
    .A2(_03583_));
 sg13g2_buf_1 _23526_ (.A(_03089_),
    .X(_03183_));
 sg13g2_nand3_1 _23527_ (.B(_05280_),
    .C(net212),
    .A(_05278_),
    .Y(_03184_));
 sg13g2_o21ai_1 _23528_ (.B1(_03184_),
    .Y(_03185_),
    .A1(_03183_),
    .A2(_03182_));
 sg13g2_a21oi_1 _23529_ (.A1(_03185_),
    .A2(_03582_),
    .Y(_03187_),
    .B1(net186));
 sg13g2_mux2_1 _23530_ (.A0(_03182_),
    .A1(_03187_),
    .S(_03117_),
    .X(_00288_));
 sg13g2_nand2_1 _23531_ (.Y(_03188_),
    .A(_03180_),
    .B(net116));
 sg13g2_o21ai_1 _23532_ (.B1(_11042_),
    .Y(_03189_),
    .A1(_03188_),
    .A2(_03594_));
 sg13g2_nand3_1 _23533_ (.B(net116),
    .C(net212),
    .A(_04206_),
    .Y(_03190_));
 sg13g2_o21ai_1 _23534_ (.B1(_03190_),
    .Y(_03191_),
    .A1(net173),
    .A2(_03189_));
 sg13g2_a21oi_1 _23535_ (.A1(_03191_),
    .A2(_03593_),
    .Y(_03192_),
    .B1(net186));
 sg13g2_mux2_1 _23536_ (.A0(_03189_),
    .A1(_03192_),
    .S(_03117_),
    .X(_00289_));
 sg13g2_nor2_1 _23537_ (.A(_07519_),
    .B(_03159_),
    .Y(_03193_));
 sg13g2_inv_1 _23538_ (.Y(_03194_),
    .A(_11666_));
 sg13g2_a21oi_1 _23539_ (.A1(_03193_),
    .A2(_06674_),
    .Y(_03195_),
    .B1(_03194_));
 sg13g2_nand2_1 _23540_ (.Y(_03196_),
    .A(_06674_),
    .B(_03163_));
 sg13g2_a21oi_1 _23541_ (.A1(net187),
    .A2(_11614_),
    .Y(_03197_),
    .B1(_03195_));
 sg13g2_o21ai_1 _23542_ (.B1(_03169_),
    .Y(_03198_),
    .A1(_03196_),
    .A2(_03197_));
 sg13g2_o21ai_1 _23543_ (.B1(_03198_),
    .Y(_00290_),
    .A1(net111),
    .A2(_03195_));
 sg13g2_nor2_1 _23544_ (.A(_06065_),
    .B(net107),
    .Y(_03199_));
 sg13g2_a21oi_1 _23545_ (.A1(_03199_),
    .A2(_06042_),
    .Y(_03200_),
    .B1(_11876_));
 sg13g2_nand2_1 _23546_ (.Y(_03201_),
    .A(_06042_),
    .B(net155));
 sg13g2_a21oi_1 _23547_ (.A1(net187),
    .A2(_11921_),
    .Y(_03202_),
    .B1(_03200_));
 sg13g2_o21ai_1 _23548_ (.B1(net106),
    .Y(_03203_),
    .A1(_03201_),
    .A2(_03202_));
 sg13g2_o21ai_1 _23549_ (.B1(_03203_),
    .Y(_00291_),
    .A1(net111),
    .A2(_03200_));
 sg13g2_nand2_1 _23550_ (.Y(_03205_),
    .A(net138),
    .B(_05637_));
 sg13g2_o21ai_1 _23551_ (.B1(_11980_),
    .Y(_03206_),
    .A1(_03205_),
    .A2(_03625_));
 sg13g2_nand3_1 _23552_ (.B(_05637_),
    .C(net212),
    .A(_05635_),
    .Y(_03207_));
 sg13g2_o21ai_1 _23553_ (.B1(_03207_),
    .Y(_03208_),
    .A1(net173),
    .A2(_03206_));
 sg13g2_a21oi_1 _23554_ (.A1(_03208_),
    .A2(_03624_),
    .Y(_03209_),
    .B1(net186));
 sg13g2_mux2_1 _23555_ (.A0(_03206_),
    .A1(_03209_),
    .S(net108),
    .X(_00292_));
 sg13g2_nand3_1 _23556_ (.B(net127),
    .C(net139),
    .A(_06386_),
    .Y(_03210_));
 sg13g2_nand2_1 _23557_ (.Y(_03211_),
    .A(_03210_),
    .B(_11861_));
 sg13g2_nand3_1 _23558_ (.B(net127),
    .C(net212),
    .A(_06379_),
    .Y(_03212_));
 sg13g2_o21ai_1 _23559_ (.B1(_03212_),
    .Y(_03213_),
    .A1(net173),
    .A2(_03211_));
 sg13g2_a21oi_1 _23560_ (.A1(_03213_),
    .A2(_06386_),
    .Y(_03214_),
    .B1(net186));
 sg13g2_buf_1 _23561_ (.A(net124),
    .X(_03215_));
 sg13g2_mux2_1 _23562_ (.A0(_03211_),
    .A1(_03214_),
    .S(net105),
    .X(_00293_));
 sg13g2_nand2_1 _23563_ (.Y(_03216_),
    .A(net138),
    .B(_04887_));
 sg13g2_o21ai_1 _23564_ (.B1(_11794_),
    .Y(_03217_),
    .A1(_03216_),
    .A2(_03640_));
 sg13g2_nand3_1 _23565_ (.B(_04887_),
    .C(net212),
    .A(_04885_),
    .Y(_03218_));
 sg13g2_o21ai_1 _23566_ (.B1(_03218_),
    .Y(_03219_),
    .A1(net173),
    .A2(_03217_));
 sg13g2_a21oi_1 _23567_ (.A1(_03219_),
    .A2(_04892_),
    .Y(_03220_),
    .B1(net186));
 sg13g2_mux2_1 _23568_ (.A0(_03217_),
    .A1(_03220_),
    .S(net105),
    .X(_00294_));
 sg13g2_nand2_1 _23569_ (.Y(_03222_),
    .A(_03104_),
    .B(_05337_));
 sg13g2_o21ai_1 _23570_ (.B1(_00749_),
    .Y(_03223_),
    .A1(_03651_),
    .A2(_03222_));
 sg13g2_nand3_1 _23571_ (.B(_05337_),
    .C(_03173_),
    .A(_05335_),
    .Y(_03224_));
 sg13g2_o21ai_1 _23572_ (.B1(_03224_),
    .Y(_03225_),
    .A1(_03183_),
    .A2(_03223_));
 sg13g2_inv_1 _23573_ (.Y(_03226_),
    .A(_03651_));
 sg13g2_a21oi_1 _23574_ (.A1(_03225_),
    .A2(_03226_),
    .Y(_03227_),
    .B1(_03178_));
 sg13g2_mux2_1 _23575_ (.A0(_03223_),
    .A1(_03227_),
    .S(_03215_),
    .X(_00295_));
 sg13g2_nand2_1 _23576_ (.Y(_03228_),
    .A(net138),
    .B(_06177_));
 sg13g2_o21ai_1 _23577_ (.B1(_00851_),
    .Y(_03229_),
    .A1(_03228_),
    .A2(_03659_));
 sg13g2_nand3_1 _23578_ (.B(_06177_),
    .C(net212),
    .A(_06220_),
    .Y(_03230_));
 sg13g2_o21ai_1 _23579_ (.B1(_03230_),
    .Y(_03232_),
    .A1(net173),
    .A2(_03229_));
 sg13g2_inv_1 _23580_ (.Y(_03233_),
    .A(_03659_));
 sg13g2_a21oi_1 _23581_ (.A1(_03232_),
    .A2(_03233_),
    .Y(_03234_),
    .B1(net186));
 sg13g2_mux2_1 _23582_ (.A0(_03229_),
    .A1(_03234_),
    .S(net105),
    .X(_00296_));
 sg13g2_nor2_1 _23583_ (.A(_06351_),
    .B(net125),
    .Y(_03235_));
 sg13g2_inv_1 _23584_ (.Y(_03236_),
    .A(_03670_));
 sg13g2_a21oi_1 _23585_ (.A1(_03235_),
    .A2(_03236_),
    .Y(_03237_),
    .B1(_10570_));
 sg13g2_inv_1 _23586_ (.Y(_03238_),
    .A(_03237_));
 sg13g2_o21ai_1 _23587_ (.B1(_03238_),
    .Y(_03239_),
    .A1(_01664_),
    .A2(_10566_));
 sg13g2_nand3_1 _23588_ (.B(_03236_),
    .C(_03078_),
    .A(_03239_),
    .Y(_03240_));
 sg13g2_nand2_1 _23589_ (.Y(_03242_),
    .A(_03240_),
    .B(_03083_));
 sg13g2_o21ai_1 _23590_ (.B1(_03242_),
    .Y(_00297_),
    .A1(_03075_),
    .A2(_03237_));
 sg13g2_nand2_1 _23591_ (.Y(_03243_),
    .A(net138),
    .B(_04148_));
 sg13g2_o21ai_1 _23592_ (.B1(_00961_),
    .Y(_03244_),
    .A1(_03243_),
    .A2(_03678_));
 sg13g2_nand3_1 _23593_ (.B(_04148_),
    .C(net212),
    .A(_04140_),
    .Y(_03245_));
 sg13g2_o21ai_1 _23594_ (.B1(_03245_),
    .Y(_03246_),
    .A1(net173),
    .A2(_03244_));
 sg13g2_a21oi_1 _23595_ (.A1(_03246_),
    .A2(_04143_),
    .Y(_03247_),
    .B1(net186));
 sg13g2_mux2_1 _23596_ (.A0(_03244_),
    .A1(_03247_),
    .S(net105),
    .X(_00298_));
 sg13g2_inv_1 _23597_ (.Y(_03248_),
    .A(_03686_));
 sg13g2_nor2_1 _23598_ (.A(_06855_),
    .B(net125),
    .Y(_03249_));
 sg13g2_a21oi_1 _23599_ (.A1(_03248_),
    .A2(_03249_),
    .Y(_03251_),
    .B1(_01059_));
 sg13g2_nand2_1 _23600_ (.Y(_03252_),
    .A(_03248_),
    .B(net155));
 sg13g2_a21oi_1 _23601_ (.A1(net187),
    .A2(_01052_),
    .Y(_03253_),
    .B1(_03251_));
 sg13g2_o21ai_1 _23602_ (.B1(net106),
    .Y(_03254_),
    .A1(_03252_),
    .A2(_03253_));
 sg13g2_o21ai_1 _23603_ (.B1(_03254_),
    .Y(_00299_),
    .A1(net111),
    .A2(_03251_));
 sg13g2_nor2_1 _23604_ (.A(_06084_),
    .B(net107),
    .Y(_03255_));
 sg13g2_inv_1 _23605_ (.Y(_03256_),
    .A(_03698_));
 sg13g2_a21oi_1 _23606_ (.A1(_03255_),
    .A2(_03256_),
    .Y(_03257_),
    .B1(_08244_));
 sg13g2_nand2_1 _23607_ (.Y(_03258_),
    .A(_03256_),
    .B(net155));
 sg13g2_a21oi_1 _23608_ (.A1(net187),
    .A2(_08515_),
    .Y(_03259_),
    .B1(_03257_));
 sg13g2_o21ai_1 _23609_ (.B1(net106),
    .Y(_03261_),
    .A1(_03258_),
    .A2(_03259_));
 sg13g2_o21ai_1 _23610_ (.B1(_03261_),
    .Y(_00300_),
    .A1(net111),
    .A2(_03257_));
 sg13g2_nand2_1 _23611_ (.Y(_03262_),
    .A(net139),
    .B(_05668_));
 sg13g2_o21ai_1 _23612_ (.B1(_08372_),
    .Y(_03263_),
    .A1(_03706_),
    .A2(_03262_));
 sg13g2_nand3_1 _23613_ (.B(_05668_),
    .C(net212),
    .A(_05666_),
    .Y(_03264_));
 sg13g2_o21ai_1 _23614_ (.B1(_03264_),
    .Y(_03265_),
    .A1(net173),
    .A2(_03263_));
 sg13g2_inv_1 _23615_ (.Y(_03266_),
    .A(_03706_));
 sg13g2_a21oi_1 _23616_ (.A1(_03265_),
    .A2(_03266_),
    .Y(_03267_),
    .B1(net186));
 sg13g2_mux2_1 _23617_ (.A0(_03263_),
    .A1(_03267_),
    .S(net105),
    .X(_00301_));
 sg13g2_nand2_1 _23618_ (.Y(_03268_),
    .A(net139),
    .B(_05129_));
 sg13g2_o21ai_1 _23619_ (.B1(_08150_),
    .Y(_03270_),
    .A1(_03714_),
    .A2(_03268_));
 sg13g2_buf_1 _23620_ (.A(_01642_),
    .X(_03271_));
 sg13g2_nand3_1 _23621_ (.B(_05129_),
    .C(net210),
    .A(_05842_),
    .Y(_03272_));
 sg13g2_o21ai_1 _23622_ (.B1(_03272_),
    .Y(_03273_),
    .A1(net173),
    .A2(_03270_));
 sg13g2_inv_1 _23623_ (.Y(_03274_),
    .A(_03714_));
 sg13g2_buf_1 _23624_ (.A(_03177_),
    .X(_03275_));
 sg13g2_a21oi_1 _23625_ (.A1(_03273_),
    .A2(_03274_),
    .Y(_03276_),
    .B1(net185));
 sg13g2_mux2_1 _23626_ (.A0(_03270_),
    .A1(_03276_),
    .S(net105),
    .X(_00302_));
 sg13g2_nand2_1 _23627_ (.Y(_03277_),
    .A(net140),
    .B(_05368_));
 sg13g2_o21ai_1 _23628_ (.B1(_08479_),
    .Y(_03278_),
    .A1(_03722_),
    .A2(_03277_));
 sg13g2_buf_1 _23629_ (.A(net188),
    .X(_03280_));
 sg13g2_nand3_1 _23630_ (.B(_05368_),
    .C(net210),
    .A(_05366_),
    .Y(_03281_));
 sg13g2_o21ai_1 _23631_ (.B1(_03281_),
    .Y(_03282_),
    .A1(net172),
    .A2(_03278_));
 sg13g2_inv_1 _23632_ (.Y(_03283_),
    .A(_03722_));
 sg13g2_a21oi_1 _23633_ (.A1(_03282_),
    .A2(_03283_),
    .Y(_03284_),
    .B1(net185));
 sg13g2_mux2_1 _23634_ (.A0(_03278_),
    .A1(_03284_),
    .S(net105),
    .X(_00303_));
 sg13g2_nand2_1 _23635_ (.Y(_03285_),
    .A(net138),
    .B(net146));
 sg13g2_o21ai_1 _23636_ (.B1(\b.gen_square[36].sq.mask ),
    .Y(_03286_),
    .A1(_03285_),
    .A2(_03730_));
 sg13g2_nand3_1 _23637_ (.B(net146),
    .C(net210),
    .A(_04916_),
    .Y(_03287_));
 sg13g2_o21ai_1 _23638_ (.B1(_03287_),
    .Y(_03288_),
    .A1(net172),
    .A2(_03286_));
 sg13g2_inv_1 _23639_ (.Y(_03290_),
    .A(_03730_));
 sg13g2_a21oi_1 _23640_ (.A1(_03288_),
    .A2(_03290_),
    .Y(_03291_),
    .B1(net185));
 sg13g2_mux2_1 _23641_ (.A0(_03286_),
    .A1(_03291_),
    .S(net105),
    .X(_00304_));
 sg13g2_nand2_1 _23642_ (.Y(_03292_),
    .A(net138),
    .B(_04532_));
 sg13g2_o21ai_1 _23643_ (.B1(_07859_),
    .Y(_03293_),
    .A1(_03292_),
    .A2(_03742_));
 sg13g2_nand3_1 _23644_ (.B(net164),
    .C(net210),
    .A(_06694_),
    .Y(_03294_));
 sg13g2_o21ai_1 _23645_ (.B1(_03294_),
    .Y(_03295_),
    .A1(_03280_),
    .A2(_03293_));
 sg13g2_a21oi_1 _23646_ (.A1(_03295_),
    .A2(_03741_),
    .Y(_03296_),
    .B1(net185));
 sg13g2_mux2_1 _23647_ (.A0(_03293_),
    .A1(_03296_),
    .S(_03215_),
    .X(_00305_));
 sg13g2_nand2_1 _23648_ (.Y(_03297_),
    .A(net138),
    .B(_04110_));
 sg13g2_o21ai_1 _23649_ (.B1(_08757_),
    .Y(_03298_),
    .A1(_03297_),
    .A2(_03751_));
 sg13g2_nand3_1 _23650_ (.B(_04110_),
    .C(_03271_),
    .A(_04105_),
    .Y(_03299_));
 sg13g2_o21ai_1 _23651_ (.B1(_03299_),
    .Y(_03300_),
    .A1(_03280_),
    .A2(_03298_));
 sg13g2_a21oi_1 _23652_ (.A1(_03300_),
    .A2(_03750_),
    .Y(_03301_),
    .B1(_03275_));
 sg13g2_buf_1 _23653_ (.A(_03073_),
    .X(_03302_));
 sg13g2_mux2_1 _23654_ (.A0(_03298_),
    .A1(_03301_),
    .S(_03302_),
    .X(_00306_));
 sg13g2_inv_1 _23655_ (.Y(_03303_),
    .A(_03763_));
 sg13g2_nor2_1 _23656_ (.A(_07535_),
    .B(net141),
    .Y(_03304_));
 sg13g2_inv_1 _23657_ (.Y(_03305_),
    .A(_08868_));
 sg13g2_a21oi_1 _23658_ (.A1(_03303_),
    .A2(_03304_),
    .Y(_03306_),
    .B1(_03305_));
 sg13g2_inv_1 _23659_ (.Y(_03308_),
    .A(_03306_));
 sg13g2_o21ai_1 _23660_ (.B1(_03308_),
    .Y(_03309_),
    .A1(net209),
    .A2(_08879_));
 sg13g2_nand3_1 _23661_ (.B(_03303_),
    .C(net157),
    .A(_03309_),
    .Y(_03310_));
 sg13g2_nand2_1 _23662_ (.Y(_03311_),
    .A(_03310_),
    .B(net110));
 sg13g2_o21ai_1 _23663_ (.B1(_03311_),
    .Y(_00307_),
    .A1(net111),
    .A2(_03306_));
 sg13g2_nor2_1 _23664_ (.A(_06541_),
    .B(net141),
    .Y(_03312_));
 sg13g2_a21oi_1 _23665_ (.A1(_03312_),
    .A2(_03771_),
    .Y(_03313_),
    .B1(_10665_));
 sg13g2_inv_1 _23666_ (.Y(_03314_),
    .A(_03313_));
 sg13g2_o21ai_1 _23667_ (.B1(_03314_),
    .Y(_03315_),
    .A1(_01664_),
    .A2(_10681_));
 sg13g2_nand3_1 _23668_ (.B(_03771_),
    .C(_03078_),
    .A(_03315_),
    .Y(_03316_));
 sg13g2_nand2_1 _23669_ (.Y(_03317_),
    .A(_03316_),
    .B(_03083_));
 sg13g2_o21ai_1 _23670_ (.B1(_03317_),
    .Y(_00308_),
    .A1(_03075_),
    .A2(_03313_));
 sg13g2_buf_1 _23671_ (.A(net124),
    .X(_03318_));
 sg13g2_nor2_1 _23672_ (.A(_05508_),
    .B(net107),
    .Y(_03319_));
 sg13g2_inv_1 _23673_ (.Y(_03320_),
    .A(_03779_));
 sg13g2_a21oi_1 _23674_ (.A1(_03319_),
    .A2(_03320_),
    .Y(_03321_),
    .B1(_01434_));
 sg13g2_nand2_1 _23675_ (.Y(_03322_),
    .A(_03320_),
    .B(net155));
 sg13g2_nor3_1 _23676_ (.A(_01653_),
    .B(_05496_),
    .C(_05508_),
    .Y(_03323_));
 sg13g2_nor2_1 _23677_ (.A(_03323_),
    .B(_03321_),
    .Y(_03324_));
 sg13g2_o21ai_1 _23678_ (.B1(net106),
    .Y(_03325_),
    .A1(_03322_),
    .A2(_03324_));
 sg13g2_o21ai_1 _23679_ (.B1(_03325_),
    .Y(_00309_),
    .A1(net104),
    .A2(_03321_));
 sg13g2_nand2_1 _23680_ (.Y(_03327_),
    .A(net138),
    .B(net190));
 sg13g2_o21ai_1 _23681_ (.B1(\b.gen_square[41].sq.mask ),
    .Y(_03328_),
    .A1(_03327_),
    .A2(_03788_));
 sg13g2_nand3_1 _23682_ (.B(_05555_),
    .C(net210),
    .A(_05566_),
    .Y(_03329_));
 sg13g2_o21ai_1 _23683_ (.B1(_03329_),
    .Y(_03330_),
    .A1(net172),
    .A2(_03328_));
 sg13g2_a21oi_1 _23684_ (.A1(_03330_),
    .A2(_03787_),
    .Y(_03331_),
    .B1(net185));
 sg13g2_mux2_1 _23685_ (.A0(_03328_),
    .A1(_03331_),
    .S(net122),
    .X(_00310_));
 sg13g2_nand2_1 _23686_ (.Y(_03332_),
    .A(net156),
    .B(_05398_));
 sg13g2_o21ai_1 _23687_ (.B1(_01543_),
    .Y(_03333_),
    .A1(_03332_),
    .A2(_03797_));
 sg13g2_nand3_1 _23688_ (.B(_05398_),
    .C(net210),
    .A(_05396_),
    .Y(_03334_));
 sg13g2_o21ai_1 _23689_ (.B1(_03334_),
    .Y(_03335_),
    .A1(net172),
    .A2(_03333_));
 sg13g2_a21oi_1 _23690_ (.A1(_03335_),
    .A2(_03796_),
    .Y(_03336_),
    .B1(net185));
 sg13g2_mux2_1 _23691_ (.A0(_03333_),
    .A1(_03336_),
    .S(net122),
    .X(_00311_));
 sg13g2_nand2_1 _23692_ (.Y(_03337_),
    .A(net156),
    .B(_05167_));
 sg13g2_o21ai_1 _23693_ (.B1(_01633_),
    .Y(_03338_),
    .A1(_03337_),
    .A2(_03805_));
 sg13g2_nand3_1 _23694_ (.B(net94),
    .C(net210),
    .A(_06196_),
    .Y(_03339_));
 sg13g2_o21ai_1 _23695_ (.B1(_03339_),
    .Y(_03340_),
    .A1(net172),
    .A2(_03338_));
 sg13g2_inv_1 _23696_ (.Y(_03341_),
    .A(_03805_));
 sg13g2_a21oi_1 _23697_ (.A1(_03340_),
    .A2(_03341_),
    .Y(_03342_),
    .B1(net185));
 sg13g2_mux2_1 _23698_ (.A0(_03338_),
    .A1(_03342_),
    .S(net122),
    .X(_00312_));
 sg13g2_nand2_1 _23699_ (.Y(_03344_),
    .A(net140),
    .B(_04513_));
 sg13g2_o21ai_1 _23700_ (.B1(\b.gen_square[44].sq.mask ),
    .Y(_03345_),
    .A1(_03813_),
    .A2(_03344_));
 sg13g2_nand3_1 _23701_ (.B(_04513_),
    .C(net210),
    .A(_06716_),
    .Y(_03346_));
 sg13g2_o21ai_1 _23702_ (.B1(_03346_),
    .Y(_03347_),
    .A1(net172),
    .A2(_03345_));
 sg13g2_inv_1 _23703_ (.Y(_03348_),
    .A(_03813_));
 sg13g2_a21oi_1 _23704_ (.A1(_03347_),
    .A2(_03348_),
    .Y(_03349_),
    .B1(net185));
 sg13g2_mux2_1 _23705_ (.A0(_03345_),
    .A1(_03349_),
    .S(_03302_),
    .X(_00313_));
 sg13g2_nand2_1 _23706_ (.Y(_03350_),
    .A(_03085_),
    .B(_04041_));
 sg13g2_o21ai_1 _23707_ (.B1(\b.gen_square[45].sq.mask ),
    .Y(_03351_),
    .A1(_03350_),
    .A2(_03821_));
 sg13g2_nand3_1 _23708_ (.B(_04041_),
    .C(_03271_),
    .A(_04946_),
    .Y(_03352_));
 sg13g2_o21ai_1 _23709_ (.B1(_03352_),
    .Y(_03353_),
    .A1(net172),
    .A2(_03351_));
 sg13g2_inv_1 _23710_ (.Y(_03354_),
    .A(_03821_));
 sg13g2_a21oi_1 _23711_ (.A1(_03353_),
    .A2(_03354_),
    .Y(_03355_),
    .B1(_03275_));
 sg13g2_mux2_1 _23712_ (.A0(_03351_),
    .A1(_03355_),
    .S(net122),
    .X(_00314_));
 sg13g2_nand2_1 _23713_ (.Y(_03356_),
    .A(net156),
    .B(net165));
 sg13g2_o21ai_1 _23714_ (.B1(_01236_),
    .Y(_03357_),
    .A1(_03356_),
    .A2(_03829_));
 sg13g2_nand3_1 _23715_ (.B(net165),
    .C(net213),
    .A(_04235_),
    .Y(_03358_));
 sg13g2_o21ai_1 _23716_ (.B1(_03358_),
    .Y(_03359_),
    .A1(net172),
    .A2(_03357_));
 sg13g2_inv_1 _23717_ (.Y(_03360_),
    .A(_03829_));
 sg13g2_a21oi_1 _23718_ (.A1(_03359_),
    .A2(_03360_),
    .Y(_03361_),
    .B1(net211));
 sg13g2_mux2_1 _23719_ (.A0(_03357_),
    .A1(_03361_),
    .S(net122),
    .X(_00315_));
 sg13g2_nor2_1 _23720_ (.A(_04392_),
    .B(net107),
    .Y(_03363_));
 sg13g2_a21oi_1 _23721_ (.A1(_04396_),
    .A2(_03363_),
    .Y(_03364_),
    .B1(_01882_));
 sg13g2_nand2_1 _23722_ (.Y(_03365_),
    .A(_04396_),
    .B(net155));
 sg13g2_nor3_1 _23723_ (.A(_01653_),
    .B(_04403_),
    .C(_04392_),
    .Y(_03366_));
 sg13g2_nor2_1 _23724_ (.A(_03366_),
    .B(_03364_),
    .Y(_03367_));
 sg13g2_o21ai_1 _23725_ (.B1(net106),
    .Y(_03368_),
    .A1(_03365_),
    .A2(_03367_));
 sg13g2_o21ai_1 _23726_ (.B1(_03368_),
    .Y(_00316_),
    .A1(net104),
    .A2(_03364_));
 sg13g2_nor2_1 _23727_ (.A(_04732_),
    .B(net141),
    .Y(_03369_));
 sg13g2_inv_1 _23728_ (.Y(_03370_),
    .A(_03850_));
 sg13g2_a21oi_1 _23729_ (.A1(_03369_),
    .A2(_03370_),
    .Y(_03372_),
    .B1(_07326_));
 sg13g2_inv_1 _23730_ (.Y(_03373_),
    .A(_03372_));
 sg13g2_o21ai_1 _23731_ (.B1(_03373_),
    .Y(_03374_),
    .A1(net209),
    .A2(_07350_));
 sg13g2_nand3_1 _23732_ (.B(_03370_),
    .C(net157),
    .A(_03374_),
    .Y(_03375_));
 sg13g2_nand2_1 _23733_ (.Y(_03376_),
    .A(_03375_),
    .B(net110));
 sg13g2_o21ai_1 _23734_ (.B1(_03376_),
    .Y(_00317_),
    .A1(net104),
    .A2(_03372_));
 sg13g2_nand2_1 _23735_ (.Y(_03377_),
    .A(_05124_),
    .B(net156));
 sg13g2_o21ai_1 _23736_ (.B1(_05808_),
    .Y(_03378_),
    .A1(_03860_),
    .A2(_03377_));
 sg13g2_nand3_1 _23737_ (.B(_04615_),
    .C(net213),
    .A(_05124_),
    .Y(_03379_));
 sg13g2_o21ai_1 _23738_ (.B1(_03379_),
    .Y(_03380_),
    .A1(net188),
    .A2(_03378_));
 sg13g2_a21oi_1 _23739_ (.A1(_03380_),
    .A2(_04741_),
    .Y(_03382_),
    .B1(net211));
 sg13g2_mux2_1 _23740_ (.A0(_03378_),
    .A1(_03382_),
    .S(net122),
    .X(_00318_));
 sg13g2_inv_1 _23741_ (.Y(_03383_),
    .A(_03867_));
 sg13g2_nor2_1 _23742_ (.A(_06932_),
    .B(_03065_),
    .Y(_03384_));
 sg13g2_a21oi_1 _23743_ (.A1(_03383_),
    .A2(_03384_),
    .Y(_03385_),
    .B1(_10723_));
 sg13g2_nand2_1 _23744_ (.Y(_03386_),
    .A(_03383_),
    .B(_03163_));
 sg13g2_a21oi_1 _23745_ (.A1(_03166_),
    .A2(_10192_),
    .Y(_03387_),
    .B1(_03385_));
 sg13g2_o21ai_1 _23746_ (.B1(_03169_),
    .Y(_03388_),
    .A1(_03386_),
    .A2(_03387_));
 sg13g2_o21ai_1 _23747_ (.B1(_03388_),
    .Y(_00319_),
    .A1(_03318_),
    .A2(_03385_));
 sg13g2_nand2_1 _23748_ (.Y(_03389_),
    .A(net140),
    .B(_04644_));
 sg13g2_o21ai_1 _23749_ (.B1(\b.gen_square[50].sq.mask ),
    .Y(_03391_),
    .A1(_03877_),
    .A2(_03389_));
 sg13g2_nand3_1 _23750_ (.B(_04644_),
    .C(net213),
    .A(_04638_),
    .Y(_03392_));
 sg13g2_o21ai_1 _23751_ (.B1(_03392_),
    .Y(_03393_),
    .A1(net188),
    .A2(_03391_));
 sg13g2_inv_1 _23752_ (.Y(_03394_),
    .A(_03877_));
 sg13g2_a21oi_1 _23753_ (.A1(_03393_),
    .A2(_03394_),
    .Y(_03395_),
    .B1(net211));
 sg13g2_mux2_1 _23754_ (.A0(_03391_),
    .A1(_03395_),
    .S(net122),
    .X(_00320_));
 sg13g2_nand2_1 _23755_ (.Y(_03396_),
    .A(net140),
    .B(_04665_));
 sg13g2_o21ai_1 _23756_ (.B1(_06852_),
    .Y(_03397_),
    .A1(_03885_),
    .A2(_03396_));
 sg13g2_nand3_1 _23757_ (.B(_04665_),
    .C(net213),
    .A(_04663_),
    .Y(_03398_));
 sg13g2_o21ai_1 _23758_ (.B1(_03398_),
    .Y(_03399_),
    .A1(net188),
    .A2(_03397_));
 sg13g2_inv_1 _23759_ (.Y(_03401_),
    .A(_03885_));
 sg13g2_a21oi_1 _23760_ (.A1(_03399_),
    .A2(_03401_),
    .Y(_03402_),
    .B1(net211));
 sg13g2_mux2_1 _23761_ (.A0(_03397_),
    .A1(_03402_),
    .S(net122),
    .X(_00321_));
 sg13g2_nand2_1 _23762_ (.Y(_03403_),
    .A(net156),
    .B(_04689_));
 sg13g2_o21ai_1 _23763_ (.B1(\b.gen_square[52].sq.mask ),
    .Y(_03404_),
    .A1(_03403_),
    .A2(_03893_));
 sg13g2_nand3_1 _23764_ (.B(_04689_),
    .C(net213),
    .A(_04687_),
    .Y(_03405_));
 sg13g2_o21ai_1 _23765_ (.B1(_03405_),
    .Y(_03406_),
    .A1(net188),
    .A2(_03404_));
 sg13g2_inv_1 _23766_ (.Y(_03407_),
    .A(_03893_));
 sg13g2_a21oi_1 _23767_ (.A1(_03406_),
    .A2(_03407_),
    .Y(_03408_),
    .B1(net211));
 sg13g2_mux2_1 _23768_ (.A0(_03404_),
    .A1(_03408_),
    .S(net124),
    .X(_00322_));
 sg13g2_nand3_1 _23769_ (.B(net178),
    .C(net139),
    .A(_04712_),
    .Y(_03410_));
 sg13g2_nand2_1 _23770_ (.Y(_03411_),
    .A(_03410_),
    .B(_07292_));
 sg13g2_nand3_1 _23771_ (.B(net178),
    .C(net213),
    .A(_04711_),
    .Y(_03412_));
 sg13g2_o21ai_1 _23772_ (.B1(_03412_),
    .Y(_03413_),
    .A1(net188),
    .A2(_03411_));
 sg13g2_a21oi_1 _23773_ (.A1(_03413_),
    .A2(_04712_),
    .Y(_03414_),
    .B1(net211));
 sg13g2_mux2_1 _23774_ (.A0(_03411_),
    .A1(_03414_),
    .S(net124),
    .X(_00323_));
 sg13g2_nand2_1 _23775_ (.Y(_03415_),
    .A(_03592_),
    .B(_03902_));
 sg13g2_nand3_1 _23776_ (.B(net180),
    .C(net139),
    .A(_03415_),
    .Y(_03416_));
 sg13g2_nand2_1 _23777_ (.Y(_03417_),
    .A(_03416_),
    .B(_05120_));
 sg13g2_nand3_1 _23778_ (.B(net180),
    .C(_03165_),
    .A(_05037_),
    .Y(_03418_));
 sg13g2_o21ai_1 _23779_ (.B1(_03418_),
    .Y(_03420_),
    .A1(net188),
    .A2(_03417_));
 sg13g2_a21oi_1 _23780_ (.A1(_03420_),
    .A2(_03415_),
    .Y(_03421_),
    .B1(net211));
 sg13g2_mux2_1 _23781_ (.A0(_03417_),
    .A1(_03421_),
    .S(net124),
    .X(_00324_));
 sg13g2_inv_1 _23782_ (.Y(_03422_),
    .A(_03917_));
 sg13g2_nor2_1 _23783_ (.A(_04343_),
    .B(net141),
    .Y(_03423_));
 sg13g2_a21oi_1 _23784_ (.A1(_03422_),
    .A2(_03423_),
    .Y(_03424_),
    .B1(_07647_));
 sg13g2_inv_1 _23785_ (.Y(_03425_),
    .A(_03424_));
 sg13g2_o21ai_1 _23786_ (.B1(_03425_),
    .Y(_03426_),
    .A1(net209),
    .A2(_07661_));
 sg13g2_nand3_1 _23787_ (.B(_03422_),
    .C(net157),
    .A(_03426_),
    .Y(_03427_));
 sg13g2_nand2_1 _23788_ (.Y(_03428_),
    .A(_03427_),
    .B(net110));
 sg13g2_o21ai_1 _23789_ (.B1(_03428_),
    .Y(_00325_),
    .A1(net104),
    .A2(_03424_));
 sg13g2_nor2_1 _23790_ (.A(_05441_),
    .B(net107),
    .Y(_03430_));
 sg13g2_inv_1 _23791_ (.Y(_03431_),
    .A(_03927_));
 sg13g2_a21oi_1 _23792_ (.A1(_03430_),
    .A2(_03431_),
    .Y(_03432_),
    .B1(_02377_));
 sg13g2_nand2_1 _23793_ (.Y(_03433_),
    .A(_03431_),
    .B(net155));
 sg13g2_nand3_1 _23794_ (.B(_05263_),
    .C(net213),
    .A(_02347_),
    .Y(_03434_));
 sg13g2_nor2b_1 _23795_ (.A(_03432_),
    .B_N(_03434_),
    .Y(_03435_));
 sg13g2_o21ai_1 _23796_ (.B1(net106),
    .Y(_03436_),
    .A1(_03433_),
    .A2(_03435_));
 sg13g2_o21ai_1 _23797_ (.B1(_03436_),
    .Y(_00326_),
    .A1(net104),
    .A2(_03432_));
 sg13g2_nor2_1 _23798_ (.A(_02284_),
    .B(net141),
    .Y(_03437_));
 sg13g2_nand2_1 _23799_ (.Y(_03439_),
    .A(_03623_),
    .B(net169));
 sg13g2_a21oi_1 _23800_ (.A1(_03437_),
    .A2(_03439_),
    .Y(_03440_),
    .B1(_02265_));
 sg13g2_inv_1 _23801_ (.Y(_03441_),
    .A(_03440_));
 sg13g2_o21ai_1 _23802_ (.B1(_03441_),
    .Y(_03442_),
    .A1(net209),
    .A2(_02302_));
 sg13g2_nand3_1 _23803_ (.B(_03439_),
    .C(net157),
    .A(_03442_),
    .Y(_03443_));
 sg13g2_nand2_1 _23804_ (.Y(_03444_),
    .A(_03443_),
    .B(net110));
 sg13g2_o21ai_1 _23805_ (.B1(_03444_),
    .Y(_00327_),
    .A1(net104),
    .A2(_03440_));
 sg13g2_nor2_1 _23806_ (.A(_05482_),
    .B(net107),
    .Y(_03445_));
 sg13g2_a21oi_1 _23807_ (.A1(_03445_),
    .A2(_03942_),
    .Y(_03446_),
    .B1(_02419_));
 sg13g2_nand2_1 _23808_ (.Y(_03447_),
    .A(_03942_),
    .B(net175));
 sg13g2_a21oi_1 _23809_ (.A1(net187),
    .A2(_02465_),
    .Y(_03448_),
    .B1(_03446_));
 sg13g2_o21ai_1 _23810_ (.B1(net123),
    .Y(_03449_),
    .A1(_03447_),
    .A2(_03448_));
 sg13g2_o21ai_1 _23811_ (.B1(_03449_),
    .Y(_00328_),
    .A1(net104),
    .A2(_03446_));
 sg13g2_inv_1 _23812_ (.Y(_03450_),
    .A(_03951_));
 sg13g2_nor2_1 _23813_ (.A(_06254_),
    .B(net125),
    .Y(_03451_));
 sg13g2_a21oi_1 _23814_ (.A1(_03450_),
    .A2(_03451_),
    .Y(_03452_),
    .B1(_02203_));
 sg13g2_nand2_1 _23815_ (.Y(_03453_),
    .A(_03450_),
    .B(net175));
 sg13g2_a21oi_1 _23816_ (.A1(net187),
    .A2(_02258_),
    .Y(_03454_),
    .B1(_03452_));
 sg13g2_o21ai_1 _23817_ (.B1(net123),
    .Y(_03455_),
    .A1(_03453_),
    .A2(_03454_));
 sg13g2_o21ai_1 _23818_ (.B1(_03455_),
    .Y(_00329_),
    .A1(net104),
    .A2(_03452_));
 sg13g2_nor2_1 _23819_ (.A(_07082_),
    .B(_03065_),
    .Y(_03457_));
 sg13g2_a21oi_1 _23820_ (.A1(_03457_),
    .A2(_03960_),
    .Y(_03458_),
    .B1(_10759_));
 sg13g2_nand2_1 _23821_ (.Y(_03459_),
    .A(_03960_),
    .B(net175));
 sg13g2_a21oi_1 _23822_ (.A1(_03166_),
    .A2(_10106_),
    .Y(_03460_),
    .B1(_03458_));
 sg13g2_o21ai_1 _23823_ (.B1(net123),
    .Y(_03461_),
    .A1(_03459_),
    .A2(_03460_));
 sg13g2_o21ai_1 _23824_ (.B1(_03461_),
    .Y(_00330_),
    .A1(_03318_),
    .A2(_03458_));
 sg13g2_nor2_1 _23825_ (.A(_06784_),
    .B(net141),
    .Y(_03462_));
 sg13g2_inv_1 _23826_ (.Y(_03463_),
    .A(_03969_));
 sg13g2_a21oi_1 _23827_ (.A1(_03462_),
    .A2(_03463_),
    .Y(_03464_),
    .B1(_02136_));
 sg13g2_inv_1 _23828_ (.Y(_03465_),
    .A(_03464_));
 sg13g2_o21ai_1 _23829_ (.B1(_03465_),
    .Y(_03466_),
    .A1(net209),
    .A2(_02194_));
 sg13g2_nand3_1 _23830_ (.B(_03463_),
    .C(net157),
    .A(_03466_),
    .Y(_03467_));
 sg13g2_nand2_1 _23831_ (.Y(_03468_),
    .A(_03467_),
    .B(net110));
 sg13g2_o21ai_1 _23832_ (.B1(_03468_),
    .Y(_00331_),
    .A1(net109),
    .A2(_03464_));
 sg13g2_inv_1 _23833_ (.Y(_03469_),
    .A(_03977_));
 sg13g2_nor2_1 _23834_ (.A(_04362_),
    .B(net125),
    .Y(_03470_));
 sg13g2_a21oi_1 _23835_ (.A1(_03469_),
    .A2(_03470_),
    .Y(_03471_),
    .B1(_02065_));
 sg13g2_nand2_1 _23836_ (.Y(_03472_),
    .A(_03469_),
    .B(net175));
 sg13g2_a21oi_1 _23837_ (.A1(net187),
    .A2(_02129_),
    .Y(_03473_),
    .B1(_03471_));
 sg13g2_o21ai_1 _23838_ (.B1(net123),
    .Y(_03474_),
    .A1(_03472_),
    .A2(_03473_));
 sg13g2_o21ai_1 _23839_ (.B1(_03474_),
    .Y(_00332_),
    .A1(net109),
    .A2(_03471_));
 sg13g2_nor2_1 _23840_ (.A(_04452_),
    .B(net141),
    .Y(_03476_));
 sg13g2_inv_1 _23841_ (.Y(_03477_),
    .A(_03986_));
 sg13g2_a21oi_1 _23842_ (.A1(_03476_),
    .A2(_03477_),
    .Y(_03478_),
    .B1(_02603_));
 sg13g2_inv_1 _23843_ (.Y(_03479_),
    .A(_03478_));
 sg13g2_o21ai_1 _23844_ (.B1(_03479_),
    .Y(_03480_),
    .A1(_01653_),
    .A2(_02629_));
 sg13g2_nand3_1 _23845_ (.B(_03477_),
    .C(net157),
    .A(_03480_),
    .Y(_03481_));
 sg13g2_nand2_1 _23846_ (.Y(_03482_),
    .A(_03481_),
    .B(net110));
 sg13g2_o21ai_1 _23847_ (.B1(_03482_),
    .Y(_00333_),
    .A1(net109),
    .A2(_03478_));
 sg13g2_inv_1 _23848_ (.Y(_03483_),
    .A(_03994_));
 sg13g2_nor2_1 _23849_ (.A(_04427_),
    .B(net125),
    .Y(_03484_));
 sg13g2_a21oi_1 _23850_ (.A1(_03483_),
    .A2(_03484_),
    .Y(_03485_),
    .B1(_02062_));
 sg13g2_nand2_1 _23851_ (.Y(_03486_),
    .A(_03483_),
    .B(net175));
 sg13g2_a21oi_1 _23852_ (.A1(_03092_),
    .A2(_07552_),
    .Y(_03487_),
    .B1(_03485_));
 sg13g2_o21ai_1 _23853_ (.B1(net123),
    .Y(_03488_),
    .A1(_03486_),
    .A2(_03487_));
 sg13g2_o21ai_1 _23854_ (.B1(_03488_),
    .Y(_00334_),
    .A1(net109),
    .A2(_03485_));
 sg13g2_nor2_1 _23855_ (.A(_05865_),
    .B(_03064_),
    .Y(_03489_));
 sg13g2_nand2_1 _23856_ (.Y(_03490_),
    .A(_03592_),
    .B(_01814_));
 sg13g2_inv_1 _23857_ (.Y(_03491_),
    .A(_10824_));
 sg13g2_a21oi_1 _23858_ (.A1(_03489_),
    .A2(_03490_),
    .Y(_03492_),
    .B1(_03491_));
 sg13g2_inv_1 _23859_ (.Y(_03494_),
    .A(_03492_));
 sg13g2_o21ai_1 _23860_ (.B1(_03494_),
    .Y(_03495_),
    .A1(_01653_),
    .A2(_10804_));
 sg13g2_nand3_1 _23861_ (.B(_03490_),
    .C(net155),
    .A(_03495_),
    .Y(_03496_));
 sg13g2_nand2_1 _23862_ (.Y(_03497_),
    .A(_03496_),
    .B(net106));
 sg13g2_o21ai_1 _23863_ (.B1(_03497_),
    .Y(_00335_),
    .A1(net109),
    .A2(_03492_));
 sg13g2_inv_1 _23864_ (.Y(_03498_),
    .A(_04011_));
 sg13g2_nor2_1 _23865_ (.A(_10881_),
    .B(_03159_),
    .Y(_03499_));
 sg13g2_a21oi_1 _23866_ (.A1(_03498_),
    .A2(_03499_),
    .Y(_03500_),
    .B1(_10928_));
 sg13g2_nand2_1 _23867_ (.Y(_03501_),
    .A(_03498_),
    .B(_03071_));
 sg13g2_nor3_1 _23868_ (.A(_01653_),
    .B(_05518_),
    .C(_10881_),
    .Y(_03502_));
 sg13g2_nor2_1 _23869_ (.A(_03502_),
    .B(_03500_),
    .Y(_03503_));
 sg13g2_o21ai_1 _23870_ (.B1(net123),
    .Y(_03504_),
    .A1(_03501_),
    .A2(_03503_));
 sg13g2_o21ai_1 _23871_ (.B1(_03504_),
    .Y(_00336_),
    .A1(_03096_),
    .A2(_03500_));
 sg13g2_nor2_1 _23872_ (.A(_06001_),
    .B(net107),
    .Y(_03505_));
 sg13g2_inv_1 _23873_ (.Y(_03506_),
    .A(_04019_));
 sg13g2_a21oi_1 _23874_ (.A1(_03505_),
    .A2(_03506_),
    .Y(_03507_),
    .B1(_09333_));
 sg13g2_nand2_1 _23875_ (.Y(_03508_),
    .A(_03506_),
    .B(_03071_));
 sg13g2_nor3_1 _23876_ (.A(_01653_),
    .B(_05984_),
    .C(_06001_),
    .Y(_03509_));
 sg13g2_nor2_1 _23877_ (.A(_03509_),
    .B(_03507_),
    .Y(_03510_));
 sg13g2_o21ai_1 _23878_ (.B1(_03082_),
    .Y(_03511_),
    .A1(_03508_),
    .A2(_03510_));
 sg13g2_o21ai_1 _23879_ (.B1(_03511_),
    .Y(_00337_),
    .A1(_03096_),
    .A2(_03507_));
 sg13g2_nand2_1 _23880_ (.Y(_03513_),
    .A(net156),
    .B(net132));
 sg13g2_o21ai_1 _23881_ (.B1(_09461_),
    .Y(_03514_),
    .A1(_03513_),
    .A2(_04028_));
 sg13g2_nand3_1 _23882_ (.B(net132),
    .C(_03165_),
    .A(_04823_),
    .Y(_03515_));
 sg13g2_o21ai_1 _23883_ (.B1(_03515_),
    .Y(_03516_),
    .A1(net188),
    .A2(_03514_));
 sg13g2_a21oi_1 _23884_ (.A1(_03516_),
    .A2(_04027_),
    .Y(_03517_),
    .B1(_03177_));
 sg13g2_mux2_1 _23885_ (.A0(_03514_),
    .A1(_03517_),
    .S(_03074_),
    .X(_00338_));
 sg13g2_a21oi_1 _23886_ (.A1(_00805_),
    .A2(_01492_),
    .Y(_03518_),
    .B1(_03051_));
 sg13g2_nand2_1 _23887_ (.Y(_03519_),
    .A(_00838_),
    .B(_00926_));
 sg13g2_nand3_1 _23888_ (.B(_03519_),
    .C(_01417_),
    .A(_03518_),
    .Y(_03520_));
 sg13g2_o21ai_1 _23889_ (.B1(_00772_),
    .Y(_03522_),
    .A1(_01351_),
    .A2(_01373_));
 sg13g2_nand4_1 _23890_ (.B(_03001_),
    .C(_01111_),
    .A(_03520_),
    .Y(_03523_),
    .D(_03522_));
 sg13g2_a21oi_1 _23891_ (.A1(\state[10] ),
    .A2(_01198_),
    .Y(_00339_),
    .B1(_03523_));
 sg13g2_nand3_1 _23892_ (.B(data_out_valid),
    .C(_01013_),
    .A(_01002_),
    .Y(_03524_));
 sg13g2_buf_1 _23893_ (.A(_03524_),
    .X(_03525_));
 sg13g2_nor2b_1 _23894_ (.A(_03525_),
    .B_N(\data_out[0] ),
    .Y(net8));
 sg13g2_nor2b_1 _23895_ (.A(_03525_),
    .B_N(\data_out[1] ),
    .Y(net9));
 sg13g2_nor2b_1 _23896_ (.A(_03525_),
    .B_N(\data_out[2] ),
    .Y(net10));
 sg13g2_nor2_1 _23897_ (.A(_02896_),
    .B(_03525_),
    .Y(net11));
 sg13g2_dfrbp_1 _23898_ (.CLK(clknet_leaf_15_clk),
    .RESET_B(net239),
    .D(_00340_),
    .Q_N(_12056_),
    .Q(\state[8] ));
 sg13g2_dfrbp_1 _23899_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net242),
    .D(_00341_),
    .Q_N(_12055_),
    .Q(\state[2] ));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_tiehi \spi.din[0]$_DFFE_PP__313  (.L_HI(net313));
 sg13g2_buf_1 _23902_ (.A(net293),
    .X(uio_oe[0]));
 sg13g2_buf_1 _23903_ (.A(net294),
    .X(uio_oe[1]));
 sg13g2_buf_1 _23904_ (.A(net295),
    .X(uio_oe[2]));
 sg13g2_buf_1 _23905_ (.A(net296),
    .X(uio_oe[3]));
 sg13g2_buf_1 _23906_ (.A(net297),
    .X(uio_oe[4]));
 sg13g2_buf_1 _23907_ (.A(net298),
    .X(uio_oe[5]));
 sg13g2_buf_1 _23908_ (.A(net299),
    .X(uio_oe[6]));
 sg13g2_buf_1 _23909_ (.A(net300),
    .X(uio_oe[7]));
 sg13g2_buf_1 _23910_ (.A(net301),
    .X(uio_out[0]));
 sg13g2_buf_1 _23911_ (.A(net302),
    .X(uio_out[1]));
 sg13g2_buf_1 _23912_ (.A(net303),
    .X(uio_out[2]));
 sg13g2_buf_1 _23913_ (.A(net304),
    .X(uio_out[3]));
 sg13g2_buf_1 _23914_ (.A(net305),
    .X(uio_out[4]));
 sg13g2_buf_1 _23915_ (.A(net306),
    .X(uio_out[5]));
 sg13g2_buf_1 _23916_ (.A(net307),
    .X(uio_out[6]));
 sg13g2_buf_1 _23917_ (.A(net308),
    .X(uio_out[7]));
 sg13g2_buf_1 _23918_ (.A(net309),
    .X(uo_out[0]));
 sg13g2_buf_1 _23919_ (.A(net310),
    .X(uo_out[1]));
 sg13g2_buf_1 _23920_ (.A(net311),
    .X(uo_out[2]));
 sg13g2_buf_1 _23921_ (.A(net312),
    .X(uo_out[3]));
 sg13g2_dfrbp_1 \b.gen_square[0].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net279),
    .D(_00342_),
    .Q_N(_12054_),
    .Q(\b.gen_square[0].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[0].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net280),
    .D(_00275_),
    .Q_N(\b.gen_square[0].sq.mask ),
    .Q(_12066_));
 sg13g2_dfrbp_1 \b.gen_square[0].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net280),
    .D(_00343_),
    .Q_N(\b.gen_square[0].sq.piece[0] ),
    .Q(_00081_));
 sg13g2_dfrbp_1 \b.gen_square[0].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net280),
    .D(_00344_),
    .Q_N(\b.gen_square[0].sq.piece[1] ),
    .Q(_00082_));
 sg13g2_dfrbp_1 \b.gen_square[0].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net280),
    .D(_00345_),
    .Q_N(\b.gen_square[0].sq.piece[2] ),
    .Q(_00083_));
 sg13g2_dfrbp_1 \b.gen_square[10].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net283),
    .D(_00346_),
    .Q_N(_00063_),
    .Q(\b.gen_square[10].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[10].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net283),
    .D(_00276_),
    .Q_N(\b.gen_square[10].sq.mask ),
    .Q(_12067_));
 sg13g2_dfrbp_1 \b.gen_square[10].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net282),
    .D(_00347_),
    .Q_N(\b.gen_square[10].sq.piece[0] ),
    .Q(_00084_));
 sg13g2_dfrbp_1 \b.gen_square[10].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net282),
    .D(_00348_),
    .Q_N(\b.gen_square[10].sq.piece[1] ),
    .Q(_00085_));
 sg13g2_dfrbp_1 \b.gen_square[10].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net282),
    .D(_00349_),
    .Q_N(\b.gen_square[10].sq.piece[2] ),
    .Q(_00086_));
 sg13g2_dfrbp_1 \b.gen_square[11].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net283),
    .D(_00350_),
    .Q_N(_00060_),
    .Q(\b.gen_square[11].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[11].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net281),
    .D(_00277_),
    .Q_N(\b.gen_square[11].sq.mask ),
    .Q(_12068_));
 sg13g2_dfrbp_1 \b.gen_square[11].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net281),
    .D(_00351_),
    .Q_N(\b.gen_square[11].sq.piece[0] ),
    .Q(_00087_));
 sg13g2_dfrbp_1 \b.gen_square[11].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net281),
    .D(_00352_),
    .Q_N(\b.gen_square[11].sq.piece[1] ),
    .Q(_00088_));
 sg13g2_dfrbp_1 \b.gen_square[11].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net281),
    .D(_00353_),
    .Q_N(\b.gen_square[11].sq.piece[2] ),
    .Q(_00089_));
 sg13g2_dfrbp_1 \b.gen_square[12].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net288),
    .D(_00354_),
    .Q_N(_00054_),
    .Q(\b.gen_square[12].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[12].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net287),
    .D(_00278_),
    .Q_N(\b.gen_square[12].sq.mask ),
    .Q(_12069_));
 sg13g2_dfrbp_1 \b.gen_square[12].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net287),
    .D(_00355_),
    .Q_N(\b.gen_square[12].sq.piece[0] ),
    .Q(_00090_));
 sg13g2_dfrbp_1 \b.gen_square[12].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net287),
    .D(_00356_),
    .Q_N(\b.gen_square[12].sq.piece[1] ),
    .Q(_00091_));
 sg13g2_dfrbp_1 \b.gen_square[12].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net287),
    .D(_00357_),
    .Q_N(\b.gen_square[12].sq.piece[2] ),
    .Q(_00092_));
 sg13g2_dfrbp_1 \b.gen_square[13].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net289),
    .D(_00358_),
    .Q_N(_00047_),
    .Q(\b.gen_square[13].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[13].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net289),
    .D(_00279_),
    .Q_N(\b.gen_square[13].sq.mask ),
    .Q(_12070_));
 sg13g2_dfrbp_1 \b.gen_square[13].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net289),
    .D(_00359_),
    .Q_N(\b.gen_square[13].sq.piece[0] ),
    .Q(_00093_));
 sg13g2_dfrbp_1 \b.gen_square[13].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net289),
    .D(_00360_),
    .Q_N(\b.gen_square[13].sq.piece[1] ),
    .Q(_00094_));
 sg13g2_dfrbp_1 \b.gen_square[13].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net289),
    .D(_00361_),
    .Q_N(\b.gen_square[13].sq.piece[2] ),
    .Q(_00095_));
 sg13g2_dfrbp_1 \b.gen_square[14].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net285),
    .D(_00362_),
    .Q_N(_00038_),
    .Q(\b.gen_square[14].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[14].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net285),
    .D(_00280_),
    .Q_N(\b.gen_square[14].sq.mask ),
    .Q(_12071_));
 sg13g2_dfrbp_1 \b.gen_square[14].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net289),
    .D(_00363_),
    .Q_N(\b.gen_square[14].sq.piece[0] ),
    .Q(_00096_));
 sg13g2_dfrbp_1 \b.gen_square[14].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net290),
    .D(_00364_),
    .Q_N(\b.gen_square[14].sq.piece[1] ),
    .Q(_00097_));
 sg13g2_dfrbp_1 \b.gen_square[14].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net290),
    .D(_00365_),
    .Q_N(\b.gen_square[14].sq.piece[2] ),
    .Q(_00098_));
 sg13g2_dfrbp_1 \b.gen_square[15].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net277),
    .D(_00366_),
    .Q_N(_00019_),
    .Q(\b.gen_square[15].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[15].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net285),
    .D(_00281_),
    .Q_N(\b.gen_square[15].sq.mask ),
    .Q(_12072_));
 sg13g2_dfrbp_1 \b.gen_square[15].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net290),
    .D(_00367_),
    .Q_N(\b.gen_square[15].sq.piece[0] ),
    .Q(_00099_));
 sg13g2_dfrbp_1 \b.gen_square[15].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net288),
    .D(_00368_),
    .Q_N(\b.gen_square[15].sq.piece[1] ),
    .Q(_00100_));
 sg13g2_dfrbp_1 \b.gen_square[15].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net290),
    .D(_00369_),
    .Q_N(\b.gen_square[15].sq.piece[2] ),
    .Q(_00101_));
 sg13g2_dfrbp_1 \b.gen_square[16].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net267),
    .D(_00370_),
    .Q_N(_00065_),
    .Q(\b.gen_square[16].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[16].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net268),
    .D(_00282_),
    .Q_N(\b.gen_square[16].sq.mask ),
    .Q(_12073_));
 sg13g2_dfrbp_1 \b.gen_square[16].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net279),
    .D(_00371_),
    .Q_N(\b.gen_square[16].sq.piece[0] ),
    .Q(_00102_));
 sg13g2_dfrbp_1 \b.gen_square[16].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net278),
    .D(_00372_),
    .Q_N(\b.gen_square[16].sq.piece[1] ),
    .Q(_00103_));
 sg13g2_dfrbp_1 \b.gen_square[16].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net279),
    .D(_00373_),
    .Q_N(\b.gen_square[16].sq.piece[2] ),
    .Q(_00104_));
 sg13g2_dfrbp_1 \b.gen_square[17].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net268),
    .D(_00374_),
    .Q_N(_00032_),
    .Q(\b.gen_square[17].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[17].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net278),
    .D(_00283_),
    .Q_N(\b.gen_square[17].sq.mask ),
    .Q(_12074_));
 sg13g2_dfrbp_1 \b.gen_square[17].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net278),
    .D(_00375_),
    .Q_N(\b.gen_square[17].sq.piece[0] ),
    .Q(_00105_));
 sg13g2_dfrbp_1 \b.gen_square[17].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net278),
    .D(_00376_),
    .Q_N(\b.gen_square[17].sq.piece[1] ),
    .Q(_00106_));
 sg13g2_dfrbp_1 \b.gen_square[17].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net279),
    .D(_00377_),
    .Q_N(\b.gen_square[17].sq.piece[2] ),
    .Q(_00107_));
 sg13g2_dfrbp_1 \b.gen_square[18].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net269),
    .D(_00378_),
    .Q_N(_00075_),
    .Q(\b.gen_square[18].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[18].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net267),
    .D(_00284_),
    .Q_N(\b.gen_square[18].sq.mask ),
    .Q(_12075_));
 sg13g2_dfrbp_1 \b.gen_square[18].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net268),
    .D(_00379_),
    .Q_N(\b.gen_square[18].sq.piece[0] ),
    .Q(_00108_));
 sg13g2_dfrbp_1 \b.gen_square[18].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net267),
    .D(_00380_),
    .Q_N(\b.gen_square[18].sq.piece[1] ),
    .Q(_00109_));
 sg13g2_dfrbp_1 \b.gen_square[18].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net268),
    .D(_00381_),
    .Q_N(\b.gen_square[18].sq.piece[2] ),
    .Q(_00110_));
 sg13g2_dfrbp_1 \b.gen_square[19].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net269),
    .D(_00382_),
    .Q_N(_00059_),
    .Q(\b.gen_square[19].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[19].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net285),
    .D(_00285_),
    .Q_N(\b.gen_square[19].sq.mask ),
    .Q(_12076_));
 sg13g2_dfrbp_1 \b.gen_square[19].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net286),
    .D(_00383_),
    .Q_N(\b.gen_square[19].sq.piece[0] ),
    .Q(_00111_));
 sg13g2_dfrbp_1 \b.gen_square[19].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net286),
    .D(_00384_),
    .Q_N(\b.gen_square[19].sq.piece[1] ),
    .Q(_00112_));
 sg13g2_dfrbp_1 \b.gen_square[19].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net286),
    .D(_00385_),
    .Q_N(\b.gen_square[19].sq.piece[2] ),
    .Q(_00113_));
 sg13g2_dfrbp_1 \b.gen_square[1].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net278),
    .D(_00386_),
    .Q_N(_00014_),
    .Q(\b.gen_square[1].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[1].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net279),
    .D(_00286_),
    .Q_N(\b.gen_square[1].sq.mask ),
    .Q(_12077_));
 sg13g2_dfrbp_1 \b.gen_square[1].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net278),
    .D(_00387_),
    .Q_N(\b.gen_square[1].sq.piece[0] ),
    .Q(_00114_));
 sg13g2_dfrbp_1 \b.gen_square[1].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net278),
    .D(_00388_),
    .Q_N(\b.gen_square[1].sq.piece[1] ),
    .Q(_00115_));
 sg13g2_dfrbp_1 \b.gen_square[1].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net278),
    .D(_00389_),
    .Q_N(\b.gen_square[1].sq.piece[2] ),
    .Q(_00116_));
 sg13g2_dfrbp_1 \b.gen_square[20].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net269),
    .D(_00390_),
    .Q_N(_00053_),
    .Q(\b.gen_square[20].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[20].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net269),
    .D(_00287_),
    .Q_N(\b.gen_square[20].sq.mask ),
    .Q(_12078_));
 sg13g2_dfrbp_1 \b.gen_square[20].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net276),
    .D(_00391_),
    .Q_N(\b.gen_square[20].sq.piece[0] ),
    .Q(_00117_));
 sg13g2_dfrbp_1 \b.gen_square[20].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net275),
    .D(_00392_),
    .Q_N(\b.gen_square[20].sq.piece[1] ),
    .Q(_00118_));
 sg13g2_dfrbp_1 \b.gen_square[20].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net276),
    .D(_00393_),
    .Q_N(\b.gen_square[20].sq.piece[2] ),
    .Q(_00119_));
 sg13g2_dfrbp_1 \b.gen_square[21].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net277),
    .D(_00394_),
    .Q_N(_00046_),
    .Q(\b.gen_square[21].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[21].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net277),
    .D(_00288_),
    .Q_N(\b.gen_square[21].sq.mask ),
    .Q(_12079_));
 sg13g2_dfrbp_1 \b.gen_square[21].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net275),
    .D(_00395_),
    .Q_N(\b.gen_square[21].sq.piece[0] ),
    .Q(_00120_));
 sg13g2_dfrbp_1 \b.gen_square[21].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net275),
    .D(_00396_),
    .Q_N(\b.gen_square[21].sq.piece[1] ),
    .Q(_00121_));
 sg13g2_dfrbp_1 \b.gen_square[21].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net275),
    .D(_00397_),
    .Q_N(\b.gen_square[21].sq.piece[2] ),
    .Q(_00122_));
 sg13g2_dfrbp_1 \b.gen_square[22].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net276),
    .D(_00398_),
    .Q_N(_00037_),
    .Q(\b.gen_square[22].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[22].sq.mask$_DFF_PN1_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net275),
    .D(_00289_),
    .Q_N(\b.gen_square[22].sq.mask ),
    .Q(_12080_));
 sg13g2_dfrbp_1 \b.gen_square[22].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net275),
    .D(_00399_),
    .Q_N(\b.gen_square[22].sq.piece[0] ),
    .Q(_00123_));
 sg13g2_dfrbp_1 \b.gen_square[22].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net275),
    .D(_00400_),
    .Q_N(\b.gen_square[22].sq.piece[1] ),
    .Q(_00124_));
 sg13g2_dfrbp_1 \b.gen_square[22].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net276),
    .D(_00401_),
    .Q_N(\b.gen_square[22].sq.piece[2] ),
    .Q(_00125_));
 sg13g2_dfrbp_1 \b.gen_square[23].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net272),
    .D(_00402_),
    .Q_N(_00018_),
    .Q(\b.gen_square[23].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[23].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net272),
    .D(_00290_),
    .Q_N(\b.gen_square[23].sq.mask ),
    .Q(_12081_));
 sg13g2_dfrbp_1 \b.gen_square[23].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net272),
    .D(_00403_),
    .Q_N(\b.gen_square[23].sq.piece[0] ),
    .Q(_00126_));
 sg13g2_dfrbp_1 \b.gen_square[23].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net272),
    .D(_00404_),
    .Q_N(\b.gen_square[23].sq.piece[1] ),
    .Q(_00127_));
 sg13g2_dfrbp_1 \b.gen_square[23].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net272),
    .D(_00405_),
    .Q_N(\b.gen_square[23].sq.piece[2] ),
    .Q(_00128_));
 sg13g2_dfrbp_1 \b.gen_square[24].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net267),
    .D(_00406_),
    .Q_N(_00064_),
    .Q(\b.gen_square[24].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[24].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net267),
    .D(_00291_),
    .Q_N(\b.gen_square[24].sq.mask ),
    .Q(_12082_));
 sg13g2_dfrbp_1 \b.gen_square[24].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net267),
    .D(_00407_),
    .Q_N(\b.gen_square[24].sq.piece[0] ),
    .Q(_00129_));
 sg13g2_dfrbp_1 \b.gen_square[24].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net267),
    .D(_00408_),
    .Q_N(\b.gen_square[24].sq.piece[1] ),
    .Q(_00130_));
 sg13g2_dfrbp_1 \b.gen_square[24].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net267),
    .D(_00409_),
    .Q_N(\b.gen_square[24].sq.piece[2] ),
    .Q(_00131_));
 sg13g2_dfrbp_1 \b.gen_square[25].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net264),
    .D(_00410_),
    .Q_N(_00043_),
    .Q(\b.gen_square[25].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[25].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net264),
    .D(_00292_),
    .Q_N(\b.gen_square[25].sq.mask ),
    .Q(_12083_));
 sg13g2_dfrbp_1 \b.gen_square[25].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net264),
    .D(_00411_),
    .Q_N(\b.gen_square[25].sq.piece[0] ),
    .Q(_00132_));
 sg13g2_dfrbp_1 \b.gen_square[25].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net264),
    .D(_00412_),
    .Q_N(\b.gen_square[25].sq.piece[1] ),
    .Q(_00133_));
 sg13g2_dfrbp_1 \b.gen_square[25].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net264),
    .D(_00413_),
    .Q_N(\b.gen_square[25].sq.piece[2] ),
    .Q(_00134_));
 sg13g2_dfrbp_1 \b.gen_square[26].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net266),
    .D(_00414_),
    .Q_N(_00031_),
    .Q(\b.gen_square[26].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[26].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net265),
    .D(_00293_),
    .Q_N(\b.gen_square[26].sq.mask ),
    .Q(_12084_));
 sg13g2_dfrbp_1 \b.gen_square[26].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net263),
    .D(_00415_),
    .Q_N(\b.gen_square[26].sq.piece[0] ),
    .Q(_00135_));
 sg13g2_dfrbp_1 \b.gen_square[26].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net264),
    .D(_00416_),
    .Q_N(\b.gen_square[26].sq.piece[1] ),
    .Q(_00136_));
 sg13g2_dfrbp_1 \b.gen_square[26].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net264),
    .D(_00417_),
    .Q_N(\b.gen_square[26].sq.piece[2] ),
    .Q(_00137_));
 sg13g2_dfrbp_1 \b.gen_square[27].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net269),
    .D(_00418_),
    .Q_N(_00074_),
    .Q(\b.gen_square[27].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[27].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net265),
    .D(_00294_),
    .Q_N(\b.gen_square[27].sq.mask ),
    .Q(_12085_));
 sg13g2_dfrbp_1 \b.gen_square[27].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net263),
    .D(_00419_),
    .Q_N(\b.gen_square[27].sq.piece[0] ),
    .Q(_00138_));
 sg13g2_dfrbp_1 \b.gen_square[27].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net263),
    .D(_00420_),
    .Q_N(\b.gen_square[27].sq.piece[1] ),
    .Q(_00139_));
 sg13g2_dfrbp_1 \b.gen_square[27].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net263),
    .D(_00421_),
    .Q_N(\b.gen_square[27].sq.piece[2] ),
    .Q(_00140_));
 sg13g2_dfrbp_1 \b.gen_square[28].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net266),
    .D(_00422_),
    .Q_N(_00052_),
    .Q(\b.gen_square[28].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[28].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net274),
    .D(_00295_),
    .Q_N(\b.gen_square[28].sq.mask ),
    .Q(_12086_));
 sg13g2_dfrbp_1 \b.gen_square[28].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net265),
    .D(_00423_),
    .Q_N(\b.gen_square[28].sq.piece[0] ),
    .Q(_00141_));
 sg13g2_dfrbp_1 \b.gen_square[28].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net265),
    .D(_00424_),
    .Q_N(\b.gen_square[28].sq.piece[1] ),
    .Q(_00142_));
 sg13g2_dfrbp_1 \b.gen_square[28].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net265),
    .D(_00425_),
    .Q_N(\b.gen_square[28].sq.piece[2] ),
    .Q(_00143_));
 sg13g2_dfrbp_1 \b.gen_square[29].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net274),
    .D(_00426_),
    .Q_N(_00045_),
    .Q(\b.gen_square[29].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[29].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net274),
    .D(_00296_),
    .Q_N(\b.gen_square[29].sq.mask ),
    .Q(_12087_));
 sg13g2_dfrbp_1 \b.gen_square[29].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net271),
    .D(_00427_),
    .Q_N(\b.gen_square[29].sq.piece[0] ),
    .Q(_00144_));
 sg13g2_dfrbp_1 \b.gen_square[29].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net271),
    .D(_00428_),
    .Q_N(\b.gen_square[29].sq.piece[1] ),
    .Q(_00145_));
 sg13g2_dfrbp_1 \b.gen_square[29].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net271),
    .D(_00429_),
    .Q_N(\b.gen_square[29].sq.piece[2] ),
    .Q(_00146_));
 sg13g2_dfrbp_1 \b.gen_square[2].sq.color$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net284),
    .D(_00430_),
    .Q_N(_00013_),
    .Q(\b.gen_square[2].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[2].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net282),
    .D(_00297_),
    .Q_N(\b.gen_square[2].sq.mask ),
    .Q(_12088_));
 sg13g2_dfrbp_1 \b.gen_square[2].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net280),
    .D(_00431_),
    .Q_N(\b.gen_square[2].sq.piece[0] ),
    .Q(_00147_));
 sg13g2_dfrbp_1 \b.gen_square[2].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net279),
    .D(_00432_),
    .Q_N(\b.gen_square[2].sq.piece[1] ),
    .Q(_00148_));
 sg13g2_dfrbp_1 \b.gen_square[2].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net279),
    .D(_00433_),
    .Q_N(\b.gen_square[2].sq.piece[2] ),
    .Q(_00149_));
 sg13g2_dfrbp_1 \b.gen_square[30].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net274),
    .D(_00434_),
    .Q_N(_00036_),
    .Q(\b.gen_square[30].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[30].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net272),
    .D(_00298_),
    .Q_N(\b.gen_square[30].sq.mask ),
    .Q(_12089_));
 sg13g2_dfrbp_1 \b.gen_square[30].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net272),
    .D(_00435_),
    .Q_N(\b.gen_square[30].sq.piece[0] ),
    .Q(_00150_));
 sg13g2_dfrbp_1 \b.gen_square[30].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net271),
    .D(_00436_),
    .Q_N(\b.gen_square[30].sq.piece[1] ),
    .Q(_00151_));
 sg13g2_dfrbp_1 \b.gen_square[30].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net271),
    .D(_00437_),
    .Q_N(\b.gen_square[30].sq.piece[2] ),
    .Q(_00152_));
 sg13g2_dfrbp_1 \b.gen_square[31].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net260),
    .D(_00438_),
    .Q_N(_00017_),
    .Q(\b.gen_square[31].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[31].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net273),
    .D(_00299_),
    .Q_N(\b.gen_square[31].sq.mask ),
    .Q(_12090_));
 sg13g2_dfrbp_1 \b.gen_square[31].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net271),
    .D(_00439_),
    .Q_N(\b.gen_square[31].sq.piece[0] ),
    .Q(_00153_));
 sg13g2_dfrbp_1 \b.gen_square[31].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net271),
    .D(_00440_),
    .Q_N(\b.gen_square[31].sq.piece[1] ),
    .Q(_00154_));
 sg13g2_dfrbp_1 \b.gen_square[31].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net271),
    .D(_00441_),
    .Q_N(\b.gen_square[31].sq.piece[2] ),
    .Q(_00155_));
 sg13g2_dfrbp_1 \b.gen_square[32].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net253),
    .D(_00442_),
    .Q_N(_00058_),
    .Q(\b.gen_square[32].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[32].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net253),
    .D(_00300_),
    .Q_N(\b.gen_square[32].sq.mask ),
    .Q(_12091_));
 sg13g2_dfrbp_1 \b.gen_square[32].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net254),
    .D(_00443_),
    .Q_N(\b.gen_square[32].sq.piece[0] ),
    .Q(_00156_));
 sg13g2_dfrbp_1 \b.gen_square[32].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net253),
    .D(_00444_),
    .Q_N(\b.gen_square[32].sq.piece[1] ),
    .Q(_00157_));
 sg13g2_dfrbp_1 \b.gen_square[32].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net254),
    .D(_00445_),
    .Q_N(\b.gen_square[32].sq.piece[2] ),
    .Q(_00158_));
 sg13g2_dfrbp_1 \b.gen_square[33].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net263),
    .D(_00446_),
    .Q_N(_00051_),
    .Q(\b.gen_square[33].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[33].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net263),
    .D(_00301_),
    .Q_N(\b.gen_square[33].sq.mask ),
    .Q(_12092_));
 sg13g2_dfrbp_1 \b.gen_square[33].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net254),
    .D(_00447_),
    .Q_N(\b.gen_square[33].sq.piece[0] ),
    .Q(_00159_));
 sg13g2_dfrbp_1 \b.gen_square[33].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net263),
    .D(_00448_),
    .Q_N(\b.gen_square[33].sq.piece[1] ),
    .Q(_00160_));
 sg13g2_dfrbp_1 \b.gen_square[33].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net263),
    .D(_00449_),
    .Q_N(\b.gen_square[33].sq.piece[2] ),
    .Q(_00161_));
 sg13g2_dfrbp_1 \b.gen_square[34].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net254),
    .D(_00450_),
    .Q_N(_00042_),
    .Q(\b.gen_square[34].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[34].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net253),
    .D(_00302_),
    .Q_N(\b.gen_square[34].sq.mask ),
    .Q(_12093_));
 sg13g2_dfrbp_1 \b.gen_square[34].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net253),
    .D(_00451_),
    .Q_N(\b.gen_square[34].sq.piece[0] ),
    .Q(_00162_));
 sg13g2_dfrbp_1 \b.gen_square[34].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net253),
    .D(_00452_),
    .Q_N(\b.gen_square[34].sq.piece[1] ),
    .Q(_00163_));
 sg13g2_dfrbp_1 \b.gen_square[34].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net253),
    .D(_00453_),
    .Q_N(\b.gen_square[34].sq.piece[2] ),
    .Q(_00164_));
 sg13g2_dfrbp_1 \b.gen_square[35].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net265),
    .D(_00454_),
    .Q_N(_00030_),
    .Q(\b.gen_square[35].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[35].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net254),
    .D(_00303_),
    .Q_N(\b.gen_square[35].sq.mask ),
    .Q(_12094_));
 sg13g2_dfrbp_1 \b.gen_square[35].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net265),
    .D(_00455_),
    .Q_N(\b.gen_square[35].sq.piece[0] ),
    .Q(_00165_));
 sg13g2_dfrbp_1 \b.gen_square[35].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net265),
    .D(_00456_),
    .Q_N(\b.gen_square[35].sq.piece[1] ),
    .Q(_00166_));
 sg13g2_dfrbp_1 \b.gen_square[35].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net266),
    .D(_00457_),
    .Q_N(\b.gen_square[35].sq.piece[2] ),
    .Q(_00167_));
 sg13g2_dfrbp_1 \b.gen_square[36].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net254),
    .D(_00458_),
    .Q_N(_00073_),
    .Q(\b.gen_square[36].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[36].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net261),
    .D(_00304_),
    .Q_N(\b.gen_square[36].sq.mask ),
    .Q(_12095_));
 sg13g2_dfrbp_1 \b.gen_square[36].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net254),
    .D(_00459_),
    .Q_N(\b.gen_square[36].sq.piece[0] ),
    .Q(_00168_));
 sg13g2_dfrbp_1 \b.gen_square[36].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net255),
    .D(_00460_),
    .Q_N(\b.gen_square[36].sq.piece[1] ),
    .Q(_00169_));
 sg13g2_dfrbp_1 \b.gen_square[36].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net255),
    .D(_00461_),
    .Q_N(\b.gen_square[36].sq.piece[2] ),
    .Q(_00170_));
 sg13g2_dfrbp_1 \b.gen_square[37].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net261),
    .D(_00462_),
    .Q_N(_00044_),
    .Q(\b.gen_square[37].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[37].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net260),
    .D(_00305_),
    .Q_N(\b.gen_square[37].sq.mask ),
    .Q(_12096_));
 sg13g2_dfrbp_1 \b.gen_square[37].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net260),
    .D(_00463_),
    .Q_N(\b.gen_square[37].sq.piece[0] ),
    .Q(_00171_));
 sg13g2_dfrbp_1 \b.gen_square[37].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net260),
    .D(_00464_),
    .Q_N(\b.gen_square[37].sq.piece[1] ),
    .Q(_00172_));
 sg13g2_dfrbp_1 \b.gen_square[37].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net260),
    .D(_00465_),
    .Q_N(\b.gen_square[37].sq.piece[2] ),
    .Q(_00173_));
 sg13g2_dfrbp_1 \b.gen_square[38].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net261),
    .D(_00466_),
    .Q_N(_00035_),
    .Q(\b.gen_square[38].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[38].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net260),
    .D(_00306_),
    .Q_N(\b.gen_square[38].sq.mask ),
    .Q(_12097_));
 sg13g2_dfrbp_1 \b.gen_square[38].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net259),
    .D(_00467_),
    .Q_N(\b.gen_square[38].sq.piece[0] ),
    .Q(_00174_));
 sg13g2_dfrbp_1 \b.gen_square[38].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net259),
    .D(_00468_),
    .Q_N(\b.gen_square[38].sq.piece[1] ),
    .Q(_00175_));
 sg13g2_dfrbp_1 \b.gen_square[38].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net259),
    .D(_00469_),
    .Q_N(\b.gen_square[38].sq.piece[2] ),
    .Q(_00176_));
 sg13g2_dfrbp_1 \b.gen_square[39].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net256),
    .D(_00470_),
    .Q_N(_00016_),
    .Q(\b.gen_square[39].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[39].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net259),
    .D(_00307_),
    .Q_N(\b.gen_square[39].sq.mask ),
    .Q(_12098_));
 sg13g2_dfrbp_1 \b.gen_square[39].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net257),
    .D(_00471_),
    .Q_N(\b.gen_square[39].sq.piece[0] ),
    .Q(_00177_));
 sg13g2_dfrbp_1 \b.gen_square[39].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net259),
    .D(_00472_),
    .Q_N(\b.gen_square[39].sq.piece[1] ),
    .Q(_00178_));
 sg13g2_dfrbp_1 \b.gen_square[39].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net259),
    .D(_00473_),
    .Q_N(\b.gen_square[39].sq.piece[2] ),
    .Q(_00179_));
 sg13g2_dfrbp_1 \b.gen_square[3].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net285),
    .D(_00474_),
    .Q_N(_00012_),
    .Q(\b.gen_square[3].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[3].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net287),
    .D(_00308_),
    .Q_N(\b.gen_square[3].sq.mask ),
    .Q(_12099_));
 sg13g2_dfrbp_1 \b.gen_square[3].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net287),
    .D(_00475_),
    .Q_N(\b.gen_square[3].sq.piece[0] ),
    .Q(_00180_));
 sg13g2_dfrbp_1 \b.gen_square[3].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net287),
    .D(_00476_),
    .Q_N(\b.gen_square[3].sq.piece[1] ),
    .Q(_00181_));
 sg13g2_dfrbp_1 \b.gen_square[3].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net287),
    .D(_00477_),
    .Q_N(\b.gen_square[3].sq.piece[2] ),
    .Q(_00182_));
 sg13g2_dfrbp_1 \b.gen_square[40].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net250),
    .D(_00478_),
    .Q_N(_00062_),
    .Q(\b.gen_square[40].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[40].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net253),
    .D(_00309_),
    .Q_N(\b.gen_square[40].sq.mask ),
    .Q(_12100_));
 sg13g2_dfrbp_1 \b.gen_square[40].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net250),
    .D(_00479_),
    .Q_N(\b.gen_square[40].sq.piece[0] ),
    .Q(_00183_));
 sg13g2_dfrbp_1 \b.gen_square[40].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net251),
    .D(_00480_),
    .Q_N(\b.gen_square[40].sq.piece[1] ),
    .Q(_00184_));
 sg13g2_dfrbp_1 \b.gen_square[40].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net251),
    .D(_00481_),
    .Q_N(\b.gen_square[40].sq.piece[2] ),
    .Q(_00185_));
 sg13g2_dfrbp_1 \b.gen_square[41].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net250),
    .D(_00482_),
    .Q_N(_00057_),
    .Q(\b.gen_square[41].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[41].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net251),
    .D(_00310_),
    .Q_N(\b.gen_square[41].sq.mask ),
    .Q(_12101_));
 sg13g2_dfrbp_1 \b.gen_square[41].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net250),
    .D(_00483_),
    .Q_N(\b.gen_square[41].sq.piece[0] ),
    .Q(_00186_));
 sg13g2_dfrbp_1 \b.gen_square[41].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net250),
    .D(_00484_),
    .Q_N(\b.gen_square[41].sq.piece[1] ),
    .Q(_00187_));
 sg13g2_dfrbp_1 \b.gen_square[41].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net236),
    .D(_00485_),
    .Q_N(\b.gen_square[41].sq.piece[2] ),
    .Q(_00188_));
 sg13g2_dfrbp_1 \b.gen_square[42].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net255),
    .D(_00486_),
    .Q_N(_00050_),
    .Q(\b.gen_square[42].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[42].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net252),
    .D(_00311_),
    .Q_N(\b.gen_square[42].sq.mask ),
    .Q(_12102_));
 sg13g2_dfrbp_1 \b.gen_square[42].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net251),
    .D(_00487_),
    .Q_N(\b.gen_square[42].sq.piece[0] ),
    .Q(_00189_));
 sg13g2_dfrbp_1 \b.gen_square[42].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net251),
    .D(_00488_),
    .Q_N(\b.gen_square[42].sq.piece[1] ),
    .Q(_00190_));
 sg13g2_dfrbp_1 \b.gen_square[42].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net251),
    .D(_00489_),
    .Q_N(\b.gen_square[42].sq.piece[2] ),
    .Q(_00191_));
 sg13g2_dfrbp_1 \b.gen_square[43].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net252),
    .D(_00490_),
    .Q_N(_00041_),
    .Q(\b.gen_square[43].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[43].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net252),
    .D(_00312_),
    .Q_N(\b.gen_square[43].sq.mask ),
    .Q(_12103_));
 sg13g2_dfrbp_1 \b.gen_square[43].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net236),
    .D(_00491_),
    .Q_N(\b.gen_square[43].sq.piece[0] ),
    .Q(_00192_));
 sg13g2_dfrbp_1 \b.gen_square[43].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net250),
    .D(_00492_),
    .Q_N(\b.gen_square[43].sq.piece[1] ),
    .Q(_00193_));
 sg13g2_dfrbp_1 \b.gen_square[43].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net250),
    .D(_00493_),
    .Q_N(\b.gen_square[43].sq.piece[2] ),
    .Q(_00194_));
 sg13g2_dfrbp_1 \b.gen_square[44].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net252),
    .D(_00494_),
    .Q_N(_00029_),
    .Q(\b.gen_square[44].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[44].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net258),
    .D(_00313_),
    .Q_N(\b.gen_square[44].sq.mask ),
    .Q(_12104_));
 sg13g2_dfrbp_1 \b.gen_square[44].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net252),
    .D(_00495_),
    .Q_N(\b.gen_square[44].sq.piece[0] ),
    .Q(_00195_));
 sg13g2_dfrbp_1 \b.gen_square[44].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net252),
    .D(_00496_),
    .Q_N(\b.gen_square[44].sq.piece[1] ),
    .Q(_00196_));
 sg13g2_dfrbp_1 \b.gen_square[44].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net236),
    .D(_00497_),
    .Q_N(\b.gen_square[44].sq.piece[2] ),
    .Q(_00197_));
 sg13g2_dfrbp_1 \b.gen_square[45].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net258),
    .D(_00498_),
    .Q_N(_00072_),
    .Q(\b.gen_square[45].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[45].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net261),
    .D(_00314_),
    .Q_N(\b.gen_square[45].sq.mask ),
    .Q(_12105_));
 sg13g2_dfrbp_1 \b.gen_square[45].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net261),
    .D(_00499_),
    .Q_N(\b.gen_square[45].sq.piece[0] ),
    .Q(_00198_));
 sg13g2_dfrbp_1 \b.gen_square[45].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net257),
    .D(_00500_),
    .Q_N(\b.gen_square[45].sq.piece[1] ),
    .Q(_00199_));
 sg13g2_dfrbp_1 \b.gen_square[45].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net257),
    .D(_00501_),
    .Q_N(\b.gen_square[45].sq.piece[2] ),
    .Q(_00200_));
 sg13g2_dfrbp_1 \b.gen_square[46].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net258),
    .D(_00502_),
    .Q_N(_00070_),
    .Q(\b.gen_square[46].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[46].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net257),
    .D(_00315_),
    .Q_N(\b.gen_square[46].sq.mask ),
    .Q(_12106_));
 sg13g2_dfrbp_1 \b.gen_square[46].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net257),
    .D(_00503_),
    .Q_N(\b.gen_square[46].sq.piece[0] ),
    .Q(_00201_));
 sg13g2_dfrbp_1 \b.gen_square[46].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net257),
    .D(_00504_),
    .Q_N(\b.gen_square[46].sq.piece[1] ),
    .Q(_00202_));
 sg13g2_dfrbp_1 \b.gen_square[46].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net256),
    .D(_00505_),
    .Q_N(\b.gen_square[46].sq.piece[2] ),
    .Q(_00203_));
 sg13g2_dfrbp_1 \b.gen_square[47].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net256),
    .D(_00506_),
    .Q_N(_00015_),
    .Q(\b.gen_square[47].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[47].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net256),
    .D(_00316_),
    .Q_N(\b.gen_square[47].sq.mask ),
    .Q(_12107_));
 sg13g2_dfrbp_1 \b.gen_square[47].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net256),
    .D(_00507_),
    .Q_N(\b.gen_square[47].sq.piece[0] ),
    .Q(_00204_));
 sg13g2_dfrbp_1 \b.gen_square[47].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net256),
    .D(_00508_),
    .Q_N(\b.gen_square[47].sq.piece[1] ),
    .Q(_00205_));
 sg13g2_dfrbp_1 \b.gen_square[47].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net256),
    .D(_00509_),
    .Q_N(\b.gen_square[47].sq.piece[2] ),
    .Q(_00206_));
 sg13g2_dfrbp_1 \b.gen_square[48].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net236),
    .D(_00510_),
    .Q_N(_00061_),
    .Q(\b.gen_square[48].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[48].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net236),
    .D(_00317_),
    .Q_N(\b.gen_square[48].sq.mask ),
    .Q(_12108_));
 sg13g2_dfrbp_1 \b.gen_square[48].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net232),
    .D(_00511_),
    .Q_N(\b.gen_square[48].sq.piece[0] ),
    .Q(_00207_));
 sg13g2_dfrbp_1 \b.gen_square[48].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net232),
    .D(_00512_),
    .Q_N(\b.gen_square[48].sq.piece[1] ),
    .Q(_00208_));
 sg13g2_dfrbp_1 \b.gen_square[48].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net232),
    .D(_00513_),
    .Q_N(\b.gen_square[48].sq.piece[2] ),
    .Q(_00209_));
 sg13g2_dfrbp_1 \b.gen_square[49].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net232),
    .D(_00514_),
    .Q_N(_00056_),
    .Q(\b.gen_square[49].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[49].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net232),
    .D(_00318_),
    .Q_N(\b.gen_square[49].sq.mask ),
    .Q(_12109_));
 sg13g2_dfrbp_1 \b.gen_square[49].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net230),
    .D(_00515_),
    .Q_N(\b.gen_square[49].sq.piece[0] ),
    .Q(_00210_));
 sg13g2_dfrbp_1 \b.gen_square[49].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net230),
    .D(_00516_),
    .Q_N(\b.gen_square[49].sq.piece[1] ),
    .Q(_00211_));
 sg13g2_dfrbp_1 \b.gen_square[49].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net230),
    .D(_00517_),
    .Q_N(\b.gen_square[49].sq.piece[2] ),
    .Q(_00212_));
 sg13g2_dfrbp_1 \b.gen_square[4].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net285),
    .D(_00518_),
    .Q_N(_00055_),
    .Q(\b.gen_square[4].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[4].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net288),
    .D(_00319_),
    .Q_N(\b.gen_square[4].sq.mask ),
    .Q(_12110_));
 sg13g2_dfrbp_1 \b.gen_square[4].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net272),
    .D(_00519_),
    .Q_N(\b.gen_square[4].sq.piece[0] ),
    .Q(_00213_));
 sg13g2_dfrbp_1 \b.gen_square[4].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net273),
    .D(_00520_),
    .Q_N(\b.gen_square[4].sq.piece[1] ),
    .Q(_00214_));
 sg13g2_dfrbp_1 \b.gen_square[4].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net275),
    .D(_00521_),
    .Q_N(\b.gen_square[4].sq.piece[2] ),
    .Q(_00215_));
 sg13g2_dfrbp_1 \b.gen_square[50].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net255),
    .D(_00522_),
    .Q_N(_00049_),
    .Q(\b.gen_square[50].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[50].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net250),
    .D(_00320_),
    .Q_N(\b.gen_square[50].sq.mask ),
    .Q(_12111_));
 sg13g2_dfrbp_1 \b.gen_square[50].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net230),
    .D(_00523_),
    .Q_N(\b.gen_square[50].sq.piece[0] ),
    .Q(_00216_));
 sg13g2_dfrbp_1 \b.gen_square[50].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net236),
    .D(_00524_),
    .Q_N(\b.gen_square[50].sq.piece[1] ),
    .Q(_00217_));
 sg13g2_dfrbp_1 \b.gen_square[50].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net231),
    .D(_00525_),
    .Q_N(\b.gen_square[50].sq.piece[2] ),
    .Q(_00218_));
 sg13g2_dfrbp_1 \b.gen_square[51].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net249),
    .D(_00526_),
    .Q_N(_00040_),
    .Q(\b.gen_square[51].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[51].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net234),
    .D(_00321_),
    .Q_N(\b.gen_square[51].sq.mask ),
    .Q(_12112_));
 sg13g2_dfrbp_1 \b.gen_square[51].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net233),
    .D(_00527_),
    .Q_N(\b.gen_square[51].sq.piece[0] ),
    .Q(_00219_));
 sg13g2_dfrbp_1 \b.gen_square[51].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net233),
    .D(_00528_),
    .Q_N(\b.gen_square[51].sq.piece[1] ),
    .Q(_00220_));
 sg13g2_dfrbp_1 \b.gen_square[51].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net233),
    .D(_00529_),
    .Q_N(\b.gen_square[51].sq.piece[2] ),
    .Q(_00221_));
 sg13g2_dfrbp_1 \b.gen_square[52].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net249),
    .D(_00530_),
    .Q_N(_00028_),
    .Q(\b.gen_square[52].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[52].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net248),
    .D(_00322_),
    .Q_N(\b.gen_square[52].sq.mask ),
    .Q(_12113_));
 sg13g2_dfrbp_1 \b.gen_square[52].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net234),
    .D(_00531_),
    .Q_N(\b.gen_square[52].sq.piece[0] ),
    .Q(_00222_));
 sg13g2_dfrbp_1 \b.gen_square[52].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net234),
    .D(_00532_),
    .Q_N(\b.gen_square[52].sq.piece[1] ),
    .Q(_00223_));
 sg13g2_dfrbp_1 \b.gen_square[52].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net234),
    .D(_00533_),
    .Q_N(\b.gen_square[52].sq.piece[2] ),
    .Q(_00224_));
 sg13g2_dfrbp_1 \b.gen_square[53].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net258),
    .D(_00534_),
    .Q_N(_00071_),
    .Q(\b.gen_square[53].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[53].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net241),
    .D(_00323_),
    .Q_N(\b.gen_square[53].sq.mask ),
    .Q(_12114_));
 sg13g2_dfrbp_1 \b.gen_square[53].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net237),
    .D(_00535_),
    .Q_N(\b.gen_square[53].sq.piece[0] ),
    .Q(_00225_));
 sg13g2_dfrbp_1 \b.gen_square[53].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net237),
    .D(_00536_),
    .Q_N(\b.gen_square[53].sq.piece[1] ),
    .Q(_00226_));
 sg13g2_dfrbp_1 \b.gen_square[53].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net237),
    .D(_00537_),
    .Q_N(\b.gen_square[53].sq.piece[2] ),
    .Q(_00227_));
 sg13g2_dfrbp_1 \b.gen_square[54].sq.color$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net248),
    .D(_00538_),
    .Q_N(_00034_),
    .Q(\b.gen_square[54].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[54].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net248),
    .D(_00324_),
    .Q_N(\b.gen_square[54].sq.mask ),
    .Q(_12115_));
 sg13g2_dfrbp_1 \b.gen_square[54].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net246),
    .D(_00539_),
    .Q_N(\b.gen_square[54].sq.piece[0] ),
    .Q(_00228_));
 sg13g2_dfrbp_1 \b.gen_square[54].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net246),
    .D(_00540_),
    .Q_N(\b.gen_square[54].sq.piece[1] ),
    .Q(_00229_));
 sg13g2_dfrbp_1 \b.gen_square[54].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net246),
    .D(_00541_),
    .Q_N(\b.gen_square[54].sq.piece[2] ),
    .Q(_00230_));
 sg13g2_dfrbp_1 \b.gen_square[55].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net256),
    .D(_00542_),
    .Q_N(_00039_),
    .Q(\b.gen_square[55].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[55].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net246),
    .D(_00325_),
    .Q_N(\b.gen_square[55].sq.mask ),
    .Q(_12116_));
 sg13g2_dfrbp_1 \b.gen_square[55].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net246),
    .D(_00543_),
    .Q_N(\b.gen_square[55].sq.piece[0] ),
    .Q(_00231_));
 sg13g2_dfrbp_1 \b.gen_square[55].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net246),
    .D(_00544_),
    .Q_N(\b.gen_square[55].sq.piece[1] ),
    .Q(_00232_));
 sg13g2_dfrbp_1 \b.gen_square[55].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net247),
    .D(_00545_),
    .Q_N(\b.gen_square[55].sq.piece[2] ),
    .Q(_00233_));
 sg13g2_dfrbp_1 \b.gen_square[56].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net231),
    .D(_00546_),
    .Q_N(_00027_),
    .Q(\b.gen_square[56].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[56].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net230),
    .D(_00326_),
    .Q_N(\b.gen_square[56].sq.mask ),
    .Q(_12117_));
 sg13g2_dfrbp_1 \b.gen_square[56].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net230),
    .D(_00547_),
    .Q_N(\b.gen_square[56].sq.piece[0] ),
    .Q(_00234_));
 sg13g2_dfrbp_1 \b.gen_square[56].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net230),
    .D(_00548_),
    .Q_N(\b.gen_square[56].sq.piece[1] ),
    .Q(_00235_));
 sg13g2_dfrbp_1 \b.gen_square[56].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net230),
    .D(_00549_),
    .Q_N(\b.gen_square[56].sq.piece[2] ),
    .Q(_00236_));
 sg13g2_dfrbp_1 \b.gen_square[57].sq.color$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net232),
    .D(_00550_),
    .Q_N(_00026_),
    .Q(\b.gen_square[57].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[57].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net231),
    .D(_00327_),
    .Q_N(\b.gen_square[57].sq.mask ),
    .Q(_12118_));
 sg13g2_dfrbp_1 \b.gen_square[57].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net231),
    .D(_00551_),
    .Q_N(\b.gen_square[57].sq.piece[0] ),
    .Q(_00237_));
 sg13g2_dfrbp_1 \b.gen_square[57].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net231),
    .D(_00552_),
    .Q_N(\b.gen_square[57].sq.piece[1] ),
    .Q(_00238_));
 sg13g2_dfrbp_1 \b.gen_square[57].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net231),
    .D(_00553_),
    .Q_N(\b.gen_square[57].sq.piece[2] ),
    .Q(_00239_));
 sg13g2_dfrbp_1 \b.gen_square[58].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net235),
    .D(_00554_),
    .Q_N(_00025_),
    .Q(\b.gen_square[58].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[58].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net233),
    .D(_00328_),
    .Q_N(\b.gen_square[58].sq.mask ),
    .Q(_12119_));
 sg13g2_dfrbp_1 \b.gen_square[58].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net233),
    .D(_00555_),
    .Q_N(\b.gen_square[58].sq.piece[0] ),
    .Q(_00240_));
 sg13g2_dfrbp_1 \b.gen_square[58].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net233),
    .D(_00556_),
    .Q_N(\b.gen_square[58].sq.piece[1] ),
    .Q(_00241_));
 sg13g2_dfrbp_1 \b.gen_square[58].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net232),
    .D(_00557_),
    .Q_N(\b.gen_square[58].sq.piece[2] ),
    .Q(_00242_));
 sg13g2_dfrbp_1 \b.gen_square[59].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net234),
    .D(_00558_),
    .Q_N(_00024_),
    .Q(\b.gen_square[59].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[59].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net234),
    .D(_00329_),
    .Q_N(\b.gen_square[59].sq.mask ),
    .Q(_12120_));
 sg13g2_dfrbp_1 \b.gen_square[59].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net234),
    .D(_00559_),
    .Q_N(\b.gen_square[59].sq.piece[0] ),
    .Q(_00243_));
 sg13g2_dfrbp_1 \b.gen_square[59].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net233),
    .D(_00560_),
    .Q_N(\b.gen_square[59].sq.piece[1] ),
    .Q(_00244_));
 sg13g2_dfrbp_1 \b.gen_square[59].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net233),
    .D(_00561_),
    .Q_N(\b.gen_square[59].sq.piece[2] ),
    .Q(_00245_));
 sg13g2_dfrbp_1 \b.gen_square[5].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net285),
    .D(_00562_),
    .Q_N(_00048_),
    .Q(\b.gen_square[5].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[5].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net288),
    .D(_00330_),
    .Q_N(\b.gen_square[5].sq.mask ),
    .Q(_12121_));
 sg13g2_dfrbp_1 \b.gen_square[5].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net259),
    .D(_00563_),
    .Q_N(\b.gen_square[5].sq.piece[0] ),
    .Q(_00246_));
 sg13g2_dfrbp_1 \b.gen_square[5].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net259),
    .D(_00564_),
    .Q_N(\b.gen_square[5].sq.piece[1] ),
    .Q(_00247_));
 sg13g2_dfrbp_1 \b.gen_square[5].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net260),
    .D(_00565_),
    .Q_N(\b.gen_square[5].sq.piece[2] ),
    .Q(_00248_));
 sg13g2_dfrbp_1 \b.gen_square[60].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net235),
    .D(_00566_),
    .Q_N(_00023_),
    .Q(\b.gen_square[60].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[60].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net237),
    .D(_00331_),
    .Q_N(\b.gen_square[60].sq.mask ),
    .Q(_12122_));
 sg13g2_dfrbp_1 \b.gen_square[60].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net235),
    .D(_00567_),
    .Q_N(\b.gen_square[60].sq.piece[0] ),
    .Q(_00249_));
 sg13g2_dfrbp_1 \b.gen_square[60].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net235),
    .D(_00568_),
    .Q_N(\b.gen_square[60].sq.piece[1] ),
    .Q(_00250_));
 sg13g2_dfrbp_1 \b.gen_square[60].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net235),
    .D(_00569_),
    .Q_N(\b.gen_square[60].sq.piece[2] ),
    .Q(_00251_));
 sg13g2_dfrbp_1 \b.gen_square[61].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net248),
    .D(_00570_),
    .Q_N(_00022_),
    .Q(\b.gen_square[61].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[61].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net237),
    .D(_00332_),
    .Q_N(\b.gen_square[61].sq.mask ),
    .Q(_12123_));
 sg13g2_dfrbp_1 \b.gen_square[61].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net237),
    .D(_00571_),
    .Q_N(\b.gen_square[61].sq.piece[0] ),
    .Q(_00252_));
 sg13g2_dfrbp_1 \b.gen_square[61].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net238),
    .D(_00572_),
    .Q_N(\b.gen_square[61].sq.piece[1] ),
    .Q(_00253_));
 sg13g2_dfrbp_1 \b.gen_square[61].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net237),
    .D(_00573_),
    .Q_N(\b.gen_square[61].sq.piece[2] ),
    .Q(_00254_));
 sg13g2_dfrbp_1 \b.gen_square[62].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net247),
    .D(_00574_),
    .Q_N(_00021_),
    .Q(\b.gen_square[62].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[62].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net246),
    .D(_00333_),
    .Q_N(\b.gen_square[62].sq.mask ),
    .Q(_12124_));
 sg13g2_dfrbp_1 \b.gen_square[62].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net247),
    .D(_00575_),
    .Q_N(\b.gen_square[62].sq.piece[0] ),
    .Q(_00255_));
 sg13g2_dfrbp_1 \b.gen_square[62].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net247),
    .D(_00576_),
    .Q_N(\b.gen_square[62].sq.piece[1] ),
    .Q(_00256_));
 sg13g2_dfrbp_1 \b.gen_square[62].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net247),
    .D(_00577_),
    .Q_N(\b.gen_square[62].sq.piece[2] ),
    .Q(_00257_));
 sg13g2_dfrbp_1 \b.gen_square[63].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net248),
    .D(_00578_),
    .Q_N(_00033_),
    .Q(\b.gen_square[63].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[63].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net246),
    .D(_00334_),
    .Q_N(\b.gen_square[63].sq.mask ),
    .Q(_12125_));
 sg13g2_dfrbp_1 \b.gen_square[63].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net241),
    .D(_00579_),
    .Q_N(\b.gen_square[63].sq.piece[0] ),
    .Q(_00258_));
 sg13g2_dfrbp_1 \b.gen_square[63].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net241),
    .D(_00580_),
    .Q_N(\b.gen_square[63].sq.piece[1] ),
    .Q(_00259_));
 sg13g2_dfrbp_1 \b.gen_square[63].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net244),
    .D(_00581_),
    .Q_N(\b.gen_square[63].sq.piece[2] ),
    .Q(_00260_));
 sg13g2_dfrbp_1 \b.gen_square[6].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net285),
    .D(_00582_),
    .Q_N(_00077_),
    .Q(\b.gen_square[6].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[6].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net289),
    .D(_00335_),
    .Q_N(\b.gen_square[6].sq.mask ),
    .Q(_12126_));
 sg13g2_dfrbp_1 \b.gen_square[6].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net286),
    .D(_00583_),
    .Q_N(\b.gen_square[6].sq.piece[0] ),
    .Q(_00261_));
 sg13g2_dfrbp_1 \b.gen_square[6].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net286),
    .D(_00584_),
    .Q_N(\b.gen_square[6].sq.piece[1] ),
    .Q(_00262_));
 sg13g2_dfrbp_1 \b.gen_square[6].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net289),
    .D(_00585_),
    .Q_N(\b.gen_square[6].sq.piece[2] ),
    .Q(_00263_));
 sg13g2_dfrbp_1 \b.gen_square[7].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net277),
    .D(_00586_),
    .Q_N(_00020_),
    .Q(\b.gen_square[7].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[7].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net276),
    .D(_00336_),
    .Q_N(\b.gen_square[7].sq.mask ),
    .Q(_12127_));
 sg13g2_dfrbp_1 \b.gen_square[7].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net276),
    .D(_00587_),
    .Q_N(\b.gen_square[7].sq.piece[0] ),
    .Q(_00264_));
 sg13g2_dfrbp_1 \b.gen_square[7].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net276),
    .D(_00588_),
    .Q_N(\b.gen_square[7].sq.piece[1] ),
    .Q(_00265_));
 sg13g2_dfrbp_1 \b.gen_square[7].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net277),
    .D(_00589_),
    .Q_N(\b.gen_square[7].sq.piece[2] ),
    .Q(_00266_));
 sg13g2_dfrbp_1 \b.gen_square[8].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net279),
    .D(_00590_),
    .Q_N(_00066_),
    .Q(\b.gen_square[8].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[8].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net280),
    .D(_00337_),
    .Q_N(\b.gen_square[8].sq.mask ),
    .Q(_12128_));
 sg13g2_dfrbp_1 \b.gen_square[8].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net281),
    .D(_00591_),
    .Q_N(\b.gen_square[8].sq.piece[0] ),
    .Q(_00267_));
 sg13g2_dfrbp_1 \b.gen_square[8].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net281),
    .D(_00592_),
    .Q_N(\b.gen_square[8].sq.piece[1] ),
    .Q(_00268_));
 sg13g2_dfrbp_1 \b.gen_square[8].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net281),
    .D(_00593_),
    .Q_N(\b.gen_square[8].sq.piece[2] ),
    .Q(_00269_));
 sg13g2_dfrbp_1 \b.gen_square[9].sq.color$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net280),
    .D(_00594_),
    .Q_N(_00076_),
    .Q(\b.gen_square[9].sq.color ));
 sg13g2_dfrbp_1 \b.gen_square[9].sq.mask$_DFF_PN1_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net269),
    .D(_00338_),
    .Q_N(\b.gen_square[9].sq.mask ),
    .Q(_12129_));
 sg13g2_dfrbp_1 \b.gen_square[9].sq.piece[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net282),
    .D(_00595_),
    .Q_N(\b.gen_square[9].sq.piece[0] ),
    .Q(_00270_));
 sg13g2_dfrbp_1 \b.gen_square[9].sq.piece[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net282),
    .D(_00596_),
    .Q_N(\b.gen_square[9].sq.piece[1] ),
    .Q(_00271_));
 sg13g2_dfrbp_1 \b.gen_square[9].sq.piece[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net281),
    .D(_00597_),
    .Q_N(\b.gen_square[9].sq.piece[2] ),
    .Q(_00272_));
 sg13g2_dfrbp_1 \data_out[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net244),
    .D(_00598_),
    .Q_N(_12053_),
    .Q(\data_out[0] ));
 sg13g2_dfrbp_1 \data_out[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net244),
    .D(_00599_),
    .Q_N(_12052_),
    .Q(\data_out[1] ));
 sg13g2_dfrbp_1 \data_out[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net244),
    .D(_00600_),
    .Q_N(_12051_),
    .Q(\data_out[2] ));
 sg13g2_dfrbp_1 \data_out[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net245),
    .D(_00601_),
    .Q_N(_12050_),
    .Q(\data_out[3] ));
 sg13g2_dfrbp_1 \data_out_valid$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net243),
    .D(_00602_),
    .Q_N(_12057_),
    .Q(data_out_valid));
 sg13g2_dfrbp_1 \mask_mode[1]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net241),
    .D(_00001_),
    .Q_N(_00068_),
    .Q(\mask_mode[1] ));
 sg13g2_dfrbp_1 \mask_mode[2]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net239),
    .D(_00002_),
    .Q_N(_12058_),
    .Q(\mask_mode[2] ));
 sg13g2_dfrbp_1 \mask_mode[3]$_DFF_PN0_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net244),
    .D(_00003_),
    .Q_N(_12049_),
    .Q(\mask_mode[3] ));
 sg13g2_dfrbp_1 \spi.bit_count$_DFFE_PN1P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net243),
    .D(_00603_),
    .Q_N(\spi.bit_count ),
    .Q(_00273_));
 sg13g2_dfrbp_1 \spi.din[0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net313),
    .D(_00604_),
    .Q_N(_12048_),
    .Q(\data_in[0] ));
 sg13g2_dfrbp_1 \spi.din[1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net314),
    .D(_00605_),
    .Q_N(_12047_),
    .Q(\data_in[1] ));
 sg13g2_dfrbp_1 \spi.din[2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net315),
    .D(_00606_),
    .Q_N(_12046_),
    .Q(\data_in[2] ));
 sg13g2_dfrbp_1 \spi.din[3]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net316),
    .D(_00607_),
    .Q_N(_12059_),
    .Q(\data_in[3] ));
 sg13g2_dfrbp_1 \spi.din_valid$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net243),
    .D(_00011_),
    .Q_N(_00067_),
    .Q(data_in_valid));
 sg13g2_dfrbp_1 \spi.sck_r0$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net243),
    .D(net3),
    .Q_N(_12045_),
    .Q(\spi.sck_r0 ));
 sg13g2_dfrbp_1 \spi.sdi_r[0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net317),
    .D(_00608_),
    .Q_N(_12044_),
    .Q(\spi.sdi_r[0] ));
 sg13g2_dfrbp_1 \spi.sdi_r[1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net318),
    .D(_00609_),
    .Q_N(_12043_),
    .Q(\spi.sdi_r[1] ));
 sg13g2_dfrbp_1 \spi.sdi_r[2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net319),
    .D(_00610_),
    .Q_N(_12042_),
    .Q(\spi.sdi_r[2] ));
 sg13g2_dfrbp_1 \spi.sdi_r[3]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net320),
    .D(_00611_),
    .Q_N(_12041_),
    .Q(\spi.sdi_r[3] ));
 sg13g2_dfrbp_1 \ss1[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net244),
    .D(_00612_),
    .Q_N(_12040_),
    .Q(\b.ss1[0] ));
 sg13g2_dfrbp_1 \ss1[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net242),
    .D(_00613_),
    .Q_N(_12039_),
    .Q(\b.ss1[1] ));
 sg13g2_dfrbp_1 \ss1[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net244),
    .D(_00614_),
    .Q_N(_12038_),
    .Q(\b.ss1[2] ));
 sg13g2_dfrbp_1 \ss1[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net240),
    .D(_00615_),
    .Q_N(_12037_),
    .Q(\b.ss1[3] ));
 sg13g2_dfrbp_1 \ss1[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net240),
    .D(_00616_),
    .Q_N(_12036_),
    .Q(\b.ss1[4] ));
 sg13g2_dfrbp_1 \ss1[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net240),
    .D(_00617_),
    .Q_N(_12035_),
    .Q(\b.ss1[5] ));
 sg13g2_dfrbp_1 \ss2[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net238),
    .D(_00618_),
    .Q_N(_12034_),
    .Q(\ss2[0] ));
 sg13g2_dfrbp_1 \ss2[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net239),
    .D(_00619_),
    .Q_N(_12033_),
    .Q(\ss2[1] ));
 sg13g2_dfrbp_1 \ss2[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net240),
    .D(_00620_),
    .Q_N(_12032_),
    .Q(\ss2[2] ));
 sg13g2_dfrbp_1 \ss2[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net239),
    .D(_00621_),
    .Q_N(_12031_),
    .Q(\ss2[3] ));
 sg13g2_dfrbp_1 \ss2[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net239),
    .D(_00622_),
    .Q_N(_12030_),
    .Q(\ss2[4] ));
 sg13g2_dfrbp_1 \ss2[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net239),
    .D(_00623_),
    .Q_N(_12029_),
    .Q(\ss2[5] ));
 sg13g2_dfrbp_1 \state[0]$_DFF_PN1_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net245),
    .D(_00339_),
    .Q_N(\state[0] ),
    .Q(_12130_));
 sg13g2_dfrbp_1 \state[10]$_DFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net242),
    .D(_00004_),
    .Q_N(_12060_),
    .Q(\state[10] ));
 sg13g2_dfrbp_1 \state[1]$_DFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net242),
    .D(_00005_),
    .Q_N(_12061_),
    .Q(\state[1] ));
 sg13g2_dfrbp_1 \state[3]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net239),
    .D(_00006_),
    .Q_N(_12062_),
    .Q(\state[3] ));
 sg13g2_dfrbp_1 \state[4]$_DFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net242),
    .D(_00007_),
    .Q_N(_12063_),
    .Q(\state[4] ));
 sg13g2_dfrbp_1 \state[5]$_DFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net242),
    .D(_00008_),
    .Q_N(_00069_),
    .Q(\state[5] ));
 sg13g2_dfrbp_1 \state[6]$_DFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net242),
    .D(_00009_),
    .Q_N(_12064_),
    .Q(\state[6] ));
 sg13g2_dfrbp_1 \state[7]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net239),
    .D(net121),
    .Q_N(_12065_),
    .Q(\state[7] ));
 sg13g2_dfrbp_1 \state[9]$_DFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net242),
    .D(_00010_),
    .Q_N(_12028_),
    .Q(\state[9] ));
 sg13g2_dfrbp_1 \state_mode[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net237),
    .D(_00624_),
    .Q_N(_12027_),
    .Q(\b.gen_square[0].sq.state_mode[0] ));
 sg13g2_dfrbp_1 \state_mode[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net238),
    .D(_00625_),
    .Q_N(_12026_),
    .Q(\b.gen_square[0].sq.state_mode[1] ));
 sg13g2_dfrbp_1 \state_mode[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net243),
    .D(_00626_),
    .Q_N(\b.gen_square[0].sq.state_mode[2] ),
    .Q(_00274_));
 sg13g2_dfrbp_1 \write_bus[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net245),
    .D(_00627_),
    .Q_N(_00080_),
    .Q(\b.gen_square[0].sq.write_bus[0] ));
 sg13g2_dfrbp_1 \write_bus[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net243),
    .D(_00628_),
    .Q_N(_00079_),
    .Q(\b.gen_square[0].sq.write_bus[1] ));
 sg13g2_dfrbp_1 \write_bus[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net245),
    .D(_00629_),
    .Q_N(_00078_),
    .Q(\b.gen_square[0].sq.write_bus[2] ));
 sg13g2_dfrbp_1 \write_bus[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net244),
    .D(_00630_),
    .Q_N(_12025_),
    .Q(\b.gen_square[0].sq.write_bus[3] ));
 sg13g2_dfrbp_1 \wtm$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net231),
    .D(_00631_),
    .Q_N(_12024_),
    .Q(\b.gen_square[0].sq.wtm ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[4]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[5]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[6]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout12 (.A(_01978_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_01944_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_07962_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_03851_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_03752_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_03660_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_03602_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_03538_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_02155_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_06199_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_05953_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_04699_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_02144_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_07100_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_06580_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_06186_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_05961_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_04959_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_04698_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_04675_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_04370_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_04154_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_04117_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_06579_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_06530_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_06334_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_05710_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_05408_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_05347_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_05092_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_04898_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_04835_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_04674_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_04651_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_04348_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_04217_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_02122_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_06955_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_06697_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_06392_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_05691_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_05647_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_05378_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_05346_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_05116_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_05091_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_04928_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_04834_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_04550_),
    .X(net60));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(_04347_));
 sg13g2_buf_2 fanout62 (.A(_04216_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_02111_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_07071_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_06954_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_06735_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_05115_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_05090_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_04530_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_04300_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_04129_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_02100_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_05890_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_05678_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_05114_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_05089_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_04724_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_04511_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_04313_),
    .X(net79));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_04287_));
 sg13g2_buf_2 fanout81 (.A(_04253_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_04248_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_02089_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_05727_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_05113_),
    .X(net85));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(_05088_));
 sg13g2_buf_2 fanout87 (.A(_04626_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_04510_),
    .X(net88));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(_04286_));
 sg13g2_buf_2 fanout90 (.A(_04194_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_04090_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_04086_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_02078_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_05167_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_05112_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_05087_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_05079_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_05046_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_04509_),
    .X(net99));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(_04285_));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(_04089_));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(_04085_));
 sg13g2_buf_2 fanout103 (.A(_02067_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_03318_),
    .X(net104));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(_03215_));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_03169_));
 sg13g2_buf_2 fanout107 (.A(_03159_),
    .X(net107));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(_03117_));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(_03096_));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_03083_));
 sg13g2_buf_2 fanout111 (.A(_03075_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_05111_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_05086_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_05078_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_04508_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_04211_),
    .X(net116));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(_04088_));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(_04084_));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(_04051_));
 sg13g2_buf_2 fanout120 (.A(_02056_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_00000_),
    .X(net121));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(_03302_));
 sg13g2_buf_2 fanout123 (.A(_03082_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_03074_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_03065_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_06573_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_06381_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_05110_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_05085_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_05077_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_04843_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_04825_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_04485_),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(_04087_));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(_04083_));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(_04079_));
 sg13g2_buf_2 fanout137 (.A(_02045_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_03180_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_03104_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_03086_),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(_03064_));
 sg13g2_buf_2 fanout142 (.A(_07412_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_05109_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_05084_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_05076_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_04918_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_04263_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_04243_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_04141_),
    .X(net149));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(_04078_));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(_04065_));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_04061_));
 sg13g2_buf_2 fanout153 (.A(_03521_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_02034_),
    .X(net154));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(_03163_));
 sg13g2_buf_2 fanout156 (.A(_03085_),
    .X(net156));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(_03078_));
 sg13g2_buf_2 fanout158 (.A(_07381_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_06158_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_05108_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_05083_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_05075_),
    .X(net162));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(_04642_));
 sg13g2_buf_2 fanout164 (.A(_04532_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_04241_),
    .X(net165));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(_04077_));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(_04064_));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(_04048_));
 sg13g2_buf_2 fanout169 (.A(_03902_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_03697_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_01836_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_03280_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_03183_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_03091_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_03071_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_05082_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_05074_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_04717_),
    .X(net178));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(_04076_));
 sg13g2_buf_2 fanout180 (.A(_04038_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_03876_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_03390_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_02012_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_00882_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_03275_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_03178_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_03166_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_03089_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_02798_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_05555_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_05073_),
    .X(net191));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(_04046_));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(_04039_));
 sg13g2_buf_2 fanout194 (.A(_03837_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_03835_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_03833_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_03738_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_03736_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_03734_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_03648_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_03646_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_03644_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_03546_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_03544_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_03542_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_02361_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_02307_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_02253_),
    .X(net208));
 sg13g2_buf_4 fanout209 (.X(net209),
    .A(_01664_));
 sg13g2_buf_2 fanout210 (.A(_03271_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_03177_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_03173_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_03165_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_03092_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_05072_),
    .X(net215));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(_04036_));
 sg13g2_buf_2 fanout217 (.A(_03954_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_03925_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_03923_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_03921_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_03854_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_03755_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_03663_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_03562_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_02350_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_02296_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_02242_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_02199_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_01231_),
    .X(net229));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(net231));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(net232));
 sg13g2_buf_4 fanout232 (.X(net232),
    .A(net236));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(net234));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(net235));
 sg13g2_buf_2 fanout235 (.A(net236),
    .X(net235));
 sg13g2_buf_4 fanout236 (.X(net236),
    .A(net249));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(net238));
 sg13g2_buf_2 fanout238 (.A(net241),
    .X(net238));
 sg13g2_buf_4 fanout239 (.X(net239),
    .A(net241));
 sg13g2_buf_2 fanout240 (.A(net241),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(net249),
    .X(net241));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(net243));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(net245));
 sg13g2_buf_4 fanout244 (.X(net244),
    .A(net245));
 sg13g2_buf_2 fanout245 (.A(net249),
    .X(net245));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(net248));
 sg13g2_buf_2 fanout247 (.A(net248),
    .X(net247));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(net249));
 sg13g2_buf_2 fanout249 (.A(net262),
    .X(net249));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(net252));
 sg13g2_buf_2 fanout251 (.A(net252),
    .X(net251));
 sg13g2_buf_4 fanout252 (.X(net252),
    .A(net255));
 sg13g2_buf_4 fanout253 (.X(net253),
    .A(net254));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(net255));
 sg13g2_buf_2 fanout255 (.A(net262),
    .X(net255));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(net258));
 sg13g2_buf_2 fanout257 (.A(net258),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(net262),
    .X(net258));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(net260));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(net261));
 sg13g2_buf_2 fanout261 (.A(net262),
    .X(net261));
 sg13g2_buf_1 fanout262 (.A(net1),
    .X(net262));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(net270));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(net270));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(net266));
 sg13g2_buf_2 fanout266 (.A(net270),
    .X(net266));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(net269));
 sg13g2_buf_2 fanout268 (.A(net269),
    .X(net268));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(net270));
 sg13g2_buf_1 fanout270 (.A(net292),
    .X(net270));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(net273));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(net273));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(net292),
    .X(net274));
 sg13g2_buf_4 fanout275 (.X(net275),
    .A(net276));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(net277));
 sg13g2_buf_2 fanout277 (.A(net292),
    .X(net277));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(net284));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(net280));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(net284));
 sg13g2_buf_4 fanout281 (.X(net281),
    .A(net282));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(net283));
 sg13g2_buf_2 fanout283 (.A(net284),
    .X(net283));
 sg13g2_buf_1 fanout284 (.A(net292),
    .X(net284));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(net291));
 sg13g2_buf_2 fanout286 (.A(net291),
    .X(net286));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(net288));
 sg13g2_buf_2 fanout288 (.A(net291),
    .X(net288));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(net291));
 sg13g2_buf_2 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_1 fanout291 (.A(net292),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(net1),
    .X(net292));
 sg13g2_tielo _23902__293 (.L_LO(net293));
 sg13g2_tielo _23903__294 (.L_LO(net294));
 sg13g2_tielo _23904__295 (.L_LO(net295));
 sg13g2_tielo _23905__296 (.L_LO(net296));
 sg13g2_tielo _23906__297 (.L_LO(net297));
 sg13g2_tielo _23907__298 (.L_LO(net298));
 sg13g2_tielo _23908__299 (.L_LO(net299));
 sg13g2_tielo _23909__300 (.L_LO(net300));
 sg13g2_tielo _23910__301 (.L_LO(net301));
 sg13g2_tielo _23911__302 (.L_LO(net302));
 sg13g2_tielo _23912__303 (.L_LO(net303));
 sg13g2_tielo _23913__304 (.L_LO(net304));
 sg13g2_tielo _23914__305 (.L_LO(net305));
 sg13g2_tielo _23915__306 (.L_LO(net306));
 sg13g2_tielo _23916__307 (.L_LO(net307));
 sg13g2_tielo _23917__308 (.L_LO(net308));
 sg13g2_tielo _23918__309 (.L_LO(net309));
 sg13g2_tielo _23919__310 (.L_LO(net310));
 sg13g2_tielo _23920__311 (.L_LO(net311));
 sg13g2_tielo _23921__312 (.L_LO(net312));
 sg13g2_tiehi \spi.din[1]$_DFFE_PP__314  (.L_HI(net314));
 sg13g2_tiehi \spi.din[2]$_DFFE_PP__315  (.L_HI(net315));
 sg13g2_tiehi \spi.din[3]$_DFFE_PP__316  (.L_HI(net316));
 sg13g2_tiehi \spi.sdi_r[0]$_DFFE_PP__317  (.L_HI(net317));
 sg13g2_tiehi \spi.sdi_r[1]$_DFFE_PP__318  (.L_HI(net318));
 sg13g2_tiehi \spi.sdi_r[2]$_DFFE_PP__319  (.L_HI(net319));
 sg13g2_tiehi \spi.sdi_r[3]$_DFFE_PP__320  (.L_HI(net320));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_leaf_62_clk (.X(clknet_leaf_62_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_63_clk (.X(clknet_leaf_63_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_64_clk (.X(clknet_leaf_64_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_65_clk (.X(clknet_leaf_65_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_66_clk (.X(clknet_leaf_66_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_67_clk (.X(clknet_leaf_67_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_leaf_68_clk (.X(clknet_leaf_68_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_leaf_69_clk (.X(clknet_leaf_69_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_70_clk (.X(clknet_leaf_70_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_leaf_71_clk (.X(clknet_leaf_71_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkload7 (.A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkload9 (.A(clknet_4_13_0_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_4_15_0_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_0_clk));
 sg13g2_buf_16 clkload12 (.A(clknet_leaf_69_clk));
 sg13g2_buf_16 clkload13 (.A(clknet_leaf_2_clk));
 sg13g2_buf_16 clkload14 (.A(clknet_leaf_6_clk));
 sg13g2_buf_16 clkload15 (.A(clknet_leaf_63_clk));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_64_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_66_clk));
 sg13g2_buf_16 clkload18 (.A(clknet_leaf_68_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_7_clk));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_67_clk));
 sg13g2_buf_16 clkload21 (.A(clknet_leaf_5_clk));
 sg13g2_buf_16 clkload22 (.A(clknet_leaf_12_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_17_clk));
 sg13g2_buf_8 clkload25 (.A(clknet_leaf_58_clk));
 sg13g2_inv_4 clkload26 (.A(clknet_leaf_59_clk));
 sg13g2_inv_2 clkload27 (.A(clknet_leaf_9_clk));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_47_clk));
 sg13g2_buf_8 clkload29 (.A(clknet_leaf_61_clk));
 sg13g2_buf_16 clkload30 (.A(clknet_leaf_49_clk));
 sg13g2_buf_16 clkload31 (.A(clknet_leaf_52_clk));
 sg13g2_buf_8 clkload32 (.A(clknet_leaf_43_clk));
 sg13g2_buf_16 clkload33 (.A(clknet_leaf_44_clk));
 sg13g2_inv_1 clkload34 (.A(clknet_leaf_51_clk));
 sg13g2_inv_1 clkload35 (.A(clknet_leaf_30_clk));
 sg13g2_inv_1 clkload36 (.A(clknet_leaf_31_clk));
 sg13g2_inv_2 clkload37 (.A(clknet_leaf_33_clk));
 sg13g2_inv_2 clkload38 (.A(clknet_leaf_46_clk));
 sg13g2_buf_8 clkload39 (.A(clknet_leaf_26_clk));
 sg13g2_inv_2 clkload40 (.A(clknet_leaf_27_clk));
 sg13g2_inv_4 clkload41 (.A(clknet_leaf_41_clk));
 sg13g2_buf_8 clkload42 (.A(clknet_leaf_42_clk));
 sg13g2_buf_16 clkload43 (.A(clknet_leaf_45_clk));
 sg13g2_buf_16 clkload44 (.A(clknet_leaf_32_clk));
 sg13g2_buf_8 clkload45 (.A(clknet_leaf_37_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00631_));
 sg13g2_antennanp ANTENNA_2 (.A(_01231_));
 sg13g2_antennanp ANTENNA_3 (.A(_01231_));
 sg13g2_antennanp ANTENNA_4 (.A(_01231_));
 sg13g2_antennanp ANTENNA_5 (.A(_01231_));
 sg13g2_antennanp ANTENNA_6 (.A(_01231_));
 sg13g2_antennanp ANTENNA_7 (.A(_01231_));
 sg13g2_antennanp ANTENNA_8 (.A(_01653_));
 sg13g2_antennanp ANTENNA_9 (.A(_01653_));
 sg13g2_antennanp ANTENNA_10 (.A(_01653_));
 sg13g2_antennanp ANTENNA_11 (.A(_01653_));
 sg13g2_antennanp ANTENNA_12 (.A(_01653_));
 sg13g2_antennanp ANTENNA_13 (.A(_01653_));
 sg13g2_antennanp ANTENNA_14 (.A(_01653_));
 sg13g2_antennanp ANTENNA_15 (.A(_01653_));
 sg13g2_antennanp ANTENNA_16 (.A(_01653_));
 sg13g2_antennanp ANTENNA_17 (.A(_01653_));
 sg13g2_antennanp ANTENNA_18 (.A(_01653_));
 sg13g2_antennanp ANTENNA_19 (.A(_01653_));
 sg13g2_antennanp ANTENNA_20 (.A(_01653_));
 sg13g2_antennanp ANTENNA_21 (.A(_01653_));
 sg13g2_antennanp ANTENNA_22 (.A(_01653_));
 sg13g2_antennanp ANTENNA_23 (.A(_01653_));
 sg13g2_antennanp ANTENNA_24 (.A(_01653_));
 sg13g2_antennanp ANTENNA_25 (.A(_01653_));
 sg13g2_antennanp ANTENNA_26 (.A(_01653_));
 sg13g2_antennanp ANTENNA_27 (.A(_01653_));
 sg13g2_antennanp ANTENNA_28 (.A(_01653_));
 sg13g2_antennanp ANTENNA_29 (.A(_01653_));
 sg13g2_antennanp ANTENNA_30 (.A(_01653_));
 sg13g2_antennanp ANTENNA_31 (.A(_01653_));
 sg13g2_antennanp ANTENNA_32 (.A(_01653_));
 sg13g2_antennanp ANTENNA_33 (.A(_01653_));
 sg13g2_antennanp ANTENNA_34 (.A(_01653_));
 sg13g2_antennanp ANTENNA_35 (.A(_01653_));
 sg13g2_antennanp ANTENNA_36 (.A(_01653_));
 sg13g2_antennanp ANTENNA_37 (.A(_01653_));
 sg13g2_antennanp ANTENNA_38 (.A(_01653_));
 sg13g2_antennanp ANTENNA_39 (.A(_01653_));
 sg13g2_antennanp ANTENNA_40 (.A(_02012_));
 sg13g2_antennanp ANTENNA_41 (.A(_02012_));
 sg13g2_antennanp ANTENNA_42 (.A(_02012_));
 sg13g2_antennanp ANTENNA_43 (.A(_02012_));
 sg13g2_antennanp ANTENNA_44 (.A(_02067_));
 sg13g2_antennanp ANTENNA_45 (.A(_02067_));
 sg13g2_antennanp ANTENNA_46 (.A(_02067_));
 sg13g2_antennanp ANTENNA_47 (.A(_02078_));
 sg13g2_antennanp ANTENNA_48 (.A(_02078_));
 sg13g2_antennanp ANTENNA_49 (.A(_02078_));
 sg13g2_antennanp ANTENNA_50 (.A(_02078_));
 sg13g2_antennanp ANTENNA_51 (.A(_02078_));
 sg13g2_antennanp ANTENNA_52 (.A(_02078_));
 sg13g2_antennanp ANTENNA_53 (.A(_02078_));
 sg13g2_antennanp ANTENNA_54 (.A(_02242_));
 sg13g2_antennanp ANTENNA_55 (.A(_02242_));
 sg13g2_antennanp ANTENNA_56 (.A(_02296_));
 sg13g2_antennanp ANTENNA_57 (.A(_02296_));
 sg13g2_antennanp ANTENNA_58 (.A(_02296_));
 sg13g2_antennanp ANTENNA_59 (.A(_02296_));
 sg13g2_antennanp ANTENNA_60 (.A(_02350_));
 sg13g2_antennanp ANTENNA_61 (.A(_02350_));
 sg13g2_antennanp ANTENNA_62 (.A(_02807_));
 sg13g2_antennanp ANTENNA_63 (.A(_02899_));
 sg13g2_antennanp ANTENNA_64 (.A(_02899_));
 sg13g2_antennanp ANTENNA_65 (.A(_02902_));
 sg13g2_antennanp ANTENNA_66 (.A(_02902_));
 sg13g2_antennanp ANTENNA_67 (.A(_02906_));
 sg13g2_antennanp ANTENNA_68 (.A(_02914_));
 sg13g2_antennanp ANTENNA_69 (.A(_02919_));
 sg13g2_antennanp ANTENNA_70 (.A(_02921_));
 sg13g2_antennanp ANTENNA_71 (.A(_02947_));
 sg13g2_antennanp ANTENNA_72 (.A(_02948_));
 sg13g2_antennanp ANTENNA_73 (.A(_02953_));
 sg13g2_antennanp ANTENNA_74 (.A(_02954_));
 sg13g2_antennanp ANTENNA_75 (.A(_02957_));
 sg13g2_antennanp ANTENNA_76 (.A(_02959_));
 sg13g2_antennanp ANTENNA_77 (.A(_02975_));
 sg13g2_antennanp ANTENNA_78 (.A(_02975_));
 sg13g2_antennanp ANTENNA_79 (.A(_02988_));
 sg13g2_antennanp ANTENNA_80 (.A(_02989_));
 sg13g2_antennanp ANTENNA_81 (.A(_02992_));
 sg13g2_antennanp ANTENNA_82 (.A(_02993_));
 sg13g2_antennanp ANTENNA_83 (.A(_03064_));
 sg13g2_antennanp ANTENNA_84 (.A(_03064_));
 sg13g2_antennanp ANTENNA_85 (.A(_03071_));
 sg13g2_antennanp ANTENNA_86 (.A(_03071_));
 sg13g2_antennanp ANTENNA_87 (.A(_03071_));
 sg13g2_antennanp ANTENNA_88 (.A(_03074_));
 sg13g2_antennanp ANTENNA_89 (.A(_03074_));
 sg13g2_antennanp ANTENNA_90 (.A(_03078_));
 sg13g2_antennanp ANTENNA_91 (.A(_03078_));
 sg13g2_antennanp ANTENNA_92 (.A(_03078_));
 sg13g2_antennanp ANTENNA_93 (.A(_03078_));
 sg13g2_antennanp ANTENNA_94 (.A(_03078_));
 sg13g2_antennanp ANTENNA_95 (.A(_03078_));
 sg13g2_antennanp ANTENNA_96 (.A(_03078_));
 sg13g2_antennanp ANTENNA_97 (.A(_03078_));
 sg13g2_antennanp ANTENNA_98 (.A(_03082_));
 sg13g2_antennanp ANTENNA_99 (.A(_03082_));
 sg13g2_antennanp ANTENNA_100 (.A(_03082_));
 sg13g2_antennanp ANTENNA_101 (.A(_03083_));
 sg13g2_antennanp ANTENNA_102 (.A(_03083_));
 sg13g2_antennanp ANTENNA_103 (.A(_03083_));
 sg13g2_antennanp ANTENNA_104 (.A(_03083_));
 sg13g2_antennanp ANTENNA_105 (.A(_03083_));
 sg13g2_antennanp ANTENNA_106 (.A(_03083_));
 sg13g2_antennanp ANTENNA_107 (.A(_03083_));
 sg13g2_antennanp ANTENNA_108 (.A(_03083_));
 sg13g2_antennanp ANTENNA_109 (.A(_03085_));
 sg13g2_antennanp ANTENNA_110 (.A(_03085_));
 sg13g2_antennanp ANTENNA_111 (.A(_03085_));
 sg13g2_antennanp ANTENNA_112 (.A(_03086_));
 sg13g2_antennanp ANTENNA_113 (.A(_03086_));
 sg13g2_antennanp ANTENNA_114 (.A(_03086_));
 sg13g2_antennanp ANTENNA_115 (.A(_03086_));
 sg13g2_antennanp ANTENNA_116 (.A(_03089_));
 sg13g2_antennanp ANTENNA_117 (.A(_03089_));
 sg13g2_antennanp ANTENNA_118 (.A(_03089_));
 sg13g2_antennanp ANTENNA_119 (.A(_03096_));
 sg13g2_antennanp ANTENNA_120 (.A(_03096_));
 sg13g2_antennanp ANTENNA_121 (.A(_03096_));
 sg13g2_antennanp ANTENNA_122 (.A(_03104_));
 sg13g2_antennanp ANTENNA_123 (.A(_03104_));
 sg13g2_antennanp ANTENNA_124 (.A(_03104_));
 sg13g2_antennanp ANTENNA_125 (.A(_03166_));
 sg13g2_antennanp ANTENNA_126 (.A(_03166_));
 sg13g2_antennanp ANTENNA_127 (.A(_03166_));
 sg13g2_antennanp ANTENNA_128 (.A(_03166_));
 sg13g2_antennanp ANTENNA_129 (.A(_03166_));
 sg13g2_antennanp ANTENNA_130 (.A(_03166_));
 sg13g2_antennanp ANTENNA_131 (.A(_03166_));
 sg13g2_antennanp ANTENNA_132 (.A(_03166_));
 sg13g2_antennanp ANTENNA_133 (.A(_03166_));
 sg13g2_antennanp ANTENNA_134 (.A(_03318_));
 sg13g2_antennanp ANTENNA_135 (.A(_03318_));
 sg13g2_antennanp ANTENNA_136 (.A(_03318_));
 sg13g2_antennanp ANTENNA_137 (.A(_03592_));
 sg13g2_antennanp ANTENNA_138 (.A(_03592_));
 sg13g2_antennanp ANTENNA_139 (.A(_03592_));
 sg13g2_antennanp ANTENNA_140 (.A(_03592_));
 sg13g2_antennanp ANTENNA_141 (.A(_03592_));
 sg13g2_antennanp ANTENNA_142 (.A(_03592_));
 sg13g2_antennanp ANTENNA_143 (.A(_03592_));
 sg13g2_antennanp ANTENNA_144 (.A(_03592_));
 sg13g2_antennanp ANTENNA_145 (.A(_03592_));
 sg13g2_antennanp ANTENNA_146 (.A(_03613_));
 sg13g2_antennanp ANTENNA_147 (.A(_03613_));
 sg13g2_antennanp ANTENNA_148 (.A(_03613_));
 sg13g2_antennanp ANTENNA_149 (.A(_03613_));
 sg13g2_antennanp ANTENNA_150 (.A(_03644_));
 sg13g2_antennanp ANTENNA_151 (.A(_03644_));
 sg13g2_antennanp ANTENNA_152 (.A(_03644_));
 sg13g2_antennanp ANTENNA_153 (.A(_03663_));
 sg13g2_antennanp ANTENNA_154 (.A(_03663_));
 sg13g2_antennanp ANTENNA_155 (.A(_03663_));
 sg13g2_antennanp ANTENNA_156 (.A(_03663_));
 sg13g2_antennanp ANTENNA_157 (.A(_03663_));
 sg13g2_antennanp ANTENNA_158 (.A(_03695_));
 sg13g2_antennanp ANTENNA_159 (.A(_03695_));
 sg13g2_antennanp ANTENNA_160 (.A(_03695_));
 sg13g2_antennanp ANTENNA_161 (.A(_03695_));
 sg13g2_antennanp ANTENNA_162 (.A(_03695_));
 sg13g2_antennanp ANTENNA_163 (.A(_03695_));
 sg13g2_antennanp ANTENNA_164 (.A(_03695_));
 sg13g2_antennanp ANTENNA_165 (.A(_03695_));
 sg13g2_antennanp ANTENNA_166 (.A(_03695_));
 sg13g2_antennanp ANTENNA_167 (.A(_03695_));
 sg13g2_antennanp ANTENNA_168 (.A(_03954_));
 sg13g2_antennanp ANTENNA_169 (.A(_03954_));
 sg13g2_antennanp ANTENNA_170 (.A(_03954_));
 sg13g2_antennanp ANTENNA_171 (.A(_03954_));
 sg13g2_antennanp ANTENNA_172 (.A(_04044_));
 sg13g2_antennanp ANTENNA_173 (.A(_04044_));
 sg13g2_antennanp ANTENNA_174 (.A(_04044_));
 sg13g2_antennanp ANTENNA_175 (.A(_04044_));
 sg13g2_antennanp ANTENNA_176 (.A(_04044_));
 sg13g2_antennanp ANTENNA_177 (.A(_04044_));
 sg13g2_antennanp ANTENNA_178 (.A(_04044_));
 sg13g2_antennanp ANTENNA_179 (.A(_04044_));
 sg13g2_antennanp ANTENNA_180 (.A(_04044_));
 sg13g2_antennanp ANTENNA_181 (.A(_04044_));
 sg13g2_antennanp ANTENNA_182 (.A(_04044_));
 sg13g2_antennanp ANTENNA_183 (.A(_04044_));
 sg13g2_antennanp ANTENNA_184 (.A(_04048_));
 sg13g2_antennanp ANTENNA_185 (.A(_04048_));
 sg13g2_antennanp ANTENNA_186 (.A(_04048_));
 sg13g2_antennanp ANTENNA_187 (.A(_04048_));
 sg13g2_antennanp ANTENNA_188 (.A(_04051_));
 sg13g2_antennanp ANTENNA_189 (.A(_04051_));
 sg13g2_antennanp ANTENNA_190 (.A(_04051_));
 sg13g2_antennanp ANTENNA_191 (.A(_04051_));
 sg13g2_antennanp ANTENNA_192 (.A(_04064_));
 sg13g2_antennanp ANTENNA_193 (.A(_04064_));
 sg13g2_antennanp ANTENNA_194 (.A(_04064_));
 sg13g2_antennanp ANTENNA_195 (.A(_04064_));
 sg13g2_antennanp ANTENNA_196 (.A(_04243_));
 sg13g2_antennanp ANTENNA_197 (.A(_04243_));
 sg13g2_antennanp ANTENNA_198 (.A(_04243_));
 sg13g2_antennanp ANTENNA_199 (.A(_04243_));
 sg13g2_antennanp ANTENNA_200 (.A(_04255_));
 sg13g2_antennanp ANTENNA_201 (.A(_04255_));
 sg13g2_antennanp ANTENNA_202 (.A(_04255_));
 sg13g2_antennanp ANTENNA_203 (.A(_04255_));
 sg13g2_antennanp ANTENNA_204 (.A(_04255_));
 sg13g2_antennanp ANTENNA_205 (.A(_04255_));
 sg13g2_antennanp ANTENNA_206 (.A(_04255_));
 sg13g2_antennanp ANTENNA_207 (.A(_04255_));
 sg13g2_antennanp ANTENNA_208 (.A(_04263_));
 sg13g2_antennanp ANTENNA_209 (.A(_04263_));
 sg13g2_antennanp ANTENNA_210 (.A(_04263_));
 sg13g2_antennanp ANTENNA_211 (.A(_04263_));
 sg13g2_antennanp ANTENNA_212 (.A(_04263_));
 sg13g2_antennanp ANTENNA_213 (.A(_04263_));
 sg13g2_antennanp ANTENNA_214 (.A(_04263_));
 sg13g2_antennanp ANTENNA_215 (.A(_04263_));
 sg13g2_antennanp ANTENNA_216 (.A(_04263_));
 sg13g2_antennanp ANTENNA_217 (.A(_04263_));
 sg13g2_antennanp ANTENNA_218 (.A(_04286_));
 sg13g2_antennanp ANTENNA_219 (.A(_04286_));
 sg13g2_antennanp ANTENNA_220 (.A(_04286_));
 sg13g2_antennanp ANTENNA_221 (.A(_04348_));
 sg13g2_antennanp ANTENNA_222 (.A(_04348_));
 sg13g2_antennanp ANTENNA_223 (.A(_04348_));
 sg13g2_antennanp ANTENNA_224 (.A(_04348_));
 sg13g2_antennanp ANTENNA_225 (.A(_04485_));
 sg13g2_antennanp ANTENNA_226 (.A(_04485_));
 sg13g2_antennanp ANTENNA_227 (.A(_04485_));
 sg13g2_antennanp ANTENNA_228 (.A(_04485_));
 sg13g2_antennanp ANTENNA_229 (.A(_05084_));
 sg13g2_antennanp ANTENNA_230 (.A(_05084_));
 sg13g2_antennanp ANTENNA_231 (.A(_05084_));
 sg13g2_antennanp ANTENNA_232 (.A(_05090_));
 sg13g2_antennanp ANTENNA_233 (.A(_05090_));
 sg13g2_antennanp ANTENNA_234 (.A(_05090_));
 sg13g2_antennanp ANTENNA_235 (.A(_05090_));
 sg13g2_antennanp ANTENNA_236 (.A(_05111_));
 sg13g2_antennanp ANTENNA_237 (.A(_05111_));
 sg13g2_antennanp ANTENNA_238 (.A(_05111_));
 sg13g2_antennanp ANTENNA_239 (.A(_05111_));
 sg13g2_antennanp ANTENNA_240 (.A(_05111_));
 sg13g2_antennanp ANTENNA_241 (.A(_05111_));
 sg13g2_antennanp ANTENNA_242 (.A(_05111_));
 sg13g2_antennanp ANTENNA_243 (.A(_05111_));
 sg13g2_antennanp ANTENNA_244 (.A(_05111_));
 sg13g2_antennanp ANTENNA_245 (.A(_05111_));
 sg13g2_antennanp ANTENNA_246 (.A(_05828_));
 sg13g2_antennanp ANTENNA_247 (.A(_05828_));
 sg13g2_antennanp ANTENNA_248 (.A(_05828_));
 sg13g2_antennanp ANTENNA_249 (.A(_05828_));
 sg13g2_antennanp ANTENNA_250 (.A(_05828_));
 sg13g2_antennanp ANTENNA_251 (.A(_05828_));
 sg13g2_antennanp ANTENNA_252 (.A(_05828_));
 sg13g2_antennanp ANTENNA_253 (.A(_07381_));
 sg13g2_antennanp ANTENNA_254 (.A(_07381_));
 sg13g2_antennanp ANTENNA_255 (.A(_07381_));
 sg13g2_antennanp ANTENNA_256 (.A(_07412_));
 sg13g2_antennanp ANTENNA_257 (.A(_07412_));
 sg13g2_antennanp ANTENNA_258 (.A(_07412_));
 sg13g2_antennanp ANTENNA_259 (.A(_07412_));
 sg13g2_antennanp ANTENNA_260 (.A(_08176_));
 sg13g2_antennanp ANTENNA_261 (.A(_08176_));
 sg13g2_antennanp ANTENNA_262 (.A(_08176_));
 sg13g2_antennanp ANTENNA_263 (.A(_08176_));
 sg13g2_antennanp ANTENNA_264 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_265 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_266 (.A(\b.gen_square[5].sq.piece[2] ));
 sg13g2_antennanp ANTENNA_267 (.A(\b.gen_square[5].sq.piece[2] ));
 sg13g2_antennanp ANTENNA_268 (.A(clk));
 sg13g2_antennanp ANTENNA_269 (.A(net63));
 sg13g2_antennanp ANTENNA_270 (.A(net63));
 sg13g2_antennanp ANTENNA_271 (.A(net63));
 sg13g2_antennanp ANTENNA_272 (.A(net63));
 sg13g2_antennanp ANTENNA_273 (.A(net63));
 sg13g2_antennanp ANTENNA_274 (.A(net63));
 sg13g2_antennanp ANTENNA_275 (.A(net63));
 sg13g2_antennanp ANTENNA_276 (.A(net63));
 sg13g2_antennanp ANTENNA_277 (.A(net72));
 sg13g2_antennanp ANTENNA_278 (.A(net72));
 sg13g2_antennanp ANTENNA_279 (.A(net72));
 sg13g2_antennanp ANTENNA_280 (.A(net72));
 sg13g2_antennanp ANTENNA_281 (.A(net72));
 sg13g2_antennanp ANTENNA_282 (.A(net72));
 sg13g2_antennanp ANTENNA_283 (.A(net72));
 sg13g2_antennanp ANTENNA_284 (.A(net72));
 sg13g2_antennanp ANTENNA_285 (.A(net72));
 sg13g2_antennanp ANTENNA_286 (.A(net86));
 sg13g2_antennanp ANTENNA_287 (.A(net86));
 sg13g2_antennanp ANTENNA_288 (.A(net86));
 sg13g2_antennanp ANTENNA_289 (.A(net86));
 sg13g2_antennanp ANTENNA_290 (.A(net86));
 sg13g2_antennanp ANTENNA_291 (.A(net86));
 sg13g2_antennanp ANTENNA_292 (.A(net86));
 sg13g2_antennanp ANTENNA_293 (.A(net86));
 sg13g2_antennanp ANTENNA_294 (.A(net86));
 sg13g2_antennanp ANTENNA_295 (.A(net86));
 sg13g2_antennanp ANTENNA_296 (.A(net86));
 sg13g2_antennanp ANTENNA_297 (.A(net86));
 sg13g2_antennanp ANTENNA_298 (.A(net86));
 sg13g2_antennanp ANTENNA_299 (.A(net86));
 sg13g2_antennanp ANTENNA_300 (.A(net86));
 sg13g2_antennanp ANTENNA_301 (.A(net86));
 sg13g2_antennanp ANTENNA_302 (.A(net86));
 sg13g2_antennanp ANTENNA_303 (.A(net86));
 sg13g2_antennanp ANTENNA_304 (.A(net86));
 sg13g2_antennanp ANTENNA_305 (.A(net86));
 sg13g2_antennanp ANTENNA_306 (.A(net86));
 sg13g2_antennanp ANTENNA_307 (.A(net93));
 sg13g2_antennanp ANTENNA_308 (.A(net93));
 sg13g2_antennanp ANTENNA_309 (.A(net93));
 sg13g2_antennanp ANTENNA_310 (.A(net93));
 sg13g2_antennanp ANTENNA_311 (.A(net93));
 sg13g2_antennanp ANTENNA_312 (.A(net93));
 sg13g2_antennanp ANTENNA_313 (.A(net93));
 sg13g2_antennanp ANTENNA_314 (.A(net93));
 sg13g2_antennanp ANTENNA_315 (.A(net93));
 sg13g2_antennanp ANTENNA_316 (.A(net93));
 sg13g2_antennanp ANTENNA_317 (.A(net93));
 sg13g2_antennanp ANTENNA_318 (.A(net93));
 sg13g2_antennanp ANTENNA_319 (.A(net93));
 sg13g2_antennanp ANTENNA_320 (.A(net93));
 sg13g2_antennanp ANTENNA_321 (.A(net93));
 sg13g2_antennanp ANTENNA_322 (.A(net93));
 sg13g2_antennanp ANTENNA_323 (.A(net93));
 sg13g2_antennanp ANTENNA_324 (.A(net93));
 sg13g2_antennanp ANTENNA_325 (.A(net93));
 sg13g2_antennanp ANTENNA_326 (.A(net93));
 sg13g2_antennanp ANTENNA_327 (.A(net93));
 sg13g2_antennanp ANTENNA_328 (.A(net93));
 sg13g2_antennanp ANTENNA_329 (.A(net93));
 sg13g2_antennanp ANTENNA_330 (.A(net93));
 sg13g2_antennanp ANTENNA_331 (.A(net96));
 sg13g2_antennanp ANTENNA_332 (.A(net96));
 sg13g2_antennanp ANTENNA_333 (.A(net96));
 sg13g2_antennanp ANTENNA_334 (.A(net96));
 sg13g2_antennanp ANTENNA_335 (.A(net96));
 sg13g2_antennanp ANTENNA_336 (.A(net96));
 sg13g2_antennanp ANTENNA_337 (.A(net96));
 sg13g2_antennanp ANTENNA_338 (.A(net96));
 sg13g2_antennanp ANTENNA_339 (.A(net96));
 sg13g2_antennanp ANTENNA_340 (.A(net96));
 sg13g2_antennanp ANTENNA_341 (.A(net96));
 sg13g2_antennanp ANTENNA_342 (.A(net96));
 sg13g2_antennanp ANTENNA_343 (.A(net96));
 sg13g2_antennanp ANTENNA_344 (.A(net96));
 sg13g2_antennanp ANTENNA_345 (.A(net96));
 sg13g2_antennanp ANTENNA_346 (.A(net96));
 sg13g2_antennanp ANTENNA_347 (.A(net96));
 sg13g2_antennanp ANTENNA_348 (.A(net96));
 sg13g2_antennanp ANTENNA_349 (.A(net106));
 sg13g2_antennanp ANTENNA_350 (.A(net106));
 sg13g2_antennanp ANTENNA_351 (.A(net106));
 sg13g2_antennanp ANTENNA_352 (.A(net106));
 sg13g2_antennanp ANTENNA_353 (.A(net106));
 sg13g2_antennanp ANTENNA_354 (.A(net106));
 sg13g2_antennanp ANTENNA_355 (.A(net106));
 sg13g2_antennanp ANTENNA_356 (.A(net106));
 sg13g2_antennanp ANTENNA_357 (.A(net106));
 sg13g2_antennanp ANTENNA_358 (.A(net106));
 sg13g2_antennanp ANTENNA_359 (.A(net106));
 sg13g2_antennanp ANTENNA_360 (.A(net112));
 sg13g2_antennanp ANTENNA_361 (.A(net112));
 sg13g2_antennanp ANTENNA_362 (.A(net112));
 sg13g2_antennanp ANTENNA_363 (.A(net112));
 sg13g2_antennanp ANTENNA_364 (.A(net112));
 sg13g2_antennanp ANTENNA_365 (.A(net112));
 sg13g2_antennanp ANTENNA_366 (.A(net112));
 sg13g2_antennanp ANTENNA_367 (.A(net112));
 sg13g2_antennanp ANTENNA_368 (.A(net112));
 sg13g2_antennanp ANTENNA_369 (.A(net124));
 sg13g2_antennanp ANTENNA_370 (.A(net124));
 sg13g2_antennanp ANTENNA_371 (.A(net124));
 sg13g2_antennanp ANTENNA_372 (.A(net124));
 sg13g2_antennanp ANTENNA_373 (.A(net124));
 sg13g2_antennanp ANTENNA_374 (.A(net124));
 sg13g2_antennanp ANTENNA_375 (.A(net124));
 sg13g2_antennanp ANTENNA_376 (.A(net124));
 sg13g2_antennanp ANTENNA_377 (.A(net124));
 sg13g2_antennanp ANTENNA_378 (.A(net124));
 sg13g2_antennanp ANTENNA_379 (.A(net124));
 sg13g2_antennanp ANTENNA_380 (.A(net124));
 sg13g2_antennanp ANTENNA_381 (.A(net124));
 sg13g2_antennanp ANTENNA_382 (.A(net124));
 sg13g2_antennanp ANTENNA_383 (.A(net124));
 sg13g2_antennanp ANTENNA_384 (.A(net124));
 sg13g2_antennanp ANTENNA_385 (.A(net155));
 sg13g2_antennanp ANTENNA_386 (.A(net155));
 sg13g2_antennanp ANTENNA_387 (.A(net155));
 sg13g2_antennanp ANTENNA_388 (.A(net155));
 sg13g2_antennanp ANTENNA_389 (.A(net155));
 sg13g2_antennanp ANTENNA_390 (.A(net155));
 sg13g2_antennanp ANTENNA_391 (.A(net155));
 sg13g2_antennanp ANTENNA_392 (.A(net155));
 sg13g2_antennanp ANTENNA_393 (.A(net155));
 sg13g2_antennanp ANTENNA_394 (.A(net155));
 sg13g2_antennanp ANTENNA_395 (.A(net155));
 sg13g2_antennanp ANTENNA_396 (.A(net158));
 sg13g2_antennanp ANTENNA_397 (.A(net158));
 sg13g2_antennanp ANTENNA_398 (.A(net158));
 sg13g2_antennanp ANTENNA_399 (.A(net158));
 sg13g2_antennanp ANTENNA_400 (.A(net158));
 sg13g2_antennanp ANTENNA_401 (.A(net158));
 sg13g2_antennanp ANTENNA_402 (.A(net158));
 sg13g2_antennanp ANTENNA_403 (.A(net158));
 sg13g2_antennanp ANTENNA_404 (.A(net158));
 sg13g2_antennanp ANTENNA_405 (.A(net292));
 sg13g2_antennanp ANTENNA_406 (.A(net292));
 sg13g2_antennanp ANTENNA_407 (.A(net292));
 sg13g2_antennanp ANTENNA_408 (.A(net292));
 sg13g2_antennanp ANTENNA_409 (.A(net292));
 sg13g2_antennanp ANTENNA_410 (.A(net292));
 sg13g2_antennanp ANTENNA_411 (.A(net292));
 sg13g2_antennanp ANTENNA_412 (.A(net292));
 sg13g2_antennanp ANTENNA_413 (.A(net292));
 sg13g2_antennanp ANTENNA_414 (.A(_00631_));
 sg13g2_antennanp ANTENNA_415 (.A(_01231_));
 sg13g2_antennanp ANTENNA_416 (.A(_01231_));
 sg13g2_antennanp ANTENNA_417 (.A(_01231_));
 sg13g2_antennanp ANTENNA_418 (.A(_01231_));
 sg13g2_antennanp ANTENNA_419 (.A(_01968_));
 sg13g2_antennanp ANTENNA_420 (.A(_01968_));
 sg13g2_antennanp ANTENNA_421 (.A(_01968_));
 sg13g2_antennanp ANTENNA_422 (.A(_01968_));
 sg13g2_antennanp ANTENNA_423 (.A(_01968_));
 sg13g2_antennanp ANTENNA_424 (.A(_01968_));
 sg13g2_antennanp ANTENNA_425 (.A(_01968_));
 sg13g2_antennanp ANTENNA_426 (.A(_01968_));
 sg13g2_antennanp ANTENNA_427 (.A(_01968_));
 sg13g2_antennanp ANTENNA_428 (.A(_01968_));
 sg13g2_antennanp ANTENNA_429 (.A(_01968_));
 sg13g2_antennanp ANTENNA_430 (.A(_01968_));
 sg13g2_antennanp ANTENNA_431 (.A(_01968_));
 sg13g2_antennanp ANTENNA_432 (.A(_01968_));
 sg13g2_antennanp ANTENNA_433 (.A(_01968_));
 sg13g2_antennanp ANTENNA_434 (.A(_01968_));
 sg13g2_antennanp ANTENNA_435 (.A(_02012_));
 sg13g2_antennanp ANTENNA_436 (.A(_02012_));
 sg13g2_antennanp ANTENNA_437 (.A(_02012_));
 sg13g2_antennanp ANTENNA_438 (.A(_02012_));
 sg13g2_antennanp ANTENNA_439 (.A(_02067_));
 sg13g2_antennanp ANTENNA_440 (.A(_02067_));
 sg13g2_antennanp ANTENNA_441 (.A(_02067_));
 sg13g2_antennanp ANTENNA_442 (.A(_02078_));
 sg13g2_antennanp ANTENNA_443 (.A(_02078_));
 sg13g2_antennanp ANTENNA_444 (.A(_02078_));
 sg13g2_antennanp ANTENNA_445 (.A(_02078_));
 sg13g2_antennanp ANTENNA_446 (.A(_02078_));
 sg13g2_antennanp ANTENNA_447 (.A(_02078_));
 sg13g2_antennanp ANTENNA_448 (.A(_02078_));
 sg13g2_antennanp ANTENNA_449 (.A(_02242_));
 sg13g2_antennanp ANTENNA_450 (.A(_02242_));
 sg13g2_antennanp ANTENNA_451 (.A(_02296_));
 sg13g2_antennanp ANTENNA_452 (.A(_02296_));
 sg13g2_antennanp ANTENNA_453 (.A(_02296_));
 sg13g2_antennanp ANTENNA_454 (.A(_02350_));
 sg13g2_antennanp ANTENNA_455 (.A(_02350_));
 sg13g2_antennanp ANTENNA_456 (.A(_02350_));
 sg13g2_antennanp ANTENNA_457 (.A(_02350_));
 sg13g2_antennanp ANTENNA_458 (.A(_02807_));
 sg13g2_antennanp ANTENNA_459 (.A(_02807_));
 sg13g2_antennanp ANTENNA_460 (.A(_02899_));
 sg13g2_antennanp ANTENNA_461 (.A(_02899_));
 sg13g2_antennanp ANTENNA_462 (.A(_02902_));
 sg13g2_antennanp ANTENNA_463 (.A(_02906_));
 sg13g2_antennanp ANTENNA_464 (.A(_02914_));
 sg13g2_antennanp ANTENNA_465 (.A(_02919_));
 sg13g2_antennanp ANTENNA_466 (.A(_02921_));
 sg13g2_antennanp ANTENNA_467 (.A(_02948_));
 sg13g2_antennanp ANTENNA_468 (.A(_02953_));
 sg13g2_antennanp ANTENNA_469 (.A(_02954_));
 sg13g2_antennanp ANTENNA_470 (.A(_02957_));
 sg13g2_antennanp ANTENNA_471 (.A(_02959_));
 sg13g2_antennanp ANTENNA_472 (.A(_02975_));
 sg13g2_antennanp ANTENNA_473 (.A(_02988_));
 sg13g2_antennanp ANTENNA_474 (.A(_02989_));
 sg13g2_antennanp ANTENNA_475 (.A(_02992_));
 sg13g2_antennanp ANTENNA_476 (.A(_02993_));
 sg13g2_antennanp ANTENNA_477 (.A(_03064_));
 sg13g2_antennanp ANTENNA_478 (.A(_03064_));
 sg13g2_antennanp ANTENNA_479 (.A(_03071_));
 sg13g2_antennanp ANTENNA_480 (.A(_03071_));
 sg13g2_antennanp ANTENNA_481 (.A(_03071_));
 sg13g2_antennanp ANTENNA_482 (.A(_03071_));
 sg13g2_antennanp ANTENNA_483 (.A(_03071_));
 sg13g2_antennanp ANTENNA_484 (.A(_03071_));
 sg13g2_antennanp ANTENNA_485 (.A(_03071_));
 sg13g2_antennanp ANTENNA_486 (.A(_03071_));
 sg13g2_antennanp ANTENNA_487 (.A(_03071_));
 sg13g2_antennanp ANTENNA_488 (.A(_03071_));
 sg13g2_antennanp ANTENNA_489 (.A(_03074_));
 sg13g2_antennanp ANTENNA_490 (.A(_03074_));
 sg13g2_antennanp ANTENNA_491 (.A(_03074_));
 sg13g2_antennanp ANTENNA_492 (.A(_03078_));
 sg13g2_antennanp ANTENNA_493 (.A(_03078_));
 sg13g2_antennanp ANTENNA_494 (.A(_03078_));
 sg13g2_antennanp ANTENNA_495 (.A(_03078_));
 sg13g2_antennanp ANTENNA_496 (.A(_03078_));
 sg13g2_antennanp ANTENNA_497 (.A(_03078_));
 sg13g2_antennanp ANTENNA_498 (.A(_03078_));
 sg13g2_antennanp ANTENNA_499 (.A(_03078_));
 sg13g2_antennanp ANTENNA_500 (.A(_03078_));
 sg13g2_antennanp ANTENNA_501 (.A(_03078_));
 sg13g2_antennanp ANTENNA_502 (.A(_03082_));
 sg13g2_antennanp ANTENNA_503 (.A(_03082_));
 sg13g2_antennanp ANTENNA_504 (.A(_03082_));
 sg13g2_antennanp ANTENNA_505 (.A(_03086_));
 sg13g2_antennanp ANTENNA_506 (.A(_03086_));
 sg13g2_antennanp ANTENNA_507 (.A(_03086_));
 sg13g2_antennanp ANTENNA_508 (.A(_03086_));
 sg13g2_antennanp ANTENNA_509 (.A(_03089_));
 sg13g2_antennanp ANTENNA_510 (.A(_03089_));
 sg13g2_antennanp ANTENNA_511 (.A(_03089_));
 sg13g2_antennanp ANTENNA_512 (.A(_03089_));
 sg13g2_antennanp ANTENNA_513 (.A(_03089_));
 sg13g2_antennanp ANTENNA_514 (.A(_03089_));
 sg13g2_antennanp ANTENNA_515 (.A(_03089_));
 sg13g2_antennanp ANTENNA_516 (.A(_03089_));
 sg13g2_antennanp ANTENNA_517 (.A(_03096_));
 sg13g2_antennanp ANTENNA_518 (.A(_03096_));
 sg13g2_antennanp ANTENNA_519 (.A(_03096_));
 sg13g2_antennanp ANTENNA_520 (.A(_03104_));
 sg13g2_antennanp ANTENNA_521 (.A(_03104_));
 sg13g2_antennanp ANTENNA_522 (.A(_03104_));
 sg13g2_antennanp ANTENNA_523 (.A(_03166_));
 sg13g2_antennanp ANTENNA_524 (.A(_03166_));
 sg13g2_antennanp ANTENNA_525 (.A(_03166_));
 sg13g2_antennanp ANTENNA_526 (.A(_03166_));
 sg13g2_antennanp ANTENNA_527 (.A(_03318_));
 sg13g2_antennanp ANTENNA_528 (.A(_03318_));
 sg13g2_antennanp ANTENNA_529 (.A(_03318_));
 sg13g2_antennanp ANTENNA_530 (.A(_03592_));
 sg13g2_antennanp ANTENNA_531 (.A(_03592_));
 sg13g2_antennanp ANTENNA_532 (.A(_03592_));
 sg13g2_antennanp ANTENNA_533 (.A(_03592_));
 sg13g2_antennanp ANTENNA_534 (.A(_03592_));
 sg13g2_antennanp ANTENNA_535 (.A(_03592_));
 sg13g2_antennanp ANTENNA_536 (.A(_03592_));
 sg13g2_antennanp ANTENNA_537 (.A(_03592_));
 sg13g2_antennanp ANTENNA_538 (.A(_03592_));
 sg13g2_antennanp ANTENNA_539 (.A(_03592_));
 sg13g2_antennanp ANTENNA_540 (.A(_03592_));
 sg13g2_antennanp ANTENNA_541 (.A(_03592_));
 sg13g2_antennanp ANTENNA_542 (.A(_03592_));
 sg13g2_antennanp ANTENNA_543 (.A(_03592_));
 sg13g2_antennanp ANTENNA_544 (.A(_03592_));
 sg13g2_antennanp ANTENNA_545 (.A(_03592_));
 sg13g2_antennanp ANTENNA_546 (.A(_03644_));
 sg13g2_antennanp ANTENNA_547 (.A(_03644_));
 sg13g2_antennanp ANTENNA_548 (.A(_03644_));
 sg13g2_antennanp ANTENNA_549 (.A(_03663_));
 sg13g2_antennanp ANTENNA_550 (.A(_03663_));
 sg13g2_antennanp ANTENNA_551 (.A(_03663_));
 sg13g2_antennanp ANTENNA_552 (.A(_03663_));
 sg13g2_antennanp ANTENNA_553 (.A(_03663_));
 sg13g2_antennanp ANTENNA_554 (.A(_03695_));
 sg13g2_antennanp ANTENNA_555 (.A(_03695_));
 sg13g2_antennanp ANTENNA_556 (.A(_03695_));
 sg13g2_antennanp ANTENNA_557 (.A(_03695_));
 sg13g2_antennanp ANTENNA_558 (.A(_03695_));
 sg13g2_antennanp ANTENNA_559 (.A(_03695_));
 sg13g2_antennanp ANTENNA_560 (.A(_03954_));
 sg13g2_antennanp ANTENNA_561 (.A(_03954_));
 sg13g2_antennanp ANTENNA_562 (.A(_03954_));
 sg13g2_antennanp ANTENNA_563 (.A(_04044_));
 sg13g2_antennanp ANTENNA_564 (.A(_04044_));
 sg13g2_antennanp ANTENNA_565 (.A(_04044_));
 sg13g2_antennanp ANTENNA_566 (.A(_04044_));
 sg13g2_antennanp ANTENNA_567 (.A(_04044_));
 sg13g2_antennanp ANTENNA_568 (.A(_04044_));
 sg13g2_antennanp ANTENNA_569 (.A(_04044_));
 sg13g2_antennanp ANTENNA_570 (.A(_04044_));
 sg13g2_antennanp ANTENNA_571 (.A(_04044_));
 sg13g2_antennanp ANTENNA_572 (.A(_04044_));
 sg13g2_antennanp ANTENNA_573 (.A(_04044_));
 sg13g2_antennanp ANTENNA_574 (.A(_04044_));
 sg13g2_antennanp ANTENNA_575 (.A(_04048_));
 sg13g2_antennanp ANTENNA_576 (.A(_04048_));
 sg13g2_antennanp ANTENNA_577 (.A(_04048_));
 sg13g2_antennanp ANTENNA_578 (.A(_04048_));
 sg13g2_antennanp ANTENNA_579 (.A(_04064_));
 sg13g2_antennanp ANTENNA_580 (.A(_04064_));
 sg13g2_antennanp ANTENNA_581 (.A(_04064_));
 sg13g2_antennanp ANTENNA_582 (.A(_04064_));
 sg13g2_antennanp ANTENNA_583 (.A(_04243_));
 sg13g2_antennanp ANTENNA_584 (.A(_04243_));
 sg13g2_antennanp ANTENNA_585 (.A(_04243_));
 sg13g2_antennanp ANTENNA_586 (.A(_04243_));
 sg13g2_antennanp ANTENNA_587 (.A(_04263_));
 sg13g2_antennanp ANTENNA_588 (.A(_04263_));
 sg13g2_antennanp ANTENNA_589 (.A(_04263_));
 sg13g2_antennanp ANTENNA_590 (.A(_04263_));
 sg13g2_antennanp ANTENNA_591 (.A(_04263_));
 sg13g2_antennanp ANTENNA_592 (.A(_04263_));
 sg13g2_antennanp ANTENNA_593 (.A(_04286_));
 sg13g2_antennanp ANTENNA_594 (.A(_04286_));
 sg13g2_antennanp ANTENNA_595 (.A(_04286_));
 sg13g2_antennanp ANTENNA_596 (.A(_04286_));
 sg13g2_antennanp ANTENNA_597 (.A(_04286_));
 sg13g2_antennanp ANTENNA_598 (.A(_04287_));
 sg13g2_antennanp ANTENNA_599 (.A(_04287_));
 sg13g2_antennanp ANTENNA_600 (.A(_04287_));
 sg13g2_antennanp ANTENNA_601 (.A(_04287_));
 sg13g2_antennanp ANTENNA_602 (.A(_04287_));
 sg13g2_antennanp ANTENNA_603 (.A(_04348_));
 sg13g2_antennanp ANTENNA_604 (.A(_04348_));
 sg13g2_antennanp ANTENNA_605 (.A(_04348_));
 sg13g2_antennanp ANTENNA_606 (.A(_04348_));
 sg13g2_antennanp ANTENNA_607 (.A(_04485_));
 sg13g2_antennanp ANTENNA_608 (.A(_04485_));
 sg13g2_antennanp ANTENNA_609 (.A(_04485_));
 sg13g2_antennanp ANTENNA_610 (.A(_04485_));
 sg13g2_antennanp ANTENNA_611 (.A(_04485_));
 sg13g2_antennanp ANTENNA_612 (.A(_04485_));
 sg13g2_antennanp ANTENNA_613 (.A(_04485_));
 sg13g2_antennanp ANTENNA_614 (.A(_04485_));
 sg13g2_antennanp ANTENNA_615 (.A(_05084_));
 sg13g2_antennanp ANTENNA_616 (.A(_05084_));
 sg13g2_antennanp ANTENNA_617 (.A(_05084_));
 sg13g2_antennanp ANTENNA_618 (.A(_05084_));
 sg13g2_antennanp ANTENNA_619 (.A(_05084_));
 sg13g2_antennanp ANTENNA_620 (.A(_05090_));
 sg13g2_antennanp ANTENNA_621 (.A(_05090_));
 sg13g2_antennanp ANTENNA_622 (.A(_05090_));
 sg13g2_antennanp ANTENNA_623 (.A(_05090_));
 sg13g2_antennanp ANTENNA_624 (.A(_05111_));
 sg13g2_antennanp ANTENNA_625 (.A(_05111_));
 sg13g2_antennanp ANTENNA_626 (.A(_05111_));
 sg13g2_antennanp ANTENNA_627 (.A(_05111_));
 sg13g2_antennanp ANTENNA_628 (.A(_05828_));
 sg13g2_antennanp ANTENNA_629 (.A(_05828_));
 sg13g2_antennanp ANTENNA_630 (.A(_05828_));
 sg13g2_antennanp ANTENNA_631 (.A(_05828_));
 sg13g2_antennanp ANTENNA_632 (.A(_05828_));
 sg13g2_antennanp ANTENNA_633 (.A(_05828_));
 sg13g2_antennanp ANTENNA_634 (.A(_05828_));
 sg13g2_antennanp ANTENNA_635 (.A(_07381_));
 sg13g2_antennanp ANTENNA_636 (.A(_07381_));
 sg13g2_antennanp ANTENNA_637 (.A(_07381_));
 sg13g2_antennanp ANTENNA_638 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_639 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_640 (.A(clk));
 sg13g2_antennanp ANTENNA_641 (.A(net63));
 sg13g2_antennanp ANTENNA_642 (.A(net63));
 sg13g2_antennanp ANTENNA_643 (.A(net63));
 sg13g2_antennanp ANTENNA_644 (.A(net63));
 sg13g2_antennanp ANTENNA_645 (.A(net63));
 sg13g2_antennanp ANTENNA_646 (.A(net63));
 sg13g2_antennanp ANTENNA_647 (.A(net63));
 sg13g2_antennanp ANTENNA_648 (.A(net63));
 sg13g2_antennanp ANTENNA_649 (.A(net72));
 sg13g2_antennanp ANTENNA_650 (.A(net72));
 sg13g2_antennanp ANTENNA_651 (.A(net72));
 sg13g2_antennanp ANTENNA_652 (.A(net72));
 sg13g2_antennanp ANTENNA_653 (.A(net72));
 sg13g2_antennanp ANTENNA_654 (.A(net72));
 sg13g2_antennanp ANTENNA_655 (.A(net72));
 sg13g2_antennanp ANTENNA_656 (.A(net72));
 sg13g2_antennanp ANTENNA_657 (.A(net86));
 sg13g2_antennanp ANTENNA_658 (.A(net86));
 sg13g2_antennanp ANTENNA_659 (.A(net86));
 sg13g2_antennanp ANTENNA_660 (.A(net86));
 sg13g2_antennanp ANTENNA_661 (.A(net86));
 sg13g2_antennanp ANTENNA_662 (.A(net86));
 sg13g2_antennanp ANTENNA_663 (.A(net86));
 sg13g2_antennanp ANTENNA_664 (.A(net86));
 sg13g2_antennanp ANTENNA_665 (.A(net86));
 sg13g2_antennanp ANTENNA_666 (.A(net86));
 sg13g2_antennanp ANTENNA_667 (.A(net86));
 sg13g2_antennanp ANTENNA_668 (.A(net86));
 sg13g2_antennanp ANTENNA_669 (.A(net86));
 sg13g2_antennanp ANTENNA_670 (.A(net86));
 sg13g2_antennanp ANTENNA_671 (.A(net86));
 sg13g2_antennanp ANTENNA_672 (.A(net86));
 sg13g2_antennanp ANTENNA_673 (.A(net86));
 sg13g2_antennanp ANTENNA_674 (.A(net86));
 sg13g2_antennanp ANTENNA_675 (.A(net86));
 sg13g2_antennanp ANTENNA_676 (.A(net86));
 sg13g2_antennanp ANTENNA_677 (.A(net86));
 sg13g2_antennanp ANTENNA_678 (.A(net93));
 sg13g2_antennanp ANTENNA_679 (.A(net93));
 sg13g2_antennanp ANTENNA_680 (.A(net93));
 sg13g2_antennanp ANTENNA_681 (.A(net93));
 sg13g2_antennanp ANTENNA_682 (.A(net93));
 sg13g2_antennanp ANTENNA_683 (.A(net93));
 sg13g2_antennanp ANTENNA_684 (.A(net93));
 sg13g2_antennanp ANTENNA_685 (.A(net93));
 sg13g2_antennanp ANTENNA_686 (.A(net93));
 sg13g2_antennanp ANTENNA_687 (.A(net93));
 sg13g2_antennanp ANTENNA_688 (.A(net93));
 sg13g2_antennanp ANTENNA_689 (.A(net93));
 sg13g2_antennanp ANTENNA_690 (.A(net93));
 sg13g2_antennanp ANTENNA_691 (.A(net93));
 sg13g2_antennanp ANTENNA_692 (.A(net93));
 sg13g2_antennanp ANTENNA_693 (.A(net93));
 sg13g2_antennanp ANTENNA_694 (.A(net93));
 sg13g2_antennanp ANTENNA_695 (.A(net93));
 sg13g2_antennanp ANTENNA_696 (.A(net93));
 sg13g2_antennanp ANTENNA_697 (.A(net93));
 sg13g2_antennanp ANTENNA_698 (.A(net93));
 sg13g2_antennanp ANTENNA_699 (.A(net93));
 sg13g2_antennanp ANTENNA_700 (.A(net93));
 sg13g2_antennanp ANTENNA_701 (.A(net93));
 sg13g2_antennanp ANTENNA_702 (.A(net124));
 sg13g2_antennanp ANTENNA_703 (.A(net124));
 sg13g2_antennanp ANTENNA_704 (.A(net124));
 sg13g2_antennanp ANTENNA_705 (.A(net124));
 sg13g2_antennanp ANTENNA_706 (.A(net124));
 sg13g2_antennanp ANTENNA_707 (.A(net124));
 sg13g2_antennanp ANTENNA_708 (.A(net124));
 sg13g2_antennanp ANTENNA_709 (.A(net124));
 sg13g2_antennanp ANTENNA_710 (.A(net124));
 sg13g2_antennanp ANTENNA_711 (.A(net155));
 sg13g2_antennanp ANTENNA_712 (.A(net155));
 sg13g2_antennanp ANTENNA_713 (.A(net155));
 sg13g2_antennanp ANTENNA_714 (.A(net155));
 sg13g2_antennanp ANTENNA_715 (.A(net155));
 sg13g2_antennanp ANTENNA_716 (.A(net155));
 sg13g2_antennanp ANTENNA_717 (.A(net155));
 sg13g2_antennanp ANTENNA_718 (.A(net155));
 sg13g2_antennanp ANTENNA_719 (.A(net155));
 sg13g2_antennanp ANTENNA_720 (.A(net155));
 sg13g2_antennanp ANTENNA_721 (.A(net155));
 sg13g2_antennanp ANTENNA_722 (.A(_00631_));
 sg13g2_antennanp ANTENNA_723 (.A(_01231_));
 sg13g2_antennanp ANTENNA_724 (.A(_01231_));
 sg13g2_antennanp ANTENNA_725 (.A(_01231_));
 sg13g2_antennanp ANTENNA_726 (.A(_01231_));
 sg13g2_antennanp ANTENNA_727 (.A(_01653_));
 sg13g2_antennanp ANTENNA_728 (.A(_01653_));
 sg13g2_antennanp ANTENNA_729 (.A(_01653_));
 sg13g2_antennanp ANTENNA_730 (.A(_01653_));
 sg13g2_antennanp ANTENNA_731 (.A(_01653_));
 sg13g2_antennanp ANTENNA_732 (.A(_01653_));
 sg13g2_antennanp ANTENNA_733 (.A(_01653_));
 sg13g2_antennanp ANTENNA_734 (.A(_01653_));
 sg13g2_antennanp ANTENNA_735 (.A(_02012_));
 sg13g2_antennanp ANTENNA_736 (.A(_02012_));
 sg13g2_antennanp ANTENNA_737 (.A(_02012_));
 sg13g2_antennanp ANTENNA_738 (.A(_02012_));
 sg13g2_antennanp ANTENNA_739 (.A(_02067_));
 sg13g2_antennanp ANTENNA_740 (.A(_02067_));
 sg13g2_antennanp ANTENNA_741 (.A(_02067_));
 sg13g2_antennanp ANTENNA_742 (.A(_02067_));
 sg13g2_antennanp ANTENNA_743 (.A(_02067_));
 sg13g2_antennanp ANTENNA_744 (.A(_02078_));
 sg13g2_antennanp ANTENNA_745 (.A(_02078_));
 sg13g2_antennanp ANTENNA_746 (.A(_02078_));
 sg13g2_antennanp ANTENNA_747 (.A(_02078_));
 sg13g2_antennanp ANTENNA_748 (.A(_02078_));
 sg13g2_antennanp ANTENNA_749 (.A(_02078_));
 sg13g2_antennanp ANTENNA_750 (.A(_02078_));
 sg13g2_antennanp ANTENNA_751 (.A(_02078_));
 sg13g2_antennanp ANTENNA_752 (.A(_02242_));
 sg13g2_antennanp ANTENNA_753 (.A(_02242_));
 sg13g2_antennanp ANTENNA_754 (.A(_02296_));
 sg13g2_antennanp ANTENNA_755 (.A(_02296_));
 sg13g2_antennanp ANTENNA_756 (.A(_02296_));
 sg13g2_antennanp ANTENNA_757 (.A(_02350_));
 sg13g2_antennanp ANTENNA_758 (.A(_02350_));
 sg13g2_antennanp ANTENNA_759 (.A(_02350_));
 sg13g2_antennanp ANTENNA_760 (.A(_02350_));
 sg13g2_antennanp ANTENNA_761 (.A(_02807_));
 sg13g2_antennanp ANTENNA_762 (.A(_02807_));
 sg13g2_antennanp ANTENNA_763 (.A(_02899_));
 sg13g2_antennanp ANTENNA_764 (.A(_02899_));
 sg13g2_antennanp ANTENNA_765 (.A(_02902_));
 sg13g2_antennanp ANTENNA_766 (.A(_02902_));
 sg13g2_antennanp ANTENNA_767 (.A(_02906_));
 sg13g2_antennanp ANTENNA_768 (.A(_02914_));
 sg13g2_antennanp ANTENNA_769 (.A(_02919_));
 sg13g2_antennanp ANTENNA_770 (.A(_02921_));
 sg13g2_antennanp ANTENNA_771 (.A(_02948_));
 sg13g2_antennanp ANTENNA_772 (.A(_02953_));
 sg13g2_antennanp ANTENNA_773 (.A(_02954_));
 sg13g2_antennanp ANTENNA_774 (.A(_02957_));
 sg13g2_antennanp ANTENNA_775 (.A(_02959_));
 sg13g2_antennanp ANTENNA_776 (.A(_02975_));
 sg13g2_antennanp ANTENNA_777 (.A(_02988_));
 sg13g2_antennanp ANTENNA_778 (.A(_02989_));
 sg13g2_antennanp ANTENNA_779 (.A(_02992_));
 sg13g2_antennanp ANTENNA_780 (.A(_02993_));
 sg13g2_antennanp ANTENNA_781 (.A(_03064_));
 sg13g2_antennanp ANTENNA_782 (.A(_03064_));
 sg13g2_antennanp ANTENNA_783 (.A(_03064_));
 sg13g2_antennanp ANTENNA_784 (.A(_03064_));
 sg13g2_antennanp ANTENNA_785 (.A(_03071_));
 sg13g2_antennanp ANTENNA_786 (.A(_03071_));
 sg13g2_antennanp ANTENNA_787 (.A(_03071_));
 sg13g2_antennanp ANTENNA_788 (.A(_03071_));
 sg13g2_antennanp ANTENNA_789 (.A(_03071_));
 sg13g2_antennanp ANTENNA_790 (.A(_03071_));
 sg13g2_antennanp ANTENNA_791 (.A(_03074_));
 sg13g2_antennanp ANTENNA_792 (.A(_03074_));
 sg13g2_antennanp ANTENNA_793 (.A(_03082_));
 sg13g2_antennanp ANTENNA_794 (.A(_03082_));
 sg13g2_antennanp ANTENNA_795 (.A(_03082_));
 sg13g2_antennanp ANTENNA_796 (.A(_03083_));
 sg13g2_antennanp ANTENNA_797 (.A(_03083_));
 sg13g2_antennanp ANTENNA_798 (.A(_03083_));
 sg13g2_antennanp ANTENNA_799 (.A(_03083_));
 sg13g2_antennanp ANTENNA_800 (.A(_03083_));
 sg13g2_antennanp ANTENNA_801 (.A(_03083_));
 sg13g2_antennanp ANTENNA_802 (.A(_03083_));
 sg13g2_antennanp ANTENNA_803 (.A(_03083_));
 sg13g2_antennanp ANTENNA_804 (.A(_03083_));
 sg13g2_antennanp ANTENNA_805 (.A(_03083_));
 sg13g2_antennanp ANTENNA_806 (.A(_03086_));
 sg13g2_antennanp ANTENNA_807 (.A(_03086_));
 sg13g2_antennanp ANTENNA_808 (.A(_03086_));
 sg13g2_antennanp ANTENNA_809 (.A(_03089_));
 sg13g2_antennanp ANTENNA_810 (.A(_03089_));
 sg13g2_antennanp ANTENNA_811 (.A(_03089_));
 sg13g2_antennanp ANTENNA_812 (.A(_03089_));
 sg13g2_antennanp ANTENNA_813 (.A(_03089_));
 sg13g2_antennanp ANTENNA_814 (.A(_03089_));
 sg13g2_antennanp ANTENNA_815 (.A(_03089_));
 sg13g2_antennanp ANTENNA_816 (.A(_03089_));
 sg13g2_antennanp ANTENNA_817 (.A(_03096_));
 sg13g2_antennanp ANTENNA_818 (.A(_03096_));
 sg13g2_antennanp ANTENNA_819 (.A(_03096_));
 sg13g2_antennanp ANTENNA_820 (.A(_03104_));
 sg13g2_antennanp ANTENNA_821 (.A(_03104_));
 sg13g2_antennanp ANTENNA_822 (.A(_03104_));
 sg13g2_antennanp ANTENNA_823 (.A(_03166_));
 sg13g2_antennanp ANTENNA_824 (.A(_03166_));
 sg13g2_antennanp ANTENNA_825 (.A(_03166_));
 sg13g2_antennanp ANTENNA_826 (.A(_03166_));
 sg13g2_antennanp ANTENNA_827 (.A(_03166_));
 sg13g2_antennanp ANTENNA_828 (.A(_03166_));
 sg13g2_antennanp ANTENNA_829 (.A(_03166_));
 sg13g2_antennanp ANTENNA_830 (.A(_03166_));
 sg13g2_antennanp ANTENNA_831 (.A(_03166_));
 sg13g2_antennanp ANTENNA_832 (.A(_03318_));
 sg13g2_antennanp ANTENNA_833 (.A(_03318_));
 sg13g2_antennanp ANTENNA_834 (.A(_03318_));
 sg13g2_antennanp ANTENNA_835 (.A(_03592_));
 sg13g2_antennanp ANTENNA_836 (.A(_03592_));
 sg13g2_antennanp ANTENNA_837 (.A(_03592_));
 sg13g2_antennanp ANTENNA_838 (.A(_03592_));
 sg13g2_antennanp ANTENNA_839 (.A(_03592_));
 sg13g2_antennanp ANTENNA_840 (.A(_03592_));
 sg13g2_antennanp ANTENNA_841 (.A(_03592_));
 sg13g2_antennanp ANTENNA_842 (.A(_03592_));
 sg13g2_antennanp ANTENNA_843 (.A(_03592_));
 sg13g2_antennanp ANTENNA_844 (.A(_03592_));
 sg13g2_antennanp ANTENNA_845 (.A(_03592_));
 sg13g2_antennanp ANTENNA_846 (.A(_03592_));
 sg13g2_antennanp ANTENNA_847 (.A(_03592_));
 sg13g2_antennanp ANTENNA_848 (.A(_03592_));
 sg13g2_antennanp ANTENNA_849 (.A(_03592_));
 sg13g2_antennanp ANTENNA_850 (.A(_03592_));
 sg13g2_antennanp ANTENNA_851 (.A(_03644_));
 sg13g2_antennanp ANTENNA_852 (.A(_03644_));
 sg13g2_antennanp ANTENNA_853 (.A(_03644_));
 sg13g2_antennanp ANTENNA_854 (.A(_03663_));
 sg13g2_antennanp ANTENNA_855 (.A(_03663_));
 sg13g2_antennanp ANTENNA_856 (.A(_03663_));
 sg13g2_antennanp ANTENNA_857 (.A(_03695_));
 sg13g2_antennanp ANTENNA_858 (.A(_03695_));
 sg13g2_antennanp ANTENNA_859 (.A(_03695_));
 sg13g2_antennanp ANTENNA_860 (.A(_03695_));
 sg13g2_antennanp ANTENNA_861 (.A(_03695_));
 sg13g2_antennanp ANTENNA_862 (.A(_03695_));
 sg13g2_antennanp ANTENNA_863 (.A(_03954_));
 sg13g2_antennanp ANTENNA_864 (.A(_03954_));
 sg13g2_antennanp ANTENNA_865 (.A(_03954_));
 sg13g2_antennanp ANTENNA_866 (.A(_04048_));
 sg13g2_antennanp ANTENNA_867 (.A(_04048_));
 sg13g2_antennanp ANTENNA_868 (.A(_04048_));
 sg13g2_antennanp ANTENNA_869 (.A(_04048_));
 sg13g2_antennanp ANTENNA_870 (.A(_04064_));
 sg13g2_antennanp ANTENNA_871 (.A(_04064_));
 sg13g2_antennanp ANTENNA_872 (.A(_04064_));
 sg13g2_antennanp ANTENNA_873 (.A(_04064_));
 sg13g2_antennanp ANTENNA_874 (.A(_04243_));
 sg13g2_antennanp ANTENNA_875 (.A(_04243_));
 sg13g2_antennanp ANTENNA_876 (.A(_04243_));
 sg13g2_antennanp ANTENNA_877 (.A(_04243_));
 sg13g2_antennanp ANTENNA_878 (.A(_04263_));
 sg13g2_antennanp ANTENNA_879 (.A(_04263_));
 sg13g2_antennanp ANTENNA_880 (.A(_04263_));
 sg13g2_antennanp ANTENNA_881 (.A(_04287_));
 sg13g2_antennanp ANTENNA_882 (.A(_04287_));
 sg13g2_antennanp ANTENNA_883 (.A(_04287_));
 sg13g2_antennanp ANTENNA_884 (.A(_04348_));
 sg13g2_antennanp ANTENNA_885 (.A(_04348_));
 sg13g2_antennanp ANTENNA_886 (.A(_04348_));
 sg13g2_antennanp ANTENNA_887 (.A(_04348_));
 sg13g2_antennanp ANTENNA_888 (.A(_04485_));
 sg13g2_antennanp ANTENNA_889 (.A(_04485_));
 sg13g2_antennanp ANTENNA_890 (.A(_04485_));
 sg13g2_antennanp ANTENNA_891 (.A(_04485_));
 sg13g2_antennanp ANTENNA_892 (.A(_04485_));
 sg13g2_antennanp ANTENNA_893 (.A(_05084_));
 sg13g2_antennanp ANTENNA_894 (.A(_05084_));
 sg13g2_antennanp ANTENNA_895 (.A(_05084_));
 sg13g2_antennanp ANTENNA_896 (.A(_05084_));
 sg13g2_antennanp ANTENNA_897 (.A(_05084_));
 sg13g2_antennanp ANTENNA_898 (.A(_05090_));
 sg13g2_antennanp ANTENNA_899 (.A(_05090_));
 sg13g2_antennanp ANTENNA_900 (.A(_05090_));
 sg13g2_antennanp ANTENNA_901 (.A(_05090_));
 sg13g2_antennanp ANTENNA_902 (.A(_05111_));
 sg13g2_antennanp ANTENNA_903 (.A(_05111_));
 sg13g2_antennanp ANTENNA_904 (.A(_05111_));
 sg13g2_antennanp ANTENNA_905 (.A(_05111_));
 sg13g2_antennanp ANTENNA_906 (.A(_05828_));
 sg13g2_antennanp ANTENNA_907 (.A(_05828_));
 sg13g2_antennanp ANTENNA_908 (.A(_05828_));
 sg13g2_antennanp ANTENNA_909 (.A(_05828_));
 sg13g2_antennanp ANTENNA_910 (.A(_05828_));
 sg13g2_antennanp ANTENNA_911 (.A(_05828_));
 sg13g2_antennanp ANTENNA_912 (.A(_05828_));
 sg13g2_antennanp ANTENNA_913 (.A(_07381_));
 sg13g2_antennanp ANTENNA_914 (.A(_07381_));
 sg13g2_antennanp ANTENNA_915 (.A(_07381_));
 sg13g2_antennanp ANTENNA_916 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_917 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_918 (.A(clk));
 sg13g2_antennanp ANTENNA_919 (.A(clk));
 sg13g2_antennanp ANTENNA_920 (.A(net63));
 sg13g2_antennanp ANTENNA_921 (.A(net63));
 sg13g2_antennanp ANTENNA_922 (.A(net63));
 sg13g2_antennanp ANTENNA_923 (.A(net63));
 sg13g2_antennanp ANTENNA_924 (.A(net63));
 sg13g2_antennanp ANTENNA_925 (.A(net63));
 sg13g2_antennanp ANTENNA_926 (.A(net63));
 sg13g2_antennanp ANTENNA_927 (.A(net63));
 sg13g2_antennanp ANTENNA_928 (.A(net93));
 sg13g2_antennanp ANTENNA_929 (.A(net93));
 sg13g2_antennanp ANTENNA_930 (.A(net93));
 sg13g2_antennanp ANTENNA_931 (.A(net93));
 sg13g2_antennanp ANTENNA_932 (.A(net93));
 sg13g2_antennanp ANTENNA_933 (.A(net93));
 sg13g2_antennanp ANTENNA_934 (.A(net93));
 sg13g2_antennanp ANTENNA_935 (.A(net93));
 sg13g2_antennanp ANTENNA_936 (.A(net93));
 sg13g2_antennanp ANTENNA_937 (.A(net93));
 sg13g2_antennanp ANTENNA_938 (.A(net93));
 sg13g2_antennanp ANTENNA_939 (.A(net93));
 sg13g2_antennanp ANTENNA_940 (.A(net93));
 sg13g2_antennanp ANTENNA_941 (.A(net93));
 sg13g2_antennanp ANTENNA_942 (.A(net93));
 sg13g2_antennanp ANTENNA_943 (.A(net93));
 sg13g2_antennanp ANTENNA_944 (.A(net124));
 sg13g2_antennanp ANTENNA_945 (.A(net124));
 sg13g2_antennanp ANTENNA_946 (.A(net124));
 sg13g2_antennanp ANTENNA_947 (.A(net124));
 sg13g2_antennanp ANTENNA_948 (.A(net124));
 sg13g2_antennanp ANTENNA_949 (.A(net124));
 sg13g2_antennanp ANTENNA_950 (.A(net124));
 sg13g2_antennanp ANTENNA_951 (.A(net124));
 sg13g2_antennanp ANTENNA_952 (.A(net124));
 sg13g2_antennanp ANTENNA_953 (.A(net124));
 sg13g2_antennanp ANTENNA_954 (.A(net124));
 sg13g2_antennanp ANTENNA_955 (.A(net124));
 sg13g2_antennanp ANTENNA_956 (.A(net124));
 sg13g2_antennanp ANTENNA_957 (.A(net124));
 sg13g2_antennanp ANTENNA_958 (.A(net124));
 sg13g2_antennanp ANTENNA_959 (.A(net155));
 sg13g2_antennanp ANTENNA_960 (.A(net155));
 sg13g2_antennanp ANTENNA_961 (.A(net155));
 sg13g2_antennanp ANTENNA_962 (.A(net155));
 sg13g2_antennanp ANTENNA_963 (.A(net155));
 sg13g2_antennanp ANTENNA_964 (.A(net155));
 sg13g2_antennanp ANTENNA_965 (.A(net155));
 sg13g2_antennanp ANTENNA_966 (.A(net155));
 sg13g2_antennanp ANTENNA_967 (.A(net155));
 sg13g2_antennanp ANTENNA_968 (.A(net155));
 sg13g2_antennanp ANTENNA_969 (.A(net155));
 sg13g2_antennanp ANTENNA_970 (.A(net155));
 sg13g2_antennanp ANTENNA_971 (.A(net155));
 sg13g2_antennanp ANTENNA_972 (.A(net155));
 sg13g2_antennanp ANTENNA_973 (.A(net155));
 sg13g2_antennanp ANTENNA_974 (.A(net155));
 sg13g2_antennanp ANTENNA_975 (.A(net155));
 sg13g2_antennanp ANTENNA_976 (.A(net155));
 sg13g2_antennanp ANTENNA_977 (.A(net155));
 sg13g2_antennanp ANTENNA_978 (.A(net155));
 sg13g2_antennanp ANTENNA_979 (.A(net155));
 sg13g2_antennanp ANTENNA_980 (.A(net155));
 sg13g2_antennanp ANTENNA_981 (.A(net155));
 sg13g2_antennanp ANTENNA_982 (.A(net155));
 sg13g2_antennanp ANTENNA_983 (.A(_00631_));
 sg13g2_antennanp ANTENNA_984 (.A(_01231_));
 sg13g2_antennanp ANTENNA_985 (.A(_01231_));
 sg13g2_antennanp ANTENNA_986 (.A(_01231_));
 sg13g2_antennanp ANTENNA_987 (.A(_01231_));
 sg13g2_antennanp ANTENNA_988 (.A(_01231_));
 sg13g2_antennanp ANTENNA_989 (.A(_01231_));
 sg13g2_antennanp ANTENNA_990 (.A(_01231_));
 sg13g2_antennanp ANTENNA_991 (.A(_01231_));
 sg13g2_antennanp ANTENNA_992 (.A(_01231_));
 sg13g2_antennanp ANTENNA_993 (.A(_01231_));
 sg13g2_antennanp ANTENNA_994 (.A(_01653_));
 sg13g2_antennanp ANTENNA_995 (.A(_01653_));
 sg13g2_antennanp ANTENNA_996 (.A(_01653_));
 sg13g2_antennanp ANTENNA_997 (.A(_01653_));
 sg13g2_antennanp ANTENNA_998 (.A(_01653_));
 sg13g2_antennanp ANTENNA_999 (.A(_01653_));
 sg13g2_antennanp ANTENNA_1000 (.A(_01653_));
 sg13g2_antennanp ANTENNA_1001 (.A(_01653_));
 sg13g2_antennanp ANTENNA_1002 (.A(_02012_));
 sg13g2_antennanp ANTENNA_1003 (.A(_02012_));
 sg13g2_antennanp ANTENNA_1004 (.A(_02012_));
 sg13g2_antennanp ANTENNA_1005 (.A(_02012_));
 sg13g2_antennanp ANTENNA_1006 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1007 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1008 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1009 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1010 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1011 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1012 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1013 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1014 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1015 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1016 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1017 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1018 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1019 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1020 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1021 (.A(_02242_));
 sg13g2_antennanp ANTENNA_1022 (.A(_02242_));
 sg13g2_antennanp ANTENNA_1023 (.A(_02242_));
 sg13g2_antennanp ANTENNA_1024 (.A(_02242_));
 sg13g2_antennanp ANTENNA_1025 (.A(_02350_));
 sg13g2_antennanp ANTENNA_1026 (.A(_02350_));
 sg13g2_antennanp ANTENNA_1027 (.A(_02350_));
 sg13g2_antennanp ANTENNA_1028 (.A(_02350_));
 sg13g2_antennanp ANTENNA_1029 (.A(_02807_));
 sg13g2_antennanp ANTENNA_1030 (.A(_02807_));
 sg13g2_antennanp ANTENNA_1031 (.A(_02899_));
 sg13g2_antennanp ANTENNA_1032 (.A(_02899_));
 sg13g2_antennanp ANTENNA_1033 (.A(_02902_));
 sg13g2_antennanp ANTENNA_1034 (.A(_02906_));
 sg13g2_antennanp ANTENNA_1035 (.A(_02914_));
 sg13g2_antennanp ANTENNA_1036 (.A(_02919_));
 sg13g2_antennanp ANTENNA_1037 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1038 (.A(_02948_));
 sg13g2_antennanp ANTENNA_1039 (.A(_02953_));
 sg13g2_antennanp ANTENNA_1040 (.A(_02954_));
 sg13g2_antennanp ANTENNA_1041 (.A(_02957_));
 sg13g2_antennanp ANTENNA_1042 (.A(_02959_));
 sg13g2_antennanp ANTENNA_1043 (.A(_02975_));
 sg13g2_antennanp ANTENNA_1044 (.A(_02988_));
 sg13g2_antennanp ANTENNA_1045 (.A(_02989_));
 sg13g2_antennanp ANTENNA_1046 (.A(_02992_));
 sg13g2_antennanp ANTENNA_1047 (.A(_02993_));
 sg13g2_antennanp ANTENNA_1048 (.A(_03064_));
 sg13g2_antennanp ANTENNA_1049 (.A(_03064_));
 sg13g2_antennanp ANTENNA_1050 (.A(_03064_));
 sg13g2_antennanp ANTENNA_1051 (.A(_03064_));
 sg13g2_antennanp ANTENNA_1052 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1053 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1054 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1055 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1056 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1057 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1058 (.A(_03074_));
 sg13g2_antennanp ANTENNA_1059 (.A(_03074_));
 sg13g2_antennanp ANTENNA_1060 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1061 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1062 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1063 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1064 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1065 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1066 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1067 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1068 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1069 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1070 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1071 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1072 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1073 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1074 (.A(_03082_));
 sg13g2_antennanp ANTENNA_1075 (.A(_03082_));
 sg13g2_antennanp ANTENNA_1076 (.A(_03082_));
 sg13g2_antennanp ANTENNA_1077 (.A(_03083_));
 sg13g2_antennanp ANTENNA_1078 (.A(_03083_));
 sg13g2_antennanp ANTENNA_1079 (.A(_03083_));
 sg13g2_antennanp ANTENNA_1080 (.A(_03083_));
 sg13g2_antennanp ANTENNA_1081 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1082 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1083 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1084 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1085 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1086 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1087 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1088 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1089 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1090 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1091 (.A(_03089_));
 sg13g2_antennanp ANTENNA_1092 (.A(_03089_));
 sg13g2_antennanp ANTENNA_1093 (.A(_03089_));
 sg13g2_antennanp ANTENNA_1094 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1095 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1096 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1097 (.A(_03104_));
 sg13g2_antennanp ANTENNA_1098 (.A(_03104_));
 sg13g2_antennanp ANTENNA_1099 (.A(_03104_));
 sg13g2_antennanp ANTENNA_1100 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1101 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1102 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1103 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1104 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1105 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1106 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1107 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1108 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1109 (.A(_03318_));
 sg13g2_antennanp ANTENNA_1110 (.A(_03318_));
 sg13g2_antennanp ANTENNA_1111 (.A(_03318_));
 sg13g2_antennanp ANTENNA_1112 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1113 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1114 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1115 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1116 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1117 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1118 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1119 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1120 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1121 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1122 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1123 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1124 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1125 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1126 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1127 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1128 (.A(_03644_));
 sg13g2_antennanp ANTENNA_1129 (.A(_03644_));
 sg13g2_antennanp ANTENNA_1130 (.A(_03644_));
 sg13g2_antennanp ANTENNA_1131 (.A(_03663_));
 sg13g2_antennanp ANTENNA_1132 (.A(_03663_));
 sg13g2_antennanp ANTENNA_1133 (.A(_03663_));
 sg13g2_antennanp ANTENNA_1134 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1135 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1136 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1137 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1138 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1139 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1140 (.A(_03954_));
 sg13g2_antennanp ANTENNA_1141 (.A(_03954_));
 sg13g2_antennanp ANTENNA_1142 (.A(_03954_));
 sg13g2_antennanp ANTENNA_1143 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1144 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1145 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1146 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1147 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1148 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1149 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1150 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1151 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1152 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1153 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1154 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1155 (.A(_04048_));
 sg13g2_antennanp ANTENNA_1156 (.A(_04048_));
 sg13g2_antennanp ANTENNA_1157 (.A(_04048_));
 sg13g2_antennanp ANTENNA_1158 (.A(_04048_));
 sg13g2_antennanp ANTENNA_1159 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1160 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1161 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1162 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1163 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1164 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1165 (.A(_04243_));
 sg13g2_antennanp ANTENNA_1166 (.A(_04243_));
 sg13g2_antennanp ANTENNA_1167 (.A(_04243_));
 sg13g2_antennanp ANTENNA_1168 (.A(_04243_));
 sg13g2_antennanp ANTENNA_1169 (.A(_04263_));
 sg13g2_antennanp ANTENNA_1170 (.A(_04263_));
 sg13g2_antennanp ANTENNA_1171 (.A(_04263_));
 sg13g2_antennanp ANTENNA_1172 (.A(_04348_));
 sg13g2_antennanp ANTENNA_1173 (.A(_04348_));
 sg13g2_antennanp ANTENNA_1174 (.A(_04348_));
 sg13g2_antennanp ANTENNA_1175 (.A(_04348_));
 sg13g2_antennanp ANTENNA_1176 (.A(_04485_));
 sg13g2_antennanp ANTENNA_1177 (.A(_04485_));
 sg13g2_antennanp ANTENNA_1178 (.A(_04485_));
 sg13g2_antennanp ANTENNA_1179 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1180 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1181 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1182 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1183 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1184 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1185 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1186 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1187 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1188 (.A(_05111_));
 sg13g2_antennanp ANTENNA_1189 (.A(_05111_));
 sg13g2_antennanp ANTENNA_1190 (.A(_05111_));
 sg13g2_antennanp ANTENNA_1191 (.A(_05111_));
 sg13g2_antennanp ANTENNA_1192 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1193 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1194 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1195 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1196 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1197 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1198 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1199 (.A(_07381_));
 sg13g2_antennanp ANTENNA_1200 (.A(_07381_));
 sg13g2_antennanp ANTENNA_1201 (.A(_07381_));
 sg13g2_antennanp ANTENNA_1202 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_1203 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_1204 (.A(clk));
 sg13g2_antennanp ANTENNA_1205 (.A(clk));
 sg13g2_antennanp ANTENNA_1206 (.A(net93));
 sg13g2_antennanp ANTENNA_1207 (.A(net93));
 sg13g2_antennanp ANTENNA_1208 (.A(net93));
 sg13g2_antennanp ANTENNA_1209 (.A(net93));
 sg13g2_antennanp ANTENNA_1210 (.A(net93));
 sg13g2_antennanp ANTENNA_1211 (.A(net93));
 sg13g2_antennanp ANTENNA_1212 (.A(net93));
 sg13g2_antennanp ANTENNA_1213 (.A(net93));
 sg13g2_antennanp ANTENNA_1214 (.A(net93));
 sg13g2_antennanp ANTENNA_1215 (.A(net93));
 sg13g2_antennanp ANTENNA_1216 (.A(net93));
 sg13g2_antennanp ANTENNA_1217 (.A(net109));
 sg13g2_antennanp ANTENNA_1218 (.A(net109));
 sg13g2_antennanp ANTENNA_1219 (.A(net109));
 sg13g2_antennanp ANTENNA_1220 (.A(net109));
 sg13g2_antennanp ANTENNA_1221 (.A(net109));
 sg13g2_antennanp ANTENNA_1222 (.A(net109));
 sg13g2_antennanp ANTENNA_1223 (.A(net109));
 sg13g2_antennanp ANTENNA_1224 (.A(net109));
 sg13g2_antennanp ANTENNA_1225 (.A(net109));
 sg13g2_antennanp ANTENNA_1226 (.A(net124));
 sg13g2_antennanp ANTENNA_1227 (.A(net124));
 sg13g2_antennanp ANTENNA_1228 (.A(net124));
 sg13g2_antennanp ANTENNA_1229 (.A(net124));
 sg13g2_antennanp ANTENNA_1230 (.A(net124));
 sg13g2_antennanp ANTENNA_1231 (.A(net124));
 sg13g2_antennanp ANTENNA_1232 (.A(net124));
 sg13g2_antennanp ANTENNA_1233 (.A(net124));
 sg13g2_antennanp ANTENNA_1234 (.A(net124));
 sg13g2_antennanp ANTENNA_1235 (.A(_00631_));
 sg13g2_antennanp ANTENNA_1236 (.A(_01231_));
 sg13g2_antennanp ANTENNA_1237 (.A(_01231_));
 sg13g2_antennanp ANTENNA_1238 (.A(_01231_));
 sg13g2_antennanp ANTENNA_1239 (.A(_01231_));
 sg13g2_antennanp ANTENNA_1240 (.A(_02012_));
 sg13g2_antennanp ANTENNA_1241 (.A(_02012_));
 sg13g2_antennanp ANTENNA_1242 (.A(_02012_));
 sg13g2_antennanp ANTENNA_1243 (.A(_02012_));
 sg13g2_antennanp ANTENNA_1244 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1245 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1246 (.A(_02067_));
 sg13g2_antennanp ANTENNA_1247 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1248 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1249 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1250 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1251 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1252 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1253 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1254 (.A(_02078_));
 sg13g2_antennanp ANTENNA_1255 (.A(_02242_));
 sg13g2_antennanp ANTENNA_1256 (.A(_02242_));
 sg13g2_antennanp ANTENNA_1257 (.A(_02242_));
 sg13g2_antennanp ANTENNA_1258 (.A(_02242_));
 sg13g2_antennanp ANTENNA_1259 (.A(_02807_));
 sg13g2_antennanp ANTENNA_1260 (.A(_02899_));
 sg13g2_antennanp ANTENNA_1261 (.A(_02899_));
 sg13g2_antennanp ANTENNA_1262 (.A(_02902_));
 sg13g2_antennanp ANTENNA_1263 (.A(_02902_));
 sg13g2_antennanp ANTENNA_1264 (.A(_02906_));
 sg13g2_antennanp ANTENNA_1265 (.A(_02914_));
 sg13g2_antennanp ANTENNA_1266 (.A(_02919_));
 sg13g2_antennanp ANTENNA_1267 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1268 (.A(_02948_));
 sg13g2_antennanp ANTENNA_1269 (.A(_02953_));
 sg13g2_antennanp ANTENNA_1270 (.A(_02954_));
 sg13g2_antennanp ANTENNA_1271 (.A(_02957_));
 sg13g2_antennanp ANTENNA_1272 (.A(_02959_));
 sg13g2_antennanp ANTENNA_1273 (.A(_02975_));
 sg13g2_antennanp ANTENNA_1274 (.A(_02988_));
 sg13g2_antennanp ANTENNA_1275 (.A(_02989_));
 sg13g2_antennanp ANTENNA_1276 (.A(_02992_));
 sg13g2_antennanp ANTENNA_1277 (.A(_02993_));
 sg13g2_antennanp ANTENNA_1278 (.A(_03064_));
 sg13g2_antennanp ANTENNA_1279 (.A(_03064_));
 sg13g2_antennanp ANTENNA_1280 (.A(_03064_));
 sg13g2_antennanp ANTENNA_1281 (.A(_03064_));
 sg13g2_antennanp ANTENNA_1282 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1283 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1284 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1285 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1286 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1287 (.A(_03071_));
 sg13g2_antennanp ANTENNA_1288 (.A(_03074_));
 sg13g2_antennanp ANTENNA_1289 (.A(_03074_));
 sg13g2_antennanp ANTENNA_1290 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1291 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1292 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1293 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1294 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1295 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1296 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1297 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1298 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1299 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1300 (.A(_03082_));
 sg13g2_antennanp ANTENNA_1301 (.A(_03082_));
 sg13g2_antennanp ANTENNA_1302 (.A(_03082_));
 sg13g2_antennanp ANTENNA_1303 (.A(_03083_));
 sg13g2_antennanp ANTENNA_1304 (.A(_03083_));
 sg13g2_antennanp ANTENNA_1305 (.A(_03083_));
 sg13g2_antennanp ANTENNA_1306 (.A(_03083_));
 sg13g2_antennanp ANTENNA_1307 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1308 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1309 (.A(_03086_));
 sg13g2_antennanp ANTENNA_1310 (.A(_03089_));
 sg13g2_antennanp ANTENNA_1311 (.A(_03089_));
 sg13g2_antennanp ANTENNA_1312 (.A(_03089_));
 sg13g2_antennanp ANTENNA_1313 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1314 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1315 (.A(_03096_));
 sg13g2_antennanp ANTENNA_1316 (.A(_03104_));
 sg13g2_antennanp ANTENNA_1317 (.A(_03104_));
 sg13g2_antennanp ANTENNA_1318 (.A(_03104_));
 sg13g2_antennanp ANTENNA_1319 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1320 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1321 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1322 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1323 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1324 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1325 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1326 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1327 (.A(_03166_));
 sg13g2_antennanp ANTENNA_1328 (.A(_03318_));
 sg13g2_antennanp ANTENNA_1329 (.A(_03318_));
 sg13g2_antennanp ANTENNA_1330 (.A(_03318_));
 sg13g2_antennanp ANTENNA_1331 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1332 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1333 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1334 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1335 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1336 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1337 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1338 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1339 (.A(_03592_));
 sg13g2_antennanp ANTENNA_1340 (.A(_03644_));
 sg13g2_antennanp ANTENNA_1341 (.A(_03644_));
 sg13g2_antennanp ANTENNA_1342 (.A(_03644_));
 sg13g2_antennanp ANTENNA_1343 (.A(_03663_));
 sg13g2_antennanp ANTENNA_1344 (.A(_03663_));
 sg13g2_antennanp ANTENNA_1345 (.A(_03663_));
 sg13g2_antennanp ANTENNA_1346 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1347 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1348 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1349 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1350 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1351 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1352 (.A(_03954_));
 sg13g2_antennanp ANTENNA_1353 (.A(_03954_));
 sg13g2_antennanp ANTENNA_1354 (.A(_03954_));
 sg13g2_antennanp ANTENNA_1355 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1356 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1357 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1358 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1359 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1360 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1361 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1362 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1363 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1364 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1365 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1366 (.A(_04044_));
 sg13g2_antennanp ANTENNA_1367 (.A(_04048_));
 sg13g2_antennanp ANTENNA_1368 (.A(_04048_));
 sg13g2_antennanp ANTENNA_1369 (.A(_04048_));
 sg13g2_antennanp ANTENNA_1370 (.A(_04048_));
 sg13g2_antennanp ANTENNA_1371 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1372 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1373 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1374 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1375 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1376 (.A(_04064_));
 sg13g2_antennanp ANTENNA_1377 (.A(_04243_));
 sg13g2_antennanp ANTENNA_1378 (.A(_04243_));
 sg13g2_antennanp ANTENNA_1379 (.A(_04243_));
 sg13g2_antennanp ANTENNA_1380 (.A(_04243_));
 sg13g2_antennanp ANTENNA_1381 (.A(_04263_));
 sg13g2_antennanp ANTENNA_1382 (.A(_04263_));
 sg13g2_antennanp ANTENNA_1383 (.A(_04263_));
 sg13g2_antennanp ANTENNA_1384 (.A(_04348_));
 sg13g2_antennanp ANTENNA_1385 (.A(_04348_));
 sg13g2_antennanp ANTENNA_1386 (.A(_04348_));
 sg13g2_antennanp ANTENNA_1387 (.A(_04348_));
 sg13g2_antennanp ANTENNA_1388 (.A(_04485_));
 sg13g2_antennanp ANTENNA_1389 (.A(_04485_));
 sg13g2_antennanp ANTENNA_1390 (.A(_04485_));
 sg13g2_antennanp ANTENNA_1391 (.A(_04485_));
 sg13g2_antennanp ANTENNA_1392 (.A(_04485_));
 sg13g2_antennanp ANTENNA_1393 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1394 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1395 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1396 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1397 (.A(_05084_));
 sg13g2_antennanp ANTENNA_1398 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1399 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1400 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1401 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1402 (.A(_05111_));
 sg13g2_antennanp ANTENNA_1403 (.A(_05111_));
 sg13g2_antennanp ANTENNA_1404 (.A(_05111_));
 sg13g2_antennanp ANTENNA_1405 (.A(_05111_));
 sg13g2_antennanp ANTENNA_1406 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1407 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1408 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1409 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1410 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1411 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1412 (.A(_05828_));
 sg13g2_antennanp ANTENNA_1413 (.A(_08420_));
 sg13g2_antennanp ANTENNA_1414 (.A(_08420_));
 sg13g2_antennanp ANTENNA_1415 (.A(_08420_));
 sg13g2_antennanp ANTENNA_1416 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_1417 (.A(\b.gen_square[5].sq.piece[0] ));
 sg13g2_antennanp ANTENNA_1418 (.A(clk));
 sg13g2_antennanp ANTENNA_1419 (.A(clk));
 sg13g2_antennanp ANTENNA_1420 (.A(net86));
 sg13g2_antennanp ANTENNA_1421 (.A(net86));
 sg13g2_antennanp ANTENNA_1422 (.A(net86));
 sg13g2_antennanp ANTENNA_1423 (.A(net86));
 sg13g2_antennanp ANTENNA_1424 (.A(net86));
 sg13g2_antennanp ANTENNA_1425 (.A(net86));
 sg13g2_antennanp ANTENNA_1426 (.A(net86));
 sg13g2_antennanp ANTENNA_1427 (.A(net86));
 sg13g2_antennanp ANTENNA_1428 (.A(net86));
 sg13g2_antennanp ANTENNA_1429 (.A(net86));
 sg13g2_antennanp ANTENNA_1430 (.A(net86));
 sg13g2_antennanp ANTENNA_1431 (.A(net86));
 sg13g2_antennanp ANTENNA_1432 (.A(net86));
 sg13g2_antennanp ANTENNA_1433 (.A(net86));
 sg13g2_antennanp ANTENNA_1434 (.A(net93));
 sg13g2_antennanp ANTENNA_1435 (.A(net93));
 sg13g2_antennanp ANTENNA_1436 (.A(net93));
 sg13g2_antennanp ANTENNA_1437 (.A(net93));
 sg13g2_antennanp ANTENNA_1438 (.A(net93));
 sg13g2_antennanp ANTENNA_1439 (.A(net93));
 sg13g2_antennanp ANTENNA_1440 (.A(net93));
 sg13g2_antennanp ANTENNA_1441 (.A(net93));
 sg13g2_antennanp ANTENNA_1442 (.A(net109));
 sg13g2_antennanp ANTENNA_1443 (.A(net109));
 sg13g2_antennanp ANTENNA_1444 (.A(net109));
 sg13g2_antennanp ANTENNA_1445 (.A(net109));
 sg13g2_antennanp ANTENNA_1446 (.A(net109));
 sg13g2_antennanp ANTENNA_1447 (.A(net109));
 sg13g2_antennanp ANTENNA_1448 (.A(net109));
 sg13g2_antennanp ANTENNA_1449 (.A(net109));
 sg13g2_antennanp ANTENNA_1450 (.A(net109));
 sg13g2_antennanp ANTENNA_1451 (.A(net124));
 sg13g2_antennanp ANTENNA_1452 (.A(net124));
 sg13g2_antennanp ANTENNA_1453 (.A(net124));
 sg13g2_antennanp ANTENNA_1454 (.A(net124));
 sg13g2_antennanp ANTENNA_1455 (.A(net124));
 sg13g2_antennanp ANTENNA_1456 (.A(net124));
 sg13g2_antennanp ANTENNA_1457 (.A(net124));
 sg13g2_antennanp ANTENNA_1458 (.A(net124));
 sg13g2_antennanp ANTENNA_1459 (.A(net124));
 sg13g2_antennanp ANTENNA_1460 (.A(net155));
 sg13g2_antennanp ANTENNA_1461 (.A(net155));
 sg13g2_antennanp ANTENNA_1462 (.A(net155));
 sg13g2_antennanp ANTENNA_1463 (.A(net155));
 sg13g2_antennanp ANTENNA_1464 (.A(net155));
 sg13g2_antennanp ANTENNA_1465 (.A(net155));
 sg13g2_antennanp ANTENNA_1466 (.A(net155));
 sg13g2_antennanp ANTENNA_1467 (.A(net155));
 sg13g2_antennanp ANTENNA_1468 (.A(net155));
 sg13g2_antennanp ANTENNA_1469 (.A(net155));
 sg13g2_antennanp ANTENNA_1470 (.A(net155));
 sg13g2_antennanp ANTENNA_1471 (.A(net155));
 sg13g2_antennanp ANTENNA_1472 (.A(net155));
 sg13g2_antennanp ANTENNA_1473 (.A(net155));
 sg13g2_antennanp ANTENNA_1474 (.A(net155));
 sg13g2_antennanp ANTENNA_1475 (.A(net155));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_fill_1 FILLER_0_56 ();
 sg13g2_decap_4 FILLER_0_62 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_fill_2 FILLER_0_91 ();
 sg13g2_fill_1 FILLER_0_93 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_4 FILLER_0_117 ();
 sg13g2_fill_1 FILLER_0_121 ();
 sg13g2_decap_4 FILLER_0_127 ();
 sg13g2_fill_1 FILLER_0_131 ();
 sg13g2_decap_4 FILLER_0_137 ();
 sg13g2_fill_2 FILLER_0_141 ();
 sg13g2_decap_4 FILLER_0_148 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_4 FILLER_0_186 ();
 sg13g2_fill_1 FILLER_0_238 ();
 sg13g2_fill_2 FILLER_0_267 ();
 sg13g2_fill_1 FILLER_0_269 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_311 ();
 sg13g2_decap_4 FILLER_0_318 ();
 sg13g2_fill_1 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_decap_8 FILLER_0_422 ();
 sg13g2_fill_2 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_0_435 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_decap_8 FILLER_0_459 ();
 sg13g2_fill_1 FILLER_0_466 ();
 sg13g2_decap_8 FILLER_0_472 ();
 sg13g2_decap_8 FILLER_0_487 ();
 sg13g2_decap_8 FILLER_0_494 ();
 sg13g2_decap_4 FILLER_0_501 ();
 sg13g2_fill_1 FILLER_0_505 ();
 sg13g2_decap_8 FILLER_0_510 ();
 sg13g2_fill_2 FILLER_0_517 ();
 sg13g2_fill_1 FILLER_0_549 ();
 sg13g2_decap_4 FILLER_0_555 ();
 sg13g2_decap_4 FILLER_0_564 ();
 sg13g2_fill_1 FILLER_0_572 ();
 sg13g2_decap_8 FILLER_0_578 ();
 sg13g2_decap_8 FILLER_0_585 ();
 sg13g2_fill_1 FILLER_0_592 ();
 sg13g2_decap_8 FILLER_0_597 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_620 ();
 sg13g2_decap_8 FILLER_0_627 ();
 sg13g2_decap_8 FILLER_0_634 ();
 sg13g2_decap_8 FILLER_0_641 ();
 sg13g2_fill_2 FILLER_0_648 ();
 sg13g2_fill_1 FILLER_0_650 ();
 sg13g2_decap_8 FILLER_0_661 ();
 sg13g2_decap_4 FILLER_0_668 ();
 sg13g2_decap_4 FILLER_0_677 ();
 sg13g2_fill_1 FILLER_0_681 ();
 sg13g2_decap_4 FILLER_0_687 ();
 sg13g2_decap_8 FILLER_0_695 ();
 sg13g2_decap_8 FILLER_0_702 ();
 sg13g2_decap_4 FILLER_0_709 ();
 sg13g2_fill_1 FILLER_0_713 ();
 sg13g2_decap_8 FILLER_0_719 ();
 sg13g2_fill_2 FILLER_0_730 ();
 sg13g2_fill_2 FILLER_0_736 ();
 sg13g2_fill_1 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_774 ();
 sg13g2_fill_1 FILLER_0_781 ();
 sg13g2_decap_4 FILLER_0_791 ();
 sg13g2_fill_2 FILLER_0_795 ();
 sg13g2_fill_1 FILLER_0_801 ();
 sg13g2_decap_8 FILLER_0_807 ();
 sg13g2_decap_4 FILLER_0_814 ();
 sg13g2_fill_1 FILLER_0_818 ();
 sg13g2_decap_8 FILLER_0_823 ();
 sg13g2_decap_8 FILLER_0_830 ();
 sg13g2_decap_4 FILLER_0_837 ();
 sg13g2_fill_2 FILLER_0_841 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_4 FILLER_0_864 ();
 sg13g2_fill_2 FILLER_0_868 ();
 sg13g2_fill_2 FILLER_0_875 ();
 sg13g2_fill_1 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_4 FILLER_0_901 ();
 sg13g2_fill_2 FILLER_0_909 ();
 sg13g2_decap_4 FILLER_0_916 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_fill_1 FILLER_0_931 ();
 sg13g2_decap_4 FILLER_0_958 ();
 sg13g2_decap_8 FILLER_0_988 ();
 sg13g2_decap_8 FILLER_0_995 ();
 sg13g2_decap_8 FILLER_0_1002 ();
 sg13g2_decap_8 FILLER_0_1021 ();
 sg13g2_decap_4 FILLER_0_1028 ();
 sg13g2_fill_2 FILLER_0_1032 ();
 sg13g2_decap_4 FILLER_0_1039 ();
 sg13g2_fill_1 FILLER_0_1043 ();
 sg13g2_fill_2 FILLER_0_1048 ();
 sg13g2_fill_1 FILLER_0_1058 ();
 sg13g2_decap_8 FILLER_0_1064 ();
 sg13g2_decap_8 FILLER_0_1071 ();
 sg13g2_fill_2 FILLER_0_1082 ();
 sg13g2_decap_8 FILLER_0_1089 ();
 sg13g2_decap_8 FILLER_0_1096 ();
 sg13g2_decap_8 FILLER_0_1103 ();
 sg13g2_fill_1 FILLER_0_1140 ();
 sg13g2_decap_4 FILLER_0_1146 ();
 sg13g2_decap_8 FILLER_0_1159 ();
 sg13g2_fill_1 FILLER_0_1166 ();
 sg13g2_decap_8 FILLER_0_1172 ();
 sg13g2_decap_4 FILLER_0_1179 ();
 sg13g2_fill_1 FILLER_0_1183 ();
 sg13g2_fill_1 FILLER_0_1228 ();
 sg13g2_decap_8 FILLER_0_1238 ();
 sg13g2_decap_4 FILLER_0_1245 ();
 sg13g2_decap_4 FILLER_0_1254 ();
 sg13g2_decap_8 FILLER_0_1262 ();
 sg13g2_decap_8 FILLER_0_1269 ();
 sg13g2_decap_8 FILLER_0_1276 ();
 sg13g2_decap_8 FILLER_0_1283 ();
 sg13g2_decap_8 FILLER_0_1290 ();
 sg13g2_decap_8 FILLER_0_1297 ();
 sg13g2_decap_8 FILLER_0_1304 ();
 sg13g2_decap_8 FILLER_0_1311 ();
 sg13g2_decap_8 FILLER_0_1318 ();
 sg13g2_fill_1 FILLER_0_1325 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_4 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_46 ();
 sg13g2_fill_2 FILLER_1_73 ();
 sg13g2_fill_1 FILLER_1_75 ();
 sg13g2_fill_1 FILLER_1_128 ();
 sg13g2_fill_2 FILLER_1_155 ();
 sg13g2_fill_2 FILLER_1_183 ();
 sg13g2_fill_1 FILLER_1_185 ();
 sg13g2_fill_2 FILLER_1_191 ();
 sg13g2_fill_1 FILLER_1_193 ();
 sg13g2_fill_2 FILLER_1_248 ();
 sg13g2_decap_8 FILLER_1_299 ();
 sg13g2_decap_8 FILLER_1_306 ();
 sg13g2_decap_8 FILLER_1_313 ();
 sg13g2_decap_8 FILLER_1_320 ();
 sg13g2_decap_8 FILLER_1_327 ();
 sg13g2_fill_2 FILLER_1_334 ();
 sg13g2_fill_1 FILLER_1_336 ();
 sg13g2_fill_1 FILLER_1_342 ();
 sg13g2_fill_1 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_fill_1 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_fill_1 FILLER_1_398 ();
 sg13g2_decap_8 FILLER_1_521 ();
 sg13g2_decap_8 FILLER_1_528 ();
 sg13g2_fill_2 FILLER_1_535 ();
 sg13g2_decap_4 FILLER_1_541 ();
 sg13g2_fill_2 FILLER_1_545 ();
 sg13g2_fill_1 FILLER_1_599 ();
 sg13g2_decap_8 FILLER_1_734 ();
 sg13g2_fill_1 FILLER_1_741 ();
 sg13g2_fill_1 FILLER_1_768 ();
 sg13g2_fill_2 FILLER_1_774 ();
 sg13g2_fill_1 FILLER_1_802 ();
 sg13g2_fill_1 FILLER_1_829 ();
 sg13g2_fill_2 FILLER_1_943 ();
 sg13g2_decap_8 FILLER_1_949 ();
 sg13g2_decap_8 FILLER_1_956 ();
 sg13g2_decap_8 FILLER_1_963 ();
 sg13g2_decap_4 FILLER_1_970 ();
 sg13g2_decap_8 FILLER_1_983 ();
 sg13g2_decap_4 FILLER_1_990 ();
 sg13g2_fill_2 FILLER_1_994 ();
 sg13g2_decap_4 FILLER_1_1001 ();
 sg13g2_fill_2 FILLER_1_1005 ();
 sg13g2_fill_2 FILLER_1_1015 ();
 sg13g2_fill_1 FILLER_1_1020 ();
 sg13g2_fill_1 FILLER_1_1024 ();
 sg13g2_decap_4 FILLER_1_1029 ();
 sg13g2_fill_1 FILLER_1_1033 ();
 sg13g2_fill_1 FILLER_1_1060 ();
 sg13g2_fill_1 FILLER_1_1087 ();
 sg13g2_fill_2 FILLER_1_1114 ();
 sg13g2_decap_8 FILLER_1_1146 ();
 sg13g2_decap_8 FILLER_1_1153 ();
 sg13g2_decap_8 FILLER_1_1160 ();
 sg13g2_fill_2 FILLER_1_1167 ();
 sg13g2_decap_8 FILLER_1_1195 ();
 sg13g2_decap_4 FILLER_1_1206 ();
 sg13g2_decap_8 FILLER_1_1274 ();
 sg13g2_decap_8 FILLER_1_1281 ();
 sg13g2_decap_8 FILLER_1_1288 ();
 sg13g2_decap_8 FILLER_1_1295 ();
 sg13g2_decap_8 FILLER_1_1302 ();
 sg13g2_decap_8 FILLER_1_1309 ();
 sg13g2_decap_8 FILLER_1_1316 ();
 sg13g2_fill_2 FILLER_1_1323 ();
 sg13g2_fill_1 FILLER_1_1325 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_fill_2 FILLER_2_53 ();
 sg13g2_fill_1 FILLER_2_94 ();
 sg13g2_decap_8 FILLER_2_100 ();
 sg13g2_decap_8 FILLER_2_107 ();
 sg13g2_decap_8 FILLER_2_114 ();
 sg13g2_fill_2 FILLER_2_121 ();
 sg13g2_fill_1 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_128 ();
 sg13g2_decap_4 FILLER_2_135 ();
 sg13g2_fill_1 FILLER_2_139 ();
 sg13g2_decap_8 FILLER_2_148 ();
 sg13g2_decap_8 FILLER_2_155 ();
 sg13g2_decap_8 FILLER_2_162 ();
 sg13g2_decap_4 FILLER_2_169 ();
 sg13g2_decap_4 FILLER_2_176 ();
 sg13g2_fill_1 FILLER_2_183 ();
 sg13g2_fill_1 FILLER_2_205 ();
 sg13g2_fill_1 FILLER_2_237 ();
 sg13g2_fill_1 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_4 FILLER_2_270 ();
 sg13g2_fill_1 FILLER_2_274 ();
 sg13g2_decap_4 FILLER_2_278 ();
 sg13g2_decap_4 FILLER_2_296 ();
 sg13g2_fill_2 FILLER_2_300 ();
 sg13g2_fill_1 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_4 FILLER_2_336 ();
 sg13g2_fill_2 FILLER_2_340 ();
 sg13g2_decap_4 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_355 ();
 sg13g2_decap_8 FILLER_2_362 ();
 sg13g2_fill_2 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_2 FILLER_2_429 ();
 sg13g2_fill_2 FILLER_2_436 ();
 sg13g2_decap_8 FILLER_2_443 ();
 sg13g2_fill_2 FILLER_2_450 ();
 sg13g2_decap_8 FILLER_2_460 ();
 sg13g2_decap_4 FILLER_2_467 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_fill_1 FILLER_2_496 ();
 sg13g2_decap_4 FILLER_2_505 ();
 sg13g2_fill_2 FILLER_2_509 ();
 sg13g2_decap_4 FILLER_2_537 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_fill_2 FILLER_2_564 ();
 sg13g2_fill_1 FILLER_2_566 ();
 sg13g2_fill_2 FILLER_2_571 ();
 sg13g2_fill_1 FILLER_2_573 ();
 sg13g2_decap_4 FILLER_2_578 ();
 sg13g2_fill_2 FILLER_2_601 ();
 sg13g2_fill_1 FILLER_2_610 ();
 sg13g2_fill_2 FILLER_2_614 ();
 sg13g2_fill_1 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_621 ();
 sg13g2_decap_8 FILLER_2_628 ();
 sg13g2_decap_8 FILLER_2_635 ();
 sg13g2_decap_4 FILLER_2_642 ();
 sg13g2_fill_2 FILLER_2_646 ();
 sg13g2_decap_8 FILLER_2_652 ();
 sg13g2_decap_8 FILLER_2_659 ();
 sg13g2_decap_8 FILLER_2_666 ();
 sg13g2_fill_2 FILLER_2_673 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_fill_2 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_fill_2 FILLER_2_711 ();
 sg13g2_fill_1 FILLER_2_713 ();
 sg13g2_decap_8 FILLER_2_719 ();
 sg13g2_decap_4 FILLER_2_726 ();
 sg13g2_fill_2 FILLER_2_730 ();
 sg13g2_decap_8 FILLER_2_736 ();
 sg13g2_decap_4 FILLER_2_743 ();
 sg13g2_fill_2 FILLER_2_747 ();
 sg13g2_decap_8 FILLER_2_771 ();
 sg13g2_decap_8 FILLER_2_778 ();
 sg13g2_decap_8 FILLER_2_785 ();
 sg13g2_decap_4 FILLER_2_792 ();
 sg13g2_fill_1 FILLER_2_796 ();
 sg13g2_decap_8 FILLER_2_801 ();
 sg13g2_decap_8 FILLER_2_808 ();
 sg13g2_decap_8 FILLER_2_815 ();
 sg13g2_decap_8 FILLER_2_822 ();
 sg13g2_decap_8 FILLER_2_829 ();
 sg13g2_decap_8 FILLER_2_836 ();
 sg13g2_decap_8 FILLER_2_843 ();
 sg13g2_decap_8 FILLER_2_850 ();
 sg13g2_fill_2 FILLER_2_857 ();
 sg13g2_decap_8 FILLER_2_884 ();
 sg13g2_decap_8 FILLER_2_891 ();
 sg13g2_decap_4 FILLER_2_898 ();
 sg13g2_fill_1 FILLER_2_902 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_4 FILLER_2_914 ();
 sg13g2_fill_1 FILLER_2_918 ();
 sg13g2_decap_8 FILLER_2_923 ();
 sg13g2_decap_4 FILLER_2_930 ();
 sg13g2_decap_8 FILLER_2_939 ();
 sg13g2_fill_1 FILLER_2_946 ();
 sg13g2_decap_8 FILLER_2_978 ();
 sg13g2_fill_2 FILLER_2_996 ();
 sg13g2_fill_2 FILLER_2_1010 ();
 sg13g2_fill_1 FILLER_2_1012 ();
 sg13g2_fill_2 FILLER_2_1028 ();
 sg13g2_fill_1 FILLER_2_1030 ();
 sg13g2_fill_1 FILLER_2_1043 ();
 sg13g2_decap_8 FILLER_2_1048 ();
 sg13g2_decap_4 FILLER_2_1055 ();
 sg13g2_decap_8 FILLER_2_1072 ();
 sg13g2_fill_2 FILLER_2_1079 ();
 sg13g2_fill_1 FILLER_2_1085 ();
 sg13g2_decap_8 FILLER_2_1090 ();
 sg13g2_decap_4 FILLER_2_1097 ();
 sg13g2_fill_2 FILLER_2_1101 ();
 sg13g2_decap_8 FILLER_2_1107 ();
 sg13g2_decap_8 FILLER_2_1114 ();
 sg13g2_decap_8 FILLER_2_1121 ();
 sg13g2_decap_8 FILLER_2_1128 ();
 sg13g2_fill_2 FILLER_2_1135 ();
 sg13g2_fill_1 FILLER_2_1185 ();
 sg13g2_decap_4 FILLER_2_1216 ();
 sg13g2_fill_1 FILLER_2_1220 ();
 sg13g2_decap_8 FILLER_2_1228 ();
 sg13g2_decap_8 FILLER_2_1235 ();
 sg13g2_decap_8 FILLER_2_1242 ();
 sg13g2_decap_8 FILLER_2_1249 ();
 sg13g2_decap_8 FILLER_2_1256 ();
 sg13g2_decap_4 FILLER_2_1263 ();
 sg13g2_fill_2 FILLER_2_1267 ();
 sg13g2_decap_8 FILLER_2_1278 ();
 sg13g2_decap_8 FILLER_2_1285 ();
 sg13g2_decap_8 FILLER_2_1292 ();
 sg13g2_decap_8 FILLER_2_1299 ();
 sg13g2_decap_8 FILLER_2_1306 ();
 sg13g2_decap_8 FILLER_2_1313 ();
 sg13g2_decap_4 FILLER_2_1320 ();
 sg13g2_fill_2 FILLER_2_1324 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_4 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_32 ();
 sg13g2_decap_4 FILLER_3_63 ();
 sg13g2_fill_1 FILLER_3_75 ();
 sg13g2_decap_4 FILLER_3_91 ();
 sg13g2_fill_1 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_101 ();
 sg13g2_decap_4 FILLER_3_108 ();
 sg13g2_fill_1 FILLER_3_112 ();
 sg13g2_decap_4 FILLER_3_121 ();
 sg13g2_fill_1 FILLER_3_125 ();
 sg13g2_decap_4 FILLER_3_167 ();
 sg13g2_fill_1 FILLER_3_185 ();
 sg13g2_fill_1 FILLER_3_190 ();
 sg13g2_fill_2 FILLER_3_194 ();
 sg13g2_fill_1 FILLER_3_204 ();
 sg13g2_fill_1 FILLER_3_248 ();
 sg13g2_fill_2 FILLER_3_256 ();
 sg13g2_decap_4 FILLER_3_272 ();
 sg13g2_fill_2 FILLER_3_276 ();
 sg13g2_decap_8 FILLER_3_292 ();
 sg13g2_decap_8 FILLER_3_310 ();
 sg13g2_fill_1 FILLER_3_317 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_4 FILLER_3_398 ();
 sg13g2_fill_1 FILLER_3_405 ();
 sg13g2_decap_4 FILLER_3_414 ();
 sg13g2_fill_1 FILLER_3_418 ();
 sg13g2_decap_8 FILLER_3_426 ();
 sg13g2_decap_4 FILLER_3_433 ();
 sg13g2_fill_1 FILLER_3_437 ();
 sg13g2_decap_8 FILLER_3_464 ();
 sg13g2_decap_8 FILLER_3_471 ();
 sg13g2_fill_2 FILLER_3_478 ();
 sg13g2_fill_1 FILLER_3_480 ();
 sg13g2_fill_1 FILLER_3_484 ();
 sg13g2_fill_2 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_512 ();
 sg13g2_decap_8 FILLER_3_519 ();
 sg13g2_decap_4 FILLER_3_526 ();
 sg13g2_fill_2 FILLER_3_530 ();
 sg13g2_fill_2 FILLER_3_536 ();
 sg13g2_fill_1 FILLER_3_538 ();
 sg13g2_decap_8 FILLER_3_544 ();
 sg13g2_fill_1 FILLER_3_551 ();
 sg13g2_decap_8 FILLER_3_578 ();
 sg13g2_fill_2 FILLER_3_585 ();
 sg13g2_fill_2 FILLER_3_612 ();
 sg13g2_fill_1 FILLER_3_633 ();
 sg13g2_fill_1 FILLER_3_640 ();
 sg13g2_decap_8 FILLER_3_645 ();
 sg13g2_decap_8 FILLER_3_652 ();
 sg13g2_fill_2 FILLER_3_659 ();
 sg13g2_fill_1 FILLER_3_661 ();
 sg13g2_fill_1 FILLER_3_709 ();
 sg13g2_fill_2 FILLER_3_736 ();
 sg13g2_fill_2 FILLER_3_768 ();
 sg13g2_fill_1 FILLER_3_905 ();
 sg13g2_fill_1 FILLER_3_932 ();
 sg13g2_fill_1 FILLER_3_936 ();
 sg13g2_fill_1 FILLER_3_942 ();
 sg13g2_fill_2 FILLER_3_947 ();
 sg13g2_decap_8 FILLER_3_956 ();
 sg13g2_decap_8 FILLER_3_963 ();
 sg13g2_decap_4 FILLER_3_970 ();
 sg13g2_fill_2 FILLER_3_974 ();
 sg13g2_decap_8 FILLER_3_979 ();
 sg13g2_decap_8 FILLER_3_986 ();
 sg13g2_decap_4 FILLER_3_993 ();
 sg13g2_fill_1 FILLER_3_997 ();
 sg13g2_fill_2 FILLER_3_1005 ();
 sg13g2_decap_4 FILLER_3_1021 ();
 sg13g2_fill_1 FILLER_3_1035 ();
 sg13g2_fill_2 FILLER_3_1062 ();
 sg13g2_fill_1 FILLER_3_1064 ();
 sg13g2_decap_4 FILLER_3_1078 ();
 sg13g2_decap_4 FILLER_3_1094 ();
 sg13g2_fill_1 FILLER_3_1098 ();
 sg13g2_decap_8 FILLER_3_1149 ();
 sg13g2_decap_8 FILLER_3_1156 ();
 sg13g2_decap_8 FILLER_3_1163 ();
 sg13g2_decap_8 FILLER_3_1170 ();
 sg13g2_decap_8 FILLER_3_1177 ();
 sg13g2_fill_1 FILLER_3_1184 ();
 sg13g2_decap_8 FILLER_3_1195 ();
 sg13g2_decap_8 FILLER_3_1202 ();
 sg13g2_fill_2 FILLER_3_1209 ();
 sg13g2_decap_8 FILLER_3_1250 ();
 sg13g2_decap_8 FILLER_3_1257 ();
 sg13g2_fill_2 FILLER_3_1264 ();
 sg13g2_decap_8 FILLER_3_1296 ();
 sg13g2_decap_8 FILLER_3_1303 ();
 sg13g2_decap_8 FILLER_3_1310 ();
 sg13g2_decap_8 FILLER_3_1317 ();
 sg13g2_fill_2 FILLER_3_1324 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_4 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_60 ();
 sg13g2_fill_2 FILLER_4_67 ();
 sg13g2_fill_2 FILLER_4_73 ();
 sg13g2_fill_1 FILLER_4_75 ();
 sg13g2_fill_2 FILLER_4_102 ();
 sg13g2_fill_2 FILLER_4_139 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_fill_2 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_175 ();
 sg13g2_fill_2 FILLER_4_184 ();
 sg13g2_fill_1 FILLER_4_200 ();
 sg13g2_fill_2 FILLER_4_205 ();
 sg13g2_fill_1 FILLER_4_222 ();
 sg13g2_fill_2 FILLER_4_230 ();
 sg13g2_fill_1 FILLER_4_237 ();
 sg13g2_fill_2 FILLER_4_255 ();
 sg13g2_fill_1 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_268 ();
 sg13g2_fill_2 FILLER_4_275 ();
 sg13g2_fill_1 FILLER_4_277 ();
 sg13g2_fill_1 FILLER_4_290 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_314 ();
 sg13g2_decap_8 FILLER_4_321 ();
 sg13g2_decap_8 FILLER_4_328 ();
 sg13g2_decap_8 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_355 ();
 sg13g2_decap_8 FILLER_4_362 ();
 sg13g2_decap_8 FILLER_4_369 ();
 sg13g2_decap_8 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_383 ();
 sg13g2_decap_4 FILLER_4_390 ();
 sg13g2_fill_1 FILLER_4_394 ();
 sg13g2_fill_2 FILLER_4_399 ();
 sg13g2_fill_1 FILLER_4_418 ();
 sg13g2_decap_4 FILLER_4_424 ();
 sg13g2_fill_2 FILLER_4_428 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_4 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_477 ();
 sg13g2_fill_2 FILLER_4_484 ();
 sg13g2_fill_1 FILLER_4_486 ();
 sg13g2_decap_4 FILLER_4_491 ();
 sg13g2_fill_1 FILLER_4_495 ();
 sg13g2_fill_2 FILLER_4_504 ();
 sg13g2_fill_2 FILLER_4_515 ();
 sg13g2_fill_1 FILLER_4_523 ();
 sg13g2_fill_1 FILLER_4_554 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_611 ();
 sg13g2_fill_2 FILLER_4_618 ();
 sg13g2_fill_1 FILLER_4_620 ();
 sg13g2_fill_2 FILLER_4_635 ();
 sg13g2_fill_1 FILLER_4_637 ();
 sg13g2_fill_1 FILLER_4_647 ();
 sg13g2_fill_1 FILLER_4_652 ();
 sg13g2_fill_1 FILLER_4_657 ();
 sg13g2_fill_1 FILLER_4_663 ();
 sg13g2_fill_1 FILLER_4_668 ();
 sg13g2_fill_1 FILLER_4_677 ();
 sg13g2_decap_8 FILLER_4_682 ();
 sg13g2_decap_8 FILLER_4_689 ();
 sg13g2_decap_4 FILLER_4_696 ();
 sg13g2_fill_2 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_705 ();
 sg13g2_fill_1 FILLER_4_712 ();
 sg13g2_fill_1 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_decap_8 FILLER_4_734 ();
 sg13g2_fill_2 FILLER_4_741 ();
 sg13g2_decap_8 FILLER_4_747 ();
 sg13g2_decap_8 FILLER_4_754 ();
 sg13g2_fill_2 FILLER_4_761 ();
 sg13g2_fill_1 FILLER_4_767 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_4 FILLER_4_784 ();
 sg13g2_fill_2 FILLER_4_788 ();
 sg13g2_fill_2 FILLER_4_794 ();
 sg13g2_fill_1 FILLER_4_796 ();
 sg13g2_decap_4 FILLER_4_806 ();
 sg13g2_decap_8 FILLER_4_813 ();
 sg13g2_decap_8 FILLER_4_820 ();
 sg13g2_decap_8 FILLER_4_827 ();
 sg13g2_decap_4 FILLER_4_834 ();
 sg13g2_fill_1 FILLER_4_842 ();
 sg13g2_decap_8 FILLER_4_852 ();
 sg13g2_fill_1 FILLER_4_859 ();
 sg13g2_fill_2 FILLER_4_865 ();
 sg13g2_fill_1 FILLER_4_867 ();
 sg13g2_decap_4 FILLER_4_871 ();
 sg13g2_fill_2 FILLER_4_875 ();
 sg13g2_decap_8 FILLER_4_882 ();
 sg13g2_decap_4 FILLER_4_889 ();
 sg13g2_decap_8 FILLER_4_896 ();
 sg13g2_decap_8 FILLER_4_903 ();
 sg13g2_decap_8 FILLER_4_910 ();
 sg13g2_decap_8 FILLER_4_917 ();
 sg13g2_fill_2 FILLER_4_944 ();
 sg13g2_fill_1 FILLER_4_946 ();
 sg13g2_fill_2 FILLER_4_950 ();
 sg13g2_fill_1 FILLER_4_964 ();
 sg13g2_decap_8 FILLER_4_968 ();
 sg13g2_decap_8 FILLER_4_975 ();
 sg13g2_fill_2 FILLER_4_982 ();
 sg13g2_fill_1 FILLER_4_984 ();
 sg13g2_fill_1 FILLER_4_1012 ();
 sg13g2_fill_1 FILLER_4_1017 ();
 sg13g2_decap_8 FILLER_4_1026 ();
 sg13g2_decap_8 FILLER_4_1033 ();
 sg13g2_decap_8 FILLER_4_1040 ();
 sg13g2_decap_8 FILLER_4_1047 ();
 sg13g2_decap_4 FILLER_4_1054 ();
 sg13g2_decap_4 FILLER_4_1062 ();
 sg13g2_fill_1 FILLER_4_1066 ();
 sg13g2_decap_8 FILLER_4_1070 ();
 sg13g2_fill_2 FILLER_4_1077 ();
 sg13g2_fill_2 FILLER_4_1116 ();
 sg13g2_decap_8 FILLER_4_1131 ();
 sg13g2_decap_4 FILLER_4_1138 ();
 sg13g2_decap_8 FILLER_4_1197 ();
 sg13g2_decap_8 FILLER_4_1204 ();
 sg13g2_decap_8 FILLER_4_1211 ();
 sg13g2_decap_8 FILLER_4_1218 ();
 sg13g2_decap_8 FILLER_4_1225 ();
 sg13g2_decap_8 FILLER_4_1232 ();
 sg13g2_fill_2 FILLER_4_1239 ();
 sg13g2_fill_1 FILLER_4_1241 ();
 sg13g2_decap_8 FILLER_4_1298 ();
 sg13g2_decap_8 FILLER_4_1305 ();
 sg13g2_decap_8 FILLER_4_1312 ();
 sg13g2_decap_8 FILLER_4_1319 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_33 ();
 sg13g2_decap_4 FILLER_5_45 ();
 sg13g2_fill_1 FILLER_5_49 ();
 sg13g2_fill_2 FILLER_5_76 ();
 sg13g2_fill_1 FILLER_5_78 ();
 sg13g2_fill_2 FILLER_5_87 ();
 sg13g2_fill_2 FILLER_5_99 ();
 sg13g2_fill_1 FILLER_5_101 ();
 sg13g2_decap_4 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_138 ();
 sg13g2_fill_1 FILLER_5_145 ();
 sg13g2_decap_4 FILLER_5_150 ();
 sg13g2_fill_1 FILLER_5_180 ();
 sg13g2_fill_1 FILLER_5_189 ();
 sg13g2_fill_2 FILLER_5_195 ();
 sg13g2_fill_1 FILLER_5_197 ();
 sg13g2_fill_2 FILLER_5_203 ();
 sg13g2_fill_1 FILLER_5_205 ();
 sg13g2_fill_2 FILLER_5_229 ();
 sg13g2_fill_2 FILLER_5_262 ();
 sg13g2_decap_4 FILLER_5_274 ();
 sg13g2_fill_2 FILLER_5_278 ();
 sg13g2_fill_1 FILLER_5_285 ();
 sg13g2_decap_4 FILLER_5_295 ();
 sg13g2_fill_2 FILLER_5_318 ();
 sg13g2_fill_1 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_332 ();
 sg13g2_fill_1 FILLER_5_339 ();
 sg13g2_decap_4 FILLER_5_366 ();
 sg13g2_fill_2 FILLER_5_370 ();
 sg13g2_decap_8 FILLER_5_377 ();
 sg13g2_fill_1 FILLER_5_384 ();
 sg13g2_fill_1 FILLER_5_407 ();
 sg13g2_fill_1 FILLER_5_412 ();
 sg13g2_fill_1 FILLER_5_418 ();
 sg13g2_fill_2 FILLER_5_422 ();
 sg13g2_fill_1 FILLER_5_431 ();
 sg13g2_fill_2 FILLER_5_437 ();
 sg13g2_fill_1 FILLER_5_439 ();
 sg13g2_fill_1 FILLER_5_447 ();
 sg13g2_fill_1 FILLER_5_460 ();
 sg13g2_fill_1 FILLER_5_469 ();
 sg13g2_decap_4 FILLER_5_475 ();
 sg13g2_fill_2 FILLER_5_479 ();
 sg13g2_decap_4 FILLER_5_485 ();
 sg13g2_fill_2 FILLER_5_489 ();
 sg13g2_fill_2 FILLER_5_494 ();
 sg13g2_fill_2 FILLER_5_520 ();
 sg13g2_fill_2 FILLER_5_554 ();
 sg13g2_decap_4 FILLER_5_564 ();
 sg13g2_fill_2 FILLER_5_568 ();
 sg13g2_fill_2 FILLER_5_589 ();
 sg13g2_fill_1 FILLER_5_599 ();
 sg13g2_fill_1 FILLER_5_604 ();
 sg13g2_decap_4 FILLER_5_615 ();
 sg13g2_decap_8 FILLER_5_632 ();
 sg13g2_decap_8 FILLER_5_639 ();
 sg13g2_decap_4 FILLER_5_646 ();
 sg13g2_fill_1 FILLER_5_650 ();
 sg13g2_decap_4 FILLER_5_663 ();
 sg13g2_fill_1 FILLER_5_671 ();
 sg13g2_decap_4 FILLER_5_689 ();
 sg13g2_fill_2 FILLER_5_698 ();
 sg13g2_decap_8 FILLER_5_703 ();
 sg13g2_fill_2 FILLER_5_710 ();
 sg13g2_fill_1 FILLER_5_712 ();
 sg13g2_fill_1 FILLER_5_726 ();
 sg13g2_decap_4 FILLER_5_757 ();
 sg13g2_fill_2 FILLER_5_766 ();
 sg13g2_decap_4 FILLER_5_773 ();
 sg13g2_fill_1 FILLER_5_777 ();
 sg13g2_fill_1 FILLER_5_786 ();
 sg13g2_fill_1 FILLER_5_790 ();
 sg13g2_decap_8 FILLER_5_799 ();
 sg13g2_fill_2 FILLER_5_806 ();
 sg13g2_fill_1 FILLER_5_816 ();
 sg13g2_fill_1 FILLER_5_823 ();
 sg13g2_fill_1 FILLER_5_832 ();
 sg13g2_decap_4 FILLER_5_836 ();
 sg13g2_fill_2 FILLER_5_840 ();
 sg13g2_decap_4 FILLER_5_852 ();
 sg13g2_fill_1 FILLER_5_856 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_4 FILLER_5_882 ();
 sg13g2_fill_2 FILLER_5_886 ();
 sg13g2_decap_4 FILLER_5_896 ();
 sg13g2_fill_1 FILLER_5_900 ();
 sg13g2_decap_8 FILLER_5_906 ();
 sg13g2_decap_8 FILLER_5_913 ();
 sg13g2_decap_4 FILLER_5_928 ();
 sg13g2_fill_2 FILLER_5_941 ();
 sg13g2_fill_1 FILLER_5_943 ();
 sg13g2_fill_1 FILLER_5_948 ();
 sg13g2_decap_8 FILLER_5_957 ();
 sg13g2_decap_4 FILLER_5_964 ();
 sg13g2_decap_8 FILLER_5_981 ();
 sg13g2_decap_4 FILLER_5_988 ();
 sg13g2_fill_2 FILLER_5_992 ();
 sg13g2_fill_1 FILLER_5_1011 ();
 sg13g2_fill_1 FILLER_5_1016 ();
 sg13g2_decap_8 FILLER_5_1022 ();
 sg13g2_decap_8 FILLER_5_1029 ();
 sg13g2_decap_8 FILLER_5_1036 ();
 sg13g2_decap_8 FILLER_5_1043 ();
 sg13g2_decap_8 FILLER_5_1050 ();
 sg13g2_decap_8 FILLER_5_1057 ();
 sg13g2_decap_8 FILLER_5_1064 ();
 sg13g2_fill_2 FILLER_5_1071 ();
 sg13g2_decap_4 FILLER_5_1084 ();
 sg13g2_fill_2 FILLER_5_1092 ();
 sg13g2_decap_8 FILLER_5_1105 ();
 sg13g2_fill_1 FILLER_5_1112 ();
 sg13g2_fill_2 FILLER_5_1131 ();
 sg13g2_fill_1 FILLER_5_1141 ();
 sg13g2_fill_1 FILLER_5_1150 ();
 sg13g2_fill_2 FILLER_5_1159 ();
 sg13g2_decap_8 FILLER_5_1170 ();
 sg13g2_decap_4 FILLER_5_1177 ();
 sg13g2_fill_1 FILLER_5_1181 ();
 sg13g2_decap_4 FILLER_5_1191 ();
 sg13g2_fill_2 FILLER_5_1199 ();
 sg13g2_fill_1 FILLER_5_1201 ();
 sg13g2_decap_8 FILLER_5_1207 ();
 sg13g2_decap_8 FILLER_5_1214 ();
 sg13g2_decap_8 FILLER_5_1221 ();
 sg13g2_fill_2 FILLER_5_1231 ();
 sg13g2_fill_2 FILLER_5_1238 ();
 sg13g2_fill_1 FILLER_5_1240 ();
 sg13g2_decap_8 FILLER_5_1253 ();
 sg13g2_fill_2 FILLER_5_1260 ();
 sg13g2_decap_8 FILLER_5_1279 ();
 sg13g2_decap_8 FILLER_5_1286 ();
 sg13g2_decap_8 FILLER_5_1293 ();
 sg13g2_decap_8 FILLER_5_1300 ();
 sg13g2_decap_8 FILLER_5_1307 ();
 sg13g2_decap_8 FILLER_5_1314 ();
 sg13g2_decap_4 FILLER_5_1321 ();
 sg13g2_fill_1 FILLER_5_1325 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_12 ();
 sg13g2_decap_4 FILLER_6_19 ();
 sg13g2_fill_2 FILLER_6_27 ();
 sg13g2_decap_8 FILLER_6_59 ();
 sg13g2_decap_4 FILLER_6_66 ();
 sg13g2_fill_2 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_82 ();
 sg13g2_fill_1 FILLER_6_101 ();
 sg13g2_decap_8 FILLER_6_110 ();
 sg13g2_decap_8 FILLER_6_117 ();
 sg13g2_decap_8 FILLER_6_124 ();
 sg13g2_fill_2 FILLER_6_131 ();
 sg13g2_fill_1 FILLER_6_198 ();
 sg13g2_decap_4 FILLER_6_202 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_decap_4 FILLER_6_242 ();
 sg13g2_fill_1 FILLER_6_246 ();
 sg13g2_fill_1 FILLER_6_272 ();
 sg13g2_fill_2 FILLER_6_281 ();
 sg13g2_fill_1 FILLER_6_283 ();
 sg13g2_fill_1 FILLER_6_289 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_4 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_331 ();
 sg13g2_fill_2 FILLER_6_338 ();
 sg13g2_decap_4 FILLER_6_356 ();
 sg13g2_fill_1 FILLER_6_363 ();
 sg13g2_fill_2 FILLER_6_381 ();
 sg13g2_fill_1 FILLER_6_383 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_4 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_414 ();
 sg13g2_fill_1 FILLER_6_419 ();
 sg13g2_decap_4 FILLER_6_425 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_4 FILLER_6_434 ();
 sg13g2_fill_2 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_447 ();
 sg13g2_fill_2 FILLER_6_454 ();
 sg13g2_decap_4 FILLER_6_459 ();
 sg13g2_fill_2 FILLER_6_463 ();
 sg13g2_fill_1 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_475 ();
 sg13g2_fill_1 FILLER_6_482 ();
 sg13g2_fill_1 FILLER_6_488 ();
 sg13g2_fill_2 FILLER_6_494 ();
 sg13g2_fill_1 FILLER_6_500 ();
 sg13g2_fill_2 FILLER_6_518 ();
 sg13g2_fill_2 FILLER_6_528 ();
 sg13g2_fill_2 FILLER_6_536 ();
 sg13g2_fill_1 FILLER_6_538 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_575 ();
 sg13g2_decap_4 FILLER_6_582 ();
 sg13g2_fill_1 FILLER_6_586 ();
 sg13g2_decap_4 FILLER_6_597 ();
 sg13g2_fill_1 FILLER_6_606 ();
 sg13g2_fill_2 FILLER_6_612 ();
 sg13g2_decap_8 FILLER_6_618 ();
 sg13g2_decap_8 FILLER_6_625 ();
 sg13g2_decap_8 FILLER_6_632 ();
 sg13g2_decap_8 FILLER_6_639 ();
 sg13g2_fill_2 FILLER_6_646 ();
 sg13g2_fill_1 FILLER_6_648 ();
 sg13g2_fill_1 FILLER_6_653 ();
 sg13g2_fill_1 FILLER_6_659 ();
 sg13g2_fill_1 FILLER_6_664 ();
 sg13g2_fill_2 FILLER_6_670 ();
 sg13g2_fill_2 FILLER_6_677 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_4 FILLER_6_739 ();
 sg13g2_fill_1 FILLER_6_743 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_fill_2 FILLER_6_803 ();
 sg13g2_fill_1 FILLER_6_810 ();
 sg13g2_fill_2 FILLER_6_869 ();
 sg13g2_fill_2 FILLER_6_883 ();
 sg13g2_decap_8 FILLER_6_890 ();
 sg13g2_fill_1 FILLER_6_919 ();
 sg13g2_decap_4 FILLER_6_939 ();
 sg13g2_fill_2 FILLER_6_961 ();
 sg13g2_decap_8 FILLER_6_973 ();
 sg13g2_decap_8 FILLER_6_980 ();
 sg13g2_fill_2 FILLER_6_987 ();
 sg13g2_fill_2 FILLER_6_1001 ();
 sg13g2_decap_4 FILLER_6_1006 ();
 sg13g2_fill_2 FILLER_6_1010 ();
 sg13g2_fill_1 FILLER_6_1017 ();
 sg13g2_decap_4 FILLER_6_1037 ();
 sg13g2_fill_2 FILLER_6_1121 ();
 sg13g2_fill_1 FILLER_6_1190 ();
 sg13g2_fill_2 FILLER_6_1194 ();
 sg13g2_fill_2 FILLER_6_1201 ();
 sg13g2_fill_2 FILLER_6_1206 ();
 sg13g2_fill_1 FILLER_6_1237 ();
 sg13g2_decap_4 FILLER_6_1254 ();
 sg13g2_fill_1 FILLER_6_1258 ();
 sg13g2_decap_8 FILLER_6_1272 ();
 sg13g2_decap_8 FILLER_6_1279 ();
 sg13g2_decap_8 FILLER_6_1286 ();
 sg13g2_decap_8 FILLER_6_1293 ();
 sg13g2_decap_8 FILLER_6_1300 ();
 sg13g2_decap_8 FILLER_6_1307 ();
 sg13g2_decap_8 FILLER_6_1314 ();
 sg13g2_decap_4 FILLER_6_1321 ();
 sg13g2_fill_1 FILLER_6_1325 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_12 ();
 sg13g2_decap_8 FILLER_7_17 ();
 sg13g2_decap_8 FILLER_7_24 ();
 sg13g2_decap_8 FILLER_7_31 ();
 sg13g2_decap_4 FILLER_7_38 ();
 sg13g2_fill_2 FILLER_7_42 ();
 sg13g2_fill_2 FILLER_7_47 ();
 sg13g2_fill_1 FILLER_7_49 ();
 sg13g2_decap_4 FILLER_7_57 ();
 sg13g2_fill_2 FILLER_7_61 ();
 sg13g2_decap_4 FILLER_7_92 ();
 sg13g2_decap_8 FILLER_7_100 ();
 sg13g2_decap_4 FILLER_7_107 ();
 sg13g2_fill_1 FILLER_7_111 ();
 sg13g2_fill_2 FILLER_7_115 ();
 sg13g2_fill_1 FILLER_7_120 ();
 sg13g2_fill_2 FILLER_7_141 ();
 sg13g2_decap_8 FILLER_7_151 ();
 sg13g2_decap_8 FILLER_7_158 ();
 sg13g2_decap_8 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_172 ();
 sg13g2_fill_1 FILLER_7_174 ();
 sg13g2_fill_2 FILLER_7_178 ();
 sg13g2_fill_1 FILLER_7_180 ();
 sg13g2_decap_8 FILLER_7_187 ();
 sg13g2_decap_8 FILLER_7_194 ();
 sg13g2_decap_4 FILLER_7_201 ();
 sg13g2_fill_2 FILLER_7_205 ();
 sg13g2_decap_4 FILLER_7_211 ();
 sg13g2_fill_1 FILLER_7_215 ();
 sg13g2_decap_4 FILLER_7_228 ();
 sg13g2_fill_2 FILLER_7_232 ();
 sg13g2_decap_8 FILLER_7_246 ();
 sg13g2_decap_4 FILLER_7_253 ();
 sg13g2_fill_2 FILLER_7_257 ();
 sg13g2_decap_4 FILLER_7_266 ();
 sg13g2_decap_4 FILLER_7_298 ();
 sg13g2_fill_2 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_fill_2 FILLER_7_348 ();
 sg13g2_fill_1 FILLER_7_350 ();
 sg13g2_fill_1 FILLER_7_363 ();
 sg13g2_fill_2 FILLER_7_377 ();
 sg13g2_fill_1 FILLER_7_379 ();
 sg13g2_fill_2 FILLER_7_424 ();
 sg13g2_decap_4 FILLER_7_435 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_4 FILLER_7_455 ();
 sg13g2_fill_2 FILLER_7_459 ();
 sg13g2_decap_8 FILLER_7_477 ();
 sg13g2_fill_2 FILLER_7_500 ();
 sg13g2_fill_2 FILLER_7_571 ();
 sg13g2_fill_2 FILLER_7_582 ();
 sg13g2_fill_1 FILLER_7_584 ();
 sg13g2_fill_1 FILLER_7_599 ();
 sg13g2_decap_4 FILLER_7_609 ();
 sg13g2_fill_2 FILLER_7_622 ();
 sg13g2_fill_1 FILLER_7_624 ();
 sg13g2_decap_8 FILLER_7_628 ();
 sg13g2_fill_2 FILLER_7_635 ();
 sg13g2_fill_1 FILLER_7_637 ();
 sg13g2_fill_1 FILLER_7_662 ();
 sg13g2_fill_1 FILLER_7_670 ();
 sg13g2_fill_1 FILLER_7_675 ();
 sg13g2_fill_1 FILLER_7_681 ();
 sg13g2_fill_1 FILLER_7_687 ();
 sg13g2_decap_8 FILLER_7_691 ();
 sg13g2_fill_2 FILLER_7_698 ();
 sg13g2_fill_1 FILLER_7_700 ();
 sg13g2_fill_2 FILLER_7_714 ();
 sg13g2_fill_1 FILLER_7_716 ();
 sg13g2_decap_8 FILLER_7_722 ();
 sg13g2_decap_8 FILLER_7_729 ();
 sg13g2_decap_8 FILLER_7_736 ();
 sg13g2_decap_8 FILLER_7_743 ();
 sg13g2_decap_4 FILLER_7_750 ();
 sg13g2_fill_2 FILLER_7_754 ();
 sg13g2_decap_8 FILLER_7_768 ();
 sg13g2_fill_2 FILLER_7_775 ();
 sg13g2_fill_1 FILLER_7_777 ();
 sg13g2_fill_1 FILLER_7_781 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_fill_2 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_820 ();
 sg13g2_fill_2 FILLER_7_827 ();
 sg13g2_fill_2 FILLER_7_832 ();
 sg13g2_decap_4 FILLER_7_837 ();
 sg13g2_fill_2 FILLER_7_856 ();
 sg13g2_fill_1 FILLER_7_858 ();
 sg13g2_fill_2 FILLER_7_869 ();
 sg13g2_decap_8 FILLER_7_880 ();
 sg13g2_decap_8 FILLER_7_887 ();
 sg13g2_decap_8 FILLER_7_894 ();
 sg13g2_decap_8 FILLER_7_901 ();
 sg13g2_decap_4 FILLER_7_911 ();
 sg13g2_decap_8 FILLER_7_919 ();
 sg13g2_decap_4 FILLER_7_926 ();
 sg13g2_decap_4 FILLER_7_935 ();
 sg13g2_fill_2 FILLER_7_943 ();
 sg13g2_fill_1 FILLER_7_953 ();
 sg13g2_fill_1 FILLER_7_959 ();
 sg13g2_decap_8 FILLER_7_963 ();
 sg13g2_decap_8 FILLER_7_970 ();
 sg13g2_decap_8 FILLER_7_977 ();
 sg13g2_decap_8 FILLER_7_984 ();
 sg13g2_decap_8 FILLER_7_991 ();
 sg13g2_fill_2 FILLER_7_1006 ();
 sg13g2_fill_1 FILLER_7_1021 ();
 sg13g2_decap_4 FILLER_7_1032 ();
 sg13g2_fill_2 FILLER_7_1052 ();
 sg13g2_fill_2 FILLER_7_1065 ();
 sg13g2_fill_1 FILLER_7_1067 ();
 sg13g2_decap_8 FILLER_7_1072 ();
 sg13g2_decap_4 FILLER_7_1079 ();
 sg13g2_fill_1 FILLER_7_1083 ();
 sg13g2_decap_4 FILLER_7_1093 ();
 sg13g2_decap_8 FILLER_7_1101 ();
 sg13g2_fill_1 FILLER_7_1108 ();
 sg13g2_decap_8 FILLER_7_1128 ();
 sg13g2_fill_1 FILLER_7_1144 ();
 sg13g2_fill_2 FILLER_7_1148 ();
 sg13g2_decap_8 FILLER_7_1158 ();
 sg13g2_decap_8 FILLER_7_1165 ();
 sg13g2_decap_8 FILLER_7_1172 ();
 sg13g2_decap_8 FILLER_7_1179 ();
 sg13g2_fill_2 FILLER_7_1204 ();
 sg13g2_fill_1 FILLER_7_1206 ();
 sg13g2_fill_1 FILLER_7_1212 ();
 sg13g2_fill_2 FILLER_7_1223 ();
 sg13g2_fill_2 FILLER_7_1243 ();
 sg13g2_fill_2 FILLER_7_1249 ();
 sg13g2_fill_2 FILLER_7_1254 ();
 sg13g2_fill_1 FILLER_7_1256 ();
 sg13g2_fill_2 FILLER_7_1265 ();
 sg13g2_decap_8 FILLER_7_1273 ();
 sg13g2_fill_2 FILLER_7_1280 ();
 sg13g2_fill_1 FILLER_7_1286 ();
 sg13g2_decap_8 FILLER_7_1292 ();
 sg13g2_decap_8 FILLER_7_1299 ();
 sg13g2_decap_8 FILLER_7_1306 ();
 sg13g2_decap_8 FILLER_7_1313 ();
 sg13g2_decap_4 FILLER_7_1320 ();
 sg13g2_fill_2 FILLER_7_1324 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_35 ();
 sg13g2_fill_2 FILLER_8_39 ();
 sg13g2_fill_1 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_61 ();
 sg13g2_decap_8 FILLER_8_68 ();
 sg13g2_fill_2 FILLER_8_75 ();
 sg13g2_fill_1 FILLER_8_80 ();
 sg13g2_fill_1 FILLER_8_85 ();
 sg13g2_fill_2 FILLER_8_90 ();
 sg13g2_fill_1 FILLER_8_99 ();
 sg13g2_fill_2 FILLER_8_123 ();
 sg13g2_fill_2 FILLER_8_138 ();
 sg13g2_fill_1 FILLER_8_161 ();
 sg13g2_fill_2 FILLER_8_166 ();
 sg13g2_decap_8 FILLER_8_171 ();
 sg13g2_decap_8 FILLER_8_178 ();
 sg13g2_fill_2 FILLER_8_185 ();
 sg13g2_fill_1 FILLER_8_187 ();
 sg13g2_decap_4 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_222 ();
 sg13g2_fill_2 FILLER_8_232 ();
 sg13g2_fill_1 FILLER_8_251 ();
 sg13g2_fill_2 FILLER_8_309 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_327 ();
 sg13g2_fill_2 FILLER_8_354 ();
 sg13g2_fill_1 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_fill_1 FILLER_8_377 ();
 sg13g2_decap_4 FILLER_8_384 ();
 sg13g2_fill_1 FILLER_8_409 ();
 sg13g2_fill_2 FILLER_8_426 ();
 sg13g2_fill_2 FILLER_8_433 ();
 sg13g2_fill_1 FILLER_8_435 ();
 sg13g2_decap_8 FILLER_8_444 ();
 sg13g2_decap_8 FILLER_8_451 ();
 sg13g2_decap_8 FILLER_8_458 ();
 sg13g2_fill_2 FILLER_8_465 ();
 sg13g2_decap_4 FILLER_8_476 ();
 sg13g2_fill_2 FILLER_8_480 ();
 sg13g2_fill_1 FILLER_8_504 ();
 sg13g2_fill_1 FILLER_8_515 ();
 sg13g2_fill_2 FILLER_8_534 ();
 sg13g2_fill_2 FILLER_8_551 ();
 sg13g2_fill_1 FILLER_8_553 ();
 sg13g2_fill_2 FILLER_8_566 ();
 sg13g2_fill_1 FILLER_8_577 ();
 sg13g2_decap_4 FILLER_8_593 ();
 sg13g2_decap_4 FILLER_8_610 ();
 sg13g2_decap_4 FILLER_8_640 ();
 sg13g2_fill_1 FILLER_8_644 ();
 sg13g2_fill_2 FILLER_8_657 ();
 sg13g2_decap_8 FILLER_8_668 ();
 sg13g2_decap_8 FILLER_8_675 ();
 sg13g2_fill_2 FILLER_8_682 ();
 sg13g2_fill_1 FILLER_8_684 ();
 sg13g2_fill_2 FILLER_8_688 ();
 sg13g2_fill_2 FILLER_8_695 ();
 sg13g2_fill_1 FILLER_8_697 ();
 sg13g2_fill_1 FILLER_8_702 ();
 sg13g2_decap_4 FILLER_8_722 ();
 sg13g2_decap_8 FILLER_8_730 ();
 sg13g2_decap_8 FILLER_8_737 ();
 sg13g2_decap_4 FILLER_8_744 ();
 sg13g2_fill_1 FILLER_8_748 ();
 sg13g2_decap_4 FILLER_8_757 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_fill_1 FILLER_8_791 ();
 sg13g2_fill_1 FILLER_8_797 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_fill_2 FILLER_8_826 ();
 sg13g2_fill_2 FILLER_8_835 ();
 sg13g2_fill_2 FILLER_8_842 ();
 sg13g2_fill_2 FILLER_8_853 ();
 sg13g2_fill_2 FILLER_8_875 ();
 sg13g2_fill_2 FILLER_8_897 ();
 sg13g2_fill_1 FILLER_8_899 ();
 sg13g2_fill_1 FILLER_8_904 ();
 sg13g2_decap_4 FILLER_8_914 ();
 sg13g2_fill_2 FILLER_8_918 ();
 sg13g2_decap_4 FILLER_8_926 ();
 sg13g2_decap_4 FILLER_8_939 ();
 sg13g2_fill_2 FILLER_8_962 ();
 sg13g2_fill_1 FILLER_8_964 ();
 sg13g2_decap_8 FILLER_8_974 ();
 sg13g2_decap_4 FILLER_8_981 ();
 sg13g2_fill_1 FILLER_8_985 ();
 sg13g2_decap_4 FILLER_8_995 ();
 sg13g2_fill_2 FILLER_8_1005 ();
 sg13g2_fill_1 FILLER_8_1007 ();
 sg13g2_fill_2 FILLER_8_1012 ();
 sg13g2_fill_1 FILLER_8_1014 ();
 sg13g2_fill_2 FILLER_8_1029 ();
 sg13g2_fill_2 FILLER_8_1044 ();
 sg13g2_decap_4 FILLER_8_1054 ();
 sg13g2_fill_1 FILLER_8_1064 ();
 sg13g2_fill_1 FILLER_8_1069 ();
 sg13g2_fill_2 FILLER_8_1075 ();
 sg13g2_fill_2 FILLER_8_1084 ();
 sg13g2_fill_1 FILLER_8_1086 ();
 sg13g2_fill_1 FILLER_8_1105 ();
 sg13g2_fill_2 FILLER_8_1110 ();
 sg13g2_fill_1 FILLER_8_1116 ();
 sg13g2_decap_8 FILLER_8_1121 ();
 sg13g2_decap_4 FILLER_8_1128 ();
 sg13g2_decap_8 FILLER_8_1136 ();
 sg13g2_decap_8 FILLER_8_1143 ();
 sg13g2_fill_2 FILLER_8_1150 ();
 sg13g2_fill_1 FILLER_8_1158 ();
 sg13g2_decap_8 FILLER_8_1163 ();
 sg13g2_fill_2 FILLER_8_1170 ();
 sg13g2_fill_1 FILLER_8_1172 ();
 sg13g2_decap_4 FILLER_8_1181 ();
 sg13g2_fill_2 FILLER_8_1205 ();
 sg13g2_fill_2 FILLER_8_1211 ();
 sg13g2_decap_8 FILLER_8_1230 ();
 sg13g2_fill_2 FILLER_8_1237 ();
 sg13g2_decap_8 FILLER_8_1252 ();
 sg13g2_fill_2 FILLER_8_1259 ();
 sg13g2_decap_8 FILLER_8_1266 ();
 sg13g2_fill_1 FILLER_8_1273 ();
 sg13g2_fill_1 FILLER_8_1292 ();
 sg13g2_decap_8 FILLER_8_1300 ();
 sg13g2_decap_8 FILLER_8_1307 ();
 sg13g2_decap_8 FILLER_8_1314 ();
 sg13g2_decap_4 FILLER_8_1321 ();
 sg13g2_fill_1 FILLER_8_1325 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_24 ();
 sg13g2_decap_8 FILLER_9_31 ();
 sg13g2_decap_4 FILLER_9_38 ();
 sg13g2_decap_8 FILLER_9_47 ();
 sg13g2_decap_4 FILLER_9_54 ();
 sg13g2_fill_1 FILLER_9_58 ();
 sg13g2_decap_8 FILLER_9_62 ();
 sg13g2_decap_4 FILLER_9_69 ();
 sg13g2_fill_2 FILLER_9_76 ();
 sg13g2_fill_1 FILLER_9_92 ();
 sg13g2_fill_2 FILLER_9_99 ();
 sg13g2_fill_1 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_111 ();
 sg13g2_fill_1 FILLER_9_134 ();
 sg13g2_fill_1 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_149 ();
 sg13g2_decap_8 FILLER_9_159 ();
 sg13g2_decap_8 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_173 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_fill_2 FILLER_9_182 ();
 sg13g2_fill_1 FILLER_9_184 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_decap_4 FILLER_9_228 ();
 sg13g2_fill_2 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_246 ();
 sg13g2_fill_1 FILLER_9_253 ();
 sg13g2_fill_2 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_fill_2 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_293 ();
 sg13g2_decap_4 FILLER_9_300 ();
 sg13g2_fill_2 FILLER_9_320 ();
 sg13g2_fill_2 FILLER_9_329 ();
 sg13g2_decap_4 FILLER_9_352 ();
 sg13g2_fill_2 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_4 FILLER_9_370 ();
 sg13g2_fill_1 FILLER_9_374 ();
 sg13g2_fill_1 FILLER_9_378 ();
 sg13g2_fill_1 FILLER_9_401 ();
 sg13g2_fill_2 FILLER_9_418 ();
 sg13g2_fill_2 FILLER_9_431 ();
 sg13g2_fill_1 FILLER_9_433 ();
 sg13g2_decap_8 FILLER_9_464 ();
 sg13g2_fill_2 FILLER_9_489 ();
 sg13g2_fill_2 FILLER_9_496 ();
 sg13g2_fill_1 FILLER_9_498 ();
 sg13g2_decap_8 FILLER_9_544 ();
 sg13g2_decap_8 FILLER_9_551 ();
 sg13g2_fill_1 FILLER_9_558 ();
 sg13g2_fill_1 FILLER_9_574 ();
 sg13g2_fill_2 FILLER_9_578 ();
 sg13g2_fill_1 FILLER_9_580 ();
 sg13g2_fill_1 FILLER_9_586 ();
 sg13g2_fill_1 FILLER_9_597 ();
 sg13g2_fill_2 FILLER_9_602 ();
 sg13g2_fill_2 FILLER_9_609 ();
 sg13g2_fill_1 FILLER_9_611 ();
 sg13g2_decap_4 FILLER_9_625 ();
 sg13g2_fill_2 FILLER_9_629 ();
 sg13g2_fill_2 FILLER_9_639 ();
 sg13g2_fill_1 FILLER_9_641 ();
 sg13g2_fill_1 FILLER_9_650 ();
 sg13g2_fill_1 FILLER_9_658 ();
 sg13g2_decap_4 FILLER_9_669 ();
 sg13g2_fill_2 FILLER_9_673 ();
 sg13g2_fill_2 FILLER_9_679 ();
 sg13g2_decap_4 FILLER_9_685 ();
 sg13g2_decap_4 FILLER_9_765 ();
 sg13g2_fill_2 FILLER_9_774 ();
 sg13g2_decap_4 FILLER_9_789 ();
 sg13g2_fill_1 FILLER_9_823 ();
 sg13g2_fill_1 FILLER_9_833 ();
 sg13g2_fill_1 FILLER_9_845 ();
 sg13g2_fill_1 FILLER_9_852 ();
 sg13g2_fill_2 FILLER_9_857 ();
 sg13g2_fill_1 FILLER_9_864 ();
 sg13g2_decap_4 FILLER_9_894 ();
 sg13g2_fill_2 FILLER_9_903 ();
 sg13g2_fill_1 FILLER_9_905 ();
 sg13g2_decap_4 FILLER_9_922 ();
 sg13g2_decap_8 FILLER_9_956 ();
 sg13g2_decap_4 FILLER_9_963 ();
 sg13g2_fill_2 FILLER_9_976 ();
 sg13g2_fill_1 FILLER_9_978 ();
 sg13g2_decap_8 FILLER_9_983 ();
 sg13g2_fill_1 FILLER_9_990 ();
 sg13g2_fill_2 FILLER_9_996 ();
 sg13g2_decap_8 FILLER_9_1007 ();
 sg13g2_fill_2 FILLER_9_1014 ();
 sg13g2_fill_1 FILLER_9_1016 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_fill_1 FILLER_9_1033 ();
 sg13g2_fill_1 FILLER_9_1038 ();
 sg13g2_fill_2 FILLER_9_1043 ();
 sg13g2_fill_1 FILLER_9_1045 ();
 sg13g2_decap_4 FILLER_9_1057 ();
 sg13g2_fill_2 FILLER_9_1061 ();
 sg13g2_fill_2 FILLER_9_1066 ();
 sg13g2_fill_1 FILLER_9_1068 ();
 sg13g2_decap_4 FILLER_9_1073 ();
 sg13g2_decap_4 FILLER_9_1082 ();
 sg13g2_fill_2 FILLER_9_1086 ();
 sg13g2_fill_2 FILLER_9_1106 ();
 sg13g2_decap_8 FILLER_9_1112 ();
 sg13g2_fill_2 FILLER_9_1119 ();
 sg13g2_fill_1 FILLER_9_1121 ();
 sg13g2_fill_1 FILLER_9_1135 ();
 sg13g2_decap_8 FILLER_9_1143 ();
 sg13g2_decap_4 FILLER_9_1153 ();
 sg13g2_fill_2 FILLER_9_1157 ();
 sg13g2_fill_1 FILLER_9_1169 ();
 sg13g2_decap_8 FILLER_9_1190 ();
 sg13g2_fill_2 FILLER_9_1197 ();
 sg13g2_fill_1 FILLER_9_1199 ();
 sg13g2_fill_1 FILLER_9_1204 ();
 sg13g2_fill_2 FILLER_9_1210 ();
 sg13g2_fill_1 FILLER_9_1212 ();
 sg13g2_fill_2 FILLER_9_1269 ();
 sg13g2_fill_1 FILLER_9_1275 ();
 sg13g2_decap_8 FILLER_9_1299 ();
 sg13g2_decap_8 FILLER_9_1306 ();
 sg13g2_decap_8 FILLER_9_1313 ();
 sg13g2_decap_4 FILLER_9_1320 ();
 sg13g2_fill_2 FILLER_9_1324 ();
 sg13g2_fill_1 FILLER_10_26 ();
 sg13g2_fill_1 FILLER_10_31 ();
 sg13g2_fill_1 FILLER_10_40 ();
 sg13g2_decap_4 FILLER_10_54 ();
 sg13g2_fill_1 FILLER_10_58 ();
 sg13g2_decap_4 FILLER_10_82 ();
 sg13g2_fill_1 FILLER_10_95 ();
 sg13g2_decap_4 FILLER_10_101 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_decap_4 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_fill_2 FILLER_10_167 ();
 sg13g2_decap_4 FILLER_10_250 ();
 sg13g2_fill_2 FILLER_10_254 ();
 sg13g2_decap_4 FILLER_10_264 ();
 sg13g2_fill_1 FILLER_10_268 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_decap_8 FILLER_10_279 ();
 sg13g2_decap_8 FILLER_10_286 ();
 sg13g2_fill_2 FILLER_10_328 ();
 sg13g2_fill_1 FILLER_10_330 ();
 sg13g2_decap_4 FILLER_10_374 ();
 sg13g2_fill_2 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_fill_2 FILLER_10_409 ();
 sg13g2_fill_2 FILLER_10_430 ();
 sg13g2_fill_1 FILLER_10_437 ();
 sg13g2_fill_2 FILLER_10_463 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_4 FILLER_10_483 ();
 sg13g2_fill_1 FILLER_10_495 ();
 sg13g2_fill_2 FILLER_10_501 ();
 sg13g2_fill_1 FILLER_10_516 ();
 sg13g2_fill_1 FILLER_10_522 ();
 sg13g2_fill_2 FILLER_10_527 ();
 sg13g2_fill_2 FILLER_10_533 ();
 sg13g2_fill_1 FILLER_10_535 ();
 sg13g2_decap_8 FILLER_10_544 ();
 sg13g2_decap_8 FILLER_10_551 ();
 sg13g2_fill_2 FILLER_10_558 ();
 sg13g2_fill_1 FILLER_10_560 ();
 sg13g2_fill_1 FILLER_10_564 ();
 sg13g2_fill_2 FILLER_10_579 ();
 sg13g2_fill_2 FILLER_10_587 ();
 sg13g2_fill_2 FILLER_10_593 ();
 sg13g2_fill_1 FILLER_10_595 ();
 sg13g2_fill_1 FILLER_10_601 ();
 sg13g2_fill_2 FILLER_10_608 ();
 sg13g2_decap_8 FILLER_10_613 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_decap_8 FILLER_10_634 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_652 ();
 sg13g2_fill_1 FILLER_10_659 ();
 sg13g2_fill_2 FILLER_10_683 ();
 sg13g2_decap_4 FILLER_10_691 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_fill_1 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_4 FILLER_10_732 ();
 sg13g2_fill_2 FILLER_10_761 ();
 sg13g2_fill_2 FILLER_10_767 ();
 sg13g2_fill_1 FILLER_10_769 ();
 sg13g2_decap_8 FILLER_10_775 ();
 sg13g2_fill_2 FILLER_10_782 ();
 sg13g2_fill_1 FILLER_10_784 ();
 sg13g2_fill_1 FILLER_10_789 ();
 sg13g2_fill_1 FILLER_10_818 ();
 sg13g2_fill_2 FILLER_10_832 ();
 sg13g2_fill_1 FILLER_10_834 ();
 sg13g2_fill_2 FILLER_10_840 ();
 sg13g2_fill_1 FILLER_10_842 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_10_883 ();
 sg13g2_decap_4 FILLER_10_890 ();
 sg13g2_fill_2 FILLER_10_894 ();
 sg13g2_decap_4 FILLER_10_902 ();
 sg13g2_fill_1 FILLER_10_906 ();
 sg13g2_fill_2 FILLER_10_915 ();
 sg13g2_fill_2 FILLER_10_926 ();
 sg13g2_fill_1 FILLER_10_928 ();
 sg13g2_fill_1 FILLER_10_944 ();
 sg13g2_decap_8 FILLER_10_953 ();
 sg13g2_fill_2 FILLER_10_977 ();
 sg13g2_fill_1 FILLER_10_979 ();
 sg13g2_decap_8 FILLER_10_988 ();
 sg13g2_decap_8 FILLER_10_1032 ();
 sg13g2_decap_8 FILLER_10_1039 ();
 sg13g2_decap_4 FILLER_10_1046 ();
 sg13g2_fill_2 FILLER_10_1050 ();
 sg13g2_decap_8 FILLER_10_1057 ();
 sg13g2_fill_1 FILLER_10_1064 ();
 sg13g2_decap_4 FILLER_10_1081 ();
 sg13g2_fill_2 FILLER_10_1085 ();
 sg13g2_fill_1 FILLER_10_1095 ();
 sg13g2_decap_8 FILLER_10_1100 ();
 sg13g2_decap_4 FILLER_10_1107 ();
 sg13g2_decap_8 FILLER_10_1115 ();
 sg13g2_decap_8 FILLER_10_1122 ();
 sg13g2_decap_8 FILLER_10_1129 ();
 sg13g2_decap_8 FILLER_10_1136 ();
 sg13g2_decap_4 FILLER_10_1143 ();
 sg13g2_fill_1 FILLER_10_1147 ();
 sg13g2_fill_1 FILLER_10_1154 ();
 sg13g2_decap_4 FILLER_10_1164 ();
 sg13g2_fill_1 FILLER_10_1168 ();
 sg13g2_fill_1 FILLER_10_1174 ();
 sg13g2_fill_1 FILLER_10_1179 ();
 sg13g2_decap_4 FILLER_10_1193 ();
 sg13g2_fill_1 FILLER_10_1197 ();
 sg13g2_fill_2 FILLER_10_1201 ();
 sg13g2_fill_1 FILLER_10_1203 ();
 sg13g2_fill_2 FILLER_10_1208 ();
 sg13g2_fill_1 FILLER_10_1222 ();
 sg13g2_decap_8 FILLER_10_1242 ();
 sg13g2_decap_8 FILLER_10_1249 ();
 sg13g2_decap_8 FILLER_10_1256 ();
 sg13g2_decap_8 FILLER_10_1263 ();
 sg13g2_decap_8 FILLER_10_1270 ();
 sg13g2_fill_2 FILLER_10_1287 ();
 sg13g2_decap_8 FILLER_10_1293 ();
 sg13g2_decap_8 FILLER_10_1300 ();
 sg13g2_decap_8 FILLER_10_1307 ();
 sg13g2_decap_8 FILLER_10_1314 ();
 sg13g2_decap_4 FILLER_10_1321 ();
 sg13g2_fill_1 FILLER_10_1325 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_4 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_32 ();
 sg13g2_fill_2 FILLER_11_46 ();
 sg13g2_fill_1 FILLER_11_48 ();
 sg13g2_fill_1 FILLER_11_76 ();
 sg13g2_fill_1 FILLER_11_80 ();
 sg13g2_fill_2 FILLER_11_86 ();
 sg13g2_fill_2 FILLER_11_96 ();
 sg13g2_fill_2 FILLER_11_102 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_fill_2 FILLER_11_129 ();
 sg13g2_fill_1 FILLER_11_131 ();
 sg13g2_fill_1 FILLER_11_142 ();
 sg13g2_fill_1 FILLER_11_162 ();
 sg13g2_decap_4 FILLER_11_173 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_fill_1 FILLER_11_191 ();
 sg13g2_fill_1 FILLER_11_197 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_fill_1 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_215 ();
 sg13g2_fill_1 FILLER_11_222 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_235 ();
 sg13g2_fill_1 FILLER_11_237 ();
 sg13g2_decap_4 FILLER_11_242 ();
 sg13g2_fill_1 FILLER_11_246 ();
 sg13g2_decap_4 FILLER_11_259 ();
 sg13g2_fill_1 FILLER_11_296 ();
 sg13g2_fill_2 FILLER_11_330 ();
 sg13g2_fill_1 FILLER_11_337 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_4 FILLER_11_371 ();
 sg13g2_fill_1 FILLER_11_375 ();
 sg13g2_fill_1 FILLER_11_381 ();
 sg13g2_fill_1 FILLER_11_394 ();
 sg13g2_fill_1 FILLER_11_400 ();
 sg13g2_fill_1 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_4 FILLER_11_417 ();
 sg13g2_fill_1 FILLER_11_421 ();
 sg13g2_decap_8 FILLER_11_474 ();
 sg13g2_decap_4 FILLER_11_481 ();
 sg13g2_fill_2 FILLER_11_485 ();
 sg13g2_fill_1 FILLER_11_500 ();
 sg13g2_fill_2 FILLER_11_513 ();
 sg13g2_fill_1 FILLER_11_515 ();
 sg13g2_decap_8 FILLER_11_527 ();
 sg13g2_decap_4 FILLER_11_534 ();
 sg13g2_fill_2 FILLER_11_538 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_4 FILLER_11_567 ();
 sg13g2_fill_1 FILLER_11_571 ();
 sg13g2_decap_4 FILLER_11_593 ();
 sg13g2_fill_1 FILLER_11_597 ();
 sg13g2_decap_4 FILLER_11_621 ();
 sg13g2_fill_1 FILLER_11_625 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_4 FILLER_11_641 ();
 sg13g2_fill_2 FILLER_11_645 ();
 sg13g2_decap_8 FILLER_11_653 ();
 sg13g2_decap_8 FILLER_11_660 ();
 sg13g2_decap_4 FILLER_11_667 ();
 sg13g2_fill_1 FILLER_11_671 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_fill_1 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_decap_4 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_754 ();
 sg13g2_fill_2 FILLER_11_761 ();
 sg13g2_fill_2 FILLER_11_773 ();
 sg13g2_fill_1 FILLER_11_775 ();
 sg13g2_fill_1 FILLER_11_780 ();
 sg13g2_fill_1 FILLER_11_792 ();
 sg13g2_fill_2 FILLER_11_797 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_fill_1 FILLER_11_837 ();
 sg13g2_decap_4 FILLER_11_842 ();
 sg13g2_fill_2 FILLER_11_852 ();
 sg13g2_fill_1 FILLER_11_863 ();
 sg13g2_fill_1 FILLER_11_875 ();
 sg13g2_decap_8 FILLER_11_881 ();
 sg13g2_decap_8 FILLER_11_888 ();
 sg13g2_decap_8 FILLER_11_895 ();
 sg13g2_decap_8 FILLER_11_902 ();
 sg13g2_decap_4 FILLER_11_909 ();
 sg13g2_fill_2 FILLER_11_913 ();
 sg13g2_fill_2 FILLER_11_920 ();
 sg13g2_fill_1 FILLER_11_922 ();
 sg13g2_decap_4 FILLER_11_952 ();
 sg13g2_decap_8 FILLER_11_961 ();
 sg13g2_decap_8 FILLER_11_968 ();
 sg13g2_decap_4 FILLER_11_975 ();
 sg13g2_decap_8 FILLER_11_983 ();
 sg13g2_fill_2 FILLER_11_997 ();
 sg13g2_fill_1 FILLER_11_999 ();
 sg13g2_fill_2 FILLER_11_1005 ();
 sg13g2_fill_1 FILLER_11_1007 ();
 sg13g2_fill_2 FILLER_11_1013 ();
 sg13g2_fill_1 FILLER_11_1015 ();
 sg13g2_decap_8 FILLER_11_1026 ();
 sg13g2_fill_2 FILLER_11_1033 ();
 sg13g2_fill_1 FILLER_11_1035 ();
 sg13g2_fill_2 FILLER_11_1045 ();
 sg13g2_fill_1 FILLER_11_1047 ();
 sg13g2_decap_4 FILLER_11_1051 ();
 sg13g2_fill_1 FILLER_11_1055 ();
 sg13g2_decap_4 FILLER_11_1064 ();
 sg13g2_fill_1 FILLER_11_1068 ();
 sg13g2_decap_4 FILLER_11_1076 ();
 sg13g2_fill_1 FILLER_11_1080 ();
 sg13g2_fill_2 FILLER_11_1085 ();
 sg13g2_fill_1 FILLER_11_1087 ();
 sg13g2_fill_1 FILLER_11_1096 ();
 sg13g2_decap_4 FILLER_11_1102 ();
 sg13g2_fill_2 FILLER_11_1106 ();
 sg13g2_decap_8 FILLER_11_1121 ();
 sg13g2_fill_2 FILLER_11_1128 ();
 sg13g2_fill_1 FILLER_11_1130 ();
 sg13g2_fill_1 FILLER_11_1134 ();
 sg13g2_fill_1 FILLER_11_1147 ();
 sg13g2_fill_2 FILLER_11_1157 ();
 sg13g2_fill_1 FILLER_11_1159 ();
 sg13g2_fill_2 FILLER_11_1164 ();
 sg13g2_fill_1 FILLER_11_1166 ();
 sg13g2_fill_2 FILLER_11_1170 ();
 sg13g2_fill_1 FILLER_11_1176 ();
 sg13g2_fill_1 FILLER_11_1181 ();
 sg13g2_fill_2 FILLER_11_1186 ();
 sg13g2_fill_1 FILLER_11_1194 ();
 sg13g2_fill_2 FILLER_11_1211 ();
 sg13g2_fill_1 FILLER_11_1213 ();
 sg13g2_fill_1 FILLER_11_1219 ();
 sg13g2_decap_8 FILLER_11_1225 ();
 sg13g2_decap_4 FILLER_11_1232 ();
 sg13g2_fill_1 FILLER_11_1240 ();
 sg13g2_fill_1 FILLER_11_1245 ();
 sg13g2_decap_8 FILLER_11_1250 ();
 sg13g2_fill_2 FILLER_11_1261 ();
 sg13g2_fill_1 FILLER_11_1263 ();
 sg13g2_decap_4 FILLER_11_1267 ();
 sg13g2_fill_1 FILLER_11_1280 ();
 sg13g2_fill_1 FILLER_11_1285 ();
 sg13g2_fill_1 FILLER_11_1290 ();
 sg13g2_decap_8 FILLER_11_1296 ();
 sg13g2_decap_8 FILLER_11_1303 ();
 sg13g2_decap_8 FILLER_11_1310 ();
 sg13g2_decap_8 FILLER_11_1317 ();
 sg13g2_fill_2 FILLER_11_1324 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_decap_8 FILLER_12_29 ();
 sg13g2_decap_4 FILLER_12_36 ();
 sg13g2_fill_2 FILLER_12_40 ();
 sg13g2_fill_2 FILLER_12_52 ();
 sg13g2_decap_4 FILLER_12_83 ();
 sg13g2_fill_2 FILLER_12_91 ();
 sg13g2_fill_1 FILLER_12_93 ();
 sg13g2_fill_2 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_decap_8 FILLER_12_122 ();
 sg13g2_fill_2 FILLER_12_129 ();
 sg13g2_decap_8 FILLER_12_136 ();
 sg13g2_decap_8 FILLER_12_143 ();
 sg13g2_decap_8 FILLER_12_150 ();
 sg13g2_decap_8 FILLER_12_157 ();
 sg13g2_decap_4 FILLER_12_164 ();
 sg13g2_fill_1 FILLER_12_168 ();
 sg13g2_fill_1 FILLER_12_179 ();
 sg13g2_fill_2 FILLER_12_183 ();
 sg13g2_fill_2 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_207 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_fill_2 FILLER_12_217 ();
 sg13g2_fill_1 FILLER_12_219 ();
 sg13g2_fill_2 FILLER_12_230 ();
 sg13g2_fill_1 FILLER_12_232 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_241 ();
 sg13g2_fill_2 FILLER_12_248 ();
 sg13g2_decap_4 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_280 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_fill_1 FILLER_12_308 ();
 sg13g2_fill_2 FILLER_12_318 ();
 sg13g2_fill_1 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_4 FILLER_12_364 ();
 sg13g2_fill_1 FILLER_12_373 ();
 sg13g2_fill_1 FILLER_12_383 ();
 sg13g2_fill_1 FILLER_12_389 ();
 sg13g2_fill_2 FILLER_12_396 ();
 sg13g2_fill_1 FILLER_12_410 ();
 sg13g2_decap_8 FILLER_12_418 ();
 sg13g2_decap_4 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_2 FILLER_12_451 ();
 sg13g2_decap_4 FILLER_12_457 ();
 sg13g2_fill_1 FILLER_12_467 ();
 sg13g2_fill_2 FILLER_12_476 ();
 sg13g2_fill_2 FILLER_12_483 ();
 sg13g2_fill_1 FILLER_12_485 ();
 sg13g2_fill_2 FILLER_12_491 ();
 sg13g2_fill_2 FILLER_12_496 ();
 sg13g2_fill_2 FILLER_12_527 ();
 sg13g2_decap_4 FILLER_12_533 ();
 sg13g2_fill_1 FILLER_12_537 ();
 sg13g2_decap_4 FILLER_12_576 ();
 sg13g2_fill_1 FILLER_12_580 ();
 sg13g2_decap_4 FILLER_12_599 ();
 sg13g2_fill_1 FILLER_12_603 ();
 sg13g2_decap_4 FILLER_12_612 ();
 sg13g2_decap_4 FILLER_12_620 ();
 sg13g2_fill_1 FILLER_12_627 ();
 sg13g2_decap_8 FILLER_12_636 ();
 sg13g2_fill_2 FILLER_12_643 ();
 sg13g2_fill_1 FILLER_12_655 ();
 sg13g2_decap_4 FILLER_12_661 ();
 sg13g2_fill_2 FILLER_12_673 ();
 sg13g2_decap_4 FILLER_12_679 ();
 sg13g2_fill_2 FILLER_12_683 ();
 sg13g2_decap_8 FILLER_12_713 ();
 sg13g2_fill_2 FILLER_12_720 ();
 sg13g2_fill_1 FILLER_12_722 ();
 sg13g2_decap_8 FILLER_12_741 ();
 sg13g2_decap_8 FILLER_12_748 ();
 sg13g2_fill_2 FILLER_12_755 ();
 sg13g2_fill_1 FILLER_12_780 ();
 sg13g2_fill_1 FILLER_12_786 ();
 sg13g2_fill_1 FILLER_12_799 ();
 sg13g2_fill_2 FILLER_12_807 ();
 sg13g2_decap_8 FILLER_12_814 ();
 sg13g2_decap_8 FILLER_12_821 ();
 sg13g2_decap_8 FILLER_12_828 ();
 sg13g2_decap_4 FILLER_12_835 ();
 sg13g2_fill_2 FILLER_12_839 ();
 sg13g2_decap_4 FILLER_12_846 ();
 sg13g2_decap_8 FILLER_12_855 ();
 sg13g2_fill_2 FILLER_12_871 ();
 sg13g2_fill_1 FILLER_12_873 ();
 sg13g2_decap_4 FILLER_12_884 ();
 sg13g2_fill_1 FILLER_12_888 ();
 sg13g2_fill_2 FILLER_12_893 ();
 sg13g2_fill_1 FILLER_12_898 ();
 sg13g2_decap_8 FILLER_12_905 ();
 sg13g2_fill_2 FILLER_12_912 ();
 sg13g2_fill_1 FILLER_12_914 ();
 sg13g2_fill_2 FILLER_12_920 ();
 sg13g2_fill_1 FILLER_12_922 ();
 sg13g2_decap_4 FILLER_12_938 ();
 sg13g2_fill_2 FILLER_12_947 ();
 sg13g2_decap_8 FILLER_12_968 ();
 sg13g2_decap_4 FILLER_12_975 ();
 sg13g2_fill_1 FILLER_12_979 ();
 sg13g2_decap_8 FILLER_12_998 ();
 sg13g2_fill_2 FILLER_12_1010 ();
 sg13g2_fill_1 FILLER_12_1012 ();
 sg13g2_decap_4 FILLER_12_1024 ();
 sg13g2_fill_2 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_12_1046 ();
 sg13g2_fill_2 FILLER_12_1053 ();
 sg13g2_fill_1 FILLER_12_1055 ();
 sg13g2_decap_8 FILLER_12_1059 ();
 sg13g2_decap_4 FILLER_12_1066 ();
 sg13g2_fill_2 FILLER_12_1074 ();
 sg13g2_fill_1 FILLER_12_1076 ();
 sg13g2_fill_2 FILLER_12_1091 ();
 sg13g2_fill_1 FILLER_12_1093 ();
 sg13g2_fill_2 FILLER_12_1112 ();
 sg13g2_fill_1 FILLER_12_1114 ();
 sg13g2_fill_2 FILLER_12_1128 ();
 sg13g2_fill_1 FILLER_12_1130 ();
 sg13g2_decap_8 FILLER_12_1134 ();
 sg13g2_fill_1 FILLER_12_1141 ();
 sg13g2_decap_4 FILLER_12_1156 ();
 sg13g2_fill_2 FILLER_12_1160 ();
 sg13g2_fill_1 FILLER_12_1166 ();
 sg13g2_decap_4 FILLER_12_1180 ();
 sg13g2_decap_4 FILLER_12_1192 ();
 sg13g2_fill_2 FILLER_12_1196 ();
 sg13g2_fill_2 FILLER_12_1206 ();
 sg13g2_fill_1 FILLER_12_1208 ();
 sg13g2_fill_1 FILLER_12_1222 ();
 sg13g2_decap_8 FILLER_12_1227 ();
 sg13g2_decap_8 FILLER_12_1234 ();
 sg13g2_decap_4 FILLER_12_1241 ();
 sg13g2_fill_1 FILLER_12_1245 ();
 sg13g2_decap_8 FILLER_12_1255 ();
 sg13g2_decap_4 FILLER_12_1262 ();
 sg13g2_fill_1 FILLER_12_1266 ();
 sg13g2_decap_4 FILLER_12_1273 ();
 sg13g2_decap_4 FILLER_12_1281 ();
 sg13g2_fill_2 FILLER_12_1285 ();
 sg13g2_decap_8 FILLER_12_1295 ();
 sg13g2_decap_8 FILLER_12_1302 ();
 sg13g2_decap_8 FILLER_12_1309 ();
 sg13g2_decap_8 FILLER_12_1316 ();
 sg13g2_fill_2 FILLER_12_1323 ();
 sg13g2_fill_1 FILLER_12_1325 ();
 sg13g2_decap_4 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_15 ();
 sg13g2_decap_8 FILLER_13_22 ();
 sg13g2_fill_2 FILLER_13_29 ();
 sg13g2_decap_4 FILLER_13_36 ();
 sg13g2_fill_2 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_68 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_fill_2 FILLER_13_83 ();
 sg13g2_fill_1 FILLER_13_85 ();
 sg13g2_fill_2 FILLER_13_93 ();
 sg13g2_fill_2 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_101 ();
 sg13g2_fill_1 FILLER_13_131 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_decap_4 FILLER_13_162 ();
 sg13g2_fill_1 FILLER_13_166 ();
 sg13g2_fill_1 FILLER_13_176 ();
 sg13g2_decap_8 FILLER_13_180 ();
 sg13g2_decap_4 FILLER_13_191 ();
 sg13g2_decap_8 FILLER_13_199 ();
 sg13g2_fill_1 FILLER_13_206 ();
 sg13g2_decap_4 FILLER_13_213 ();
 sg13g2_fill_1 FILLER_13_217 ();
 sg13g2_decap_4 FILLER_13_234 ();
 sg13g2_fill_1 FILLER_13_238 ();
 sg13g2_fill_2 FILLER_13_244 ();
 sg13g2_decap_8 FILLER_13_250 ();
 sg13g2_fill_2 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_263 ();
 sg13g2_decap_4 FILLER_13_287 ();
 sg13g2_fill_2 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_300 ();
 sg13g2_decap_4 FILLER_13_307 ();
 sg13g2_fill_2 FILLER_13_311 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_fill_1 FILLER_13_332 ();
 sg13g2_fill_1 FILLER_13_337 ();
 sg13g2_fill_2 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_fill_1 FILLER_13_360 ();
 sg13g2_fill_2 FILLER_13_380 ();
 sg13g2_fill_2 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_411 ();
 sg13g2_decap_4 FILLER_13_421 ();
 sg13g2_fill_1 FILLER_13_425 ();
 sg13g2_decap_4 FILLER_13_441 ();
 sg13g2_decap_4 FILLER_13_476 ();
 sg13g2_fill_1 FILLER_13_485 ();
 sg13g2_fill_2 FILLER_13_491 ();
 sg13g2_decap_8 FILLER_13_540 ();
 sg13g2_fill_2 FILLER_13_547 ();
 sg13g2_fill_1 FILLER_13_549 ();
 sg13g2_decap_4 FILLER_13_558 ();
 sg13g2_fill_1 FILLER_13_562 ();
 sg13g2_fill_2 FILLER_13_567 ();
 sg13g2_fill_1 FILLER_13_569 ();
 sg13g2_fill_2 FILLER_13_590 ();
 sg13g2_fill_1 FILLER_13_601 ();
 sg13g2_decap_8 FILLER_13_607 ();
 sg13g2_fill_1 FILLER_13_614 ();
 sg13g2_fill_2 FILLER_13_654 ();
 sg13g2_decap_4 FILLER_13_663 ();
 sg13g2_fill_2 FILLER_13_667 ();
 sg13g2_fill_2 FILLER_13_681 ();
 sg13g2_fill_1 FILLER_13_683 ();
 sg13g2_fill_1 FILLER_13_697 ();
 sg13g2_decap_8 FILLER_13_708 ();
 sg13g2_decap_8 FILLER_13_715 ();
 sg13g2_fill_1 FILLER_13_722 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_fill_2 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_769 ();
 sg13g2_decap_8 FILLER_13_776 ();
 sg13g2_decap_8 FILLER_13_783 ();
 sg13g2_decap_8 FILLER_13_790 ();
 sg13g2_decap_8 FILLER_13_797 ();
 sg13g2_decap_8 FILLER_13_804 ();
 sg13g2_fill_2 FILLER_13_811 ();
 sg13g2_decap_4 FILLER_13_835 ();
 sg13g2_fill_1 FILLER_13_839 ();
 sg13g2_decap_4 FILLER_13_852 ();
 sg13g2_decap_8 FILLER_13_860 ();
 sg13g2_decap_4 FILLER_13_867 ();
 sg13g2_fill_2 FILLER_13_899 ();
 sg13g2_decap_8 FILLER_13_908 ();
 sg13g2_decap_8 FILLER_13_915 ();
 sg13g2_fill_1 FILLER_13_922 ();
 sg13g2_fill_2 FILLER_13_934 ();
 sg13g2_fill_1 FILLER_13_950 ();
 sg13g2_decap_4 FILLER_13_954 ();
 sg13g2_fill_2 FILLER_13_966 ();
 sg13g2_fill_1 FILLER_13_968 ();
 sg13g2_decap_8 FILLER_13_974 ();
 sg13g2_decap_8 FILLER_13_981 ();
 sg13g2_decap_8 FILLER_13_988 ();
 sg13g2_fill_1 FILLER_13_995 ();
 sg13g2_fill_2 FILLER_13_1001 ();
 sg13g2_decap_4 FILLER_13_1007 ();
 sg13g2_fill_1 FILLER_13_1011 ();
 sg13g2_fill_2 FILLER_13_1017 ();
 sg13g2_fill_1 FILLER_13_1019 ();
 sg13g2_decap_8 FILLER_13_1023 ();
 sg13g2_fill_2 FILLER_13_1030 ();
 sg13g2_fill_1 FILLER_13_1032 ();
 sg13g2_fill_2 FILLER_13_1038 ();
 sg13g2_decap_4 FILLER_13_1044 ();
 sg13g2_decap_4 FILLER_13_1052 ();
 sg13g2_fill_1 FILLER_13_1072 ();
 sg13g2_fill_2 FILLER_13_1088 ();
 sg13g2_fill_1 FILLER_13_1090 ();
 sg13g2_decap_4 FILLER_13_1096 ();
 sg13g2_fill_1 FILLER_13_1100 ();
 sg13g2_fill_2 FILLER_13_1106 ();
 sg13g2_fill_1 FILLER_13_1114 ();
 sg13g2_decap_4 FILLER_13_1118 ();
 sg13g2_fill_2 FILLER_13_1131 ();
 sg13g2_fill_1 FILLER_13_1133 ();
 sg13g2_fill_1 FILLER_13_1143 ();
 sg13g2_fill_2 FILLER_13_1151 ();
 sg13g2_fill_1 FILLER_13_1186 ();
 sg13g2_decap_8 FILLER_13_1191 ();
 sg13g2_decap_8 FILLER_13_1201 ();
 sg13g2_fill_2 FILLER_13_1208 ();
 sg13g2_fill_1 FILLER_13_1216 ();
 sg13g2_fill_1 FILLER_13_1222 ();
 sg13g2_decap_4 FILLER_13_1228 ();
 sg13g2_fill_2 FILLER_13_1253 ();
 sg13g2_fill_1 FILLER_13_1255 ();
 sg13g2_fill_1 FILLER_13_1280 ();
 sg13g2_fill_1 FILLER_13_1297 ();
 sg13g2_decap_8 FILLER_13_1310 ();
 sg13g2_decap_8 FILLER_13_1317 ();
 sg13g2_fill_2 FILLER_13_1324 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_43 ();
 sg13g2_fill_1 FILLER_14_45 ();
 sg13g2_decap_8 FILLER_14_50 ();
 sg13g2_decap_8 FILLER_14_57 ();
 sg13g2_fill_1 FILLER_14_64 ();
 sg13g2_fill_1 FILLER_14_69 ();
 sg13g2_fill_2 FILLER_14_75 ();
 sg13g2_fill_1 FILLER_14_77 ();
 sg13g2_fill_2 FILLER_14_82 ();
 sg13g2_decap_8 FILLER_14_87 ();
 sg13g2_decap_4 FILLER_14_94 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_115 ();
 sg13g2_fill_1 FILLER_14_121 ();
 sg13g2_fill_2 FILLER_14_131 ();
 sg13g2_fill_1 FILLER_14_141 ();
 sg13g2_decap_8 FILLER_14_169 ();
 sg13g2_fill_2 FILLER_14_176 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_fill_2 FILLER_14_204 ();
 sg13g2_fill_1 FILLER_14_206 ();
 sg13g2_decap_8 FILLER_14_244 ();
 sg13g2_fill_2 FILLER_14_263 ();
 sg13g2_fill_1 FILLER_14_265 ();
 sg13g2_fill_1 FILLER_14_270 ();
 sg13g2_fill_1 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_4 FILLER_14_308 ();
 sg13g2_fill_2 FILLER_14_312 ();
 sg13g2_fill_2 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_332 ();
 sg13g2_decap_8 FILLER_14_339 ();
 sg13g2_decap_4 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_350 ();
 sg13g2_fill_2 FILLER_14_356 ();
 sg13g2_fill_1 FILLER_14_358 ();
 sg13g2_fill_2 FILLER_14_370 ();
 sg13g2_fill_1 FILLER_14_372 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_decap_4 FILLER_14_381 ();
 sg13g2_fill_1 FILLER_14_385 ();
 sg13g2_decap_4 FILLER_14_391 ();
 sg13g2_fill_2 FILLER_14_398 ();
 sg13g2_fill_2 FILLER_14_421 ();
 sg13g2_fill_1 FILLER_14_423 ();
 sg13g2_fill_1 FILLER_14_442 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_4 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_470 ();
 sg13g2_fill_1 FILLER_14_477 ();
 sg13g2_fill_1 FILLER_14_496 ();
 sg13g2_decap_8 FILLER_14_522 ();
 sg13g2_decap_4 FILLER_14_529 ();
 sg13g2_decap_8 FILLER_14_558 ();
 sg13g2_fill_2 FILLER_14_565 ();
 sg13g2_fill_1 FILLER_14_567 ();
 sg13g2_fill_1 FILLER_14_573 ();
 sg13g2_fill_1 FILLER_14_580 ();
 sg13g2_fill_2 FILLER_14_585 ();
 sg13g2_fill_1 FILLER_14_592 ();
 sg13g2_fill_2 FILLER_14_596 ();
 sg13g2_fill_2 FILLER_14_627 ();
 sg13g2_fill_2 FILLER_14_639 ();
 sg13g2_fill_1 FILLER_14_646 ();
 sg13g2_decap_8 FILLER_14_653 ();
 sg13g2_fill_2 FILLER_14_660 ();
 sg13g2_fill_1 FILLER_14_662 ();
 sg13g2_fill_2 FILLER_14_666 ();
 sg13g2_decap_4 FILLER_14_672 ();
 sg13g2_decap_4 FILLER_14_683 ();
 sg13g2_fill_1 FILLER_14_696 ();
 sg13g2_decap_4 FILLER_14_735 ();
 sg13g2_fill_2 FILLER_14_747 ();
 sg13g2_fill_2 FILLER_14_752 ();
 sg13g2_fill_2 FILLER_14_772 ();
 sg13g2_fill_2 FILLER_14_778 ();
 sg13g2_fill_1 FILLER_14_780 ();
 sg13g2_fill_2 FILLER_14_786 ();
 sg13g2_fill_1 FILLER_14_788 ();
 sg13g2_decap_4 FILLER_14_795 ();
 sg13g2_fill_1 FILLER_14_799 ();
 sg13g2_fill_2 FILLER_14_805 ();
 sg13g2_fill_1 FILLER_14_807 ();
 sg13g2_fill_1 FILLER_14_830 ();
 sg13g2_decap_4 FILLER_14_836 ();
 sg13g2_fill_1 FILLER_14_840 ();
 sg13g2_fill_2 FILLER_14_849 ();
 sg13g2_decap_8 FILLER_14_861 ();
 sg13g2_fill_2 FILLER_14_872 ();
 sg13g2_decap_8 FILLER_14_887 ();
 sg13g2_fill_1 FILLER_14_894 ();
 sg13g2_decap_8 FILLER_14_903 ();
 sg13g2_decap_4 FILLER_14_910 ();
 sg13g2_fill_2 FILLER_14_914 ();
 sg13g2_fill_1 FILLER_14_919 ();
 sg13g2_decap_4 FILLER_14_925 ();
 sg13g2_fill_1 FILLER_14_929 ();
 sg13g2_decap_8 FILLER_14_944 ();
 sg13g2_decap_4 FILLER_14_951 ();
 sg13g2_fill_2 FILLER_14_963 ();
 sg13g2_fill_2 FILLER_14_998 ();
 sg13g2_fill_1 FILLER_14_1009 ();
 sg13g2_fill_2 FILLER_14_1014 ();
 sg13g2_decap_8 FILLER_14_1026 ();
 sg13g2_decap_8 FILLER_14_1046 ();
 sg13g2_decap_8 FILLER_14_1053 ();
 sg13g2_decap_8 FILLER_14_1069 ();
 sg13g2_fill_1 FILLER_14_1081 ();
 sg13g2_fill_1 FILLER_14_1090 ();
 sg13g2_decap_4 FILLER_14_1095 ();
 sg13g2_fill_1 FILLER_14_1099 ();
 sg13g2_decap_8 FILLER_14_1135 ();
 sg13g2_fill_1 FILLER_14_1147 ();
 sg13g2_decap_4 FILLER_14_1152 ();
 sg13g2_fill_2 FILLER_14_1156 ();
 sg13g2_fill_1 FILLER_14_1166 ();
 sg13g2_fill_1 FILLER_14_1174 ();
 sg13g2_fill_1 FILLER_14_1180 ();
 sg13g2_fill_1 FILLER_14_1227 ();
 sg13g2_decap_4 FILLER_14_1247 ();
 sg13g2_fill_1 FILLER_14_1251 ();
 sg13g2_decap_4 FILLER_14_1261 ();
 sg13g2_fill_1 FILLER_14_1265 ();
 sg13g2_fill_2 FILLER_14_1270 ();
 sg13g2_decap_4 FILLER_14_1284 ();
 sg13g2_fill_1 FILLER_14_1288 ();
 sg13g2_fill_2 FILLER_14_1294 ();
 sg13g2_fill_1 FILLER_14_1296 ();
 sg13g2_decap_8 FILLER_14_1302 ();
 sg13g2_decap_8 FILLER_14_1309 ();
 sg13g2_decap_8 FILLER_14_1316 ();
 sg13g2_fill_2 FILLER_14_1323 ();
 sg13g2_fill_1 FILLER_14_1325 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_41 ();
 sg13g2_fill_1 FILLER_15_48 ();
 sg13g2_fill_1 FILLER_15_53 ();
 sg13g2_fill_2 FILLER_15_62 ();
 sg13g2_fill_1 FILLER_15_72 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_1 FILLER_15_88 ();
 sg13g2_decap_8 FILLER_15_99 ();
 sg13g2_decap_4 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_110 ();
 sg13g2_fill_2 FILLER_15_148 ();
 sg13g2_fill_2 FILLER_15_160 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_171 ();
 sg13g2_decap_8 FILLER_15_181 ();
 sg13g2_fill_1 FILLER_15_197 ();
 sg13g2_fill_1 FILLER_15_202 ();
 sg13g2_decap_8 FILLER_15_219 ();
 sg13g2_fill_1 FILLER_15_226 ();
 sg13g2_fill_2 FILLER_15_233 ();
 sg13g2_fill_1 FILLER_15_240 ();
 sg13g2_fill_2 FILLER_15_244 ();
 sg13g2_decap_8 FILLER_15_264 ();
 sg13g2_decap_8 FILLER_15_271 ();
 sg13g2_decap_4 FILLER_15_278 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_decap_4 FILLER_15_292 ();
 sg13g2_fill_2 FILLER_15_296 ();
 sg13g2_decap_4 FILLER_15_310 ();
 sg13g2_fill_2 FILLER_15_314 ();
 sg13g2_fill_2 FILLER_15_331 ();
 sg13g2_fill_1 FILLER_15_333 ();
 sg13g2_decap_4 FILLER_15_340 ();
 sg13g2_fill_1 FILLER_15_344 ();
 sg13g2_decap_4 FILLER_15_352 ();
 sg13g2_fill_2 FILLER_15_356 ();
 sg13g2_decap_4 FILLER_15_362 ();
 sg13g2_fill_2 FILLER_15_366 ();
 sg13g2_fill_1 FILLER_15_373 ();
 sg13g2_decap_4 FILLER_15_392 ();
 sg13g2_fill_2 FILLER_15_409 ();
 sg13g2_fill_2 FILLER_15_416 ();
 sg13g2_fill_1 FILLER_15_418 ();
 sg13g2_fill_1 FILLER_15_428 ();
 sg13g2_fill_2 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_446 ();
 sg13g2_decap_8 FILLER_15_453 ();
 sg13g2_fill_2 FILLER_15_460 ();
 sg13g2_fill_1 FILLER_15_462 ();
 sg13g2_fill_1 FILLER_15_467 ();
 sg13g2_fill_2 FILLER_15_484 ();
 sg13g2_fill_2 FILLER_15_494 ();
 sg13g2_decap_4 FILLER_15_500 ();
 sg13g2_decap_8 FILLER_15_516 ();
 sg13g2_fill_1 FILLER_15_523 ();
 sg13g2_decap_4 FILLER_15_532 ();
 sg13g2_fill_2 FILLER_15_536 ();
 sg13g2_decap_4 FILLER_15_542 ();
 sg13g2_fill_1 FILLER_15_546 ();
 sg13g2_fill_2 FILLER_15_554 ();
 sg13g2_fill_1 FILLER_15_556 ();
 sg13g2_decap_8 FILLER_15_562 ();
 sg13g2_fill_2 FILLER_15_569 ();
 sg13g2_fill_1 FILLER_15_571 ();
 sg13g2_decap_8 FILLER_15_578 ();
 sg13g2_fill_1 FILLER_15_585 ();
 sg13g2_fill_1 FILLER_15_590 ();
 sg13g2_fill_2 FILLER_15_603 ();
 sg13g2_fill_1 FILLER_15_605 ();
 sg13g2_decap_4 FILLER_15_611 ();
 sg13g2_fill_1 FILLER_15_615 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_4 FILLER_15_637 ();
 sg13g2_fill_1 FILLER_15_641 ();
 sg13g2_decap_4 FILLER_15_658 ();
 sg13g2_fill_1 FILLER_15_662 ();
 sg13g2_fill_2 FILLER_15_667 ();
 sg13g2_fill_1 FILLER_15_669 ();
 sg13g2_decap_4 FILLER_15_675 ();
 sg13g2_fill_2 FILLER_15_693 ();
 sg13g2_decap_4 FILLER_15_713 ();
 sg13g2_fill_2 FILLER_15_717 ();
 sg13g2_fill_1 FILLER_15_725 ();
 sg13g2_fill_1 FILLER_15_742 ();
 sg13g2_fill_1 FILLER_15_765 ();
 sg13g2_fill_2 FILLER_15_778 ();
 sg13g2_decap_4 FILLER_15_786 ();
 sg13g2_fill_1 FILLER_15_790 ();
 sg13g2_fill_2 FILLER_15_796 ();
 sg13g2_fill_1 FILLER_15_798 ();
 sg13g2_fill_2 FILLER_15_811 ();
 sg13g2_fill_1 FILLER_15_813 ();
 sg13g2_fill_1 FILLER_15_840 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_4 FILLER_15_888 ();
 sg13g2_fill_2 FILLER_15_892 ();
 sg13g2_decap_4 FILLER_15_902 ();
 sg13g2_decap_4 FILLER_15_910 ();
 sg13g2_fill_2 FILLER_15_914 ();
 sg13g2_fill_2 FILLER_15_921 ();
 sg13g2_decap_4 FILLER_15_933 ();
 sg13g2_decap_8 FILLER_15_947 ();
 sg13g2_decap_8 FILLER_15_962 ();
 sg13g2_decap_4 FILLER_15_969 ();
 sg13g2_fill_2 FILLER_15_978 ();
 sg13g2_fill_2 FILLER_15_983 ();
 sg13g2_fill_1 FILLER_15_985 ();
 sg13g2_decap_4 FILLER_15_994 ();
 sg13g2_fill_1 FILLER_15_998 ();
 sg13g2_fill_1 FILLER_15_1006 ();
 sg13g2_decap_4 FILLER_15_1015 ();
 sg13g2_decap_8 FILLER_15_1025 ();
 sg13g2_fill_2 FILLER_15_1032 ();
 sg13g2_decap_4 FILLER_15_1043 ();
 sg13g2_fill_1 FILLER_15_1072 ();
 sg13g2_decap_8 FILLER_15_1093 ();
 sg13g2_decap_8 FILLER_15_1104 ();
 sg13g2_fill_2 FILLER_15_1111 ();
 sg13g2_decap_8 FILLER_15_1120 ();
 sg13g2_decap_8 FILLER_15_1127 ();
 sg13g2_decap_8 FILLER_15_1134 ();
 sg13g2_fill_1 FILLER_15_1141 ();
 sg13g2_fill_1 FILLER_15_1150 ();
 sg13g2_fill_1 FILLER_15_1156 ();
 sg13g2_decap_8 FILLER_15_1172 ();
 sg13g2_decap_4 FILLER_15_1179 ();
 sg13g2_fill_2 FILLER_15_1183 ();
 sg13g2_fill_2 FILLER_15_1189 ();
 sg13g2_fill_1 FILLER_15_1191 ();
 sg13g2_fill_1 FILLER_15_1196 ();
 sg13g2_fill_1 FILLER_15_1240 ();
 sg13g2_decap_8 FILLER_15_1249 ();
 sg13g2_decap_8 FILLER_15_1256 ();
 sg13g2_fill_2 FILLER_15_1263 ();
 sg13g2_fill_1 FILLER_15_1265 ();
 sg13g2_decap_8 FILLER_15_1274 ();
 sg13g2_decap_4 FILLER_15_1281 ();
 sg13g2_fill_2 FILLER_15_1285 ();
 sg13g2_decap_8 FILLER_15_1317 ();
 sg13g2_fill_2 FILLER_15_1324 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_4 FILLER_16_14 ();
 sg13g2_decap_4 FILLER_16_30 ();
 sg13g2_fill_1 FILLER_16_34 ();
 sg13g2_decap_8 FILLER_16_40 ();
 sg13g2_fill_2 FILLER_16_47 ();
 sg13g2_fill_2 FILLER_16_62 ();
 sg13g2_fill_1 FILLER_16_64 ();
 sg13g2_fill_1 FILLER_16_71 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_fill_1 FILLER_16_95 ();
 sg13g2_fill_1 FILLER_16_127 ();
 sg13g2_fill_1 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_1 FILLER_16_161 ();
 sg13g2_fill_1 FILLER_16_167 ();
 sg13g2_decap_4 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_fill_2 FILLER_16_198 ();
 sg13g2_decap_4 FILLER_16_209 ();
 sg13g2_fill_2 FILLER_16_213 ();
 sg13g2_decap_4 FILLER_16_220 ();
 sg13g2_fill_1 FILLER_16_233 ();
 sg13g2_fill_2 FILLER_16_243 ();
 sg13g2_fill_1 FILLER_16_259 ();
 sg13g2_fill_1 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_fill_2 FILLER_16_304 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_fill_2 FILLER_16_317 ();
 sg13g2_fill_2 FILLER_16_324 ();
 sg13g2_fill_2 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_decap_4 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_390 ();
 sg13g2_fill_2 FILLER_16_397 ();
 sg13g2_fill_1 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_434 ();
 sg13g2_fill_1 FILLER_16_442 ();
 sg13g2_decap_4 FILLER_16_447 ();
 sg13g2_fill_2 FILLER_16_451 ();
 sg13g2_fill_2 FILLER_16_459 ();
 sg13g2_fill_1 FILLER_16_461 ();
 sg13g2_fill_1 FILLER_16_470 ();
 sg13g2_fill_2 FILLER_16_484 ();
 sg13g2_fill_1 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_495 ();
 sg13g2_decap_8 FILLER_16_502 ();
 sg13g2_decap_8 FILLER_16_509 ();
 sg13g2_decap_4 FILLER_16_516 ();
 sg13g2_fill_2 FILLER_16_523 ();
 sg13g2_fill_1 FILLER_16_525 ();
 sg13g2_fill_1 FILLER_16_529 ();
 sg13g2_fill_1 FILLER_16_549 ();
 sg13g2_fill_2 FILLER_16_564 ();
 sg13g2_decap_8 FILLER_16_570 ();
 sg13g2_decap_8 FILLER_16_577 ();
 sg13g2_decap_4 FILLER_16_584 ();
 sg13g2_fill_1 FILLER_16_592 ();
 sg13g2_decap_4 FILLER_16_598 ();
 sg13g2_fill_2 FILLER_16_607 ();
 sg13g2_decap_4 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_624 ();
 sg13g2_decap_4 FILLER_16_631 ();
 sg13g2_fill_2 FILLER_16_640 ();
 sg13g2_fill_1 FILLER_16_642 ();
 sg13g2_fill_2 FILLER_16_651 ();
 sg13g2_fill_1 FILLER_16_653 ();
 sg13g2_fill_1 FILLER_16_659 ();
 sg13g2_fill_1 FILLER_16_673 ();
 sg13g2_decap_4 FILLER_16_683 ();
 sg13g2_fill_2 FILLER_16_693 ();
 sg13g2_fill_1 FILLER_16_695 ();
 sg13g2_fill_1 FILLER_16_701 ();
 sg13g2_fill_1 FILLER_16_706 ();
 sg13g2_fill_1 FILLER_16_711 ();
 sg13g2_fill_1 FILLER_16_769 ();
 sg13g2_fill_1 FILLER_16_801 ();
 sg13g2_fill_2 FILLER_16_808 ();
 sg13g2_fill_2 FILLER_16_820 ();
 sg13g2_decap_4 FILLER_16_825 ();
 sg13g2_fill_2 FILLER_16_829 ();
 sg13g2_fill_2 FILLER_16_843 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_866 ();
 sg13g2_fill_2 FILLER_16_883 ();
 sg13g2_decap_4 FILLER_16_889 ();
 sg13g2_fill_2 FILLER_16_893 ();
 sg13g2_fill_2 FILLER_16_912 ();
 sg13g2_fill_1 FILLER_16_914 ();
 sg13g2_decap_8 FILLER_16_919 ();
 sg13g2_decap_8 FILLER_16_926 ();
 sg13g2_decap_4 FILLER_16_933 ();
 sg13g2_fill_2 FILLER_16_937 ();
 sg13g2_decap_8 FILLER_16_962 ();
 sg13g2_decap_4 FILLER_16_969 ();
 sg13g2_fill_1 FILLER_16_973 ();
 sg13g2_fill_1 FILLER_16_987 ();
 sg13g2_decap_8 FILLER_16_998 ();
 sg13g2_fill_2 FILLER_16_1009 ();
 sg13g2_fill_1 FILLER_16_1011 ();
 sg13g2_fill_1 FILLER_16_1015 ();
 sg13g2_fill_1 FILLER_16_1020 ();
 sg13g2_fill_2 FILLER_16_1025 ();
 sg13g2_fill_1 FILLER_16_1027 ();
 sg13g2_fill_2 FILLER_16_1036 ();
 sg13g2_fill_1 FILLER_16_1038 ();
 sg13g2_decap_8 FILLER_16_1043 ();
 sg13g2_fill_2 FILLER_16_1050 ();
 sg13g2_decap_8 FILLER_16_1061 ();
 sg13g2_decap_8 FILLER_16_1081 ();
 sg13g2_decap_4 FILLER_16_1088 ();
 sg13g2_fill_1 FILLER_16_1092 ();
 sg13g2_fill_2 FILLER_16_1106 ();
 sg13g2_fill_1 FILLER_16_1108 ();
 sg13g2_decap_4 FILLER_16_1118 ();
 sg13g2_fill_1 FILLER_16_1134 ();
 sg13g2_decap_8 FILLER_16_1141 ();
 sg13g2_fill_1 FILLER_16_1160 ();
 sg13g2_fill_1 FILLER_16_1165 ();
 sg13g2_fill_2 FILLER_16_1171 ();
 sg13g2_fill_2 FILLER_16_1181 ();
 sg13g2_fill_1 FILLER_16_1188 ();
 sg13g2_fill_1 FILLER_16_1213 ();
 sg13g2_fill_1 FILLER_16_1217 ();
 sg13g2_fill_2 FILLER_16_1267 ();
 sg13g2_fill_1 FILLER_16_1274 ();
 sg13g2_fill_1 FILLER_16_1283 ();
 sg13g2_decap_8 FILLER_16_1287 ();
 sg13g2_decap_4 FILLER_16_1294 ();
 sg13g2_decap_8 FILLER_16_1312 ();
 sg13g2_decap_8 FILLER_16_1319 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_decap_4 FILLER_17_11 ();
 sg13g2_fill_2 FILLER_17_15 ();
 sg13g2_decap_4 FILLER_17_55 ();
 sg13g2_fill_1 FILLER_17_59 ();
 sg13g2_fill_2 FILLER_17_86 ();
 sg13g2_fill_1 FILLER_17_103 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_decap_4 FILLER_17_116 ();
 sg13g2_decap_4 FILLER_17_139 ();
 sg13g2_fill_1 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_174 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_206 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_decap_4 FILLER_17_246 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_decap_4 FILLER_17_269 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_292 ();
 sg13g2_decap_8 FILLER_17_304 ();
 sg13g2_fill_1 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_fill_2 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_fill_1 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_fill_2 FILLER_17_363 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_fill_2 FILLER_17_376 ();
 sg13g2_decap_4 FILLER_17_400 ();
 sg13g2_decap_8 FILLER_17_409 ();
 sg13g2_decap_4 FILLER_17_416 ();
 sg13g2_fill_1 FILLER_17_420 ();
 sg13g2_fill_1 FILLER_17_424 ();
 sg13g2_decap_4 FILLER_17_433 ();
 sg13g2_decap_8 FILLER_17_449 ();
 sg13g2_decap_4 FILLER_17_456 ();
 sg13g2_fill_2 FILLER_17_473 ();
 sg13g2_decap_8 FILLER_17_495 ();
 sg13g2_fill_2 FILLER_17_502 ();
 sg13g2_fill_1 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_508 ();
 sg13g2_decap_8 FILLER_17_515 ();
 sg13g2_decap_8 FILLER_17_522 ();
 sg13g2_fill_2 FILLER_17_529 ();
 sg13g2_fill_1 FILLER_17_531 ();
 sg13g2_fill_2 FILLER_17_537 ();
 sg13g2_fill_1 FILLER_17_543 ();
 sg13g2_fill_2 FILLER_17_552 ();
 sg13g2_fill_1 FILLER_17_554 ();
 sg13g2_fill_1 FILLER_17_573 ();
 sg13g2_fill_2 FILLER_17_578 ();
 sg13g2_fill_1 FILLER_17_580 ();
 sg13g2_decap_8 FILLER_17_586 ();
 sg13g2_fill_2 FILLER_17_593 ();
 sg13g2_decap_8 FILLER_17_600 ();
 sg13g2_decap_8 FILLER_17_607 ();
 sg13g2_decap_8 FILLER_17_614 ();
 sg13g2_decap_8 FILLER_17_625 ();
 sg13g2_decap_4 FILLER_17_643 ();
 sg13g2_fill_1 FILLER_17_651 ();
 sg13g2_fill_1 FILLER_17_658 ();
 sg13g2_fill_1 FILLER_17_669 ();
 sg13g2_fill_2 FILLER_17_673 ();
 sg13g2_fill_1 FILLER_17_685 ();
 sg13g2_decap_8 FILLER_17_694 ();
 sg13g2_decap_8 FILLER_17_701 ();
 sg13g2_decap_8 FILLER_17_708 ();
 sg13g2_fill_2 FILLER_17_715 ();
 sg13g2_fill_1 FILLER_17_717 ();
 sg13g2_decap_4 FILLER_17_722 ();
 sg13g2_fill_1 FILLER_17_730 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_fill_2 FILLER_17_749 ();
 sg13g2_fill_1 FILLER_17_751 ();
 sg13g2_decap_8 FILLER_17_757 ();
 sg13g2_decap_4 FILLER_17_771 ();
 sg13g2_fill_1 FILLER_17_775 ();
 sg13g2_fill_2 FILLER_17_780 ();
 sg13g2_fill_2 FILLER_17_791 ();
 sg13g2_fill_2 FILLER_17_802 ();
 sg13g2_fill_1 FILLER_17_814 ();
 sg13g2_fill_2 FILLER_17_819 ();
 sg13g2_fill_1 FILLER_17_825 ();
 sg13g2_fill_1 FILLER_17_836 ();
 sg13g2_fill_2 FILLER_17_846 ();
 sg13g2_fill_1 FILLER_17_853 ();
 sg13g2_fill_1 FILLER_17_865 ();
 sg13g2_fill_2 FILLER_17_871 ();
 sg13g2_decap_8 FILLER_17_878 ();
 sg13g2_fill_1 FILLER_17_885 ();
 sg13g2_decap_4 FILLER_17_890 ();
 sg13g2_fill_1 FILLER_17_894 ();
 sg13g2_decap_8 FILLER_17_898 ();
 sg13g2_decap_8 FILLER_17_905 ();
 sg13g2_decap_4 FILLER_17_912 ();
 sg13g2_decap_8 FILLER_17_925 ();
 sg13g2_decap_8 FILLER_17_932 ();
 sg13g2_decap_8 FILLER_17_943 ();
 sg13g2_fill_1 FILLER_17_950 ();
 sg13g2_fill_2 FILLER_17_969 ();
 sg13g2_fill_1 FILLER_17_976 ();
 sg13g2_fill_1 FILLER_17_981 ();
 sg13g2_fill_1 FILLER_17_987 ();
 sg13g2_decap_8 FILLER_17_993 ();
 sg13g2_decap_4 FILLER_17_1000 ();
 sg13g2_fill_2 FILLER_17_1008 ();
 sg13g2_fill_1 FILLER_17_1010 ();
 sg13g2_fill_2 FILLER_17_1019 ();
 sg13g2_decap_8 FILLER_17_1025 ();
 sg13g2_fill_2 FILLER_17_1032 ();
 sg13g2_fill_1 FILLER_17_1046 ();
 sg13g2_fill_2 FILLER_17_1054 ();
 sg13g2_fill_1 FILLER_17_1056 ();
 sg13g2_decap_8 FILLER_17_1065 ();
 sg13g2_decap_8 FILLER_17_1072 ();
 sg13g2_decap_8 FILLER_17_1079 ();
 sg13g2_fill_1 FILLER_17_1086 ();
 sg13g2_decap_8 FILLER_17_1090 ();
 sg13g2_decap_8 FILLER_17_1097 ();
 sg13g2_fill_2 FILLER_17_1104 ();
 sg13g2_fill_1 FILLER_17_1106 ();
 sg13g2_fill_1 FILLER_17_1116 ();
 sg13g2_fill_1 FILLER_17_1126 ();
 sg13g2_decap_8 FILLER_17_1134 ();
 sg13g2_decap_8 FILLER_17_1141 ();
 sg13g2_decap_8 FILLER_17_1148 ();
 sg13g2_decap_4 FILLER_17_1155 ();
 sg13g2_fill_1 FILLER_17_1159 ();
 sg13g2_decap_4 FILLER_17_1169 ();
 sg13g2_fill_1 FILLER_17_1173 ();
 sg13g2_decap_8 FILLER_17_1185 ();
 sg13g2_fill_2 FILLER_17_1192 ();
 sg13g2_fill_1 FILLER_17_1194 ();
 sg13g2_fill_1 FILLER_17_1225 ();
 sg13g2_decap_8 FILLER_17_1251 ();
 sg13g2_decap_8 FILLER_17_1258 ();
 sg13g2_decap_8 FILLER_17_1265 ();
 sg13g2_decap_8 FILLER_17_1272 ();
 sg13g2_decap_8 FILLER_17_1279 ();
 sg13g2_decap_8 FILLER_17_1286 ();
 sg13g2_decap_8 FILLER_17_1293 ();
 sg13g2_decap_8 FILLER_17_1300 ();
 sg13g2_fill_1 FILLER_17_1307 ();
 sg13g2_fill_1 FILLER_17_1316 ();
 sg13g2_decap_4 FILLER_17_1320 ();
 sg13g2_fill_2 FILLER_17_1324 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_4 FILLER_18_35 ();
 sg13g2_fill_1 FILLER_18_39 ();
 sg13g2_fill_2 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_70 ();
 sg13g2_fill_1 FILLER_18_101 ();
 sg13g2_decap_8 FILLER_18_106 ();
 sg13g2_decap_8 FILLER_18_113 ();
 sg13g2_decap_4 FILLER_18_120 ();
 sg13g2_fill_1 FILLER_18_124 ();
 sg13g2_decap_8 FILLER_18_138 ();
 sg13g2_decap_8 FILLER_18_145 ();
 sg13g2_decap_8 FILLER_18_152 ();
 sg13g2_decap_8 FILLER_18_159 ();
 sg13g2_decap_4 FILLER_18_166 ();
 sg13g2_fill_1 FILLER_18_170 ();
 sg13g2_decap_4 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_212 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_fill_2 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_235 ();
 sg13g2_decap_4 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_261 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_decap_4 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_296 ();
 sg13g2_decap_4 FILLER_18_300 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_2 FILLER_18_331 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_367 ();
 sg13g2_fill_1 FILLER_18_374 ();
 sg13g2_decap_4 FILLER_18_389 ();
 sg13g2_decap_4 FILLER_18_397 ();
 sg13g2_fill_2 FILLER_18_401 ();
 sg13g2_decap_8 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_18_426 ();
 sg13g2_fill_1 FILLER_18_433 ();
 sg13g2_decap_8 FILLER_18_437 ();
 sg13g2_decap_8 FILLER_18_444 ();
 sg13g2_decap_4 FILLER_18_451 ();
 sg13g2_fill_1 FILLER_18_455 ();
 sg13g2_fill_1 FILLER_18_468 ();
 sg13g2_fill_1 FILLER_18_474 ();
 sg13g2_decap_8 FILLER_18_493 ();
 sg13g2_decap_4 FILLER_18_500 ();
 sg13g2_fill_1 FILLER_18_509 ();
 sg13g2_decap_4 FILLER_18_514 ();
 sg13g2_decap_4 FILLER_18_529 ();
 sg13g2_fill_1 FILLER_18_543 ();
 sg13g2_fill_1 FILLER_18_548 ();
 sg13g2_fill_1 FILLER_18_553 ();
 sg13g2_fill_1 FILLER_18_559 ();
 sg13g2_fill_1 FILLER_18_565 ();
 sg13g2_decap_8 FILLER_18_575 ();
 sg13g2_fill_2 FILLER_18_582 ();
 sg13g2_fill_1 FILLER_18_584 ();
 sg13g2_fill_1 FILLER_18_602 ();
 sg13g2_fill_1 FILLER_18_609 ();
 sg13g2_fill_1 FILLER_18_614 ();
 sg13g2_fill_2 FILLER_18_620 ();
 sg13g2_fill_1 FILLER_18_627 ();
 sg13g2_fill_1 FILLER_18_637 ();
 sg13g2_fill_1 FILLER_18_643 ();
 sg13g2_fill_1 FILLER_18_650 ();
 sg13g2_decap_8 FILLER_18_657 ();
 sg13g2_fill_2 FILLER_18_664 ();
 sg13g2_fill_1 FILLER_18_674 ();
 sg13g2_decap_8 FILLER_18_680 ();
 sg13g2_decap_8 FILLER_18_687 ();
 sg13g2_fill_1 FILLER_18_702 ();
 sg13g2_fill_1 FILLER_18_706 ();
 sg13g2_decap_8 FILLER_18_739 ();
 sg13g2_fill_1 FILLER_18_756 ();
 sg13g2_decap_4 FILLER_18_760 ();
 sg13g2_fill_2 FILLER_18_764 ();
 sg13g2_decap_8 FILLER_18_772 ();
 sg13g2_decap_8 FILLER_18_779 ();
 sg13g2_fill_1 FILLER_18_786 ();
 sg13g2_decap_8 FILLER_18_790 ();
 sg13g2_decap_8 FILLER_18_867 ();
 sg13g2_decap_8 FILLER_18_874 ();
 sg13g2_decap_8 FILLER_18_881 ();
 sg13g2_decap_4 FILLER_18_888 ();
 sg13g2_fill_2 FILLER_18_892 ();
 sg13g2_fill_2 FILLER_18_902 ();
 sg13g2_fill_1 FILLER_18_904 ();
 sg13g2_fill_2 FILLER_18_912 ();
 sg13g2_fill_2 FILLER_18_918 ();
 sg13g2_fill_1 FILLER_18_920 ();
 sg13g2_fill_2 FILLER_18_926 ();
 sg13g2_fill_1 FILLER_18_928 ();
 sg13g2_decap_8 FILLER_18_933 ();
 sg13g2_decap_8 FILLER_18_940 ();
 sg13g2_decap_8 FILLER_18_947 ();
 sg13g2_fill_2 FILLER_18_954 ();
 sg13g2_fill_1 FILLER_18_956 ();
 sg13g2_decap_8 FILLER_18_966 ();
 sg13g2_decap_8 FILLER_18_973 ();
 sg13g2_decap_4 FILLER_18_980 ();
 sg13g2_fill_2 FILLER_18_984 ();
 sg13g2_fill_2 FILLER_18_1009 ();
 sg13g2_fill_1 FILLER_18_1011 ();
 sg13g2_fill_1 FILLER_18_1027 ();
 sg13g2_decap_8 FILLER_18_1033 ();
 sg13g2_decap_8 FILLER_18_1040 ();
 sg13g2_decap_4 FILLER_18_1047 ();
 sg13g2_fill_2 FILLER_18_1051 ();
 sg13g2_fill_1 FILLER_18_1069 ();
 sg13g2_fill_1 FILLER_18_1076 ();
 sg13g2_fill_1 FILLER_18_1085 ();
 sg13g2_decap_8 FILLER_18_1089 ();
 sg13g2_fill_2 FILLER_18_1101 ();
 sg13g2_fill_1 FILLER_18_1103 ();
 sg13g2_decap_4 FILLER_18_1108 ();
 sg13g2_fill_1 FILLER_18_1112 ();
 sg13g2_decap_4 FILLER_18_1118 ();
 sg13g2_fill_1 FILLER_18_1122 ();
 sg13g2_decap_8 FILLER_18_1140 ();
 sg13g2_fill_2 FILLER_18_1147 ();
 sg13g2_fill_1 FILLER_18_1149 ();
 sg13g2_decap_4 FILLER_18_1153 ();
 sg13g2_fill_2 FILLER_18_1157 ();
 sg13g2_fill_1 FILLER_18_1163 ();
 sg13g2_fill_1 FILLER_18_1168 ();
 sg13g2_decap_4 FILLER_18_1185 ();
 sg13g2_fill_2 FILLER_18_1194 ();
 sg13g2_fill_1 FILLER_18_1196 ();
 sg13g2_fill_2 FILLER_18_1205 ();
 sg13g2_fill_1 FILLER_18_1213 ();
 sg13g2_fill_2 FILLER_18_1220 ();
 sg13g2_fill_1 FILLER_18_1225 ();
 sg13g2_fill_1 FILLER_18_1233 ();
 sg13g2_fill_1 FILLER_18_1242 ();
 sg13g2_fill_2 FILLER_18_1246 ();
 sg13g2_fill_2 FILLER_18_1256 ();
 sg13g2_fill_1 FILLER_18_1258 ();
 sg13g2_fill_1 FILLER_18_1267 ();
 sg13g2_fill_2 FILLER_18_1274 ();
 sg13g2_fill_2 FILLER_18_1280 ();
 sg13g2_fill_2 FILLER_18_1286 ();
 sg13g2_fill_1 FILLER_18_1288 ();
 sg13g2_decap_8 FILLER_18_1293 ();
 sg13g2_decap_4 FILLER_18_1300 ();
 sg13g2_fill_1 FILLER_18_1304 ();
 sg13g2_fill_2 FILLER_18_1313 ();
 sg13g2_fill_2 FILLER_18_1324 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_fill_1 FILLER_19_10 ();
 sg13g2_decap_8 FILLER_19_16 ();
 sg13g2_fill_2 FILLER_19_23 ();
 sg13g2_decap_8 FILLER_19_29 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_fill_2 FILLER_19_59 ();
 sg13g2_decap_8 FILLER_19_71 ();
 sg13g2_decap_8 FILLER_19_78 ();
 sg13g2_fill_1 FILLER_19_89 ();
 sg13g2_fill_1 FILLER_19_94 ();
 sg13g2_fill_1 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_107 ();
 sg13g2_decap_4 FILLER_19_114 ();
 sg13g2_fill_2 FILLER_19_118 ();
 sg13g2_fill_2 FILLER_19_124 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_141 ();
 sg13g2_fill_2 FILLER_19_148 ();
 sg13g2_fill_1 FILLER_19_150 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_decap_4 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_180 ();
 sg13g2_fill_2 FILLER_19_187 ();
 sg13g2_decap_4 FILLER_19_202 ();
 sg13g2_fill_2 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_220 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_236 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_fill_2 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_fill_2 FILLER_19_277 ();
 sg13g2_fill_1 FILLER_19_283 ();
 sg13g2_fill_2 FILLER_19_295 ();
 sg13g2_decap_4 FILLER_19_302 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_324 ();
 sg13g2_fill_1 FILLER_19_330 ();
 sg13g2_fill_1 FILLER_19_336 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_347 ();
 sg13g2_decap_4 FILLER_19_354 ();
 sg13g2_fill_1 FILLER_19_358 ();
 sg13g2_decap_8 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_decap_4 FILLER_19_388 ();
 sg13g2_fill_1 FILLER_19_392 ();
 sg13g2_decap_4 FILLER_19_411 ();
 sg13g2_decap_4 FILLER_19_420 ();
 sg13g2_decap_4 FILLER_19_430 ();
 sg13g2_fill_1 FILLER_19_434 ();
 sg13g2_fill_2 FILLER_19_462 ();
 sg13g2_fill_2 FILLER_19_469 ();
 sg13g2_fill_1 FILLER_19_471 ();
 sg13g2_fill_2 FILLER_19_484 ();
 sg13g2_fill_1 FILLER_19_496 ();
 sg13g2_decap_8 FILLER_19_502 ();
 sg13g2_decap_8 FILLER_19_509 ();
 sg13g2_fill_2 FILLER_19_516 ();
 sg13g2_fill_1 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_523 ();
 sg13g2_fill_2 FILLER_19_555 ();
 sg13g2_fill_2 FILLER_19_561 ();
 sg13g2_fill_2 FILLER_19_568 ();
 sg13g2_fill_1 FILLER_19_570 ();
 sg13g2_decap_4 FILLER_19_576 ();
 sg13g2_fill_1 FILLER_19_580 ();
 sg13g2_fill_1 FILLER_19_589 ();
 sg13g2_decap_8 FILLER_19_607 ();
 sg13g2_fill_2 FILLER_19_614 ();
 sg13g2_decap_8 FILLER_19_624 ();
 sg13g2_decap_4 FILLER_19_631 ();
 sg13g2_fill_2 FILLER_19_635 ();
 sg13g2_fill_1 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_655 ();
 sg13g2_decap_8 FILLER_19_662 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_decap_8 FILLER_19_676 ();
 sg13g2_decap_4 FILLER_19_683 ();
 sg13g2_fill_2 FILLER_19_691 ();
 sg13g2_fill_2 FILLER_19_709 ();
 sg13g2_fill_1 FILLER_19_711 ();
 sg13g2_fill_2 FILLER_19_716 ();
 sg13g2_fill_2 FILLER_19_722 ();
 sg13g2_decap_4 FILLER_19_759 ();
 sg13g2_fill_2 FILLER_19_766 ();
 sg13g2_decap_8 FILLER_19_773 ();
 sg13g2_decap_8 FILLER_19_780 ();
 sg13g2_decap_8 FILLER_19_787 ();
 sg13g2_decap_8 FILLER_19_794 ();
 sg13g2_fill_1 FILLER_19_801 ();
 sg13g2_decap_8 FILLER_19_806 ();
 sg13g2_fill_2 FILLER_19_813 ();
 sg13g2_decap_4 FILLER_19_818 ();
 sg13g2_fill_1 FILLER_19_822 ();
 sg13g2_fill_1 FILLER_19_831 ();
 sg13g2_fill_1 FILLER_19_850 ();
 sg13g2_decap_4 FILLER_19_873 ();
 sg13g2_fill_2 FILLER_19_877 ();
 sg13g2_decap_8 FILLER_19_883 ();
 sg13g2_decap_4 FILLER_19_890 ();
 sg13g2_fill_1 FILLER_19_894 ();
 sg13g2_fill_2 FILLER_19_899 ();
 sg13g2_fill_1 FILLER_19_901 ();
 sg13g2_decap_4 FILLER_19_906 ();
 sg13g2_fill_1 FILLER_19_913 ();
 sg13g2_fill_1 FILLER_19_918 ();
 sg13g2_decap_8 FILLER_19_942 ();
 sg13g2_decap_4 FILLER_19_949 ();
 sg13g2_fill_2 FILLER_19_953 ();
 sg13g2_decap_4 FILLER_19_967 ();
 sg13g2_fill_1 FILLER_19_985 ();
 sg13g2_fill_2 FILLER_19_992 ();
 sg13g2_fill_1 FILLER_19_994 ();
 sg13g2_fill_2 FILLER_19_1004 ();
 sg13g2_fill_1 FILLER_19_1006 ();
 sg13g2_decap_4 FILLER_19_1014 ();
 sg13g2_fill_1 FILLER_19_1018 ();
 sg13g2_fill_2 FILLER_19_1023 ();
 sg13g2_fill_2 FILLER_19_1033 ();
 sg13g2_fill_1 FILLER_19_1035 ();
 sg13g2_decap_4 FILLER_19_1041 ();
 sg13g2_fill_2 FILLER_19_1045 ();
 sg13g2_fill_1 FILLER_19_1052 ();
 sg13g2_decap_4 FILLER_19_1067 ();
 sg13g2_fill_1 FILLER_19_1071 ();
 sg13g2_fill_1 FILLER_19_1083 ();
 sg13g2_decap_4 FILLER_19_1088 ();
 sg13g2_fill_2 FILLER_19_1117 ();
 sg13g2_fill_1 FILLER_19_1124 ();
 sg13g2_fill_1 FILLER_19_1130 ();
 sg13g2_fill_1 FILLER_19_1148 ();
 sg13g2_fill_1 FILLER_19_1171 ();
 sg13g2_fill_1 FILLER_19_1175 ();
 sg13g2_fill_2 FILLER_19_1206 ();
 sg13g2_fill_1 FILLER_19_1222 ();
 sg13g2_fill_1 FILLER_19_1230 ();
 sg13g2_fill_1 FILLER_19_1235 ();
 sg13g2_decap_4 FILLER_19_1248 ();
 sg13g2_fill_2 FILLER_19_1252 ();
 sg13g2_fill_1 FILLER_19_1258 ();
 sg13g2_fill_2 FILLER_19_1277 ();
 sg13g2_fill_1 FILLER_19_1283 ();
 sg13g2_fill_2 FILLER_19_1304 ();
 sg13g2_fill_1 FILLER_19_1306 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_33 ();
 sg13g2_fill_1 FILLER_20_39 ();
 sg13g2_fill_2 FILLER_20_44 ();
 sg13g2_fill_1 FILLER_20_46 ();
 sg13g2_fill_2 FILLER_20_59 ();
 sg13g2_fill_1 FILLER_20_64 ();
 sg13g2_decap_4 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_76 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_fill_1 FILLER_20_83 ();
 sg13g2_fill_2 FILLER_20_93 ();
 sg13g2_fill_1 FILLER_20_106 ();
 sg13g2_fill_1 FILLER_20_118 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_fill_1 FILLER_20_130 ();
 sg13g2_fill_2 FILLER_20_169 ();
 sg13g2_decap_8 FILLER_20_181 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_decap_4 FILLER_20_265 ();
 sg13g2_fill_2 FILLER_20_269 ();
 sg13g2_fill_1 FILLER_20_276 ();
 sg13g2_fill_1 FILLER_20_280 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_292 ();
 sg13g2_fill_1 FILLER_20_296 ();
 sg13g2_fill_1 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_fill_2 FILLER_20_382 ();
 sg13g2_fill_1 FILLER_20_384 ();
 sg13g2_fill_1 FILLER_20_399 ();
 sg13g2_fill_1 FILLER_20_403 ();
 sg13g2_decap_4 FILLER_20_409 ();
 sg13g2_fill_1 FILLER_20_413 ();
 sg13g2_fill_1 FILLER_20_436 ();
 sg13g2_fill_1 FILLER_20_443 ();
 sg13g2_fill_1 FILLER_20_449 ();
 sg13g2_fill_2 FILLER_20_455 ();
 sg13g2_fill_1 FILLER_20_457 ();
 sg13g2_decap_8 FILLER_20_463 ();
 sg13g2_decap_4 FILLER_20_495 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_4 FILLER_20_539 ();
 sg13g2_fill_1 FILLER_20_543 ();
 sg13g2_fill_2 FILLER_20_581 ();
 sg13g2_fill_2 FILLER_20_588 ();
 sg13g2_fill_1 FILLER_20_590 ();
 sg13g2_fill_2 FILLER_20_605 ();
 sg13g2_fill_2 FILLER_20_612 ();
 sg13g2_decap_8 FILLER_20_622 ();
 sg13g2_decap_4 FILLER_20_629 ();
 sg13g2_fill_2 FILLER_20_633 ();
 sg13g2_fill_2 FILLER_20_638 ();
 sg13g2_fill_1 FILLER_20_649 ();
 sg13g2_decap_8 FILLER_20_654 ();
 sg13g2_decap_8 FILLER_20_661 ();
 sg13g2_decap_8 FILLER_20_668 ();
 sg13g2_decap_4 FILLER_20_675 ();
 sg13g2_fill_2 FILLER_20_692 ();
 sg13g2_fill_1 FILLER_20_694 ();
 sg13g2_fill_2 FILLER_20_702 ();
 sg13g2_fill_1 FILLER_20_707 ();
 sg13g2_fill_2 FILLER_20_713 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_decap_4 FILLER_20_726 ();
 sg13g2_fill_1 FILLER_20_730 ();
 sg13g2_fill_2 FILLER_20_743 ();
 sg13g2_fill_1 FILLER_20_745 ();
 sg13g2_fill_1 FILLER_20_754 ();
 sg13g2_fill_2 FILLER_20_775 ();
 sg13g2_fill_1 FILLER_20_777 ();
 sg13g2_decap_4 FILLER_20_782 ();
 sg13g2_decap_4 FILLER_20_807 ();
 sg13g2_fill_2 FILLER_20_817 ();
 sg13g2_fill_1 FILLER_20_827 ();
 sg13g2_fill_2 FILLER_20_831 ();
 sg13g2_fill_2 FILLER_20_838 ();
 sg13g2_decap_8 FILLER_20_857 ();
 sg13g2_decap_4 FILLER_20_864 ();
 sg13g2_fill_2 FILLER_20_868 ();
 sg13g2_fill_1 FILLER_20_875 ();
 sg13g2_fill_2 FILLER_20_902 ();
 sg13g2_fill_1 FILLER_20_904 ();
 sg13g2_fill_1 FILLER_20_932 ();
 sg13g2_fill_2 FILLER_20_954 ();
 sg13g2_fill_2 FILLER_20_965 ();
 sg13g2_fill_2 FILLER_20_970 ();
 sg13g2_decap_8 FILLER_20_975 ();
 sg13g2_decap_8 FILLER_20_982 ();
 sg13g2_fill_2 FILLER_20_989 ();
 sg13g2_decap_8 FILLER_20_1007 ();
 sg13g2_fill_2 FILLER_20_1014 ();
 sg13g2_decap_8 FILLER_20_1026 ();
 sg13g2_fill_1 FILLER_20_1033 ();
 sg13g2_fill_1 FILLER_20_1038 ();
 sg13g2_fill_2 FILLER_20_1044 ();
 sg13g2_fill_1 FILLER_20_1050 ();
 sg13g2_fill_1 FILLER_20_1057 ();
 sg13g2_fill_1 FILLER_20_1067 ();
 sg13g2_fill_2 FILLER_20_1085 ();
 sg13g2_decap_8 FILLER_20_1092 ();
 sg13g2_decap_4 FILLER_20_1099 ();
 sg13g2_decap_4 FILLER_20_1107 ();
 sg13g2_fill_2 FILLER_20_1111 ();
 sg13g2_fill_1 FILLER_20_1117 ();
 sg13g2_fill_1 FILLER_20_1128 ();
 sg13g2_fill_1 FILLER_20_1134 ();
 sg13g2_fill_1 FILLER_20_1139 ();
 sg13g2_decap_8 FILLER_20_1149 ();
 sg13g2_decap_4 FILLER_20_1156 ();
 sg13g2_fill_2 FILLER_20_1175 ();
 sg13g2_decap_4 FILLER_20_1185 ();
 sg13g2_fill_1 FILLER_20_1189 ();
 sg13g2_decap_8 FILLER_20_1193 ();
 sg13g2_fill_1 FILLER_20_1200 ();
 sg13g2_fill_1 FILLER_20_1249 ();
 sg13g2_fill_1 FILLER_20_1267 ();
 sg13g2_decap_8 FILLER_20_1272 ();
 sg13g2_decap_8 FILLER_20_1279 ();
 sg13g2_decap_8 FILLER_20_1286 ();
 sg13g2_decap_8 FILLER_20_1293 ();
 sg13g2_decap_8 FILLER_20_1300 ();
 sg13g2_fill_1 FILLER_20_1307 ();
 sg13g2_decap_8 FILLER_20_1312 ();
 sg13g2_decap_8 FILLER_20_1319 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_40 ();
 sg13g2_decap_4 FILLER_21_47 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_decap_8 FILLER_21_57 ();
 sg13g2_decap_8 FILLER_21_64 ();
 sg13g2_fill_2 FILLER_21_71 ();
 sg13g2_fill_1 FILLER_21_73 ();
 sg13g2_fill_2 FILLER_21_83 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_fill_2 FILLER_21_103 ();
 sg13g2_fill_2 FILLER_21_109 ();
 sg13g2_fill_2 FILLER_21_117 ();
 sg13g2_decap_4 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_fill_1 FILLER_21_207 ();
 sg13g2_fill_2 FILLER_21_219 ();
 sg13g2_decap_8 FILLER_21_229 ();
 sg13g2_fill_2 FILLER_21_236 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_244 ();
 sg13g2_fill_2 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_282 ();
 sg13g2_fill_1 FILLER_21_288 ();
 sg13g2_decap_8 FILLER_21_303 ();
 sg13g2_fill_1 FILLER_21_310 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_decap_4 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_fill_2 FILLER_21_365 ();
 sg13g2_fill_2 FILLER_21_371 ();
 sg13g2_fill_2 FILLER_21_378 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_405 ();
 sg13g2_fill_1 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_21_421 ();
 sg13g2_decap_8 FILLER_21_428 ();
 sg13g2_decap_4 FILLER_21_435 ();
 sg13g2_decap_8 FILLER_21_444 ();
 sg13g2_fill_2 FILLER_21_451 ();
 sg13g2_fill_1 FILLER_21_453 ();
 sg13g2_decap_8 FILLER_21_464 ();
 sg13g2_fill_1 FILLER_21_471 ();
 sg13g2_fill_2 FILLER_21_490 ();
 sg13g2_fill_1 FILLER_21_492 ();
 sg13g2_decap_4 FILLER_21_501 ();
 sg13g2_fill_2 FILLER_21_505 ();
 sg13g2_fill_2 FILLER_21_513 ();
 sg13g2_fill_1 FILLER_21_515 ();
 sg13g2_decap_8 FILLER_21_524 ();
 sg13g2_decap_4 FILLER_21_531 ();
 sg13g2_fill_2 FILLER_21_535 ();
 sg13g2_fill_2 FILLER_21_543 ();
 sg13g2_fill_2 FILLER_21_554 ();
 sg13g2_fill_1 FILLER_21_556 ();
 sg13g2_fill_1 FILLER_21_562 ();
 sg13g2_fill_2 FILLER_21_568 ();
 sg13g2_fill_2 FILLER_21_574 ();
 sg13g2_fill_2 FILLER_21_604 ();
 sg13g2_fill_1 FILLER_21_618 ();
 sg13g2_fill_1 FILLER_21_631 ();
 sg13g2_fill_2 FILLER_21_636 ();
 sg13g2_fill_1 FILLER_21_638 ();
 sg13g2_fill_1 FILLER_21_647 ();
 sg13g2_decap_4 FILLER_21_653 ();
 sg13g2_fill_1 FILLER_21_657 ();
 sg13g2_decap_8 FILLER_21_689 ();
 sg13g2_fill_1 FILLER_21_696 ();
 sg13g2_fill_2 FILLER_21_725 ();
 sg13g2_fill_2 FILLER_21_731 ();
 sg13g2_fill_1 FILLER_21_733 ();
 sg13g2_fill_1 FILLER_21_738 ();
 sg13g2_fill_2 FILLER_21_744 ();
 sg13g2_fill_1 FILLER_21_746 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_fill_2 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_769 ();
 sg13g2_decap_8 FILLER_21_776 ();
 sg13g2_decap_4 FILLER_21_783 ();
 sg13g2_fill_1 FILLER_21_787 ();
 sg13g2_fill_2 FILLER_21_804 ();
 sg13g2_fill_2 FILLER_21_823 ();
 sg13g2_fill_1 FILLER_21_852 ();
 sg13g2_decap_8 FILLER_21_879 ();
 sg13g2_decap_4 FILLER_21_886 ();
 sg13g2_fill_2 FILLER_21_893 ();
 sg13g2_fill_1 FILLER_21_895 ();
 sg13g2_fill_2 FILLER_21_905 ();
 sg13g2_fill_1 FILLER_21_907 ();
 sg13g2_fill_1 FILLER_21_913 ();
 sg13g2_fill_1 FILLER_21_917 ();
 sg13g2_fill_1 FILLER_21_921 ();
 sg13g2_fill_1 FILLER_21_927 ();
 sg13g2_fill_2 FILLER_21_931 ();
 sg13g2_fill_2 FILLER_21_941 ();
 sg13g2_fill_1 FILLER_21_943 ();
 sg13g2_decap_8 FILLER_21_948 ();
 sg13g2_fill_2 FILLER_21_955 ();
 sg13g2_fill_1 FILLER_21_957 ();
 sg13g2_decap_8 FILLER_21_979 ();
 sg13g2_fill_1 FILLER_21_986 ();
 sg13g2_fill_2 FILLER_21_1000 ();
 sg13g2_fill_1 FILLER_21_1002 ();
 sg13g2_decap_8 FILLER_21_1008 ();
 sg13g2_decap_4 FILLER_21_1015 ();
 sg13g2_fill_2 FILLER_21_1019 ();
 sg13g2_fill_1 FILLER_21_1025 ();
 sg13g2_decap_8 FILLER_21_1032 ();
 sg13g2_fill_2 FILLER_21_1039 ();
 sg13g2_decap_8 FILLER_21_1044 ();
 sg13g2_fill_2 FILLER_21_1055 ();
 sg13g2_decap_4 FILLER_21_1061 ();
 sg13g2_fill_2 FILLER_21_1081 ();
 sg13g2_fill_2 FILLER_21_1108 ();
 sg13g2_fill_2 FILLER_21_1114 ();
 sg13g2_fill_2 FILLER_21_1120 ();
 sg13g2_decap_4 FILLER_21_1129 ();
 sg13g2_fill_1 FILLER_21_1137 ();
 sg13g2_decap_8 FILLER_21_1144 ();
 sg13g2_fill_2 FILLER_21_1151 ();
 sg13g2_fill_1 FILLER_21_1153 ();
 sg13g2_fill_1 FILLER_21_1183 ();
 sg13g2_fill_1 FILLER_21_1189 ();
 sg13g2_fill_2 FILLER_21_1194 ();
 sg13g2_fill_1 FILLER_21_1196 ();
 sg13g2_fill_1 FILLER_21_1205 ();
 sg13g2_fill_1 FILLER_21_1215 ();
 sg13g2_fill_2 FILLER_21_1232 ();
 sg13g2_fill_2 FILLER_21_1238 ();
 sg13g2_fill_1 FILLER_21_1265 ();
 sg13g2_fill_2 FILLER_21_1270 ();
 sg13g2_decap_8 FILLER_21_1276 ();
 sg13g2_decap_8 FILLER_21_1283 ();
 sg13g2_decap_4 FILLER_21_1290 ();
 sg13g2_fill_2 FILLER_21_1294 ();
 sg13g2_fill_2 FILLER_21_1312 ();
 sg13g2_fill_2 FILLER_21_1323 ();
 sg13g2_fill_1 FILLER_21_1325 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_13 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_57 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_2 FILLER_22_75 ();
 sg13g2_decap_4 FILLER_22_122 ();
 sg13g2_decap_8 FILLER_22_139 ();
 sg13g2_decap_8 FILLER_22_146 ();
 sg13g2_decap_4 FILLER_22_153 ();
 sg13g2_fill_2 FILLER_22_157 ();
 sg13g2_fill_2 FILLER_22_162 ();
 sg13g2_fill_1 FILLER_22_164 ();
 sg13g2_decap_8 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_fill_2 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_fill_1 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_251 ();
 sg13g2_fill_1 FILLER_22_258 ();
 sg13g2_decap_4 FILLER_22_263 ();
 sg13g2_fill_1 FILLER_22_267 ();
 sg13g2_decap_8 FILLER_22_279 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_313 ();
 sg13g2_fill_2 FILLER_22_320 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_fill_2 FILLER_22_329 ();
 sg13g2_fill_1 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_8 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_351 ();
 sg13g2_decap_4 FILLER_22_358 ();
 sg13g2_fill_1 FILLER_22_362 ();
 sg13g2_fill_2 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_398 ();
 sg13g2_fill_1 FILLER_22_407 ();
 sg13g2_fill_1 FILLER_22_417 ();
 sg13g2_decap_4 FILLER_22_426 ();
 sg13g2_fill_1 FILLER_22_430 ();
 sg13g2_decap_8 FILLER_22_436 ();
 sg13g2_fill_1 FILLER_22_443 ();
 sg13g2_fill_2 FILLER_22_448 ();
 sg13g2_fill_1 FILLER_22_450 ();
 sg13g2_fill_1 FILLER_22_461 ();
 sg13g2_fill_1 FILLER_22_466 ();
 sg13g2_fill_1 FILLER_22_477 ();
 sg13g2_fill_1 FILLER_22_482 ();
 sg13g2_decap_4 FILLER_22_491 ();
 sg13g2_fill_1 FILLER_22_500 ();
 sg13g2_fill_2 FILLER_22_507 ();
 sg13g2_decap_8 FILLER_22_513 ();
 sg13g2_decap_8 FILLER_22_520 ();
 sg13g2_decap_4 FILLER_22_527 ();
 sg13g2_fill_2 FILLER_22_531 ();
 sg13g2_fill_1 FILLER_22_538 ();
 sg13g2_fill_1 FILLER_22_543 ();
 sg13g2_fill_1 FILLER_22_567 ();
 sg13g2_decap_4 FILLER_22_577 ();
 sg13g2_fill_1 FILLER_22_585 ();
 sg13g2_decap_8 FILLER_22_591 ();
 sg13g2_fill_1 FILLER_22_601 ();
 sg13g2_fill_1 FILLER_22_610 ();
 sg13g2_decap_8 FILLER_22_624 ();
 sg13g2_decap_4 FILLER_22_631 ();
 sg13g2_fill_1 FILLER_22_635 ();
 sg13g2_fill_1 FILLER_22_643 ();
 sg13g2_decap_4 FILLER_22_649 ();
 sg13g2_decap_4 FILLER_22_663 ();
 sg13g2_decap_4 FILLER_22_675 ();
 sg13g2_fill_2 FILLER_22_683 ();
 sg13g2_fill_2 FILLER_22_699 ();
 sg13g2_fill_1 FILLER_22_701 ();
 sg13g2_fill_2 FILLER_22_706 ();
 sg13g2_fill_2 FILLER_22_712 ();
 sg13g2_decap_8 FILLER_22_719 ();
 sg13g2_fill_1 FILLER_22_726 ();
 sg13g2_fill_1 FILLER_22_737 ();
 sg13g2_decap_8 FILLER_22_741 ();
 sg13g2_decap_8 FILLER_22_760 ();
 sg13g2_fill_2 FILLER_22_767 ();
 sg13g2_decap_8 FILLER_22_778 ();
 sg13g2_fill_2 FILLER_22_785 ();
 sg13g2_fill_1 FILLER_22_787 ();
 sg13g2_fill_1 FILLER_22_800 ();
 sg13g2_fill_2 FILLER_22_805 ();
 sg13g2_decap_4 FILLER_22_810 ();
 sg13g2_fill_2 FILLER_22_819 ();
 sg13g2_decap_4 FILLER_22_826 ();
 sg13g2_fill_1 FILLER_22_835 ();
 sg13g2_decap_8 FILLER_22_846 ();
 sg13g2_decap_4 FILLER_22_856 ();
 sg13g2_decap_8 FILLER_22_865 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_fill_1 FILLER_22_879 ();
 sg13g2_decap_4 FILLER_22_890 ();
 sg13g2_fill_1 FILLER_22_894 ();
 sg13g2_decap_4 FILLER_22_905 ();
 sg13g2_fill_1 FILLER_22_919 ();
 sg13g2_fill_1 FILLER_22_938 ();
 sg13g2_decap_8 FILLER_22_953 ();
 sg13g2_decap_4 FILLER_22_964 ();
 sg13g2_decap_8 FILLER_22_977 ();
 sg13g2_decap_8 FILLER_22_984 ();
 sg13g2_decap_4 FILLER_22_991 ();
 sg13g2_fill_2 FILLER_22_995 ();
 sg13g2_fill_2 FILLER_22_1007 ();
 sg13g2_fill_2 FILLER_22_1029 ();
 sg13g2_fill_1 FILLER_22_1040 ();
 sg13g2_decap_8 FILLER_22_1047 ();
 sg13g2_decap_4 FILLER_22_1054 ();
 sg13g2_decap_4 FILLER_22_1066 ();
 sg13g2_fill_2 FILLER_22_1070 ();
 sg13g2_decap_8 FILLER_22_1081 ();
 sg13g2_decap_8 FILLER_22_1092 ();
 sg13g2_decap_8 FILLER_22_1099 ();
 sg13g2_fill_2 FILLER_22_1106 ();
 sg13g2_fill_1 FILLER_22_1120 ();
 sg13g2_fill_1 FILLER_22_1125 ();
 sg13g2_fill_2 FILLER_22_1133 ();
 sg13g2_decap_8 FILLER_22_1145 ();
 sg13g2_fill_2 FILLER_22_1152 ();
 sg13g2_decap_8 FILLER_22_1162 ();
 sg13g2_fill_2 FILLER_22_1169 ();
 sg13g2_decap_8 FILLER_22_1174 ();
 sg13g2_decap_8 FILLER_22_1181 ();
 sg13g2_fill_2 FILLER_22_1188 ();
 sg13g2_fill_1 FILLER_22_1190 ();
 sg13g2_fill_2 FILLER_22_1196 ();
 sg13g2_fill_1 FILLER_22_1213 ();
 sg13g2_fill_1 FILLER_22_1218 ();
 sg13g2_fill_2 FILLER_22_1223 ();
 sg13g2_decap_8 FILLER_22_1243 ();
 sg13g2_fill_2 FILLER_22_1250 ();
 sg13g2_fill_1 FILLER_22_1252 ();
 sg13g2_fill_2 FILLER_22_1256 ();
 sg13g2_fill_1 FILLER_22_1258 ();
 sg13g2_decap_8 FILLER_22_1262 ();
 sg13g2_decap_4 FILLER_22_1269 ();
 sg13g2_fill_1 FILLER_22_1273 ();
 sg13g2_decap_8 FILLER_22_1281 ();
 sg13g2_decap_8 FILLER_22_1288 ();
 sg13g2_decap_8 FILLER_22_1295 ();
 sg13g2_decap_4 FILLER_22_1302 ();
 sg13g2_fill_2 FILLER_22_1306 ();
 sg13g2_decap_8 FILLER_22_1319 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_51 ();
 sg13g2_decap_4 FILLER_23_73 ();
 sg13g2_fill_1 FILLER_23_120 ();
 sg13g2_fill_1 FILLER_23_159 ();
 sg13g2_decap_8 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_4 FILLER_23_224 ();
 sg13g2_fill_2 FILLER_23_228 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_2 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_249 ();
 sg13g2_decap_4 FILLER_23_255 ();
 sg13g2_decap_4 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_272 ();
 sg13g2_decap_4 FILLER_23_279 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_4 FILLER_23_298 ();
 sg13g2_fill_2 FILLER_23_302 ();
 sg13g2_fill_2 FILLER_23_338 ();
 sg13g2_fill_2 FILLER_23_366 ();
 sg13g2_fill_1 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_fill_1 FILLER_23_384 ();
 sg13g2_fill_2 FILLER_23_389 ();
 sg13g2_fill_1 FILLER_23_394 ();
 sg13g2_fill_2 FILLER_23_400 ();
 sg13g2_decap_8 FILLER_23_424 ();
 sg13g2_decap_8 FILLER_23_431 ();
 sg13g2_fill_2 FILLER_23_438 ();
 sg13g2_fill_1 FILLER_23_440 ();
 sg13g2_fill_1 FILLER_23_450 ();
 sg13g2_fill_1 FILLER_23_456 ();
 sg13g2_fill_2 FILLER_23_468 ();
 sg13g2_fill_1 FILLER_23_470 ();
 sg13g2_decap_4 FILLER_23_484 ();
 sg13g2_fill_2 FILLER_23_488 ();
 sg13g2_decap_4 FILLER_23_535 ();
 sg13g2_fill_1 FILLER_23_539 ();
 sg13g2_fill_1 FILLER_23_547 ();
 sg13g2_decap_8 FILLER_23_552 ();
 sg13g2_fill_2 FILLER_23_559 ();
 sg13g2_fill_1 FILLER_23_561 ();
 sg13g2_fill_1 FILLER_23_574 ();
 sg13g2_fill_2 FILLER_23_584 ();
 sg13g2_decap_4 FILLER_23_591 ();
 sg13g2_fill_1 FILLER_23_595 ();
 sg13g2_fill_2 FILLER_23_609 ();
 sg13g2_fill_1 FILLER_23_620 ();
 sg13g2_fill_2 FILLER_23_627 ();
 sg13g2_decap_4 FILLER_23_637 ();
 sg13g2_decap_4 FILLER_23_645 ();
 sg13g2_fill_1 FILLER_23_649 ();
 sg13g2_decap_8 FILLER_23_655 ();
 sg13g2_decap_8 FILLER_23_662 ();
 sg13g2_decap_8 FILLER_23_669 ();
 sg13g2_fill_2 FILLER_23_676 ();
 sg13g2_decap_4 FILLER_23_694 ();
 sg13g2_fill_1 FILLER_23_698 ();
 sg13g2_fill_2 FILLER_23_714 ();
 sg13g2_fill_1 FILLER_23_726 ();
 sg13g2_fill_1 FILLER_23_738 ();
 sg13g2_fill_1 FILLER_23_744 ();
 sg13g2_fill_2 FILLER_23_749 ();
 sg13g2_fill_1 FILLER_23_751 ();
 sg13g2_fill_1 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_765 ();
 sg13g2_fill_2 FILLER_23_772 ();
 sg13g2_decap_4 FILLER_23_777 ();
 sg13g2_fill_2 FILLER_23_781 ();
 sg13g2_fill_2 FILLER_23_786 ();
 sg13g2_fill_1 FILLER_23_788 ();
 sg13g2_fill_1 FILLER_23_811 ();
 sg13g2_decap_4 FILLER_23_829 ();
 sg13g2_fill_2 FILLER_23_851 ();
 sg13g2_fill_1 FILLER_23_853 ();
 sg13g2_decap_8 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_decap_8 FILLER_23_875 ();
 sg13g2_fill_2 FILLER_23_891 ();
 sg13g2_fill_1 FILLER_23_893 ();
 sg13g2_fill_1 FILLER_23_898 ();
 sg13g2_decap_4 FILLER_23_912 ();
 sg13g2_fill_2 FILLER_23_916 ();
 sg13g2_fill_1 FILLER_23_921 ();
 sg13g2_decap_8 FILLER_23_933 ();
 sg13g2_decap_4 FILLER_23_940 ();
 sg13g2_decap_8 FILLER_23_949 ();
 sg13g2_fill_2 FILLER_23_956 ();
 sg13g2_fill_1 FILLER_23_958 ();
 sg13g2_decap_4 FILLER_23_971 ();
 sg13g2_fill_2 FILLER_23_979 ();
 sg13g2_decap_8 FILLER_23_989 ();
 sg13g2_decap_8 FILLER_23_996 ();
 sg13g2_decap_8 FILLER_23_1003 ();
 sg13g2_decap_4 FILLER_23_1010 ();
 sg13g2_fill_2 FILLER_23_1026 ();
 sg13g2_decap_8 FILLER_23_1040 ();
 sg13g2_fill_1 FILLER_23_1054 ();
 sg13g2_decap_8 FILLER_23_1061 ();
 sg13g2_decap_8 FILLER_23_1068 ();
 sg13g2_decap_4 FILLER_23_1075 ();
 sg13g2_fill_1 FILLER_23_1079 ();
 sg13g2_fill_2 FILLER_23_1119 ();
 sg13g2_fill_1 FILLER_23_1121 ();
 sg13g2_decap_8 FILLER_23_1135 ();
 sg13g2_decap_4 FILLER_23_1142 ();
 sg13g2_fill_1 FILLER_23_1146 ();
 sg13g2_fill_2 FILLER_23_1155 ();
 sg13g2_fill_1 FILLER_23_1157 ();
 sg13g2_fill_1 FILLER_23_1162 ();
 sg13g2_fill_2 FILLER_23_1179 ();
 sg13g2_fill_1 FILLER_23_1181 ();
 sg13g2_fill_1 FILLER_23_1206 ();
 sg13g2_fill_1 FILLER_23_1211 ();
 sg13g2_fill_1 FILLER_23_1225 ();
 sg13g2_fill_1 FILLER_23_1234 ();
 sg13g2_decap_8 FILLER_23_1239 ();
 sg13g2_decap_8 FILLER_23_1246 ();
 sg13g2_decap_4 FILLER_23_1253 ();
 sg13g2_fill_1 FILLER_23_1257 ();
 sg13g2_fill_1 FILLER_23_1262 ();
 sg13g2_decap_8 FILLER_23_1297 ();
 sg13g2_fill_2 FILLER_23_1304 ();
 sg13g2_fill_1 FILLER_23_1306 ();
 sg13g2_decap_8 FILLER_23_1319 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_25 ();
 sg13g2_decap_4 FILLER_24_31 ();
 sg13g2_decap_4 FILLER_24_44 ();
 sg13g2_fill_1 FILLER_24_48 ();
 sg13g2_decap_8 FILLER_24_66 ();
 sg13g2_decap_8 FILLER_24_73 ();
 sg13g2_decap_4 FILLER_24_80 ();
 sg13g2_fill_2 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_114 ();
 sg13g2_fill_1 FILLER_24_121 ();
 sg13g2_fill_1 FILLER_24_163 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_4 FILLER_24_182 ();
 sg13g2_fill_2 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_218 ();
 sg13g2_decap_8 FILLER_24_225 ();
 sg13g2_decap_4 FILLER_24_232 ();
 sg13g2_decap_8 FILLER_24_239 ();
 sg13g2_decap_8 FILLER_24_246 ();
 sg13g2_decap_8 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_260 ();
 sg13g2_fill_1 FILLER_24_267 ();
 sg13g2_fill_1 FILLER_24_272 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_fill_1 FILLER_24_281 ();
 sg13g2_decap_4 FILLER_24_286 ();
 sg13g2_fill_1 FILLER_24_290 ();
 sg13g2_fill_2 FILLER_24_300 ();
 sg13g2_fill_1 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_309 ();
 sg13g2_fill_2 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_fill_2 FILLER_24_363 ();
 sg13g2_fill_1 FILLER_24_373 ();
 sg13g2_fill_2 FILLER_24_379 ();
 sg13g2_fill_2 FILLER_24_386 ();
 sg13g2_decap_4 FILLER_24_393 ();
 sg13g2_decap_4 FILLER_24_402 ();
 sg13g2_fill_2 FILLER_24_410 ();
 sg13g2_fill_1 FILLER_24_412 ();
 sg13g2_fill_2 FILLER_24_418 ();
 sg13g2_decap_4 FILLER_24_423 ();
 sg13g2_fill_2 FILLER_24_427 ();
 sg13g2_fill_1 FILLER_24_446 ();
 sg13g2_fill_1 FILLER_24_455 ();
 sg13g2_fill_2 FILLER_24_468 ();
 sg13g2_fill_1 FILLER_24_470 ();
 sg13g2_fill_1 FILLER_24_476 ();
 sg13g2_fill_2 FILLER_24_480 ();
 sg13g2_decap_8 FILLER_24_487 ();
 sg13g2_decap_8 FILLER_24_494 ();
 sg13g2_decap_8 FILLER_24_501 ();
 sg13g2_fill_2 FILLER_24_508 ();
 sg13g2_decap_4 FILLER_24_519 ();
 sg13g2_fill_1 FILLER_24_523 ();
 sg13g2_fill_2 FILLER_24_544 ();
 sg13g2_decap_4 FILLER_24_558 ();
 sg13g2_fill_1 FILLER_24_562 ();
 sg13g2_fill_2 FILLER_24_566 ();
 sg13g2_fill_1 FILLER_24_568 ();
 sg13g2_fill_2 FILLER_24_574 ();
 sg13g2_fill_1 FILLER_24_576 ();
 sg13g2_decap_8 FILLER_24_585 ();
 sg13g2_decap_4 FILLER_24_592 ();
 sg13g2_fill_1 FILLER_24_596 ();
 sg13g2_fill_2 FILLER_24_620 ();
 sg13g2_decap_4 FILLER_24_625 ();
 sg13g2_fill_1 FILLER_24_629 ();
 sg13g2_decap_8 FILLER_24_661 ();
 sg13g2_fill_2 FILLER_24_668 ();
 sg13g2_fill_1 FILLER_24_670 ();
 sg13g2_decap_4 FILLER_24_701 ();
 sg13g2_fill_2 FILLER_24_720 ();
 sg13g2_fill_1 FILLER_24_722 ();
 sg13g2_decap_8 FILLER_24_734 ();
 sg13g2_decap_4 FILLER_24_741 ();
 sg13g2_fill_1 FILLER_24_745 ();
 sg13g2_fill_2 FILLER_24_757 ();
 sg13g2_fill_1 FILLER_24_759 ();
 sg13g2_decap_4 FILLER_24_796 ();
 sg13g2_decap_4 FILLER_24_805 ();
 sg13g2_decap_4 FILLER_24_826 ();
 sg13g2_fill_1 FILLER_24_830 ();
 sg13g2_decap_8 FILLER_24_839 ();
 sg13g2_decap_8 FILLER_24_846 ();
 sg13g2_decap_8 FILLER_24_871 ();
 sg13g2_decap_4 FILLER_24_878 ();
 sg13g2_fill_1 FILLER_24_882 ();
 sg13g2_fill_2 FILLER_24_888 ();
 sg13g2_decap_4 FILLER_24_893 ();
 sg13g2_decap_8 FILLER_24_908 ();
 sg13g2_fill_2 FILLER_24_915 ();
 sg13g2_fill_1 FILLER_24_917 ();
 sg13g2_fill_1 FILLER_24_938 ();
 sg13g2_decap_4 FILLER_24_948 ();
 sg13g2_decap_8 FILLER_24_956 ();
 sg13g2_decap_4 FILLER_24_963 ();
 sg13g2_fill_1 FILLER_24_967 ();
 sg13g2_decap_8 FILLER_24_973 ();
 sg13g2_decap_8 FILLER_24_980 ();
 sg13g2_decap_4 FILLER_24_987 ();
 sg13g2_fill_2 FILLER_24_991 ();
 sg13g2_decap_8 FILLER_24_998 ();
 sg13g2_fill_2 FILLER_24_1005 ();
 sg13g2_fill_2 FILLER_24_1011 ();
 sg13g2_fill_2 FILLER_24_1018 ();
 sg13g2_fill_1 FILLER_24_1033 ();
 sg13g2_decap_8 FILLER_24_1047 ();
 sg13g2_decap_4 FILLER_24_1054 ();
 sg13g2_decap_8 FILLER_24_1062 ();
 sg13g2_decap_8 FILLER_24_1069 ();
 sg13g2_fill_1 FILLER_24_1076 ();
 sg13g2_fill_2 FILLER_24_1081 ();
 sg13g2_fill_1 FILLER_24_1088 ();
 sg13g2_decap_8 FILLER_24_1093 ();
 sg13g2_decap_8 FILLER_24_1100 ();
 sg13g2_decap_4 FILLER_24_1107 ();
 sg13g2_fill_2 FILLER_24_1129 ();
 sg13g2_decap_8 FILLER_24_1141 ();
 sg13g2_fill_2 FILLER_24_1148 ();
 sg13g2_fill_2 FILLER_24_1165 ();
 sg13g2_fill_1 FILLER_24_1167 ();
 sg13g2_fill_2 FILLER_24_1177 ();
 sg13g2_fill_1 FILLER_24_1200 ();
 sg13g2_fill_2 FILLER_24_1229 ();
 sg13g2_decap_4 FILLER_24_1252 ();
 sg13g2_decap_4 FILLER_24_1265 ();
 sg13g2_fill_2 FILLER_24_1269 ();
 sg13g2_decap_8 FILLER_24_1292 ();
 sg13g2_decap_4 FILLER_24_1299 ();
 sg13g2_fill_2 FILLER_24_1303 ();
 sg13g2_fill_2 FILLER_24_1323 ();
 sg13g2_fill_1 FILLER_24_1325 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_4 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_31 ();
 sg13g2_decap_4 FILLER_25_38 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_2 FILLER_25_48 ();
 sg13g2_fill_1 FILLER_25_50 ();
 sg13g2_fill_1 FILLER_25_55 ();
 sg13g2_decap_4 FILLER_25_63 ();
 sg13g2_decap_4 FILLER_25_70 ();
 sg13g2_fill_1 FILLER_25_74 ();
 sg13g2_fill_1 FILLER_25_87 ();
 sg13g2_fill_2 FILLER_25_93 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_114 ();
 sg13g2_fill_1 FILLER_25_118 ();
 sg13g2_decap_4 FILLER_25_156 ();
 sg13g2_decap_4 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_243 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_296 ();
 sg13g2_decap_8 FILLER_25_303 ();
 sg13g2_decap_8 FILLER_25_310 ();
 sg13g2_decap_8 FILLER_25_317 ();
 sg13g2_fill_2 FILLER_25_324 ();
 sg13g2_fill_1 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_4 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_fill_2 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_4 FILLER_25_436 ();
 sg13g2_fill_2 FILLER_25_440 ();
 sg13g2_decap_8 FILLER_25_463 ();
 sg13g2_decap_4 FILLER_25_470 ();
 sg13g2_fill_1 FILLER_25_474 ();
 sg13g2_fill_2 FILLER_25_479 ();
 sg13g2_fill_1 FILLER_25_481 ();
 sg13g2_decap_4 FILLER_25_496 ();
 sg13g2_fill_2 FILLER_25_500 ();
 sg13g2_fill_2 FILLER_25_513 ();
 sg13g2_fill_1 FILLER_25_515 ();
 sg13g2_decap_8 FILLER_25_519 ();
 sg13g2_decap_8 FILLER_25_526 ();
 sg13g2_fill_2 FILLER_25_533 ();
 sg13g2_fill_1 FILLER_25_535 ();
 sg13g2_decap_8 FILLER_25_541 ();
 sg13g2_decap_8 FILLER_25_548 ();
 sg13g2_fill_1 FILLER_25_564 ();
 sg13g2_decap_4 FILLER_25_578 ();
 sg13g2_fill_2 FILLER_25_603 ();
 sg13g2_fill_2 FILLER_25_628 ();
 sg13g2_fill_1 FILLER_25_630 ();
 sg13g2_fill_2 FILLER_25_640 ();
 sg13g2_fill_2 FILLER_25_653 ();
 sg13g2_decap_4 FILLER_25_688 ();
 sg13g2_fill_2 FILLER_25_692 ();
 sg13g2_decap_8 FILLER_25_699 ();
 sg13g2_decap_8 FILLER_25_706 ();
 sg13g2_decap_4 FILLER_25_713 ();
 sg13g2_fill_2 FILLER_25_721 ();
 sg13g2_fill_1 FILLER_25_723 ();
 sg13g2_decap_8 FILLER_25_727 ();
 sg13g2_decap_8 FILLER_25_734 ();
 sg13g2_fill_2 FILLER_25_741 ();
 sg13g2_fill_1 FILLER_25_747 ();
 sg13g2_fill_1 FILLER_25_754 ();
 sg13g2_decap_8 FILLER_25_760 ();
 sg13g2_fill_2 FILLER_25_767 ();
 sg13g2_decap_8 FILLER_25_775 ();
 sg13g2_decap_8 FILLER_25_782 ();
 sg13g2_decap_8 FILLER_25_789 ();
 sg13g2_fill_2 FILLER_25_796 ();
 sg13g2_decap_8 FILLER_25_801 ();
 sg13g2_decap_4 FILLER_25_808 ();
 sg13g2_fill_1 FILLER_25_812 ();
 sg13g2_fill_2 FILLER_25_817 ();
 sg13g2_decap_8 FILLER_25_845 ();
 sg13g2_fill_2 FILLER_25_852 ();
 sg13g2_fill_1 FILLER_25_854 ();
 sg13g2_decap_4 FILLER_25_858 ();
 sg13g2_fill_2 FILLER_25_874 ();
 sg13g2_decap_8 FILLER_25_900 ();
 sg13g2_fill_1 FILLER_25_907 ();
 sg13g2_fill_1 FILLER_25_939 ();
 sg13g2_fill_1 FILLER_25_957 ();
 sg13g2_fill_1 FILLER_25_966 ();
 sg13g2_decap_8 FILLER_25_975 ();
 sg13g2_decap_4 FILLER_25_982 ();
 sg13g2_decap_4 FILLER_25_1009 ();
 sg13g2_fill_1 FILLER_25_1017 ();
 sg13g2_fill_2 FILLER_25_1069 ();
 sg13g2_fill_1 FILLER_25_1071 ();
 sg13g2_fill_2 FILLER_25_1078 ();
 sg13g2_fill_1 FILLER_25_1080 ();
 sg13g2_decap_8 FILLER_25_1084 ();
 sg13g2_decap_8 FILLER_25_1091 ();
 sg13g2_decap_4 FILLER_25_1098 ();
 sg13g2_fill_2 FILLER_25_1102 ();
 sg13g2_decap_8 FILLER_25_1111 ();
 sg13g2_fill_2 FILLER_25_1118 ();
 sg13g2_fill_1 FILLER_25_1120 ();
 sg13g2_decap_8 FILLER_25_1135 ();
 sg13g2_decap_4 FILLER_25_1180 ();
 sg13g2_fill_2 FILLER_25_1184 ();
 sg13g2_fill_1 FILLER_25_1191 ();
 sg13g2_fill_1 FILLER_25_1196 ();
 sg13g2_fill_1 FILLER_25_1200 ();
 sg13g2_fill_2 FILLER_25_1204 ();
 sg13g2_fill_1 FILLER_25_1211 ();
 sg13g2_fill_1 FILLER_25_1217 ();
 sg13g2_fill_1 FILLER_25_1223 ();
 sg13g2_fill_1 FILLER_25_1228 ();
 sg13g2_decap_8 FILLER_25_1258 ();
 sg13g2_fill_2 FILLER_25_1265 ();
 sg13g2_fill_1 FILLER_25_1267 ();
 sg13g2_fill_2 FILLER_25_1272 ();
 sg13g2_fill_1 FILLER_25_1274 ();
 sg13g2_decap_8 FILLER_25_1292 ();
 sg13g2_decap_4 FILLER_25_1299 ();
 sg13g2_decap_8 FILLER_25_1306 ();
 sg13g2_decap_8 FILLER_25_1316 ();
 sg13g2_fill_2 FILLER_25_1323 ();
 sg13g2_fill_1 FILLER_25_1325 ();
 sg13g2_fill_2 FILLER_26_31 ();
 sg13g2_decap_8 FILLER_26_59 ();
 sg13g2_fill_2 FILLER_26_66 ();
 sg13g2_fill_1 FILLER_26_68 ();
 sg13g2_decap_8 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_84 ();
 sg13g2_decap_4 FILLER_26_100 ();
 sg13g2_decap_4 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_170 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_fill_2 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_221 ();
 sg13g2_decap_4 FILLER_26_240 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_264 ();
 sg13g2_fill_2 FILLER_26_269 ();
 sg13g2_fill_2 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_fill_2 FILLER_26_319 ();
 sg13g2_decap_4 FILLER_26_324 ();
 sg13g2_decap_8 FILLER_26_332 ();
 sg13g2_decap_8 FILLER_26_339 ();
 sg13g2_decap_4 FILLER_26_346 ();
 sg13g2_fill_2 FILLER_26_350 ();
 sg13g2_decap_4 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_370 ();
 sg13g2_fill_1 FILLER_26_372 ();
 sg13g2_fill_2 FILLER_26_378 ();
 sg13g2_fill_1 FILLER_26_380 ();
 sg13g2_fill_1 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_4 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_409 ();
 sg13g2_fill_2 FILLER_26_414 ();
 sg13g2_decap_4 FILLER_26_420 ();
 sg13g2_fill_2 FILLER_26_424 ();
 sg13g2_decap_4 FILLER_26_438 ();
 sg13g2_fill_2 FILLER_26_442 ();
 sg13g2_fill_1 FILLER_26_448 ();
 sg13g2_fill_2 FILLER_26_488 ();
 sg13g2_fill_2 FILLER_26_516 ();
 sg13g2_decap_8 FILLER_26_528 ();
 sg13g2_fill_2 FILLER_26_535 ();
 sg13g2_fill_2 FILLER_26_547 ();
 sg13g2_fill_1 FILLER_26_549 ();
 sg13g2_decap_8 FILLER_26_568 ();
 sg13g2_decap_4 FILLER_26_581 ();
 sg13g2_fill_1 FILLER_26_585 ();
 sg13g2_fill_1 FILLER_26_590 ();
 sg13g2_fill_1 FILLER_26_595 ();
 sg13g2_fill_1 FILLER_26_605 ();
 sg13g2_fill_2 FILLER_26_611 ();
 sg13g2_decap_8 FILLER_26_624 ();
 sg13g2_decap_8 FILLER_26_631 ();
 sg13g2_decap_4 FILLER_26_638 ();
 sg13g2_fill_2 FILLER_26_642 ();
 sg13g2_fill_2 FILLER_26_652 ();
 sg13g2_fill_1 FILLER_26_654 ();
 sg13g2_decap_4 FILLER_26_660 ();
 sg13g2_fill_2 FILLER_26_664 ();
 sg13g2_decap_8 FILLER_26_688 ();
 sg13g2_fill_2 FILLER_26_712 ();
 sg13g2_fill_2 FILLER_26_738 ();
 sg13g2_fill_1 FILLER_26_745 ();
 sg13g2_fill_1 FILLER_26_750 ();
 sg13g2_decap_4 FILLER_26_764 ();
 sg13g2_fill_2 FILLER_26_768 ();
 sg13g2_fill_2 FILLER_26_775 ();
 sg13g2_fill_1 FILLER_26_777 ();
 sg13g2_fill_2 FILLER_26_784 ();
 sg13g2_fill_2 FILLER_26_800 ();
 sg13g2_fill_1 FILLER_26_808 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_fill_2 FILLER_26_831 ();
 sg13g2_fill_2 FILLER_26_836 ();
 sg13g2_decap_4 FILLER_26_845 ();
 sg13g2_fill_2 FILLER_26_857 ();
 sg13g2_fill_1 FILLER_26_877 ();
 sg13g2_fill_1 FILLER_26_892 ();
 sg13g2_fill_1 FILLER_26_902 ();
 sg13g2_fill_2 FILLER_26_910 ();
 sg13g2_fill_1 FILLER_26_921 ();
 sg13g2_fill_2 FILLER_26_936 ();
 sg13g2_fill_2 FILLER_26_941 ();
 sg13g2_decap_4 FILLER_26_957 ();
 sg13g2_fill_1 FILLER_26_961 ();
 sg13g2_decap_4 FILLER_26_968 ();
 sg13g2_fill_1 FILLER_26_984 ();
 sg13g2_fill_2 FILLER_26_1014 ();
 sg13g2_fill_1 FILLER_26_1016 ();
 sg13g2_decap_4 FILLER_26_1024 ();
 sg13g2_decap_8 FILLER_26_1034 ();
 sg13g2_decap_4 FILLER_26_1044 ();
 sg13g2_fill_1 FILLER_26_1048 ();
 sg13g2_decap_8 FILLER_26_1058 ();
 sg13g2_decap_4 FILLER_26_1065 ();
 sg13g2_fill_2 FILLER_26_1073 ();
 sg13g2_decap_4 FILLER_26_1081 ();
 sg13g2_fill_1 FILLER_26_1085 ();
 sg13g2_fill_1 FILLER_26_1092 ();
 sg13g2_decap_8 FILLER_26_1097 ();
 sg13g2_decap_8 FILLER_26_1113 ();
 sg13g2_fill_2 FILLER_26_1120 ();
 sg13g2_decap_8 FILLER_26_1141 ();
 sg13g2_decap_8 FILLER_26_1148 ();
 sg13g2_decap_8 FILLER_26_1159 ();
 sg13g2_decap_4 FILLER_26_1166 ();
 sg13g2_fill_1 FILLER_26_1170 ();
 sg13g2_decap_8 FILLER_26_1177 ();
 sg13g2_fill_1 FILLER_26_1184 ();
 sg13g2_fill_2 FILLER_26_1189 ();
 sg13g2_fill_1 FILLER_26_1200 ();
 sg13g2_fill_1 FILLER_26_1211 ();
 sg13g2_fill_2 FILLER_26_1223 ();
 sg13g2_fill_1 FILLER_26_1325 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_fill_1 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_19 ();
 sg13g2_fill_2 FILLER_27_30 ();
 sg13g2_fill_1 FILLER_27_32 ();
 sg13g2_decap_4 FILLER_27_41 ();
 sg13g2_fill_1 FILLER_27_45 ();
 sg13g2_decap_8 FILLER_27_50 ();
 sg13g2_decap_8 FILLER_27_57 ();
 sg13g2_decap_8 FILLER_27_64 ();
 sg13g2_decap_8 FILLER_27_71 ();
 sg13g2_decap_4 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_92 ();
 sg13g2_fill_1 FILLER_27_102 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_fill_1 FILLER_27_113 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_150 ();
 sg13g2_fill_2 FILLER_27_154 ();
 sg13g2_fill_1 FILLER_27_165 ();
 sg13g2_decap_4 FILLER_27_179 ();
 sg13g2_fill_2 FILLER_27_183 ();
 sg13g2_fill_2 FILLER_27_218 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_decap_4 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_286 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_decap_8 FILLER_27_313 ();
 sg13g2_decap_8 FILLER_27_331 ();
 sg13g2_fill_1 FILLER_27_338 ();
 sg13g2_decap_4 FILLER_27_351 ();
 sg13g2_fill_1 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_fill_2 FILLER_27_375 ();
 sg13g2_fill_1 FILLER_27_382 ();
 sg13g2_fill_2 FILLER_27_393 ();
 sg13g2_fill_1 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_444 ();
 sg13g2_decap_8 FILLER_27_451 ();
 sg13g2_decap_4 FILLER_27_458 ();
 sg13g2_fill_1 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_471 ();
 sg13g2_decap_8 FILLER_27_478 ();
 sg13g2_decap_4 FILLER_27_485 ();
 sg13g2_fill_2 FILLER_27_489 ();
 sg13g2_fill_1 FILLER_27_515 ();
 sg13g2_decap_8 FILLER_27_522 ();
 sg13g2_fill_2 FILLER_27_536 ();
 sg13g2_decap_4 FILLER_27_543 ();
 sg13g2_decap_4 FILLER_27_558 ();
 sg13g2_decap_8 FILLER_27_573 ();
 sg13g2_fill_2 FILLER_27_580 ();
 sg13g2_fill_1 FILLER_27_591 ();
 sg13g2_fill_1 FILLER_27_595 ();
 sg13g2_fill_2 FILLER_27_602 ();
 sg13g2_fill_1 FILLER_27_607 ();
 sg13g2_fill_1 FILLER_27_613 ();
 sg13g2_fill_1 FILLER_27_617 ();
 sg13g2_decap_8 FILLER_27_622 ();
 sg13g2_fill_2 FILLER_27_634 ();
 sg13g2_fill_1 FILLER_27_640 ();
 sg13g2_decap_4 FILLER_27_644 ();
 sg13g2_fill_2 FILLER_27_648 ();
 sg13g2_decap_8 FILLER_27_689 ();
 sg13g2_decap_4 FILLER_27_696 ();
 sg13g2_fill_2 FILLER_27_713 ();
 sg13g2_fill_1 FILLER_27_715 ();
 sg13g2_fill_2 FILLER_27_719 ();
 sg13g2_decap_8 FILLER_27_739 ();
 sg13g2_fill_1 FILLER_27_746 ();
 sg13g2_decap_8 FILLER_27_751 ();
 sg13g2_fill_2 FILLER_27_758 ();
 sg13g2_fill_1 FILLER_27_760 ();
 sg13g2_decap_8 FILLER_27_765 ();
 sg13g2_fill_1 FILLER_27_772 ();
 sg13g2_fill_1 FILLER_27_781 ();
 sg13g2_fill_1 FILLER_27_791 ();
 sg13g2_fill_1 FILLER_27_802 ();
 sg13g2_fill_1 FILLER_27_812 ();
 sg13g2_fill_1 FILLER_27_821 ();
 sg13g2_fill_2 FILLER_27_826 ();
 sg13g2_fill_1 FILLER_27_847 ();
 sg13g2_fill_1 FILLER_27_852 ();
 sg13g2_decap_4 FILLER_27_858 ();
 sg13g2_fill_2 FILLER_27_866 ();
 sg13g2_fill_1 FILLER_27_868 ();
 sg13g2_fill_2 FILLER_27_878 ();
 sg13g2_decap_4 FILLER_27_903 ();
 sg13g2_fill_1 FILLER_27_907 ();
 sg13g2_fill_2 FILLER_27_926 ();
 sg13g2_decap_4 FILLER_27_949 ();
 sg13g2_fill_1 FILLER_27_953 ();
 sg13g2_fill_2 FILLER_27_983 ();
 sg13g2_fill_1 FILLER_27_985 ();
 sg13g2_fill_2 FILLER_27_1003 ();
 sg13g2_fill_1 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1014 ();
 sg13g2_decap_8 FILLER_27_1021 ();
 sg13g2_decap_8 FILLER_27_1028 ();
 sg13g2_fill_2 FILLER_27_1040 ();
 sg13g2_fill_1 FILLER_27_1042 ();
 sg13g2_fill_1 FILLER_27_1053 ();
 sg13g2_fill_1 FILLER_27_1062 ();
 sg13g2_fill_1 FILLER_27_1068 ();
 sg13g2_fill_2 FILLER_27_1073 ();
 sg13g2_fill_2 FILLER_27_1107 ();
 sg13g2_decap_8 FILLER_27_1113 ();
 sg13g2_decap_4 FILLER_27_1120 ();
 sg13g2_fill_2 FILLER_27_1124 ();
 sg13g2_decap_8 FILLER_27_1131 ();
 sg13g2_decap_8 FILLER_27_1138 ();
 sg13g2_decap_8 FILLER_27_1145 ();
 sg13g2_decap_8 FILLER_27_1152 ();
 sg13g2_decap_4 FILLER_27_1159 ();
 sg13g2_decap_8 FILLER_27_1170 ();
 sg13g2_decap_8 FILLER_27_1177 ();
 sg13g2_decap_8 FILLER_27_1184 ();
 sg13g2_fill_1 FILLER_27_1214 ();
 sg13g2_fill_2 FILLER_27_1225 ();
 sg13g2_fill_1 FILLER_27_1250 ();
 sg13g2_decap_8 FILLER_27_1255 ();
 sg13g2_decap_8 FILLER_27_1262 ();
 sg13g2_fill_1 FILLER_27_1275 ();
 sg13g2_decap_4 FILLER_27_1284 ();
 sg13g2_fill_2 FILLER_27_1288 ();
 sg13g2_decap_4 FILLER_27_1294 ();
 sg13g2_fill_2 FILLER_27_1298 ();
 sg13g2_decap_4 FILLER_27_1304 ();
 sg13g2_fill_1 FILLER_27_1308 ();
 sg13g2_decap_8 FILLER_27_1314 ();
 sg13g2_decap_4 FILLER_27_1321 ();
 sg13g2_fill_1 FILLER_27_1325 ();
 sg13g2_fill_1 FILLER_28_26 ();
 sg13g2_decap_4 FILLER_28_53 ();
 sg13g2_decap_4 FILLER_28_83 ();
 sg13g2_fill_2 FILLER_28_87 ();
 sg13g2_decap_8 FILLER_28_96 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_110 ();
 sg13g2_decap_4 FILLER_28_117 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_137 ();
 sg13g2_fill_2 FILLER_28_147 ();
 sg13g2_fill_2 FILLER_28_164 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_fill_1 FILLER_28_186 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_2 FILLER_28_225 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_decap_4 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_237 ();
 sg13g2_decap_4 FILLER_28_246 ();
 sg13g2_fill_1 FILLER_28_260 ();
 sg13g2_fill_1 FILLER_28_264 ();
 sg13g2_fill_1 FILLER_28_276 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_fill_2 FILLER_28_299 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_decap_4 FILLER_28_319 ();
 sg13g2_fill_1 FILLER_28_323 ();
 sg13g2_decap_8 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_decap_4 FILLER_28_343 ();
 sg13g2_decap_4 FILLER_28_355 ();
 sg13g2_fill_1 FILLER_28_376 ();
 sg13g2_decap_4 FILLER_28_396 ();
 sg13g2_fill_2 FILLER_28_417 ();
 sg13g2_fill_2 FILLER_28_424 ();
 sg13g2_fill_1 FILLER_28_426 ();
 sg13g2_fill_1 FILLER_28_447 ();
 sg13g2_decap_4 FILLER_28_456 ();
 sg13g2_fill_2 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_487 ();
 sg13g2_fill_2 FILLER_28_494 ();
 sg13g2_fill_1 FILLER_28_496 ();
 sg13g2_fill_2 FILLER_28_501 ();
 sg13g2_decap_8 FILLER_28_521 ();
 sg13g2_decap_4 FILLER_28_535 ();
 sg13g2_decap_4 FILLER_28_543 ();
 sg13g2_fill_1 FILLER_28_547 ();
 sg13g2_fill_1 FILLER_28_552 ();
 sg13g2_decap_4 FILLER_28_559 ();
 sg13g2_fill_2 FILLER_28_563 ();
 sg13g2_fill_2 FILLER_28_573 ();
 sg13g2_decap_8 FILLER_28_589 ();
 sg13g2_decap_8 FILLER_28_596 ();
 sg13g2_fill_2 FILLER_28_617 ();
 sg13g2_fill_1 FILLER_28_619 ();
 sg13g2_decap_8 FILLER_28_623 ();
 sg13g2_decap_4 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_657 ();
 sg13g2_fill_1 FILLER_28_664 ();
 sg13g2_fill_2 FILLER_28_676 ();
 sg13g2_fill_1 FILLER_28_678 ();
 sg13g2_fill_2 FILLER_28_682 ();
 sg13g2_fill_1 FILLER_28_684 ();
 sg13g2_decap_8 FILLER_28_688 ();
 sg13g2_decap_8 FILLER_28_695 ();
 sg13g2_decap_8 FILLER_28_702 ();
 sg13g2_decap_4 FILLER_28_709 ();
 sg13g2_fill_1 FILLER_28_726 ();
 sg13g2_fill_2 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_4 FILLER_28_749 ();
 sg13g2_decap_4 FILLER_28_766 ();
 sg13g2_fill_2 FILLER_28_817 ();
 sg13g2_decap_8 FILLER_28_832 ();
 sg13g2_decap_4 FILLER_28_839 ();
 sg13g2_decap_8 FILLER_28_850 ();
 sg13g2_fill_2 FILLER_28_857 ();
 sg13g2_decap_8 FILLER_28_875 ();
 sg13g2_decap_4 FILLER_28_882 ();
 sg13g2_decap_8 FILLER_28_894 ();
 sg13g2_decap_4 FILLER_28_901 ();
 sg13g2_decap_8 FILLER_28_919 ();
 sg13g2_fill_2 FILLER_28_926 ();
 sg13g2_fill_1 FILLER_28_928 ();
 sg13g2_decap_4 FILLER_28_942 ();
 sg13g2_decap_8 FILLER_28_951 ();
 sg13g2_fill_2 FILLER_28_962 ();
 sg13g2_fill_2 FILLER_28_967 ();
 sg13g2_fill_1 FILLER_28_969 ();
 sg13g2_fill_1 FILLER_28_977 ();
 sg13g2_decap_8 FILLER_28_981 ();
 sg13g2_fill_1 FILLER_28_988 ();
 sg13g2_fill_2 FILLER_28_992 ();
 sg13g2_fill_1 FILLER_28_994 ();
 sg13g2_decap_4 FILLER_28_1018 ();
 sg13g2_fill_2 FILLER_28_1022 ();
 sg13g2_decap_8 FILLER_28_1027 ();
 sg13g2_fill_1 FILLER_28_1034 ();
 sg13g2_decap_8 FILLER_28_1040 ();
 sg13g2_fill_2 FILLER_28_1047 ();
 sg13g2_fill_1 FILLER_28_1049 ();
 sg13g2_fill_1 FILLER_28_1065 ();
 sg13g2_fill_2 FILLER_28_1075 ();
 sg13g2_decap_8 FILLER_28_1080 ();
 sg13g2_decap_4 FILLER_28_1087 ();
 sg13g2_fill_1 FILLER_28_1099 ();
 sg13g2_fill_2 FILLER_28_1119 ();
 sg13g2_fill_1 FILLER_28_1126 ();
 sg13g2_decap_8 FILLER_28_1132 ();
 sg13g2_decap_8 FILLER_28_1139 ();
 sg13g2_fill_1 FILLER_28_1146 ();
 sg13g2_fill_1 FILLER_28_1159 ();
 sg13g2_fill_1 FILLER_28_1164 ();
 sg13g2_fill_2 FILLER_28_1179 ();
 sg13g2_fill_1 FILLER_28_1181 ();
 sg13g2_fill_2 FILLER_28_1195 ();
 sg13g2_fill_2 FILLER_28_1203 ();
 sg13g2_fill_2 FILLER_28_1230 ();
 sg13g2_fill_1 FILLER_28_1245 ();
 sg13g2_fill_1 FILLER_28_1250 ();
 sg13g2_fill_1 FILLER_28_1264 ();
 sg13g2_decap_8 FILLER_28_1317 ();
 sg13g2_fill_2 FILLER_28_1324 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_4 FILLER_29_47 ();
 sg13g2_decap_4 FILLER_29_60 ();
 sg13g2_decap_4 FILLER_29_72 ();
 sg13g2_fill_2 FILLER_29_76 ();
 sg13g2_decap_8 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_122 ();
 sg13g2_decap_8 FILLER_29_136 ();
 sg13g2_decap_4 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_150 ();
 sg13g2_decap_4 FILLER_29_157 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_165 ();
 sg13g2_fill_1 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_179 ();
 sg13g2_decap_8 FILLER_29_187 ();
 sg13g2_fill_2 FILLER_29_194 ();
 sg13g2_decap_4 FILLER_29_203 ();
 sg13g2_fill_2 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_212 ();
 sg13g2_decap_4 FILLER_29_219 ();
 sg13g2_fill_1 FILLER_29_231 ();
 sg13g2_fill_2 FILLER_29_237 ();
 sg13g2_decap_4 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_261 ();
 sg13g2_decap_4 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_fill_2 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_293 ();
 sg13g2_fill_2 FILLER_29_303 ();
 sg13g2_decap_4 FILLER_29_311 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_353 ();
 sg13g2_fill_2 FILLER_29_388 ();
 sg13g2_fill_1 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_401 ();
 sg13g2_fill_2 FILLER_29_411 ();
 sg13g2_fill_2 FILLER_29_454 ();
 sg13g2_fill_1 FILLER_29_456 ();
 sg13g2_fill_2 FILLER_29_462 ();
 sg13g2_fill_1 FILLER_29_464 ();
 sg13g2_fill_1 FILLER_29_469 ();
 sg13g2_fill_2 FILLER_29_479 ();
 sg13g2_fill_1 FILLER_29_481 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_fill_2 FILLER_29_518 ();
 sg13g2_fill_1 FILLER_29_520 ();
 sg13g2_decap_8 FILLER_29_530 ();
 sg13g2_decap_4 FILLER_29_537 ();
 sg13g2_fill_1 FILLER_29_541 ();
 sg13g2_fill_2 FILLER_29_545 ();
 sg13g2_fill_1 FILLER_29_547 ();
 sg13g2_decap_4 FILLER_29_560 ();
 sg13g2_fill_1 FILLER_29_564 ();
 sg13g2_decap_4 FILLER_29_569 ();
 sg13g2_fill_2 FILLER_29_577 ();
 sg13g2_fill_1 FILLER_29_584 ();
 sg13g2_fill_2 FILLER_29_588 ();
 sg13g2_fill_2 FILLER_29_593 ();
 sg13g2_fill_2 FILLER_29_632 ();
 sg13g2_fill_2 FILLER_29_638 ();
 sg13g2_fill_1 FILLER_29_640 ();
 sg13g2_fill_1 FILLER_29_645 ();
 sg13g2_fill_2 FILLER_29_652 ();
 sg13g2_decap_8 FILLER_29_678 ();
 sg13g2_decap_8 FILLER_29_685 ();
 sg13g2_fill_2 FILLER_29_692 ();
 sg13g2_decap_8 FILLER_29_702 ();
 sg13g2_decap_8 FILLER_29_709 ();
 sg13g2_fill_2 FILLER_29_716 ();
 sg13g2_decap_4 FILLER_29_736 ();
 sg13g2_fill_1 FILLER_29_740 ();
 sg13g2_decap_4 FILLER_29_803 ();
 sg13g2_fill_2 FILLER_29_807 ();
 sg13g2_decap_4 FILLER_29_818 ();
 sg13g2_fill_2 FILLER_29_825 ();
 sg13g2_fill_2 FILLER_29_836 ();
 sg13g2_fill_1 FILLER_29_838 ();
 sg13g2_fill_2 FILLER_29_843 ();
 sg13g2_decap_8 FILLER_29_854 ();
 sg13g2_fill_1 FILLER_29_861 ();
 sg13g2_fill_1 FILLER_29_876 ();
 sg13g2_fill_2 FILLER_29_897 ();
 sg13g2_decap_4 FILLER_29_903 ();
 sg13g2_fill_1 FILLER_29_907 ();
 sg13g2_fill_2 FILLER_29_922 ();
 sg13g2_fill_1 FILLER_29_924 ();
 sg13g2_fill_2 FILLER_29_929 ();
 sg13g2_fill_1 FILLER_29_931 ();
 sg13g2_decap_8 FILLER_29_943 ();
 sg13g2_decap_8 FILLER_29_950 ();
 sg13g2_decap_4 FILLER_29_957 ();
 sg13g2_fill_2 FILLER_29_961 ();
 sg13g2_fill_2 FILLER_29_968 ();
 sg13g2_fill_1 FILLER_29_970 ();
 sg13g2_fill_1 FILLER_29_977 ();
 sg13g2_fill_2 FILLER_29_983 ();
 sg13g2_fill_1 FILLER_29_985 ();
 sg13g2_fill_1 FILLER_29_991 ();
 sg13g2_fill_2 FILLER_29_997 ();
 sg13g2_fill_2 FILLER_29_1002 ();
 sg13g2_fill_2 FILLER_29_1009 ();
 sg13g2_fill_2 FILLER_29_1015 ();
 sg13g2_fill_1 FILLER_29_1017 ();
 sg13g2_fill_2 FILLER_29_1023 ();
 sg13g2_fill_1 FILLER_29_1025 ();
 sg13g2_fill_1 FILLER_29_1057 ();
 sg13g2_fill_2 FILLER_29_1061 ();
 sg13g2_decap_4 FILLER_29_1083 ();
 sg13g2_fill_2 FILLER_29_1092 ();
 sg13g2_fill_1 FILLER_29_1094 ();
 sg13g2_decap_8 FILLER_29_1098 ();
 sg13g2_decap_4 FILLER_29_1105 ();
 sg13g2_fill_1 FILLER_29_1114 ();
 sg13g2_fill_1 FILLER_29_1119 ();
 sg13g2_fill_1 FILLER_29_1133 ();
 sg13g2_fill_2 FILLER_29_1142 ();
 sg13g2_fill_2 FILLER_29_1153 ();
 sg13g2_fill_2 FILLER_29_1168 ();
 sg13g2_fill_1 FILLER_29_1170 ();
 sg13g2_fill_2 FILLER_29_1184 ();
 sg13g2_fill_1 FILLER_29_1186 ();
 sg13g2_decap_8 FILLER_29_1191 ();
 sg13g2_fill_2 FILLER_29_1198 ();
 sg13g2_fill_1 FILLER_29_1250 ();
 sg13g2_fill_2 FILLER_29_1257 ();
 sg13g2_fill_1 FILLER_29_1285 ();
 sg13g2_decap_8 FILLER_29_1294 ();
 sg13g2_decap_8 FILLER_29_1301 ();
 sg13g2_decap_4 FILLER_29_1308 ();
 sg13g2_fill_1 FILLER_29_1312 ();
 sg13g2_decap_4 FILLER_29_1322 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_21 ();
 sg13g2_fill_1 FILLER_30_23 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_46 ();
 sg13g2_fill_2 FILLER_30_57 ();
 sg13g2_fill_1 FILLER_30_59 ();
 sg13g2_decap_4 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_86 ();
 sg13g2_decap_4 FILLER_30_96 ();
 sg13g2_fill_2 FILLER_30_100 ();
 sg13g2_fill_2 FILLER_30_154 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_185 ();
 sg13g2_fill_1 FILLER_30_216 ();
 sg13g2_fill_1 FILLER_30_222 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_fill_2 FILLER_30_245 ();
 sg13g2_fill_1 FILLER_30_247 ();
 sg13g2_decap_8 FILLER_30_256 ();
 sg13g2_fill_2 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_decap_8 FILLER_30_281 ();
 sg13g2_decap_4 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_300 ();
 sg13g2_fill_1 FILLER_30_307 ();
 sg13g2_decap_8 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_327 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_fill_2 FILLER_30_338 ();
 sg13g2_fill_2 FILLER_30_344 ();
 sg13g2_fill_2 FILLER_30_355 ();
 sg13g2_fill_2 FILLER_30_370 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_decap_4 FILLER_30_390 ();
 sg13g2_fill_2 FILLER_30_394 ();
 sg13g2_fill_2 FILLER_30_405 ();
 sg13g2_fill_2 FILLER_30_421 ();
 sg13g2_fill_1 FILLER_30_440 ();
 sg13g2_decap_4 FILLER_30_446 ();
 sg13g2_fill_2 FILLER_30_450 ();
 sg13g2_fill_2 FILLER_30_456 ();
 sg13g2_fill_1 FILLER_30_458 ();
 sg13g2_decap_8 FILLER_30_465 ();
 sg13g2_decap_4 FILLER_30_472 ();
 sg13g2_decap_8 FILLER_30_489 ();
 sg13g2_decap_4 FILLER_30_496 ();
 sg13g2_fill_2 FILLER_30_500 ();
 sg13g2_decap_4 FILLER_30_516 ();
 sg13g2_fill_1 FILLER_30_520 ();
 sg13g2_decap_4 FILLER_30_547 ();
 sg13g2_fill_2 FILLER_30_563 ();
 sg13g2_fill_1 FILLER_30_576 ();
 sg13g2_decap_4 FILLER_30_587 ();
 sg13g2_fill_1 FILLER_30_591 ();
 sg13g2_fill_2 FILLER_30_600 ();
 sg13g2_fill_1 FILLER_30_619 ();
 sg13g2_fill_1 FILLER_30_631 ();
 sg13g2_fill_1 FILLER_30_638 ();
 sg13g2_fill_1 FILLER_30_653 ();
 sg13g2_fill_1 FILLER_30_659 ();
 sg13g2_decap_8 FILLER_30_673 ();
 sg13g2_decap_8 FILLER_30_680 ();
 sg13g2_decap_8 FILLER_30_687 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_4 FILLER_30_739 ();
 sg13g2_fill_1 FILLER_30_743 ();
 sg13g2_fill_1 FILLER_30_757 ();
 sg13g2_fill_2 FILLER_30_770 ();
 sg13g2_fill_1 FILLER_30_779 ();
 sg13g2_fill_1 FILLER_30_785 ();
 sg13g2_fill_2 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_810 ();
 sg13g2_fill_1 FILLER_30_817 ();
 sg13g2_fill_1 FILLER_30_822 ();
 sg13g2_fill_2 FILLER_30_833 ();
 sg13g2_fill_2 FILLER_30_838 ();
 sg13g2_decap_4 FILLER_30_848 ();
 sg13g2_fill_1 FILLER_30_855 ();
 sg13g2_fill_1 FILLER_30_874 ();
 sg13g2_fill_2 FILLER_30_881 ();
 sg13g2_fill_1 FILLER_30_883 ();
 sg13g2_decap_8 FILLER_30_888 ();
 sg13g2_fill_1 FILLER_30_895 ();
 sg13g2_fill_2 FILLER_30_901 ();
 sg13g2_fill_2 FILLER_30_907 ();
 sg13g2_fill_1 FILLER_30_909 ();
 sg13g2_decap_8 FILLER_30_939 ();
 sg13g2_fill_2 FILLER_30_946 ();
 sg13g2_decap_8 FILLER_30_957 ();
 sg13g2_decap_4 FILLER_30_964 ();
 sg13g2_fill_2 FILLER_30_968 ();
 sg13g2_decap_4 FILLER_30_978 ();
 sg13g2_fill_1 FILLER_30_982 ();
 sg13g2_decap_8 FILLER_30_994 ();
 sg13g2_decap_8 FILLER_30_1001 ();
 sg13g2_fill_1 FILLER_30_1008 ();
 sg13g2_decap_8 FILLER_30_1013 ();
 sg13g2_decap_8 FILLER_30_1020 ();
 sg13g2_decap_4 FILLER_30_1027 ();
 sg13g2_fill_1 FILLER_30_1031 ();
 sg13g2_fill_1 FILLER_30_1048 ();
 sg13g2_fill_1 FILLER_30_1068 ();
 sg13g2_fill_2 FILLER_30_1073 ();
 sg13g2_fill_1 FILLER_30_1075 ();
 sg13g2_fill_2 FILLER_30_1081 ();
 sg13g2_fill_1 FILLER_30_1083 ();
 sg13g2_fill_2 FILLER_30_1089 ();
 sg13g2_fill_1 FILLER_30_1091 ();
 sg13g2_fill_1 FILLER_30_1099 ();
 sg13g2_decap_4 FILLER_30_1104 ();
 sg13g2_fill_1 FILLER_30_1115 ();
 sg13g2_fill_2 FILLER_30_1124 ();
 sg13g2_decap_4 FILLER_30_1131 ();
 sg13g2_fill_2 FILLER_30_1144 ();
 sg13g2_fill_1 FILLER_30_1146 ();
 sg13g2_fill_2 FILLER_30_1171 ();
 sg13g2_fill_2 FILLER_30_1178 ();
 sg13g2_fill_1 FILLER_30_1180 ();
 sg13g2_decap_4 FILLER_30_1187 ();
 sg13g2_fill_2 FILLER_30_1191 ();
 sg13g2_fill_1 FILLER_30_1197 ();
 sg13g2_fill_2 FILLER_30_1217 ();
 sg13g2_fill_1 FILLER_30_1228 ();
 sg13g2_fill_2 FILLER_30_1242 ();
 sg13g2_fill_1 FILLER_30_1252 ();
 sg13g2_fill_2 FILLER_30_1262 ();
 sg13g2_decap_4 FILLER_30_1277 ();
 sg13g2_fill_1 FILLER_30_1281 ();
 sg13g2_fill_2 FILLER_30_1286 ();
 sg13g2_fill_1 FILLER_30_1288 ();
 sg13g2_decap_4 FILLER_30_1293 ();
 sg13g2_decap_4 FILLER_30_1301 ();
 sg13g2_fill_1 FILLER_30_1305 ();
 sg13g2_decap_4 FILLER_30_1320 ();
 sg13g2_fill_2 FILLER_30_1324 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_27 ();
 sg13g2_fill_2 FILLER_31_54 ();
 sg13g2_fill_2 FILLER_31_60 ();
 sg13g2_decap_8 FILLER_31_73 ();
 sg13g2_decap_4 FILLER_31_88 ();
 sg13g2_fill_2 FILLER_31_102 ();
 sg13g2_fill_1 FILLER_31_119 ();
 sg13g2_fill_2 FILLER_31_145 ();
 sg13g2_decap_4 FILLER_31_151 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_176 ();
 sg13g2_decap_8 FILLER_31_181 ();
 sg13g2_decap_8 FILLER_31_188 ();
 sg13g2_fill_2 FILLER_31_195 ();
 sg13g2_fill_2 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_207 ();
 sg13g2_decap_8 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_224 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_248 ();
 sg13g2_fill_2 FILLER_31_258 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_fill_2 FILLER_31_281 ();
 sg13g2_fill_2 FILLER_31_288 ();
 sg13g2_fill_2 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_decap_4 FILLER_31_314 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_fill_2 FILLER_31_329 ();
 sg13g2_fill_1 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_decap_4 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_385 ();
 sg13g2_fill_1 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_416 ();
 sg13g2_fill_2 FILLER_31_453 ();
 sg13g2_fill_1 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_fill_1 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_485 ();
 sg13g2_decap_8 FILLER_31_492 ();
 sg13g2_fill_2 FILLER_31_499 ();
 sg13g2_decap_8 FILLER_31_509 ();
 sg13g2_fill_1 FILLER_31_516 ();
 sg13g2_fill_1 FILLER_31_522 ();
 sg13g2_decap_8 FILLER_31_527 ();
 sg13g2_decap_8 FILLER_31_534 ();
 sg13g2_decap_4 FILLER_31_546 ();
 sg13g2_fill_1 FILLER_31_560 ();
 sg13g2_fill_1 FILLER_31_564 ();
 sg13g2_fill_2 FILLER_31_573 ();
 sg13g2_fill_1 FILLER_31_580 ();
 sg13g2_decap_8 FILLER_31_597 ();
 sg13g2_fill_1 FILLER_31_604 ();
 sg13g2_decap_4 FILLER_31_610 ();
 sg13g2_fill_1 FILLER_31_614 ();
 sg13g2_fill_1 FILLER_31_626 ();
 sg13g2_fill_1 FILLER_31_648 ();
 sg13g2_fill_2 FILLER_31_652 ();
 sg13g2_fill_1 FILLER_31_670 ();
 sg13g2_decap_8 FILLER_31_706 ();
 sg13g2_decap_8 FILLER_31_713 ();
 sg13g2_decap_4 FILLER_31_720 ();
 sg13g2_fill_2 FILLER_31_724 ();
 sg13g2_fill_1 FILLER_31_731 ();
 sg13g2_decap_4 FILLER_31_740 ();
 sg13g2_fill_2 FILLER_31_744 ();
 sg13g2_decap_4 FILLER_31_754 ();
 sg13g2_fill_2 FILLER_31_758 ();
 sg13g2_fill_1 FILLER_31_768 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_fill_2 FILLER_31_835 ();
 sg13g2_fill_1 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_31_867 ();
 sg13g2_fill_2 FILLER_31_877 ();
 sg13g2_fill_2 FILLER_31_883 ();
 sg13g2_decap_8 FILLER_31_890 ();
 sg13g2_decap_8 FILLER_31_902 ();
 sg13g2_decap_4 FILLER_31_909 ();
 sg13g2_fill_2 FILLER_31_920 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_4 FILLER_31_952 ();
 sg13g2_decap_8 FILLER_31_961 ();
 sg13g2_fill_2 FILLER_31_968 ();
 sg13g2_decap_4 FILLER_31_976 ();
 sg13g2_fill_2 FILLER_31_988 ();
 sg13g2_decap_8 FILLER_31_993 ();
 sg13g2_decap_8 FILLER_31_1000 ();
 sg13g2_decap_8 FILLER_31_1007 ();
 sg13g2_decap_8 FILLER_31_1014 ();
 sg13g2_decap_8 FILLER_31_1021 ();
 sg13g2_decap_8 FILLER_31_1028 ();
 sg13g2_decap_4 FILLER_31_1035 ();
 sg13g2_fill_1 FILLER_31_1039 ();
 sg13g2_decap_8 FILLER_31_1044 ();
 sg13g2_decap_8 FILLER_31_1051 ();
 sg13g2_decap_8 FILLER_31_1058 ();
 sg13g2_decap_8 FILLER_31_1069 ();
 sg13g2_decap_4 FILLER_31_1076 ();
 sg13g2_decap_4 FILLER_31_1084 ();
 sg13g2_decap_4 FILLER_31_1092 ();
 sg13g2_fill_2 FILLER_31_1096 ();
 sg13g2_decap_8 FILLER_31_1106 ();
 sg13g2_decap_8 FILLER_31_1113 ();
 sg13g2_decap_8 FILLER_31_1120 ();
 sg13g2_decap_4 FILLER_31_1130 ();
 sg13g2_fill_2 FILLER_31_1134 ();
 sg13g2_fill_1 FILLER_31_1173 ();
 sg13g2_decap_4 FILLER_31_1183 ();
 sg13g2_fill_1 FILLER_31_1187 ();
 sg13g2_decap_8 FILLER_31_1202 ();
 sg13g2_fill_2 FILLER_31_1209 ();
 sg13g2_fill_1 FILLER_31_1211 ();
 sg13g2_fill_1 FILLER_31_1230 ();
 sg13g2_decap_8 FILLER_31_1240 ();
 sg13g2_fill_2 FILLER_31_1250 ();
 sg13g2_fill_1 FILLER_31_1252 ();
 sg13g2_decap_8 FILLER_31_1257 ();
 sg13g2_decap_8 FILLER_31_1264 ();
 sg13g2_decap_8 FILLER_31_1271 ();
 sg13g2_decap_4 FILLER_31_1278 ();
 sg13g2_fill_2 FILLER_31_1282 ();
 sg13g2_decap_8 FILLER_31_1288 ();
 sg13g2_fill_1 FILLER_31_1295 ();
 sg13g2_fill_2 FILLER_31_1304 ();
 sg13g2_fill_1 FILLER_31_1306 ();
 sg13g2_fill_2 FILLER_31_1312 ();
 sg13g2_fill_2 FILLER_31_1323 ();
 sg13g2_fill_1 FILLER_31_1325 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_decap_4 FILLER_32_25 ();
 sg13g2_fill_1 FILLER_32_29 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_75 ();
 sg13g2_decap_4 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_84 ();
 sg13g2_fill_1 FILLER_32_89 ();
 sg13g2_decap_4 FILLER_32_102 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_fill_2 FILLER_32_122 ();
 sg13g2_fill_1 FILLER_32_129 ();
 sg13g2_fill_2 FILLER_32_146 ();
 sg13g2_fill_1 FILLER_32_148 ();
 sg13g2_fill_2 FILLER_32_186 ();
 sg13g2_decap_4 FILLER_32_192 ();
 sg13g2_fill_1 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_238 ();
 sg13g2_decap_4 FILLER_32_244 ();
 sg13g2_fill_1 FILLER_32_252 ();
 sg13g2_decap_4 FILLER_32_258 ();
 sg13g2_decap_4 FILLER_32_265 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_2 FILLER_32_276 ();
 sg13g2_decap_8 FILLER_32_293 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_fill_2 FILLER_32_313 ();
 sg13g2_decap_4 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_fill_1 FILLER_32_335 ();
 sg13g2_fill_1 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_345 ();
 sg13g2_decap_8 FILLER_32_352 ();
 sg13g2_fill_2 FILLER_32_359 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_decap_4 FILLER_32_387 ();
 sg13g2_fill_2 FILLER_32_391 ();
 sg13g2_fill_2 FILLER_32_404 ();
 sg13g2_decap_4 FILLER_32_411 ();
 sg13g2_fill_2 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_421 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_fill_1 FILLER_32_430 ();
 sg13g2_decap_4 FILLER_32_454 ();
 sg13g2_fill_2 FILLER_32_458 ();
 sg13g2_decap_8 FILLER_32_464 ();
 sg13g2_fill_2 FILLER_32_471 ();
 sg13g2_decap_4 FILLER_32_490 ();
 sg13g2_fill_1 FILLER_32_507 ();
 sg13g2_fill_1 FILLER_32_512 ();
 sg13g2_fill_1 FILLER_32_539 ();
 sg13g2_fill_1 FILLER_32_544 ();
 sg13g2_fill_1 FILLER_32_550 ();
 sg13g2_fill_2 FILLER_32_555 ();
 sg13g2_decap_8 FILLER_32_573 ();
 sg13g2_fill_1 FILLER_32_588 ();
 sg13g2_fill_1 FILLER_32_592 ();
 sg13g2_fill_1 FILLER_32_596 ();
 sg13g2_fill_1 FILLER_32_602 ();
 sg13g2_fill_2 FILLER_32_607 ();
 sg13g2_fill_2 FILLER_32_620 ();
 sg13g2_fill_1 FILLER_32_626 ();
 sg13g2_fill_2 FILLER_32_642 ();
 sg13g2_fill_1 FILLER_32_654 ();
 sg13g2_fill_2 FILLER_32_674 ();
 sg13g2_fill_1 FILLER_32_676 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_4 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_701 ();
 sg13g2_decap_8 FILLER_32_708 ();
 sg13g2_decap_8 FILLER_32_733 ();
 sg13g2_fill_2 FILLER_32_740 ();
 sg13g2_fill_2 FILLER_32_745 ();
 sg13g2_fill_1 FILLER_32_754 ();
 sg13g2_fill_2 FILLER_32_759 ();
 sg13g2_fill_1 FILLER_32_761 ();
 sg13g2_fill_2 FILLER_32_766 ();
 sg13g2_fill_1 FILLER_32_768 ();
 sg13g2_fill_2 FILLER_32_783 ();
 sg13g2_fill_2 FILLER_32_795 ();
 sg13g2_fill_1 FILLER_32_802 ();
 sg13g2_fill_1 FILLER_32_807 ();
 sg13g2_fill_1 FILLER_32_813 ();
 sg13g2_fill_1 FILLER_32_820 ();
 sg13g2_fill_1 FILLER_32_824 ();
 sg13g2_fill_2 FILLER_32_836 ();
 sg13g2_decap_4 FILLER_32_841 ();
 sg13g2_fill_1 FILLER_32_845 ();
 sg13g2_decap_8 FILLER_32_867 ();
 sg13g2_decap_8 FILLER_32_878 ();
 sg13g2_decap_4 FILLER_32_885 ();
 sg13g2_fill_2 FILLER_32_889 ();
 sg13g2_fill_1 FILLER_32_898 ();
 sg13g2_fill_2 FILLER_32_902 ();
 sg13g2_fill_1 FILLER_32_912 ();
 sg13g2_fill_2 FILLER_32_921 ();
 sg13g2_decap_4 FILLER_32_932 ();
 sg13g2_fill_2 FILLER_32_936 ();
 sg13g2_fill_2 FILLER_32_943 ();
 sg13g2_fill_1 FILLER_32_945 ();
 sg13g2_fill_1 FILLER_32_955 ();
 sg13g2_fill_1 FILLER_32_960 ();
 sg13g2_fill_1 FILLER_32_964 ();
 sg13g2_fill_2 FILLER_32_973 ();
 sg13g2_fill_2 FILLER_32_998 ();
 sg13g2_fill_1 FILLER_32_1009 ();
 sg13g2_fill_1 FILLER_32_1014 ();
 sg13g2_decap_8 FILLER_32_1025 ();
 sg13g2_fill_2 FILLER_32_1032 ();
 sg13g2_decap_8 FILLER_32_1051 ();
 sg13g2_fill_1 FILLER_32_1058 ();
 sg13g2_decap_8 FILLER_32_1062 ();
 sg13g2_fill_1 FILLER_32_1069 ();
 sg13g2_decap_4 FILLER_32_1075 ();
 sg13g2_decap_8 FILLER_32_1086 ();
 sg13g2_fill_2 FILLER_32_1093 ();
 sg13g2_fill_1 FILLER_32_1095 ();
 sg13g2_decap_4 FILLER_32_1100 ();
 sg13g2_fill_1 FILLER_32_1104 ();
 sg13g2_decap_4 FILLER_32_1112 ();
 sg13g2_decap_8 FILLER_32_1121 ();
 sg13g2_decap_4 FILLER_32_1128 ();
 sg13g2_decap_8 FILLER_32_1137 ();
 sg13g2_decap_8 FILLER_32_1144 ();
 sg13g2_decap_8 FILLER_32_1151 ();
 sg13g2_decap_8 FILLER_32_1158 ();
 sg13g2_decap_8 FILLER_32_1165 ();
 sg13g2_decap_8 FILLER_32_1172 ();
 sg13g2_fill_2 FILLER_32_1179 ();
 sg13g2_decap_4 FILLER_32_1184 ();
 sg13g2_fill_2 FILLER_32_1188 ();
 sg13g2_fill_1 FILLER_32_1211 ();
 sg13g2_decap_4 FILLER_32_1220 ();
 sg13g2_fill_2 FILLER_32_1224 ();
 sg13g2_fill_2 FILLER_32_1248 ();
 sg13g2_fill_1 FILLER_32_1250 ();
 sg13g2_decap_4 FILLER_32_1260 ();
 sg13g2_decap_8 FILLER_32_1290 ();
 sg13g2_decap_8 FILLER_32_1297 ();
 sg13g2_decap_4 FILLER_32_1304 ();
 sg13g2_fill_2 FILLER_32_1308 ();
 sg13g2_decap_8 FILLER_32_1314 ();
 sg13g2_decap_4 FILLER_32_1321 ();
 sg13g2_fill_1 FILLER_32_1325 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_27 ();
 sg13g2_fill_1 FILLER_33_29 ();
 sg13g2_decap_4 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_decap_8 FILLER_33_73 ();
 sg13g2_decap_8 FILLER_33_80 ();
 sg13g2_fill_2 FILLER_33_87 ();
 sg13g2_decap_8 FILLER_33_117 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_4 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_162 ();
 sg13g2_decap_8 FILLER_33_167 ();
 sg13g2_decap_8 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_185 ();
 sg13g2_decap_8 FILLER_33_192 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_229 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_decap_8 FILLER_33_247 ();
 sg13g2_fill_2 FILLER_33_254 ();
 sg13g2_decap_4 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_263 ();
 sg13g2_decap_4 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_281 ();
 sg13g2_fill_2 FILLER_33_287 ();
 sg13g2_decap_4 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_296 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_2 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_316 ();
 sg13g2_decap_8 FILLER_33_327 ();
 sg13g2_fill_1 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_fill_2 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_33_389 ();
 sg13g2_fill_1 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_33_411 ();
 sg13g2_fill_2 FILLER_33_417 ();
 sg13g2_fill_1 FILLER_33_423 ();
 sg13g2_fill_2 FILLER_33_430 ();
 sg13g2_fill_1 FILLER_33_435 ();
 sg13g2_decap_8 FILLER_33_446 ();
 sg13g2_decap_8 FILLER_33_453 ();
 sg13g2_fill_2 FILLER_33_460 ();
 sg13g2_decap_8 FILLER_33_466 ();
 sg13g2_fill_2 FILLER_33_473 ();
 sg13g2_decap_4 FILLER_33_482 ();
 sg13g2_fill_2 FILLER_33_491 ();
 sg13g2_fill_1 FILLER_33_493 ();
 sg13g2_fill_1 FILLER_33_497 ();
 sg13g2_fill_2 FILLER_33_504 ();
 sg13g2_fill_1 FILLER_33_506 ();
 sg13g2_decap_8 FILLER_33_526 ();
 sg13g2_fill_1 FILLER_33_533 ();
 sg13g2_decap_4 FILLER_33_538 ();
 sg13g2_decap_8 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_decap_4 FILLER_33_567 ();
 sg13g2_fill_1 FILLER_33_594 ();
 sg13g2_fill_1 FILLER_33_606 ();
 sg13g2_fill_1 FILLER_33_611 ();
 sg13g2_fill_2 FILLER_33_621 ();
 sg13g2_fill_2 FILLER_33_626 ();
 sg13g2_fill_1 FILLER_33_638 ();
 sg13g2_fill_1 FILLER_33_678 ();
 sg13g2_fill_1 FILLER_33_683 ();
 sg13g2_decap_4 FILLER_33_710 ();
 sg13g2_fill_2 FILLER_33_714 ();
 sg13g2_decap_4 FILLER_33_720 ();
 sg13g2_decap_8 FILLER_33_747 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_fill_2 FILLER_33_770 ();
 sg13g2_fill_1 FILLER_33_776 ();
 sg13g2_fill_2 FILLER_33_789 ();
 sg13g2_fill_2 FILLER_33_801 ();
 sg13g2_fill_1 FILLER_33_803 ();
 sg13g2_decap_4 FILLER_33_815 ();
 sg13g2_fill_2 FILLER_33_819 ();
 sg13g2_fill_2 FILLER_33_831 ();
 sg13g2_fill_1 FILLER_33_833 ();
 sg13g2_fill_2 FILLER_33_837 ();
 sg13g2_decap_8 FILLER_33_859 ();
 sg13g2_decap_8 FILLER_33_870 ();
 sg13g2_decap_4 FILLER_33_877 ();
 sg13g2_fill_2 FILLER_33_881 ();
 sg13g2_decap_8 FILLER_33_892 ();
 sg13g2_decap_8 FILLER_33_899 ();
 sg13g2_fill_2 FILLER_33_906 ();
 sg13g2_fill_1 FILLER_33_913 ();
 sg13g2_decap_8 FILLER_33_927 ();
 sg13g2_fill_2 FILLER_33_939 ();
 sg13g2_fill_1 FILLER_33_941 ();
 sg13g2_fill_1 FILLER_33_958 ();
 sg13g2_fill_1 FILLER_33_964 ();
 sg13g2_fill_2 FILLER_33_974 ();
 sg13g2_fill_1 FILLER_33_976 ();
 sg13g2_decap_8 FILLER_33_983 ();
 sg13g2_fill_1 FILLER_33_990 ();
 sg13g2_decap_4 FILLER_33_1001 ();
 sg13g2_fill_2 FILLER_33_1014 ();
 sg13g2_fill_2 FILLER_33_1020 ();
 sg13g2_fill_1 FILLER_33_1022 ();
 sg13g2_fill_2 FILLER_33_1029 ();
 sg13g2_fill_1 FILLER_33_1031 ();
 sg13g2_fill_1 FILLER_33_1038 ();
 sg13g2_decap_4 FILLER_33_1044 ();
 sg13g2_fill_2 FILLER_33_1056 ();
 sg13g2_fill_1 FILLER_33_1058 ();
 sg13g2_fill_2 FILLER_33_1081 ();
 sg13g2_fill_2 FILLER_33_1091 ();
 sg13g2_decap_4 FILLER_33_1103 ();
 sg13g2_fill_2 FILLER_33_1111 ();
 sg13g2_fill_1 FILLER_33_1113 ();
 sg13g2_decap_4 FILLER_33_1123 ();
 sg13g2_fill_2 FILLER_33_1127 ();
 sg13g2_fill_1 FILLER_33_1134 ();
 sg13g2_decap_8 FILLER_33_1138 ();
 sg13g2_fill_1 FILLER_33_1182 ();
 sg13g2_fill_2 FILLER_33_1192 ();
 sg13g2_fill_1 FILLER_33_1208 ();
 sg13g2_decap_8 FILLER_33_1282 ();
 sg13g2_fill_2 FILLER_33_1298 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_11 ();
 sg13g2_fill_2 FILLER_34_17 ();
 sg13g2_decap_8 FILLER_34_23 ();
 sg13g2_fill_1 FILLER_34_30 ();
 sg13g2_decap_4 FILLER_34_39 ();
 sg13g2_fill_1 FILLER_34_43 ();
 sg13g2_decap_4 FILLER_34_48 ();
 sg13g2_decap_4 FILLER_34_61 ();
 sg13g2_fill_1 FILLER_34_65 ();
 sg13g2_fill_2 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_fill_2 FILLER_34_117 ();
 sg13g2_decap_8 FILLER_34_127 ();
 sg13g2_fill_2 FILLER_34_134 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_decap_8 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_167 ();
 sg13g2_fill_2 FILLER_34_171 ();
 sg13g2_decap_8 FILLER_34_180 ();
 sg13g2_fill_2 FILLER_34_187 ();
 sg13g2_decap_8 FILLER_34_194 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_fill_2 FILLER_34_208 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_290 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_fill_2 FILLER_34_304 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_fill_1 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_366 ();
 sg13g2_decap_8 FILLER_34_373 ();
 sg13g2_fill_2 FILLER_34_380 ();
 sg13g2_decap_4 FILLER_34_391 ();
 sg13g2_decap_4 FILLER_34_399 ();
 sg13g2_fill_1 FILLER_34_403 ();
 sg13g2_decap_4 FILLER_34_410 ();
 sg13g2_fill_1 FILLER_34_414 ();
 sg13g2_decap_8 FILLER_34_442 ();
 sg13g2_decap_8 FILLER_34_449 ();
 sg13g2_decap_4 FILLER_34_456 ();
 sg13g2_decap_4 FILLER_34_464 ();
 sg13g2_fill_1 FILLER_34_468 ();
 sg13g2_decap_8 FILLER_34_489 ();
 sg13g2_decap_8 FILLER_34_496 ();
 sg13g2_decap_4 FILLER_34_503 ();
 sg13g2_fill_2 FILLER_34_507 ();
 sg13g2_fill_1 FILLER_34_520 ();
 sg13g2_decap_4 FILLER_34_526 ();
 sg13g2_fill_1 FILLER_34_530 ();
 sg13g2_decap_8 FILLER_34_535 ();
 sg13g2_fill_2 FILLER_34_545 ();
 sg13g2_decap_8 FILLER_34_552 ();
 sg13g2_decap_4 FILLER_34_559 ();
 sg13g2_decap_8 FILLER_34_570 ();
 sg13g2_decap_8 FILLER_34_577 ();
 sg13g2_fill_1 FILLER_34_584 ();
 sg13g2_fill_2 FILLER_34_588 ();
 sg13g2_fill_2 FILLER_34_618 ();
 sg13g2_fill_1 FILLER_34_664 ();
 sg13g2_decap_8 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_691 ();
 sg13g2_fill_2 FILLER_34_698 ();
 sg13g2_fill_2 FILLER_34_731 ();
 sg13g2_fill_1 FILLER_34_733 ();
 sg13g2_decap_4 FILLER_34_738 ();
 sg13g2_fill_2 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_fill_1 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_779 ();
 sg13g2_decap_8 FILLER_34_786 ();
 sg13g2_fill_2 FILLER_34_793 ();
 sg13g2_decap_8 FILLER_34_799 ();
 sg13g2_fill_2 FILLER_34_806 ();
 sg13g2_decap_8 FILLER_34_811 ();
 sg13g2_fill_2 FILLER_34_818 ();
 sg13g2_decap_4 FILLER_34_829 ();
 sg13g2_decap_4 FILLER_34_845 ();
 sg13g2_fill_1 FILLER_34_849 ();
 sg13g2_fill_2 FILLER_34_853 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_fill_1 FILLER_34_867 ();
 sg13g2_fill_2 FILLER_34_873 ();
 sg13g2_fill_1 FILLER_34_875 ();
 sg13g2_fill_1 FILLER_34_881 ();
 sg13g2_decap_8 FILLER_34_904 ();
 sg13g2_fill_2 FILLER_34_931 ();
 sg13g2_decap_4 FILLER_34_938 ();
 sg13g2_fill_2 FILLER_34_957 ();
 sg13g2_fill_1 FILLER_34_959 ();
 sg13g2_fill_1 FILLER_34_990 ();
 sg13g2_decap_4 FILLER_34_1008 ();
 sg13g2_fill_2 FILLER_34_1023 ();
 sg13g2_fill_1 FILLER_34_1030 ();
 sg13g2_decap_4 FILLER_34_1044 ();
 sg13g2_fill_2 FILLER_34_1048 ();
 sg13g2_fill_1 FILLER_34_1083 ();
 sg13g2_fill_1 FILLER_34_1087 ();
 sg13g2_decap_8 FILLER_34_1101 ();
 sg13g2_fill_1 FILLER_34_1112 ();
 sg13g2_fill_1 FILLER_34_1117 ();
 sg13g2_fill_2 FILLER_34_1123 ();
 sg13g2_decap_4 FILLER_34_1129 ();
 sg13g2_fill_1 FILLER_34_1133 ();
 sg13g2_fill_1 FILLER_34_1160 ();
 sg13g2_decap_8 FILLER_34_1166 ();
 sg13g2_fill_2 FILLER_34_1173 ();
 sg13g2_fill_1 FILLER_34_1180 ();
 sg13g2_fill_2 FILLER_34_1202 ();
 sg13g2_fill_1 FILLER_34_1208 ();
 sg13g2_fill_1 FILLER_34_1213 ();
 sg13g2_decap_8 FILLER_34_1222 ();
 sg13g2_fill_2 FILLER_34_1229 ();
 sg13g2_decap_8 FILLER_34_1239 ();
 sg13g2_fill_1 FILLER_34_1246 ();
 sg13g2_fill_1 FILLER_34_1254 ();
 sg13g2_fill_1 FILLER_34_1269 ();
 sg13g2_fill_1 FILLER_34_1277 ();
 sg13g2_decap_8 FILLER_34_1317 ();
 sg13g2_fill_2 FILLER_34_1324 ();
 sg13g2_decap_8 FILLER_35_26 ();
 sg13g2_fill_1 FILLER_35_38 ();
 sg13g2_fill_2 FILLER_35_65 ();
 sg13g2_fill_1 FILLER_35_67 ();
 sg13g2_fill_2 FILLER_35_80 ();
 sg13g2_fill_1 FILLER_35_82 ();
 sg13g2_fill_2 FILLER_35_88 ();
 sg13g2_decap_8 FILLER_35_94 ();
 sg13g2_fill_2 FILLER_35_101 ();
 sg13g2_fill_1 FILLER_35_115 ();
 sg13g2_fill_2 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_130 ();
 sg13g2_decap_4 FILLER_35_145 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_181 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_fill_1 FILLER_35_204 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_fill_1 FILLER_35_215 ();
 sg13g2_fill_1 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_225 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_fill_1 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_1 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_decap_8 FILLER_35_260 ();
 sg13g2_fill_2 FILLER_35_267 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_fill_1 FILLER_35_312 ();
 sg13g2_decap_8 FILLER_35_321 ();
 sg13g2_fill_2 FILLER_35_328 ();
 sg13g2_decap_8 FILLER_35_356 ();
 sg13g2_decap_8 FILLER_35_363 ();
 sg13g2_decap_8 FILLER_35_370 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_393 ();
 sg13g2_decap_8 FILLER_35_403 ();
 sg13g2_decap_4 FILLER_35_410 ();
 sg13g2_fill_2 FILLER_35_414 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_decap_8 FILLER_35_426 ();
 sg13g2_fill_1 FILLER_35_433 ();
 sg13g2_decap_4 FILLER_35_470 ();
 sg13g2_fill_1 FILLER_35_474 ();
 sg13g2_decap_8 FILLER_35_488 ();
 sg13g2_fill_1 FILLER_35_495 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_decap_4 FILLER_35_511 ();
 sg13g2_decap_8 FILLER_35_555 ();
 sg13g2_decap_8 FILLER_35_562 ();
 sg13g2_fill_2 FILLER_35_569 ();
 sg13g2_decap_8 FILLER_35_579 ();
 sg13g2_decap_8 FILLER_35_586 ();
 sg13g2_decap_4 FILLER_35_593 ();
 sg13g2_fill_2 FILLER_35_610 ();
 sg13g2_fill_1 FILLER_35_612 ();
 sg13g2_fill_2 FILLER_35_638 ();
 sg13g2_fill_1 FILLER_35_652 ();
 sg13g2_fill_2 FILLER_35_669 ();
 sg13g2_decap_8 FILLER_35_685 ();
 sg13g2_decap_8 FILLER_35_692 ();
 sg13g2_decap_8 FILLER_35_699 ();
 sg13g2_fill_1 FILLER_35_706 ();
 sg13g2_fill_2 FILLER_35_716 ();
 sg13g2_decap_4 FILLER_35_722 ();
 sg13g2_decap_8 FILLER_35_730 ();
 sg13g2_decap_8 FILLER_35_741 ();
 sg13g2_decap_8 FILLER_35_748 ();
 sg13g2_fill_1 FILLER_35_755 ();
 sg13g2_decap_8 FILLER_35_761 ();
 sg13g2_decap_8 FILLER_35_768 ();
 sg13g2_decap_8 FILLER_35_775 ();
 sg13g2_decap_4 FILLER_35_782 ();
 sg13g2_decap_8 FILLER_35_790 ();
 sg13g2_fill_1 FILLER_35_797 ();
 sg13g2_decap_4 FILLER_35_810 ();
 sg13g2_decap_4 FILLER_35_830 ();
 sg13g2_fill_1 FILLER_35_839 ();
 sg13g2_fill_2 FILLER_35_844 ();
 sg13g2_fill_1 FILLER_35_846 ();
 sg13g2_fill_2 FILLER_35_852 ();
 sg13g2_fill_1 FILLER_35_854 ();
 sg13g2_decap_8 FILLER_35_860 ();
 sg13g2_decap_8 FILLER_35_867 ();
 sg13g2_decap_8 FILLER_35_874 ();
 sg13g2_fill_2 FILLER_35_881 ();
 sg13g2_fill_1 FILLER_35_883 ();
 sg13g2_fill_1 FILLER_35_887 ();
 sg13g2_decap_4 FILLER_35_891 ();
 sg13g2_fill_1 FILLER_35_895 ();
 sg13g2_decap_8 FILLER_35_905 ();
 sg13g2_decap_4 FILLER_35_912 ();
 sg13g2_fill_2 FILLER_35_916 ();
 sg13g2_decap_8 FILLER_35_930 ();
 sg13g2_decap_4 FILLER_35_945 ();
 sg13g2_fill_1 FILLER_35_949 ();
 sg13g2_fill_1 FILLER_35_965 ();
 sg13g2_fill_2 FILLER_35_971 ();
 sg13g2_decap_4 FILLER_35_976 ();
 sg13g2_fill_1 FILLER_35_980 ();
 sg13g2_fill_1 FILLER_35_986 ();
 sg13g2_fill_1 FILLER_35_992 ();
 sg13g2_decap_8 FILLER_35_996 ();
 sg13g2_decap_8 FILLER_35_1029 ();
 sg13g2_decap_8 FILLER_35_1036 ();
 sg13g2_decap_8 FILLER_35_1043 ();
 sg13g2_fill_2 FILLER_35_1050 ();
 sg13g2_fill_2 FILLER_35_1056 ();
 sg13g2_fill_1 FILLER_35_1058 ();
 sg13g2_fill_1 FILLER_35_1062 ();
 sg13g2_decap_8 FILLER_35_1067 ();
 sg13g2_decap_4 FILLER_35_1074 ();
 sg13g2_fill_2 FILLER_35_1087 ();
 sg13g2_fill_1 FILLER_35_1098 ();
 sg13g2_decap_4 FILLER_35_1104 ();
 sg13g2_fill_1 FILLER_35_1108 ();
 sg13g2_decap_8 FILLER_35_1121 ();
 sg13g2_decap_8 FILLER_35_1128 ();
 sg13g2_decap_8 FILLER_35_1135 ();
 sg13g2_decap_8 FILLER_35_1142 ();
 sg13g2_decap_4 FILLER_35_1149 ();
 sg13g2_fill_2 FILLER_35_1179 ();
 sg13g2_fill_1 FILLER_35_1228 ();
 sg13g2_fill_2 FILLER_35_1240 ();
 sg13g2_fill_1 FILLER_35_1248 ();
 sg13g2_fill_2 FILLER_35_1254 ();
 sg13g2_fill_1 FILLER_35_1259 ();
 sg13g2_decap_8 FILLER_35_1286 ();
 sg13g2_fill_2 FILLER_35_1293 ();
 sg13g2_decap_8 FILLER_35_1300 ();
 sg13g2_decap_8 FILLER_35_1307 ();
 sg13g2_decap_8 FILLER_35_1314 ();
 sg13g2_decap_4 FILLER_35_1321 ();
 sg13g2_fill_1 FILLER_35_1325 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_31 ();
 sg13g2_fill_1 FILLER_36_33 ();
 sg13g2_decap_4 FILLER_36_48 ();
 sg13g2_decap_4 FILLER_36_56 ();
 sg13g2_fill_1 FILLER_36_60 ();
 sg13g2_fill_2 FILLER_36_77 ();
 sg13g2_fill_1 FILLER_36_79 ();
 sg13g2_fill_1 FILLER_36_90 ();
 sg13g2_fill_1 FILLER_36_94 ();
 sg13g2_fill_1 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_111 ();
 sg13g2_fill_1 FILLER_36_117 ();
 sg13g2_fill_1 FILLER_36_123 ();
 sg13g2_fill_1 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_150 ();
 sg13g2_fill_1 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_183 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_4 FILLER_36_238 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_decap_8 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_fill_2 FILLER_36_316 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_331 ();
 sg13g2_decap_4 FILLER_36_338 ();
 sg13g2_fill_1 FILLER_36_351 ();
 sg13g2_fill_1 FILLER_36_357 ();
 sg13g2_decap_4 FILLER_36_368 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_2 FILLER_36_417 ();
 sg13g2_decap_8 FILLER_36_431 ();
 sg13g2_decap_8 FILLER_36_438 ();
 sg13g2_decap_8 FILLER_36_445 ();
 sg13g2_decap_8 FILLER_36_452 ();
 sg13g2_decap_8 FILLER_36_459 ();
 sg13g2_decap_4 FILLER_36_466 ();
 sg13g2_fill_1 FILLER_36_470 ();
 sg13g2_decap_4 FILLER_36_485 ();
 sg13g2_fill_2 FILLER_36_530 ();
 sg13g2_fill_1 FILLER_36_544 ();
 sg13g2_fill_1 FILLER_36_554 ();
 sg13g2_fill_2 FILLER_36_564 ();
 sg13g2_fill_1 FILLER_36_569 ();
 sg13g2_fill_1 FILLER_36_575 ();
 sg13g2_fill_2 FILLER_36_580 ();
 sg13g2_fill_2 FILLER_36_586 ();
 sg13g2_fill_1 FILLER_36_588 ();
 sg13g2_decap_8 FILLER_36_593 ();
 sg13g2_fill_1 FILLER_36_600 ();
 sg13g2_fill_2 FILLER_36_615 ();
 sg13g2_fill_2 FILLER_36_633 ();
 sg13g2_fill_1 FILLER_36_641 ();
 sg13g2_fill_2 FILLER_36_650 ();
 sg13g2_fill_2 FILLER_36_661 ();
 sg13g2_fill_2 FILLER_36_675 ();
 sg13g2_fill_2 FILLER_36_687 ();
 sg13g2_fill_1 FILLER_36_689 ();
 sg13g2_fill_1 FILLER_36_716 ();
 sg13g2_fill_2 FILLER_36_752 ();
 sg13g2_fill_1 FILLER_36_754 ();
 sg13g2_fill_2 FILLER_36_758 ();
 sg13g2_fill_1 FILLER_36_760 ();
 sg13g2_decap_4 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_788 ();
 sg13g2_decap_4 FILLER_36_795 ();
 sg13g2_fill_1 FILLER_36_799 ();
 sg13g2_decap_8 FILLER_36_836 ();
 sg13g2_decap_8 FILLER_36_843 ();
 sg13g2_decap_8 FILLER_36_850 ();
 sg13g2_decap_4 FILLER_36_857 ();
 sg13g2_fill_2 FILLER_36_865 ();
 sg13g2_fill_2 FILLER_36_872 ();
 sg13g2_fill_1 FILLER_36_883 ();
 sg13g2_decap_4 FILLER_36_887 ();
 sg13g2_fill_1 FILLER_36_891 ();
 sg13g2_fill_2 FILLER_36_921 ();
 sg13g2_decap_4 FILLER_36_931 ();
 sg13g2_fill_2 FILLER_36_935 ();
 sg13g2_fill_1 FILLER_36_946 ();
 sg13g2_decap_8 FILLER_36_965 ();
 sg13g2_decap_4 FILLER_36_972 ();
 sg13g2_fill_2 FILLER_36_986 ();
 sg13g2_decap_4 FILLER_36_1002 ();
 sg13g2_fill_1 FILLER_36_1006 ();
 sg13g2_fill_1 FILLER_36_1011 ();
 sg13g2_fill_2 FILLER_36_1020 ();
 sg13g2_fill_1 FILLER_36_1022 ();
 sg13g2_fill_2 FILLER_36_1030 ();
 sg13g2_fill_2 FILLER_36_1037 ();
 sg13g2_fill_1 FILLER_36_1039 ();
 sg13g2_fill_1 FILLER_36_1045 ();
 sg13g2_fill_2 FILLER_36_1062 ();
 sg13g2_fill_1 FILLER_36_1064 ();
 sg13g2_fill_2 FILLER_36_1070 ();
 sg13g2_fill_1 FILLER_36_1113 ();
 sg13g2_decap_8 FILLER_36_1118 ();
 sg13g2_fill_2 FILLER_36_1134 ();
 sg13g2_fill_1 FILLER_36_1136 ();
 sg13g2_fill_2 FILLER_36_1142 ();
 sg13g2_fill_1 FILLER_36_1148 ();
 sg13g2_fill_2 FILLER_36_1158 ();
 sg13g2_fill_1 FILLER_36_1179 ();
 sg13g2_fill_1 FILLER_36_1221 ();
 sg13g2_fill_2 FILLER_36_1246 ();
 sg13g2_decap_8 FILLER_36_1257 ();
 sg13g2_decap_4 FILLER_36_1264 ();
 sg13g2_decap_4 FILLER_36_1276 ();
 sg13g2_fill_2 FILLER_36_1280 ();
 sg13g2_fill_2 FILLER_36_1286 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_37 ();
 sg13g2_fill_2 FILLER_37_44 ();
 sg13g2_decap_8 FILLER_37_60 ();
 sg13g2_decap_8 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_74 ();
 sg13g2_fill_1 FILLER_37_81 ();
 sg13g2_fill_1 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_138 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_fill_2 FILLER_37_154 ();
 sg13g2_fill_1 FILLER_37_156 ();
 sg13g2_fill_2 FILLER_37_162 ();
 sg13g2_fill_2 FILLER_37_168 ();
 sg13g2_fill_1 FILLER_37_170 ();
 sg13g2_fill_2 FILLER_37_176 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_decap_4 FILLER_37_240 ();
 sg13g2_fill_2 FILLER_37_244 ();
 sg13g2_decap_8 FILLER_37_251 ();
 sg13g2_decap_4 FILLER_37_258 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_268 ();
 sg13g2_fill_1 FILLER_37_278 ();
 sg13g2_fill_2 FILLER_37_296 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_350 ();
 sg13g2_fill_1 FILLER_37_352 ();
 sg13g2_decap_4 FILLER_37_379 ();
 sg13g2_fill_1 FILLER_37_383 ();
 sg13g2_fill_1 FILLER_37_392 ();
 sg13g2_fill_2 FILLER_37_402 ();
 sg13g2_fill_1 FILLER_37_415 ();
 sg13g2_fill_1 FILLER_37_439 ();
 sg13g2_fill_1 FILLER_37_444 ();
 sg13g2_fill_1 FILLER_37_450 ();
 sg13g2_decap_8 FILLER_37_459 ();
 sg13g2_decap_8 FILLER_37_466 ();
 sg13g2_decap_4 FILLER_37_473 ();
 sg13g2_fill_2 FILLER_37_481 ();
 sg13g2_decap_4 FILLER_37_487 ();
 sg13g2_fill_2 FILLER_37_491 ();
 sg13g2_decap_4 FILLER_37_499 ();
 sg13g2_fill_2 FILLER_37_503 ();
 sg13g2_fill_2 FILLER_37_513 ();
 sg13g2_fill_2 FILLER_37_524 ();
 sg13g2_decap_4 FILLER_37_537 ();
 sg13g2_fill_1 FILLER_37_541 ();
 sg13g2_fill_2 FILLER_37_549 ();
 sg13g2_fill_1 FILLER_37_551 ();
 sg13g2_fill_1 FILLER_37_560 ();
 sg13g2_fill_2 FILLER_37_565 ();
 sg13g2_fill_1 FILLER_37_567 ();
 sg13g2_fill_2 FILLER_37_577 ();
 sg13g2_decap_8 FILLER_37_583 ();
 sg13g2_decap_4 FILLER_37_590 ();
 sg13g2_fill_2 FILLER_37_594 ();
 sg13g2_decap_8 FILLER_37_611 ();
 sg13g2_decap_8 FILLER_37_618 ();
 sg13g2_fill_2 FILLER_37_625 ();
 sg13g2_fill_1 FILLER_37_627 ();
 sg13g2_decap_8 FILLER_37_682 ();
 sg13g2_decap_8 FILLER_37_695 ();
 sg13g2_decap_4 FILLER_37_702 ();
 sg13g2_fill_2 FILLER_37_706 ();
 sg13g2_fill_1 FILLER_37_745 ();
 sg13g2_fill_1 FILLER_37_754 ();
 sg13g2_fill_2 FILLER_37_779 ();
 sg13g2_fill_1 FILLER_37_781 ();
 sg13g2_fill_2 FILLER_37_794 ();
 sg13g2_fill_1 FILLER_37_796 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_4 FILLER_37_819 ();
 sg13g2_fill_1 FILLER_37_823 ();
 sg13g2_fill_1 FILLER_37_845 ();
 sg13g2_fill_2 FILLER_37_863 ();
 sg13g2_decap_8 FILLER_37_899 ();
 sg13g2_decap_8 FILLER_37_906 ();
 sg13g2_fill_2 FILLER_37_913 ();
 sg13g2_fill_1 FILLER_37_915 ();
 sg13g2_fill_2 FILLER_37_936 ();
 sg13g2_decap_8 FILLER_37_947 ();
 sg13g2_fill_2 FILLER_37_954 ();
 sg13g2_fill_1 FILLER_37_956 ();
 sg13g2_fill_2 FILLER_37_963 ();
 sg13g2_decap_4 FILLER_37_969 ();
 sg13g2_decap_4 FILLER_37_984 ();
 sg13g2_decap_4 FILLER_37_993 ();
 sg13g2_fill_1 FILLER_37_997 ();
 sg13g2_fill_2 FILLER_37_1028 ();
 sg13g2_fill_1 FILLER_37_1030 ();
 sg13g2_fill_2 FILLER_37_1036 ();
 sg13g2_decap_8 FILLER_37_1042 ();
 sg13g2_fill_2 FILLER_37_1049 ();
 sg13g2_fill_1 FILLER_37_1051 ();
 sg13g2_decap_8 FILLER_37_1055 ();
 sg13g2_decap_8 FILLER_37_1062 ();
 sg13g2_decap_4 FILLER_37_1074 ();
 sg13g2_fill_1 FILLER_37_1078 ();
 sg13g2_decap_4 FILLER_37_1085 ();
 sg13g2_fill_1 FILLER_37_1089 ();
 sg13g2_fill_1 FILLER_37_1100 ();
 sg13g2_fill_1 FILLER_37_1106 ();
 sg13g2_decap_8 FILLER_37_1110 ();
 sg13g2_decap_8 FILLER_37_1120 ();
 sg13g2_decap_8 FILLER_37_1127 ();
 sg13g2_decap_8 FILLER_37_1134 ();
 sg13g2_decap_8 FILLER_37_1141 ();
 sg13g2_fill_1 FILLER_37_1148 ();
 sg13g2_decap_8 FILLER_37_1159 ();
 sg13g2_decap_4 FILLER_37_1166 ();
 sg13g2_fill_2 FILLER_37_1170 ();
 sg13g2_decap_4 FILLER_37_1180 ();
 sg13g2_fill_1 FILLER_37_1184 ();
 sg13g2_fill_1 FILLER_37_1197 ();
 sg13g2_decap_8 FILLER_37_1209 ();
 sg13g2_decap_4 FILLER_37_1216 ();
 sg13g2_fill_1 FILLER_37_1220 ();
 sg13g2_decap_8 FILLER_37_1225 ();
 sg13g2_fill_2 FILLER_37_1232 ();
 sg13g2_decap_8 FILLER_37_1245 ();
 sg13g2_decap_8 FILLER_37_1252 ();
 sg13g2_decap_8 FILLER_37_1299 ();
 sg13g2_decap_8 FILLER_37_1306 ();
 sg13g2_decap_8 FILLER_37_1313 ();
 sg13g2_decap_4 FILLER_37_1320 ();
 sg13g2_fill_2 FILLER_37_1324 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_4 ();
 sg13g2_fill_1 FILLER_38_41 ();
 sg13g2_fill_1 FILLER_38_46 ();
 sg13g2_fill_1 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_69 ();
 sg13g2_decap_4 FILLER_38_77 ();
 sg13g2_fill_1 FILLER_38_89 ();
 sg13g2_fill_1 FILLER_38_98 ();
 sg13g2_fill_2 FILLER_38_106 ();
 sg13g2_decap_4 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_146 ();
 sg13g2_fill_2 FILLER_38_153 ();
 sg13g2_fill_1 FILLER_38_155 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_fill_1 FILLER_38_200 ();
 sg13g2_fill_2 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_fill_1 FILLER_38_225 ();
 sg13g2_decap_4 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_251 ();
 sg13g2_decap_4 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_4 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_decap_8 FILLER_38_323 ();
 sg13g2_decap_8 FILLER_38_330 ();
 sg13g2_decap_4 FILLER_38_337 ();
 sg13g2_decap_8 FILLER_38_346 ();
 sg13g2_decap_4 FILLER_38_353 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_fill_1 FILLER_38_363 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_fill_1 FILLER_38_405 ();
 sg13g2_fill_1 FILLER_38_411 ();
 sg13g2_fill_1 FILLER_38_419 ();
 sg13g2_fill_2 FILLER_38_437 ();
 sg13g2_fill_1 FILLER_38_443 ();
 sg13g2_decap_8 FILLER_38_454 ();
 sg13g2_fill_1 FILLER_38_461 ();
 sg13g2_fill_2 FILLER_38_466 ();
 sg13g2_fill_1 FILLER_38_468 ();
 sg13g2_fill_1 FILLER_38_472 ();
 sg13g2_decap_8 FILLER_38_478 ();
 sg13g2_fill_2 FILLER_38_485 ();
 sg13g2_fill_1 FILLER_38_492 ();
 sg13g2_fill_2 FILLER_38_505 ();
 sg13g2_fill_1 FILLER_38_519 ();
 sg13g2_decap_4 FILLER_38_529 ();
 sg13g2_fill_1 FILLER_38_533 ();
 sg13g2_fill_1 FILLER_38_538 ();
 sg13g2_fill_2 FILLER_38_544 ();
 sg13g2_fill_1 FILLER_38_546 ();
 sg13g2_decap_4 FILLER_38_550 ();
 sg13g2_fill_1 FILLER_38_554 ();
 sg13g2_decap_4 FILLER_38_597 ();
 sg13g2_fill_2 FILLER_38_601 ();
 sg13g2_fill_2 FILLER_38_648 ();
 sg13g2_fill_2 FILLER_38_656 ();
 sg13g2_fill_2 FILLER_38_695 ();
 sg13g2_decap_4 FILLER_38_712 ();
 sg13g2_fill_2 FILLER_38_722 ();
 sg13g2_fill_2 FILLER_38_732 ();
 sg13g2_decap_4 FILLER_38_742 ();
 sg13g2_fill_2 FILLER_38_746 ();
 sg13g2_fill_2 FILLER_38_757 ();
 sg13g2_fill_1 FILLER_38_776 ();
 sg13g2_fill_1 FILLER_38_788 ();
 sg13g2_fill_2 FILLER_38_800 ();
 sg13g2_fill_2 FILLER_38_818 ();
 sg13g2_fill_1 FILLER_38_820 ();
 sg13g2_fill_2 FILLER_38_825 ();
 sg13g2_fill_1 FILLER_38_827 ();
 sg13g2_decap_8 FILLER_38_839 ();
 sg13g2_decap_8 FILLER_38_846 ();
 sg13g2_fill_1 FILLER_38_853 ();
 sg13g2_decap_8 FILLER_38_862 ();
 sg13g2_decap_4 FILLER_38_869 ();
 sg13g2_fill_2 FILLER_38_873 ();
 sg13g2_decap_8 FILLER_38_879 ();
 sg13g2_decap_8 FILLER_38_892 ();
 sg13g2_decap_8 FILLER_38_899 ();
 sg13g2_decap_8 FILLER_38_906 ();
 sg13g2_decap_8 FILLER_38_913 ();
 sg13g2_fill_2 FILLER_38_920 ();
 sg13g2_fill_1 FILLER_38_922 ();
 sg13g2_fill_1 FILLER_38_926 ();
 sg13g2_fill_1 FILLER_38_935 ();
 sg13g2_decap_4 FILLER_38_962 ();
 sg13g2_decap_4 FILLER_38_970 ();
 sg13g2_decap_8 FILLER_38_978 ();
 sg13g2_decap_8 FILLER_38_985 ();
 sg13g2_fill_2 FILLER_38_992 ();
 sg13g2_decap_4 FILLER_38_1003 ();
 sg13g2_fill_2 FILLER_38_1033 ();
 sg13g2_decap_4 FILLER_38_1048 ();
 sg13g2_decap_8 FILLER_38_1056 ();
 sg13g2_decap_4 FILLER_38_1063 ();
 sg13g2_fill_1 FILLER_38_1067 ();
 sg13g2_decap_4 FILLER_38_1073 ();
 sg13g2_decap_8 FILLER_38_1082 ();
 sg13g2_fill_2 FILLER_38_1089 ();
 sg13g2_fill_1 FILLER_38_1091 ();
 sg13g2_fill_1 FILLER_38_1104 ();
 sg13g2_fill_1 FILLER_38_1109 ();
 sg13g2_fill_1 FILLER_38_1113 ();
 sg13g2_fill_1 FILLER_38_1124 ();
 sg13g2_fill_1 FILLER_38_1135 ();
 sg13g2_decap_8 FILLER_38_1146 ();
 sg13g2_fill_2 FILLER_38_1153 ();
 sg13g2_decap_8 FILLER_38_1160 ();
 sg13g2_decap_4 FILLER_38_1167 ();
 sg13g2_fill_1 FILLER_38_1171 ();
 sg13g2_decap_8 FILLER_38_1176 ();
 sg13g2_fill_2 FILLER_38_1183 ();
 sg13g2_fill_1 FILLER_38_1185 ();
 sg13g2_fill_1 FILLER_38_1191 ();
 sg13g2_fill_1 FILLER_38_1197 ();
 sg13g2_decap_8 FILLER_38_1208 ();
 sg13g2_decap_4 FILLER_38_1215 ();
 sg13g2_fill_2 FILLER_38_1219 ();
 sg13g2_decap_8 FILLER_38_1229 ();
 sg13g2_decap_4 FILLER_38_1236 ();
 sg13g2_decap_8 FILLER_38_1266 ();
 sg13g2_decap_8 FILLER_38_1273 ();
 sg13g2_fill_2 FILLER_38_1280 ();
 sg13g2_fill_1 FILLER_38_1282 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_37 ();
 sg13g2_decap_4 FILLER_39_44 ();
 sg13g2_fill_2 FILLER_39_54 ();
 sg13g2_fill_1 FILLER_39_56 ();
 sg13g2_decap_4 FILLER_39_60 ();
 sg13g2_fill_1 FILLER_39_64 ();
 sg13g2_fill_1 FILLER_39_74 ();
 sg13g2_fill_2 FILLER_39_114 ();
 sg13g2_fill_1 FILLER_39_137 ();
 sg13g2_fill_1 FILLER_39_143 ();
 sg13g2_fill_2 FILLER_39_148 ();
 sg13g2_fill_2 FILLER_39_154 ();
 sg13g2_fill_2 FILLER_39_171 ();
 sg13g2_fill_2 FILLER_39_176 ();
 sg13g2_fill_1 FILLER_39_178 ();
 sg13g2_fill_2 FILLER_39_183 ();
 sg13g2_decap_4 FILLER_39_214 ();
 sg13g2_fill_1 FILLER_39_218 ();
 sg13g2_fill_1 FILLER_39_256 ();
 sg13g2_fill_1 FILLER_39_270 ();
 sg13g2_decap_4 FILLER_39_274 ();
 sg13g2_fill_2 FILLER_39_278 ();
 sg13g2_decap_8 FILLER_39_317 ();
 sg13g2_decap_8 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_347 ();
 sg13g2_fill_2 FILLER_39_354 ();
 sg13g2_fill_1 FILLER_39_367 ();
 sg13g2_fill_2 FILLER_39_390 ();
 sg13g2_fill_1 FILLER_39_392 ();
 sg13g2_fill_1 FILLER_39_407 ();
 sg13g2_fill_1 FILLER_39_413 ();
 sg13g2_fill_1 FILLER_39_424 ();
 sg13g2_decap_8 FILLER_39_437 ();
 sg13g2_fill_1 FILLER_39_444 ();
 sg13g2_decap_4 FILLER_39_459 ();
 sg13g2_fill_2 FILLER_39_471 ();
 sg13g2_fill_2 FILLER_39_483 ();
 sg13g2_fill_2 FILLER_39_490 ();
 sg13g2_fill_1 FILLER_39_492 ();
 sg13g2_decap_4 FILLER_39_503 ();
 sg13g2_fill_1 FILLER_39_511 ();
 sg13g2_decap_4 FILLER_39_530 ();
 sg13g2_fill_2 FILLER_39_549 ();
 sg13g2_fill_1 FILLER_39_551 ();
 sg13g2_decap_4 FILLER_39_557 ();
 sg13g2_fill_2 FILLER_39_570 ();
 sg13g2_fill_1 FILLER_39_572 ();
 sg13g2_decap_8 FILLER_39_581 ();
 sg13g2_fill_1 FILLER_39_588 ();
 sg13g2_fill_2 FILLER_39_592 ();
 sg13g2_fill_2 FILLER_39_598 ();
 sg13g2_decap_8 FILLER_39_620 ();
 sg13g2_fill_1 FILLER_39_644 ();
 sg13g2_fill_2 FILLER_39_656 ();
 sg13g2_decap_8 FILLER_39_674 ();
 sg13g2_fill_2 FILLER_39_681 ();
 sg13g2_fill_1 FILLER_39_683 ();
 sg13g2_decap_4 FILLER_39_688 ();
 sg13g2_fill_2 FILLER_39_692 ();
 sg13g2_decap_8 FILLER_39_736 ();
 sg13g2_fill_2 FILLER_39_759 ();
 sg13g2_fill_1 FILLER_39_780 ();
 sg13g2_fill_1 FILLER_39_791 ();
 sg13g2_decap_4 FILLER_39_796 ();
 sg13g2_fill_1 FILLER_39_805 ();
 sg13g2_decap_8 FILLER_39_810 ();
 sg13g2_fill_2 FILLER_39_817 ();
 sg13g2_fill_2 FILLER_39_824 ();
 sg13g2_fill_1 FILLER_39_826 ();
 sg13g2_decap_8 FILLER_39_834 ();
 sg13g2_decap_4 FILLER_39_841 ();
 sg13g2_fill_2 FILLER_39_881 ();
 sg13g2_fill_2 FILLER_39_889 ();
 sg13g2_fill_2 FILLER_39_901 ();
 sg13g2_fill_1 FILLER_39_922 ();
 sg13g2_fill_2 FILLER_39_927 ();
 sg13g2_decap_8 FILLER_39_950 ();
 sg13g2_decap_8 FILLER_39_957 ();
 sg13g2_decap_8 FILLER_39_964 ();
 sg13g2_decap_4 FILLER_39_980 ();
 sg13g2_fill_2 FILLER_39_984 ();
 sg13g2_fill_2 FILLER_39_995 ();
 sg13g2_fill_2 FILLER_39_1002 ();
 sg13g2_fill_1 FILLER_39_1017 ();
 sg13g2_fill_2 FILLER_39_1030 ();
 sg13g2_fill_1 FILLER_39_1032 ();
 sg13g2_decap_8 FILLER_39_1037 ();
 sg13g2_decap_8 FILLER_39_1048 ();
 sg13g2_decap_8 FILLER_39_1069 ();
 sg13g2_fill_2 FILLER_39_1076 ();
 sg13g2_decap_8 FILLER_39_1090 ();
 sg13g2_decap_8 FILLER_39_1097 ();
 sg13g2_fill_1 FILLER_39_1104 ();
 sg13g2_fill_1 FILLER_39_1108 ();
 sg13g2_fill_2 FILLER_39_1113 ();
 sg13g2_fill_1 FILLER_39_1120 ();
 sg13g2_fill_1 FILLER_39_1126 ();
 sg13g2_fill_2 FILLER_39_1151 ();
 sg13g2_fill_1 FILLER_39_1163 ();
 sg13g2_fill_1 FILLER_39_1190 ();
 sg13g2_fill_1 FILLER_39_1200 ();
 sg13g2_decap_4 FILLER_39_1222 ();
 sg13g2_decap_8 FILLER_39_1249 ();
 sg13g2_decap_4 FILLER_39_1264 ();
 sg13g2_fill_2 FILLER_39_1272 ();
 sg13g2_fill_1 FILLER_39_1274 ();
 sg13g2_decap_8 FILLER_39_1288 ();
 sg13g2_decap_8 FILLER_39_1295 ();
 sg13g2_decap_8 FILLER_39_1302 ();
 sg13g2_decap_8 FILLER_39_1309 ();
 sg13g2_decap_8 FILLER_39_1316 ();
 sg13g2_fill_2 FILLER_39_1323 ();
 sg13g2_fill_1 FILLER_39_1325 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_59 ();
 sg13g2_fill_2 FILLER_40_63 ();
 sg13g2_fill_1 FILLER_40_80 ();
 sg13g2_fill_2 FILLER_40_110 ();
 sg13g2_fill_1 FILLER_40_130 ();
 sg13g2_fill_1 FILLER_40_143 ();
 sg13g2_fill_1 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_186 ();
 sg13g2_decap_8 FILLER_40_191 ();
 sg13g2_decap_8 FILLER_40_198 ();
 sg13g2_fill_2 FILLER_40_214 ();
 sg13g2_fill_1 FILLER_40_216 ();
 sg13g2_decap_4 FILLER_40_230 ();
 sg13g2_fill_2 FILLER_40_253 ();
 sg13g2_decap_4 FILLER_40_258 ();
 sg13g2_decap_4 FILLER_40_267 ();
 sg13g2_decap_8 FILLER_40_275 ();
 sg13g2_fill_2 FILLER_40_282 ();
 sg13g2_fill_1 FILLER_40_284 ();
 sg13g2_fill_2 FILLER_40_294 ();
 sg13g2_fill_1 FILLER_40_296 ();
 sg13g2_decap_8 FILLER_40_316 ();
 sg13g2_decap_8 FILLER_40_323 ();
 sg13g2_decap_4 FILLER_40_337 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_fill_1 FILLER_40_405 ();
 sg13g2_decap_8 FILLER_40_418 ();
 sg13g2_fill_2 FILLER_40_459 ();
 sg13g2_fill_1 FILLER_40_465 ();
 sg13g2_fill_1 FILLER_40_474 ();
 sg13g2_fill_1 FILLER_40_479 ();
 sg13g2_fill_1 FILLER_40_484 ();
 sg13g2_fill_1 FILLER_40_490 ();
 sg13g2_fill_1 FILLER_40_495 ();
 sg13g2_fill_2 FILLER_40_514 ();
 sg13g2_fill_1 FILLER_40_516 ();
 sg13g2_decap_4 FILLER_40_525 ();
 sg13g2_fill_2 FILLER_40_542 ();
 sg13g2_fill_1 FILLER_40_552 ();
 sg13g2_fill_1 FILLER_40_557 ();
 sg13g2_fill_2 FILLER_40_579 ();
 sg13g2_fill_2 FILLER_40_589 ();
 sg13g2_fill_1 FILLER_40_591 ();
 sg13g2_fill_1 FILLER_40_597 ();
 sg13g2_fill_2 FILLER_40_603 ();
 sg13g2_decap_8 FILLER_40_611 ();
 sg13g2_decap_4 FILLER_40_618 ();
 sg13g2_fill_2 FILLER_40_622 ();
 sg13g2_decap_4 FILLER_40_629 ();
 sg13g2_decap_8 FILLER_40_670 ();
 sg13g2_fill_1 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_696 ();
 sg13g2_fill_2 FILLER_40_721 ();
 sg13g2_fill_1 FILLER_40_729 ();
 sg13g2_fill_2 FILLER_40_734 ();
 sg13g2_decap_4 FILLER_40_740 ();
 sg13g2_fill_1 FILLER_40_744 ();
 sg13g2_fill_2 FILLER_40_749 ();
 sg13g2_fill_2 FILLER_40_773 ();
 sg13g2_decap_8 FILLER_40_792 ();
 sg13g2_decap_8 FILLER_40_799 ();
 sg13g2_fill_2 FILLER_40_806 ();
 sg13g2_fill_2 FILLER_40_836 ();
 sg13g2_fill_1 FILLER_40_838 ();
 sg13g2_fill_1 FILLER_40_848 ();
 sg13g2_fill_1 FILLER_40_854 ();
 sg13g2_fill_2 FILLER_40_861 ();
 sg13g2_fill_2 FILLER_40_893 ();
 sg13g2_fill_2 FILLER_40_959 ();
 sg13g2_fill_2 FILLER_40_966 ();
 sg13g2_fill_1 FILLER_40_968 ();
 sg13g2_decap_4 FILLER_40_973 ();
 sg13g2_fill_1 FILLER_40_980 ();
 sg13g2_decap_8 FILLER_40_989 ();
 sg13g2_decap_4 FILLER_40_1004 ();
 sg13g2_fill_1 FILLER_40_1008 ();
 sg13g2_decap_8 FILLER_40_1018 ();
 sg13g2_fill_1 FILLER_40_1042 ();
 sg13g2_decap_8 FILLER_40_1047 ();
 sg13g2_decap_4 FILLER_40_1057 ();
 sg13g2_decap_8 FILLER_40_1064 ();
 sg13g2_decap_8 FILLER_40_1071 ();
 sg13g2_decap_4 FILLER_40_1078 ();
 sg13g2_fill_1 FILLER_40_1082 ();
 sg13g2_fill_2 FILLER_40_1087 ();
 sg13g2_fill_2 FILLER_40_1126 ();
 sg13g2_decap_8 FILLER_40_1131 ();
 sg13g2_decap_4 FILLER_40_1138 ();
 sg13g2_fill_1 FILLER_40_1142 ();
 sg13g2_decap_8 FILLER_40_1147 ();
 sg13g2_decap_4 FILLER_40_1154 ();
 sg13g2_fill_1 FILLER_40_1158 ();
 sg13g2_fill_1 FILLER_40_1164 ();
 sg13g2_fill_2 FILLER_40_1178 ();
 sg13g2_fill_1 FILLER_40_1185 ();
 sg13g2_fill_1 FILLER_40_1190 ();
 sg13g2_fill_1 FILLER_40_1199 ();
 sg13g2_fill_1 FILLER_40_1224 ();
 sg13g2_fill_2 FILLER_40_1232 ();
 sg13g2_fill_1 FILLER_40_1234 ();
 sg13g2_decap_4 FILLER_40_1239 ();
 sg13g2_fill_2 FILLER_40_1251 ();
 sg13g2_decap_4 FILLER_40_1258 ();
 sg13g2_fill_2 FILLER_40_1262 ();
 sg13g2_fill_1 FILLER_40_1272 ();
 sg13g2_fill_2 FILLER_40_1303 ();
 sg13g2_fill_1 FILLER_40_1305 ();
 sg13g2_decap_8 FILLER_40_1310 ();
 sg13g2_decap_8 FILLER_40_1317 ();
 sg13g2_fill_2 FILLER_40_1324 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_55 ();
 sg13g2_fill_2 FILLER_41_62 ();
 sg13g2_fill_1 FILLER_41_64 ();
 sg13g2_fill_1 FILLER_41_68 ();
 sg13g2_fill_2 FILLER_41_78 ();
 sg13g2_fill_1 FILLER_41_94 ();
 sg13g2_fill_1 FILLER_41_157 ();
 sg13g2_fill_2 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_fill_1 FILLER_41_228 ();
 sg13g2_decap_4 FILLER_41_234 ();
 sg13g2_fill_2 FILLER_41_251 ();
 sg13g2_fill_1 FILLER_41_253 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_fill_2 FILLER_41_280 ();
 sg13g2_decap_4 FILLER_41_296 ();
 sg13g2_fill_2 FILLER_41_300 ();
 sg13g2_decap_8 FILLER_41_305 ();
 sg13g2_decap_4 FILLER_41_312 ();
 sg13g2_fill_1 FILLER_41_319 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_4 FILLER_41_339 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_fill_2 FILLER_41_375 ();
 sg13g2_fill_1 FILLER_41_377 ();
 sg13g2_fill_2 FILLER_41_382 ();
 sg13g2_fill_1 FILLER_41_384 ();
 sg13g2_decap_4 FILLER_41_388 ();
 sg13g2_fill_2 FILLER_41_392 ();
 sg13g2_fill_2 FILLER_41_401 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_fill_2 FILLER_41_421 ();
 sg13g2_decap_4 FILLER_41_438 ();
 sg13g2_fill_1 FILLER_41_442 ();
 sg13g2_fill_2 FILLER_41_454 ();
 sg13g2_decap_8 FILLER_41_459 ();
 sg13g2_decap_8 FILLER_41_466 ();
 sg13g2_fill_2 FILLER_41_473 ();
 sg13g2_fill_1 FILLER_41_475 ();
 sg13g2_fill_1 FILLER_41_485 ();
 sg13g2_decap_8 FILLER_41_496 ();
 sg13g2_decap_8 FILLER_41_503 ();
 sg13g2_decap_4 FILLER_41_510 ();
 sg13g2_fill_1 FILLER_41_514 ();
 sg13g2_decap_8 FILLER_41_528 ();
 sg13g2_fill_2 FILLER_41_535 ();
 sg13g2_fill_1 FILLER_41_537 ();
 sg13g2_fill_1 FILLER_41_549 ();
 sg13g2_decap_8 FILLER_41_554 ();
 sg13g2_decap_8 FILLER_41_565 ();
 sg13g2_fill_1 FILLER_41_581 ();
 sg13g2_fill_2 FILLER_41_586 ();
 sg13g2_fill_2 FILLER_41_598 ();
 sg13g2_fill_1 FILLER_41_600 ();
 sg13g2_decap_4 FILLER_41_624 ();
 sg13g2_fill_1 FILLER_41_649 ();
 sg13g2_decap_8 FILLER_41_662 ();
 sg13g2_decap_8 FILLER_41_669 ();
 sg13g2_fill_2 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_716 ();
 sg13g2_fill_1 FILLER_41_722 ();
 sg13g2_fill_1 FILLER_41_731 ();
 sg13g2_fill_2 FILLER_41_737 ();
 sg13g2_fill_1 FILLER_41_739 ();
 sg13g2_decap_4 FILLER_41_744 ();
 sg13g2_fill_1 FILLER_41_748 ();
 sg13g2_decap_4 FILLER_41_764 ();
 sg13g2_fill_1 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_796 ();
 sg13g2_fill_2 FILLER_41_803 ();
 sg13g2_fill_1 FILLER_41_805 ();
 sg13g2_fill_2 FILLER_41_828 ();
 sg13g2_fill_2 FILLER_41_834 ();
 sg13g2_fill_1 FILLER_41_836 ();
 sg13g2_decap_4 FILLER_41_842 ();
 sg13g2_fill_1 FILLER_41_854 ();
 sg13g2_fill_2 FILLER_41_882 ();
 sg13g2_fill_1 FILLER_41_893 ();
 sg13g2_decap_4 FILLER_41_913 ();
 sg13g2_fill_1 FILLER_41_926 ();
 sg13g2_decap_4 FILLER_41_930 ();
 sg13g2_decap_8 FILLER_41_938 ();
 sg13g2_decap_4 FILLER_41_945 ();
 sg13g2_fill_2 FILLER_41_949 ();
 sg13g2_fill_1 FILLER_41_956 ();
 sg13g2_decap_4 FILLER_41_965 ();
 sg13g2_fill_2 FILLER_41_969 ();
 sg13g2_fill_1 FILLER_41_1010 ();
 sg13g2_fill_2 FILLER_41_1015 ();
 sg13g2_fill_1 FILLER_41_1025 ();
 sg13g2_fill_1 FILLER_41_1031 ();
 sg13g2_fill_1 FILLER_41_1037 ();
 sg13g2_decap_4 FILLER_41_1046 ();
 sg13g2_fill_1 FILLER_41_1050 ();
 sg13g2_fill_2 FILLER_41_1063 ();
 sg13g2_decap_4 FILLER_41_1071 ();
 sg13g2_fill_1 FILLER_41_1075 ();
 sg13g2_decap_4 FILLER_41_1105 ();
 sg13g2_fill_1 FILLER_41_1109 ();
 sg13g2_decap_4 FILLER_41_1113 ();
 sg13g2_fill_2 FILLER_41_1117 ();
 sg13g2_decap_4 FILLER_41_1148 ();
 sg13g2_fill_2 FILLER_41_1157 ();
 sg13g2_fill_1 FILLER_41_1159 ();
 sg13g2_fill_1 FILLER_41_1175 ();
 sg13g2_fill_2 FILLER_41_1185 ();
 sg13g2_fill_1 FILLER_41_1211 ();
 sg13g2_fill_2 FILLER_41_1217 ();
 sg13g2_fill_2 FILLER_41_1224 ();
 sg13g2_fill_2 FILLER_41_1230 ();
 sg13g2_decap_8 FILLER_41_1237 ();
 sg13g2_decap_4 FILLER_41_1244 ();
 sg13g2_fill_2 FILLER_41_1248 ();
 sg13g2_decap_8 FILLER_41_1270 ();
 sg13g2_fill_1 FILLER_41_1277 ();
 sg13g2_fill_1 FILLER_41_1309 ();
 sg13g2_decap_8 FILLER_41_1314 ();
 sg13g2_decap_4 FILLER_41_1321 ();
 sg13g2_fill_1 FILLER_41_1325 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_decap_4 FILLER_42_30 ();
 sg13g2_decap_8 FILLER_42_39 ();
 sg13g2_decap_4 FILLER_42_46 ();
 sg13g2_fill_1 FILLER_42_50 ();
 sg13g2_decap_4 FILLER_42_55 ();
 sg13g2_fill_1 FILLER_42_59 ();
 sg13g2_fill_2 FILLER_42_69 ();
 sg13g2_decap_8 FILLER_42_75 ();
 sg13g2_decap_4 FILLER_42_82 ();
 sg13g2_fill_1 FILLER_42_95 ();
 sg13g2_fill_1 FILLER_42_106 ();
 sg13g2_fill_1 FILLER_42_155 ();
 sg13g2_decap_8 FILLER_42_165 ();
 sg13g2_fill_2 FILLER_42_172 ();
 sg13g2_decap_8 FILLER_42_177 ();
 sg13g2_fill_2 FILLER_42_184 ();
 sg13g2_fill_1 FILLER_42_186 ();
 sg13g2_fill_2 FILLER_42_203 ();
 sg13g2_fill_2 FILLER_42_217 ();
 sg13g2_fill_1 FILLER_42_219 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_fill_1 FILLER_42_231 ();
 sg13g2_fill_2 FILLER_42_235 ();
 sg13g2_fill_1 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_255 ();
 sg13g2_decap_4 FILLER_42_262 ();
 sg13g2_decap_8 FILLER_42_281 ();
 sg13g2_decap_8 FILLER_42_288 ();
 sg13g2_fill_2 FILLER_42_295 ();
 sg13g2_fill_1 FILLER_42_310 ();
 sg13g2_fill_2 FILLER_42_317 ();
 sg13g2_decap_8 FILLER_42_323 ();
 sg13g2_decap_4 FILLER_42_330 ();
 sg13g2_decap_8 FILLER_42_337 ();
 sg13g2_fill_2 FILLER_42_344 ();
 sg13g2_fill_1 FILLER_42_346 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_fill_2 FILLER_42_375 ();
 sg13g2_fill_1 FILLER_42_393 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_414 ();
 sg13g2_decap_4 FILLER_42_421 ();
 sg13g2_fill_2 FILLER_42_431 ();
 sg13g2_fill_2 FILLER_42_441 ();
 sg13g2_fill_2 FILLER_42_448 ();
 sg13g2_fill_2 FILLER_42_455 ();
 sg13g2_fill_1 FILLER_42_457 ();
 sg13g2_decap_4 FILLER_42_463 ();
 sg13g2_decap_8 FILLER_42_482 ();
 sg13g2_decap_8 FILLER_42_489 ();
 sg13g2_decap_8 FILLER_42_496 ();
 sg13g2_decap_8 FILLER_42_503 ();
 sg13g2_fill_1 FILLER_42_510 ();
 sg13g2_fill_2 FILLER_42_519 ();
 sg13g2_fill_1 FILLER_42_521 ();
 sg13g2_decap_8 FILLER_42_527 ();
 sg13g2_fill_2 FILLER_42_534 ();
 sg13g2_fill_1 FILLER_42_536 ();
 sg13g2_fill_1 FILLER_42_542 ();
 sg13g2_fill_2 FILLER_42_548 ();
 sg13g2_fill_1 FILLER_42_550 ();
 sg13g2_decap_8 FILLER_42_556 ();
 sg13g2_decap_8 FILLER_42_563 ();
 sg13g2_fill_1 FILLER_42_570 ();
 sg13g2_fill_2 FILLER_42_581 ();
 sg13g2_decap_4 FILLER_42_592 ();
 sg13g2_fill_2 FILLER_42_601 ();
 sg13g2_fill_1 FILLER_42_603 ();
 sg13g2_decap_8 FILLER_42_610 ();
 sg13g2_decap_8 FILLER_42_621 ();
 sg13g2_decap_4 FILLER_42_628 ();
 sg13g2_fill_2 FILLER_42_632 ();
 sg13g2_fill_2 FILLER_42_644 ();
 sg13g2_fill_2 FILLER_42_651 ();
 sg13g2_fill_1 FILLER_42_653 ();
 sg13g2_decap_4 FILLER_42_661 ();
 sg13g2_decap_8 FILLER_42_704 ();
 sg13g2_decap_8 FILLER_42_711 ();
 sg13g2_decap_8 FILLER_42_718 ();
 sg13g2_fill_2 FILLER_42_725 ();
 sg13g2_fill_1 FILLER_42_731 ();
 sg13g2_decap_8 FILLER_42_744 ();
 sg13g2_decap_4 FILLER_42_751 ();
 sg13g2_fill_1 FILLER_42_755 ();
 sg13g2_fill_2 FILLER_42_772 ();
 sg13g2_decap_8 FILLER_42_796 ();
 sg13g2_decap_4 FILLER_42_803 ();
 sg13g2_fill_2 FILLER_42_807 ();
 sg13g2_fill_2 FILLER_42_836 ();
 sg13g2_decap_8 FILLER_42_847 ();
 sg13g2_decap_4 FILLER_42_854 ();
 sg13g2_fill_1 FILLER_42_897 ();
 sg13g2_fill_1 FILLER_42_901 ();
 sg13g2_fill_1 FILLER_42_911 ();
 sg13g2_fill_2 FILLER_42_934 ();
 sg13g2_fill_1 FILLER_42_939 ();
 sg13g2_decap_8 FILLER_42_953 ();
 sg13g2_decap_8 FILLER_42_960 ();
 sg13g2_fill_2 FILLER_42_967 ();
 sg13g2_fill_1 FILLER_42_978 ();
 sg13g2_fill_2 FILLER_42_996 ();
 sg13g2_decap_8 FILLER_42_1015 ();
 sg13g2_decap_4 FILLER_42_1022 ();
 sg13g2_fill_1 FILLER_42_1026 ();
 sg13g2_decap_8 FILLER_42_1030 ();
 sg13g2_fill_2 FILLER_42_1037 ();
 sg13g2_decap_8 FILLER_42_1044 ();
 sg13g2_decap_4 FILLER_42_1051 ();
 sg13g2_fill_2 FILLER_42_1055 ();
 sg13g2_fill_2 FILLER_42_1061 ();
 sg13g2_decap_8 FILLER_42_1072 ();
 sg13g2_decap_8 FILLER_42_1079 ();
 sg13g2_fill_1 FILLER_42_1086 ();
 sg13g2_decap_4 FILLER_42_1091 ();
 sg13g2_fill_2 FILLER_42_1095 ();
 sg13g2_fill_2 FILLER_42_1102 ();
 sg13g2_fill_2 FILLER_42_1109 ();
 sg13g2_fill_2 FILLER_42_1115 ();
 sg13g2_fill_1 FILLER_42_1117 ();
 sg13g2_decap_8 FILLER_42_1123 ();
 sg13g2_fill_2 FILLER_42_1130 ();
 sg13g2_fill_1 FILLER_42_1168 ();
 sg13g2_decap_8 FILLER_42_1173 ();
 sg13g2_decap_8 FILLER_42_1180 ();
 sg13g2_fill_1 FILLER_42_1193 ();
 sg13g2_fill_1 FILLER_42_1210 ();
 sg13g2_decap_4 FILLER_42_1232 ();
 sg13g2_fill_1 FILLER_42_1236 ();
 sg13g2_decap_4 FILLER_42_1245 ();
 sg13g2_fill_2 FILLER_42_1263 ();
 sg13g2_fill_2 FILLER_42_1282 ();
 sg13g2_decap_8 FILLER_42_1288 ();
 sg13g2_fill_1 FILLER_42_1295 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_24 ();
 sg13g2_fill_1 FILLER_43_51 ();
 sg13g2_fill_1 FILLER_43_78 ();
 sg13g2_fill_1 FILLER_43_94 ();
 sg13g2_fill_2 FILLER_43_105 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_decap_8 FILLER_43_180 ();
 sg13g2_fill_1 FILLER_43_187 ();
 sg13g2_fill_1 FILLER_43_205 ();
 sg13g2_fill_2 FILLER_43_212 ();
 sg13g2_fill_2 FILLER_43_230 ();
 sg13g2_fill_2 FILLER_43_241 ();
 sg13g2_decap_8 FILLER_43_248 ();
 sg13g2_fill_1 FILLER_43_258 ();
 sg13g2_decap_8 FILLER_43_268 ();
 sg13g2_decap_8 FILLER_43_275 ();
 sg13g2_decap_4 FILLER_43_282 ();
 sg13g2_decap_8 FILLER_43_289 ();
 sg13g2_decap_8 FILLER_43_296 ();
 sg13g2_decap_8 FILLER_43_303 ();
 sg13g2_fill_1 FILLER_43_310 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_4 FILLER_43_322 ();
 sg13g2_fill_2 FILLER_43_345 ();
 sg13g2_fill_1 FILLER_43_347 ();
 sg13g2_fill_2 FILLER_43_359 ();
 sg13g2_decap_4 FILLER_43_364 ();
 sg13g2_fill_1 FILLER_43_368 ();
 sg13g2_decap_8 FILLER_43_374 ();
 sg13g2_fill_1 FILLER_43_381 ();
 sg13g2_decap_8 FILLER_43_394 ();
 sg13g2_decap_8 FILLER_43_401 ();
 sg13g2_decap_4 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_43_417 ();
 sg13g2_fill_2 FILLER_43_430 ();
 sg13g2_decap_4 FILLER_43_438 ();
 sg13g2_fill_1 FILLER_43_442 ();
 sg13g2_fill_1 FILLER_43_449 ();
 sg13g2_fill_1 FILLER_43_470 ();
 sg13g2_decap_4 FILLER_43_504 ();
 sg13g2_fill_1 FILLER_43_508 ();
 sg13g2_decap_4 FILLER_43_519 ();
 sg13g2_fill_2 FILLER_43_523 ();
 sg13g2_decap_8 FILLER_43_536 ();
 sg13g2_decap_4 FILLER_43_543 ();
 sg13g2_fill_1 FILLER_43_547 ();
 sg13g2_fill_1 FILLER_43_555 ();
 sg13g2_fill_2 FILLER_43_561 ();
 sg13g2_fill_1 FILLER_43_563 ();
 sg13g2_fill_1 FILLER_43_587 ();
 sg13g2_fill_2 FILLER_43_592 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_4 FILLER_43_609 ();
 sg13g2_fill_2 FILLER_43_613 ();
 sg13g2_fill_1 FILLER_43_619 ();
 sg13g2_fill_1 FILLER_43_623 ();
 sg13g2_fill_1 FILLER_43_628 ();
 sg13g2_fill_1 FILLER_43_634 ();
 sg13g2_fill_2 FILLER_43_640 ();
 sg13g2_fill_2 FILLER_43_646 ();
 sg13g2_fill_1 FILLER_43_648 ();
 sg13g2_decap_8 FILLER_43_653 ();
 sg13g2_decap_8 FILLER_43_673 ();
 sg13g2_fill_2 FILLER_43_680 ();
 sg13g2_decap_8 FILLER_43_690 ();
 sg13g2_decap_8 FILLER_43_697 ();
 sg13g2_decap_8 FILLER_43_704 ();
 sg13g2_decap_4 FILLER_43_711 ();
 sg13g2_fill_1 FILLER_43_715 ();
 sg13g2_decap_8 FILLER_43_728 ();
 sg13g2_decap_4 FILLER_43_735 ();
 sg13g2_fill_2 FILLER_43_739 ();
 sg13g2_decap_8 FILLER_43_744 ();
 sg13g2_decap_8 FILLER_43_751 ();
 sg13g2_fill_2 FILLER_43_758 ();
 sg13g2_fill_1 FILLER_43_760 ();
 sg13g2_fill_1 FILLER_43_767 ();
 sg13g2_fill_1 FILLER_43_779 ();
 sg13g2_decap_4 FILLER_43_793 ();
 sg13g2_fill_2 FILLER_43_797 ();
 sg13g2_fill_1 FILLER_43_819 ();
 sg13g2_fill_2 FILLER_43_825 ();
 sg13g2_decap_8 FILLER_43_846 ();
 sg13g2_fill_2 FILLER_43_857 ();
 sg13g2_fill_1 FILLER_43_859 ();
 sg13g2_fill_2 FILLER_43_864 ();
 sg13g2_fill_1 FILLER_43_866 ();
 sg13g2_decap_4 FILLER_43_870 ();
 sg13g2_fill_2 FILLER_43_878 ();
 sg13g2_fill_1 FILLER_43_880 ();
 sg13g2_fill_1 FILLER_43_884 ();
 sg13g2_decap_4 FILLER_43_889 ();
 sg13g2_fill_1 FILLER_43_916 ();
 sg13g2_fill_2 FILLER_43_942 ();
 sg13g2_fill_1 FILLER_43_944 ();
 sg13g2_decap_4 FILLER_43_950 ();
 sg13g2_fill_1 FILLER_43_954 ();
 sg13g2_decap_8 FILLER_43_960 ();
 sg13g2_decap_8 FILLER_43_967 ();
 sg13g2_fill_2 FILLER_43_974 ();
 sg13g2_fill_1 FILLER_43_976 ();
 sg13g2_fill_1 FILLER_43_990 ();
 sg13g2_fill_1 FILLER_43_996 ();
 sg13g2_fill_1 FILLER_43_1007 ();
 sg13g2_decap_8 FILLER_43_1034 ();
 sg13g2_decap_8 FILLER_43_1041 ();
 sg13g2_decap_4 FILLER_43_1048 ();
 sg13g2_fill_1 FILLER_43_1052 ();
 sg13g2_decap_4 FILLER_43_1079 ();
 sg13g2_decap_8 FILLER_43_1088 ();
 sg13g2_fill_2 FILLER_43_1095 ();
 sg13g2_fill_1 FILLER_43_1104 ();
 sg13g2_decap_8 FILLER_43_1115 ();
 sg13g2_fill_1 FILLER_43_1122 ();
 sg13g2_decap_8 FILLER_43_1152 ();
 sg13g2_fill_2 FILLER_43_1159 ();
 sg13g2_decap_8 FILLER_43_1164 ();
 sg13g2_decap_8 FILLER_43_1171 ();
 sg13g2_decap_4 FILLER_43_1178 ();
 sg13g2_fill_2 FILLER_43_1200 ();
 sg13g2_fill_2 FILLER_43_1218 ();
 sg13g2_fill_1 FILLER_43_1220 ();
 sg13g2_decap_4 FILLER_43_1247 ();
 sg13g2_fill_1 FILLER_43_1251 ();
 sg13g2_fill_2 FILLER_43_1256 ();
 sg13g2_decap_4 FILLER_43_1290 ();
 sg13g2_fill_1 FILLER_43_1294 ();
 sg13g2_decap_8 FILLER_43_1300 ();
 sg13g2_decap_8 FILLER_43_1307 ();
 sg13g2_decap_8 FILLER_43_1314 ();
 sg13g2_decap_4 FILLER_43_1321 ();
 sg13g2_fill_1 FILLER_43_1325 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_7 ();
 sg13g2_fill_1 FILLER_44_9 ();
 sg13g2_decap_8 FILLER_44_19 ();
 sg13g2_decap_4 FILLER_44_26 ();
 sg13g2_fill_2 FILLER_44_30 ();
 sg13g2_fill_2 FILLER_44_37 ();
 sg13g2_decap_8 FILLER_44_43 ();
 sg13g2_decap_8 FILLER_44_50 ();
 sg13g2_fill_1 FILLER_44_57 ();
 sg13g2_fill_1 FILLER_44_62 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_4 FILLER_44_84 ();
 sg13g2_fill_1 FILLER_44_95 ();
 sg13g2_fill_1 FILLER_44_118 ();
 sg13g2_fill_2 FILLER_44_125 ();
 sg13g2_fill_2 FILLER_44_132 ();
 sg13g2_fill_1 FILLER_44_134 ();
 sg13g2_fill_2 FILLER_44_146 ();
 sg13g2_fill_2 FILLER_44_166 ();
 sg13g2_fill_1 FILLER_44_168 ();
 sg13g2_fill_1 FILLER_44_190 ();
 sg13g2_fill_1 FILLER_44_200 ();
 sg13g2_fill_1 FILLER_44_214 ();
 sg13g2_fill_1 FILLER_44_223 ();
 sg13g2_fill_2 FILLER_44_235 ();
 sg13g2_fill_2 FILLER_44_244 ();
 sg13g2_decap_8 FILLER_44_251 ();
 sg13g2_fill_1 FILLER_44_258 ();
 sg13g2_fill_2 FILLER_44_270 ();
 sg13g2_fill_2 FILLER_44_277 ();
 sg13g2_decap_4 FILLER_44_292 ();
 sg13g2_decap_4 FILLER_44_300 ();
 sg13g2_decap_8 FILLER_44_321 ();
 sg13g2_decap_8 FILLER_44_328 ();
 sg13g2_decap_4 FILLER_44_335 ();
 sg13g2_fill_2 FILLER_44_344 ();
 sg13g2_fill_1 FILLER_44_346 ();
 sg13g2_decap_4 FILLER_44_352 ();
 sg13g2_fill_2 FILLER_44_356 ();
 sg13g2_fill_2 FILLER_44_373 ();
 sg13g2_fill_2 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_44_416 ();
 sg13g2_decap_8 FILLER_44_423 ();
 sg13g2_decap_8 FILLER_44_430 ();
 sg13g2_decap_8 FILLER_44_437 ();
 sg13g2_fill_2 FILLER_44_448 ();
 sg13g2_fill_2 FILLER_44_454 ();
 sg13g2_fill_2 FILLER_44_476 ();
 sg13g2_fill_1 FILLER_44_487 ();
 sg13g2_decap_8 FILLER_44_497 ();
 sg13g2_fill_2 FILLER_44_504 ();
 sg13g2_fill_1 FILLER_44_506 ();
 sg13g2_fill_1 FILLER_44_519 ();
 sg13g2_fill_1 FILLER_44_533 ();
 sg13g2_decap_4 FILLER_44_544 ();
 sg13g2_fill_1 FILLER_44_548 ();
 sg13g2_decap_4 FILLER_44_554 ();
 sg13g2_fill_2 FILLER_44_558 ();
 sg13g2_fill_2 FILLER_44_565 ();
 sg13g2_fill_1 FILLER_44_567 ();
 sg13g2_fill_2 FILLER_44_575 ();
 sg13g2_fill_1 FILLER_44_577 ();
 sg13g2_fill_1 FILLER_44_588 ();
 sg13g2_fill_1 FILLER_44_592 ();
 sg13g2_decap_8 FILLER_44_606 ();
 sg13g2_decap_4 FILLER_44_613 ();
 sg13g2_fill_1 FILLER_44_621 ();
 sg13g2_fill_1 FILLER_44_627 ();
 sg13g2_fill_1 FILLER_44_634 ();
 sg13g2_decap_8 FILLER_44_648 ();
 sg13g2_decap_8 FILLER_44_655 ();
 sg13g2_decap_8 FILLER_44_701 ();
 sg13g2_decap_4 FILLER_44_708 ();
 sg13g2_fill_2 FILLER_44_712 ();
 sg13g2_fill_2 FILLER_44_727 ();
 sg13g2_decap_8 FILLER_44_751 ();
 sg13g2_decap_8 FILLER_44_764 ();
 sg13g2_decap_8 FILLER_44_780 ();
 sg13g2_decap_8 FILLER_44_787 ();
 sg13g2_fill_2 FILLER_44_794 ();
 sg13g2_fill_1 FILLER_44_796 ();
 sg13g2_decap_4 FILLER_44_806 ();
 sg13g2_fill_2 FILLER_44_813 ();
 sg13g2_fill_1 FILLER_44_815 ();
 sg13g2_decap_4 FILLER_44_820 ();
 sg13g2_decap_8 FILLER_44_829 ();
 sg13g2_decap_4 FILLER_44_839 ();
 sg13g2_fill_2 FILLER_44_848 ();
 sg13g2_fill_1 FILLER_44_850 ();
 sg13g2_decap_4 FILLER_44_855 ();
 sg13g2_decap_8 FILLER_44_865 ();
 sg13g2_decap_8 FILLER_44_872 ();
 sg13g2_decap_8 FILLER_44_879 ();
 sg13g2_decap_8 FILLER_44_886 ();
 sg13g2_fill_2 FILLER_44_893 ();
 sg13g2_fill_1 FILLER_44_895 ();
 sg13g2_decap_8 FILLER_44_913 ();
 sg13g2_decap_8 FILLER_44_920 ();
 sg13g2_fill_1 FILLER_44_927 ();
 sg13g2_decap_8 FILLER_44_937 ();
 sg13g2_fill_1 FILLER_44_944 ();
 sg13g2_fill_1 FILLER_44_952 ();
 sg13g2_fill_2 FILLER_44_964 ();
 sg13g2_decap_8 FILLER_44_973 ();
 sg13g2_decap_4 FILLER_44_980 ();
 sg13g2_fill_1 FILLER_44_988 ();
 sg13g2_decap_4 FILLER_44_998 ();
 sg13g2_fill_1 FILLER_44_1002 ();
 sg13g2_fill_1 FILLER_44_1006 ();
 sg13g2_decap_4 FILLER_44_1026 ();
 sg13g2_decap_4 FILLER_44_1034 ();
 sg13g2_fill_1 FILLER_44_1038 ();
 sg13g2_fill_1 FILLER_44_1044 ();
 sg13g2_decap_4 FILLER_44_1091 ();
 sg13g2_fill_1 FILLER_44_1095 ();
 sg13g2_fill_1 FILLER_44_1104 ();
 sg13g2_fill_1 FILLER_44_1125 ();
 sg13g2_fill_1 FILLER_44_1134 ();
 sg13g2_fill_2 FILLER_44_1138 ();
 sg13g2_fill_1 FILLER_44_1140 ();
 sg13g2_fill_2 FILLER_44_1167 ();
 sg13g2_fill_1 FILLER_44_1169 ();
 sg13g2_decap_4 FILLER_44_1175 ();
 sg13g2_fill_1 FILLER_44_1179 ();
 sg13g2_fill_2 FILLER_44_1185 ();
 sg13g2_fill_2 FILLER_44_1191 ();
 sg13g2_fill_1 FILLER_44_1196 ();
 sg13g2_fill_2 FILLER_44_1224 ();
 sg13g2_fill_1 FILLER_44_1226 ();
 sg13g2_decap_4 FILLER_44_1232 ();
 sg13g2_decap_8 FILLER_44_1239 ();
 sg13g2_decap_8 FILLER_44_1246 ();
 sg13g2_fill_1 FILLER_44_1275 ();
 sg13g2_decap_4 FILLER_44_1281 ();
 sg13g2_decap_4 FILLER_44_1290 ();
 sg13g2_fill_2 FILLER_44_1294 ();
 sg13g2_decap_8 FILLER_44_1305 ();
 sg13g2_decap_8 FILLER_44_1312 ();
 sg13g2_decap_8 FILLER_44_1319 ();
 sg13g2_decap_4 FILLER_45_26 ();
 sg13g2_decap_4 FILLER_45_56 ();
 sg13g2_fill_1 FILLER_45_60 ();
 sg13g2_fill_2 FILLER_45_72 ();
 sg13g2_decap_8 FILLER_45_78 ();
 sg13g2_decap_4 FILLER_45_85 ();
 sg13g2_fill_2 FILLER_45_89 ();
 sg13g2_fill_1 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_101 ();
 sg13g2_fill_1 FILLER_45_103 ();
 sg13g2_fill_2 FILLER_45_117 ();
 sg13g2_fill_1 FILLER_45_123 ();
 sg13g2_fill_2 FILLER_45_129 ();
 sg13g2_fill_1 FILLER_45_136 ();
 sg13g2_fill_2 FILLER_45_143 ();
 sg13g2_fill_2 FILLER_45_155 ();
 sg13g2_fill_2 FILLER_45_163 ();
 sg13g2_fill_1 FILLER_45_165 ();
 sg13g2_decap_8 FILLER_45_170 ();
 sg13g2_fill_2 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_234 ();
 sg13g2_fill_2 FILLER_45_238 ();
 sg13g2_fill_1 FILLER_45_240 ();
 sg13g2_fill_1 FILLER_45_246 ();
 sg13g2_fill_1 FILLER_45_252 ();
 sg13g2_fill_1 FILLER_45_262 ();
 sg13g2_fill_2 FILLER_45_272 ();
 sg13g2_fill_1 FILLER_45_279 ();
 sg13g2_decap_8 FILLER_45_289 ();
 sg13g2_decap_4 FILLER_45_296 ();
 sg13g2_fill_2 FILLER_45_300 ();
 sg13g2_fill_2 FILLER_45_310 ();
 sg13g2_fill_2 FILLER_45_325 ();
 sg13g2_decap_8 FILLER_45_335 ();
 sg13g2_fill_1 FILLER_45_342 ();
 sg13g2_decap_8 FILLER_45_347 ();
 sg13g2_decap_4 FILLER_45_354 ();
 sg13g2_fill_1 FILLER_45_358 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_382 ();
 sg13g2_decap_4 FILLER_45_389 ();
 sg13g2_fill_2 FILLER_45_393 ();
 sg13g2_decap_4 FILLER_45_400 ();
 sg13g2_fill_1 FILLER_45_404 ();
 sg13g2_decap_8 FILLER_45_415 ();
 sg13g2_decap_4 FILLER_45_422 ();
 sg13g2_fill_2 FILLER_45_437 ();
 sg13g2_fill_1 FILLER_45_439 ();
 sg13g2_decap_8 FILLER_45_445 ();
 sg13g2_decap_8 FILLER_45_452 ();
 sg13g2_fill_2 FILLER_45_474 ();
 sg13g2_fill_1 FILLER_45_476 ();
 sg13g2_fill_2 FILLER_45_486 ();
 sg13g2_fill_1 FILLER_45_488 ();
 sg13g2_decap_4 FILLER_45_508 ();
 sg13g2_fill_2 FILLER_45_517 ();
 sg13g2_decap_4 FILLER_45_528 ();
 sg13g2_fill_2 FILLER_45_543 ();
 sg13g2_decap_4 FILLER_45_548 ();
 sg13g2_fill_1 FILLER_45_567 ();
 sg13g2_fill_1 FILLER_45_574 ();
 sg13g2_fill_1 FILLER_45_580 ();
 sg13g2_fill_1 FILLER_45_589 ();
 sg13g2_fill_2 FILLER_45_595 ();
 sg13g2_decap_8 FILLER_45_605 ();
 sg13g2_decap_8 FILLER_45_612 ();
 sg13g2_decap_8 FILLER_45_619 ();
 sg13g2_decap_8 FILLER_45_626 ();
 sg13g2_decap_8 FILLER_45_633 ();
 sg13g2_fill_2 FILLER_45_640 ();
 sg13g2_fill_1 FILLER_45_642 ();
 sg13g2_decap_8 FILLER_45_647 ();
 sg13g2_decap_8 FILLER_45_654 ();
 sg13g2_decap_8 FILLER_45_661 ();
 sg13g2_decap_4 FILLER_45_671 ();
 sg13g2_fill_2 FILLER_45_675 ();
 sg13g2_decap_8 FILLER_45_687 ();
 sg13g2_fill_1 FILLER_45_694 ();
 sg13g2_decap_8 FILLER_45_699 ();
 sg13g2_fill_1 FILLER_45_706 ();
 sg13g2_fill_1 FILLER_45_718 ();
 sg13g2_decap_8 FILLER_45_730 ();
 sg13g2_fill_1 FILLER_45_737 ();
 sg13g2_decap_8 FILLER_45_747 ();
 sg13g2_fill_2 FILLER_45_754 ();
 sg13g2_decap_8 FILLER_45_762 ();
 sg13g2_decap_4 FILLER_45_769 ();
 sg13g2_fill_1 FILLER_45_773 ();
 sg13g2_decap_8 FILLER_45_790 ();
 sg13g2_decap_8 FILLER_45_797 ();
 sg13g2_decap_8 FILLER_45_804 ();
 sg13g2_fill_2 FILLER_45_811 ();
 sg13g2_fill_1 FILLER_45_825 ();
 sg13g2_fill_2 FILLER_45_830 ();
 sg13g2_fill_1 FILLER_45_836 ();
 sg13g2_fill_2 FILLER_45_841 ();
 sg13g2_fill_1 FILLER_45_847 ();
 sg13g2_decap_8 FILLER_45_854 ();
 sg13g2_fill_2 FILLER_45_861 ();
 sg13g2_fill_1 FILLER_45_863 ();
 sg13g2_fill_2 FILLER_45_871 ();
 sg13g2_fill_2 FILLER_45_879 ();
 sg13g2_fill_1 FILLER_45_881 ();
 sg13g2_decap_4 FILLER_45_888 ();
 sg13g2_fill_1 FILLER_45_892 ();
 sg13g2_fill_2 FILLER_45_898 ();
 sg13g2_fill_1 FILLER_45_900 ();
 sg13g2_fill_1 FILLER_45_907 ();
 sg13g2_fill_1 FILLER_45_913 ();
 sg13g2_fill_1 FILLER_45_928 ();
 sg13g2_decap_8 FILLER_45_933 ();
 sg13g2_fill_2 FILLER_45_940 ();
 sg13g2_decap_8 FILLER_45_945 ();
 sg13g2_fill_2 FILLER_45_952 ();
 sg13g2_fill_1 FILLER_45_954 ();
 sg13g2_decap_8 FILLER_45_965 ();
 sg13g2_fill_2 FILLER_45_972 ();
 sg13g2_decap_4 FILLER_45_985 ();
 sg13g2_decap_8 FILLER_45_1008 ();
 sg13g2_decap_8 FILLER_45_1015 ();
 sg13g2_decap_4 FILLER_45_1022 ();
 sg13g2_decap_8 FILLER_45_1030 ();
 sg13g2_fill_2 FILLER_45_1037 ();
 sg13g2_decap_4 FILLER_45_1044 ();
 sg13g2_fill_2 FILLER_45_1056 ();
 sg13g2_fill_1 FILLER_45_1058 ();
 sg13g2_decap_8 FILLER_45_1076 ();
 sg13g2_fill_2 FILLER_45_1083 ();
 sg13g2_fill_2 FILLER_45_1091 ();
 sg13g2_decap_8 FILLER_45_1112 ();
 sg13g2_decap_4 FILLER_45_1119 ();
 sg13g2_decap_4 FILLER_45_1130 ();
 sg13g2_fill_1 FILLER_45_1134 ();
 sg13g2_decap_8 FILLER_45_1143 ();
 sg13g2_decap_8 FILLER_45_1150 ();
 sg13g2_decap_4 FILLER_45_1157 ();
 sg13g2_decap_8 FILLER_45_1168 ();
 sg13g2_decap_8 FILLER_45_1175 ();
 sg13g2_fill_1 FILLER_45_1182 ();
 sg13g2_fill_1 FILLER_45_1200 ();
 sg13g2_fill_1 FILLER_45_1236 ();
 sg13g2_fill_1 FILLER_45_1243 ();
 sg13g2_fill_1 FILLER_45_1251 ();
 sg13g2_fill_2 FILLER_45_1260 ();
 sg13g2_decap_8 FILLER_45_1279 ();
 sg13g2_fill_2 FILLER_45_1286 ();
 sg13g2_fill_1 FILLER_45_1288 ();
 sg13g2_decap_4 FILLER_45_1293 ();
 sg13g2_fill_1 FILLER_45_1297 ();
 sg13g2_fill_2 FILLER_45_1324 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_14 ();
 sg13g2_fill_1 FILLER_46_16 ();
 sg13g2_fill_1 FILLER_46_22 ();
 sg13g2_fill_2 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_37 ();
 sg13g2_decap_8 FILLER_46_50 ();
 sg13g2_decap_4 FILLER_46_57 ();
 sg13g2_fill_1 FILLER_46_69 ();
 sg13g2_fill_2 FILLER_46_73 ();
 sg13g2_fill_1 FILLER_46_75 ();
 sg13g2_decap_4 FILLER_46_105 ();
 sg13g2_fill_2 FILLER_46_109 ();
 sg13g2_fill_2 FILLER_46_121 ();
 sg13g2_fill_1 FILLER_46_123 ();
 sg13g2_decap_8 FILLER_46_128 ();
 sg13g2_fill_1 FILLER_46_144 ();
 sg13g2_decap_8 FILLER_46_157 ();
 sg13g2_fill_1 FILLER_46_164 ();
 sg13g2_fill_2 FILLER_46_169 ();
 sg13g2_fill_1 FILLER_46_171 ();
 sg13g2_decap_8 FILLER_46_181 ();
 sg13g2_decap_8 FILLER_46_188 ();
 sg13g2_fill_1 FILLER_46_195 ();
 sg13g2_decap_4 FILLER_46_200 ();
 sg13g2_fill_2 FILLER_46_204 ();
 sg13g2_fill_2 FILLER_46_212 ();
 sg13g2_fill_1 FILLER_46_214 ();
 sg13g2_fill_1 FILLER_46_220 ();
 sg13g2_decap_4 FILLER_46_225 ();
 sg13g2_fill_2 FILLER_46_229 ();
 sg13g2_decap_4 FILLER_46_244 ();
 sg13g2_decap_4 FILLER_46_262 ();
 sg13g2_fill_1 FILLER_46_266 ();
 sg13g2_fill_1 FILLER_46_275 ();
 sg13g2_fill_1 FILLER_46_280 ();
 sg13g2_fill_1 FILLER_46_286 ();
 sg13g2_fill_1 FILLER_46_291 ();
 sg13g2_fill_1 FILLER_46_297 ();
 sg13g2_fill_1 FILLER_46_307 ();
 sg13g2_fill_2 FILLER_46_315 ();
 sg13g2_fill_2 FILLER_46_322 ();
 sg13g2_fill_1 FILLER_46_324 ();
 sg13g2_fill_2 FILLER_46_341 ();
 sg13g2_fill_2 FILLER_46_347 ();
 sg13g2_fill_1 FILLER_46_349 ();
 sg13g2_fill_2 FILLER_46_359 ();
 sg13g2_decap_8 FILLER_46_369 ();
 sg13g2_decap_8 FILLER_46_376 ();
 sg13g2_decap_4 FILLER_46_383 ();
 sg13g2_fill_2 FILLER_46_390 ();
 sg13g2_fill_1 FILLER_46_392 ();
 sg13g2_decap_4 FILLER_46_400 ();
 sg13g2_fill_2 FILLER_46_404 ();
 sg13g2_fill_2 FILLER_46_422 ();
 sg13g2_fill_1 FILLER_46_424 ();
 sg13g2_fill_2 FILLER_46_450 ();
 sg13g2_fill_1 FILLER_46_478 ();
 sg13g2_fill_2 FILLER_46_482 ();
 sg13g2_fill_2 FILLER_46_489 ();
 sg13g2_fill_2 FILLER_46_495 ();
 sg13g2_fill_1 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_510 ();
 sg13g2_fill_2 FILLER_46_517 ();
 sg13g2_fill_1 FILLER_46_519 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_4 FILLER_46_539 ();
 sg13g2_fill_1 FILLER_46_543 ();
 sg13g2_fill_1 FILLER_46_549 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_fill_2 FILLER_46_567 ();
 sg13g2_fill_1 FILLER_46_569 ();
 sg13g2_decap_8 FILLER_46_573 ();
 sg13g2_fill_1 FILLER_46_580 ();
 sg13g2_fill_1 FILLER_46_586 ();
 sg13g2_fill_2 FILLER_46_592 ();
 sg13g2_fill_2 FILLER_46_599 ();
 sg13g2_fill_2 FILLER_46_606 ();
 sg13g2_decap_4 FILLER_46_641 ();
 sg13g2_decap_4 FILLER_46_648 ();
 sg13g2_fill_2 FILLER_46_652 ();
 sg13g2_fill_1 FILLER_46_662 ();
 sg13g2_decap_4 FILLER_46_693 ();
 sg13g2_fill_2 FILLER_46_707 ();
 sg13g2_fill_1 FILLER_46_709 ();
 sg13g2_fill_1 FILLER_46_713 ();
 sg13g2_decap_8 FILLER_46_718 ();
 sg13g2_decap_4 FILLER_46_725 ();
 sg13g2_decap_4 FILLER_46_734 ();
 sg13g2_decap_8 FILLER_46_747 ();
 sg13g2_fill_2 FILLER_46_754 ();
 sg13g2_decap_8 FILLER_46_764 ();
 sg13g2_fill_2 FILLER_46_771 ();
 sg13g2_fill_1 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_837 ();
 sg13g2_decap_8 FILLER_46_844 ();
 sg13g2_decap_8 FILLER_46_851 ();
 sg13g2_decap_8 FILLER_46_858 ();
 sg13g2_decap_8 FILLER_46_872 ();
 sg13g2_decap_8 FILLER_46_879 ();
 sg13g2_decap_8 FILLER_46_886 ();
 sg13g2_fill_2 FILLER_46_893 ();
 sg13g2_fill_1 FILLER_46_895 ();
 sg13g2_fill_2 FILLER_46_905 ();
 sg13g2_decap_8 FILLER_46_919 ();
 sg13g2_fill_2 FILLER_46_926 ();
 sg13g2_fill_1 FILLER_46_928 ();
 sg13g2_decap_4 FILLER_46_935 ();
 sg13g2_fill_2 FILLER_46_946 ();
 sg13g2_fill_2 FILLER_46_957 ();
 sg13g2_fill_2 FILLER_46_969 ();
 sg13g2_fill_2 FILLER_46_974 ();
 sg13g2_fill_1 FILLER_46_983 ();
 sg13g2_fill_1 FILLER_46_988 ();
 sg13g2_decap_8 FILLER_46_993 ();
 sg13g2_fill_1 FILLER_46_1039 ();
 sg13g2_fill_1 FILLER_46_1045 ();
 sg13g2_fill_1 FILLER_46_1051 ();
 sg13g2_decap_8 FILLER_46_1055 ();
 sg13g2_decap_4 FILLER_46_1066 ();
 sg13g2_fill_2 FILLER_46_1075 ();
 sg13g2_fill_1 FILLER_46_1077 ();
 sg13g2_decap_4 FILLER_46_1089 ();
 sg13g2_fill_1 FILLER_46_1093 ();
 sg13g2_fill_2 FILLER_46_1099 ();
 sg13g2_fill_1 FILLER_46_1101 ();
 sg13g2_fill_1 FILLER_46_1111 ();
 sg13g2_fill_2 FILLER_46_1119 ();
 sg13g2_fill_2 FILLER_46_1125 ();
 sg13g2_fill_1 FILLER_46_1127 ();
 sg13g2_fill_1 FILLER_46_1131 ();
 sg13g2_fill_1 FILLER_46_1136 ();
 sg13g2_fill_1 FILLER_46_1147 ();
 sg13g2_fill_1 FILLER_46_1158 ();
 sg13g2_decap_8 FILLER_46_1166 ();
 sg13g2_fill_2 FILLER_46_1181 ();
 sg13g2_fill_2 FILLER_46_1188 ();
 sg13g2_fill_1 FILLER_46_1190 ();
 sg13g2_fill_2 FILLER_46_1196 ();
 sg13g2_fill_1 FILLER_46_1203 ();
 sg13g2_fill_1 FILLER_46_1216 ();
 sg13g2_fill_2 FILLER_46_1242 ();
 sg13g2_decap_8 FILLER_46_1263 ();
 sg13g2_decap_4 FILLER_46_1270 ();
 sg13g2_decap_4 FILLER_46_1291 ();
 sg13g2_fill_2 FILLER_46_1295 ();
 sg13g2_decap_8 FILLER_46_1301 ();
 sg13g2_decap_8 FILLER_46_1312 ();
 sg13g2_decap_8 FILLER_46_1319 ();
 sg13g2_decap_8 FILLER_47_26 ();
 sg13g2_fill_2 FILLER_47_33 ();
 sg13g2_fill_1 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_40 ();
 sg13g2_decap_8 FILLER_47_47 ();
 sg13g2_decap_8 FILLER_47_54 ();
 sg13g2_fill_1 FILLER_47_61 ();
 sg13g2_fill_2 FILLER_47_75 ();
 sg13g2_fill_2 FILLER_47_80 ();
 sg13g2_fill_1 FILLER_47_86 ();
 sg13g2_fill_2 FILLER_47_114 ();
 sg13g2_fill_1 FILLER_47_116 ();
 sg13g2_fill_1 FILLER_47_131 ();
 sg13g2_fill_2 FILLER_47_147 ();
 sg13g2_fill_1 FILLER_47_149 ();
 sg13g2_fill_2 FILLER_47_157 ();
 sg13g2_fill_1 FILLER_47_159 ();
 sg13g2_decap_8 FILLER_47_163 ();
 sg13g2_decap_4 FILLER_47_170 ();
 sg13g2_decap_4 FILLER_47_179 ();
 sg13g2_fill_1 FILLER_47_183 ();
 sg13g2_fill_1 FILLER_47_188 ();
 sg13g2_fill_1 FILLER_47_197 ();
 sg13g2_fill_1 FILLER_47_201 ();
 sg13g2_fill_1 FILLER_47_207 ();
 sg13g2_decap_4 FILLER_47_211 ();
 sg13g2_decap_8 FILLER_47_219 ();
 sg13g2_decap_8 FILLER_47_226 ();
 sg13g2_decap_4 FILLER_47_237 ();
 sg13g2_fill_2 FILLER_47_241 ();
 sg13g2_decap_4 FILLER_47_253 ();
 sg13g2_decap_4 FILLER_47_267 ();
 sg13g2_fill_2 FILLER_47_276 ();
 sg13g2_decap_8 FILLER_47_282 ();
 sg13g2_decap_8 FILLER_47_289 ();
 sg13g2_decap_4 FILLER_47_296 ();
 sg13g2_fill_2 FILLER_47_300 ();
 sg13g2_fill_2 FILLER_47_305 ();
 sg13g2_fill_1 FILLER_47_307 ();
 sg13g2_decap_4 FILLER_47_318 ();
 sg13g2_fill_2 FILLER_47_322 ();
 sg13g2_fill_2 FILLER_47_333 ();
 sg13g2_fill_1 FILLER_47_347 ();
 sg13g2_decap_8 FILLER_47_352 ();
 sg13g2_decap_4 FILLER_47_359 ();
 sg13g2_fill_2 FILLER_47_363 ();
 sg13g2_decap_4 FILLER_47_370 ();
 sg13g2_fill_1 FILLER_47_374 ();
 sg13g2_decap_4 FILLER_47_383 ();
 sg13g2_fill_2 FILLER_47_387 ();
 sg13g2_decap_8 FILLER_47_396 ();
 sg13g2_decap_4 FILLER_47_403 ();
 sg13g2_fill_1 FILLER_47_416 ();
 sg13g2_fill_2 FILLER_47_433 ();
 sg13g2_fill_2 FILLER_47_438 ();
 sg13g2_decap_8 FILLER_47_443 ();
 sg13g2_decap_8 FILLER_47_450 ();
 sg13g2_decap_8 FILLER_47_457 ();
 sg13g2_decap_8 FILLER_47_464 ();
 sg13g2_fill_2 FILLER_47_471 ();
 sg13g2_decap_8 FILLER_47_481 ();
 sg13g2_decap_8 FILLER_47_488 ();
 sg13g2_decap_4 FILLER_47_495 ();
 sg13g2_decap_8 FILLER_47_521 ();
 sg13g2_decap_8 FILLER_47_528 ();
 sg13g2_fill_1 FILLER_47_535 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_fill_1 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_593 ();
 sg13g2_decap_4 FILLER_47_600 ();
 sg13g2_fill_2 FILLER_47_604 ();
 sg13g2_decap_8 FILLER_47_615 ();
 sg13g2_fill_2 FILLER_47_648 ();
 sg13g2_fill_1 FILLER_47_650 ();
 sg13g2_fill_2 FILLER_47_656 ();
 sg13g2_decap_8 FILLER_47_664 ();
 sg13g2_decap_4 FILLER_47_671 ();
 sg13g2_fill_1 FILLER_47_675 ();
 sg13g2_fill_2 FILLER_47_681 ();
 sg13g2_fill_1 FILLER_47_683 ();
 sg13g2_decap_8 FILLER_47_689 ();
 sg13g2_fill_2 FILLER_47_696 ();
 sg13g2_fill_2 FILLER_47_702 ();
 sg13g2_fill_1 FILLER_47_704 ();
 sg13g2_decap_8 FILLER_47_747 ();
 sg13g2_decap_4 FILLER_47_754 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_fill_1 FILLER_47_777 ();
 sg13g2_fill_1 FILLER_47_782 ();
 sg13g2_fill_2 FILLER_47_789 ();
 sg13g2_fill_2 FILLER_47_823 ();
 sg13g2_decap_4 FILLER_47_840 ();
 sg13g2_decap_4 FILLER_47_851 ();
 sg13g2_fill_1 FILLER_47_855 ();
 sg13g2_fill_2 FILLER_47_881 ();
 sg13g2_decap_8 FILLER_47_892 ();
 sg13g2_fill_2 FILLER_47_899 ();
 sg13g2_decap_8 FILLER_47_914 ();
 sg13g2_decap_4 FILLER_47_921 ();
 sg13g2_fill_1 FILLER_47_955 ();
 sg13g2_fill_2 FILLER_47_959 ();
 sg13g2_decap_4 FILLER_47_970 ();
 sg13g2_fill_1 FILLER_47_982 ();
 sg13g2_fill_1 FILLER_47_988 ();
 sg13g2_fill_1 FILLER_47_997 ();
 sg13g2_decap_4 FILLER_47_1012 ();
 sg13g2_decap_4 FILLER_47_1020 ();
 sg13g2_decap_8 FILLER_47_1027 ();
 sg13g2_decap_4 FILLER_47_1034 ();
 sg13g2_fill_2 FILLER_47_1038 ();
 sg13g2_fill_1 FILLER_47_1046 ();
 sg13g2_fill_1 FILLER_47_1051 ();
 sg13g2_fill_1 FILLER_47_1058 ();
 sg13g2_fill_2 FILLER_47_1062 ();
 sg13g2_fill_2 FILLER_47_1069 ();
 sg13g2_fill_1 FILLER_47_1071 ();
 sg13g2_decap_8 FILLER_47_1075 ();
 sg13g2_fill_1 FILLER_47_1088 ();
 sg13g2_fill_2 FILLER_47_1094 ();
 sg13g2_fill_1 FILLER_47_1096 ();
 sg13g2_decap_8 FILLER_47_1112 ();
 sg13g2_fill_1 FILLER_47_1122 ();
 sg13g2_decap_8 FILLER_47_1130 ();
 sg13g2_fill_2 FILLER_47_1137 ();
 sg13g2_decap_8 FILLER_47_1150 ();
 sg13g2_fill_2 FILLER_47_1157 ();
 sg13g2_fill_2 FILLER_47_1174 ();
 sg13g2_fill_1 FILLER_47_1180 ();
 sg13g2_fill_1 FILLER_47_1186 ();
 sg13g2_fill_2 FILLER_47_1218 ();
 sg13g2_fill_2 FILLER_47_1225 ();
 sg13g2_fill_2 FILLER_47_1232 ();
 sg13g2_decap_8 FILLER_47_1259 ();
 sg13g2_decap_8 FILLER_47_1266 ();
 sg13g2_decap_8 FILLER_47_1273 ();
 sg13g2_decap_4 FILLER_47_1280 ();
 sg13g2_fill_2 FILLER_47_1284 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_68 ();
 sg13g2_fill_2 FILLER_48_75 ();
 sg13g2_fill_1 FILLER_48_77 ();
 sg13g2_decap_4 FILLER_48_82 ();
 sg13g2_fill_2 FILLER_48_86 ();
 sg13g2_decap_8 FILLER_48_94 ();
 sg13g2_fill_2 FILLER_48_101 ();
 sg13g2_fill_1 FILLER_48_109 ();
 sg13g2_decap_4 FILLER_48_117 ();
 sg13g2_fill_2 FILLER_48_121 ();
 sg13g2_fill_2 FILLER_48_128 ();
 sg13g2_fill_1 FILLER_48_130 ();
 sg13g2_decap_8 FILLER_48_136 ();
 sg13g2_decap_4 FILLER_48_143 ();
 sg13g2_decap_4 FILLER_48_157 ();
 sg13g2_fill_1 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_170 ();
 sg13g2_decap_4 FILLER_48_177 ();
 sg13g2_fill_2 FILLER_48_194 ();
 sg13g2_fill_2 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_250 ();
 sg13g2_fill_1 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_277 ();
 sg13g2_fill_1 FILLER_48_283 ();
 sg13g2_fill_1 FILLER_48_289 ();
 sg13g2_fill_1 FILLER_48_295 ();
 sg13g2_decap_4 FILLER_48_313 ();
 sg13g2_fill_2 FILLER_48_322 ();
 sg13g2_fill_2 FILLER_48_333 ();
 sg13g2_decap_8 FILLER_48_339 ();
 sg13g2_fill_1 FILLER_48_346 ();
 sg13g2_decap_8 FILLER_48_373 ();
 sg13g2_decap_4 FILLER_48_380 ();
 sg13g2_fill_2 FILLER_48_388 ();
 sg13g2_fill_1 FILLER_48_398 ();
 sg13g2_decap_4 FILLER_48_402 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_fill_2 FILLER_48_420 ();
 sg13g2_fill_1 FILLER_48_433 ();
 sg13g2_fill_1 FILLER_48_456 ();
 sg13g2_fill_1 FILLER_48_462 ();
 sg13g2_fill_1 FILLER_48_466 ();
 sg13g2_fill_2 FILLER_48_472 ();
 sg13g2_decap_8 FILLER_48_479 ();
 sg13g2_fill_1 FILLER_48_497 ();
 sg13g2_fill_2 FILLER_48_503 ();
 sg13g2_fill_1 FILLER_48_505 ();
 sg13g2_fill_2 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_534 ();
 sg13g2_decap_4 FILLER_48_541 ();
 sg13g2_fill_2 FILLER_48_545 ();
 sg13g2_decap_8 FILLER_48_552 ();
 sg13g2_fill_2 FILLER_48_559 ();
 sg13g2_fill_1 FILLER_48_561 ();
 sg13g2_fill_2 FILLER_48_581 ();
 sg13g2_fill_2 FILLER_48_592 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_fill_1 FILLER_48_609 ();
 sg13g2_decap_4 FILLER_48_622 ();
 sg13g2_fill_1 FILLER_48_626 ();
 sg13g2_decap_8 FILLER_48_636 ();
 sg13g2_decap_8 FILLER_48_643 ();
 sg13g2_decap_8 FILLER_48_650 ();
 sg13g2_decap_4 FILLER_48_657 ();
 sg13g2_fill_2 FILLER_48_672 ();
 sg13g2_fill_2 FILLER_48_678 ();
 sg13g2_fill_1 FILLER_48_695 ();
 sg13g2_fill_2 FILLER_48_701 ();
 sg13g2_decap_4 FILLER_48_717 ();
 sg13g2_fill_1 FILLER_48_721 ();
 sg13g2_decap_4 FILLER_48_728 ();
 sg13g2_fill_2 FILLER_48_732 ();
 sg13g2_fill_1 FILLER_48_742 ();
 sg13g2_fill_2 FILLER_48_747 ();
 sg13g2_decap_4 FILLER_48_753 ();
 sg13g2_fill_2 FILLER_48_757 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_fill_2 FILLER_48_786 ();
 sg13g2_fill_2 FILLER_48_804 ();
 sg13g2_fill_1 FILLER_48_806 ();
 sg13g2_fill_2 FILLER_48_810 ();
 sg13g2_fill_1 FILLER_48_812 ();
 sg13g2_fill_1 FILLER_48_819 ();
 sg13g2_fill_2 FILLER_48_823 ();
 sg13g2_decap_8 FILLER_48_829 ();
 sg13g2_decap_8 FILLER_48_836 ();
 sg13g2_fill_2 FILLER_48_850 ();
 sg13g2_decap_4 FILLER_48_859 ();
 sg13g2_fill_2 FILLER_48_867 ();
 sg13g2_fill_1 FILLER_48_869 ();
 sg13g2_fill_2 FILLER_48_877 ();
 sg13g2_fill_1 FILLER_48_879 ();
 sg13g2_decap_8 FILLER_48_899 ();
 sg13g2_decap_4 FILLER_48_906 ();
 sg13g2_decap_4 FILLER_48_920 ();
 sg13g2_fill_1 FILLER_48_928 ();
 sg13g2_fill_2 FILLER_48_944 ();
 sg13g2_fill_2 FILLER_48_951 ();
 sg13g2_decap_8 FILLER_48_956 ();
 sg13g2_decap_8 FILLER_48_963 ();
 sg13g2_fill_2 FILLER_48_970 ();
 sg13g2_fill_1 FILLER_48_972 ();
 sg13g2_fill_1 FILLER_48_982 ();
 sg13g2_decap_8 FILLER_48_992 ();
 sg13g2_fill_1 FILLER_48_999 ();
 sg13g2_fill_2 FILLER_48_1004 ();
 sg13g2_fill_1 FILLER_48_1006 ();
 sg13g2_fill_1 FILLER_48_1012 ();
 sg13g2_fill_2 FILLER_48_1021 ();
 sg13g2_decap_8 FILLER_48_1029 ();
 sg13g2_fill_2 FILLER_48_1036 ();
 sg13g2_fill_2 FILLER_48_1050 ();
 sg13g2_fill_1 FILLER_48_1052 ();
 sg13g2_fill_2 FILLER_48_1057 ();
 sg13g2_fill_1 FILLER_48_1110 ();
 sg13g2_fill_1 FILLER_48_1116 ();
 sg13g2_fill_1 FILLER_48_1123 ();
 sg13g2_fill_1 FILLER_48_1132 ();
 sg13g2_fill_1 FILLER_48_1137 ();
 sg13g2_decap_8 FILLER_48_1146 ();
 sg13g2_decap_8 FILLER_48_1153 ();
 sg13g2_fill_1 FILLER_48_1160 ();
 sg13g2_decap_8 FILLER_48_1168 ();
 sg13g2_fill_1 FILLER_48_1175 ();
 sg13g2_decap_8 FILLER_48_1180 ();
 sg13g2_fill_1 FILLER_48_1187 ();
 sg13g2_decap_8 FILLER_48_1219 ();
 sg13g2_fill_2 FILLER_48_1226 ();
 sg13g2_decap_8 FILLER_48_1233 ();
 sg13g2_decap_8 FILLER_48_1240 ();
 sg13g2_fill_2 FILLER_48_1247 ();
 sg13g2_decap_4 FILLER_48_1257 ();
 sg13g2_decap_4 FILLER_48_1265 ();
 sg13g2_fill_2 FILLER_48_1269 ();
 sg13g2_decap_8 FILLER_48_1305 ();
 sg13g2_fill_2 FILLER_48_1312 ();
 sg13g2_decap_8 FILLER_48_1318 ();
 sg13g2_fill_1 FILLER_48_1325 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_4 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_27 ();
 sg13g2_decap_8 FILLER_49_34 ();
 sg13g2_decap_8 FILLER_49_41 ();
 sg13g2_decap_4 FILLER_49_48 ();
 sg13g2_decap_4 FILLER_49_66 ();
 sg13g2_decap_8 FILLER_49_75 ();
 sg13g2_decap_8 FILLER_49_82 ();
 sg13g2_decap_8 FILLER_49_89 ();
 sg13g2_fill_1 FILLER_49_96 ();
 sg13g2_decap_4 FILLER_49_116 ();
 sg13g2_fill_1 FILLER_49_120 ();
 sg13g2_decap_4 FILLER_49_129 ();
 sg13g2_fill_2 FILLER_49_133 ();
 sg13g2_fill_2 FILLER_49_139 ();
 sg13g2_fill_1 FILLER_49_141 ();
 sg13g2_fill_2 FILLER_49_158 ();
 sg13g2_fill_2 FILLER_49_164 ();
 sg13g2_fill_1 FILLER_49_166 ();
 sg13g2_decap_8 FILLER_49_177 ();
 sg13g2_fill_2 FILLER_49_184 ();
 sg13g2_fill_1 FILLER_49_186 ();
 sg13g2_decap_8 FILLER_49_191 ();
 sg13g2_fill_1 FILLER_49_198 ();
 sg13g2_decap_8 FILLER_49_202 ();
 sg13g2_fill_2 FILLER_49_213 ();
 sg13g2_fill_1 FILLER_49_215 ();
 sg13g2_fill_2 FILLER_49_225 ();
 sg13g2_fill_2 FILLER_49_240 ();
 sg13g2_fill_1 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_253 ();
 sg13g2_decap_8 FILLER_49_260 ();
 sg13g2_fill_1 FILLER_49_267 ();
 sg13g2_fill_2 FILLER_49_271 ();
 sg13g2_fill_1 FILLER_49_273 ();
 sg13g2_fill_2 FILLER_49_281 ();
 sg13g2_fill_2 FILLER_49_296 ();
 sg13g2_fill_1 FILLER_49_316 ();
 sg13g2_decap_4 FILLER_49_353 ();
 sg13g2_fill_1 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_fill_1 FILLER_49_396 ();
 sg13g2_fill_1 FILLER_49_403 ();
 sg13g2_fill_1 FILLER_49_419 ();
 sg13g2_decap_8 FILLER_49_430 ();
 sg13g2_decap_4 FILLER_49_437 ();
 sg13g2_fill_1 FILLER_49_445 ();
 sg13g2_fill_1 FILLER_49_458 ();
 sg13g2_decap_8 FILLER_49_464 ();
 sg13g2_fill_2 FILLER_49_471 ();
 sg13g2_fill_1 FILLER_49_488 ();
 sg13g2_fill_1 FILLER_49_508 ();
 sg13g2_decap_8 FILLER_49_513 ();
 sg13g2_fill_1 FILLER_49_537 ();
 sg13g2_fill_2 FILLER_49_542 ();
 sg13g2_fill_1 FILLER_49_544 ();
 sg13g2_fill_1 FILLER_49_574 ();
 sg13g2_fill_1 FILLER_49_585 ();
 sg13g2_fill_1 FILLER_49_591 ();
 sg13g2_fill_1 FILLER_49_596 ();
 sg13g2_fill_1 FILLER_49_612 ();
 sg13g2_decap_4 FILLER_49_617 ();
 sg13g2_fill_2 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_666 ();
 sg13g2_fill_1 FILLER_49_673 ();
 sg13g2_decap_8 FILLER_49_692 ();
 sg13g2_fill_2 FILLER_49_699 ();
 sg13g2_fill_1 FILLER_49_705 ();
 sg13g2_fill_1 FILLER_49_709 ();
 sg13g2_fill_1 FILLER_49_722 ();
 sg13g2_fill_1 FILLER_49_735 ();
 sg13g2_fill_2 FILLER_49_741 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_fill_2 FILLER_49_756 ();
 sg13g2_fill_1 FILLER_49_758 ();
 sg13g2_decap_8 FILLER_49_776 ();
 sg13g2_decap_4 FILLER_49_783 ();
 sg13g2_fill_1 FILLER_49_798 ();
 sg13g2_decap_4 FILLER_49_804 ();
 sg13g2_fill_1 FILLER_49_808 ();
 sg13g2_decap_8 FILLER_49_816 ();
 sg13g2_fill_1 FILLER_49_823 ();
 sg13g2_fill_1 FILLER_49_837 ();
 sg13g2_decap_4 FILLER_49_853 ();
 sg13g2_fill_1 FILLER_49_864 ();
 sg13g2_fill_2 FILLER_49_874 ();
 sg13g2_fill_1 FILLER_49_880 ();
 sg13g2_decap_8 FILLER_49_890 ();
 sg13g2_decap_4 FILLER_49_897 ();
 sg13g2_fill_2 FILLER_49_901 ();
 sg13g2_decap_8 FILLER_49_908 ();
 sg13g2_fill_2 FILLER_49_915 ();
 sg13g2_fill_1 FILLER_49_917 ();
 sg13g2_fill_2 FILLER_49_924 ();
 sg13g2_fill_1 FILLER_49_926 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_941 ();
 sg13g2_decap_8 FILLER_49_948 ();
 sg13g2_decap_4 FILLER_49_963 ();
 sg13g2_fill_2 FILLER_49_967 ();
 sg13g2_decap_4 FILLER_49_972 ();
 sg13g2_fill_1 FILLER_49_989 ();
 sg13g2_decap_8 FILLER_49_995 ();
 sg13g2_fill_2 FILLER_49_1002 ();
 sg13g2_fill_2 FILLER_49_1017 ();
 sg13g2_fill_1 FILLER_49_1024 ();
 sg13g2_decap_8 FILLER_49_1031 ();
 sg13g2_decap_8 FILLER_49_1038 ();
 sg13g2_decap_4 FILLER_49_1045 ();
 sg13g2_fill_2 FILLER_49_1065 ();
 sg13g2_fill_1 FILLER_49_1067 ();
 sg13g2_fill_2 FILLER_49_1073 ();
 sg13g2_fill_1 FILLER_49_1075 ();
 sg13g2_fill_1 FILLER_49_1079 ();
 sg13g2_decap_8 FILLER_49_1096 ();
 sg13g2_decap_4 FILLER_49_1107 ();
 sg13g2_fill_2 FILLER_49_1116 ();
 sg13g2_fill_1 FILLER_49_1118 ();
 sg13g2_decap_8 FILLER_49_1138 ();
 sg13g2_fill_1 FILLER_49_1145 ();
 sg13g2_fill_1 FILLER_49_1152 ();
 sg13g2_decap_8 FILLER_49_1164 ();
 sg13g2_decap_8 FILLER_49_1171 ();
 sg13g2_fill_1 FILLER_49_1178 ();
 sg13g2_fill_1 FILLER_49_1184 ();
 sg13g2_fill_2 FILLER_49_1195 ();
 sg13g2_decap_8 FILLER_49_1226 ();
 sg13g2_decap_4 FILLER_49_1259 ();
 sg13g2_decap_8 FILLER_49_1271 ();
 sg13g2_decap_8 FILLER_49_1278 ();
 sg13g2_decap_8 FILLER_49_1285 ();
 sg13g2_decap_8 FILLER_49_1292 ();
 sg13g2_decap_4 FILLER_49_1299 ();
 sg13g2_fill_1 FILLER_49_1303 ();
 sg13g2_decap_4 FILLER_49_1308 ();
 sg13g2_fill_1 FILLER_49_1312 ();
 sg13g2_decap_8 FILLER_49_1317 ();
 sg13g2_fill_2 FILLER_49_1324 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_fill_1 FILLER_50_28 ();
 sg13g2_fill_2 FILLER_50_104 ();
 sg13g2_fill_1 FILLER_50_112 ();
 sg13g2_decap_4 FILLER_50_137 ();
 sg13g2_fill_2 FILLER_50_141 ();
 sg13g2_fill_1 FILLER_50_166 ();
 sg13g2_fill_1 FILLER_50_178 ();
 sg13g2_fill_1 FILLER_50_183 ();
 sg13g2_fill_1 FILLER_50_189 ();
 sg13g2_fill_2 FILLER_50_195 ();
 sg13g2_fill_1 FILLER_50_205 ();
 sg13g2_decap_4 FILLER_50_217 ();
 sg13g2_fill_2 FILLER_50_221 ();
 sg13g2_fill_1 FILLER_50_236 ();
 sg13g2_decap_4 FILLER_50_242 ();
 sg13g2_fill_2 FILLER_50_246 ();
 sg13g2_decap_8 FILLER_50_253 ();
 sg13g2_decap_8 FILLER_50_260 ();
 sg13g2_decap_4 FILLER_50_267 ();
 sg13g2_decap_4 FILLER_50_276 ();
 sg13g2_fill_2 FILLER_50_280 ();
 sg13g2_fill_2 FILLER_50_287 ();
 sg13g2_fill_1 FILLER_50_289 ();
 sg13g2_fill_1 FILLER_50_293 ();
 sg13g2_fill_1 FILLER_50_302 ();
 sg13g2_fill_1 FILLER_50_306 ();
 sg13g2_fill_2 FILLER_50_317 ();
 sg13g2_fill_1 FILLER_50_340 ();
 sg13g2_fill_2 FILLER_50_345 ();
 sg13g2_decap_8 FILLER_50_355 ();
 sg13g2_fill_1 FILLER_50_362 ();
 sg13g2_fill_2 FILLER_50_367 ();
 sg13g2_fill_1 FILLER_50_369 ();
 sg13g2_decap_8 FILLER_50_383 ();
 sg13g2_fill_2 FILLER_50_390 ();
 sg13g2_fill_1 FILLER_50_392 ();
 sg13g2_fill_1 FILLER_50_398 ();
 sg13g2_fill_2 FILLER_50_402 ();
 sg13g2_fill_2 FILLER_50_418 ();
 sg13g2_fill_1 FILLER_50_430 ();
 sg13g2_decap_8 FILLER_50_438 ();
 sg13g2_fill_1 FILLER_50_445 ();
 sg13g2_fill_1 FILLER_50_459 ();
 sg13g2_fill_2 FILLER_50_472 ();
 sg13g2_decap_8 FILLER_50_481 ();
 sg13g2_fill_2 FILLER_50_492 ();
 sg13g2_decap_4 FILLER_50_499 ();
 sg13g2_fill_2 FILLER_50_503 ();
 sg13g2_decap_8 FILLER_50_509 ();
 sg13g2_fill_2 FILLER_50_516 ();
 sg13g2_decap_4 FILLER_50_524 ();
 sg13g2_decap_8 FILLER_50_538 ();
 sg13g2_decap_4 FILLER_50_545 ();
 sg13g2_fill_1 FILLER_50_549 ();
 sg13g2_decap_4 FILLER_50_554 ();
 sg13g2_fill_1 FILLER_50_558 ();
 sg13g2_fill_2 FILLER_50_563 ();
 sg13g2_fill_1 FILLER_50_568 ();
 sg13g2_fill_2 FILLER_50_594 ();
 sg13g2_fill_1 FILLER_50_596 ();
 sg13g2_fill_1 FILLER_50_608 ();
 sg13g2_fill_1 FILLER_50_622 ();
 sg13g2_decap_4 FILLER_50_632 ();
 sg13g2_fill_1 FILLER_50_641 ();
 sg13g2_decap_8 FILLER_50_657 ();
 sg13g2_decap_4 FILLER_50_664 ();
 sg13g2_fill_2 FILLER_50_668 ();
 sg13g2_fill_2 FILLER_50_673 ();
 sg13g2_fill_1 FILLER_50_683 ();
 sg13g2_fill_1 FILLER_50_705 ();
 sg13g2_fill_1 FILLER_50_711 ();
 sg13g2_fill_1 FILLER_50_715 ();
 sg13g2_fill_2 FILLER_50_721 ();
 sg13g2_decap_8 FILLER_50_738 ();
 sg13g2_fill_1 FILLER_50_745 ();
 sg13g2_decap_4 FILLER_50_756 ();
 sg13g2_fill_1 FILLER_50_760 ();
 sg13g2_fill_1 FILLER_50_767 ();
 sg13g2_fill_2 FILLER_50_786 ();
 sg13g2_decap_4 FILLER_50_796 ();
 sg13g2_fill_1 FILLER_50_800 ();
 sg13g2_decap_8 FILLER_50_806 ();
 sg13g2_decap_8 FILLER_50_813 ();
 sg13g2_fill_1 FILLER_50_846 ();
 sg13g2_fill_1 FILLER_50_850 ();
 sg13g2_fill_2 FILLER_50_855 ();
 sg13g2_decap_4 FILLER_50_862 ();
 sg13g2_fill_1 FILLER_50_866 ();
 sg13g2_decap_8 FILLER_50_871 ();
 sg13g2_decap_8 FILLER_50_887 ();
 sg13g2_fill_1 FILLER_50_894 ();
 sg13g2_fill_1 FILLER_50_900 ();
 sg13g2_decap_8 FILLER_50_906 ();
 sg13g2_decap_4 FILLER_50_913 ();
 sg13g2_fill_1 FILLER_50_921 ();
 sg13g2_fill_1 FILLER_50_926 ();
 sg13g2_decap_8 FILLER_50_931 ();
 sg13g2_decap_8 FILLER_50_938 ();
 sg13g2_decap_4 FILLER_50_945 ();
 sg13g2_decap_8 FILLER_50_958 ();
 sg13g2_fill_2 FILLER_50_965 ();
 sg13g2_fill_1 FILLER_50_967 ();
 sg13g2_fill_2 FILLER_50_987 ();
 sg13g2_decap_8 FILLER_50_995 ();
 sg13g2_decap_8 FILLER_50_1002 ();
 sg13g2_decap_8 FILLER_50_1009 ();
 sg13g2_decap_8 FILLER_50_1016 ();
 sg13g2_fill_2 FILLER_50_1023 ();
 sg13g2_fill_1 FILLER_50_1025 ();
 sg13g2_decap_4 FILLER_50_1035 ();
 sg13g2_fill_1 FILLER_50_1039 ();
 sg13g2_decap_8 FILLER_50_1052 ();
 sg13g2_decap_4 FILLER_50_1059 ();
 sg13g2_fill_1 FILLER_50_1063 ();
 sg13g2_fill_2 FILLER_50_1070 ();
 sg13g2_decap_8 FILLER_50_1076 ();
 sg13g2_fill_2 FILLER_50_1083 ();
 sg13g2_fill_1 FILLER_50_1090 ();
 sg13g2_fill_2 FILLER_50_1100 ();
 sg13g2_fill_1 FILLER_50_1106 ();
 sg13g2_decap_4 FILLER_50_1112 ();
 sg13g2_fill_1 FILLER_50_1116 ();
 sg13g2_fill_1 FILLER_50_1121 ();
 sg13g2_fill_2 FILLER_50_1127 ();
 sg13g2_fill_2 FILLER_50_1134 ();
 sg13g2_fill_2 FILLER_50_1141 ();
 sg13g2_decap_8 FILLER_50_1148 ();
 sg13g2_fill_1 FILLER_50_1155 ();
 sg13g2_fill_1 FILLER_50_1159 ();
 sg13g2_fill_1 FILLER_50_1164 ();
 sg13g2_fill_2 FILLER_50_1169 ();
 sg13g2_fill_1 FILLER_50_1175 ();
 sg13g2_fill_2 FILLER_50_1195 ();
 sg13g2_fill_1 FILLER_50_1197 ();
 sg13g2_fill_1 FILLER_50_1201 ();
 sg13g2_fill_2 FILLER_50_1224 ();
 sg13g2_fill_2 FILLER_50_1236 ();
 sg13g2_decap_8 FILLER_50_1241 ();
 sg13g2_decap_8 FILLER_50_1252 ();
 sg13g2_fill_2 FILLER_50_1259 ();
 sg13g2_fill_1 FILLER_50_1269 ();
 sg13g2_fill_2 FILLER_50_1275 ();
 sg13g2_fill_1 FILLER_50_1277 ();
 sg13g2_fill_2 FILLER_50_1286 ();
 sg13g2_decap_8 FILLER_50_1301 ();
 sg13g2_fill_1 FILLER_50_1312 ();
 sg13g2_fill_1 FILLER_50_1325 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_36 ();
 sg13g2_decap_4 FILLER_51_43 ();
 sg13g2_fill_1 FILLER_51_47 ();
 sg13g2_decap_8 FILLER_51_78 ();
 sg13g2_fill_1 FILLER_51_85 ();
 sg13g2_fill_2 FILLER_51_112 ();
 sg13g2_fill_2 FILLER_51_118 ();
 sg13g2_fill_1 FILLER_51_120 ();
 sg13g2_fill_1 FILLER_51_125 ();
 sg13g2_fill_1 FILLER_51_132 ();
 sg13g2_fill_1 FILLER_51_137 ();
 sg13g2_fill_1 FILLER_51_172 ();
 sg13g2_fill_1 FILLER_51_182 ();
 sg13g2_fill_1 FILLER_51_229 ();
 sg13g2_fill_1 FILLER_51_238 ();
 sg13g2_decap_4 FILLER_51_252 ();
 sg13g2_fill_1 FILLER_51_256 ();
 sg13g2_decap_4 FILLER_51_264 ();
 sg13g2_fill_2 FILLER_51_268 ();
 sg13g2_fill_2 FILLER_51_284 ();
 sg13g2_decap_8 FILLER_51_291 ();
 sg13g2_fill_2 FILLER_51_298 ();
 sg13g2_fill_1 FILLER_51_300 ();
 sg13g2_fill_1 FILLER_51_313 ();
 sg13g2_fill_1 FILLER_51_323 ();
 sg13g2_fill_2 FILLER_51_328 ();
 sg13g2_fill_2 FILLER_51_334 ();
 sg13g2_decap_8 FILLER_51_345 ();
 sg13g2_decap_4 FILLER_51_352 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_decap_8 FILLER_51_363 ();
 sg13g2_decap_4 FILLER_51_370 ();
 sg13g2_fill_2 FILLER_51_374 ();
 sg13g2_decap_4 FILLER_51_387 ();
 sg13g2_fill_2 FILLER_51_394 ();
 sg13g2_fill_1 FILLER_51_396 ();
 sg13g2_decap_8 FILLER_51_410 ();
 sg13g2_decap_8 FILLER_51_421 ();
 sg13g2_fill_2 FILLER_51_428 ();
 sg13g2_decap_4 FILLER_51_440 ();
 sg13g2_fill_1 FILLER_51_444 ();
 sg13g2_fill_1 FILLER_51_457 ();
 sg13g2_decap_4 FILLER_51_461 ();
 sg13g2_fill_2 FILLER_51_465 ();
 sg13g2_fill_1 FILLER_51_486 ();
 sg13g2_fill_2 FILLER_51_496 ();
 sg13g2_fill_1 FILLER_51_498 ();
 sg13g2_decap_4 FILLER_51_504 ();
 sg13g2_fill_1 FILLER_51_508 ();
 sg13g2_fill_1 FILLER_51_516 ();
 sg13g2_decap_4 FILLER_51_522 ();
 sg13g2_decap_8 FILLER_51_536 ();
 sg13g2_fill_1 FILLER_51_543 ();
 sg13g2_decap_8 FILLER_51_549 ();
 sg13g2_decap_8 FILLER_51_556 ();
 sg13g2_fill_1 FILLER_51_563 ();
 sg13g2_fill_1 FILLER_51_576 ();
 sg13g2_fill_1 FILLER_51_582 ();
 sg13g2_fill_2 FILLER_51_588 ();
 sg13g2_fill_2 FILLER_51_595 ();
 sg13g2_fill_2 FILLER_51_600 ();
 sg13g2_fill_2 FILLER_51_610 ();
 sg13g2_fill_1 FILLER_51_612 ();
 sg13g2_fill_2 FILLER_51_618 ();
 sg13g2_fill_1 FILLER_51_620 ();
 sg13g2_fill_2 FILLER_51_624 ();
 sg13g2_fill_1 FILLER_51_626 ();
 sg13g2_fill_2 FILLER_51_640 ();
 sg13g2_fill_1 FILLER_51_642 ();
 sg13g2_decap_4 FILLER_51_647 ();
 sg13g2_decap_8 FILLER_51_656 ();
 sg13g2_decap_8 FILLER_51_663 ();
 sg13g2_fill_1 FILLER_51_699 ();
 sg13g2_fill_2 FILLER_51_708 ();
 sg13g2_decap_8 FILLER_51_748 ();
 sg13g2_fill_1 FILLER_51_755 ();
 sg13g2_decap_8 FILLER_51_805 ();
 sg13g2_decap_8 FILLER_51_812 ();
 sg13g2_decap_8 FILLER_51_819 ();
 sg13g2_decap_8 FILLER_51_826 ();
 sg13g2_fill_2 FILLER_51_833 ();
 sg13g2_fill_1 FILLER_51_835 ();
 sg13g2_fill_1 FILLER_51_857 ();
 sg13g2_decap_4 FILLER_51_864 ();
 sg13g2_fill_2 FILLER_51_868 ();
 sg13g2_fill_2 FILLER_51_876 ();
 sg13g2_fill_1 FILLER_51_878 ();
 sg13g2_fill_1 FILLER_51_884 ();
 sg13g2_fill_1 FILLER_51_894 ();
 sg13g2_fill_2 FILLER_51_904 ();
 sg13g2_fill_1 FILLER_51_906 ();
 sg13g2_fill_2 FILLER_51_915 ();
 sg13g2_decap_8 FILLER_51_930 ();
 sg13g2_decap_8 FILLER_51_937 ();
 sg13g2_decap_4 FILLER_51_944 ();
 sg13g2_fill_2 FILLER_51_951 ();
 sg13g2_fill_1 FILLER_51_953 ();
 sg13g2_fill_2 FILLER_51_957 ();
 sg13g2_fill_1 FILLER_51_959 ();
 sg13g2_decap_4 FILLER_51_965 ();
 sg13g2_fill_1 FILLER_51_969 ();
 sg13g2_decap_8 FILLER_51_974 ();
 sg13g2_fill_1 FILLER_51_981 ();
 sg13g2_fill_2 FILLER_51_986 ();
 sg13g2_decap_8 FILLER_51_1001 ();
 sg13g2_decap_4 FILLER_51_1008 ();
 sg13g2_fill_2 FILLER_51_1023 ();
 sg13g2_fill_1 FILLER_51_1025 ();
 sg13g2_decap_4 FILLER_51_1057 ();
 sg13g2_fill_1 FILLER_51_1065 ();
 sg13g2_decap_4 FILLER_51_1071 ();
 sg13g2_decap_8 FILLER_51_1078 ();
 sg13g2_fill_2 FILLER_51_1085 ();
 sg13g2_fill_1 FILLER_51_1087 ();
 sg13g2_decap_4 FILLER_51_1095 ();
 sg13g2_fill_1 FILLER_51_1099 ();
 sg13g2_decap_8 FILLER_51_1110 ();
 sg13g2_decap_4 FILLER_51_1117 ();
 sg13g2_fill_1 FILLER_51_1126 ();
 sg13g2_fill_1 FILLER_51_1131 ();
 sg13g2_fill_1 FILLER_51_1139 ();
 sg13g2_decap_4 FILLER_51_1145 ();
 sg13g2_fill_1 FILLER_51_1149 ();
 sg13g2_fill_2 FILLER_51_1158 ();
 sg13g2_fill_1 FILLER_51_1160 ();
 sg13g2_decap_8 FILLER_51_1171 ();
 sg13g2_fill_1 FILLER_51_1178 ();
 sg13g2_decap_8 FILLER_51_1192 ();
 sg13g2_fill_2 FILLER_51_1199 ();
 sg13g2_fill_1 FILLER_51_1201 ();
 sg13g2_fill_2 FILLER_51_1210 ();
 sg13g2_fill_2 FILLER_51_1231 ();
 sg13g2_decap_4 FILLER_51_1267 ();
 sg13g2_fill_2 FILLER_51_1275 ();
 sg13g2_fill_1 FILLER_51_1277 ();
 sg13g2_fill_2 FILLER_51_1291 ();
 sg13g2_decap_8 FILLER_51_1315 ();
 sg13g2_decap_4 FILLER_51_1322 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_14 ();
 sg13g2_fill_2 FILLER_52_41 ();
 sg13g2_fill_2 FILLER_52_56 ();
 sg13g2_fill_1 FILLER_52_58 ();
 sg13g2_decap_4 FILLER_52_102 ();
 sg13g2_decap_8 FILLER_52_122 ();
 sg13g2_decap_8 FILLER_52_143 ();
 sg13g2_decap_8 FILLER_52_150 ();
 sg13g2_fill_2 FILLER_52_177 ();
 sg13g2_fill_2 FILLER_52_200 ();
 sg13g2_fill_1 FILLER_52_219 ();
 sg13g2_fill_1 FILLER_52_243 ();
 sg13g2_fill_2 FILLER_52_256 ();
 sg13g2_decap_4 FILLER_52_272 ();
 sg13g2_fill_1 FILLER_52_276 ();
 sg13g2_decap_4 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_286 ();
 sg13g2_decap_8 FILLER_52_292 ();
 sg13g2_decap_8 FILLER_52_299 ();
 sg13g2_decap_8 FILLER_52_306 ();
 sg13g2_decap_8 FILLER_52_313 ();
 sg13g2_decap_8 FILLER_52_320 ();
 sg13g2_decap_8 FILLER_52_327 ();
 sg13g2_decap_4 FILLER_52_342 ();
 sg13g2_fill_2 FILLER_52_346 ();
 sg13g2_decap_4 FILLER_52_354 ();
 sg13g2_decap_8 FILLER_52_367 ();
 sg13g2_decap_8 FILLER_52_374 ();
 sg13g2_decap_8 FILLER_52_381 ();
 sg13g2_decap_4 FILLER_52_388 ();
 sg13g2_fill_2 FILLER_52_392 ();
 sg13g2_fill_2 FILLER_52_411 ();
 sg13g2_fill_1 FILLER_52_413 ();
 sg13g2_fill_1 FILLER_52_423 ();
 sg13g2_fill_2 FILLER_52_429 ();
 sg13g2_fill_1 FILLER_52_440 ();
 sg13g2_fill_1 FILLER_52_455 ();
 sg13g2_fill_1 FILLER_52_465 ();
 sg13g2_fill_1 FILLER_52_473 ();
 sg13g2_decap_8 FILLER_52_477 ();
 sg13g2_fill_1 FILLER_52_484 ();
 sg13g2_decap_8 FILLER_52_490 ();
 sg13g2_decap_8 FILLER_52_497 ();
 sg13g2_decap_8 FILLER_52_504 ();
 sg13g2_decap_4 FILLER_52_511 ();
 sg13g2_decap_4 FILLER_52_560 ();
 sg13g2_fill_2 FILLER_52_575 ();
 sg13g2_fill_1 FILLER_52_577 ();
 sg13g2_fill_2 FILLER_52_583 ();
 sg13g2_decap_8 FILLER_52_591 ();
 sg13g2_decap_4 FILLER_52_605 ();
 sg13g2_fill_1 FILLER_52_619 ();
 sg13g2_fill_2 FILLER_52_625 ();
 sg13g2_decap_4 FILLER_52_632 ();
 sg13g2_decap_8 FILLER_52_651 ();
 sg13g2_fill_2 FILLER_52_658 ();
 sg13g2_fill_1 FILLER_52_660 ();
 sg13g2_decap_4 FILLER_52_665 ();
 sg13g2_fill_1 FILLER_52_669 ();
 sg13g2_decap_4 FILLER_52_674 ();
 sg13g2_fill_2 FILLER_52_685 ();
 sg13g2_fill_2 FILLER_52_695 ();
 sg13g2_fill_1 FILLER_52_697 ();
 sg13g2_fill_2 FILLER_52_705 ();
 sg13g2_fill_2 FILLER_52_724 ();
 sg13g2_fill_2 FILLER_52_734 ();
 sg13g2_fill_2 FILLER_52_755 ();
 sg13g2_fill_1 FILLER_52_757 ();
 sg13g2_decap_4 FILLER_52_768 ();
 sg13g2_decap_4 FILLER_52_784 ();
 sg13g2_fill_1 FILLER_52_793 ();
 sg13g2_fill_1 FILLER_52_797 ();
 sg13g2_fill_1 FILLER_52_801 ();
 sg13g2_fill_2 FILLER_52_808 ();
 sg13g2_fill_1 FILLER_52_810 ();
 sg13g2_fill_2 FILLER_52_820 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_fill_1 FILLER_52_833 ();
 sg13g2_fill_2 FILLER_52_842 ();
 sg13g2_decap_4 FILLER_52_849 ();
 sg13g2_decap_8 FILLER_52_898 ();
 sg13g2_decap_8 FILLER_52_905 ();
 sg13g2_decap_4 FILLER_52_912 ();
 sg13g2_fill_2 FILLER_52_916 ();
 sg13g2_decap_4 FILLER_52_926 ();
 sg13g2_fill_1 FILLER_52_930 ();
 sg13g2_fill_2 FILLER_52_959 ();
 sg13g2_decap_4 FILLER_52_966 ();
 sg13g2_fill_2 FILLER_52_970 ();
 sg13g2_decap_4 FILLER_52_976 ();
 sg13g2_fill_2 FILLER_52_980 ();
 sg13g2_decap_8 FILLER_52_991 ();
 sg13g2_fill_2 FILLER_52_998 ();
 sg13g2_fill_1 FILLER_52_1026 ();
 sg13g2_decap_8 FILLER_52_1030 ();
 sg13g2_decap_8 FILLER_52_1037 ();
 sg13g2_decap_8 FILLER_52_1044 ();
 sg13g2_decap_8 FILLER_52_1051 ();
 sg13g2_fill_1 FILLER_52_1058 ();
 sg13g2_fill_1 FILLER_52_1062 ();
 sg13g2_fill_1 FILLER_52_1068 ();
 sg13g2_fill_1 FILLER_52_1075 ();
 sg13g2_decap_8 FILLER_52_1080 ();
 sg13g2_fill_2 FILLER_52_1087 ();
 sg13g2_decap_8 FILLER_52_1092 ();
 sg13g2_fill_2 FILLER_52_1099 ();
 sg13g2_fill_1 FILLER_52_1132 ();
 sg13g2_decap_8 FILLER_52_1142 ();
 sg13g2_fill_1 FILLER_52_1149 ();
 sg13g2_fill_1 FILLER_52_1178 ();
 sg13g2_fill_2 FILLER_52_1184 ();
 sg13g2_fill_2 FILLER_52_1190 ();
 sg13g2_fill_1 FILLER_52_1198 ();
 sg13g2_fill_2 FILLER_52_1212 ();
 sg13g2_fill_1 FILLER_52_1220 ();
 sg13g2_fill_1 FILLER_52_1234 ();
 sg13g2_fill_1 FILLER_52_1249 ();
 sg13g2_decap_4 FILLER_52_1254 ();
 sg13g2_fill_2 FILLER_52_1262 ();
 sg13g2_fill_1 FILLER_52_1264 ();
 sg13g2_fill_1 FILLER_52_1271 ();
 sg13g2_decap_8 FILLER_52_1285 ();
 sg13g2_decap_4 FILLER_52_1292 ();
 sg13g2_fill_1 FILLER_52_1296 ();
 sg13g2_fill_2 FILLER_52_1302 ();
 sg13g2_fill_1 FILLER_52_1304 ();
 sg13g2_fill_1 FILLER_52_1325 ();
 sg13g2_decap_8 FILLER_53_26 ();
 sg13g2_decap_8 FILLER_53_33 ();
 sg13g2_decap_8 FILLER_53_53 ();
 sg13g2_decap_8 FILLER_53_60 ();
 sg13g2_decap_8 FILLER_53_67 ();
 sg13g2_decap_8 FILLER_53_74 ();
 sg13g2_decap_8 FILLER_53_81 ();
 sg13g2_decap_8 FILLER_53_88 ();
 sg13g2_fill_2 FILLER_53_95 ();
 sg13g2_fill_1 FILLER_53_97 ();
 sg13g2_decap_8 FILLER_53_115 ();
 sg13g2_decap_4 FILLER_53_122 ();
 sg13g2_fill_1 FILLER_53_143 ();
 sg13g2_fill_2 FILLER_53_148 ();
 sg13g2_fill_1 FILLER_53_154 ();
 sg13g2_fill_2 FILLER_53_174 ();
 sg13g2_fill_2 FILLER_53_192 ();
 sg13g2_fill_1 FILLER_53_201 ();
 sg13g2_fill_2 FILLER_53_224 ();
 sg13g2_fill_1 FILLER_53_226 ();
 sg13g2_decap_8 FILLER_53_268 ();
 sg13g2_decap_8 FILLER_53_275 ();
 sg13g2_fill_2 FILLER_53_282 ();
 sg13g2_fill_1 FILLER_53_284 ();
 sg13g2_fill_1 FILLER_53_296 ();
 sg13g2_fill_2 FILLER_53_304 ();
 sg13g2_fill_1 FILLER_53_306 ();
 sg13g2_fill_2 FILLER_53_339 ();
 sg13g2_decap_8 FILLER_53_348 ();
 sg13g2_fill_2 FILLER_53_355 ();
 sg13g2_fill_1 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_362 ();
 sg13g2_decap_8 FILLER_53_369 ();
 sg13g2_decap_8 FILLER_53_376 ();
 sg13g2_decap_8 FILLER_53_383 ();
 sg13g2_decap_8 FILLER_53_390 ();
 sg13g2_decap_8 FILLER_53_407 ();
 sg13g2_decap_4 FILLER_53_431 ();
 sg13g2_fill_1 FILLER_53_435 ();
 sg13g2_fill_2 FILLER_53_445 ();
 sg13g2_fill_1 FILLER_53_447 ();
 sg13g2_fill_2 FILLER_53_463 ();
 sg13g2_fill_1 FILLER_53_474 ();
 sg13g2_fill_1 FILLER_53_483 ();
 sg13g2_fill_1 FILLER_53_497 ();
 sg13g2_fill_1 FILLER_53_501 ();
 sg13g2_fill_2 FILLER_53_532 ();
 sg13g2_decap_8 FILLER_53_544 ();
 sg13g2_decap_8 FILLER_53_551 ();
 sg13g2_decap_4 FILLER_53_558 ();
 sg13g2_decap_8 FILLER_53_571 ();
 sg13g2_decap_8 FILLER_53_578 ();
 sg13g2_fill_1 FILLER_53_588 ();
 sg13g2_fill_2 FILLER_53_594 ();
 sg13g2_decap_4 FILLER_53_607 ();
 sg13g2_fill_2 FILLER_53_611 ();
 sg13g2_decap_4 FILLER_53_635 ();
 sg13g2_fill_2 FILLER_53_643 ();
 sg13g2_decap_8 FILLER_53_650 ();
 sg13g2_decap_8 FILLER_53_657 ();
 sg13g2_decap_8 FILLER_53_664 ();
 sg13g2_decap_4 FILLER_53_680 ();
 sg13g2_decap_4 FILLER_53_690 ();
 sg13g2_fill_1 FILLER_53_694 ();
 sg13g2_fill_1 FILLER_53_762 ();
 sg13g2_fill_1 FILLER_53_767 ();
 sg13g2_decap_8 FILLER_53_773 ();
 sg13g2_fill_1 FILLER_53_780 ();
 sg13g2_fill_2 FILLER_53_798 ();
 sg13g2_fill_1 FILLER_53_800 ();
 sg13g2_decap_8 FILLER_53_804 ();
 sg13g2_decap_8 FILLER_53_811 ();
 sg13g2_fill_1 FILLER_53_818 ();
 sg13g2_fill_2 FILLER_53_825 ();
 sg13g2_fill_1 FILLER_53_832 ();
 sg13g2_fill_1 FILLER_53_866 ();
 sg13g2_fill_1 FILLER_53_874 ();
 sg13g2_decap_4 FILLER_53_911 ();
 sg13g2_fill_2 FILLER_53_915 ();
 sg13g2_fill_1 FILLER_53_939 ();
 sg13g2_fill_2 FILLER_53_944 ();
 sg13g2_fill_1 FILLER_53_946 ();
 sg13g2_decap_8 FILLER_53_968 ();
 sg13g2_fill_1 FILLER_53_975 ();
 sg13g2_decap_8 FILLER_53_994 ();
 sg13g2_fill_2 FILLER_53_1001 ();
 sg13g2_fill_2 FILLER_53_1011 ();
 sg13g2_fill_1 FILLER_53_1013 ();
 sg13g2_decap_8 FILLER_53_1026 ();
 sg13g2_fill_1 FILLER_53_1048 ();
 sg13g2_fill_1 FILLER_53_1054 ();
 sg13g2_fill_1 FILLER_53_1073 ();
 sg13g2_fill_2 FILLER_53_1090 ();
 sg13g2_decap_4 FILLER_53_1101 ();
 sg13g2_fill_1 FILLER_53_1114 ();
 sg13g2_fill_1 FILLER_53_1120 ();
 sg13g2_fill_1 FILLER_53_1124 ();
 sg13g2_fill_2 FILLER_53_1130 ();
 sg13g2_fill_1 FILLER_53_1132 ();
 sg13g2_decap_8 FILLER_53_1138 ();
 sg13g2_fill_2 FILLER_53_1145 ();
 sg13g2_fill_1 FILLER_53_1147 ();
 sg13g2_decap_8 FILLER_53_1151 ();
 sg13g2_decap_8 FILLER_53_1158 ();
 sg13g2_decap_4 FILLER_53_1165 ();
 sg13g2_fill_2 FILLER_53_1169 ();
 sg13g2_decap_8 FILLER_53_1179 ();
 sg13g2_fill_2 FILLER_53_1186 ();
 sg13g2_fill_2 FILLER_53_1212 ();
 sg13g2_decap_8 FILLER_53_1241 ();
 sg13g2_decap_4 FILLER_53_1248 ();
 sg13g2_fill_1 FILLER_53_1252 ();
 sg13g2_decap_8 FILLER_53_1257 ();
 sg13g2_fill_2 FILLER_53_1264 ();
 sg13g2_fill_1 FILLER_53_1266 ();
 sg13g2_decap_8 FILLER_53_1276 ();
 sg13g2_decap_8 FILLER_53_1283 ();
 sg13g2_decap_4 FILLER_53_1290 ();
 sg13g2_fill_1 FILLER_53_1303 ();
 sg13g2_decap_4 FILLER_53_1309 ();
 sg13g2_decap_8 FILLER_53_1316 ();
 sg13g2_fill_2 FILLER_53_1323 ();
 sg13g2_fill_1 FILLER_53_1325 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_fill_2 FILLER_54_21 ();
 sg13g2_fill_2 FILLER_54_53 ();
 sg13g2_decap_8 FILLER_54_60 ();
 sg13g2_decap_8 FILLER_54_67 ();
 sg13g2_decap_8 FILLER_54_74 ();
 sg13g2_decap_8 FILLER_54_81 ();
 sg13g2_decap_4 FILLER_54_88 ();
 sg13g2_decap_8 FILLER_54_108 ();
 sg13g2_decap_8 FILLER_54_115 ();
 sg13g2_fill_2 FILLER_54_122 ();
 sg13g2_decap_8 FILLER_54_128 ();
 sg13g2_fill_2 FILLER_54_135 ();
 sg13g2_fill_1 FILLER_54_168 ();
 sg13g2_fill_2 FILLER_54_185 ();
 sg13g2_fill_2 FILLER_54_207 ();
 sg13g2_decap_4 FILLER_54_230 ();
 sg13g2_fill_2 FILLER_54_234 ();
 sg13g2_decap_8 FILLER_54_240 ();
 sg13g2_decap_8 FILLER_54_247 ();
 sg13g2_decap_8 FILLER_54_254 ();
 sg13g2_decap_8 FILLER_54_261 ();
 sg13g2_decap_8 FILLER_54_268 ();
 sg13g2_fill_2 FILLER_54_275 ();
 sg13g2_fill_2 FILLER_54_281 ();
 sg13g2_fill_1 FILLER_54_288 ();
 sg13g2_fill_1 FILLER_54_294 ();
 sg13g2_fill_1 FILLER_54_300 ();
 sg13g2_decap_4 FILLER_54_306 ();
 sg13g2_decap_4 FILLER_54_314 ();
 sg13g2_fill_2 FILLER_54_318 ();
 sg13g2_fill_2 FILLER_54_323 ();
 sg13g2_fill_1 FILLER_54_325 ();
 sg13g2_fill_1 FILLER_54_330 ();
 sg13g2_fill_2 FILLER_54_348 ();
 sg13g2_fill_1 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_358 ();
 sg13g2_decap_8 FILLER_54_365 ();
 sg13g2_fill_2 FILLER_54_372 ();
 sg13g2_decap_8 FILLER_54_382 ();
 sg13g2_fill_2 FILLER_54_389 ();
 sg13g2_fill_1 FILLER_54_391 ();
 sg13g2_decap_8 FILLER_54_402 ();
 sg13g2_fill_2 FILLER_54_409 ();
 sg13g2_fill_1 FILLER_54_411 ();
 sg13g2_decap_8 FILLER_54_416 ();
 sg13g2_fill_2 FILLER_54_423 ();
 sg13g2_decap_8 FILLER_54_428 ();
 sg13g2_decap_4 FILLER_54_435 ();
 sg13g2_fill_1 FILLER_54_439 ();
 sg13g2_fill_1 FILLER_54_444 ();
 sg13g2_fill_1 FILLER_54_453 ();
 sg13g2_fill_1 FILLER_54_458 ();
 sg13g2_fill_1 FILLER_54_465 ();
 sg13g2_fill_1 FILLER_54_470 ();
 sg13g2_fill_1 FILLER_54_476 ();
 sg13g2_fill_1 FILLER_54_482 ();
 sg13g2_decap_8 FILLER_54_488 ();
 sg13g2_decap_4 FILLER_54_495 ();
 sg13g2_fill_2 FILLER_54_502 ();
 sg13g2_fill_1 FILLER_54_504 ();
 sg13g2_decap_4 FILLER_54_510 ();
 sg13g2_decap_8 FILLER_54_517 ();
 sg13g2_decap_4 FILLER_54_524 ();
 sg13g2_fill_1 FILLER_54_528 ();
 sg13g2_fill_2 FILLER_54_533 ();
 sg13g2_fill_2 FILLER_54_538 ();
 sg13g2_fill_1 FILLER_54_540 ();
 sg13g2_fill_2 FILLER_54_554 ();
 sg13g2_fill_1 FILLER_54_556 ();
 sg13g2_fill_2 FILLER_54_562 ();
 sg13g2_fill_1 FILLER_54_564 ();
 sg13g2_decap_4 FILLER_54_570 ();
 sg13g2_fill_2 FILLER_54_574 ();
 sg13g2_fill_2 FILLER_54_607 ();
 sg13g2_fill_1 FILLER_54_613 ();
 sg13g2_fill_2 FILLER_54_622 ();
 sg13g2_decap_4 FILLER_54_629 ();
 sg13g2_fill_2 FILLER_54_633 ();
 sg13g2_decap_8 FILLER_54_668 ();
 sg13g2_decap_4 FILLER_54_675 ();
 sg13g2_fill_2 FILLER_54_679 ();
 sg13g2_fill_1 FILLER_54_703 ();
 sg13g2_fill_2 FILLER_54_708 ();
 sg13g2_fill_1 FILLER_54_753 ();
 sg13g2_fill_2 FILLER_54_759 ();
 sg13g2_fill_2 FILLER_54_775 ();
 sg13g2_fill_1 FILLER_54_777 ();
 sg13g2_fill_1 FILLER_54_783 ();
 sg13g2_decap_8 FILLER_54_808 ();
 sg13g2_decap_4 FILLER_54_815 ();
 sg13g2_fill_1 FILLER_54_819 ();
 sg13g2_decap_4 FILLER_54_824 ();
 sg13g2_fill_2 FILLER_54_828 ();
 sg13g2_decap_8 FILLER_54_833 ();
 sg13g2_decap_8 FILLER_54_840 ();
 sg13g2_fill_2 FILLER_54_847 ();
 sg13g2_fill_1 FILLER_54_854 ();
 sg13g2_decap_4 FILLER_54_860 ();
 sg13g2_fill_2 FILLER_54_871 ();
 sg13g2_fill_1 FILLER_54_886 ();
 sg13g2_fill_2 FILLER_54_892 ();
 sg13g2_fill_2 FILLER_54_898 ();
 sg13g2_fill_2 FILLER_54_905 ();
 sg13g2_fill_1 FILLER_54_907 ();
 sg13g2_decap_8 FILLER_54_916 ();
 sg13g2_decap_4 FILLER_54_923 ();
 sg13g2_fill_1 FILLER_54_930 ();
 sg13g2_fill_1 FILLER_54_935 ();
 sg13g2_fill_1 FILLER_54_939 ();
 sg13g2_decap_4 FILLER_54_943 ();
 sg13g2_fill_1 FILLER_54_947 ();
 sg13g2_fill_2 FILLER_54_953 ();
 sg13g2_decap_4 FILLER_54_965 ();
 sg13g2_fill_2 FILLER_54_981 ();
 sg13g2_fill_1 FILLER_54_983 ();
 sg13g2_fill_1 FILLER_54_996 ();
 sg13g2_fill_1 FILLER_54_1002 ();
 sg13g2_fill_2 FILLER_54_1036 ();
 sg13g2_decap_8 FILLER_54_1043 ();
 sg13g2_fill_2 FILLER_54_1050 ();
 sg13g2_fill_1 FILLER_54_1052 ();
 sg13g2_fill_1 FILLER_54_1064 ();
 sg13g2_fill_2 FILLER_54_1071 ();
 sg13g2_decap_8 FILLER_54_1077 ();
 sg13g2_decap_8 FILLER_54_1084 ();
 sg13g2_decap_4 FILLER_54_1091 ();
 sg13g2_fill_2 FILLER_54_1100 ();
 sg13g2_fill_1 FILLER_54_1102 ();
 sg13g2_fill_1 FILLER_54_1115 ();
 sg13g2_fill_1 FILLER_54_1120 ();
 sg13g2_fill_1 FILLER_54_1129 ();
 sg13g2_fill_1 FILLER_54_1134 ();
 sg13g2_decap_4 FILLER_54_1138 ();
 sg13g2_fill_1 FILLER_54_1142 ();
 sg13g2_decap_8 FILLER_54_1160 ();
 sg13g2_decap_8 FILLER_54_1167 ();
 sg13g2_decap_8 FILLER_54_1174 ();
 sg13g2_decap_8 FILLER_54_1181 ();
 sg13g2_fill_1 FILLER_54_1188 ();
 sg13g2_fill_2 FILLER_54_1193 ();
 sg13g2_decap_4 FILLER_54_1199 ();
 sg13g2_fill_2 FILLER_54_1203 ();
 sg13g2_fill_1 FILLER_54_1223 ();
 sg13g2_fill_1 FILLER_54_1234 ();
 sg13g2_fill_2 FILLER_54_1244 ();
 sg13g2_decap_4 FILLER_54_1251 ();
 sg13g2_fill_2 FILLER_54_1259 ();
 sg13g2_fill_1 FILLER_54_1261 ();
 sg13g2_decap_8 FILLER_54_1276 ();
 sg13g2_decap_4 FILLER_54_1283 ();
 sg13g2_fill_2 FILLER_54_1287 ();
 sg13g2_fill_2 FILLER_54_1298 ();
 sg13g2_fill_2 FILLER_54_1308 ();
 sg13g2_fill_1 FILLER_54_1310 ();
 sg13g2_decap_8 FILLER_54_1316 ();
 sg13g2_fill_2 FILLER_54_1323 ();
 sg13g2_fill_1 FILLER_54_1325 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_4 FILLER_55_21 ();
 sg13g2_fill_1 FILLER_55_25 ();
 sg13g2_fill_2 FILLER_55_31 ();
 sg13g2_decap_8 FILLER_55_47 ();
 sg13g2_decap_4 FILLER_55_54 ();
 sg13g2_fill_2 FILLER_55_58 ();
 sg13g2_decap_8 FILLER_55_103 ();
 sg13g2_decap_8 FILLER_55_110 ();
 sg13g2_fill_2 FILLER_55_117 ();
 sg13g2_decap_8 FILLER_55_132 ();
 sg13g2_decap_4 FILLER_55_139 ();
 sg13g2_fill_1 FILLER_55_143 ();
 sg13g2_fill_1 FILLER_55_200 ();
 sg13g2_fill_1 FILLER_55_206 ();
 sg13g2_decap_8 FILLER_55_251 ();
 sg13g2_fill_2 FILLER_55_273 ();
 sg13g2_fill_1 FILLER_55_275 ();
 sg13g2_fill_2 FILLER_55_281 ();
 sg13g2_fill_1 FILLER_55_283 ();
 sg13g2_decap_4 FILLER_55_306 ();
 sg13g2_fill_2 FILLER_55_310 ();
 sg13g2_decap_4 FILLER_55_316 ();
 sg13g2_fill_2 FILLER_55_326 ();
 sg13g2_fill_1 FILLER_55_337 ();
 sg13g2_fill_2 FILLER_55_364 ();
 sg13g2_fill_2 FILLER_55_372 ();
 sg13g2_fill_1 FILLER_55_374 ();
 sg13g2_fill_1 FILLER_55_382 ();
 sg13g2_decap_8 FILLER_55_387 ();
 sg13g2_fill_1 FILLER_55_394 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_fill_1 FILLER_55_409 ();
 sg13g2_fill_2 FILLER_55_418 ();
 sg13g2_fill_2 FILLER_55_424 ();
 sg13g2_fill_1 FILLER_55_440 ();
 sg13g2_decap_8 FILLER_55_447 ();
 sg13g2_decap_8 FILLER_55_454 ();
 sg13g2_fill_2 FILLER_55_461 ();
 sg13g2_fill_1 FILLER_55_463 ();
 sg13g2_decap_4 FILLER_55_478 ();
 sg13g2_decap_8 FILLER_55_486 ();
 sg13g2_decap_8 FILLER_55_493 ();
 sg13g2_decap_4 FILLER_55_500 ();
 sg13g2_fill_1 FILLER_55_508 ();
 sg13g2_fill_1 FILLER_55_513 ();
 sg13g2_decap_8 FILLER_55_540 ();
 sg13g2_decap_4 FILLER_55_547 ();
 sg13g2_fill_1 FILLER_55_571 ();
 sg13g2_fill_2 FILLER_55_577 ();
 sg13g2_decap_8 FILLER_55_614 ();
 sg13g2_decap_8 FILLER_55_630 ();
 sg13g2_fill_2 FILLER_55_637 ();
 sg13g2_decap_8 FILLER_55_660 ();
 sg13g2_decap_4 FILLER_55_667 ();
 sg13g2_decap_4 FILLER_55_680 ();
 sg13g2_fill_2 FILLER_55_692 ();
 sg13g2_fill_2 FILLER_55_698 ();
 sg13g2_fill_1 FILLER_55_700 ();
 sg13g2_fill_1 FILLER_55_706 ();
 sg13g2_fill_2 FILLER_55_711 ();
 sg13g2_fill_2 FILLER_55_720 ();
 sg13g2_fill_1 FILLER_55_725 ();
 sg13g2_decap_8 FILLER_55_761 ();
 sg13g2_fill_2 FILLER_55_768 ();
 sg13g2_fill_1 FILLER_55_770 ();
 sg13g2_decap_4 FILLER_55_787 ();
 sg13g2_fill_2 FILLER_55_796 ();
 sg13g2_decap_8 FILLER_55_815 ();
 sg13g2_fill_2 FILLER_55_822 ();
 sg13g2_fill_1 FILLER_55_824 ();
 sg13g2_fill_2 FILLER_55_845 ();
 sg13g2_fill_1 FILLER_55_851 ();
 sg13g2_fill_1 FILLER_55_855 ();
 sg13g2_fill_1 FILLER_55_860 ();
 sg13g2_fill_1 FILLER_55_868 ();
 sg13g2_fill_2 FILLER_55_881 ();
 sg13g2_fill_2 FILLER_55_887 ();
 sg13g2_decap_8 FILLER_55_895 ();
 sg13g2_decap_8 FILLER_55_902 ();
 sg13g2_fill_1 FILLER_55_915 ();
 sg13g2_fill_2 FILLER_55_958 ();
 sg13g2_fill_1 FILLER_55_960 ();
 sg13g2_decap_8 FILLER_55_965 ();
 sg13g2_decap_4 FILLER_55_972 ();
 sg13g2_fill_2 FILLER_55_981 ();
 sg13g2_fill_1 FILLER_55_983 ();
 sg13g2_fill_2 FILLER_55_996 ();
 sg13g2_fill_1 FILLER_55_998 ();
 sg13g2_decap_8 FILLER_55_1003 ();
 sg13g2_decap_4 FILLER_55_1010 ();
 sg13g2_fill_2 FILLER_55_1018 ();
 sg13g2_fill_1 FILLER_55_1024 ();
 sg13g2_fill_2 FILLER_55_1029 ();
 sg13g2_fill_1 FILLER_55_1036 ();
 sg13g2_decap_8 FILLER_55_1043 ();
 sg13g2_fill_1 FILLER_55_1069 ();
 sg13g2_decap_8 FILLER_55_1075 ();
 sg13g2_fill_2 FILLER_55_1082 ();
 sg13g2_fill_1 FILLER_55_1084 ();
 sg13g2_fill_1 FILLER_55_1096 ();
 sg13g2_decap_4 FILLER_55_1103 ();
 sg13g2_fill_2 FILLER_55_1110 ();
 sg13g2_fill_1 FILLER_55_1112 ();
 sg13g2_decap_8 FILLER_55_1121 ();
 sg13g2_fill_1 FILLER_55_1128 ();
 sg13g2_decap_8 FILLER_55_1137 ();
 sg13g2_fill_2 FILLER_55_1144 ();
 sg13g2_fill_1 FILLER_55_1146 ();
 sg13g2_decap_4 FILLER_55_1152 ();
 sg13g2_fill_1 FILLER_55_1161 ();
 sg13g2_fill_2 FILLER_55_1167 ();
 sg13g2_fill_2 FILLER_55_1172 ();
 sg13g2_fill_2 FILLER_55_1180 ();
 sg13g2_fill_2 FILLER_55_1186 ();
 sg13g2_fill_1 FILLER_55_1188 ();
 sg13g2_fill_2 FILLER_55_1194 ();
 sg13g2_fill_1 FILLER_55_1196 ();
 sg13g2_fill_2 FILLER_55_1202 ();
 sg13g2_fill_2 FILLER_55_1212 ();
 sg13g2_decap_8 FILLER_55_1258 ();
 sg13g2_decap_4 FILLER_55_1265 ();
 sg13g2_decap_8 FILLER_55_1277 ();
 sg13g2_fill_2 FILLER_55_1284 ();
 sg13g2_fill_1 FILLER_55_1290 ();
 sg13g2_decap_4 FILLER_55_1295 ();
 sg13g2_fill_2 FILLER_55_1299 ();
 sg13g2_decap_8 FILLER_55_1305 ();
 sg13g2_decap_8 FILLER_55_1312 ();
 sg13g2_decap_8 FILLER_55_1319 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_4 FILLER_56_44 ();
 sg13g2_fill_1 FILLER_56_48 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_fill_1 FILLER_56_80 ();
 sg13g2_fill_2 FILLER_56_169 ();
 sg13g2_fill_2 FILLER_56_185 ();
 sg13g2_fill_2 FILLER_56_219 ();
 sg13g2_decap_8 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_238 ();
 sg13g2_fill_2 FILLER_56_245 ();
 sg13g2_fill_2 FILLER_56_258 ();
 sg13g2_fill_2 FILLER_56_274 ();
 sg13g2_fill_1 FILLER_56_276 ();
 sg13g2_fill_1 FILLER_56_282 ();
 sg13g2_fill_1 FILLER_56_289 ();
 sg13g2_fill_1 FILLER_56_295 ();
 sg13g2_fill_1 FILLER_56_300 ();
 sg13g2_fill_1 FILLER_56_307 ();
 sg13g2_fill_1 FILLER_56_313 ();
 sg13g2_decap_8 FILLER_56_318 ();
 sg13g2_fill_1 FILLER_56_325 ();
 sg13g2_fill_2 FILLER_56_344 ();
 sg13g2_fill_1 FILLER_56_346 ();
 sg13g2_fill_1 FILLER_56_352 ();
 sg13g2_decap_8 FILLER_56_371 ();
 sg13g2_decap_8 FILLER_56_385 ();
 sg13g2_decap_8 FILLER_56_395 ();
 sg13g2_fill_1 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_411 ();
 sg13g2_decap_8 FILLER_56_418 ();
 sg13g2_decap_4 FILLER_56_437 ();
 sg13g2_decap_4 FILLER_56_445 ();
 sg13g2_decap_4 FILLER_56_459 ();
 sg13g2_fill_1 FILLER_56_463 ();
 sg13g2_fill_2 FILLER_56_469 ();
 sg13g2_fill_1 FILLER_56_471 ();
 sg13g2_decap_8 FILLER_56_476 ();
 sg13g2_fill_1 FILLER_56_483 ();
 sg13g2_fill_2 FILLER_56_500 ();
 sg13g2_fill_2 FILLER_56_518 ();
 sg13g2_fill_1 FILLER_56_520 ();
 sg13g2_fill_1 FILLER_56_525 ();
 sg13g2_decap_8 FILLER_56_534 ();
 sg13g2_decap_8 FILLER_56_541 ();
 sg13g2_decap_4 FILLER_56_548 ();
 sg13g2_fill_2 FILLER_56_566 ();
 sg13g2_fill_1 FILLER_56_574 ();
 sg13g2_fill_2 FILLER_56_585 ();
 sg13g2_fill_1 FILLER_56_595 ();
 sg13g2_fill_1 FILLER_56_605 ();
 sg13g2_fill_2 FILLER_56_654 ();
 sg13g2_fill_1 FILLER_56_662 ();
 sg13g2_decap_8 FILLER_56_666 ();
 sg13g2_fill_2 FILLER_56_673 ();
 sg13g2_fill_1 FILLER_56_675 ();
 sg13g2_decap_4 FILLER_56_679 ();
 sg13g2_fill_2 FILLER_56_687 ();
 sg13g2_fill_1 FILLER_56_718 ();
 sg13g2_fill_1 FILLER_56_737 ();
 sg13g2_decap_8 FILLER_56_784 ();
 sg13g2_decap_8 FILLER_56_791 ();
 sg13g2_fill_2 FILLER_56_798 ();
 sg13g2_fill_1 FILLER_56_800 ();
 sg13g2_fill_1 FILLER_56_804 ();
 sg13g2_decap_8 FILLER_56_817 ();
 sg13g2_fill_1 FILLER_56_824 ();
 sg13g2_decap_4 FILLER_56_835 ();
 sg13g2_decap_8 FILLER_56_843 ();
 sg13g2_decap_4 FILLER_56_850 ();
 sg13g2_fill_2 FILLER_56_854 ();
 sg13g2_fill_2 FILLER_56_861 ();
 sg13g2_fill_2 FILLER_56_867 ();
 sg13g2_fill_1 FILLER_56_869 ();
 sg13g2_fill_2 FILLER_56_874 ();
 sg13g2_fill_1 FILLER_56_876 ();
 sg13g2_fill_2 FILLER_56_882 ();
 sg13g2_fill_1 FILLER_56_901 ();
 sg13g2_decap_8 FILLER_56_922 ();
 sg13g2_decap_8 FILLER_56_939 ();
 sg13g2_decap_8 FILLER_56_946 ();
 sg13g2_decap_4 FILLER_56_953 ();
 sg13g2_decap_4 FILLER_56_966 ();
 sg13g2_decap_8 FILLER_56_973 ();
 sg13g2_fill_2 FILLER_56_980 ();
 sg13g2_decap_8 FILLER_56_988 ();
 sg13g2_decap_8 FILLER_56_995 ();
 sg13g2_decap_4 FILLER_56_1002 ();
 sg13g2_fill_2 FILLER_56_1006 ();
 sg13g2_fill_2 FILLER_56_1017 ();
 sg13g2_fill_2 FILLER_56_1023 ();
 sg13g2_fill_2 FILLER_56_1029 ();
 sg13g2_fill_2 FILLER_56_1035 ();
 sg13g2_decap_8 FILLER_56_1042 ();
 sg13g2_decap_4 FILLER_56_1055 ();
 sg13g2_fill_1 FILLER_56_1059 ();
 sg13g2_fill_1 FILLER_56_1071 ();
 sg13g2_fill_2 FILLER_56_1085 ();
 sg13g2_decap_4 FILLER_56_1100 ();
 sg13g2_decap_8 FILLER_56_1128 ();
 sg13g2_fill_2 FILLER_56_1135 ();
 sg13g2_decap_8 FILLER_56_1151 ();
 sg13g2_fill_1 FILLER_56_1158 ();
 sg13g2_fill_2 FILLER_56_1175 ();
 sg13g2_fill_2 FILLER_56_1181 ();
 sg13g2_fill_1 FILLER_56_1183 ();
 sg13g2_fill_1 FILLER_56_1188 ();
 sg13g2_fill_2 FILLER_56_1193 ();
 sg13g2_fill_1 FILLER_56_1195 ();
 sg13g2_decap_4 FILLER_56_1200 ();
 sg13g2_fill_1 FILLER_56_1218 ();
 sg13g2_fill_2 FILLER_56_1242 ();
 sg13g2_decap_4 FILLER_56_1277 ();
 sg13g2_fill_2 FILLER_56_1281 ();
 sg13g2_decap_8 FILLER_56_1305 ();
 sg13g2_decap_8 FILLER_56_1312 ();
 sg13g2_decap_8 FILLER_56_1319 ();
 sg13g2_decap_8 FILLER_57_26 ();
 sg13g2_fill_2 FILLER_57_37 ();
 sg13g2_fill_2 FILLER_57_47 ();
 sg13g2_fill_2 FILLER_57_71 ();
 sg13g2_fill_2 FILLER_57_79 ();
 sg13g2_fill_1 FILLER_57_81 ();
 sg13g2_decap_8 FILLER_57_87 ();
 sg13g2_decap_8 FILLER_57_94 ();
 sg13g2_decap_8 FILLER_57_101 ();
 sg13g2_decap_8 FILLER_57_108 ();
 sg13g2_decap_8 FILLER_57_115 ();
 sg13g2_decap_8 FILLER_57_122 ();
 sg13g2_decap_4 FILLER_57_129 ();
 sg13g2_fill_1 FILLER_57_133 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_decap_4 FILLER_57_152 ();
 sg13g2_fill_1 FILLER_57_156 ();
 sg13g2_decap_8 FILLER_57_163 ();
 sg13g2_fill_1 FILLER_57_170 ();
 sg13g2_decap_4 FILLER_57_177 ();
 sg13g2_fill_1 FILLER_57_181 ();
 sg13g2_fill_2 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_220 ();
 sg13g2_decap_8 FILLER_57_227 ();
 sg13g2_fill_1 FILLER_57_234 ();
 sg13g2_fill_1 FILLER_57_238 ();
 sg13g2_decap_8 FILLER_57_248 ();
 sg13g2_decap_8 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_267 ();
 sg13g2_decap_4 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_277 ();
 sg13g2_decap_4 FILLER_57_283 ();
 sg13g2_fill_1 FILLER_57_294 ();
 sg13g2_decap_4 FILLER_57_301 ();
 sg13g2_fill_2 FILLER_57_305 ();
 sg13g2_fill_1 FILLER_57_310 ();
 sg13g2_fill_2 FILLER_57_315 ();
 sg13g2_fill_2 FILLER_57_320 ();
 sg13g2_fill_2 FILLER_57_328 ();
 sg13g2_fill_1 FILLER_57_338 ();
 sg13g2_fill_1 FILLER_57_342 ();
 sg13g2_fill_1 FILLER_57_347 ();
 sg13g2_fill_1 FILLER_57_352 ();
 sg13g2_fill_1 FILLER_57_366 ();
 sg13g2_fill_2 FILLER_57_376 ();
 sg13g2_fill_1 FILLER_57_378 ();
 sg13g2_fill_2 FILLER_57_383 ();
 sg13g2_fill_1 FILLER_57_385 ();
 sg13g2_fill_1 FILLER_57_390 ();
 sg13g2_fill_2 FILLER_57_409 ();
 sg13g2_decap_4 FILLER_57_416 ();
 sg13g2_fill_1 FILLER_57_435 ();
 sg13g2_decap_4 FILLER_57_459 ();
 sg13g2_fill_1 FILLER_57_463 ();
 sg13g2_decap_8 FILLER_57_488 ();
 sg13g2_fill_2 FILLER_57_495 ();
 sg13g2_fill_1 FILLER_57_497 ();
 sg13g2_decap_8 FILLER_57_504 ();
 sg13g2_decap_8 FILLER_57_511 ();
 sg13g2_decap_8 FILLER_57_518 ();
 sg13g2_fill_2 FILLER_57_525 ();
 sg13g2_fill_1 FILLER_57_527 ();
 sg13g2_fill_1 FILLER_57_532 ();
 sg13g2_decap_4 FILLER_57_547 ();
 sg13g2_fill_1 FILLER_57_559 ();
 sg13g2_decap_4 FILLER_57_573 ();
 sg13g2_decap_4 FILLER_57_582 ();
 sg13g2_fill_1 FILLER_57_586 ();
 sg13g2_decap_8 FILLER_57_601 ();
 sg13g2_decap_4 FILLER_57_608 ();
 sg13g2_fill_1 FILLER_57_616 ();
 sg13g2_decap_4 FILLER_57_621 ();
 sg13g2_fill_1 FILLER_57_643 ();
 sg13g2_fill_1 FILLER_57_649 ();
 sg13g2_fill_2 FILLER_57_654 ();
 sg13g2_decap_8 FILLER_57_660 ();
 sg13g2_decap_8 FILLER_57_667 ();
 sg13g2_fill_2 FILLER_57_674 ();
 sg13g2_fill_2 FILLER_57_680 ();
 sg13g2_decap_8 FILLER_57_685 ();
 sg13g2_fill_2 FILLER_57_692 ();
 sg13g2_fill_1 FILLER_57_694 ();
 sg13g2_decap_4 FILLER_57_699 ();
 sg13g2_decap_4 FILLER_57_711 ();
 sg13g2_fill_1 FILLER_57_715 ();
 sg13g2_fill_1 FILLER_57_722 ();
 sg13g2_decap_8 FILLER_57_741 ();
 sg13g2_decap_8 FILLER_57_748 ();
 sg13g2_decap_8 FILLER_57_755 ();
 sg13g2_decap_8 FILLER_57_762 ();
 sg13g2_decap_8 FILLER_57_769 ();
 sg13g2_fill_1 FILLER_57_776 ();
 sg13g2_decap_8 FILLER_57_789 ();
 sg13g2_fill_1 FILLER_57_796 ();
 sg13g2_decap_8 FILLER_57_803 ();
 sg13g2_fill_2 FILLER_57_816 ();
 sg13g2_fill_1 FILLER_57_818 ();
 sg13g2_decap_4 FILLER_57_845 ();
 sg13g2_fill_1 FILLER_57_849 ();
 sg13g2_decap_4 FILLER_57_858 ();
 sg13g2_decap_8 FILLER_57_886 ();
 sg13g2_decap_8 FILLER_57_893 ();
 sg13g2_decap_8 FILLER_57_900 ();
 sg13g2_decap_8 FILLER_57_907 ();
 sg13g2_decap_8 FILLER_57_914 ();
 sg13g2_decap_4 FILLER_57_921 ();
 sg13g2_fill_1 FILLER_57_925 ();
 sg13g2_decap_8 FILLER_57_935 ();
 sg13g2_decap_8 FILLER_57_942 ();
 sg13g2_fill_1 FILLER_57_957 ();
 sg13g2_decap_4 FILLER_57_961 ();
 sg13g2_fill_2 FILLER_57_965 ();
 sg13g2_decap_8 FILLER_57_998 ();
 sg13g2_fill_1 FILLER_57_1005 ();
 sg13g2_decap_8 FILLER_57_1015 ();
 sg13g2_decap_4 FILLER_57_1022 ();
 sg13g2_decap_8 FILLER_57_1036 ();
 sg13g2_decap_4 FILLER_57_1043 ();
 sg13g2_decap_8 FILLER_57_1060 ();
 sg13g2_decap_4 FILLER_57_1067 ();
 sg13g2_fill_1 FILLER_57_1074 ();
 sg13g2_fill_2 FILLER_57_1083 ();
 sg13g2_fill_1 FILLER_57_1088 ();
 sg13g2_decap_4 FILLER_57_1101 ();
 sg13g2_fill_1 FILLER_57_1115 ();
 sg13g2_fill_1 FILLER_57_1120 ();
 sg13g2_fill_1 FILLER_57_1142 ();
 sg13g2_fill_1 FILLER_57_1147 ();
 sg13g2_fill_1 FILLER_57_1156 ();
 sg13g2_fill_2 FILLER_57_1162 ();
 sg13g2_fill_2 FILLER_57_1173 ();
 sg13g2_fill_2 FILLER_57_1185 ();
 sg13g2_decap_8 FILLER_57_1197 ();
 sg13g2_decap_8 FILLER_57_1204 ();
 sg13g2_fill_2 FILLER_57_1225 ();
 sg13g2_decap_4 FILLER_57_1232 ();
 sg13g2_fill_1 FILLER_57_1236 ();
 sg13g2_decap_8 FILLER_57_1257 ();
 sg13g2_fill_2 FILLER_57_1264 ();
 sg13g2_fill_1 FILLER_57_1266 ();
 sg13g2_decap_4 FILLER_57_1271 ();
 sg13g2_fill_1 FILLER_57_1279 ();
 sg13g2_fill_2 FILLER_57_1296 ();
 sg13g2_decap_8 FILLER_57_1303 ();
 sg13g2_decap_8 FILLER_57_1310 ();
 sg13g2_decap_8 FILLER_57_1317 ();
 sg13g2_fill_2 FILLER_57_1324 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_4 FILLER_58_14 ();
 sg13g2_fill_2 FILLER_58_18 ();
 sg13g2_fill_1 FILLER_58_23 ();
 sg13g2_fill_1 FILLER_58_29 ();
 sg13g2_fill_1 FILLER_58_39 ();
 sg13g2_fill_1 FILLER_58_58 ();
 sg13g2_decap_8 FILLER_58_75 ();
 sg13g2_decap_8 FILLER_58_82 ();
 sg13g2_decap_8 FILLER_58_89 ();
 sg13g2_decap_8 FILLER_58_96 ();
 sg13g2_decap_8 FILLER_58_103 ();
 sg13g2_decap_4 FILLER_58_110 ();
 sg13g2_fill_1 FILLER_58_114 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_4 FILLER_58_126 ();
 sg13g2_fill_2 FILLER_58_130 ();
 sg13g2_fill_2 FILLER_58_146 ();
 sg13g2_fill_2 FILLER_58_153 ();
 sg13g2_fill_1 FILLER_58_155 ();
 sg13g2_fill_1 FILLER_58_161 ();
 sg13g2_fill_2 FILLER_58_167 ();
 sg13g2_fill_1 FILLER_58_169 ();
 sg13g2_decap_4 FILLER_58_185 ();
 sg13g2_fill_1 FILLER_58_189 ();
 sg13g2_decap_4 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_212 ();
 sg13g2_fill_1 FILLER_58_219 ();
 sg13g2_fill_2 FILLER_58_228 ();
 sg13g2_fill_2 FILLER_58_240 ();
 sg13g2_fill_2 FILLER_58_259 ();
 sg13g2_decap_4 FILLER_58_270 ();
 sg13g2_fill_1 FILLER_58_274 ();
 sg13g2_fill_1 FILLER_58_278 ();
 sg13g2_fill_2 FILLER_58_285 ();
 sg13g2_decap_8 FILLER_58_291 ();
 sg13g2_fill_1 FILLER_58_298 ();
 sg13g2_fill_1 FILLER_58_304 ();
 sg13g2_decap_4 FILLER_58_317 ();
 sg13g2_fill_2 FILLER_58_321 ();
 sg13g2_decap_8 FILLER_58_332 ();
 sg13g2_decap_4 FILLER_58_339 ();
 sg13g2_fill_2 FILLER_58_347 ();
 sg13g2_decap_8 FILLER_58_363 ();
 sg13g2_decap_8 FILLER_58_370 ();
 sg13g2_decap_4 FILLER_58_377 ();
 sg13g2_decap_8 FILLER_58_388 ();
 sg13g2_decap_4 FILLER_58_395 ();
 sg13g2_fill_1 FILLER_58_399 ();
 sg13g2_decap_8 FILLER_58_403 ();
 sg13g2_decap_8 FILLER_58_410 ();
 sg13g2_decap_4 FILLER_58_434 ();
 sg13g2_fill_2 FILLER_58_438 ();
 sg13g2_fill_2 FILLER_58_451 ();
 sg13g2_fill_1 FILLER_58_453 ();
 sg13g2_decap_8 FILLER_58_480 ();
 sg13g2_decap_8 FILLER_58_487 ();
 sg13g2_fill_1 FILLER_58_494 ();
 sg13g2_decap_8 FILLER_58_499 ();
 sg13g2_decap_4 FILLER_58_506 ();
 sg13g2_fill_2 FILLER_58_523 ();
 sg13g2_fill_1 FILLER_58_525 ();
 sg13g2_decap_4 FILLER_58_531 ();
 sg13g2_fill_2 FILLER_58_540 ();
 sg13g2_fill_2 FILLER_58_550 ();
 sg13g2_fill_2 FILLER_58_557 ();
 sg13g2_fill_2 FILLER_58_573 ();
 sg13g2_fill_2 FILLER_58_579 ();
 sg13g2_fill_1 FILLER_58_585 ();
 sg13g2_decap_8 FILLER_58_622 ();
 sg13g2_decap_4 FILLER_58_629 ();
 sg13g2_fill_1 FILLER_58_637 ();
 sg13g2_fill_1 FILLER_58_642 ();
 sg13g2_fill_1 FILLER_58_654 ();
 sg13g2_fill_1 FILLER_58_661 ();
 sg13g2_decap_8 FILLER_58_666 ();
 sg13g2_decap_8 FILLER_58_673 ();
 sg13g2_decap_8 FILLER_58_680 ();
 sg13g2_decap_8 FILLER_58_687 ();
 sg13g2_decap_8 FILLER_58_694 ();
 sg13g2_decap_4 FILLER_58_701 ();
 sg13g2_fill_1 FILLER_58_705 ();
 sg13g2_fill_1 FILLER_58_709 ();
 sg13g2_decap_4 FILLER_58_714 ();
 sg13g2_fill_2 FILLER_58_718 ();
 sg13g2_fill_2 FILLER_58_729 ();
 sg13g2_fill_1 FILLER_58_731 ();
 sg13g2_fill_1 FILLER_58_738 ();
 sg13g2_fill_1 FILLER_58_744 ();
 sg13g2_fill_2 FILLER_58_749 ();
 sg13g2_fill_1 FILLER_58_754 ();
 sg13g2_decap_4 FILLER_58_760 ();
 sg13g2_fill_2 FILLER_58_774 ();
 sg13g2_fill_1 FILLER_58_776 ();
 sg13g2_decap_4 FILLER_58_793 ();
 sg13g2_fill_1 FILLER_58_797 ();
 sg13g2_fill_1 FILLER_58_825 ();
 sg13g2_fill_2 FILLER_58_832 ();
 sg13g2_fill_2 FILLER_58_840 ();
 sg13g2_fill_1 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_846 ();
 sg13g2_fill_1 FILLER_58_853 ();
 sg13g2_fill_1 FILLER_58_867 ();
 sg13g2_fill_2 FILLER_58_874 ();
 sg13g2_fill_1 FILLER_58_876 ();
 sg13g2_decap_8 FILLER_58_905 ();
 sg13g2_decap_8 FILLER_58_912 ();
 sg13g2_decap_4 FILLER_58_919 ();
 sg13g2_fill_2 FILLER_58_927 ();
 sg13g2_fill_2 FILLER_58_971 ();
 sg13g2_fill_1 FILLER_58_973 ();
 sg13g2_decap_4 FILLER_58_982 ();
 sg13g2_fill_1 FILLER_58_986 ();
 sg13g2_decap_4 FILLER_58_990 ();
 sg13g2_decap_8 FILLER_58_1001 ();
 sg13g2_decap_8 FILLER_58_1008 ();
 sg13g2_fill_2 FILLER_58_1015 ();
 sg13g2_fill_1 FILLER_58_1020 ();
 sg13g2_fill_2 FILLER_58_1026 ();
 sg13g2_decap_4 FILLER_58_1033 ();
 sg13g2_fill_1 FILLER_58_1037 ();
 sg13g2_decap_4 FILLER_58_1048 ();
 sg13g2_decap_4 FILLER_58_1064 ();
 sg13g2_fill_1 FILLER_58_1068 ();
 sg13g2_fill_1 FILLER_58_1077 ();
 sg13g2_decap_4 FILLER_58_1086 ();
 sg13g2_fill_2 FILLER_58_1090 ();
 sg13g2_decap_4 FILLER_58_1096 ();
 sg13g2_fill_1 FILLER_58_1100 ();
 sg13g2_decap_4 FILLER_58_1106 ();
 sg13g2_fill_1 FILLER_58_1110 ();
 sg13g2_decap_4 FILLER_58_1121 ();
 sg13g2_fill_2 FILLER_58_1129 ();
 sg13g2_fill_2 FILLER_58_1134 ();
 sg13g2_decap_8 FILLER_58_1144 ();
 sg13g2_decap_4 FILLER_58_1155 ();
 sg13g2_decap_8 FILLER_58_1162 ();
 sg13g2_decap_4 FILLER_58_1169 ();
 sg13g2_fill_1 FILLER_58_1173 ();
 sg13g2_fill_1 FILLER_58_1201 ();
 sg13g2_fill_1 FILLER_58_1205 ();
 sg13g2_decap_4 FILLER_58_1210 ();
 sg13g2_fill_2 FILLER_58_1222 ();
 sg13g2_decap_4 FILLER_58_1239 ();
 sg13g2_fill_1 FILLER_58_1243 ();
 sg13g2_fill_2 FILLER_58_1252 ();
 sg13g2_decap_8 FILLER_58_1258 ();
 sg13g2_fill_1 FILLER_58_1269 ();
 sg13g2_decap_4 FILLER_58_1273 ();
 sg13g2_fill_1 FILLER_58_1277 ();
 sg13g2_decap_8 FILLER_58_1284 ();
 sg13g2_fill_2 FILLER_58_1291 ();
 sg13g2_fill_1 FILLER_58_1293 ();
 sg13g2_fill_2 FILLER_58_1298 ();
 sg13g2_decap_4 FILLER_59_39 ();
 sg13g2_decap_4 FILLER_59_51 ();
 sg13g2_fill_1 FILLER_59_55 ();
 sg13g2_decap_8 FILLER_59_75 ();
 sg13g2_decap_4 FILLER_59_82 ();
 sg13g2_fill_2 FILLER_59_112 ();
 sg13g2_fill_2 FILLER_59_143 ();
 sg13g2_fill_1 FILLER_59_156 ();
 sg13g2_decap_4 FILLER_59_185 ();
 sg13g2_fill_1 FILLER_59_189 ();
 sg13g2_decap_4 FILLER_59_198 ();
 sg13g2_fill_1 FILLER_59_202 ();
 sg13g2_decap_8 FILLER_59_207 ();
 sg13g2_fill_2 FILLER_59_214 ();
 sg13g2_fill_1 FILLER_59_216 ();
 sg13g2_fill_2 FILLER_59_233 ();
 sg13g2_decap_8 FILLER_59_252 ();
 sg13g2_fill_1 FILLER_59_259 ();
 sg13g2_decap_4 FILLER_59_263 ();
 sg13g2_fill_1 FILLER_59_267 ();
 sg13g2_fill_2 FILLER_59_286 ();
 sg13g2_fill_1 FILLER_59_291 ();
 sg13g2_fill_1 FILLER_59_297 ();
 sg13g2_fill_1 FILLER_59_304 ();
 sg13g2_decap_8 FILLER_59_313 ();
 sg13g2_fill_2 FILLER_59_345 ();
 sg13g2_decap_4 FILLER_59_357 ();
 sg13g2_fill_2 FILLER_59_361 ();
 sg13g2_fill_2 FILLER_59_367 ();
 sg13g2_decap_8 FILLER_59_372 ();
 sg13g2_decap_4 FILLER_59_379 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_fill_2 FILLER_59_399 ();
 sg13g2_fill_1 FILLER_59_401 ();
 sg13g2_fill_1 FILLER_59_413 ();
 sg13g2_decap_4 FILLER_59_419 ();
 sg13g2_fill_2 FILLER_59_423 ();
 sg13g2_fill_2 FILLER_59_433 ();
 sg13g2_decap_4 FILLER_59_455 ();
 sg13g2_fill_1 FILLER_59_459 ();
 sg13g2_decap_8 FILLER_59_465 ();
 sg13g2_decap_4 FILLER_59_472 ();
 sg13g2_fill_2 FILLER_59_476 ();
 sg13g2_decap_4 FILLER_59_481 ();
 sg13g2_fill_2 FILLER_59_485 ();
 sg13g2_decap_8 FILLER_59_499 ();
 sg13g2_fill_2 FILLER_59_511 ();
 sg13g2_fill_1 FILLER_59_513 ();
 sg13g2_decap_8 FILLER_59_523 ();
 sg13g2_decap_8 FILLER_59_530 ();
 sg13g2_decap_4 FILLER_59_537 ();
 sg13g2_fill_2 FILLER_59_541 ();
 sg13g2_decap_4 FILLER_59_546 ();
 sg13g2_fill_1 FILLER_59_555 ();
 sg13g2_fill_1 FILLER_59_561 ();
 sg13g2_decap_4 FILLER_59_567 ();
 sg13g2_fill_1 FILLER_59_591 ();
 sg13g2_decap_4 FILLER_59_603 ();
 sg13g2_fill_2 FILLER_59_607 ();
 sg13g2_fill_1 FILLER_59_614 ();
 sg13g2_fill_2 FILLER_59_620 ();
 sg13g2_fill_1 FILLER_59_635 ();
 sg13g2_fill_1 FILLER_59_647 ();
 sg13g2_fill_2 FILLER_59_653 ();
 sg13g2_decap_4 FILLER_59_664 ();
 sg13g2_fill_2 FILLER_59_668 ();
 sg13g2_fill_1 FILLER_59_703 ();
 sg13g2_decap_4 FILLER_59_708 ();
 sg13g2_fill_1 FILLER_59_716 ();
 sg13g2_fill_1 FILLER_59_738 ();
 sg13g2_fill_2 FILLER_59_742 ();
 sg13g2_fill_1 FILLER_59_744 ();
 sg13g2_decap_8 FILLER_59_750 ();
 sg13g2_fill_1 FILLER_59_757 ();
 sg13g2_fill_1 FILLER_59_761 ();
 sg13g2_fill_1 FILLER_59_767 ();
 sg13g2_fill_1 FILLER_59_781 ();
 sg13g2_fill_2 FILLER_59_787 ();
 sg13g2_fill_1 FILLER_59_789 ();
 sg13g2_decap_8 FILLER_59_795 ();
 sg13g2_decap_8 FILLER_59_802 ();
 sg13g2_decap_8 FILLER_59_809 ();
 sg13g2_decap_4 FILLER_59_816 ();
 sg13g2_fill_2 FILLER_59_820 ();
 sg13g2_decap_4 FILLER_59_826 ();
 sg13g2_fill_2 FILLER_59_830 ();
 sg13g2_fill_2 FILLER_59_842 ();
 sg13g2_fill_1 FILLER_59_844 ();
 sg13g2_decap_8 FILLER_59_862 ();
 sg13g2_decap_8 FILLER_59_869 ();
 sg13g2_fill_2 FILLER_59_876 ();
 sg13g2_fill_1 FILLER_59_878 ();
 sg13g2_decap_4 FILLER_59_895 ();
 sg13g2_decap_8 FILLER_59_924 ();
 sg13g2_decap_4 FILLER_59_931 ();
 sg13g2_fill_2 FILLER_59_939 ();
 sg13g2_decap_4 FILLER_59_945 ();
 sg13g2_fill_1 FILLER_59_952 ();
 sg13g2_fill_1 FILLER_59_957 ();
 sg13g2_decap_4 FILLER_59_963 ();
 sg13g2_fill_1 FILLER_59_967 ();
 sg13g2_decap_4 FILLER_59_972 ();
 sg13g2_decap_4 FILLER_59_985 ();
 sg13g2_fill_2 FILLER_59_997 ();
 sg13g2_fill_1 FILLER_59_999 ();
 sg13g2_fill_1 FILLER_59_1005 ();
 sg13g2_decap_4 FILLER_59_1059 ();
 sg13g2_fill_2 FILLER_59_1063 ();
 sg13g2_fill_1 FILLER_59_1070 ();
 sg13g2_decap_4 FILLER_59_1075 ();
 sg13g2_decap_8 FILLER_59_1084 ();
 sg13g2_fill_2 FILLER_59_1091 ();
 sg13g2_fill_2 FILLER_59_1138 ();
 sg13g2_fill_1 FILLER_59_1140 ();
 sg13g2_decap_8 FILLER_59_1146 ();
 sg13g2_decap_8 FILLER_59_1153 ();
 sg13g2_decap_4 FILLER_59_1160 ();
 sg13g2_decap_8 FILLER_59_1174 ();
 sg13g2_decap_8 FILLER_59_1181 ();
 sg13g2_decap_8 FILLER_59_1188 ();
 sg13g2_decap_8 FILLER_59_1195 ();
 sg13g2_fill_2 FILLER_59_1202 ();
 sg13g2_fill_1 FILLER_59_1204 ();
 sg13g2_fill_2 FILLER_59_1209 ();
 sg13g2_fill_1 FILLER_59_1211 ();
 sg13g2_fill_1 FILLER_59_1219 ();
 sg13g2_decap_8 FILLER_59_1225 ();
 sg13g2_decap_8 FILLER_59_1232 ();
 sg13g2_decap_8 FILLER_59_1239 ();
 sg13g2_decap_8 FILLER_59_1246 ();
 sg13g2_decap_4 FILLER_59_1253 ();
 sg13g2_fill_1 FILLER_59_1262 ();
 sg13g2_fill_2 FILLER_59_1267 ();
 sg13g2_fill_1 FILLER_59_1274 ();
 sg13g2_fill_1 FILLER_59_1279 ();
 sg13g2_fill_1 FILLER_59_1289 ();
 sg13g2_fill_1 FILLER_59_1294 ();
 sg13g2_fill_2 FILLER_59_1300 ();
 sg13g2_fill_1 FILLER_59_1302 ();
 sg13g2_decap_8 FILLER_59_1311 ();
 sg13g2_decap_8 FILLER_59_1318 ();
 sg13g2_fill_1 FILLER_59_1325 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_4 FILLER_60_31 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_fill_1 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_83 ();
 sg13g2_decap_8 FILLER_60_90 ();
 sg13g2_decap_8 FILLER_60_97 ();
 sg13g2_fill_2 FILLER_60_104 ();
 sg13g2_fill_1 FILLER_60_119 ();
 sg13g2_fill_1 FILLER_60_152 ();
 sg13g2_fill_1 FILLER_60_163 ();
 sg13g2_fill_1 FILLER_60_170 ();
 sg13g2_fill_1 FILLER_60_178 ();
 sg13g2_fill_1 FILLER_60_184 ();
 sg13g2_fill_2 FILLER_60_211 ();
 sg13g2_fill_2 FILLER_60_228 ();
 sg13g2_fill_2 FILLER_60_242 ();
 sg13g2_decap_4 FILLER_60_249 ();
 sg13g2_fill_1 FILLER_60_265 ();
 sg13g2_fill_1 FILLER_60_280 ();
 sg13g2_decap_4 FILLER_60_289 ();
 sg13g2_decap_4 FILLER_60_296 ();
 sg13g2_fill_2 FILLER_60_305 ();
 sg13g2_fill_1 FILLER_60_307 ();
 sg13g2_decap_8 FILLER_60_314 ();
 sg13g2_decap_8 FILLER_60_321 ();
 sg13g2_decap_8 FILLER_60_328 ();
 sg13g2_decap_8 FILLER_60_335 ();
 sg13g2_fill_2 FILLER_60_342 ();
 sg13g2_fill_1 FILLER_60_344 ();
 sg13g2_decap_8 FILLER_60_355 ();
 sg13g2_fill_2 FILLER_60_370 ();
 sg13g2_fill_1 FILLER_60_372 ();
 sg13g2_decap_4 FILLER_60_382 ();
 sg13g2_fill_2 FILLER_60_390 ();
 sg13g2_fill_1 FILLER_60_430 ();
 sg13g2_fill_1 FILLER_60_434 ();
 sg13g2_decap_8 FILLER_60_439 ();
 sg13g2_fill_1 FILLER_60_446 ();
 sg13g2_fill_2 FILLER_60_455 ();
 sg13g2_fill_1 FILLER_60_457 ();
 sg13g2_decap_8 FILLER_60_462 ();
 sg13g2_decap_8 FILLER_60_480 ();
 sg13g2_decap_8 FILLER_60_487 ();
 sg13g2_decap_8 FILLER_60_494 ();
 sg13g2_decap_4 FILLER_60_508 ();
 sg13g2_fill_2 FILLER_60_512 ();
 sg13g2_fill_2 FILLER_60_526 ();
 sg13g2_fill_2 FILLER_60_551 ();
 sg13g2_fill_2 FILLER_60_558 ();
 sg13g2_fill_2 FILLER_60_568 ();
 sg13g2_decap_8 FILLER_60_587 ();
 sg13g2_decap_8 FILLER_60_594 ();
 sg13g2_decap_4 FILLER_60_601 ();
 sg13g2_fill_1 FILLER_60_605 ();
 sg13g2_decap_8 FILLER_60_616 ();
 sg13g2_decap_8 FILLER_60_628 ();
 sg13g2_decap_8 FILLER_60_635 ();
 sg13g2_decap_4 FILLER_60_642 ();
 sg13g2_fill_1 FILLER_60_646 ();
 sg13g2_decap_8 FILLER_60_655 ();
 sg13g2_decap_8 FILLER_60_662 ();
 sg13g2_fill_2 FILLER_60_669 ();
 sg13g2_decap_8 FILLER_60_684 ();
 sg13g2_decap_4 FILLER_60_691 ();
 sg13g2_fill_1 FILLER_60_695 ();
 sg13g2_decap_8 FILLER_60_703 ();
 sg13g2_fill_2 FILLER_60_710 ();
 sg13g2_fill_1 FILLER_60_712 ();
 sg13g2_decap_4 FILLER_60_725 ();
 sg13g2_fill_1 FILLER_60_746 ();
 sg13g2_decap_8 FILLER_60_752 ();
 sg13g2_fill_1 FILLER_60_764 ();
 sg13g2_fill_2 FILLER_60_778 ();
 sg13g2_fill_1 FILLER_60_780 ();
 sg13g2_decap_8 FILLER_60_790 ();
 sg13g2_decap_8 FILLER_60_797 ();
 sg13g2_fill_2 FILLER_60_804 ();
 sg13g2_fill_1 FILLER_60_806 ();
 sg13g2_decap_4 FILLER_60_812 ();
 sg13g2_decap_4 FILLER_60_819 ();
 sg13g2_fill_1 FILLER_60_823 ();
 sg13g2_fill_1 FILLER_60_856 ();
 sg13g2_fill_1 FILLER_60_864 ();
 sg13g2_decap_8 FILLER_60_869 ();
 sg13g2_fill_2 FILLER_60_876 ();
 sg13g2_fill_1 FILLER_60_878 ();
 sg13g2_fill_2 FILLER_60_887 ();
 sg13g2_fill_2 FILLER_60_894 ();
 sg13g2_fill_1 FILLER_60_896 ();
 sg13g2_fill_1 FILLER_60_902 ();
 sg13g2_fill_2 FILLER_60_907 ();
 sg13g2_fill_1 FILLER_60_909 ();
 sg13g2_fill_2 FILLER_60_926 ();
 sg13g2_fill_2 FILLER_60_933 ();
 sg13g2_fill_1 FILLER_60_935 ();
 sg13g2_decap_8 FILLER_60_940 ();
 sg13g2_fill_2 FILLER_60_947 ();
 sg13g2_decap_8 FILLER_60_953 ();
 sg13g2_decap_4 FILLER_60_960 ();
 sg13g2_fill_1 FILLER_60_964 ();
 sg13g2_decap_4 FILLER_60_968 ();
 sg13g2_fill_2 FILLER_60_980 ();
 sg13g2_decap_8 FILLER_60_986 ();
 sg13g2_fill_1 FILLER_60_997 ();
 sg13g2_fill_2 FILLER_60_1007 ();
 sg13g2_fill_2 FILLER_60_1014 ();
 sg13g2_fill_2 FILLER_60_1028 ();
 sg13g2_decap_8 FILLER_60_1037 ();
 sg13g2_decap_8 FILLER_60_1044 ();
 sg13g2_decap_8 FILLER_60_1051 ();
 sg13g2_decap_8 FILLER_60_1070 ();
 sg13g2_decap_8 FILLER_60_1077 ();
 sg13g2_decap_8 FILLER_60_1084 ();
 sg13g2_fill_1 FILLER_60_1091 ();
 sg13g2_decap_8 FILLER_60_1104 ();
 sg13g2_fill_2 FILLER_60_1111 ();
 sg13g2_decap_4 FILLER_60_1118 ();
 sg13g2_fill_2 FILLER_60_1122 ();
 sg13g2_fill_2 FILLER_60_1128 ();
 sg13g2_fill_1 FILLER_60_1130 ();
 sg13g2_decap_8 FILLER_60_1136 ();
 sg13g2_decap_8 FILLER_60_1143 ();
 sg13g2_decap_4 FILLER_60_1150 ();
 sg13g2_fill_2 FILLER_60_1154 ();
 sg13g2_decap_8 FILLER_60_1165 ();
 sg13g2_decap_4 FILLER_60_1172 ();
 sg13g2_fill_2 FILLER_60_1176 ();
 sg13g2_fill_1 FILLER_60_1186 ();
 sg13g2_fill_2 FILLER_60_1191 ();
 sg13g2_fill_2 FILLER_60_1197 ();
 sg13g2_decap_4 FILLER_60_1209 ();
 sg13g2_fill_1 FILLER_60_1245 ();
 sg13g2_decap_8 FILLER_60_1267 ();
 sg13g2_fill_2 FILLER_60_1274 ();
 sg13g2_fill_1 FILLER_60_1276 ();
 sg13g2_fill_2 FILLER_60_1284 ();
 sg13g2_decap_8 FILLER_60_1290 ();
 sg13g2_decap_8 FILLER_60_1297 ();
 sg13g2_decap_8 FILLER_60_1304 ();
 sg13g2_decap_8 FILLER_60_1311 ();
 sg13g2_decap_8 FILLER_60_1318 ();
 sg13g2_fill_1 FILLER_60_1325 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_fill_1 FILLER_61_54 ();
 sg13g2_fill_1 FILLER_61_80 ();
 sg13g2_fill_2 FILLER_61_140 ();
 sg13g2_fill_1 FILLER_61_149 ();
 sg13g2_decap_8 FILLER_61_178 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_decap_4 FILLER_61_202 ();
 sg13g2_decap_8 FILLER_61_209 ();
 sg13g2_decap_4 FILLER_61_216 ();
 sg13g2_fill_1 FILLER_61_220 ();
 sg13g2_fill_2 FILLER_61_229 ();
 sg13g2_fill_2 FILLER_61_235 ();
 sg13g2_decap_4 FILLER_61_242 ();
 sg13g2_fill_2 FILLER_61_246 ();
 sg13g2_fill_2 FILLER_61_258 ();
 sg13g2_fill_1 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_267 ();
 sg13g2_fill_1 FILLER_61_271 ();
 sg13g2_decap_8 FILLER_61_275 ();
 sg13g2_fill_2 FILLER_61_282 ();
 sg13g2_fill_1 FILLER_61_284 ();
 sg13g2_fill_1 FILLER_61_299 ();
 sg13g2_fill_1 FILLER_61_305 ();
 sg13g2_fill_1 FILLER_61_316 ();
 sg13g2_decap_8 FILLER_61_321 ();
 sg13g2_decap_4 FILLER_61_339 ();
 sg13g2_fill_2 FILLER_61_343 ();
 sg13g2_fill_1 FILLER_61_349 ();
 sg13g2_decap_4 FILLER_61_355 ();
 sg13g2_fill_1 FILLER_61_359 ();
 sg13g2_decap_8 FILLER_61_372 ();
 sg13g2_decap_4 FILLER_61_379 ();
 sg13g2_fill_2 FILLER_61_386 ();
 sg13g2_fill_1 FILLER_61_388 ();
 sg13g2_decap_4 FILLER_61_396 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_fill_2 FILLER_61_409 ();
 sg13g2_decap_4 FILLER_61_414 ();
 sg13g2_fill_2 FILLER_61_418 ();
 sg13g2_fill_2 FILLER_61_441 ();
 sg13g2_decap_4 FILLER_61_448 ();
 sg13g2_fill_2 FILLER_61_452 ();
 sg13g2_decap_4 FILLER_61_462 ();
 sg13g2_fill_1 FILLER_61_470 ();
 sg13g2_decap_8 FILLER_61_475 ();
 sg13g2_decap_4 FILLER_61_482 ();
 sg13g2_fill_1 FILLER_61_486 ();
 sg13g2_decap_4 FILLER_61_494 ();
 sg13g2_fill_1 FILLER_61_498 ();
 sg13g2_fill_2 FILLER_61_508 ();
 sg13g2_fill_1 FILLER_61_533 ();
 sg13g2_fill_1 FILLER_61_544 ();
 sg13g2_fill_2 FILLER_61_548 ();
 sg13g2_fill_2 FILLER_61_565 ();
 sg13g2_fill_2 FILLER_61_572 ();
 sg13g2_fill_2 FILLER_61_580 ();
 sg13g2_decap_8 FILLER_61_588 ();
 sg13g2_fill_2 FILLER_61_595 ();
 sg13g2_decap_4 FILLER_61_602 ();
 sg13g2_fill_1 FILLER_61_606 ();
 sg13g2_fill_2 FILLER_61_637 ();
 sg13g2_fill_1 FILLER_61_642 ();
 sg13g2_fill_2 FILLER_61_668 ();
 sg13g2_fill_2 FILLER_61_674 ();
 sg13g2_fill_1 FILLER_61_676 ();
 sg13g2_fill_2 FILLER_61_702 ();
 sg13g2_decap_4 FILLER_61_707 ();
 sg13g2_decap_4 FILLER_61_722 ();
 sg13g2_fill_1 FILLER_61_726 ();
 sg13g2_fill_1 FILLER_61_768 ();
 sg13g2_decap_4 FILLER_61_777 ();
 sg13g2_decap_8 FILLER_61_786 ();
 sg13g2_decap_8 FILLER_61_793 ();
 sg13g2_fill_2 FILLER_61_800 ();
 sg13g2_fill_1 FILLER_61_802 ();
 sg13g2_decap_4 FILLER_61_807 ();
 sg13g2_decap_8 FILLER_61_819 ();
 sg13g2_fill_1 FILLER_61_829 ();
 sg13g2_fill_2 FILLER_61_836 ();
 sg13g2_fill_2 FILLER_61_843 ();
 sg13g2_fill_2 FILLER_61_849 ();
 sg13g2_fill_1 FILLER_61_851 ();
 sg13g2_decap_4 FILLER_61_857 ();
 sg13g2_fill_1 FILLER_61_861 ();
 sg13g2_decap_8 FILLER_61_868 ();
 sg13g2_fill_1 FILLER_61_875 ();
 sg13g2_decap_4 FILLER_61_886 ();
 sg13g2_fill_2 FILLER_61_894 ();
 sg13g2_fill_1 FILLER_61_896 ();
 sg13g2_fill_2 FILLER_61_900 ();
 sg13g2_fill_2 FILLER_61_905 ();
 sg13g2_fill_1 FILLER_61_907 ();
 sg13g2_fill_2 FILLER_61_949 ();
 sg13g2_fill_2 FILLER_61_959 ();
 sg13g2_fill_1 FILLER_61_961 ();
 sg13g2_decap_4 FILLER_61_967 ();
 sg13g2_fill_2 FILLER_61_971 ();
 sg13g2_fill_2 FILLER_61_983 ();
 sg13g2_decap_4 FILLER_61_988 ();
 sg13g2_fill_2 FILLER_61_992 ();
 sg13g2_fill_1 FILLER_61_999 ();
 sg13g2_fill_1 FILLER_61_1012 ();
 sg13g2_decap_4 FILLER_61_1019 ();
 sg13g2_fill_2 FILLER_61_1026 ();
 sg13g2_fill_1 FILLER_61_1028 ();
 sg13g2_fill_1 FILLER_61_1033 ();
 sg13g2_decap_4 FILLER_61_1048 ();
 sg13g2_fill_2 FILLER_61_1055 ();
 sg13g2_fill_1 FILLER_61_1057 ();
 sg13g2_fill_2 FILLER_61_1072 ();
 sg13g2_fill_1 FILLER_61_1088 ();
 sg13g2_decap_4 FILLER_61_1092 ();
 sg13g2_fill_1 FILLER_61_1096 ();
 sg13g2_decap_8 FILLER_61_1116 ();
 sg13g2_decap_4 FILLER_61_1123 ();
 sg13g2_fill_2 FILLER_61_1127 ();
 sg13g2_decap_4 FILLER_61_1136 ();
 sg13g2_fill_2 FILLER_61_1140 ();
 sg13g2_fill_1 FILLER_61_1147 ();
 sg13g2_fill_2 FILLER_61_1151 ();
 sg13g2_fill_1 FILLER_61_1153 ();
 sg13g2_fill_1 FILLER_61_1183 ();
 sg13g2_fill_1 FILLER_61_1198 ();
 sg13g2_decap_8 FILLER_61_1213 ();
 sg13g2_fill_1 FILLER_61_1220 ();
 sg13g2_decap_4 FILLER_61_1233 ();
 sg13g2_fill_2 FILLER_61_1237 ();
 sg13g2_decap_8 FILLER_61_1256 ();
 sg13g2_fill_1 FILLER_61_1263 ();
 sg13g2_fill_2 FILLER_61_1281 ();
 sg13g2_fill_1 FILLER_61_1283 ();
 sg13g2_decap_8 FILLER_61_1292 ();
 sg13g2_fill_2 FILLER_61_1299 ();
 sg13g2_decap_4 FILLER_61_1306 ();
 sg13g2_fill_1 FILLER_61_1310 ();
 sg13g2_decap_8 FILLER_61_1315 ();
 sg13g2_decap_4 FILLER_61_1322 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_4 FILLER_62_14 ();
 sg13g2_fill_1 FILLER_62_18 ();
 sg13g2_fill_1 FILLER_62_23 ();
 sg13g2_fill_2 FILLER_62_47 ();
 sg13g2_fill_1 FILLER_62_49 ();
 sg13g2_fill_1 FILLER_62_54 ();
 sg13g2_decap_8 FILLER_62_58 ();
 sg13g2_fill_2 FILLER_62_65 ();
 sg13g2_fill_1 FILLER_62_76 ();
 sg13g2_fill_1 FILLER_62_81 ();
 sg13g2_fill_2 FILLER_62_93 ();
 sg13g2_fill_2 FILLER_62_146 ();
 sg13g2_fill_1 FILLER_62_155 ();
 sg13g2_fill_1 FILLER_62_162 ();
 sg13g2_fill_2 FILLER_62_168 ();
 sg13g2_fill_2 FILLER_62_183 ();
 sg13g2_decap_8 FILLER_62_213 ();
 sg13g2_fill_2 FILLER_62_220 ();
 sg13g2_fill_1 FILLER_62_222 ();
 sg13g2_decap_4 FILLER_62_257 ();
 sg13g2_fill_1 FILLER_62_261 ();
 sg13g2_decap_8 FILLER_62_265 ();
 sg13g2_decap_4 FILLER_62_272 ();
 sg13g2_fill_2 FILLER_62_276 ();
 sg13g2_decap_4 FILLER_62_287 ();
 sg13g2_fill_2 FILLER_62_291 ();
 sg13g2_decap_4 FILLER_62_309 ();
 sg13g2_fill_1 FILLER_62_313 ();
 sg13g2_decap_8 FILLER_62_352 ();
 sg13g2_decap_4 FILLER_62_359 ();
 sg13g2_decap_8 FILLER_62_367 ();
 sg13g2_decap_8 FILLER_62_388 ();
 sg13g2_decap_8 FILLER_62_395 ();
 sg13g2_decap_4 FILLER_62_402 ();
 sg13g2_decap_8 FILLER_62_419 ();
 sg13g2_decap_8 FILLER_62_426 ();
 sg13g2_fill_2 FILLER_62_443 ();
 sg13g2_fill_1 FILLER_62_445 ();
 sg13g2_fill_1 FILLER_62_451 ();
 sg13g2_fill_2 FILLER_62_456 ();
 sg13g2_fill_1 FILLER_62_458 ();
 sg13g2_fill_1 FILLER_62_476 ();
 sg13g2_decap_8 FILLER_62_482 ();
 sg13g2_decap_8 FILLER_62_489 ();
 sg13g2_fill_1 FILLER_62_529 ();
 sg13g2_fill_1 FILLER_62_551 ();
 sg13g2_fill_1 FILLER_62_565 ();
 sg13g2_decap_4 FILLER_62_574 ();
 sg13g2_fill_2 FILLER_62_582 ();
 sg13g2_fill_1 FILLER_62_584 ();
 sg13g2_fill_1 FILLER_62_599 ();
 sg13g2_decap_8 FILLER_62_604 ();
 sg13g2_decap_4 FILLER_62_611 ();
 sg13g2_fill_1 FILLER_62_615 ();
 sg13g2_decap_8 FILLER_62_620 ();
 sg13g2_fill_1 FILLER_62_631 ();
 sg13g2_fill_1 FILLER_62_639 ();
 sg13g2_fill_1 FILLER_62_645 ();
 sg13g2_decap_8 FILLER_62_650 ();
 sg13g2_decap_8 FILLER_62_657 ();
 sg13g2_fill_1 FILLER_62_664 ();
 sg13g2_fill_1 FILLER_62_674 ();
 sg13g2_fill_1 FILLER_62_695 ();
 sg13g2_fill_1 FILLER_62_709 ();
 sg13g2_fill_1 FILLER_62_715 ();
 sg13g2_decap_8 FILLER_62_722 ();
 sg13g2_fill_1 FILLER_62_729 ();
 sg13g2_fill_2 FILLER_62_736 ();
 sg13g2_fill_1 FILLER_62_738 ();
 sg13g2_decap_8 FILLER_62_742 ();
 sg13g2_decap_8 FILLER_62_749 ();
 sg13g2_fill_2 FILLER_62_756 ();
 sg13g2_decap_4 FILLER_62_761 ();
 sg13g2_fill_2 FILLER_62_765 ();
 sg13g2_fill_2 FILLER_62_788 ();
 sg13g2_fill_1 FILLER_62_790 ();
 sg13g2_fill_1 FILLER_62_796 ();
 sg13g2_fill_1 FILLER_62_801 ();
 sg13g2_fill_1 FILLER_62_808 ();
 sg13g2_fill_2 FILLER_62_812 ();
 sg13g2_fill_1 FILLER_62_828 ();
 sg13g2_decap_4 FILLER_62_845 ();
 sg13g2_fill_2 FILLER_62_866 ();
 sg13g2_fill_1 FILLER_62_868 ();
 sg13g2_fill_2 FILLER_62_915 ();
 sg13g2_fill_1 FILLER_62_926 ();
 sg13g2_decap_8 FILLER_62_933 ();
 sg13g2_decap_8 FILLER_62_940 ();
 sg13g2_fill_2 FILLER_62_951 ();
 sg13g2_fill_1 FILLER_62_953 ();
 sg13g2_decap_4 FILLER_62_959 ();
 sg13g2_fill_1 FILLER_62_972 ();
 sg13g2_decap_8 FILLER_62_978 ();
 sg13g2_decap_4 FILLER_62_985 ();
 sg13g2_fill_2 FILLER_62_989 ();
 sg13g2_fill_1 FILLER_62_1015 ();
 sg13g2_fill_1 FILLER_62_1021 ();
 sg13g2_fill_1 FILLER_62_1026 ();
 sg13g2_decap_8 FILLER_62_1031 ();
 sg13g2_fill_1 FILLER_62_1038 ();
 sg13g2_fill_2 FILLER_62_1045 ();
 sg13g2_fill_1 FILLER_62_1050 ();
 sg13g2_fill_1 FILLER_62_1063 ();
 sg13g2_fill_1 FILLER_62_1073 ();
 sg13g2_fill_1 FILLER_62_1089 ();
 sg13g2_fill_2 FILLER_62_1119 ();
 sg13g2_fill_1 FILLER_62_1162 ();
 sg13g2_decap_4 FILLER_62_1166 ();
 sg13g2_fill_1 FILLER_62_1170 ();
 sg13g2_decap_4 FILLER_62_1179 ();
 sg13g2_decap_8 FILLER_62_1188 ();
 sg13g2_fill_2 FILLER_62_1195 ();
 sg13g2_fill_2 FILLER_62_1205 ();
 sg13g2_fill_1 FILLER_62_1207 ();
 sg13g2_fill_1 FILLER_62_1220 ();
 sg13g2_fill_2 FILLER_62_1226 ();
 sg13g2_fill_1 FILLER_62_1228 ();
 sg13g2_decap_4 FILLER_62_1233 ();
 sg13g2_fill_2 FILLER_62_1237 ();
 sg13g2_fill_2 FILLER_62_1243 ();
 sg13g2_fill_1 FILLER_62_1245 ();
 sg13g2_decap_4 FILLER_62_1251 ();
 sg13g2_fill_2 FILLER_62_1255 ();
 sg13g2_decap_8 FILLER_62_1270 ();
 sg13g2_fill_1 FILLER_62_1277 ();
 sg13g2_decap_8 FILLER_62_1313 ();
 sg13g2_decap_4 FILLER_62_1320 ();
 sg13g2_fill_2 FILLER_62_1324 ();
 sg13g2_fill_1 FILLER_63_26 ();
 sg13g2_fill_2 FILLER_63_33 ();
 sg13g2_fill_1 FILLER_63_35 ();
 sg13g2_fill_2 FILLER_63_67 ();
 sg13g2_fill_2 FILLER_63_90 ();
 sg13g2_fill_2 FILLER_63_103 ();
 sg13g2_fill_2 FILLER_63_170 ();
 sg13g2_fill_1 FILLER_63_210 ();
 sg13g2_fill_1 FILLER_63_223 ();
 sg13g2_fill_1 FILLER_63_229 ();
 sg13g2_decap_8 FILLER_63_241 ();
 sg13g2_fill_2 FILLER_63_248 ();
 sg13g2_fill_1 FILLER_63_254 ();
 sg13g2_decap_8 FILLER_63_260 ();
 sg13g2_decap_4 FILLER_63_267 ();
 sg13g2_fill_1 FILLER_63_271 ();
 sg13g2_decap_8 FILLER_63_280 ();
 sg13g2_fill_2 FILLER_63_287 ();
 sg13g2_fill_1 FILLER_63_304 ();
 sg13g2_fill_2 FILLER_63_314 ();
 sg13g2_fill_1 FILLER_63_316 ();
 sg13g2_decap_4 FILLER_63_329 ();
 sg13g2_fill_1 FILLER_63_333 ();
 sg13g2_decap_8 FILLER_63_337 ();
 sg13g2_decap_8 FILLER_63_344 ();
 sg13g2_decap_8 FILLER_63_351 ();
 sg13g2_decap_4 FILLER_63_368 ();
 sg13g2_fill_2 FILLER_63_372 ();
 sg13g2_fill_2 FILLER_63_403 ();
 sg13g2_fill_2 FILLER_63_419 ();
 sg13g2_decap_8 FILLER_63_424 ();
 sg13g2_fill_2 FILLER_63_431 ();
 sg13g2_fill_1 FILLER_63_433 ();
 sg13g2_decap_8 FILLER_63_448 ();
 sg13g2_decap_8 FILLER_63_460 ();
 sg13g2_decap_4 FILLER_63_485 ();
 sg13g2_fill_1 FILLER_63_489 ();
 sg13g2_decap_4 FILLER_63_493 ();
 sg13g2_fill_2 FILLER_63_497 ();
 sg13g2_decap_4 FILLER_63_523 ();
 sg13g2_fill_1 FILLER_63_527 ();
 sg13g2_fill_1 FILLER_63_535 ();
 sg13g2_fill_2 FILLER_63_558 ();
 sg13g2_fill_2 FILLER_63_585 ();
 sg13g2_fill_1 FILLER_63_587 ();
 sg13g2_fill_1 FILLER_63_603 ();
 sg13g2_decap_8 FILLER_63_608 ();
 sg13g2_decap_8 FILLER_63_615 ();
 sg13g2_decap_8 FILLER_63_622 ();
 sg13g2_decap_4 FILLER_63_629 ();
 sg13g2_fill_1 FILLER_63_637 ();
 sg13g2_fill_1 FILLER_63_642 ();
 sg13g2_decap_8 FILLER_63_653 ();
 sg13g2_decap_8 FILLER_63_660 ();
 sg13g2_fill_2 FILLER_63_667 ();
 sg13g2_fill_1 FILLER_63_669 ();
 sg13g2_decap_8 FILLER_63_678 ();
 sg13g2_fill_1 FILLER_63_685 ();
 sg13g2_fill_2 FILLER_63_693 ();
 sg13g2_fill_1 FILLER_63_704 ();
 sg13g2_fill_2 FILLER_63_713 ();
 sg13g2_decap_4 FILLER_63_720 ();
 sg13g2_fill_1 FILLER_63_734 ();
 sg13g2_fill_2 FILLER_63_749 ();
 sg13g2_fill_1 FILLER_63_755 ();
 sg13g2_fill_2 FILLER_63_765 ();
 sg13g2_fill_1 FILLER_63_767 ();
 sg13g2_decap_8 FILLER_63_772 ();
 sg13g2_decap_8 FILLER_63_779 ();
 sg13g2_decap_8 FILLER_63_786 ();
 sg13g2_decap_4 FILLER_63_793 ();
 sg13g2_fill_2 FILLER_63_797 ();
 sg13g2_fill_1 FILLER_63_814 ();
 sg13g2_fill_2 FILLER_63_824 ();
 sg13g2_fill_1 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_842 ();
 sg13g2_fill_2 FILLER_63_849 ();
 sg13g2_fill_1 FILLER_63_851 ();
 sg13g2_decap_8 FILLER_63_855 ();
 sg13g2_decap_8 FILLER_63_862 ();
 sg13g2_decap_8 FILLER_63_869 ();
 sg13g2_fill_1 FILLER_63_879 ();
 sg13g2_fill_1 FILLER_63_885 ();
 sg13g2_fill_2 FILLER_63_891 ();
 sg13g2_fill_1 FILLER_63_902 ();
 sg13g2_fill_1 FILLER_63_931 ();
 sg13g2_decap_8 FILLER_63_938 ();
 sg13g2_decap_8 FILLER_63_945 ();
 sg13g2_decap_4 FILLER_63_952 ();
 sg13g2_fill_2 FILLER_63_956 ();
 sg13g2_fill_1 FILLER_63_961 ();
 sg13g2_decap_4 FILLER_63_965 ();
 sg13g2_fill_1 FILLER_63_969 ();
 sg13g2_fill_2 FILLER_63_976 ();
 sg13g2_fill_1 FILLER_63_978 ();
 sg13g2_fill_1 FILLER_63_993 ();
 sg13g2_fill_2 FILLER_63_1004 ();
 sg13g2_fill_1 FILLER_63_1011 ();
 sg13g2_fill_1 FILLER_63_1020 ();
 sg13g2_fill_2 FILLER_63_1040 ();
 sg13g2_fill_1 FILLER_63_1052 ();
 sg13g2_fill_2 FILLER_63_1061 ();
 sg13g2_fill_1 FILLER_63_1067 ();
 sg13g2_fill_1 FILLER_63_1107 ();
 sg13g2_decap_8 FILLER_63_1135 ();
 sg13g2_decap_4 FILLER_63_1142 ();
 sg13g2_fill_2 FILLER_63_1154 ();
 sg13g2_fill_1 FILLER_63_1156 ();
 sg13g2_decap_4 FILLER_63_1161 ();
 sg13g2_fill_1 FILLER_63_1165 ();
 sg13g2_fill_1 FILLER_63_1175 ();
 sg13g2_fill_2 FILLER_63_1185 ();
 sg13g2_fill_2 FILLER_63_1191 ();
 sg13g2_decap_4 FILLER_63_1197 ();
 sg13g2_fill_2 FILLER_63_1206 ();
 sg13g2_fill_2 FILLER_63_1218 ();
 sg13g2_fill_1 FILLER_63_1223 ();
 sg13g2_fill_1 FILLER_63_1242 ();
 sg13g2_decap_8 FILLER_63_1247 ();
 sg13g2_decap_4 FILLER_63_1254 ();
 sg13g2_fill_1 FILLER_63_1258 ();
 sg13g2_decap_4 FILLER_63_1263 ();
 sg13g2_decap_8 FILLER_63_1270 ();
 sg13g2_decap_8 FILLER_63_1277 ();
 sg13g2_fill_2 FILLER_63_1289 ();
 sg13g2_decap_8 FILLER_63_1295 ();
 sg13g2_decap_8 FILLER_63_1307 ();
 sg13g2_decap_8 FILLER_63_1314 ();
 sg13g2_decap_4 FILLER_63_1321 ();
 sg13g2_fill_1 FILLER_63_1325 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_14 ();
 sg13g2_fill_2 FILLER_64_40 ();
 sg13g2_fill_1 FILLER_64_42 ();
 sg13g2_fill_2 FILLER_64_48 ();
 sg13g2_fill_1 FILLER_64_50 ();
 sg13g2_fill_2 FILLER_64_65 ();
 sg13g2_fill_2 FILLER_64_111 ();
 sg13g2_decap_4 FILLER_64_117 ();
 sg13g2_fill_1 FILLER_64_121 ();
 sg13g2_fill_1 FILLER_64_127 ();
 sg13g2_fill_1 FILLER_64_173 ();
 sg13g2_fill_2 FILLER_64_193 ();
 sg13g2_fill_1 FILLER_64_200 ();
 sg13g2_fill_1 FILLER_64_219 ();
 sg13g2_fill_2 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_237 ();
 sg13g2_decap_4 FILLER_64_243 ();
 sg13g2_decap_4 FILLER_64_250 ();
 sg13g2_fill_1 FILLER_64_254 ();
 sg13g2_decap_8 FILLER_64_285 ();
 sg13g2_decap_4 FILLER_64_292 ();
 sg13g2_fill_1 FILLER_64_296 ();
 sg13g2_fill_2 FILLER_64_300 ();
 sg13g2_fill_1 FILLER_64_302 ();
 sg13g2_decap_8 FILLER_64_307 ();
 sg13g2_fill_2 FILLER_64_314 ();
 sg13g2_fill_1 FILLER_64_316 ();
 sg13g2_decap_4 FILLER_64_330 ();
 sg13g2_fill_2 FILLER_64_334 ();
 sg13g2_decap_8 FILLER_64_362 ();
 sg13g2_decap_8 FILLER_64_369 ();
 sg13g2_fill_2 FILLER_64_376 ();
 sg13g2_decap_8 FILLER_64_383 ();
 sg13g2_decap_8 FILLER_64_390 ();
 sg13g2_fill_2 FILLER_64_397 ();
 sg13g2_fill_1 FILLER_64_399 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_64_421 ();
 sg13g2_fill_1 FILLER_64_428 ();
 sg13g2_fill_2 FILLER_64_465 ();
 sg13g2_decap_8 FILLER_64_486 ();
 sg13g2_decap_8 FILLER_64_493 ();
 sg13g2_fill_1 FILLER_64_506 ();
 sg13g2_fill_1 FILLER_64_510 ();
 sg13g2_decap_8 FILLER_64_520 ();
 sg13g2_fill_2 FILLER_64_527 ();
 sg13g2_fill_1 FILLER_64_529 ();
 sg13g2_fill_1 FILLER_64_539 ();
 sg13g2_fill_2 FILLER_64_562 ();
 sg13g2_decap_8 FILLER_64_577 ();
 sg13g2_fill_1 FILLER_64_584 ();
 sg13g2_fill_1 FILLER_64_598 ();
 sg13g2_decap_8 FILLER_64_606 ();
 sg13g2_decap_8 FILLER_64_613 ();
 sg13g2_decap_8 FILLER_64_620 ();
 sg13g2_fill_1 FILLER_64_627 ();
 sg13g2_decap_4 FILLER_64_636 ();
 sg13g2_fill_2 FILLER_64_640 ();
 sg13g2_decap_4 FILLER_64_649 ();
 sg13g2_decap_4 FILLER_64_657 ();
 sg13g2_fill_1 FILLER_64_661 ();
 sg13g2_fill_2 FILLER_64_665 ();
 sg13g2_fill_1 FILLER_64_667 ();
 sg13g2_fill_1 FILLER_64_692 ();
 sg13g2_decap_4 FILLER_64_696 ();
 sg13g2_fill_2 FILLER_64_700 ();
 sg13g2_fill_1 FILLER_64_707 ();
 sg13g2_fill_1 FILLER_64_712 ();
 sg13g2_fill_2 FILLER_64_718 ();
 sg13g2_fill_1 FILLER_64_728 ();
 sg13g2_fill_2 FILLER_64_739 ();
 sg13g2_fill_1 FILLER_64_741 ();
 sg13g2_decap_4 FILLER_64_745 ();
 sg13g2_fill_2 FILLER_64_749 ();
 sg13g2_fill_1 FILLER_64_758 ();
 sg13g2_decap_8 FILLER_64_763 ();
 sg13g2_fill_2 FILLER_64_770 ();
 sg13g2_fill_1 FILLER_64_772 ();
 sg13g2_decap_4 FILLER_64_778 ();
 sg13g2_fill_1 FILLER_64_782 ();
 sg13g2_fill_1 FILLER_64_809 ();
 sg13g2_fill_2 FILLER_64_815 ();
 sg13g2_decap_8 FILLER_64_820 ();
 sg13g2_decap_4 FILLER_64_827 ();
 sg13g2_fill_2 FILLER_64_831 ();
 sg13g2_decap_8 FILLER_64_843 ();
 sg13g2_fill_1 FILLER_64_850 ();
 sg13g2_decap_8 FILLER_64_857 ();
 sg13g2_decap_8 FILLER_64_864 ();
 sg13g2_decap_8 FILLER_64_871 ();
 sg13g2_decap_8 FILLER_64_878 ();
 sg13g2_fill_2 FILLER_64_885 ();
 sg13g2_fill_1 FILLER_64_887 ();
 sg13g2_fill_2 FILLER_64_897 ();
 sg13g2_fill_1 FILLER_64_899 ();
 sg13g2_fill_2 FILLER_64_912 ();
 sg13g2_fill_1 FILLER_64_938 ();
 sg13g2_fill_2 FILLER_64_943 ();
 sg13g2_fill_2 FILLER_64_949 ();
 sg13g2_fill_1 FILLER_64_951 ();
 sg13g2_fill_1 FILLER_64_966 ();
 sg13g2_fill_2 FILLER_64_975 ();
 sg13g2_fill_1 FILLER_64_977 ();
 sg13g2_decap_4 FILLER_64_987 ();
 sg13g2_fill_2 FILLER_64_991 ();
 sg13g2_decap_8 FILLER_64_996 ();
 sg13g2_decap_4 FILLER_64_1003 ();
 sg13g2_fill_1 FILLER_64_1007 ();
 sg13g2_decap_4 FILLER_64_1013 ();
 sg13g2_fill_2 FILLER_64_1017 ();
 sg13g2_decap_4 FILLER_64_1027 ();
 sg13g2_fill_2 FILLER_64_1035 ();
 sg13g2_fill_1 FILLER_64_1037 ();
 sg13g2_fill_1 FILLER_64_1047 ();
 sg13g2_fill_1 FILLER_64_1052 ();
 sg13g2_fill_2 FILLER_64_1058 ();
 sg13g2_fill_1 FILLER_64_1089 ();
 sg13g2_fill_2 FILLER_64_1096 ();
 sg13g2_fill_1 FILLER_64_1102 ();
 sg13g2_fill_2 FILLER_64_1122 ();
 sg13g2_fill_1 FILLER_64_1129 ();
 sg13g2_decap_4 FILLER_64_1138 ();
 sg13g2_fill_2 FILLER_64_1142 ();
 sg13g2_fill_2 FILLER_64_1149 ();
 sg13g2_fill_1 FILLER_64_1151 ();
 sg13g2_decap_8 FILLER_64_1156 ();
 sg13g2_decap_4 FILLER_64_1163 ();
 sg13g2_fill_2 FILLER_64_1170 ();
 sg13g2_decap_8 FILLER_64_1181 ();
 sg13g2_fill_2 FILLER_64_1195 ();
 sg13g2_fill_2 FILLER_64_1205 ();
 sg13g2_fill_1 FILLER_64_1207 ();
 sg13g2_decap_8 FILLER_64_1211 ();
 sg13g2_decap_8 FILLER_64_1218 ();
 sg13g2_decap_8 FILLER_64_1225 ();
 sg13g2_decap_8 FILLER_64_1232 ();
 sg13g2_fill_2 FILLER_64_1239 ();
 sg13g2_fill_1 FILLER_64_1241 ();
 sg13g2_fill_2 FILLER_64_1249 ();
 sg13g2_fill_1 FILLER_64_1251 ();
 sg13g2_decap_4 FILLER_64_1264 ();
 sg13g2_fill_1 FILLER_64_1268 ();
 sg13g2_decap_8 FILLER_64_1274 ();
 sg13g2_fill_1 FILLER_64_1290 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_fill_1 FILLER_65_16 ();
 sg13g2_fill_1 FILLER_65_21 ();
 sg13g2_fill_2 FILLER_65_30 ();
 sg13g2_fill_1 FILLER_65_32 ();
 sg13g2_fill_1 FILLER_65_38 ();
 sg13g2_decap_4 FILLER_65_48 ();
 sg13g2_fill_1 FILLER_65_57 ();
 sg13g2_decap_8 FILLER_65_74 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_4 FILLER_65_105 ();
 sg13g2_fill_2 FILLER_65_114 ();
 sg13g2_fill_2 FILLER_65_165 ();
 sg13g2_fill_1 FILLER_65_178 ();
 sg13g2_fill_1 FILLER_65_184 ();
 sg13g2_fill_2 FILLER_65_190 ();
 sg13g2_fill_2 FILLER_65_197 ();
 sg13g2_fill_1 FILLER_65_220 ();
 sg13g2_fill_2 FILLER_65_226 ();
 sg13g2_fill_1 FILLER_65_228 ();
 sg13g2_fill_1 FILLER_65_243 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_decap_8 FILLER_65_258 ();
 sg13g2_decap_4 FILLER_65_265 ();
 sg13g2_fill_2 FILLER_65_269 ();
 sg13g2_fill_2 FILLER_65_275 ();
 sg13g2_fill_1 FILLER_65_289 ();
 sg13g2_fill_1 FILLER_65_299 ();
 sg13g2_fill_2 FILLER_65_309 ();
 sg13g2_decap_4 FILLER_65_316 ();
 sg13g2_decap_4 FILLER_65_333 ();
 sg13g2_decap_4 FILLER_65_342 ();
 sg13g2_fill_1 FILLER_65_346 ();
 sg13g2_decap_8 FILLER_65_373 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_4 FILLER_65_421 ();
 sg13g2_fill_2 FILLER_65_425 ();
 sg13g2_decap_8 FILLER_65_430 ();
 sg13g2_decap_4 FILLER_65_437 ();
 sg13g2_decap_8 FILLER_65_444 ();
 sg13g2_decap_4 FILLER_65_451 ();
 sg13g2_fill_1 FILLER_65_464 ();
 sg13g2_decap_8 FILLER_65_473 ();
 sg13g2_decap_8 FILLER_65_480 ();
 sg13g2_decap_8 FILLER_65_487 ();
 sg13g2_fill_1 FILLER_65_500 ();
 sg13g2_decap_4 FILLER_65_510 ();
 sg13g2_fill_2 FILLER_65_514 ();
 sg13g2_decap_8 FILLER_65_519 ();
 sg13g2_fill_2 FILLER_65_526 ();
 sg13g2_fill_1 FILLER_65_528 ();
 sg13g2_fill_2 FILLER_65_537 ();
 sg13g2_fill_1 FILLER_65_539 ();
 sg13g2_decap_4 FILLER_65_556 ();
 sg13g2_fill_2 FILLER_65_560 ();
 sg13g2_fill_1 FILLER_65_565 ();
 sg13g2_fill_2 FILLER_65_592 ();
 sg13g2_fill_1 FILLER_65_594 ();
 sg13g2_fill_1 FILLER_65_599 ();
 sg13g2_decap_8 FILLER_65_605 ();
 sg13g2_fill_2 FILLER_65_612 ();
 sg13g2_fill_1 FILLER_65_614 ();
 sg13g2_decap_8 FILLER_65_642 ();
 sg13g2_decap_4 FILLER_65_649 ();
 sg13g2_fill_1 FILLER_65_653 ();
 sg13g2_decap_4 FILLER_65_659 ();
 sg13g2_fill_1 FILLER_65_663 ();
 sg13g2_fill_2 FILLER_65_676 ();
 sg13g2_fill_1 FILLER_65_678 ();
 sg13g2_decap_8 FILLER_65_695 ();
 sg13g2_fill_1 FILLER_65_702 ();
 sg13g2_decap_8 FILLER_65_707 ();
 sg13g2_fill_1 FILLER_65_714 ();
 sg13g2_decap_8 FILLER_65_742 ();
 sg13g2_fill_2 FILLER_65_760 ();
 sg13g2_fill_1 FILLER_65_762 ();
 sg13g2_decap_4 FILLER_65_772 ();
 sg13g2_fill_1 FILLER_65_776 ();
 sg13g2_fill_2 FILLER_65_784 ();
 sg13g2_fill_1 FILLER_65_786 ();
 sg13g2_fill_1 FILLER_65_805 ();
 sg13g2_decap_4 FILLER_65_814 ();
 sg13g2_fill_2 FILLER_65_828 ();
 sg13g2_decap_4 FILLER_65_835 ();
 sg13g2_fill_1 FILLER_65_839 ();
 sg13g2_fill_2 FILLER_65_849 ();
 sg13g2_fill_2 FILLER_65_868 ();
 sg13g2_fill_1 FILLER_65_870 ();
 sg13g2_fill_1 FILLER_65_874 ();
 sg13g2_fill_2 FILLER_65_881 ();
 sg13g2_fill_2 FILLER_65_896 ();
 sg13g2_decap_8 FILLER_65_908 ();
 sg13g2_decap_8 FILLER_65_915 ();
 sg13g2_fill_2 FILLER_65_922 ();
 sg13g2_fill_1 FILLER_65_924 ();
 sg13g2_fill_1 FILLER_65_931 ();
 sg13g2_fill_2 FILLER_65_941 ();
 sg13g2_fill_1 FILLER_65_966 ();
 sg13g2_fill_2 FILLER_65_973 ();
 sg13g2_decap_8 FILLER_65_984 ();
 sg13g2_fill_1 FILLER_65_991 ();
 sg13g2_fill_1 FILLER_65_1012 ();
 sg13g2_fill_2 FILLER_65_1018 ();
 sg13g2_fill_1 FILLER_65_1023 ();
 sg13g2_fill_2 FILLER_65_1033 ();
 sg13g2_fill_1 FILLER_65_1039 ();
 sg13g2_fill_2 FILLER_65_1062 ();
 sg13g2_fill_1 FILLER_65_1064 ();
 sg13g2_fill_1 FILLER_65_1071 ();
 sg13g2_fill_1 FILLER_65_1077 ();
 sg13g2_fill_1 FILLER_65_1085 ();
 sg13g2_fill_1 FILLER_65_1098 ();
 sg13g2_fill_1 FILLER_65_1132 ();
 sg13g2_fill_2 FILLER_65_1149 ();
 sg13g2_fill_1 FILLER_65_1151 ();
 sg13g2_fill_2 FILLER_65_1157 ();
 sg13g2_fill_1 FILLER_65_1159 ();
 sg13g2_fill_2 FILLER_65_1191 ();
 sg13g2_decap_8 FILLER_65_1208 ();
 sg13g2_decap_8 FILLER_65_1215 ();
 sg13g2_decap_4 FILLER_65_1222 ();
 sg13g2_fill_2 FILLER_65_1230 ();
 sg13g2_fill_1 FILLER_65_1232 ();
 sg13g2_fill_1 FILLER_65_1241 ();
 sg13g2_fill_2 FILLER_65_1248 ();
 sg13g2_fill_1 FILLER_65_1250 ();
 sg13g2_fill_2 FILLER_65_1261 ();
 sg13g2_fill_2 FILLER_65_1289 ();
 sg13g2_decap_4 FILLER_65_1321 ();
 sg13g2_fill_1 FILLER_65_1325 ();
 sg13g2_fill_2 FILLER_66_30 ();
 sg13g2_fill_1 FILLER_66_32 ();
 sg13g2_fill_2 FILLER_66_51 ();
 sg13g2_fill_1 FILLER_66_53 ();
 sg13g2_fill_1 FILLER_66_58 ();
 sg13g2_decap_4 FILLER_66_63 ();
 sg13g2_fill_1 FILLER_66_67 ();
 sg13g2_decap_8 FILLER_66_73 ();
 sg13g2_fill_2 FILLER_66_80 ();
 sg13g2_fill_1 FILLER_66_82 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_fill_1 FILLER_66_93 ();
 sg13g2_decap_4 FILLER_66_107 ();
 sg13g2_fill_1 FILLER_66_111 ();
 sg13g2_decap_4 FILLER_66_136 ();
 sg13g2_decap_4 FILLER_66_143 ();
 sg13g2_fill_2 FILLER_66_151 ();
 sg13g2_fill_2 FILLER_66_165 ();
 sg13g2_decap_4 FILLER_66_178 ();
 sg13g2_fill_2 FILLER_66_182 ();
 sg13g2_fill_1 FILLER_66_201 ();
 sg13g2_fill_1 FILLER_66_215 ();
 sg13g2_fill_1 FILLER_66_224 ();
 sg13g2_fill_1 FILLER_66_230 ();
 sg13g2_fill_1 FILLER_66_236 ();
 sg13g2_fill_1 FILLER_66_240 ();
 sg13g2_fill_1 FILLER_66_244 ();
 sg13g2_fill_2 FILLER_66_249 ();
 sg13g2_decap_4 FILLER_66_267 ();
 sg13g2_fill_1 FILLER_66_287 ();
 sg13g2_fill_1 FILLER_66_292 ();
 sg13g2_fill_1 FILLER_66_300 ();
 sg13g2_decap_8 FILLER_66_306 ();
 sg13g2_fill_2 FILLER_66_313 ();
 sg13g2_decap_8 FILLER_66_323 ();
 sg13g2_decap_8 FILLER_66_330 ();
 sg13g2_decap_4 FILLER_66_337 ();
 sg13g2_fill_2 FILLER_66_366 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_fill_2 FILLER_66_407 ();
 sg13g2_fill_2 FILLER_66_414 ();
 sg13g2_decap_8 FILLER_66_420 ();
 sg13g2_fill_1 FILLER_66_427 ();
 sg13g2_fill_2 FILLER_66_437 ();
 sg13g2_decap_8 FILLER_66_444 ();
 sg13g2_fill_1 FILLER_66_456 ();
 sg13g2_fill_1 FILLER_66_471 ();
 sg13g2_decap_8 FILLER_66_516 ();
 sg13g2_decap_4 FILLER_66_533 ();
 sg13g2_fill_2 FILLER_66_537 ();
 sg13g2_decap_8 FILLER_66_543 ();
 sg13g2_decap_8 FILLER_66_550 ();
 sg13g2_fill_2 FILLER_66_557 ();
 sg13g2_fill_1 FILLER_66_559 ();
 sg13g2_fill_2 FILLER_66_566 ();
 sg13g2_fill_2 FILLER_66_571 ();
 sg13g2_fill_1 FILLER_66_573 ();
 sg13g2_fill_2 FILLER_66_577 ();
 sg13g2_fill_1 FILLER_66_579 ();
 sg13g2_fill_2 FILLER_66_587 ();
 sg13g2_fill_1 FILLER_66_589 ();
 sg13g2_fill_2 FILLER_66_593 ();
 sg13g2_fill_1 FILLER_66_595 ();
 sg13g2_fill_2 FILLER_66_600 ();
 sg13g2_decap_8 FILLER_66_607 ();
 sg13g2_fill_2 FILLER_66_614 ();
 sg13g2_decap_8 FILLER_66_620 ();
 sg13g2_decap_4 FILLER_66_627 ();
 sg13g2_fill_1 FILLER_66_631 ();
 sg13g2_decap_4 FILLER_66_637 ();
 sg13g2_decap_4 FILLER_66_667 ();
 sg13g2_decap_4 FILLER_66_679 ();
 sg13g2_fill_1 FILLER_66_687 ();
 sg13g2_fill_1 FILLER_66_705 ();
 sg13g2_decap_8 FILLER_66_712 ();
 sg13g2_fill_1 FILLER_66_719 ();
 sg13g2_fill_1 FILLER_66_736 ();
 sg13g2_fill_1 FILLER_66_745 ();
 sg13g2_decap_8 FILLER_66_754 ();
 sg13g2_decap_4 FILLER_66_761 ();
 sg13g2_fill_2 FILLER_66_765 ();
 sg13g2_decap_8 FILLER_66_772 ();
 sg13g2_decap_8 FILLER_66_779 ();
 sg13g2_fill_1 FILLER_66_791 ();
 sg13g2_fill_2 FILLER_66_805 ();
 sg13g2_fill_2 FILLER_66_812 ();
 sg13g2_fill_1 FILLER_66_823 ();
 sg13g2_fill_1 FILLER_66_828 ();
 sg13g2_fill_2 FILLER_66_832 ();
 sg13g2_fill_2 FILLER_66_849 ();
 sg13g2_fill_1 FILLER_66_864 ();
 sg13g2_fill_2 FILLER_66_869 ();
 sg13g2_decap_8 FILLER_66_876 ();
 sg13g2_fill_2 FILLER_66_883 ();
 sg13g2_decap_4 FILLER_66_890 ();
 sg13g2_fill_1 FILLER_66_894 ();
 sg13g2_decap_8 FILLER_66_903 ();
 sg13g2_decap_8 FILLER_66_910 ();
 sg13g2_fill_2 FILLER_66_917 ();
 sg13g2_fill_2 FILLER_66_952 ();
 sg13g2_fill_2 FILLER_66_961 ();
 sg13g2_fill_1 FILLER_66_974 ();
 sg13g2_decap_8 FILLER_66_979 ();
 sg13g2_fill_2 FILLER_66_1046 ();
 sg13g2_fill_2 FILLER_66_1052 ();
 sg13g2_fill_1 FILLER_66_1054 ();
 sg13g2_fill_1 FILLER_66_1069 ();
 sg13g2_fill_1 FILLER_66_1085 ();
 sg13g2_fill_1 FILLER_66_1090 ();
 sg13g2_fill_1 FILLER_66_1095 ();
 sg13g2_fill_1 FILLER_66_1101 ();
 sg13g2_fill_2 FILLER_66_1106 ();
 sg13g2_fill_1 FILLER_66_1112 ();
 sg13g2_fill_2 FILLER_66_1121 ();
 sg13g2_fill_2 FILLER_66_1127 ();
 sg13g2_fill_2 FILLER_66_1154 ();
 sg13g2_fill_1 FILLER_66_1187 ();
 sg13g2_fill_1 FILLER_66_1194 ();
 sg13g2_fill_1 FILLER_66_1205 ();
 sg13g2_decap_8 FILLER_66_1232 ();
 sg13g2_decap_8 FILLER_66_1239 ();
 sg13g2_fill_1 FILLER_66_1246 ();
 sg13g2_fill_1 FILLER_66_1252 ();
 sg13g2_fill_2 FILLER_66_1264 ();
 sg13g2_fill_2 FILLER_66_1270 ();
 sg13g2_fill_1 FILLER_66_1272 ();
 sg13g2_decap_8 FILLER_66_1288 ();
 sg13g2_decap_8 FILLER_66_1304 ();
 sg13g2_decap_8 FILLER_66_1311 ();
 sg13g2_decap_8 FILLER_66_1318 ();
 sg13g2_fill_1 FILLER_66_1325 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_41 ();
 sg13g2_fill_1 FILLER_67_68 ();
 sg13g2_decap_4 FILLER_67_74 ();
 sg13g2_decap_8 FILLER_67_104 ();
 sg13g2_decap_8 FILLER_67_116 ();
 sg13g2_decap_8 FILLER_67_123 ();
 sg13g2_decap_8 FILLER_67_130 ();
 sg13g2_fill_1 FILLER_67_140 ();
 sg13g2_fill_2 FILLER_67_144 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_decap_8 FILLER_67_172 ();
 sg13g2_decap_4 FILLER_67_179 ();
 sg13g2_decap_8 FILLER_67_213 ();
 sg13g2_decap_4 FILLER_67_225 ();
 sg13g2_fill_1 FILLER_67_229 ();
 sg13g2_fill_1 FILLER_67_243 ();
 sg13g2_decap_4 FILLER_67_252 ();
 sg13g2_fill_2 FILLER_67_256 ();
 sg13g2_fill_2 FILLER_67_263 ();
 sg13g2_fill_2 FILLER_67_279 ();
 sg13g2_fill_1 FILLER_67_285 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_fill_1 FILLER_67_301 ();
 sg13g2_decap_4 FILLER_67_306 ();
 sg13g2_decap_8 FILLER_67_315 ();
 sg13g2_fill_1 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_332 ();
 sg13g2_decap_4 FILLER_67_339 ();
 sg13g2_decap_8 FILLER_67_349 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_fill_1 FILLER_67_363 ();
 sg13g2_fill_1 FILLER_67_368 ();
 sg13g2_fill_1 FILLER_67_410 ();
 sg13g2_decap_8 FILLER_67_418 ();
 sg13g2_fill_1 FILLER_67_425 ();
 sg13g2_decap_8 FILLER_67_443 ();
 sg13g2_decap_4 FILLER_67_450 ();
 sg13g2_fill_1 FILLER_67_454 ();
 sg13g2_fill_2 FILLER_67_459 ();
 sg13g2_fill_1 FILLER_67_473 ();
 sg13g2_decap_4 FILLER_67_486 ();
 sg13g2_fill_1 FILLER_67_495 ();
 sg13g2_fill_1 FILLER_67_500 ();
 sg13g2_fill_2 FILLER_67_506 ();
 sg13g2_fill_2 FILLER_67_517 ();
 sg13g2_fill_1 FILLER_67_519 ();
 sg13g2_decap_4 FILLER_67_525 ();
 sg13g2_fill_2 FILLER_67_540 ();
 sg13g2_fill_1 FILLER_67_542 ();
 sg13g2_decap_8 FILLER_67_546 ();
 sg13g2_decap_8 FILLER_67_553 ();
 sg13g2_fill_2 FILLER_67_560 ();
 sg13g2_fill_1 FILLER_67_562 ();
 sg13g2_fill_2 FILLER_67_576 ();
 sg13g2_fill_1 FILLER_67_578 ();
 sg13g2_fill_1 FILLER_67_583 ();
 sg13g2_decap_8 FILLER_67_608 ();
 sg13g2_fill_2 FILLER_67_615 ();
 sg13g2_fill_1 FILLER_67_617 ();
 sg13g2_decap_4 FILLER_67_621 ();
 sg13g2_fill_2 FILLER_67_665 ();
 sg13g2_fill_1 FILLER_67_670 ();
 sg13g2_decap_8 FILLER_67_678 ();
 sg13g2_decap_8 FILLER_67_685 ();
 sg13g2_decap_4 FILLER_67_692 ();
 sg13g2_fill_1 FILLER_67_696 ();
 sg13g2_fill_2 FILLER_67_709 ();
 sg13g2_fill_1 FILLER_67_715 ();
 sg13g2_fill_2 FILLER_67_755 ();
 sg13g2_fill_1 FILLER_67_761 ();
 sg13g2_fill_1 FILLER_67_772 ();
 sg13g2_fill_2 FILLER_67_778 ();
 sg13g2_decap_4 FILLER_67_784 ();
 sg13g2_fill_2 FILLER_67_797 ();
 sg13g2_fill_1 FILLER_67_799 ();
 sg13g2_fill_1 FILLER_67_813 ();
 sg13g2_fill_2 FILLER_67_834 ();
 sg13g2_fill_2 FILLER_67_844 ();
 sg13g2_fill_2 FILLER_67_852 ();
 sg13g2_fill_2 FILLER_67_898 ();
 sg13g2_fill_1 FILLER_67_910 ();
 sg13g2_fill_2 FILLER_67_924 ();
 sg13g2_fill_1 FILLER_67_934 ();
 sg13g2_fill_2 FILLER_67_997 ();
 sg13g2_fill_2 FILLER_67_1007 ();
 sg13g2_fill_2 FILLER_67_1022 ();
 sg13g2_fill_1 FILLER_67_1040 ();
 sg13g2_fill_2 FILLER_67_1069 ();
 sg13g2_fill_1 FILLER_67_1083 ();
 sg13g2_fill_2 FILLER_67_1099 ();
 sg13g2_fill_2 FILLER_67_1106 ();
 sg13g2_fill_1 FILLER_67_1135 ();
 sg13g2_fill_1 FILLER_67_1150 ();
 sg13g2_fill_1 FILLER_67_1169 ();
 sg13g2_fill_1 FILLER_67_1178 ();
 sg13g2_fill_1 FILLER_67_1185 ();
 sg13g2_decap_8 FILLER_67_1214 ();
 sg13g2_decap_4 FILLER_67_1221 ();
 sg13g2_fill_2 FILLER_67_1225 ();
 sg13g2_decap_8 FILLER_67_1236 ();
 sg13g2_decap_4 FILLER_67_1243 ();
 sg13g2_fill_1 FILLER_67_1247 ();
 sg13g2_fill_1 FILLER_67_1256 ();
 sg13g2_decap_4 FILLER_67_1266 ();
 sg13g2_fill_1 FILLER_67_1270 ();
 sg13g2_decap_8 FILLER_67_1313 ();
 sg13g2_decap_4 FILLER_67_1320 ();
 sg13g2_fill_2 FILLER_67_1324 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_4 FILLER_68_21 ();
 sg13g2_fill_2 FILLER_68_25 ();
 sg13g2_decap_4 FILLER_68_31 ();
 sg13g2_fill_1 FILLER_68_35 ();
 sg13g2_decap_4 FILLER_68_79 ();
 sg13g2_fill_2 FILLER_68_83 ();
 sg13g2_decap_8 FILLER_68_89 ();
 sg13g2_decap_8 FILLER_68_96 ();
 sg13g2_decap_8 FILLER_68_129 ();
 sg13g2_fill_2 FILLER_68_136 ();
 sg13g2_fill_1 FILLER_68_141 ();
 sg13g2_decap_4 FILLER_68_158 ();
 sg13g2_fill_1 FILLER_68_162 ();
 sg13g2_decap_8 FILLER_68_172 ();
 sg13g2_decap_8 FILLER_68_179 ();
 sg13g2_decap_8 FILLER_68_186 ();
 sg13g2_decap_8 FILLER_68_193 ();
 sg13g2_decap_8 FILLER_68_200 ();
 sg13g2_decap_4 FILLER_68_207 ();
 sg13g2_fill_2 FILLER_68_211 ();
 sg13g2_fill_1 FILLER_68_217 ();
 sg13g2_fill_1 FILLER_68_263 ();
 sg13g2_fill_2 FILLER_68_284 ();
 sg13g2_fill_1 FILLER_68_286 ();
 sg13g2_fill_1 FILLER_68_295 ();
 sg13g2_fill_1 FILLER_68_299 ();
 sg13g2_fill_2 FILLER_68_308 ();
 sg13g2_decap_4 FILLER_68_315 ();
 sg13g2_decap_4 FILLER_68_322 ();
 sg13g2_fill_2 FILLER_68_373 ();
 sg13g2_fill_1 FILLER_68_386 ();
 sg13g2_fill_2 FILLER_68_394 ();
 sg13g2_decap_8 FILLER_68_413 ();
 sg13g2_decap_8 FILLER_68_420 ();
 sg13g2_decap_4 FILLER_68_427 ();
 sg13g2_fill_1 FILLER_68_446 ();
 sg13g2_fill_1 FILLER_68_451 ();
 sg13g2_fill_1 FILLER_68_459 ();
 sg13g2_decap_8 FILLER_68_465 ();
 sg13g2_fill_2 FILLER_68_472 ();
 sg13g2_fill_1 FILLER_68_474 ();
 sg13g2_decap_4 FILLER_68_479 ();
 sg13g2_decap_8 FILLER_68_488 ();
 sg13g2_fill_2 FILLER_68_495 ();
 sg13g2_fill_1 FILLER_68_497 ();
 sg13g2_fill_2 FILLER_68_506 ();
 sg13g2_fill_1 FILLER_68_508 ();
 sg13g2_fill_2 FILLER_68_513 ();
 sg13g2_fill_1 FILLER_68_520 ();
 sg13g2_fill_1 FILLER_68_525 ();
 sg13g2_fill_2 FILLER_68_530 ();
 sg13g2_fill_1 FILLER_68_541 ();
 sg13g2_decap_8 FILLER_68_550 ();
 sg13g2_decap_4 FILLER_68_557 ();
 sg13g2_fill_1 FILLER_68_572 ();
 sg13g2_fill_2 FILLER_68_577 ();
 sg13g2_fill_1 FILLER_68_582 ();
 sg13g2_fill_1 FILLER_68_589 ();
 sg13g2_fill_2 FILLER_68_594 ();
 sg13g2_fill_2 FILLER_68_601 ();
 sg13g2_fill_2 FILLER_68_608 ();
 sg13g2_fill_1 FILLER_68_610 ();
 sg13g2_fill_1 FILLER_68_622 ();
 sg13g2_fill_2 FILLER_68_628 ();
 sg13g2_fill_1 FILLER_68_630 ();
 sg13g2_decap_4 FILLER_68_645 ();
 sg13g2_fill_2 FILLER_68_649 ();
 sg13g2_fill_1 FILLER_68_655 ();
 sg13g2_fill_1 FILLER_68_674 ();
 sg13g2_fill_1 FILLER_68_687 ();
 sg13g2_fill_2 FILLER_68_702 ();
 sg13g2_fill_1 FILLER_68_741 ();
 sg13g2_fill_1 FILLER_68_747 ();
 sg13g2_fill_2 FILLER_68_760 ();
 sg13g2_fill_1 FILLER_68_762 ();
 sg13g2_decap_8 FILLER_68_773 ();
 sg13g2_fill_2 FILLER_68_796 ();
 sg13g2_fill_2 FILLER_68_823 ();
 sg13g2_fill_1 FILLER_68_841 ();
 sg13g2_fill_1 FILLER_68_847 ();
 sg13g2_fill_2 FILLER_68_858 ();
 sg13g2_decap_4 FILLER_68_881 ();
 sg13g2_decap_8 FILLER_68_889 ();
 sg13g2_decap_8 FILLER_68_896 ();
 sg13g2_fill_1 FILLER_68_903 ();
 sg13g2_fill_1 FILLER_68_912 ();
 sg13g2_fill_1 FILLER_68_932 ();
 sg13g2_fill_2 FILLER_68_975 ();
 sg13g2_fill_1 FILLER_68_977 ();
 sg13g2_fill_2 FILLER_68_983 ();
 sg13g2_fill_2 FILLER_68_1003 ();
 sg13g2_fill_2 FILLER_68_1014 ();
 sg13g2_fill_2 FILLER_68_1019 ();
 sg13g2_fill_1 FILLER_68_1029 ();
 sg13g2_fill_2 FILLER_68_1044 ();
 sg13g2_fill_2 FILLER_68_1059 ();
 sg13g2_fill_1 FILLER_68_1065 ();
 sg13g2_fill_2 FILLER_68_1077 ();
 sg13g2_fill_1 FILLER_68_1093 ();
 sg13g2_fill_2 FILLER_68_1114 ();
 sg13g2_fill_1 FILLER_68_1131 ();
 sg13g2_fill_1 FILLER_68_1136 ();
 sg13g2_fill_1 FILLER_68_1152 ();
 sg13g2_fill_1 FILLER_68_1159 ();
 sg13g2_fill_2 FILLER_68_1165 ();
 sg13g2_fill_2 FILLER_68_1180 ();
 sg13g2_fill_2 FILLER_68_1196 ();
 sg13g2_fill_1 FILLER_68_1209 ();
 sg13g2_fill_2 FILLER_68_1219 ();
 sg13g2_fill_1 FILLER_68_1221 ();
 sg13g2_fill_2 FILLER_68_1226 ();
 sg13g2_decap_8 FILLER_68_1232 ();
 sg13g2_decap_8 FILLER_68_1239 ();
 sg13g2_fill_2 FILLER_68_1246 ();
 sg13g2_fill_2 FILLER_68_1260 ();
 sg13g2_fill_1 FILLER_68_1262 ();
 sg13g2_decap_8 FILLER_68_1267 ();
 sg13g2_decap_4 FILLER_68_1274 ();
 sg13g2_fill_1 FILLER_68_1283 ();
 sg13g2_fill_2 FILLER_68_1288 ();
 sg13g2_fill_1 FILLER_68_1290 ();
 sg13g2_fill_1 FILLER_68_1296 ();
 sg13g2_decap_8 FILLER_68_1302 ();
 sg13g2_decap_8 FILLER_68_1309 ();
 sg13g2_decap_8 FILLER_68_1316 ();
 sg13g2_fill_2 FILLER_68_1323 ();
 sg13g2_fill_1 FILLER_68_1325 ();
 sg13g2_decap_8 FILLER_69_47 ();
 sg13g2_decap_8 FILLER_69_54 ();
 sg13g2_fill_2 FILLER_69_61 ();
 sg13g2_fill_1 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_67 ();
 sg13g2_fill_1 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_110 ();
 sg13g2_fill_1 FILLER_69_117 ();
 sg13g2_decap_4 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_127 ();
 sg13g2_fill_2 FILLER_69_138 ();
 sg13g2_fill_2 FILLER_69_157 ();
 sg13g2_decap_8 FILLER_69_177 ();
 sg13g2_decap_4 FILLER_69_188 ();
 sg13g2_fill_1 FILLER_69_192 ();
 sg13g2_fill_1 FILLER_69_201 ();
 sg13g2_decap_4 FILLER_69_207 ();
 sg13g2_fill_2 FILLER_69_211 ();
 sg13g2_decap_4 FILLER_69_221 ();
 sg13g2_decap_8 FILLER_69_240 ();
 sg13g2_fill_2 FILLER_69_247 ();
 sg13g2_fill_1 FILLER_69_254 ();
 sg13g2_fill_1 FILLER_69_260 ();
 sg13g2_fill_2 FILLER_69_281 ();
 sg13g2_fill_1 FILLER_69_283 ();
 sg13g2_fill_1 FILLER_69_293 ();
 sg13g2_decap_4 FILLER_69_306 ();
 sg13g2_fill_1 FILLER_69_310 ();
 sg13g2_decap_8 FILLER_69_330 ();
 sg13g2_fill_1 FILLER_69_337 ();
 sg13g2_decap_8 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_350 ();
 sg13g2_decap_8 FILLER_69_357 ();
 sg13g2_decap_4 FILLER_69_364 ();
 sg13g2_fill_2 FILLER_69_368 ();
 sg13g2_fill_1 FILLER_69_381 ();
 sg13g2_fill_1 FILLER_69_390 ();
 sg13g2_fill_1 FILLER_69_415 ();
 sg13g2_fill_2 FILLER_69_425 ();
 sg13g2_fill_1 FILLER_69_427 ();
 sg13g2_fill_1 FILLER_69_433 ();
 sg13g2_fill_2 FILLER_69_441 ();
 sg13g2_fill_1 FILLER_69_448 ();
 sg13g2_fill_1 FILLER_69_453 ();
 sg13g2_decap_8 FILLER_69_459 ();
 sg13g2_decap_8 FILLER_69_466 ();
 sg13g2_decap_8 FILLER_69_473 ();
 sg13g2_decap_4 FILLER_69_480 ();
 sg13g2_decap_8 FILLER_69_489 ();
 sg13g2_decap_8 FILLER_69_496 ();
 sg13g2_fill_2 FILLER_69_503 ();
 sg13g2_fill_2 FILLER_69_536 ();
 sg13g2_fill_1 FILLER_69_538 ();
 sg13g2_fill_1 FILLER_69_544 ();
 sg13g2_fill_2 FILLER_69_550 ();
 sg13g2_fill_2 FILLER_69_556 ();
 sg13g2_fill_2 FILLER_69_563 ();
 sg13g2_fill_1 FILLER_69_565 ();
 sg13g2_fill_1 FILLER_69_588 ();
 sg13g2_fill_2 FILLER_69_604 ();
 sg13g2_decap_4 FILLER_69_610 ();
 sg13g2_fill_1 FILLER_69_618 ();
 sg13g2_decap_4 FILLER_69_624 ();
 sg13g2_fill_2 FILLER_69_643 ();
 sg13g2_fill_2 FILLER_69_650 ();
 sg13g2_fill_1 FILLER_69_652 ();
 sg13g2_fill_2 FILLER_69_668 ();
 sg13g2_fill_1 FILLER_69_670 ();
 sg13g2_fill_1 FILLER_69_678 ();
 sg13g2_fill_1 FILLER_69_712 ();
 sg13g2_fill_1 FILLER_69_733 ();
 sg13g2_fill_1 FILLER_69_746 ();
 sg13g2_fill_1 FILLER_69_752 ();
 sg13g2_fill_2 FILLER_69_771 ();
 sg13g2_fill_1 FILLER_69_773 ();
 sg13g2_decap_8 FILLER_69_777 ();
 sg13g2_decap_4 FILLER_69_784 ();
 sg13g2_fill_1 FILLER_69_788 ();
 sg13g2_fill_2 FILLER_69_803 ();
 sg13g2_fill_2 FILLER_69_822 ();
 sg13g2_fill_1 FILLER_69_849 ();
 sg13g2_fill_2 FILLER_69_874 ();
 sg13g2_fill_1 FILLER_69_881 ();
 sg13g2_fill_1 FILLER_69_887 ();
 sg13g2_fill_2 FILLER_69_892 ();
 sg13g2_decap_8 FILLER_69_898 ();
 sg13g2_decap_4 FILLER_69_909 ();
 sg13g2_fill_2 FILLER_69_925 ();
 sg13g2_fill_2 FILLER_69_942 ();
 sg13g2_fill_1 FILLER_69_982 ();
 sg13g2_fill_2 FILLER_69_994 ();
 sg13g2_fill_1 FILLER_69_1010 ();
 sg13g2_fill_1 FILLER_69_1042 ();
 sg13g2_decap_8 FILLER_69_1062 ();
 sg13g2_fill_1 FILLER_69_1069 ();
 sg13g2_decap_4 FILLER_69_1100 ();
 sg13g2_fill_1 FILLER_69_1108 ();
 sg13g2_fill_1 FILLER_69_1119 ();
 sg13g2_decap_8 FILLER_69_1123 ();
 sg13g2_decap_4 FILLER_69_1130 ();
 sg13g2_fill_2 FILLER_69_1134 ();
 sg13g2_fill_1 FILLER_69_1152 ();
 sg13g2_fill_1 FILLER_69_1202 ();
 sg13g2_fill_1 FILLER_69_1208 ();
 sg13g2_fill_1 FILLER_69_1215 ();
 sg13g2_fill_1 FILLER_69_1223 ();
 sg13g2_decap_8 FILLER_69_1228 ();
 sg13g2_decap_8 FILLER_69_1235 ();
 sg13g2_decap_4 FILLER_69_1242 ();
 sg13g2_fill_1 FILLER_69_1250 ();
 sg13g2_decap_4 FILLER_69_1268 ();
 sg13g2_fill_1 FILLER_69_1272 ();
 sg13g2_fill_1 FILLER_69_1278 ();
 sg13g2_decap_8 FILLER_69_1305 ();
 sg13g2_decap_8 FILLER_69_1312 ();
 sg13g2_decap_8 FILLER_69_1319 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_4 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_25 ();
 sg13g2_decap_8 FILLER_70_32 ();
 sg13g2_decap_4 FILLER_70_39 ();
 sg13g2_fill_1 FILLER_70_62 ();
 sg13g2_decap_4 FILLER_70_71 ();
 sg13g2_fill_2 FILLER_70_75 ();
 sg13g2_decap_8 FILLER_70_80 ();
 sg13g2_decap_8 FILLER_70_87 ();
 sg13g2_decap_8 FILLER_70_94 ();
 sg13g2_decap_8 FILLER_70_101 ();
 sg13g2_decap_8 FILLER_70_108 ();
 sg13g2_fill_2 FILLER_70_115 ();
 sg13g2_decap_8 FILLER_70_121 ();
 sg13g2_decap_4 FILLER_70_128 ();
 sg13g2_fill_2 FILLER_70_132 ();
 sg13g2_fill_2 FILLER_70_154 ();
 sg13g2_fill_1 FILLER_70_156 ();
 sg13g2_fill_1 FILLER_70_161 ();
 sg13g2_fill_2 FILLER_70_165 ();
 sg13g2_decap_8 FILLER_70_172 ();
 sg13g2_fill_2 FILLER_70_179 ();
 sg13g2_fill_2 FILLER_70_201 ();
 sg13g2_decap_4 FILLER_70_206 ();
 sg13g2_fill_1 FILLER_70_210 ();
 sg13g2_decap_4 FILLER_70_216 ();
 sg13g2_fill_2 FILLER_70_220 ();
 sg13g2_fill_1 FILLER_70_232 ();
 sg13g2_decap_8 FILLER_70_262 ();
 sg13g2_fill_2 FILLER_70_269 ();
 sg13g2_decap_4 FILLER_70_274 ();
 sg13g2_fill_2 FILLER_70_288 ();
 sg13g2_fill_1 FILLER_70_290 ();
 sg13g2_decap_4 FILLER_70_296 ();
 sg13g2_fill_1 FILLER_70_300 ();
 sg13g2_decap_4 FILLER_70_305 ();
 sg13g2_fill_1 FILLER_70_309 ();
 sg13g2_fill_2 FILLER_70_315 ();
 sg13g2_fill_1 FILLER_70_317 ();
 sg13g2_decap_8 FILLER_70_321 ();
 sg13g2_decap_4 FILLER_70_328 ();
 sg13g2_fill_2 FILLER_70_335 ();
 sg13g2_decap_8 FILLER_70_357 ();
 sg13g2_fill_2 FILLER_70_372 ();
 sg13g2_decap_4 FILLER_70_404 ();
 sg13g2_fill_2 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_70_419 ();
 sg13g2_fill_2 FILLER_70_426 ();
 sg13g2_fill_2 FILLER_70_432 ();
 sg13g2_fill_1 FILLER_70_434 ();
 sg13g2_fill_1 FILLER_70_484 ();
 sg13g2_decap_4 FILLER_70_489 ();
 sg13g2_fill_2 FILLER_70_493 ();
 sg13g2_fill_2 FILLER_70_500 ();
 sg13g2_fill_2 FILLER_70_510 ();
 sg13g2_decap_8 FILLER_70_533 ();
 sg13g2_decap_4 FILLER_70_540 ();
 sg13g2_fill_2 FILLER_70_547 ();
 sg13g2_fill_1 FILLER_70_549 ();
 sg13g2_fill_1 FILLER_70_555 ();
 sg13g2_decap_4 FILLER_70_560 ();
 sg13g2_fill_2 FILLER_70_564 ();
 sg13g2_decap_8 FILLER_70_596 ();
 sg13g2_decap_8 FILLER_70_603 ();
 sg13g2_decap_8 FILLER_70_610 ();
 sg13g2_fill_2 FILLER_70_624 ();
 sg13g2_fill_1 FILLER_70_626 ();
 sg13g2_decap_4 FILLER_70_636 ();
 sg13g2_fill_1 FILLER_70_640 ();
 sg13g2_fill_2 FILLER_70_646 ();
 sg13g2_fill_1 FILLER_70_648 ();
 sg13g2_decap_8 FILLER_70_653 ();
 sg13g2_decap_8 FILLER_70_660 ();
 sg13g2_decap_4 FILLER_70_667 ();
 sg13g2_fill_2 FILLER_70_671 ();
 sg13g2_decap_8 FILLER_70_680 ();
 sg13g2_fill_1 FILLER_70_687 ();
 sg13g2_decap_8 FILLER_70_692 ();
 sg13g2_decap_4 FILLER_70_699 ();
 sg13g2_fill_2 FILLER_70_703 ();
 sg13g2_fill_1 FILLER_70_711 ();
 sg13g2_fill_1 FILLER_70_715 ();
 sg13g2_fill_1 FILLER_70_722 ();
 sg13g2_fill_1 FILLER_70_729 ();
 sg13g2_fill_2 FILLER_70_734 ();
 sg13g2_fill_2 FILLER_70_744 ();
 sg13g2_fill_1 FILLER_70_746 ();
 sg13g2_fill_1 FILLER_70_758 ();
 sg13g2_decap_8 FILLER_70_764 ();
 sg13g2_decap_8 FILLER_70_771 ();
 sg13g2_decap_8 FILLER_70_778 ();
 sg13g2_fill_2 FILLER_70_785 ();
 sg13g2_fill_1 FILLER_70_787 ();
 sg13g2_decap_4 FILLER_70_801 ();
 sg13g2_fill_1 FILLER_70_818 ();
 sg13g2_decap_4 FILLER_70_830 ();
 sg13g2_fill_2 FILLER_70_839 ();
 sg13g2_fill_1 FILLER_70_845 ();
 sg13g2_decap_8 FILLER_70_850 ();
 sg13g2_decap_8 FILLER_70_857 ();
 sg13g2_decap_4 FILLER_70_864 ();
 sg13g2_fill_2 FILLER_70_868 ();
 sg13g2_decap_8 FILLER_70_874 ();
 sg13g2_decap_8 FILLER_70_881 ();
 sg13g2_fill_2 FILLER_70_893 ();
 sg13g2_fill_1 FILLER_70_917 ();
 sg13g2_fill_2 FILLER_70_935 ();
 sg13g2_fill_1 FILLER_70_943 ();
 sg13g2_fill_2 FILLER_70_954 ();
 sg13g2_fill_2 FILLER_70_971 ();
 sg13g2_fill_1 FILLER_70_983 ();
 sg13g2_fill_1 FILLER_70_1018 ();
 sg13g2_fill_2 FILLER_70_1026 ();
 sg13g2_decap_8 FILLER_70_1063 ();
 sg13g2_fill_2 FILLER_70_1070 ();
 sg13g2_fill_1 FILLER_70_1072 ();
 sg13g2_decap_4 FILLER_70_1088 ();
 sg13g2_decap_8 FILLER_70_1102 ();
 sg13g2_decap_8 FILLER_70_1117 ();
 sg13g2_decap_4 FILLER_70_1124 ();
 sg13g2_fill_2 FILLER_70_1132 ();
 sg13g2_fill_1 FILLER_70_1134 ();
 sg13g2_fill_2 FILLER_70_1144 ();
 sg13g2_fill_2 FILLER_70_1161 ();
 sg13g2_fill_2 FILLER_70_1187 ();
 sg13g2_decap_4 FILLER_70_1205 ();
 sg13g2_fill_1 FILLER_70_1209 ();
 sg13g2_fill_2 FILLER_70_1214 ();
 sg13g2_fill_2 FILLER_70_1220 ();
 sg13g2_fill_1 FILLER_70_1222 ();
 sg13g2_fill_1 FILLER_70_1227 ();
 sg13g2_fill_1 FILLER_70_1235 ();
 sg13g2_fill_1 FILLER_70_1244 ();
 sg13g2_fill_1 FILLER_70_1254 ();
 sg13g2_decap_4 FILLER_70_1259 ();
 sg13g2_fill_2 FILLER_70_1272 ();
 sg13g2_fill_1 FILLER_70_1274 ();
 sg13g2_decap_8 FILLER_70_1279 ();
 sg13g2_decap_8 FILLER_70_1286 ();
 sg13g2_decap_8 FILLER_70_1293 ();
 sg13g2_decap_8 FILLER_70_1300 ();
 sg13g2_decap_8 FILLER_70_1307 ();
 sg13g2_decap_8 FILLER_70_1314 ();
 sg13g2_decap_4 FILLER_70_1321 ();
 sg13g2_fill_1 FILLER_70_1325 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_2 FILLER_71_29 ();
 sg13g2_fill_1 FILLER_71_31 ();
 sg13g2_decap_8 FILLER_71_36 ();
 sg13g2_decap_4 FILLER_71_43 ();
 sg13g2_decap_4 FILLER_71_64 ();
 sg13g2_fill_1 FILLER_71_74 ();
 sg13g2_decap_8 FILLER_71_83 ();
 sg13g2_fill_2 FILLER_71_90 ();
 sg13g2_fill_2 FILLER_71_101 ();
 sg13g2_fill_2 FILLER_71_117 ();
 sg13g2_fill_1 FILLER_71_119 ();
 sg13g2_decap_4 FILLER_71_125 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_fill_2 FILLER_71_140 ();
 sg13g2_decap_4 FILLER_71_151 ();
 sg13g2_fill_1 FILLER_71_170 ();
 sg13g2_decap_4 FILLER_71_181 ();
 sg13g2_fill_2 FILLER_71_200 ();
 sg13g2_fill_1 FILLER_71_202 ();
 sg13g2_fill_2 FILLER_71_207 ();
 sg13g2_decap_8 FILLER_71_214 ();
 sg13g2_decap_4 FILLER_71_221 ();
 sg13g2_fill_2 FILLER_71_228 ();
 sg13g2_fill_1 FILLER_71_230 ();
 sg13g2_fill_2 FILLER_71_235 ();
 sg13g2_fill_1 FILLER_71_237 ();
 sg13g2_decap_4 FILLER_71_251 ();
 sg13g2_fill_1 FILLER_71_255 ();
 sg13g2_decap_4 FILLER_71_259 ();
 sg13g2_fill_2 FILLER_71_272 ();
 sg13g2_fill_1 FILLER_71_274 ();
 sg13g2_decap_4 FILLER_71_278 ();
 sg13g2_fill_1 FILLER_71_282 ();
 sg13g2_fill_1 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_307 ();
 sg13g2_fill_2 FILLER_71_314 ();
 sg13g2_decap_4 FILLER_71_319 ();
 sg13g2_fill_1 FILLER_71_323 ();
 sg13g2_fill_1 FILLER_71_341 ();
 sg13g2_decap_8 FILLER_71_355 ();
 sg13g2_decap_8 FILLER_71_362 ();
 sg13g2_fill_2 FILLER_71_395 ();
 sg13g2_fill_2 FILLER_71_406 ();
 sg13g2_decap_8 FILLER_71_416 ();
 sg13g2_decap_8 FILLER_71_458 ();
 sg13g2_decap_8 FILLER_71_465 ();
 sg13g2_fill_2 FILLER_71_472 ();
 sg13g2_decap_8 FILLER_71_484 ();
 sg13g2_decap_4 FILLER_71_491 ();
 sg13g2_fill_1 FILLER_71_495 ();
 sg13g2_fill_2 FILLER_71_508 ();
 sg13g2_fill_2 FILLER_71_528 ();
 sg13g2_fill_2 FILLER_71_534 ();
 sg13g2_fill_1 FILLER_71_536 ();
 sg13g2_decap_8 FILLER_71_541 ();
 sg13g2_fill_2 FILLER_71_548 ();
 sg13g2_fill_1 FILLER_71_550 ();
 sg13g2_decap_8 FILLER_71_585 ();
 sg13g2_decap_8 FILLER_71_592 ();
 sg13g2_fill_1 FILLER_71_611 ();
 sg13g2_fill_1 FILLER_71_629 ();
 sg13g2_decap_4 FILLER_71_634 ();
 sg13g2_decap_8 FILLER_71_659 ();
 sg13g2_fill_1 FILLER_71_666 ();
 sg13g2_fill_1 FILLER_71_690 ();
 sg13g2_fill_2 FILLER_71_695 ();
 sg13g2_fill_2 FILLER_71_700 ();
 sg13g2_decap_4 FILLER_71_718 ();
 sg13g2_fill_2 FILLER_71_725 ();
 sg13g2_fill_2 FILLER_71_735 ();
 sg13g2_fill_1 FILLER_71_741 ();
 sg13g2_fill_2 FILLER_71_746 ();
 sg13g2_fill_1 FILLER_71_752 ();
 sg13g2_fill_2 FILLER_71_765 ();
 sg13g2_fill_1 FILLER_71_767 ();
 sg13g2_decap_8 FILLER_71_794 ();
 sg13g2_decap_8 FILLER_71_801 ();
 sg13g2_decap_4 FILLER_71_808 ();
 sg13g2_fill_2 FILLER_71_812 ();
 sg13g2_decap_4 FILLER_71_817 ();
 sg13g2_decap_4 FILLER_71_830 ();
 sg13g2_fill_1 FILLER_71_843 ();
 sg13g2_decap_4 FILLER_71_849 ();
 sg13g2_decap_4 FILLER_71_884 ();
 sg13g2_fill_1 FILLER_71_888 ();
 sg13g2_fill_2 FILLER_71_900 ();
 sg13g2_fill_1 FILLER_71_902 ();
 sg13g2_fill_2 FILLER_71_915 ();
 sg13g2_fill_2 FILLER_71_925 ();
 sg13g2_fill_1 FILLER_71_940 ();
 sg13g2_fill_1 FILLER_71_960 ();
 sg13g2_fill_2 FILLER_71_966 ();
 sg13g2_fill_2 FILLER_71_973 ();
 sg13g2_fill_2 FILLER_71_980 ();
 sg13g2_decap_8 FILLER_71_986 ();
 sg13g2_fill_2 FILLER_71_993 ();
 sg13g2_fill_2 FILLER_71_998 ();
 sg13g2_fill_1 FILLER_71_1000 ();
 sg13g2_fill_1 FILLER_71_1041 ();
 sg13g2_decap_8 FILLER_71_1055 ();
 sg13g2_fill_1 FILLER_71_1070 ();
 sg13g2_decap_8 FILLER_71_1074 ();
 sg13g2_fill_2 FILLER_71_1086 ();
 sg13g2_decap_8 FILLER_71_1102 ();
 sg13g2_fill_2 FILLER_71_1109 ();
 sg13g2_fill_1 FILLER_71_1140 ();
 sg13g2_fill_2 FILLER_71_1144 ();
 sg13g2_fill_2 FILLER_71_1152 ();
 sg13g2_decap_8 FILLER_71_1170 ();
 sg13g2_decap_4 FILLER_71_1177 ();
 sg13g2_fill_2 FILLER_71_1185 ();
 sg13g2_fill_1 FILLER_71_1187 ();
 sg13g2_decap_4 FILLER_71_1195 ();
 sg13g2_fill_2 FILLER_71_1199 ();
 sg13g2_decap_8 FILLER_71_1218 ();
 sg13g2_decap_8 FILLER_71_1225 ();
 sg13g2_fill_1 FILLER_71_1232 ();
 sg13g2_decap_4 FILLER_71_1237 ();
 sg13g2_fill_1 FILLER_71_1241 ();
 sg13g2_fill_2 FILLER_71_1251 ();
 sg13g2_fill_1 FILLER_71_1253 ();
 sg13g2_fill_2 FILLER_71_1257 ();
 sg13g2_fill_1 FILLER_71_1290 ();
 sg13g2_decap_8 FILLER_71_1300 ();
 sg13g2_decap_8 FILLER_71_1307 ();
 sg13g2_decap_8 FILLER_71_1314 ();
 sg13g2_decap_4 FILLER_71_1321 ();
 sg13g2_fill_1 FILLER_71_1325 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_fill_1 FILLER_72_33 ();
 sg13g2_fill_2 FILLER_72_68 ();
 sg13g2_fill_2 FILLER_72_96 ();
 sg13g2_fill_2 FILLER_72_102 ();
 sg13g2_fill_2 FILLER_72_110 ();
 sg13g2_fill_1 FILLER_72_112 ();
 sg13g2_decap_4 FILLER_72_118 ();
 sg13g2_fill_1 FILLER_72_122 ();
 sg13g2_decap_8 FILLER_72_150 ();
 sg13g2_decap_8 FILLER_72_157 ();
 sg13g2_decap_8 FILLER_72_164 ();
 sg13g2_decap_4 FILLER_72_181 ();
 sg13g2_fill_2 FILLER_72_185 ();
 sg13g2_fill_1 FILLER_72_197 ();
 sg13g2_decap_8 FILLER_72_226 ();
 sg13g2_decap_8 FILLER_72_233 ();
 sg13g2_fill_1 FILLER_72_240 ();
 sg13g2_fill_2 FILLER_72_266 ();
 sg13g2_fill_2 FILLER_72_302 ();
 sg13g2_decap_8 FILLER_72_307 ();
 sg13g2_decap_4 FILLER_72_314 ();
 sg13g2_fill_1 FILLER_72_318 ();
 sg13g2_fill_2 FILLER_72_339 ();
 sg13g2_fill_2 FILLER_72_346 ();
 sg13g2_fill_1 FILLER_72_348 ();
 sg13g2_decap_4 FILLER_72_358 ();
 sg13g2_fill_2 FILLER_72_362 ();
 sg13g2_fill_2 FILLER_72_382 ();
 sg13g2_fill_2 FILLER_72_398 ();
 sg13g2_fill_1 FILLER_72_400 ();
 sg13g2_decap_8 FILLER_72_418 ();
 sg13g2_fill_1 FILLER_72_432 ();
 sg13g2_fill_2 FILLER_72_461 ();
 sg13g2_fill_1 FILLER_72_471 ();
 sg13g2_fill_1 FILLER_72_476 ();
 sg13g2_fill_1 FILLER_72_486 ();
 sg13g2_decap_8 FILLER_72_497 ();
 sg13g2_fill_1 FILLER_72_504 ();
 sg13g2_fill_1 FILLER_72_518 ();
 sg13g2_fill_1 FILLER_72_523 ();
 sg13g2_fill_2 FILLER_72_529 ();
 sg13g2_fill_1 FILLER_72_531 ();
 sg13g2_decap_8 FILLER_72_541 ();
 sg13g2_decap_4 FILLER_72_548 ();
 sg13g2_fill_2 FILLER_72_560 ();
 sg13g2_decap_4 FILLER_72_567 ();
 sg13g2_fill_1 FILLER_72_571 ();
 sg13g2_fill_2 FILLER_72_576 ();
 sg13g2_decap_8 FILLER_72_583 ();
 sg13g2_fill_2 FILLER_72_633 ();
 sg13g2_decap_8 FILLER_72_639 ();
 sg13g2_fill_2 FILLER_72_646 ();
 sg13g2_fill_2 FILLER_72_652 ();
 sg13g2_decap_8 FILLER_72_663 ();
 sg13g2_fill_2 FILLER_72_710 ();
 sg13g2_decap_8 FILLER_72_716 ();
 sg13g2_decap_4 FILLER_72_723 ();
 sg13g2_fill_2 FILLER_72_727 ();
 sg13g2_decap_8 FILLER_72_751 ();
 sg13g2_decap_8 FILLER_72_758 ();
 sg13g2_decap_8 FILLER_72_765 ();
 sg13g2_decap_8 FILLER_72_772 ();
 sg13g2_decap_8 FILLER_72_779 ();
 sg13g2_fill_2 FILLER_72_786 ();
 sg13g2_decap_8 FILLER_72_792 ();
 sg13g2_decap_8 FILLER_72_799 ();
 sg13g2_decap_8 FILLER_72_806 ();
 sg13g2_fill_1 FILLER_72_836 ();
 sg13g2_fill_1 FILLER_72_842 ();
 sg13g2_decap_8 FILLER_72_847 ();
 sg13g2_decap_8 FILLER_72_854 ();
 sg13g2_decap_8 FILLER_72_861 ();
 sg13g2_decap_8 FILLER_72_868 ();
 sg13g2_fill_2 FILLER_72_875 ();
 sg13g2_fill_1 FILLER_72_877 ();
 sg13g2_decap_4 FILLER_72_882 ();
 sg13g2_fill_2 FILLER_72_886 ();
 sg13g2_fill_2 FILLER_72_902 ();
 sg13g2_fill_1 FILLER_72_908 ();
 sg13g2_fill_1 FILLER_72_916 ();
 sg13g2_fill_2 FILLER_72_920 ();
 sg13g2_fill_1 FILLER_72_922 ();
 sg13g2_decap_4 FILLER_72_931 ();
 sg13g2_fill_2 FILLER_72_954 ();
 sg13g2_fill_1 FILLER_72_956 ();
 sg13g2_fill_1 FILLER_72_967 ();
 sg13g2_fill_1 FILLER_72_986 ();
 sg13g2_decap_4 FILLER_72_996 ();
 sg13g2_decap_4 FILLER_72_1008 ();
 sg13g2_fill_1 FILLER_72_1012 ();
 sg13g2_fill_1 FILLER_72_1046 ();
 sg13g2_decap_8 FILLER_72_1055 ();
 sg13g2_fill_2 FILLER_72_1091 ();
 sg13g2_fill_1 FILLER_72_1103 ();
 sg13g2_fill_2 FILLER_72_1117 ();
 sg13g2_fill_1 FILLER_72_1119 ();
 sg13g2_decap_8 FILLER_72_1133 ();
 sg13g2_fill_2 FILLER_72_1140 ();
 sg13g2_fill_1 FILLER_72_1142 ();
 sg13g2_fill_1 FILLER_72_1161 ();
 sg13g2_fill_2 FILLER_72_1192 ();
 sg13g2_fill_2 FILLER_72_1198 ();
 sg13g2_decap_4 FILLER_72_1209 ();
 sg13g2_fill_2 FILLER_72_1213 ();
 sg13g2_decap_4 FILLER_72_1220 ();
 sg13g2_decap_8 FILLER_72_1234 ();
 sg13g2_decap_8 FILLER_72_1241 ();
 sg13g2_fill_1 FILLER_72_1248 ();
 sg13g2_fill_2 FILLER_72_1268 ();
 sg13g2_decap_8 FILLER_72_1275 ();
 sg13g2_decap_8 FILLER_72_1282 ();
 sg13g2_fill_1 FILLER_72_1289 ();
 sg13g2_decap_4 FILLER_72_1320 ();
 sg13g2_fill_2 FILLER_72_1324 ();
 sg13g2_fill_1 FILLER_73_26 ();
 sg13g2_decap_8 FILLER_73_36 ();
 sg13g2_decap_8 FILLER_73_43 ();
 sg13g2_fill_2 FILLER_73_50 ();
 sg13g2_decap_4 FILLER_73_56 ();
 sg13g2_fill_2 FILLER_73_60 ();
 sg13g2_fill_2 FILLER_73_66 ();
 sg13g2_decap_4 FILLER_73_73 ();
 sg13g2_fill_2 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_83 ();
 sg13g2_decap_8 FILLER_73_90 ();
 sg13g2_decap_8 FILLER_73_106 ();
 sg13g2_fill_2 FILLER_73_113 ();
 sg13g2_fill_1 FILLER_73_115 ();
 sg13g2_fill_1 FILLER_73_128 ();
 sg13g2_decap_8 FILLER_73_134 ();
 sg13g2_decap_4 FILLER_73_164 ();
 sg13g2_decap_4 FILLER_73_173 ();
 sg13g2_fill_1 FILLER_73_195 ();
 sg13g2_decap_4 FILLER_73_201 ();
 sg13g2_fill_2 FILLER_73_221 ();
 sg13g2_decap_8 FILLER_73_227 ();
 sg13g2_decap_4 FILLER_73_234 ();
 sg13g2_fill_2 FILLER_73_238 ();
 sg13g2_fill_1 FILLER_73_249 ();
 sg13g2_decap_8 FILLER_73_291 ();
 sg13g2_decap_8 FILLER_73_298 ();
 sg13g2_decap_4 FILLER_73_305 ();
 sg13g2_fill_2 FILLER_73_326 ();
 sg13g2_fill_1 FILLER_73_344 ();
 sg13g2_fill_2 FILLER_73_350 ();
 sg13g2_fill_1 FILLER_73_352 ();
 sg13g2_decap_4 FILLER_73_362 ();
 sg13g2_fill_2 FILLER_73_366 ();
 sg13g2_fill_1 FILLER_73_373 ();
 sg13g2_fill_2 FILLER_73_379 ();
 sg13g2_fill_2 FILLER_73_388 ();
 sg13g2_fill_1 FILLER_73_390 ();
 sg13g2_fill_2 FILLER_73_395 ();
 sg13g2_fill_1 FILLER_73_401 ();
 sg13g2_fill_2 FILLER_73_410 ();
 sg13g2_decap_8 FILLER_73_417 ();
 sg13g2_decap_4 FILLER_73_424 ();
 sg13g2_decap_4 FILLER_73_437 ();
 sg13g2_decap_4 FILLER_73_450 ();
 sg13g2_fill_2 FILLER_73_458 ();
 sg13g2_fill_2 FILLER_73_468 ();
 sg13g2_fill_1 FILLER_73_470 ();
 sg13g2_fill_2 FILLER_73_475 ();
 sg13g2_decap_8 FILLER_73_492 ();
 sg13g2_decap_8 FILLER_73_499 ();
 sg13g2_fill_2 FILLER_73_506 ();
 sg13g2_fill_1 FILLER_73_513 ();
 sg13g2_fill_1 FILLER_73_529 ();
 sg13g2_fill_2 FILLER_73_560 ();
 sg13g2_fill_1 FILLER_73_562 ();
 sg13g2_decap_4 FILLER_73_589 ();
 sg13g2_fill_1 FILLER_73_593 ();
 sg13g2_decap_8 FILLER_73_598 ();
 sg13g2_decap_8 FILLER_73_605 ();
 sg13g2_decap_8 FILLER_73_612 ();
 sg13g2_decap_8 FILLER_73_619 ();
 sg13g2_fill_1 FILLER_73_626 ();
 sg13g2_decap_8 FILLER_73_642 ();
 sg13g2_fill_1 FILLER_73_649 ();
 sg13g2_fill_1 FILLER_73_680 ();
 sg13g2_fill_1 FILLER_73_685 ();
 sg13g2_fill_1 FILLER_73_690 ();
 sg13g2_fill_1 FILLER_73_694 ();
 sg13g2_decap_8 FILLER_73_700 ();
 sg13g2_decap_4 FILLER_73_707 ();
 sg13g2_fill_2 FILLER_73_711 ();
 sg13g2_decap_8 FILLER_73_717 ();
 sg13g2_decap_4 FILLER_73_724 ();
 sg13g2_fill_2 FILLER_73_731 ();
 sg13g2_fill_1 FILLER_73_733 ();
 sg13g2_decap_8 FILLER_73_741 ();
 sg13g2_decap_8 FILLER_73_748 ();
 sg13g2_decap_4 FILLER_73_755 ();
 sg13g2_fill_2 FILLER_73_759 ();
 sg13g2_decap_8 FILLER_73_769 ();
 sg13g2_decap_4 FILLER_73_776 ();
 sg13g2_fill_1 FILLER_73_780 ();
 sg13g2_decap_4 FILLER_73_811 ();
 sg13g2_fill_2 FILLER_73_815 ();
 sg13g2_fill_2 FILLER_73_821 ();
 sg13g2_fill_1 FILLER_73_823 ();
 sg13g2_fill_2 FILLER_73_832 ();
 sg13g2_fill_2 FILLER_73_839 ();
 sg13g2_fill_1 FILLER_73_841 ();
 sg13g2_fill_2 FILLER_73_846 ();
 sg13g2_fill_1 FILLER_73_848 ();
 sg13g2_decap_8 FILLER_73_855 ();
 sg13g2_decap_4 FILLER_73_862 ();
 sg13g2_fill_2 FILLER_73_866 ();
 sg13g2_decap_8 FILLER_73_877 ();
 sg13g2_decap_4 FILLER_73_884 ();
 sg13g2_fill_1 FILLER_73_905 ();
 sg13g2_fill_1 FILLER_73_911 ();
 sg13g2_fill_1 FILLER_73_915 ();
 sg13g2_fill_1 FILLER_73_920 ();
 sg13g2_decap_8 FILLER_73_932 ();
 sg13g2_decap_8 FILLER_73_939 ();
 sg13g2_fill_2 FILLER_73_946 ();
 sg13g2_fill_1 FILLER_73_948 ();
 sg13g2_decap_4 FILLER_73_953 ();
 sg13g2_decap_4 FILLER_73_967 ();
 sg13g2_fill_1 FILLER_73_971 ();
 sg13g2_fill_2 FILLER_73_980 ();
 sg13g2_fill_1 FILLER_73_982 ();
 sg13g2_decap_4 FILLER_73_989 ();
 sg13g2_fill_2 FILLER_73_996 ();
 sg13g2_decap_8 FILLER_73_1002 ();
 sg13g2_decap_8 FILLER_73_1009 ();
 sg13g2_decap_8 FILLER_73_1016 ();
 sg13g2_fill_2 FILLER_73_1033 ();
 sg13g2_fill_1 FILLER_73_1043 ();
 sg13g2_fill_2 FILLER_73_1048 ();
 sg13g2_fill_1 FILLER_73_1050 ();
 sg13g2_decap_8 FILLER_73_1055 ();
 sg13g2_decap_4 FILLER_73_1062 ();
 sg13g2_fill_2 FILLER_73_1066 ();
 sg13g2_decap_4 FILLER_73_1076 ();
 sg13g2_decap_8 FILLER_73_1085 ();
 sg13g2_decap_8 FILLER_73_1092 ();
 sg13g2_decap_4 FILLER_73_1099 ();
 sg13g2_fill_2 FILLER_73_1120 ();
 sg13g2_fill_2 FILLER_73_1126 ();
 sg13g2_decap_8 FILLER_73_1136 ();
 sg13g2_fill_1 FILLER_73_1143 ();
 sg13g2_decap_8 FILLER_73_1163 ();
 sg13g2_decap_8 FILLER_73_1170 ();
 sg13g2_decap_8 FILLER_73_1177 ();
 sg13g2_decap_4 FILLER_73_1184 ();
 sg13g2_decap_4 FILLER_73_1192 ();
 sg13g2_fill_2 FILLER_73_1196 ();
 sg13g2_decap_8 FILLER_73_1201 ();
 sg13g2_fill_1 FILLER_73_1208 ();
 sg13g2_fill_1 FILLER_73_1218 ();
 sg13g2_fill_2 FILLER_73_1234 ();
 sg13g2_fill_1 FILLER_73_1236 ();
 sg13g2_fill_1 FILLER_73_1240 ();
 sg13g2_fill_2 FILLER_73_1250 ();
 sg13g2_fill_1 FILLER_73_1262 ();
 sg13g2_decap_8 FILLER_73_1268 ();
 sg13g2_decap_8 FILLER_73_1275 ();
 sg13g2_decap_8 FILLER_73_1282 ();
 sg13g2_decap_8 FILLER_73_1289 ();
 sg13g2_decap_8 FILLER_73_1296 ();
 sg13g2_decap_8 FILLER_73_1303 ();
 sg13g2_decap_8 FILLER_73_1310 ();
 sg13g2_decap_8 FILLER_73_1317 ();
 sg13g2_fill_2 FILLER_73_1324 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_4 FILLER_74_21 ();
 sg13g2_fill_2 FILLER_74_56 ();
 sg13g2_fill_1 FILLER_74_58 ();
 sg13g2_fill_1 FILLER_74_67 ();
 sg13g2_fill_1 FILLER_74_73 ();
 sg13g2_fill_1 FILLER_74_100 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_fill_1 FILLER_74_121 ();
 sg13g2_fill_1 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_132 ();
 sg13g2_decap_4 FILLER_74_139 ();
 sg13g2_decap_8 FILLER_74_164 ();
 sg13g2_fill_1 FILLER_74_185 ();
 sg13g2_decap_8 FILLER_74_207 ();
 sg13g2_fill_2 FILLER_74_214 ();
 sg13g2_fill_1 FILLER_74_216 ();
 sg13g2_fill_2 FILLER_74_251 ();
 sg13g2_fill_1 FILLER_74_259 ();
 sg13g2_fill_1 FILLER_74_263 ();
 sg13g2_fill_1 FILLER_74_269 ();
 sg13g2_fill_1 FILLER_74_273 ();
 sg13g2_fill_1 FILLER_74_278 ();
 sg13g2_fill_1 FILLER_74_283 ();
 sg13g2_fill_2 FILLER_74_290 ();
 sg13g2_fill_2 FILLER_74_350 ();
 sg13g2_fill_1 FILLER_74_361 ();
 sg13g2_decap_4 FILLER_74_367 ();
 sg13g2_decap_4 FILLER_74_375 ();
 sg13g2_fill_1 FILLER_74_379 ();
 sg13g2_fill_1 FILLER_74_391 ();
 sg13g2_fill_2 FILLER_74_400 ();
 sg13g2_decap_8 FILLER_74_417 ();
 sg13g2_fill_1 FILLER_74_424 ();
 sg13g2_decap_8 FILLER_74_437 ();
 sg13g2_decap_8 FILLER_74_444 ();
 sg13g2_decap_8 FILLER_74_451 ();
 sg13g2_fill_2 FILLER_74_458 ();
 sg13g2_decap_8 FILLER_74_465 ();
 sg13g2_decap_8 FILLER_74_472 ();
 sg13g2_fill_2 FILLER_74_489 ();
 sg13g2_fill_1 FILLER_74_496 ();
 sg13g2_decap_4 FILLER_74_502 ();
 sg13g2_fill_2 FILLER_74_509 ();
 sg13g2_fill_1 FILLER_74_524 ();
 sg13g2_decap_8 FILLER_74_528 ();
 sg13g2_decap_4 FILLER_74_535 ();
 sg13g2_fill_1 FILLER_74_539 ();
 sg13g2_decap_4 FILLER_74_550 ();
 sg13g2_fill_2 FILLER_74_558 ();
 sg13g2_decap_8 FILLER_74_568 ();
 sg13g2_decap_8 FILLER_74_575 ();
 sg13g2_decap_8 FILLER_74_582 ();
 sg13g2_decap_8 FILLER_74_589 ();
 sg13g2_decap_8 FILLER_74_596 ();
 sg13g2_fill_1 FILLER_74_603 ();
 sg13g2_decap_4 FILLER_74_609 ();
 sg13g2_fill_2 FILLER_74_613 ();
 sg13g2_fill_2 FILLER_74_619 ();
 sg13g2_fill_1 FILLER_74_621 ();
 sg13g2_decap_4 FILLER_74_627 ();
 sg13g2_fill_1 FILLER_74_636 ();
 sg13g2_fill_2 FILLER_74_641 ();
 sg13g2_fill_1 FILLER_74_647 ();
 sg13g2_fill_2 FILLER_74_653 ();
 sg13g2_decap_8 FILLER_74_660 ();
 sg13g2_fill_2 FILLER_74_667 ();
 sg13g2_decap_8 FILLER_74_673 ();
 sg13g2_decap_8 FILLER_74_680 ();
 sg13g2_decap_4 FILLER_74_687 ();
 sg13g2_fill_2 FILLER_74_691 ();
 sg13g2_fill_1 FILLER_74_697 ();
 sg13g2_fill_2 FILLER_74_724 ();
 sg13g2_fill_1 FILLER_74_726 ();
 sg13g2_decap_8 FILLER_74_755 ();
 sg13g2_fill_1 FILLER_74_762 ();
 sg13g2_fill_2 FILLER_74_781 ();
 sg13g2_fill_1 FILLER_74_813 ();
 sg13g2_decap_8 FILLER_74_837 ();
 sg13g2_decap_8 FILLER_74_844 ();
 sg13g2_decap_4 FILLER_74_851 ();
 sg13g2_fill_2 FILLER_74_855 ();
 sg13g2_fill_2 FILLER_74_904 ();
 sg13g2_fill_1 FILLER_74_906 ();
 sg13g2_fill_1 FILLER_74_915 ();
 sg13g2_fill_1 FILLER_74_921 ();
 sg13g2_fill_1 FILLER_74_926 ();
 sg13g2_fill_2 FILLER_74_935 ();
 sg13g2_decap_4 FILLER_74_941 ();
 sg13g2_fill_1 FILLER_74_945 ();
 sg13g2_fill_1 FILLER_74_971 ();
 sg13g2_fill_2 FILLER_74_975 ();
 sg13g2_decap_4 FILLER_74_1017 ();
 sg13g2_fill_1 FILLER_74_1021 ();
 sg13g2_fill_1 FILLER_74_1025 ();
 sg13g2_decap_4 FILLER_74_1041 ();
 sg13g2_decap_8 FILLER_74_1050 ();
 sg13g2_fill_2 FILLER_74_1057 ();
 sg13g2_decap_4 FILLER_74_1085 ();
 sg13g2_decap_8 FILLER_74_1094 ();
 sg13g2_decap_8 FILLER_74_1101 ();
 sg13g2_decap_8 FILLER_74_1108 ();
 sg13g2_fill_2 FILLER_74_1115 ();
 sg13g2_fill_1 FILLER_74_1117 ();
 sg13g2_decap_8 FILLER_74_1126 ();
 sg13g2_fill_2 FILLER_74_1133 ();
 sg13g2_decap_8 FILLER_74_1139 ();
 sg13g2_decap_8 FILLER_74_1146 ();
 sg13g2_decap_4 FILLER_74_1153 ();
 sg13g2_fill_1 FILLER_74_1162 ();
 sg13g2_fill_2 FILLER_74_1167 ();
 sg13g2_fill_1 FILLER_74_1169 ();
 sg13g2_fill_2 FILLER_74_1173 ();
 sg13g2_decap_8 FILLER_74_1179 ();
 sg13g2_decap_4 FILLER_74_1186 ();
 sg13g2_fill_1 FILLER_74_1190 ();
 sg13g2_fill_1 FILLER_74_1206 ();
 sg13g2_decap_4 FILLER_74_1215 ();
 sg13g2_decap_8 FILLER_74_1224 ();
 sg13g2_decap_8 FILLER_74_1231 ();
 sg13g2_fill_2 FILLER_74_1238 ();
 sg13g2_fill_1 FILLER_74_1240 ();
 sg13g2_fill_1 FILLER_74_1254 ();
 sg13g2_decap_8 FILLER_74_1260 ();
 sg13g2_decap_8 FILLER_74_1267 ();
 sg13g2_decap_8 FILLER_74_1274 ();
 sg13g2_decap_8 FILLER_74_1281 ();
 sg13g2_decap_8 FILLER_74_1288 ();
 sg13g2_decap_8 FILLER_74_1295 ();
 sg13g2_decap_8 FILLER_74_1302 ();
 sg13g2_decap_8 FILLER_74_1309 ();
 sg13g2_decap_8 FILLER_74_1316 ();
 sg13g2_fill_2 FILLER_74_1323 ();
 sg13g2_fill_1 FILLER_74_1325 ();
 sg13g2_fill_1 FILLER_75_30 ();
 sg13g2_decap_8 FILLER_75_36 ();
 sg13g2_decap_4 FILLER_75_43 ();
 sg13g2_fill_2 FILLER_75_78 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_98 ();
 sg13g2_decap_4 FILLER_75_103 ();
 sg13g2_fill_2 FILLER_75_107 ();
 sg13g2_fill_1 FILLER_75_113 ();
 sg13g2_decap_4 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_149 ();
 sg13g2_fill_2 FILLER_75_156 ();
 sg13g2_fill_2 FILLER_75_163 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_decap_4 FILLER_75_176 ();
 sg13g2_fill_1 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_207 ();
 sg13g2_fill_1 FILLER_75_211 ();
 sg13g2_fill_1 FILLER_75_216 ();
 sg13g2_fill_1 FILLER_75_221 ();
 sg13g2_fill_2 FILLER_75_229 ();
 sg13g2_decap_8 FILLER_75_235 ();
 sg13g2_decap_8 FILLER_75_242 ();
 sg13g2_fill_1 FILLER_75_249 ();
 sg13g2_fill_2 FILLER_75_262 ();
 sg13g2_fill_2 FILLER_75_274 ();
 sg13g2_fill_1 FILLER_75_276 ();
 sg13g2_decap_8 FILLER_75_289 ();
 sg13g2_decap_8 FILLER_75_296 ();
 sg13g2_decap_8 FILLER_75_303 ();
 sg13g2_decap_8 FILLER_75_310 ();
 sg13g2_fill_2 FILLER_75_317 ();
 sg13g2_fill_2 FILLER_75_336 ();
 sg13g2_fill_2 FILLER_75_343 ();
 sg13g2_fill_1 FILLER_75_353 ();
 sg13g2_decap_8 FILLER_75_358 ();
 sg13g2_decap_8 FILLER_75_365 ();
 sg13g2_fill_2 FILLER_75_372 ();
 sg13g2_fill_1 FILLER_75_374 ();
 sg13g2_fill_1 FILLER_75_395 ();
 sg13g2_fill_2 FILLER_75_401 ();
 sg13g2_fill_2 FILLER_75_410 ();
 sg13g2_decap_8 FILLER_75_419 ();
 sg13g2_fill_2 FILLER_75_426 ();
 sg13g2_fill_1 FILLER_75_432 ();
 sg13g2_fill_2 FILLER_75_441 ();
 sg13g2_decap_4 FILLER_75_447 ();
 sg13g2_decap_4 FILLER_75_455 ();
 sg13g2_fill_2 FILLER_75_459 ();
 sg13g2_decap_4 FILLER_75_466 ();
 sg13g2_fill_2 FILLER_75_477 ();
 sg13g2_decap_4 FILLER_75_489 ();
 sg13g2_decap_8 FILLER_75_498 ();
 sg13g2_fill_1 FILLER_75_505 ();
 sg13g2_decap_8 FILLER_75_519 ();
 sg13g2_decap_4 FILLER_75_526 ();
 sg13g2_fill_1 FILLER_75_530 ();
 sg13g2_decap_4 FILLER_75_540 ();
 sg13g2_fill_2 FILLER_75_544 ();
 sg13g2_decap_4 FILLER_75_572 ();
 sg13g2_fill_2 FILLER_75_576 ();
 sg13g2_fill_2 FILLER_75_591 ();
 sg13g2_fill_2 FILLER_75_617 ();
 sg13g2_decap_8 FILLER_75_622 ();
 sg13g2_decap_8 FILLER_75_629 ();
 sg13g2_decap_8 FILLER_75_636 ();
 sg13g2_decap_4 FILLER_75_643 ();
 sg13g2_fill_2 FILLER_75_647 ();
 sg13g2_fill_2 FILLER_75_675 ();
 sg13g2_fill_1 FILLER_75_677 ();
 sg13g2_decap_8 FILLER_75_709 ();
 sg13g2_fill_1 FILLER_75_716 ();
 sg13g2_fill_2 FILLER_75_721 ();
 sg13g2_decap_8 FILLER_75_732 ();
 sg13g2_fill_1 FILLER_75_739 ();
 sg13g2_fill_2 FILLER_75_764 ();
 sg13g2_fill_2 FILLER_75_770 ();
 sg13g2_fill_1 FILLER_75_772 ();
 sg13g2_decap_8 FILLER_75_778 ();
 sg13g2_fill_2 FILLER_75_785 ();
 sg13g2_decap_4 FILLER_75_792 ();
 sg13g2_decap_4 FILLER_75_826 ();
 sg13g2_fill_1 FILLER_75_830 ();
 sg13g2_decap_8 FILLER_75_866 ();
 sg13g2_decap_8 FILLER_75_873 ();
 sg13g2_decap_4 FILLER_75_880 ();
 sg13g2_fill_1 FILLER_75_884 ();
 sg13g2_decap_4 FILLER_75_889 ();
 sg13g2_fill_2 FILLER_75_893 ();
 sg13g2_decap_8 FILLER_75_900 ();
 sg13g2_decap_4 FILLER_75_907 ();
 sg13g2_fill_1 FILLER_75_911 ();
 sg13g2_decap_8 FILLER_75_917 ();
 sg13g2_decap_4 FILLER_75_924 ();
 sg13g2_decap_8 FILLER_75_937 ();
 sg13g2_fill_1 FILLER_75_955 ();
 sg13g2_fill_1 FILLER_75_960 ();
 sg13g2_fill_1 FILLER_75_965 ();
 sg13g2_fill_1 FILLER_75_971 ();
 sg13g2_fill_2 FILLER_75_992 ();
 sg13g2_fill_1 FILLER_75_994 ();
 sg13g2_decap_4 FILLER_75_999 ();
 sg13g2_decap_4 FILLER_75_1007 ();
 sg13g2_fill_2 FILLER_75_1011 ();
 sg13g2_decap_4 FILLER_75_1017 ();
 sg13g2_fill_2 FILLER_75_1021 ();
 sg13g2_fill_1 FILLER_75_1027 ();
 sg13g2_fill_1 FILLER_75_1032 ();
 sg13g2_fill_2 FILLER_75_1037 ();
 sg13g2_fill_1 FILLER_75_1044 ();
 sg13g2_fill_1 FILLER_75_1050 ();
 sg13g2_decap_4 FILLER_75_1055 ();
 sg13g2_decap_4 FILLER_75_1064 ();
 sg13g2_fill_1 FILLER_75_1068 ();
 sg13g2_decap_4 FILLER_75_1073 ();
 sg13g2_decap_8 FILLER_75_1082 ();
 sg13g2_decap_8 FILLER_75_1093 ();
 sg13g2_fill_1 FILLER_75_1100 ();
 sg13g2_fill_2 FILLER_75_1127 ();
 sg13g2_fill_2 FILLER_75_1133 ();
 sg13g2_fill_1 FILLER_75_1166 ();
 sg13g2_fill_1 FILLER_75_1174 ();
 sg13g2_fill_1 FILLER_75_1183 ();
 sg13g2_decap_8 FILLER_75_1189 ();
 sg13g2_decap_8 FILLER_75_1214 ();
 sg13g2_decap_8 FILLER_75_1221 ();
 sg13g2_decap_4 FILLER_75_1228 ();
 sg13g2_fill_2 FILLER_75_1232 ();
 sg13g2_decap_8 FILLER_75_1239 ();
 sg13g2_decap_8 FILLER_75_1246 ();
 sg13g2_decap_8 FILLER_75_1253 ();
 sg13g2_decap_8 FILLER_75_1260 ();
 sg13g2_decap_8 FILLER_75_1267 ();
 sg13g2_decap_8 FILLER_75_1274 ();
 sg13g2_decap_8 FILLER_75_1281 ();
 sg13g2_decap_8 FILLER_75_1288 ();
 sg13g2_decap_8 FILLER_75_1295 ();
 sg13g2_decap_8 FILLER_75_1302 ();
 sg13g2_decap_8 FILLER_75_1309 ();
 sg13g2_decap_8 FILLER_75_1316 ();
 sg13g2_fill_2 FILLER_75_1323 ();
 sg13g2_fill_1 FILLER_75_1325 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_16 ();
 sg13g2_fill_2 FILLER_76_29 ();
 sg13g2_fill_2 FILLER_76_37 ();
 sg13g2_fill_1 FILLER_76_39 ();
 sg13g2_fill_1 FILLER_76_44 ();
 sg13g2_fill_2 FILLER_76_50 ();
 sg13g2_fill_1 FILLER_76_52 ();
 sg13g2_fill_2 FILLER_76_61 ();
 sg13g2_decap_8 FILLER_76_67 ();
 sg13g2_fill_1 FILLER_76_74 ();
 sg13g2_decap_8 FILLER_76_110 ();
 sg13g2_decap_4 FILLER_76_117 ();
 sg13g2_fill_1 FILLER_76_121 ();
 sg13g2_decap_4 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_fill_1 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_152 ();
 sg13g2_fill_2 FILLER_76_159 ();
 sg13g2_fill_2 FILLER_76_180 ();
 sg13g2_fill_2 FILLER_76_194 ();
 sg13g2_fill_2 FILLER_76_208 ();
 sg13g2_fill_1 FILLER_76_222 ();
 sg13g2_decap_8 FILLER_76_227 ();
 sg13g2_decap_4 FILLER_76_234 ();
 sg13g2_fill_1 FILLER_76_238 ();
 sg13g2_fill_2 FILLER_76_243 ();
 sg13g2_decap_8 FILLER_76_292 ();
 sg13g2_decap_8 FILLER_76_299 ();
 sg13g2_decap_4 FILLER_76_306 ();
 sg13g2_fill_1 FILLER_76_310 ();
 sg13g2_fill_2 FILLER_76_320 ();
 sg13g2_fill_1 FILLER_76_330 ();
 sg13g2_decap_8 FILLER_76_352 ();
 sg13g2_decap_4 FILLER_76_359 ();
 sg13g2_fill_2 FILLER_76_363 ();
 sg13g2_decap_8 FILLER_76_370 ();
 sg13g2_decap_4 FILLER_76_381 ();
 sg13g2_fill_2 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_419 ();
 sg13g2_fill_1 FILLER_76_426 ();
 sg13g2_fill_1 FILLER_76_457 ();
 sg13g2_fill_1 FILLER_76_491 ();
 sg13g2_decap_4 FILLER_76_497 ();
 sg13g2_decap_4 FILLER_76_509 ();
 sg13g2_fill_1 FILLER_76_513 ();
 sg13g2_fill_2 FILLER_76_518 ();
 sg13g2_decap_8 FILLER_76_525 ();
 sg13g2_decap_4 FILLER_76_532 ();
 sg13g2_decap_4 FILLER_76_562 ();
 sg13g2_decap_4 FILLER_76_570 ();
 sg13g2_fill_1 FILLER_76_574 ();
 sg13g2_decap_8 FILLER_76_589 ();
 sg13g2_decap_8 FILLER_76_607 ();
 sg13g2_fill_1 FILLER_76_614 ();
 sg13g2_fill_2 FILLER_76_624 ();
 sg13g2_fill_2 FILLER_76_630 ();
 sg13g2_fill_1 FILLER_76_632 ();
 sg13g2_decap_8 FILLER_76_646 ();
 sg13g2_decap_4 FILLER_76_653 ();
 sg13g2_fill_2 FILLER_76_657 ();
 sg13g2_decap_8 FILLER_76_663 ();
 sg13g2_decap_4 FILLER_76_670 ();
 sg13g2_fill_1 FILLER_76_674 ();
 sg13g2_decap_8 FILLER_76_705 ();
 sg13g2_decap_8 FILLER_76_712 ();
 sg13g2_fill_1 FILLER_76_719 ();
 sg13g2_fill_2 FILLER_76_724 ();
 sg13g2_fill_1 FILLER_76_731 ();
 sg13g2_fill_1 FILLER_76_745 ();
 sg13g2_decap_8 FILLER_76_759 ();
 sg13g2_fill_2 FILLER_76_766 ();
 sg13g2_decap_8 FILLER_76_772 ();
 sg13g2_decap_8 FILLER_76_779 ();
 sg13g2_decap_8 FILLER_76_786 ();
 sg13g2_decap_4 FILLER_76_793 ();
 sg13g2_fill_1 FILLER_76_797 ();
 sg13g2_decap_8 FILLER_76_807 ();
 sg13g2_decap_8 FILLER_76_826 ();
 sg13g2_decap_8 FILLER_76_838 ();
 sg13g2_decap_4 FILLER_76_845 ();
 sg13g2_fill_1 FILLER_76_849 ();
 sg13g2_fill_2 FILLER_76_858 ();
 sg13g2_fill_2 FILLER_76_891 ();
 sg13g2_fill_1 FILLER_76_893 ();
 sg13g2_fill_2 FILLER_76_950 ();
 sg13g2_fill_1 FILLER_76_952 ();
 sg13g2_fill_1 FILLER_76_957 ();
 sg13g2_decap_8 FILLER_76_970 ();
 sg13g2_decap_8 FILLER_76_977 ();
 sg13g2_decap_8 FILLER_76_984 ();
 sg13g2_decap_8 FILLER_76_991 ();
 sg13g2_fill_1 FILLER_76_998 ();
 sg13g2_fill_2 FILLER_76_1016 ();
 sg13g2_decap_8 FILLER_76_1023 ();
 sg13g2_decap_8 FILLER_76_1030 ();
 sg13g2_fill_1 FILLER_76_1037 ();
 sg13g2_decap_8 FILLER_76_1043 ();
 sg13g2_decap_4 FILLER_76_1050 ();
 sg13g2_fill_2 FILLER_76_1054 ();
 sg13g2_decap_8 FILLER_76_1091 ();
 sg13g2_decap_8 FILLER_76_1098 ();
 sg13g2_fill_2 FILLER_76_1105 ();
 sg13g2_fill_2 FILLER_76_1115 ();
 sg13g2_decap_4 FILLER_76_1122 ();
 sg13g2_decap_8 FILLER_76_1130 ();
 sg13g2_decap_8 FILLER_76_1137 ();
 sg13g2_decap_8 FILLER_76_1144 ();
 sg13g2_decap_8 FILLER_76_1151 ();
 sg13g2_decap_8 FILLER_76_1158 ();
 sg13g2_decap_8 FILLER_76_1165 ();
 sg13g2_fill_1 FILLER_76_1172 ();
 sg13g2_decap_8 FILLER_76_1177 ();
 sg13g2_decap_8 FILLER_76_1184 ();
 sg13g2_decap_8 FILLER_76_1191 ();
 sg13g2_decap_8 FILLER_76_1198 ();
 sg13g2_fill_2 FILLER_76_1205 ();
 sg13g2_decap_8 FILLER_76_1214 ();
 sg13g2_decap_8 FILLER_76_1221 ();
 sg13g2_fill_2 FILLER_76_1228 ();
 sg13g2_fill_1 FILLER_76_1230 ();
 sg13g2_fill_1 FILLER_76_1247 ();
 sg13g2_decap_8 FILLER_76_1253 ();
 sg13g2_decap_8 FILLER_76_1260 ();
 sg13g2_decap_8 FILLER_76_1267 ();
 sg13g2_decap_8 FILLER_76_1274 ();
 sg13g2_decap_8 FILLER_76_1281 ();
 sg13g2_decap_8 FILLER_76_1288 ();
 sg13g2_decap_8 FILLER_76_1295 ();
 sg13g2_decap_8 FILLER_76_1302 ();
 sg13g2_decap_8 FILLER_76_1309 ();
 sg13g2_decap_8 FILLER_76_1316 ();
 sg13g2_fill_2 FILLER_76_1323 ();
 sg13g2_fill_1 FILLER_76_1325 ();
 sg13g2_decap_4 FILLER_77_26 ();
 sg13g2_fill_2 FILLER_77_35 ();
 sg13g2_fill_1 FILLER_77_37 ();
 sg13g2_decap_4 FILLER_77_50 ();
 sg13g2_fill_2 FILLER_77_94 ();
 sg13g2_fill_1 FILLER_77_96 ();
 sg13g2_decap_8 FILLER_77_101 ();
 sg13g2_fill_2 FILLER_77_108 ();
 sg13g2_decap_4 FILLER_77_118 ();
 sg13g2_fill_2 FILLER_77_126 ();
 sg13g2_fill_1 FILLER_77_133 ();
 sg13g2_fill_1 FILLER_77_160 ();
 sg13g2_decap_4 FILLER_77_164 ();
 sg13g2_decap_8 FILLER_77_172 ();
 sg13g2_fill_1 FILLER_77_179 ();
 sg13g2_fill_1 FILLER_77_204 ();
 sg13g2_decap_8 FILLER_77_209 ();
 sg13g2_fill_1 FILLER_77_216 ();
 sg13g2_decap_8 FILLER_77_221 ();
 sg13g2_decap_8 FILLER_77_228 ();
 sg13g2_decap_4 FILLER_77_235 ();
 sg13g2_fill_2 FILLER_77_250 ();
 sg13g2_fill_2 FILLER_77_273 ();
 sg13g2_decap_4 FILLER_77_314 ();
 sg13g2_fill_1 FILLER_77_343 ();
 sg13g2_fill_2 FILLER_77_349 ();
 sg13g2_fill_1 FILLER_77_351 ();
 sg13g2_fill_1 FILLER_77_382 ();
 sg13g2_fill_1 FILLER_77_398 ();
 sg13g2_decap_8 FILLER_77_438 ();
 sg13g2_decap_8 FILLER_77_445 ();
 sg13g2_decap_8 FILLER_77_452 ();
 sg13g2_fill_2 FILLER_77_459 ();
 sg13g2_decap_8 FILLER_77_474 ();
 sg13g2_decap_8 FILLER_77_481 ();
 sg13g2_fill_1 FILLER_77_488 ();
 sg13g2_decap_8 FILLER_77_524 ();
 sg13g2_decap_8 FILLER_77_531 ();
 sg13g2_decap_8 FILLER_77_538 ();
 sg13g2_decap_4 FILLER_77_545 ();
 sg13g2_fill_2 FILLER_77_549 ();
 sg13g2_decap_8 FILLER_77_563 ();
 sg13g2_fill_2 FILLER_77_570 ();
 sg13g2_fill_2 FILLER_77_580 ();
 sg13g2_fill_1 FILLER_77_582 ();
 sg13g2_decap_8 FILLER_77_609 ();
 sg13g2_decap_8 FILLER_77_616 ();
 sg13g2_decap_4 FILLER_77_623 ();
 sg13g2_decap_8 FILLER_77_653 ();
 sg13g2_decap_8 FILLER_77_660 ();
 sg13g2_decap_8 FILLER_77_667 ();
 sg13g2_decap_8 FILLER_77_674 ();
 sg13g2_decap_4 FILLER_77_681 ();
 sg13g2_fill_1 FILLER_77_685 ();
 sg13g2_decap_8 FILLER_77_694 ();
 sg13g2_fill_1 FILLER_77_758 ();
 sg13g2_fill_1 FILLER_77_764 ();
 sg13g2_fill_2 FILLER_77_770 ();
 sg13g2_fill_2 FILLER_77_777 ();
 sg13g2_decap_8 FILLER_77_784 ();
 sg13g2_decap_4 FILLER_77_791 ();
 sg13g2_fill_2 FILLER_77_795 ();
 sg13g2_decap_8 FILLER_77_806 ();
 sg13g2_decap_8 FILLER_77_813 ();
 sg13g2_decap_8 FILLER_77_820 ();
 sg13g2_decap_4 FILLER_77_827 ();
 sg13g2_fill_2 FILLER_77_831 ();
 sg13g2_fill_2 FILLER_77_859 ();
 sg13g2_decap_8 FILLER_77_887 ();
 sg13g2_decap_4 FILLER_77_894 ();
 sg13g2_fill_2 FILLER_77_898 ();
 sg13g2_decap_4 FILLER_77_904 ();
 sg13g2_fill_2 FILLER_77_913 ();
 sg13g2_decap_8 FILLER_77_919 ();
 sg13g2_decap_8 FILLER_77_926 ();
 sg13g2_decap_8 FILLER_77_933 ();
 sg13g2_decap_8 FILLER_77_940 ();
 sg13g2_decap_8 FILLER_77_947 ();
 sg13g2_decap_8 FILLER_77_954 ();
 sg13g2_decap_4 FILLER_77_961 ();
 sg13g2_decap_8 FILLER_77_969 ();
 sg13g2_decap_8 FILLER_77_976 ();
 sg13g2_fill_1 FILLER_77_983 ();
 sg13g2_fill_1 FILLER_77_993 ();
 sg13g2_fill_2 FILLER_77_998 ();
 sg13g2_fill_1 FILLER_77_1000 ();
 sg13g2_decap_4 FILLER_77_1010 ();
 sg13g2_fill_1 FILLER_77_1014 ();
 sg13g2_fill_1 FILLER_77_1028 ();
 sg13g2_decap_8 FILLER_77_1034 ();
 sg13g2_fill_1 FILLER_77_1041 ();
 sg13g2_fill_1 FILLER_77_1059 ();
 sg13g2_fill_2 FILLER_77_1064 ();
 sg13g2_decap_8 FILLER_77_1070 ();
 sg13g2_fill_2 FILLER_77_1077 ();
 sg13g2_decap_8 FILLER_77_1083 ();
 sg13g2_decap_8 FILLER_77_1090 ();
 sg13g2_decap_8 FILLER_77_1097 ();
 sg13g2_decap_4 FILLER_77_1104 ();
 sg13g2_fill_1 FILLER_77_1108 ();
 sg13g2_fill_2 FILLER_77_1135 ();
 sg13g2_decap_8 FILLER_77_1142 ();
 sg13g2_fill_2 FILLER_77_1149 ();
 sg13g2_decap_8 FILLER_77_1173 ();
 sg13g2_fill_2 FILLER_77_1180 ();
 sg13g2_fill_1 FILLER_77_1182 ();
 sg13g2_fill_1 FILLER_77_1214 ();
 sg13g2_decap_8 FILLER_77_1221 ();
 sg13g2_fill_2 FILLER_77_1228 ();
 sg13g2_fill_2 FILLER_77_1253 ();
 sg13g2_decap_8 FILLER_77_1268 ();
 sg13g2_decap_8 FILLER_77_1275 ();
 sg13g2_decap_8 FILLER_77_1282 ();
 sg13g2_decap_8 FILLER_77_1289 ();
 sg13g2_decap_8 FILLER_77_1296 ();
 sg13g2_decap_8 FILLER_77_1303 ();
 sg13g2_decap_8 FILLER_77_1310 ();
 sg13g2_decap_8 FILLER_77_1317 ();
 sg13g2_fill_2 FILLER_77_1324 ();
 sg13g2_decap_8 FILLER_78_26 ();
 sg13g2_decap_8 FILLER_78_69 ();
 sg13g2_decap_8 FILLER_78_76 ();
 sg13g2_decap_8 FILLER_78_83 ();
 sg13g2_decap_8 FILLER_78_90 ();
 sg13g2_fill_2 FILLER_78_97 ();
 sg13g2_decap_8 FILLER_78_129 ();
 sg13g2_decap_8 FILLER_78_136 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_4 FILLER_78_175 ();
 sg13g2_fill_1 FILLER_78_179 ();
 sg13g2_fill_1 FILLER_78_208 ();
 sg13g2_fill_2 FILLER_78_218 ();
 sg13g2_fill_2 FILLER_78_225 ();
 sg13g2_fill_2 FILLER_78_232 ();
 sg13g2_fill_1 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_243 ();
 sg13g2_decap_8 FILLER_78_286 ();
 sg13g2_decap_8 FILLER_78_293 ();
 sg13g2_decap_4 FILLER_78_300 ();
 sg13g2_fill_2 FILLER_78_304 ();
 sg13g2_decap_4 FILLER_78_311 ();
 sg13g2_fill_1 FILLER_78_325 ();
 sg13g2_fill_2 FILLER_78_341 ();
 sg13g2_fill_1 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_349 ();
 sg13g2_fill_1 FILLER_78_360 ();
 sg13g2_decap_8 FILLER_78_366 ();
 sg13g2_decap_8 FILLER_78_373 ();
 sg13g2_decap_4 FILLER_78_380 ();
 sg13g2_fill_1 FILLER_78_384 ();
 sg13g2_fill_2 FILLER_78_406 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_fill_2 FILLER_78_413 ();
 sg13g2_fill_2 FILLER_78_420 ();
 sg13g2_fill_1 FILLER_78_422 ();
 sg13g2_fill_2 FILLER_78_427 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_fill_2 FILLER_78_434 ();
 sg13g2_fill_1 FILLER_78_436 ();
 sg13g2_fill_2 FILLER_78_441 ();
 sg13g2_fill_1 FILLER_78_443 ();
 sg13g2_decap_8 FILLER_78_474 ();
 sg13g2_fill_2 FILLER_78_481 ();
 sg13g2_decap_4 FILLER_78_488 ();
 sg13g2_fill_2 FILLER_78_492 ();
 sg13g2_fill_1 FILLER_78_498 ();
 sg13g2_decap_8 FILLER_78_508 ();
 sg13g2_fill_2 FILLER_78_515 ();
 sg13g2_fill_1 FILLER_78_521 ();
 sg13g2_fill_2 FILLER_78_526 ();
 sg13g2_fill_1 FILLER_78_528 ();
 sg13g2_decap_8 FILLER_78_534 ();
 sg13g2_fill_1 FILLER_78_541 ();
 sg13g2_decap_8 FILLER_78_547 ();
 sg13g2_decap_8 FILLER_78_558 ();
 sg13g2_fill_1 FILLER_78_565 ();
 sg13g2_decap_8 FILLER_78_570 ();
 sg13g2_fill_1 FILLER_78_577 ();
 sg13g2_fill_1 FILLER_78_583 ();
 sg13g2_fill_2 FILLER_78_597 ();
 sg13g2_fill_1 FILLER_78_599 ();
 sg13g2_decap_4 FILLER_78_612 ();
 sg13g2_fill_1 FILLER_78_616 ();
 sg13g2_fill_1 FILLER_78_635 ();
 sg13g2_fill_1 FILLER_78_640 ();
 sg13g2_fill_1 FILLER_78_659 ();
 sg13g2_fill_1 FILLER_78_665 ();
 sg13g2_fill_1 FILLER_78_671 ();
 sg13g2_fill_2 FILLER_78_676 ();
 sg13g2_decap_4 FILLER_78_682 ();
 sg13g2_fill_2 FILLER_78_691 ();
 sg13g2_fill_1 FILLER_78_693 ();
 sg13g2_fill_1 FILLER_78_699 ();
 sg13g2_decap_4 FILLER_78_716 ();
 sg13g2_fill_2 FILLER_78_720 ();
 sg13g2_fill_1 FILLER_78_727 ();
 sg13g2_fill_2 FILLER_78_762 ();
 sg13g2_decap_4 FILLER_78_790 ();
 sg13g2_fill_1 FILLER_78_794 ();
 sg13g2_decap_4 FILLER_78_821 ();
 sg13g2_fill_2 FILLER_78_825 ();
 sg13g2_fill_1 FILLER_78_858 ();
 sg13g2_fill_2 FILLER_78_868 ();
 sg13g2_decap_8 FILLER_78_922 ();
 sg13g2_decap_8 FILLER_78_929 ();
 sg13g2_fill_1 FILLER_78_936 ();
 sg13g2_decap_4 FILLER_78_972 ();
 sg13g2_decap_8 FILLER_78_980 ();
 sg13g2_decap_4 FILLER_78_987 ();
 sg13g2_decap_4 FILLER_78_997 ();
 sg13g2_fill_1 FILLER_78_1001 ();
 sg13g2_fill_2 FILLER_78_1026 ();
 sg13g2_fill_1 FILLER_78_1048 ();
 sg13g2_fill_1 FILLER_78_1067 ();
 sg13g2_decap_8 FILLER_78_1073 ();
 sg13g2_fill_2 FILLER_78_1080 ();
 sg13g2_decap_8 FILLER_78_1091 ();
 sg13g2_decap_4 FILLER_78_1107 ();
 sg13g2_fill_1 FILLER_78_1111 ();
 sg13g2_fill_2 FILLER_78_1121 ();
 sg13g2_fill_1 FILLER_78_1123 ();
 sg13g2_fill_2 FILLER_78_1137 ();
 sg13g2_fill_1 FILLER_78_1139 ();
 sg13g2_fill_1 FILLER_78_1167 ();
 sg13g2_fill_2 FILLER_78_1182 ();
 sg13g2_fill_2 FILLER_78_1188 ();
 sg13g2_fill_1 FILLER_78_1190 ();
 sg13g2_fill_1 FILLER_78_1195 ();
 sg13g2_decap_8 FILLER_78_1216 ();
 sg13g2_decap_4 FILLER_78_1223 ();
 sg13g2_fill_2 FILLER_78_1227 ();
 sg13g2_fill_1 FILLER_78_1233 ();
 sg13g2_decap_8 FILLER_78_1238 ();
 sg13g2_decap_8 FILLER_78_1249 ();
 sg13g2_decap_8 FILLER_78_1256 ();
 sg13g2_decap_8 FILLER_78_1263 ();
 sg13g2_decap_8 FILLER_78_1270 ();
 sg13g2_decap_8 FILLER_78_1277 ();
 sg13g2_decap_8 FILLER_78_1284 ();
 sg13g2_decap_8 FILLER_78_1291 ();
 sg13g2_decap_8 FILLER_78_1298 ();
 sg13g2_decap_8 FILLER_78_1305 ();
 sg13g2_decap_8 FILLER_78_1312 ();
 sg13g2_decap_8 FILLER_78_1319 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_2 FILLER_79_11 ();
 sg13g2_decap_8 FILLER_79_20 ();
 sg13g2_fill_1 FILLER_79_31 ();
 sg13g2_decap_8 FILLER_79_37 ();
 sg13g2_decap_4 FILLER_79_44 ();
 sg13g2_fill_1 FILLER_79_92 ();
 sg13g2_fill_2 FILLER_79_97 ();
 sg13g2_fill_2 FILLER_79_103 ();
 sg13g2_fill_2 FILLER_79_113 ();
 sg13g2_fill_1 FILLER_79_115 ();
 sg13g2_decap_4 FILLER_79_120 ();
 sg13g2_fill_1 FILLER_79_159 ();
 sg13g2_decap_8 FILLER_79_165 ();
 sg13g2_decap_8 FILLER_79_172 ();
 sg13g2_fill_1 FILLER_79_179 ();
 sg13g2_decap_4 FILLER_79_184 ();
 sg13g2_fill_2 FILLER_79_188 ();
 sg13g2_fill_2 FILLER_79_220 ();
 sg13g2_fill_1 FILLER_79_222 ();
 sg13g2_decap_8 FILLER_79_249 ();
 sg13g2_decap_8 FILLER_79_443 ();
 sg13g2_decap_8 FILLER_79_450 ();
 sg13g2_fill_2 FILLER_79_457 ();
 sg13g2_fill_1 FILLER_79_459 ();
 sg13g2_fill_1 FILLER_79_474 ();
 sg13g2_fill_2 FILLER_79_501 ();
 sg13g2_fill_2 FILLER_79_529 ();
 sg13g2_fill_2 FILLER_79_557 ();
 sg13g2_decap_4 FILLER_79_603 ();
 sg13g2_fill_1 FILLER_79_607 ();
 sg13g2_decap_8 FILLER_79_612 ();
 sg13g2_decap_8 FILLER_79_619 ();
 sg13g2_decap_4 FILLER_79_626 ();
 sg13g2_fill_2 FILLER_79_641 ();
 sg13g2_decap_8 FILLER_79_646 ();
 sg13g2_fill_2 FILLER_79_653 ();
 sg13g2_fill_1 FILLER_79_655 ();
 sg13g2_decap_8 FILLER_79_665 ();
 sg13g2_decap_8 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_679 ();
 sg13g2_decap_4 FILLER_79_738 ();
 sg13g2_fill_1 FILLER_79_742 ();
 sg13g2_decap_8 FILLER_79_772 ();
 sg13g2_fill_1 FILLER_79_805 ();
 sg13g2_decap_8 FILLER_79_832 ();
 sg13g2_decap_4 FILLER_79_839 ();
 sg13g2_fill_2 FILLER_79_843 ();
 sg13g2_decap_8 FILLER_79_848 ();
 sg13g2_fill_2 FILLER_79_855 ();
 sg13g2_fill_1 FILLER_79_857 ();
 sg13g2_decap_4 FILLER_79_884 ();
 sg13g2_fill_2 FILLER_79_888 ();
 sg13g2_decap_8 FILLER_79_894 ();
 sg13g2_decap_4 FILLER_79_901 ();
 sg13g2_decap_8 FILLER_79_923 ();
 sg13g2_fill_2 FILLER_79_930 ();
 sg13g2_fill_1 FILLER_79_932 ();
 sg13g2_fill_2 FILLER_79_1014 ();
 sg13g2_fill_1 FILLER_79_1032 ();
 sg13g2_decap_4 FILLER_79_1038 ();
 sg13g2_fill_2 FILLER_79_1042 ();
 sg13g2_fill_1 FILLER_79_1057 ();
 sg13g2_fill_2 FILLER_79_1075 ();
 sg13g2_fill_1 FILLER_79_1077 ();
 sg13g2_fill_2 FILLER_79_1109 ();
 sg13g2_fill_2 FILLER_79_1142 ();
 sg13g2_fill_2 FILLER_79_1156 ();
 sg13g2_fill_1 FILLER_79_1166 ();
 sg13g2_decap_8 FILLER_79_1175 ();
 sg13g2_decap_4 FILLER_79_1182 ();
 sg13g2_fill_2 FILLER_79_1186 ();
 sg13g2_fill_2 FILLER_79_1195 ();
 sg13g2_decap_4 FILLER_79_1201 ();
 sg13g2_fill_2 FILLER_79_1205 ();
 sg13g2_decap_4 FILLER_79_1224 ();
 sg13g2_decap_8 FILLER_79_1239 ();
 sg13g2_decap_8 FILLER_79_1246 ();
 sg13g2_decap_8 FILLER_79_1253 ();
 sg13g2_decap_8 FILLER_79_1260 ();
 sg13g2_decap_8 FILLER_79_1267 ();
 sg13g2_decap_8 FILLER_79_1274 ();
 sg13g2_decap_8 FILLER_79_1281 ();
 sg13g2_decap_8 FILLER_79_1288 ();
 sg13g2_decap_8 FILLER_79_1295 ();
 sg13g2_decap_8 FILLER_79_1302 ();
 sg13g2_decap_8 FILLER_79_1309 ();
 sg13g2_decap_8 FILLER_79_1316 ();
 sg13g2_fill_2 FILLER_79_1323 ();
 sg13g2_fill_1 FILLER_79_1325 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_4 FILLER_80_14 ();
 sg13g2_fill_2 FILLER_80_18 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_4 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_74 ();
 sg13g2_fill_1 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_128 ();
 sg13g2_fill_2 FILLER_80_133 ();
 sg13g2_fill_2 FILLER_80_140 ();
 sg13g2_fill_2 FILLER_80_146 ();
 sg13g2_fill_1 FILLER_80_160 ();
 sg13g2_fill_2 FILLER_80_169 ();
 sg13g2_fill_1 FILLER_80_171 ();
 sg13g2_fill_2 FILLER_80_192 ();
 sg13g2_decap_8 FILLER_80_206 ();
 sg13g2_fill_1 FILLER_80_213 ();
 sg13g2_decap_4 FILLER_80_218 ();
 sg13g2_decap_4 FILLER_80_250 ();
 sg13g2_fill_1 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_289 ();
 sg13g2_fill_1 FILLER_80_296 ();
 sg13g2_decap_4 FILLER_80_318 ();
 sg13g2_decap_4 FILLER_80_326 ();
 sg13g2_decap_4 FILLER_80_334 ();
 sg13g2_fill_1 FILLER_80_338 ();
 sg13g2_fill_2 FILLER_80_352 ();
 sg13g2_decap_4 FILLER_80_359 ();
 sg13g2_decap_8 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_378 ();
 sg13g2_fill_1 FILLER_80_385 ();
 sg13g2_decap_8 FILLER_80_396 ();
 sg13g2_decap_8 FILLER_80_403 ();
 sg13g2_decap_4 FILLER_80_410 ();
 sg13g2_fill_1 FILLER_80_414 ();
 sg13g2_decap_4 FILLER_80_419 ();
 sg13g2_decap_8 FILLER_80_435 ();
 sg13g2_decap_8 FILLER_80_442 ();
 sg13g2_decap_8 FILLER_80_480 ();
 sg13g2_decap_8 FILLER_80_487 ();
 sg13g2_decap_8 FILLER_80_494 ();
 sg13g2_decap_8 FILLER_80_501 ();
 sg13g2_decap_4 FILLER_80_508 ();
 sg13g2_fill_1 FILLER_80_512 ();
 sg13g2_decap_8 FILLER_80_518 ();
 sg13g2_decap_8 FILLER_80_525 ();
 sg13g2_decap_4 FILLER_80_532 ();
 sg13g2_fill_1 FILLER_80_544 ();
 sg13g2_decap_8 FILLER_80_571 ();
 sg13g2_decap_4 FILLER_80_578 ();
 sg13g2_fill_2 FILLER_80_582 ();
 sg13g2_decap_8 FILLER_80_592 ();
 sg13g2_decap_8 FILLER_80_629 ();
 sg13g2_fill_1 FILLER_80_636 ();
 sg13g2_decap_8 FILLER_80_645 ();
 sg13g2_decap_8 FILLER_80_652 ();
 sg13g2_decap_4 FILLER_80_690 ();
 sg13g2_fill_2 FILLER_80_699 ();
 sg13g2_fill_1 FILLER_80_701 ();
 sg13g2_fill_2 FILLER_80_707 ();
 sg13g2_decap_8 FILLER_80_719 ();
 sg13g2_decap_8 FILLER_80_726 ();
 sg13g2_decap_8 FILLER_80_733 ();
 sg13g2_decap_8 FILLER_80_740 ();
 sg13g2_decap_8 FILLER_80_773 ();
 sg13g2_decap_8 FILLER_80_780 ();
 sg13g2_decap_8 FILLER_80_787 ();
 sg13g2_decap_8 FILLER_80_794 ();
 sg13g2_fill_2 FILLER_80_801 ();
 sg13g2_fill_1 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_809 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_fill_2 FILLER_80_823 ();
 sg13g2_decap_8 FILLER_80_829 ();
 sg13g2_decap_8 FILLER_80_836 ();
 sg13g2_fill_2 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_850 ();
 sg13g2_decap_8 FILLER_80_857 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_fill_2 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_893 ();
 sg13g2_decap_4 FILLER_80_926 ();
 sg13g2_decap_8 FILLER_80_939 ();
 sg13g2_decap_4 FILLER_80_946 ();
 sg13g2_fill_2 FILLER_80_950 ();
 sg13g2_decap_8 FILLER_80_982 ();
 sg13g2_decap_8 FILLER_80_989 ();
 sg13g2_decap_8 FILLER_80_996 ();
 sg13g2_decap_8 FILLER_80_1003 ();
 sg13g2_decap_4 FILLER_80_1010 ();
 sg13g2_fill_2 FILLER_80_1014 ();
 sg13g2_decap_8 FILLER_80_1020 ();
 sg13g2_fill_2 FILLER_80_1027 ();
 sg13g2_fill_1 FILLER_80_1029 ();
 sg13g2_decap_8 FILLER_80_1042 ();
 sg13g2_decap_8 FILLER_80_1049 ();
 sg13g2_decap_8 FILLER_80_1064 ();
 sg13g2_fill_2 FILLER_80_1071 ();
 sg13g2_decap_8 FILLER_80_1078 ();
 sg13g2_decap_8 FILLER_80_1085 ();
 sg13g2_decap_8 FILLER_80_1092 ();
 sg13g2_decap_8 FILLER_80_1099 ();
 sg13g2_decap_8 FILLER_80_1106 ();
 sg13g2_decap_8 FILLER_80_1113 ();
 sg13g2_decap_8 FILLER_80_1120 ();
 sg13g2_decap_4 FILLER_80_1127 ();
 sg13g2_fill_1 FILLER_80_1131 ();
 sg13g2_decap_8 FILLER_80_1172 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_decap_8 FILLER_80_1186 ();
 sg13g2_fill_2 FILLER_80_1193 ();
 sg13g2_fill_1 FILLER_80_1195 ();
 sg13g2_decap_8 FILLER_80_1202 ();
 sg13g2_decap_8 FILLER_80_1209 ();
 sg13g2_decap_8 FILLER_80_1216 ();
 sg13g2_decap_8 FILLER_80_1223 ();
 sg13g2_decap_8 FILLER_80_1230 ();
 sg13g2_decap_8 FILLER_80_1237 ();
 sg13g2_decap_8 FILLER_80_1244 ();
 sg13g2_decap_8 FILLER_80_1251 ();
 sg13g2_decap_8 FILLER_80_1258 ();
 sg13g2_decap_8 FILLER_80_1265 ();
 sg13g2_decap_8 FILLER_80_1272 ();
 sg13g2_decap_8 FILLER_80_1279 ();
 sg13g2_decap_8 FILLER_80_1286 ();
 sg13g2_decap_8 FILLER_80_1293 ();
 sg13g2_decap_8 FILLER_80_1300 ();
 sg13g2_decap_8 FILLER_80_1307 ();
 sg13g2_decap_8 FILLER_80_1314 ();
 sg13g2_decap_4 FILLER_80_1321 ();
 sg13g2_fill_1 FILLER_80_1325 ();
endmodule
