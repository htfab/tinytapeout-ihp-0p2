module tt_um_calonso88_rsa (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire clknet_leaf_0_clk;
 wire net155;
 wire cpha_sync;
 wire cpol_sync;
 wire eoc_rsa;
 wire \gpio_wrapper_i.gpio_start_cmd_i.data ;
 wire \gpio_wrapper_i.gpio_start_cmd_i.data_dly ;
 wire \gpio_wrapper_i.gpio_stop_cmd_i.data ;
 wire \gpio_wrapper_i.gpio_stop_cmd_i.data_dly ;
 wire \gpio_wrapper_i.sync_gpio_start.data_sync[1] ;
 wire \gpio_wrapper_i.sync_gpio_stop.data_sync[1] ;
 wire irq;
 wire \rsa_c[0] ;
 wire \rsa_c[1] ;
 wire \rsa_c[2] ;
 wire \rsa_c[3] ;
 wire \rsa_c[4] ;
 wire \rsa_c[5] ;
 wire \rsa_c[6] ;
 wire \rsa_c[7] ;
 wire \rsa_const[0] ;
 wire \rsa_const[1] ;
 wire \rsa_const[2] ;
 wire \rsa_const[3] ;
 wire \rsa_const[4] ;
 wire \rsa_const[5] ;
 wire \rsa_const[6] ;
 wire \rsa_const[7] ;
 wire \rsa_e[0] ;
 wire \rsa_e[1] ;
 wire \rsa_e[2] ;
 wire \rsa_e[3] ;
 wire \rsa_e[4] ;
 wire \rsa_e[5] ;
 wire \rsa_e[6] ;
 wire \rsa_e[7] ;
 wire \rsa_en_logic_i.state[0] ;
 wire \rsa_en_logic_i.state[1] ;
 wire \rsa_en_logic_i.state[2] ;
 wire \rsa_en_logic_i.state[3] ;
 wire \rsa_en_logic_i.state[4] ;
 wire \rsa_en_logic_i.state[5] ;
 wire \rsa_p[0] ;
 wire \rsa_p[1] ;
 wire \rsa_p[2] ;
 wire \rsa_p[3] ;
 wire \rsa_p[4] ;
 wire \rsa_p[5] ;
 wire \rsa_p[6] ;
 wire \rsa_p[7] ;
 wire \rsa_spi_wrapper_i.config_regs[0] ;
 wire \rsa_spi_wrapper_i.config_regs[10] ;
 wire \rsa_spi_wrapper_i.config_regs[11] ;
 wire \rsa_spi_wrapper_i.config_regs[12] ;
 wire \rsa_spi_wrapper_i.config_regs[13] ;
 wire \rsa_spi_wrapper_i.config_regs[14] ;
 wire \rsa_spi_wrapper_i.config_regs[15] ;
 wire \rsa_spi_wrapper_i.config_regs[1] ;
 wire \rsa_spi_wrapper_i.config_regs[2] ;
 wire \rsa_spi_wrapper_i.config_regs[32] ;
 wire \rsa_spi_wrapper_i.config_regs[33] ;
 wire \rsa_spi_wrapper_i.config_regs[34] ;
 wire \rsa_spi_wrapper_i.config_regs[35] ;
 wire \rsa_spi_wrapper_i.config_regs[36] ;
 wire \rsa_spi_wrapper_i.config_regs[37] ;
 wire \rsa_spi_wrapper_i.config_regs[38] ;
 wire \rsa_spi_wrapper_i.config_regs[39] ;
 wire \rsa_spi_wrapper_i.config_regs[3] ;
 wire \rsa_spi_wrapper_i.config_regs[48] ;
 wire \rsa_spi_wrapper_i.config_regs[49] ;
 wire \rsa_spi_wrapper_i.config_regs[4] ;
 wire \rsa_spi_wrapper_i.config_regs[50] ;
 wire \rsa_spi_wrapper_i.config_regs[51] ;
 wire \rsa_spi_wrapper_i.config_regs[52] ;
 wire \rsa_spi_wrapper_i.config_regs[53] ;
 wire \rsa_spi_wrapper_i.config_regs[54] ;
 wire \rsa_spi_wrapper_i.config_regs[55] ;
 wire \rsa_spi_wrapper_i.config_regs[56] ;
 wire \rsa_spi_wrapper_i.config_regs[57] ;
 wire \rsa_spi_wrapper_i.config_regs[58] ;
 wire \rsa_spi_wrapper_i.config_regs[59] ;
 wire \rsa_spi_wrapper_i.config_regs[5] ;
 wire \rsa_spi_wrapper_i.config_regs[60] ;
 wire \rsa_spi_wrapper_i.config_regs[61] ;
 wire \rsa_spi_wrapper_i.config_regs[62] ;
 wire \rsa_spi_wrapper_i.config_regs[63] ;
 wire \rsa_spi_wrapper_i.config_regs[6] ;
 wire \rsa_spi_wrapper_i.config_regs[7] ;
 wire \rsa_spi_wrapper_i.config_regs[8] ;
 wire \rsa_spi_wrapper_i.config_regs[9] ;
 wire \rsa_spi_wrapper_i.spi_clk ;
 wire \rsa_spi_wrapper_i.spi_cs_n ;
 wire \rsa_spi_wrapper_i.spi_miso ;
 wire \rsa_spi_wrapper_i.spi_mosi ;
 wire \rsa_spi_wrapper_i.spi_start_cmd_i.data_dly ;
 wire \rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[4] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[5] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[6] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[7] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o_vld ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[3] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[4] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[5] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[6] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ;
 wire \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ;
 wire \rsa_unit_i.P_i[0] ;
 wire \rsa_unit_i.P_i[1] ;
 wire \rsa_unit_i.P_i[2] ;
 wire \rsa_unit_i.P_i[3] ;
 wire \rsa_unit_i.P_i[4] ;
 wire \rsa_unit_i.P_i[5] ;
 wire \rsa_unit_i.P_i[6] ;
 wire \rsa_unit_i.P_i[7] ;
 wire \rsa_unit_i.P_i[8] ;
 wire \rsa_unit_i.P_i[9] ;
 wire \rsa_unit_i.R_i[0] ;
 wire \rsa_unit_i.R_i[1] ;
 wire \rsa_unit_i.R_i[2] ;
 wire \rsa_unit_i.R_i[3] ;
 wire \rsa_unit_i.R_i[4] ;
 wire \rsa_unit_i.R_i[5] ;
 wire \rsa_unit_i.R_i[6] ;
 wire \rsa_unit_i.R_i[7] ;
 wire \rsa_unit_i.R_i[8] ;
 wire \rsa_unit_i.R_i[9] ;
 wire \rsa_unit_i.mmm_multiply.A_bit ;
 wire \rsa_unit_i.mmm_multiply.adder2.fa_bit0.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[1].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[2].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[3].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[4].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[5].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[6].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[7].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.adder2.gen_fa[8].fa.HA1.a ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[1] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[2] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[3] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[4] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[5] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[6] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[7] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[8] ;
 wire \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[9] ;
 wire \rsa_unit_i.mmm_square.A_bit ;
 wire \rsa_unit_i.mmm_square.adder2.fa_bit0.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[1].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[2].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[3].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[4].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[5].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[6].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[7].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.adder2.gen_fa[8].fa.HA1.a ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[1] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[2] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[3] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[4] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[5] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[6] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[7] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[8] ;
 wire \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[9] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_rounds[0] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_rounds[1] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_rounds[2] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_rounds[3] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_steps[0] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_steps[1] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_steps[2] ;
 wire \rsa_unit_i.rsa_control_fsm.counter_steps[3] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[0] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[1] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[2] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[3] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[4] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[5] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[6] ;
 wire \rsa_unit_i.rsa_control_fsm.exp[7] ;
 wire \rsa_unit_i.rsa_control_fsm.increment_rounds ;
 wire \rsa_unit_i.rsa_control_fsm.load_exp ;
 wire \rsa_unit_i.rsa_control_fsm.state[0] ;
 wire \rsa_unit_i.rsa_control_fsm.state[10] ;
 wire \rsa_unit_i.rsa_control_fsm.state[11] ;
 wire \rsa_unit_i.rsa_control_fsm.state[1] ;
 wire \rsa_unit_i.rsa_control_fsm.state[2] ;
 wire \rsa_unit_i.rsa_control_fsm.state[3] ;
 wire \rsa_unit_i.rsa_control_fsm.state[6] ;
 wire \rsa_unit_i.rsa_control_fsm.state[7] ;
 wire \rsa_unit_i.rsa_control_fsm.state[8] ;
 wire \synchronizer_spi_clk_inst.data_sync[1] ;
 wire \synchronizer_spi_cs_n_inst.data_sync[1] ;
 wire \synchronizer_spi_mode_cpha.data_sync[1] ;
 wire \synchronizer_spi_mode_cpol.data_sync[1] ;
 wire \synchronizer_spi_mosi_inst.data_sync[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_1 _1595_ (.A(ena),
    .X(_1155_));
 sg13g2_inv_1 _1596_ (.Y(_1156_),
    .A(_1155_));
 sg13g2_inv_1 _1597_ (.Y(_1157_),
    .A(\gpio_wrapper_i.gpio_start_cmd_i.data_dly ));
 sg13g2_inv_1 _1598_ (.Y(_1158_),
    .A(\rsa_spi_wrapper_i.spi_start_cmd_i.data_dly ));
 sg13g2_a22oi_1 _1599_ (.Y(_1159_),
    .B1(\rsa_spi_wrapper_i.config_regs[8] ),
    .B2(_1158_),
    .A2(_1157_),
    .A1(\gpio_wrapper_i.gpio_start_cmd_i.data ));
 sg13g2_nor2_1 _1600_ (.A(_1156_),
    .B(_1159_),
    .Y(_1160_));
 sg13g2_a22oi_1 _1601_ (.Y(_1161_),
    .B1(\rsa_en_logic_i.state[3] ),
    .B2(_1160_),
    .A2(_1156_),
    .A1(\rsa_en_logic_i.state[2] ));
 sg13g2_inv_1 _1602_ (.Y(_0001_),
    .A(_1161_));
 sg13g2_buf_1 _1603_ (.A(_1155_),
    .X(_1162_));
 sg13g2_buf_1 _1604_ (.A(net111),
    .X(_1163_));
 sg13g2_nand2_1 _1605_ (.Y(_1164_),
    .A(net88),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_buf_1 _1606_ (.A(\rsa_spi_wrapper_i.spi_cs_n ),
    .X(_1165_));
 sg13g2_nor2b_1 _1607_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .B_N(_1165_),
    .Y(_1166_));
 sg13g2_buf_2 _1608_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ),
    .X(_1167_));
 sg13g2_nor3_2 _1609_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .B(_1167_),
    .C(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .Y(_1168_));
 sg13g2_mux2_1 _1610_ (.A0(_1166_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .S(_1168_),
    .X(_1169_));
 sg13g2_nand2_1 _1611_ (.Y(_1170_),
    .A(net88),
    .B(_1169_));
 sg13g2_nand2_1 _1612_ (.Y(_1171_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ),
    .B(_1170_));
 sg13g2_o21ai_1 _1613_ (.B1(_1171_),
    .Y(_0005_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ),
    .A2(_1164_));
 sg13g2_buf_8 _1614_ (.A(\rsa_unit_i.rsa_control_fsm.state[1] ),
    .X(_1172_));
 sg13g2_buf_2 _1615_ (.A(\rsa_en_logic_i.state[4] ),
    .X(_1173_));
 sg13g2_nand2b_1 _1616_ (.Y(_1174_),
    .B(_0056_),
    .A_N(\rsa_en_logic_i.state[1] ));
 sg13g2_nor2_2 _1617_ (.A(_1173_),
    .B(_1174_),
    .Y(_1175_));
 sg13g2_buf_2 _1618_ (.A(\rsa_unit_i.rsa_control_fsm.counter_steps[0] ),
    .X(_1176_));
 sg13g2_nand2b_1 _1619_ (.Y(_1177_),
    .B(_1176_),
    .A_N(\rsa_unit_i.rsa_control_fsm.counter_steps[1] ));
 sg13g2_nor2b_1 _1620_ (.A(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ),
    .B_N(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ),
    .Y(_1178_));
 sg13g2_nand2b_1 _1621_ (.Y(_1179_),
    .B(_1178_),
    .A_N(_1177_));
 sg13g2_inv_1 _1622_ (.Y(_1180_),
    .A(_1179_));
 sg13g2_or2_1 _1623_ (.X(_1181_),
    .B(\rsa_en_logic_i.state[5] ),
    .A(\rsa_en_logic_i.state[2] ));
 sg13g2_buf_1 _1624_ (.A(_1181_),
    .X(_1182_));
 sg13g2_or3_1 _1625_ (.A(\rsa_en_logic_i.state[1] ),
    .B(_1173_),
    .C(_1182_),
    .X(_1183_));
 sg13g2_buf_1 _1626_ (.A(_1183_),
    .X(_1184_));
 sg13g2_o21ai_1 _1627_ (.B1(net65),
    .Y(_1185_),
    .A1(_1175_),
    .A2(_1180_));
 sg13g2_nor3_2 _1628_ (.A(\rsa_en_logic_i.state[1] ),
    .B(_1173_),
    .C(_1182_),
    .Y(_1186_));
 sg13g2_buf_1 _1629_ (.A(_1186_),
    .X(_1187_));
 sg13g2_or2_1 _1630_ (.X(_1188_),
    .B(_1175_),
    .A(net64));
 sg13g2_nor2_1 _1631_ (.A(_0055_),
    .B(_1188_),
    .Y(_1189_));
 sg13g2_a21o_1 _1632_ (.A2(_1185_),
    .A1(_1172_),
    .B1(_1189_),
    .X(_0011_));
 sg13g2_inv_1 _1633_ (.Y(_1190_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_buf_1 _1634_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ),
    .X(_1191_));
 sg13g2_inv_1 _1635_ (.Y(_1192_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_nor4_2 _1636_ (.A(_1191_),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .C(_1192_),
    .Y(_1193_),
    .D(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ));
 sg13g2_o21ai_1 _1637_ (.B1(net111),
    .Y(_1194_),
    .A1(_1166_),
    .A2(_1193_));
 sg13g2_nand2_1 _1638_ (.Y(_1195_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ),
    .B(_1194_));
 sg13g2_o21ai_1 _1639_ (.B1(_1195_),
    .Y(_0008_),
    .A1(_1190_),
    .A2(_1164_));
 sg13g2_o21ai_1 _1640_ (.B1(net88),
    .Y(_1196_),
    .A1(_1165_),
    .A2(_1193_));
 sg13g2_inv_1 _1641_ (.Y(_1197_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_nand3b_1 _1642_ (.B(net111),
    .C(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0] ),
    .Y(_1198_),
    .A_N(_1165_));
 sg13g2_o21ai_1 _1643_ (.B1(_1198_),
    .Y(_1199_),
    .A1(_1197_),
    .A2(_1193_));
 sg13g2_a22oi_1 _1644_ (.Y(_1200_),
    .B1(_1199_),
    .B2(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .A2(_1196_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_inv_1 _1645_ (.Y(_0007_),
    .A(_1200_));
 sg13g2_buf_1 _1646_ (.A(net88),
    .X(_1201_));
 sg13g2_inv_1 _1647_ (.Y(_1202_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_nand3_1 _1648_ (.B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ),
    .C(_1193_),
    .A(_1162_),
    .Y(_1203_));
 sg13g2_buf_2 _1649_ (.A(_1203_),
    .X(_1204_));
 sg13g2_o21ai_1 _1650_ (.B1(_1204_),
    .Y(_0006_),
    .A1(net73),
    .A2(_1202_));
 sg13g2_nor2_1 _1651_ (.A(_1188_),
    .B(_1179_),
    .Y(_1205_));
 sg13g2_nand2_1 _1652_ (.Y(_1206_),
    .A(\rsa_unit_i.rsa_control_fsm.state[3] ),
    .B(_1205_));
 sg13g2_o21ai_1 _1653_ (.B1(_1206_),
    .Y(_0019_),
    .A1(_0054_),
    .A2(net65));
 sg13g2_buf_1 _1654_ (.A(eoc_rsa),
    .X(_1207_));
 sg13g2_nand2_1 _1655_ (.Y(_1208_),
    .A(net110),
    .B(net65));
 sg13g2_buf_1 _1656_ (.A(_1208_),
    .X(_1209_));
 sg13g2_inv_1 _1657_ (.Y(_1210_),
    .A(\rsa_unit_i.rsa_control_fsm.state[10] ));
 sg13g2_a22oi_1 _1658_ (.Y(_0009_),
    .B1(_1209_),
    .B2(_1210_),
    .A2(_1175_),
    .A1(_1182_));
 sg13g2_buf_1 _1659_ (.A(\rsa_unit_i.rsa_control_fsm.increment_rounds ),
    .X(_1211_));
 sg13g2_nor2_2 _1660_ (.A(net64),
    .B(_1175_),
    .Y(_1212_));
 sg13g2_inv_1 _1661_ (.Y(_1213_),
    .A(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ));
 sg13g2_buf_2 _1662_ (.A(\rsa_unit_i.rsa_control_fsm.counter_rounds[0] ),
    .X(_1214_));
 sg13g2_nand2b_1 _1663_ (.Y(_1215_),
    .B(_1214_),
    .A_N(\rsa_unit_i.rsa_control_fsm.counter_rounds[1] ));
 sg13g2_nor3_1 _1664_ (.A(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ),
    .B(_1213_),
    .C(_1215_),
    .Y(_1216_));
 sg13g2_nand3_1 _1665_ (.B(_1212_),
    .C(_1216_),
    .A(net109),
    .Y(_1217_));
 sg13g2_o21ai_1 _1666_ (.B1(_1217_),
    .Y(_0010_),
    .A1(_0055_),
    .A2(net65));
 sg13g2_inv_1 _1667_ (.Y(_1218_),
    .A(\gpio_wrapper_i.gpio_stop_cmd_i.data ));
 sg13g2_nand2b_1 _1668_ (.Y(_1219_),
    .B(\rsa_spi_wrapper_i.config_regs[9] ),
    .A_N(\rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly ));
 sg13g2_o21ai_1 _1669_ (.B1(_1219_),
    .Y(_1220_),
    .A1(_1218_),
    .A2(\gpio_wrapper_i.gpio_stop_cmd_i.data_dly ));
 sg13g2_buf_1 _1670_ (.A(_1220_),
    .X(_1221_));
 sg13g2_buf_1 _1671_ (.A(net111),
    .X(_1222_));
 sg13g2_nand2_1 _1672_ (.Y(_1223_),
    .A(\rsa_en_logic_i.state[5] ),
    .B(net87));
 sg13g2_o21ai_1 _1673_ (.B1(_1163_),
    .Y(_1224_),
    .A1(net110),
    .A2(_1221_));
 sg13g2_nand2_1 _1674_ (.Y(_1225_),
    .A(\rsa_en_logic_i.state[1] ),
    .B(_1224_));
 sg13g2_o21ai_1 _1675_ (.B1(_1225_),
    .Y(_0000_),
    .A1(_1221_),
    .A2(_1223_));
 sg13g2_buf_1 _1676_ (.A(net64),
    .X(_1226_));
 sg13g2_a22oi_1 _1677_ (.Y(_1227_),
    .B1(_1205_),
    .B2(\rsa_unit_i.rsa_control_fsm.state[8] ),
    .A2(net59),
    .A1(_1211_));
 sg13g2_inv_1 _1678_ (.Y(_0015_),
    .A(_1227_));
 sg13g2_a22oi_1 _1679_ (.Y(_1228_),
    .B1(_1212_),
    .B2(\rsa_unit_i.rsa_control_fsm.state[0] ),
    .A2(net59),
    .A1(\rsa_unit_i.rsa_control_fsm.state[6] ));
 sg13g2_inv_1 _1680_ (.Y(_0016_),
    .A(_1228_));
 sg13g2_buf_8 _1681_ (.A(\rsa_unit_i.rsa_control_fsm.state[7] ),
    .X(_1229_));
 sg13g2_a22oi_1 _1682_ (.Y(_1230_),
    .B1(_1205_),
    .B2(_1172_),
    .A2(net59),
    .A1(_1229_));
 sg13g2_inv_1 _1683_ (.Y(_0017_),
    .A(_1230_));
 sg13g2_a21oi_1 _1684_ (.A1(\rsa_unit_i.rsa_control_fsm.state[8] ),
    .A2(_1179_),
    .Y(_1231_),
    .B1(\rsa_unit_i.rsa_control_fsm.state[2] ));
 sg13g2_buf_1 _1685_ (.A(_0057_),
    .X(_1232_));
 sg13g2_nand2b_1 _1686_ (.Y(_1233_),
    .B(_1226_),
    .A_N(_1232_));
 sg13g2_o21ai_1 _1687_ (.B1(_1233_),
    .Y(_0018_),
    .A1(_1188_),
    .A2(_1231_));
 sg13g2_inv_1 _1688_ (.Y(_1234_),
    .A(net109));
 sg13g2_o21ai_1 _1689_ (.B1(_0054_),
    .Y(_1235_),
    .A1(_1234_),
    .A2(_1216_));
 sg13g2_a22oi_1 _1690_ (.Y(_1236_),
    .B1(_1212_),
    .B2(_1235_),
    .A2(_1226_),
    .A1(\rsa_unit_i.rsa_control_fsm.state[2] ));
 sg13g2_inv_1 _1691_ (.Y(_0012_),
    .A(_1236_));
 sg13g2_a22oi_1 _1692_ (.Y(_1237_),
    .B1(_1185_),
    .B2(\rsa_unit_i.rsa_control_fsm.state[3] ),
    .A2(_1212_),
    .A1(\rsa_unit_i.rsa_control_fsm.state[6] ));
 sg13g2_inv_1 _1693_ (.Y(_0013_),
    .A(_1237_));
 sg13g2_nand2_1 _1694_ (.Y(_1238_),
    .A(_1229_),
    .B(_1212_));
 sg13g2_o21ai_1 _1695_ (.B1(_1238_),
    .Y(_0014_),
    .A1(_0058_),
    .A2(_1184_));
 sg13g2_nand2_1 _1696_ (.Y(_1239_),
    .A(\rsa_en_logic_i.state[2] ),
    .B(net87));
 sg13g2_nand2_1 _1697_ (.Y(_1240_),
    .A(\rsa_en_logic_i.state[5] ),
    .B(_1156_));
 sg13g2_o21ai_1 _1698_ (.B1(_1240_),
    .Y(_0004_),
    .A1(_1221_),
    .A2(_1239_));
 sg13g2_nand3_1 _1699_ (.B(net87),
    .C(net110),
    .A(\rsa_en_logic_i.state[1] ),
    .Y(_1241_));
 sg13g2_nand2_1 _1700_ (.Y(_1242_),
    .A(_1173_),
    .B(_1156_));
 sg13g2_o21ai_1 _1701_ (.B1(_1242_),
    .Y(_0003_),
    .A1(_1221_),
    .A2(_1241_));
 sg13g2_inv_1 _1702_ (.Y(_1243_),
    .A(_1160_));
 sg13g2_nor2_1 _1703_ (.A(_1173_),
    .B(\rsa_en_logic_i.state[0] ),
    .Y(_1244_));
 sg13g2_o21ai_1 _1704_ (.B1(_1221_),
    .Y(_1245_),
    .A1(\rsa_en_logic_i.state[2] ),
    .A2(_1174_));
 sg13g2_nand2_1 _1705_ (.Y(_1246_),
    .A(_1244_),
    .B(_1245_));
 sg13g2_a22oi_1 _1706_ (.Y(_1247_),
    .B1(_1246_),
    .B2(net73),
    .A2(_1243_),
    .A1(\rsa_en_logic_i.state[3] ));
 sg13g2_inv_1 _1707_ (.Y(_0002_),
    .A(_1247_));
 sg13g2_nand2_1 _1708_ (.Y(_1248_),
    .A(net73),
    .B(\gpio_wrapper_i.gpio_start_cmd_i.data ));
 sg13g2_o21ai_1 _1709_ (.B1(_1248_),
    .Y(_0122_),
    .A1(net73),
    .A2(_1157_));
 sg13g2_buf_1 _1710_ (.A(net88),
    .X(_1249_));
 sg13g2_mux2_1 _1711_ (.A0(\gpio_wrapper_i.gpio_stop_cmd_i.data_dly ),
    .A1(\gpio_wrapper_i.gpio_stop_cmd_i.data ),
    .S(net72),
    .X(_0123_));
 sg13g2_mux2_1 _1712_ (.A0(\gpio_wrapper_i.sync_gpio_start.data_sync[1] ),
    .A1(net2),
    .S(net72),
    .X(_0124_));
 sg13g2_mux2_1 _1713_ (.A0(\gpio_wrapper_i.gpio_start_cmd_i.data ),
    .A1(\gpio_wrapper_i.sync_gpio_start.data_sync[1] ),
    .S(_1249_),
    .X(_0125_));
 sg13g2_mux2_1 _1714_ (.A0(\gpio_wrapper_i.sync_gpio_stop.data_sync[1] ),
    .A1(net3),
    .S(_1249_),
    .X(_0126_));
 sg13g2_nand2_1 _1715_ (.Y(_1250_),
    .A(net73),
    .B(\gpio_wrapper_i.sync_gpio_stop.data_sync[1] ));
 sg13g2_o21ai_1 _1716_ (.B1(_1250_),
    .Y(_0127_),
    .A1(_1201_),
    .A2(_1218_));
 sg13g2_a21oi_1 _1717_ (.A1(_1173_),
    .A2(net111),
    .Y(_1251_),
    .B1(irq));
 sg13g2_a21oi_1 _1718_ (.A1(net88),
    .A2(_1221_),
    .Y(_1252_),
    .B1(_1251_));
 sg13g2_nor2b_1 _1719_ (.A(_1160_),
    .B_N(_1252_),
    .Y(_0128_));
 sg13g2_nand2_1 _1720_ (.Y(_1253_),
    .A(net73),
    .B(\rsa_spi_wrapper_i.config_regs[8] ));
 sg13g2_o21ai_1 _1721_ (.B1(_1253_),
    .Y(_0129_),
    .A1(net73),
    .A2(_1158_));
 sg13g2_mux2_1 _1722_ (.A0(\rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly ),
    .A1(\rsa_spi_wrapper_i.config_regs[9] ),
    .S(net72),
    .X(_0130_));
 sg13g2_buf_1 _1723_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[0] ),
    .X(_1254_));
 sg13g2_buf_1 _1724_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[0] ),
    .X(_1255_));
 sg13g2_buf_1 _1725_ (.A(net106),
    .X(_1256_));
 sg13g2_buf_1 _1726_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[1] ),
    .X(_1257_));
 sg13g2_buf_1 _1727_ (.A(net105),
    .X(_1258_));
 sg13g2_buf_1 _1728_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[2] ),
    .X(_1259_));
 sg13g2_buf_1 _1729_ (.A(_1259_),
    .X(_1260_));
 sg13g2_nand2_2 _1730_ (.Y(_1261_),
    .A(_1155_),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o_vld ));
 sg13g2_nor4_1 _1731_ (.A(net86),
    .B(_1258_),
    .C(net84),
    .D(_1261_),
    .Y(_1262_));
 sg13g2_buf_4 _1732_ (.X(_1263_),
    .A(_1262_));
 sg13g2_mux2_1 _1733_ (.A0(\rsa_spi_wrapper_i.config_regs[0] ),
    .A1(net107),
    .S(_1263_),
    .X(_0131_));
 sg13g2_buf_1 _1734_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[1] ),
    .X(_1264_));
 sg13g2_mux2_1 _1735_ (.A0(\rsa_spi_wrapper_i.config_regs[1] ),
    .A1(net104),
    .S(_1263_),
    .X(_0132_));
 sg13g2_buf_1 _1736_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[2] ),
    .X(_1265_));
 sg13g2_mux2_1 _1737_ (.A0(\rsa_spi_wrapper_i.config_regs[2] ),
    .A1(net103),
    .S(_1263_),
    .X(_0133_));
 sg13g2_buf_1 _1738_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[3] ),
    .X(_1266_));
 sg13g2_mux2_1 _1739_ (.A0(\rsa_spi_wrapper_i.config_regs[3] ),
    .A1(net102),
    .S(_1263_),
    .X(_0134_));
 sg13g2_buf_1 _1740_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[4] ),
    .X(_1267_));
 sg13g2_mux2_1 _1741_ (.A0(\rsa_spi_wrapper_i.config_regs[4] ),
    .A1(net101),
    .S(_1263_),
    .X(_0135_));
 sg13g2_buf_1 _1742_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[5] ),
    .X(_1268_));
 sg13g2_mux2_1 _1743_ (.A0(\rsa_spi_wrapper_i.config_regs[5] ),
    .A1(net100),
    .S(_1263_),
    .X(_0136_));
 sg13g2_buf_1 _1744_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[6] ),
    .X(_1269_));
 sg13g2_mux2_1 _1745_ (.A0(\rsa_spi_wrapper_i.config_regs[6] ),
    .A1(net99),
    .S(_1263_),
    .X(_0137_));
 sg13g2_buf_1 _1746_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[7] ),
    .X(_1270_));
 sg13g2_mux2_1 _1747_ (.A0(\rsa_spi_wrapper_i.config_regs[7] ),
    .A1(net98),
    .S(_1263_),
    .X(_0138_));
 sg13g2_buf_1 _1748_ (.A(_0053_),
    .X(_1271_));
 sg13g2_nor2b_1 _1749_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[1] ),
    .B_N(_1271_),
    .Y(_1272_));
 sg13g2_and2_1 _1750_ (.A(_1255_),
    .B(_1272_),
    .X(_1273_));
 sg13g2_buf_2 _1751_ (.A(_1273_),
    .X(_1274_));
 sg13g2_nor2b_1 _1752_ (.A(_1261_),
    .B_N(_1274_),
    .Y(_1275_));
 sg13g2_buf_4 _1753_ (.X(_1276_),
    .A(_1275_));
 sg13g2_mux2_1 _1754_ (.A0(\rsa_spi_wrapper_i.config_regs[8] ),
    .A1(net107),
    .S(_1276_),
    .X(_0139_));
 sg13g2_mux2_1 _1755_ (.A0(\rsa_spi_wrapper_i.config_regs[9] ),
    .A1(net104),
    .S(_1276_),
    .X(_0140_));
 sg13g2_mux2_1 _1756_ (.A0(\rsa_spi_wrapper_i.config_regs[10] ),
    .A1(net103),
    .S(_1276_),
    .X(_0141_));
 sg13g2_mux2_1 _1757_ (.A0(\rsa_spi_wrapper_i.config_regs[11] ),
    .A1(net102),
    .S(_1276_),
    .X(_0142_));
 sg13g2_mux2_1 _1758_ (.A0(\rsa_spi_wrapper_i.config_regs[12] ),
    .A1(net101),
    .S(_1276_),
    .X(_0143_));
 sg13g2_mux2_1 _1759_ (.A0(\rsa_spi_wrapper_i.config_regs[13] ),
    .A1(net100),
    .S(_1276_),
    .X(_0144_));
 sg13g2_mux2_1 _1760_ (.A0(\rsa_spi_wrapper_i.config_regs[14] ),
    .A1(net99),
    .S(_1276_),
    .X(_0145_));
 sg13g2_mux2_1 _1761_ (.A0(\rsa_spi_wrapper_i.config_regs[15] ),
    .A1(net98),
    .S(_1276_),
    .X(_0146_));
 sg13g2_inv_2 _1762_ (.Y(_1277_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[1] ));
 sg13g2_nor4_1 _1763_ (.A(net86),
    .B(_1277_),
    .C(net84),
    .D(_1261_),
    .Y(_1278_));
 sg13g2_buf_1 _1764_ (.A(_1278_),
    .X(_1279_));
 sg13g2_mux2_1 _1765_ (.A0(\rsa_p[0] ),
    .A1(net107),
    .S(net63),
    .X(_0147_));
 sg13g2_buf_2 _1766_ (.A(\rsa_p[1] ),
    .X(_1280_));
 sg13g2_inv_1 _1767_ (.Y(_1281_),
    .A(_1280_));
 sg13g2_nand2_1 _1768_ (.Y(_1282_),
    .A(net104),
    .B(net63));
 sg13g2_o21ai_1 _1769_ (.B1(_1282_),
    .Y(_0148_),
    .A1(_1281_),
    .A2(net63));
 sg13g2_mux2_1 _1770_ (.A0(\rsa_p[2] ),
    .A1(net103),
    .S(net63),
    .X(_0149_));
 sg13g2_mux2_1 _1771_ (.A0(\rsa_p[3] ),
    .A1(net102),
    .S(net63),
    .X(_0150_));
 sg13g2_mux2_1 _1772_ (.A0(\rsa_p[4] ),
    .A1(net101),
    .S(_1279_),
    .X(_0151_));
 sg13g2_mux2_1 _1773_ (.A0(\rsa_p[5] ),
    .A1(net100),
    .S(net63),
    .X(_0152_));
 sg13g2_mux2_1 _1774_ (.A0(\rsa_p[6] ),
    .A1(net99),
    .S(net63),
    .X(_0153_));
 sg13g2_mux2_1 _1775_ (.A0(\rsa_p[7] ),
    .A1(net98),
    .S(net63),
    .X(_0154_));
 sg13g2_nand2_1 _1776_ (.Y(_1283_),
    .A(net106),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[1] ));
 sg13g2_nor3_1 _1777_ (.A(_1260_),
    .B(_1261_),
    .C(_1283_),
    .Y(_1284_));
 sg13g2_buf_4 _1778_ (.X(_1285_),
    .A(_1284_));
 sg13g2_mux2_1 _1779_ (.A0(\rsa_e[0] ),
    .A1(_1254_),
    .S(_1285_),
    .X(_0155_));
 sg13g2_mux2_1 _1780_ (.A0(\rsa_e[1] ),
    .A1(net104),
    .S(_1285_),
    .X(_0156_));
 sg13g2_mux2_1 _1781_ (.A0(\rsa_e[2] ),
    .A1(net103),
    .S(_1285_),
    .X(_0157_));
 sg13g2_mux2_1 _1782_ (.A0(\rsa_e[3] ),
    .A1(net102),
    .S(_1285_),
    .X(_0158_));
 sg13g2_mux2_1 _1783_ (.A0(\rsa_e[4] ),
    .A1(net101),
    .S(_1285_),
    .X(_0159_));
 sg13g2_mux2_1 _1784_ (.A0(\rsa_e[5] ),
    .A1(net100),
    .S(_1285_),
    .X(_0160_));
 sg13g2_mux2_1 _1785_ (.A0(\rsa_e[6] ),
    .A1(net99),
    .S(_1285_),
    .X(_0161_));
 sg13g2_mux2_1 _1786_ (.A0(\rsa_e[7] ),
    .A1(net98),
    .S(_1285_),
    .X(_0162_));
 sg13g2_buf_8 _1787_ (.A(\rsa_spi_wrapper_i.config_regs[32] ),
    .X(_1286_));
 sg13g2_buf_1 _1788_ (.A(_1286_),
    .X(_1287_));
 sg13g2_inv_1 _1789_ (.Y(_1288_),
    .A(net106));
 sg13g2_buf_1 _1790_ (.A(_1288_),
    .X(_1289_));
 sg13g2_nand2_1 _1791_ (.Y(_1290_),
    .A(net71),
    .B(net84));
 sg13g2_nor3_1 _1792_ (.A(net85),
    .B(_1261_),
    .C(_1290_),
    .Y(_1291_));
 sg13g2_buf_1 _1793_ (.A(_1291_),
    .X(_1292_));
 sg13g2_mux2_1 _1794_ (.A0(net83),
    .A1(net107),
    .S(net47),
    .X(_0163_));
 sg13g2_inv_2 _1795_ (.Y(_1293_),
    .A(\rsa_spi_wrapper_i.config_regs[33] ));
 sg13g2_nand2_1 _1796_ (.Y(_1294_),
    .A(net104),
    .B(net47));
 sg13g2_o21ai_1 _1797_ (.B1(_1294_),
    .Y(_0164_),
    .A1(_1293_),
    .A2(_1292_));
 sg13g2_mux2_1 _1798_ (.A0(\rsa_spi_wrapper_i.config_regs[34] ),
    .A1(net103),
    .S(net47),
    .X(_0165_));
 sg13g2_mux2_1 _1799_ (.A0(\rsa_spi_wrapper_i.config_regs[35] ),
    .A1(net102),
    .S(net47),
    .X(_0166_));
 sg13g2_mux2_1 _1800_ (.A0(\rsa_spi_wrapper_i.config_regs[36] ),
    .A1(net101),
    .S(net47),
    .X(_0167_));
 sg13g2_mux2_1 _1801_ (.A0(\rsa_spi_wrapper_i.config_regs[37] ),
    .A1(net100),
    .S(net47),
    .X(_0168_));
 sg13g2_mux2_1 _1802_ (.A0(\rsa_spi_wrapper_i.config_regs[38] ),
    .A1(net99),
    .S(net47),
    .X(_0169_));
 sg13g2_mux2_1 _1803_ (.A0(\rsa_spi_wrapper_i.config_regs[39] ),
    .A1(net98),
    .S(net47),
    .X(_0170_));
 sg13g2_buf_1 _1804_ (.A(_1271_),
    .X(_1295_));
 sg13g2_nor4_1 _1805_ (.A(_1289_),
    .B(net85),
    .C(net82),
    .D(_1261_),
    .Y(_1296_));
 sg13g2_buf_1 _1806_ (.A(_1296_),
    .X(_1297_));
 sg13g2_mux2_1 _1807_ (.A0(\rsa_const[0] ),
    .A1(net107),
    .S(net58),
    .X(_0171_));
 sg13g2_mux2_1 _1808_ (.A0(\rsa_const[1] ),
    .A1(_1264_),
    .S(net58),
    .X(_0172_));
 sg13g2_inv_1 _1809_ (.Y(_1298_),
    .A(\rsa_const[2] ));
 sg13g2_nand2_1 _1810_ (.Y(_1299_),
    .A(net103),
    .B(net58));
 sg13g2_o21ai_1 _1811_ (.B1(_1299_),
    .Y(_0173_),
    .A1(_1298_),
    .A2(net58));
 sg13g2_mux2_1 _1812_ (.A0(\rsa_const[3] ),
    .A1(_1266_),
    .S(net58),
    .X(_0174_));
 sg13g2_mux2_1 _1813_ (.A0(\rsa_const[4] ),
    .A1(_1267_),
    .S(net58),
    .X(_0175_));
 sg13g2_mux2_1 _1814_ (.A0(\rsa_const[5] ),
    .A1(net100),
    .S(_1297_),
    .X(_0176_));
 sg13g2_mux2_1 _1815_ (.A0(\rsa_const[6] ),
    .A1(_1269_),
    .S(net58),
    .X(_0177_));
 sg13g2_mux2_1 _1816_ (.A0(\rsa_const[7] ),
    .A1(net98),
    .S(net58),
    .X(_0178_));
 sg13g2_nor3_2 _1817_ (.A(net106),
    .B(_1277_),
    .C(_1271_),
    .Y(_1300_));
 sg13g2_nor2b_1 _1818_ (.A(_1261_),
    .B_N(_1300_),
    .Y(_1301_));
 sg13g2_buf_4 _1819_ (.X(_1302_),
    .A(_1301_));
 sg13g2_mux2_1 _1820_ (.A0(\rsa_spi_wrapper_i.config_regs[48] ),
    .A1(net107),
    .S(_1302_),
    .X(_0179_));
 sg13g2_mux2_1 _1821_ (.A0(\rsa_spi_wrapper_i.config_regs[49] ),
    .A1(net104),
    .S(_1302_),
    .X(_0180_));
 sg13g2_mux2_1 _1822_ (.A0(\rsa_spi_wrapper_i.config_regs[50] ),
    .A1(net103),
    .S(_1302_),
    .X(_0181_));
 sg13g2_mux2_1 _1823_ (.A0(\rsa_spi_wrapper_i.config_regs[51] ),
    .A1(net102),
    .S(_1302_),
    .X(_0182_));
 sg13g2_mux2_1 _1824_ (.A0(\rsa_spi_wrapper_i.config_regs[52] ),
    .A1(net101),
    .S(_1302_),
    .X(_0183_));
 sg13g2_mux2_1 _1825_ (.A0(\rsa_spi_wrapper_i.config_regs[53] ),
    .A1(net100),
    .S(_1302_),
    .X(_0184_));
 sg13g2_mux2_1 _1826_ (.A0(\rsa_spi_wrapper_i.config_regs[54] ),
    .A1(net99),
    .S(_1302_),
    .X(_0185_));
 sg13g2_mux2_1 _1827_ (.A0(\rsa_spi_wrapper_i.config_regs[55] ),
    .A1(net98),
    .S(_1302_),
    .X(_0186_));
 sg13g2_nand3_1 _1828_ (.B(net85),
    .C(_1260_),
    .A(_1256_),
    .Y(_1303_));
 sg13g2_nor2_1 _1829_ (.A(_1261_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_buf_4 _1830_ (.X(_1305_),
    .A(_1304_));
 sg13g2_mux2_1 _1831_ (.A0(\rsa_spi_wrapper_i.config_regs[56] ),
    .A1(net107),
    .S(_1305_),
    .X(_0187_));
 sg13g2_mux2_1 _1832_ (.A0(\rsa_spi_wrapper_i.config_regs[57] ),
    .A1(net104),
    .S(_1305_),
    .X(_0188_));
 sg13g2_mux2_1 _1833_ (.A0(\rsa_spi_wrapper_i.config_regs[58] ),
    .A1(_1265_),
    .S(_1305_),
    .X(_0189_));
 sg13g2_mux2_1 _1834_ (.A0(\rsa_spi_wrapper_i.config_regs[59] ),
    .A1(net102),
    .S(_1305_),
    .X(_0190_));
 sg13g2_mux2_1 _1835_ (.A0(\rsa_spi_wrapper_i.config_regs[60] ),
    .A1(net101),
    .S(_1305_),
    .X(_0191_));
 sg13g2_mux2_1 _1836_ (.A0(\rsa_spi_wrapper_i.config_regs[61] ),
    .A1(_1268_),
    .S(_1305_),
    .X(_0192_));
 sg13g2_mux2_1 _1837_ (.A0(\rsa_spi_wrapper_i.config_regs[62] ),
    .A1(net99),
    .S(_1305_),
    .X(_0193_));
 sg13g2_mux2_1 _1838_ (.A0(\rsa_spi_wrapper_i.config_regs[63] ),
    .A1(_1270_),
    .S(_1305_),
    .X(_0194_));
 sg13g2_mux2_1 _1839_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .A1(net86),
    .S(_1204_),
    .X(_0195_));
 sg13g2_mux2_1 _1840_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .A1(net85),
    .S(_1204_),
    .X(_0196_));
 sg13g2_mux2_1 _1841_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .A1(net84),
    .S(_1204_),
    .X(_0197_));
 sg13g2_buf_2 _1842_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[3] ),
    .X(_1306_));
 sg13g2_buf_1 _1843_ (.A(_1306_),
    .X(_1307_));
 sg13g2_mux2_1 _1844_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .A1(_1307_),
    .S(_1204_),
    .X(_0198_));
 sg13g2_nand3_1 _1845_ (.B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ),
    .C(_1193_),
    .A(_1162_),
    .Y(_1308_));
 sg13g2_buf_1 _1846_ (.A(_1308_),
    .X(_1309_));
 sg13g2_mux2_1 _1847_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .A1(net107),
    .S(net62),
    .X(_0199_));
 sg13g2_mux2_1 _1848_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .A1(net104),
    .S(net62),
    .X(_0200_));
 sg13g2_mux2_1 _1849_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .A1(net103),
    .S(net62),
    .X(_0201_));
 sg13g2_mux2_1 _1850_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .A1(net102),
    .S(net62),
    .X(_0202_));
 sg13g2_mux2_1 _1851_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .A1(net101),
    .S(net62),
    .X(_0203_));
 sg13g2_mux2_1 _1852_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .A1(net100),
    .S(net62),
    .X(_0204_));
 sg13g2_mux2_1 _1853_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .A1(net99),
    .S(net62),
    .X(_0205_));
 sg13g2_mux2_1 _1854_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .A1(net98),
    .S(net62),
    .X(_0206_));
 sg13g2_nand2_1 _1855_ (.Y(_1310_),
    .A(_1156_),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o_vld ));
 sg13g2_o21ai_1 _1856_ (.B1(_1310_),
    .Y(_0207_),
    .A1(_1190_),
    .A2(_1309_));
 sg13g2_mux2_1 _1857_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ),
    .S(_1204_),
    .X(_0208_));
 sg13g2_inv_1 _1858_ (.Y(_1311_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ));
 sg13g2_nand2_1 _1859_ (.Y(_1312_),
    .A(_1165_),
    .B(_1155_));
 sg13g2_o21ai_1 _1860_ (.B1(_1312_),
    .Y(_0209_),
    .A1(_1311_),
    .A2(_1201_));
 sg13g2_mux2_1 _1861_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .A1(\rsa_spi_wrapper_i.spi_clk ),
    .S(net72),
    .X(_0210_));
 sg13g2_nor2b_1 _1862_ (.A(\rsa_spi_wrapper_i.spi_clk ),
    .B_N(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .Y(_1313_));
 sg13g2_nor2b_1 _1863_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ),
    .B_N(\rsa_spi_wrapper_i.spi_clk ),
    .Y(_1314_));
 sg13g2_xnor2_1 _1864_ (.Y(_1315_),
    .A(cpha_sync),
    .B(cpol_sync));
 sg13g2_mux2_1 _1865_ (.A0(_1313_),
    .A1(_1314_),
    .S(_1315_),
    .X(_1316_));
 sg13g2_and3_1 _1866_ (.X(_1317_),
    .A(_0052_),
    .B(_1155_),
    .C(_1316_));
 sg13g2_buf_1 _1867_ (.A(_1317_),
    .X(_1318_));
 sg13g2_buf_1 _1868_ (.A(_1318_),
    .X(_1319_));
 sg13g2_mux2_1 _1869_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .A1(\rsa_spi_wrapper_i.spi_mosi ),
    .S(net57),
    .X(_0211_));
 sg13g2_mux2_1 _1870_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ),
    .S(net57),
    .X(_0212_));
 sg13g2_mux2_1 _1871_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ),
    .S(net57),
    .X(_0213_));
 sg13g2_mux2_1 _1872_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ),
    .S(net57),
    .X(_0214_));
 sg13g2_mux2_1 _1873_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ),
    .S(net57),
    .X(_0215_));
 sg13g2_mux2_1 _1874_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ),
    .S(net57),
    .X(_0216_));
 sg13g2_mux2_1 _1875_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ),
    .S(net57),
    .X(_0217_));
 sg13g2_mux2_1 _1876_ (.A0(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ),
    .S(net57),
    .X(_0218_));
 sg13g2_xnor2_1 _1877_ (.Y(_1320_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .B(_1319_));
 sg13g2_a21oi_1 _1878_ (.A1(net73),
    .A2(_1193_),
    .Y(_0219_),
    .B1(_1320_));
 sg13g2_and2_1 _1879_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .B(_1318_),
    .X(_1321_));
 sg13g2_buf_1 _1880_ (.A(_1321_),
    .X(_1322_));
 sg13g2_xor2_1 _1881_ (.B(_1322_),
    .A(_1191_),
    .X(_0220_));
 sg13g2_nand2_1 _1882_ (.Y(_1323_),
    .A(_1191_),
    .B(_1322_));
 sg13g2_xnor2_1 _1883_ (.Y(_0221_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .B(_1323_));
 sg13g2_a21oi_1 _1884_ (.A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .A2(_1322_),
    .Y(_1324_),
    .B1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_nor2_1 _1885_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .Y(_1325_));
 sg13g2_a21oi_1 _1886_ (.A1(net88),
    .A2(_1325_),
    .Y(_1326_),
    .B1(_1192_));
 sg13g2_nand4_1 _1887_ (.B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ),
    .C(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ),
    .A(_1191_),
    .Y(_1327_),
    .D(_1322_));
 sg13g2_o21ai_1 _1888_ (.B1(_1327_),
    .Y(_1328_),
    .A1(_1191_),
    .A2(_1326_));
 sg13g2_nor2_1 _1889_ (.A(_1324_),
    .B(_1328_),
    .Y(_0222_));
 sg13g2_nor3_2 _1890_ (.A(_1257_),
    .B(net84),
    .C(_1274_),
    .Y(_1329_));
 sg13g2_buf_1 _1891_ (.A(_1329_),
    .X(_1330_));
 sg13g2_nand2b_1 _1892_ (.Y(_1331_),
    .B(_1306_),
    .A_N(_0061_));
 sg13g2_o21ai_1 _1893_ (.B1(_1331_),
    .Y(_1332_),
    .A1(_0059_),
    .A2(net81));
 sg13g2_nor2_1 _1894_ (.A(_1277_),
    .B(_1271_),
    .Y(_1333_));
 sg13g2_nor2b_2 _1895_ (.A(_1257_),
    .B_N(_1259_),
    .Y(_1334_));
 sg13g2_a21oi_1 _1896_ (.A1(\rsa_c[0] ),
    .A2(_1333_),
    .Y(_1335_),
    .B1(_1334_));
 sg13g2_or2_1 _1897_ (.X(_1336_),
    .B(_1335_),
    .A(net86));
 sg13g2_and2_1 _1898_ (.A(_1306_),
    .B(_1303_),
    .X(_1337_));
 sg13g2_and2_1 _1899_ (.A(net105),
    .B(_1259_),
    .X(_1338_));
 sg13g2_mux2_1 _1900_ (.A0(\rsa_const[0] ),
    .A1(\rsa_spi_wrapper_i.config_regs[8] ),
    .S(net82),
    .X(_1339_));
 sg13g2_a22oi_1 _1901_ (.Y(_1340_),
    .B1(_1339_),
    .B2(_1277_),
    .A2(_1338_),
    .A1(\rsa_spi_wrapper_i.config_regs[56] ));
 sg13g2_nor2_1 _1902_ (.A(_1277_),
    .B(_1259_),
    .Y(_1341_));
 sg13g2_buf_2 _1903_ (.A(_0060_),
    .X(_1342_));
 sg13g2_inv_1 _1904_ (.Y(_1343_),
    .A(_1342_));
 sg13g2_a22oi_1 _1905_ (.Y(_1344_),
    .B1(_1334_),
    .B2(_1343_),
    .A2(_1341_),
    .A1(\rsa_p[0] ));
 sg13g2_mux2_1 _1906_ (.A0(_1340_),
    .A1(_1344_),
    .S(net71),
    .X(_1345_));
 sg13g2_nor2_2 _1907_ (.A(net84),
    .B(_1283_),
    .Y(_1346_));
 sg13g2_a221oi_1 _1908_ (.B2(\rsa_spi_wrapper_i.config_regs[48] ),
    .C1(_1306_),
    .B1(_1300_),
    .A1(\rsa_e[0] ),
    .Y(_1347_),
    .A2(_1346_));
 sg13g2_a221oi_1 _1909_ (.B2(_1347_),
    .C1(net46),
    .B1(_1345_),
    .A1(_1336_),
    .Y(_1348_),
    .A2(_1337_));
 sg13g2_a21oi_1 _1910_ (.A1(_1330_),
    .A2(_1332_),
    .Y(_1349_),
    .B1(_1348_));
 sg13g2_inv_1 _1911_ (.Y(_1350_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ));
 sg13g2_nand2b_1 _1912_ (.Y(_1351_),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ),
    .A_N(_1165_));
 sg13g2_and2_1 _1913_ (.A(net111),
    .B(_1168_),
    .X(_1352_));
 sg13g2_nand4_1 _1914_ (.B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ),
    .C(_1351_),
    .A(_1350_),
    .Y(_1353_),
    .D(_1352_));
 sg13g2_mux2_1 _1915_ (.A0(_1314_),
    .A1(_1313_),
    .S(_1315_),
    .X(_1354_));
 sg13g2_nand2_1 _1916_ (.Y(_1355_),
    .A(_0052_),
    .B(_1354_));
 sg13g2_nand3_1 _1917_ (.B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ),
    .C(_1168_),
    .A(_1350_),
    .Y(_1356_));
 sg13g2_buf_1 _1918_ (.A(_1356_),
    .X(_1357_));
 sg13g2_nand3_1 _1919_ (.B(_1351_),
    .C(_1357_),
    .A(_1355_),
    .Y(_1358_));
 sg13g2_nand2_2 _1920_ (.Y(_1359_),
    .A(net111),
    .B(_1358_));
 sg13g2_nand2_1 _1921_ (.Y(_1360_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[0] ),
    .B(_1359_));
 sg13g2_o21ai_1 _1922_ (.B1(_1360_),
    .Y(_0223_),
    .A1(_1349_),
    .A2(_1353_));
 sg13g2_buf_1 _1923_ (.A(_1357_),
    .X(_1361_));
 sg13g2_buf_1 _1924_ (.A(_0064_),
    .X(_1362_));
 sg13g2_inv_1 _1925_ (.Y(_1363_),
    .A(net97));
 sg13g2_a22oi_1 _1926_ (.Y(_1364_),
    .B1(_1334_),
    .B2(_1363_),
    .A2(_1341_),
    .A1(_1280_));
 sg13g2_a221oi_1 _1927_ (.B2(\rsa_spi_wrapper_i.config_regs[57] ),
    .C1(net71),
    .B1(_1338_),
    .A1(\rsa_spi_wrapper_i.config_regs[9] ),
    .Y(_1365_),
    .A2(_1272_));
 sg13g2_a21oi_1 _1928_ (.A1(net71),
    .A2(_1364_),
    .Y(_1366_),
    .B1(_1365_));
 sg13g2_nor2_1 _1929_ (.A(_1288_),
    .B(net105),
    .Y(_1367_));
 sg13g2_nor2_2 _1930_ (.A(net106),
    .B(_1277_),
    .Y(_1368_));
 sg13g2_a22oi_1 _1931_ (.Y(_1369_),
    .B1(_1368_),
    .B2(\rsa_spi_wrapper_i.config_regs[49] ),
    .A2(_1367_),
    .A1(\rsa_const[1] ));
 sg13g2_nand2_1 _1932_ (.Y(_1370_),
    .A(\rsa_e[1] ),
    .B(_1346_));
 sg13g2_o21ai_1 _1933_ (.B1(_1370_),
    .Y(_1371_),
    .A1(net82),
    .A2(_1369_));
 sg13g2_nor3_1 _1934_ (.A(_1329_),
    .B(_1366_),
    .C(_1371_),
    .Y(_1372_));
 sg13g2_a21o_1 _1935_ (.A2(net46),
    .A1(_0063_),
    .B1(_1372_),
    .X(_1373_));
 sg13g2_nor2b_1 _1936_ (.A(net82),
    .B_N(\rsa_c[1] ),
    .Y(_1374_));
 sg13g2_nor2_1 _1937_ (.A(net105),
    .B(net82),
    .Y(_1375_));
 sg13g2_nor2b_1 _1938_ (.A(_1375_),
    .B_N(_1306_),
    .Y(_1376_));
 sg13g2_o21ai_1 _1939_ (.B1(_1376_),
    .Y(_1377_),
    .A1(net86),
    .A2(_1374_));
 sg13g2_o21ai_1 _1940_ (.B1(_1377_),
    .Y(_1378_),
    .A1(net81),
    .A2(_1373_));
 sg13g2_nand2_1 _1941_ (.Y(_1379_),
    .A(_0062_),
    .B(_1357_));
 sg13g2_o21ai_1 _1942_ (.B1(_1379_),
    .Y(_1380_),
    .A1(net56),
    .A2(_1378_));
 sg13g2_nand3_1 _1943_ (.B(_1351_),
    .C(_1358_),
    .A(net111),
    .Y(_1381_));
 sg13g2_buf_2 _1944_ (.A(_1381_),
    .X(_1382_));
 sg13g2_nand2_1 _1945_ (.Y(_1383_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[1] ),
    .B(_1359_));
 sg13g2_o21ai_1 _1946_ (.B1(_1383_),
    .Y(_0224_),
    .A1(_1380_),
    .A2(_1382_));
 sg13g2_nand2b_1 _1947_ (.Y(_1384_),
    .B(\rsa_c[2] ),
    .A_N(net82));
 sg13g2_a22oi_1 _1948_ (.Y(_1385_),
    .B1(_1368_),
    .B2(_1384_),
    .A2(_1290_),
    .A1(_1277_));
 sg13g2_buf_8 _1949_ (.A(_0067_),
    .X(_1386_));
 sg13g2_nor2b_2 _1950_ (.A(net106),
    .B_N(_1259_),
    .Y(_1387_));
 sg13g2_a21o_1 _1951_ (.A2(_1298_),
    .A1(net84),
    .B1(_1271_),
    .X(_1388_));
 sg13g2_a22oi_1 _1952_ (.Y(_1389_),
    .B1(_1388_),
    .B2(_1256_),
    .A2(_1387_),
    .A1(_1386_));
 sg13g2_nor2_1 _1953_ (.A(net106),
    .B(_1259_),
    .Y(_1390_));
 sg13g2_mux2_1 _1954_ (.A0(\rsa_e[2] ),
    .A1(\rsa_spi_wrapper_i.config_regs[58] ),
    .S(net84),
    .X(_1391_));
 sg13g2_a22oi_1 _1955_ (.Y(_1392_),
    .B1(_1391_),
    .B2(net86),
    .A2(_1390_),
    .A1(\rsa_p[2] ));
 sg13g2_nand2_1 _1956_ (.Y(_1393_),
    .A(net85),
    .B(_1392_));
 sg13g2_o21ai_1 _1957_ (.B1(_1393_),
    .Y(_1394_),
    .A1(net85),
    .A2(_1389_));
 sg13g2_a22oi_1 _1958_ (.Y(_1395_),
    .B1(_1300_),
    .B2(\rsa_spi_wrapper_i.config_regs[50] ),
    .A2(_1274_),
    .A1(\rsa_spi_wrapper_i.config_regs[10] ));
 sg13g2_a221oi_1 _1959_ (.B2(_1395_),
    .C1(_1306_),
    .B1(_1394_),
    .A1(_0066_),
    .Y(_1396_),
    .A2(net46));
 sg13g2_a21oi_1 _1960_ (.A1(net81),
    .A2(_1385_),
    .Y(_1397_),
    .B1(_1396_));
 sg13g2_mux2_1 _1961_ (.A0(_1397_),
    .A1(_0065_),
    .S(_1357_),
    .X(_1398_));
 sg13g2_nand2_1 _1962_ (.Y(_1399_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[2] ),
    .B(_1359_));
 sg13g2_o21ai_1 _1963_ (.B1(_1399_),
    .Y(_0225_),
    .A1(_1382_),
    .A2(_1398_));
 sg13g2_and2_1 _1964_ (.A(net106),
    .B(_1259_),
    .X(_1400_));
 sg13g2_a22oi_1 _1965_ (.Y(_1401_),
    .B1(_1400_),
    .B2(\rsa_spi_wrapper_i.config_regs[59] ),
    .A2(_1390_),
    .A1(\rsa_p[3] ));
 sg13g2_inv_1 _1966_ (.Y(_1402_),
    .A(_0070_));
 sg13g2_nor2_1 _1967_ (.A(_1288_),
    .B(_1271_),
    .Y(_1403_));
 sg13g2_a221oi_1 _1968_ (.B2(\rsa_const[3] ),
    .C1(net105),
    .B1(_1403_),
    .A1(_1402_),
    .Y(_1404_),
    .A2(_1387_));
 sg13g2_a21o_1 _1969_ (.A2(_1401_),
    .A1(net85),
    .B1(_1404_),
    .X(_1405_));
 sg13g2_nand2_1 _1970_ (.Y(_1406_),
    .A(\rsa_e[3] ),
    .B(_1346_));
 sg13g2_a22oi_1 _1971_ (.Y(_1407_),
    .B1(_1300_),
    .B2(\rsa_spi_wrapper_i.config_regs[51] ),
    .A2(_1274_),
    .A1(\rsa_spi_wrapper_i.config_regs[11] ));
 sg13g2_nand3_1 _1972_ (.B(_1406_),
    .C(_1407_),
    .A(_1405_),
    .Y(_1408_));
 sg13g2_nand2_1 _1973_ (.Y(_1409_),
    .A(_0069_),
    .B(net46));
 sg13g2_o21ai_1 _1974_ (.B1(_1409_),
    .Y(_1410_),
    .A1(net46),
    .A2(_1408_));
 sg13g2_nand2_1 _1975_ (.Y(_1411_),
    .A(_1277_),
    .B(_1387_));
 sg13g2_o21ai_1 _1976_ (.B1(_1411_),
    .Y(_1412_),
    .A1(net71),
    .A2(_1375_));
 sg13g2_and2_1 _1977_ (.A(\rsa_c[3] ),
    .B(_1333_),
    .X(_1413_));
 sg13g2_o21ai_1 _1978_ (.B1(net81),
    .Y(_1414_),
    .A1(_1412_),
    .A2(_1413_));
 sg13g2_o21ai_1 _1979_ (.B1(_1414_),
    .Y(_1415_),
    .A1(net81),
    .A2(_1410_));
 sg13g2_nand2_1 _1980_ (.Y(_1416_),
    .A(_0068_),
    .B(net56));
 sg13g2_o21ai_1 _1981_ (.B1(_1416_),
    .Y(_1417_),
    .A1(net56),
    .A2(_1415_));
 sg13g2_nand2_1 _1982_ (.Y(_1418_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[3] ),
    .B(_1359_));
 sg13g2_o21ai_1 _1983_ (.B1(_1418_),
    .Y(_0226_),
    .A1(_1382_),
    .A2(_1417_));
 sg13g2_buf_1 _1984_ (.A(_0073_),
    .X(_1419_));
 sg13g2_inv_2 _1985_ (.Y(_1420_),
    .A(_1419_));
 sg13g2_a22oi_1 _1986_ (.Y(_1421_),
    .B1(_1334_),
    .B2(_1420_),
    .A2(_1341_),
    .A1(\rsa_p[4] ));
 sg13g2_a221oi_1 _1987_ (.B2(\rsa_spi_wrapper_i.config_regs[60] ),
    .C1(_1289_),
    .B1(_1338_),
    .A1(\rsa_spi_wrapper_i.config_regs[12] ),
    .Y(_1422_),
    .A2(_1272_));
 sg13g2_a21oi_1 _1988_ (.A1(net71),
    .A2(_1421_),
    .Y(_1423_),
    .B1(_1422_));
 sg13g2_a22oi_1 _1989_ (.Y(_1424_),
    .B1(_1368_),
    .B2(\rsa_spi_wrapper_i.config_regs[52] ),
    .A2(_1367_),
    .A1(\rsa_const[4] ));
 sg13g2_nand2_1 _1990_ (.Y(_1425_),
    .A(\rsa_e[4] ),
    .B(_1346_));
 sg13g2_o21ai_1 _1991_ (.B1(_1425_),
    .Y(_1426_),
    .A1(_1295_),
    .A2(_1424_));
 sg13g2_nor3_1 _1992_ (.A(_1329_),
    .B(_1423_),
    .C(_1426_),
    .Y(_1427_));
 sg13g2_a21o_1 _1993_ (.A2(net46),
    .A1(_0072_),
    .B1(_1427_),
    .X(_1428_));
 sg13g2_inv_1 _1994_ (.Y(_1429_),
    .A(\rsa_c[4] ));
 sg13g2_o21ai_1 _1995_ (.B1(_1387_),
    .Y(_1430_),
    .A1(net82),
    .A2(_1429_));
 sg13g2_nand3_1 _1996_ (.B(_1306_),
    .C(_1430_),
    .A(_1258_),
    .Y(_1431_));
 sg13g2_o21ai_1 _1997_ (.B1(_1431_),
    .Y(_1432_),
    .A1(net81),
    .A2(_1428_));
 sg13g2_nand2_1 _1998_ (.Y(_1433_),
    .A(_0071_),
    .B(net56));
 sg13g2_o21ai_1 _1999_ (.B1(_1433_),
    .Y(_1434_),
    .A1(net56),
    .A2(_1432_));
 sg13g2_nand2_1 _2000_ (.Y(_1435_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[4] ),
    .B(_1359_));
 sg13g2_o21ai_1 _2001_ (.B1(_1435_),
    .Y(_0227_),
    .A1(_1382_),
    .A2(_1434_));
 sg13g2_a22oi_1 _2002_ (.Y(_1436_),
    .B1(_1400_),
    .B2(\rsa_spi_wrapper_i.config_regs[61] ),
    .A2(_1390_),
    .A1(\rsa_p[5] ));
 sg13g2_buf_8 _2003_ (.A(_0076_),
    .X(_1437_));
 sg13g2_inv_1 _2004_ (.Y(_1438_),
    .A(_1437_));
 sg13g2_a221oi_1 _2005_ (.B2(\rsa_const[5] ),
    .C1(net105),
    .B1(_1403_),
    .A1(_1438_),
    .Y(_1439_),
    .A2(_1387_));
 sg13g2_a21oi_1 _2006_ (.A1(net85),
    .A2(_1436_),
    .Y(_1440_),
    .B1(_1439_));
 sg13g2_nand2_1 _2007_ (.Y(_1441_),
    .A(\rsa_e[5] ),
    .B(_1346_));
 sg13g2_a22oi_1 _2008_ (.Y(_1442_),
    .B1(_1300_),
    .B2(\rsa_spi_wrapper_i.config_regs[53] ),
    .A2(_1274_),
    .A1(\rsa_spi_wrapper_i.config_regs[13] ));
 sg13g2_nand2_1 _2009_ (.Y(_1443_),
    .A(_1441_),
    .B(_1442_));
 sg13g2_nor3_1 _2010_ (.A(_1329_),
    .B(_1440_),
    .C(_1443_),
    .Y(_1444_));
 sg13g2_a21oi_1 _2011_ (.A1(_0075_),
    .A2(net46),
    .Y(_1445_),
    .B1(_1444_));
 sg13g2_a21oi_1 _2012_ (.A1(\rsa_c[5] ),
    .A2(_1333_),
    .Y(_1446_),
    .B1(_1334_));
 sg13g2_o21ai_1 _2013_ (.B1(_1303_),
    .Y(_1447_),
    .A1(net86),
    .A2(_1446_));
 sg13g2_mux2_1 _2014_ (.A0(_1445_),
    .A1(_1447_),
    .S(_1306_),
    .X(_1448_));
 sg13g2_nand2_1 _2015_ (.Y(_1449_),
    .A(_0074_),
    .B(net56));
 sg13g2_o21ai_1 _2016_ (.B1(_1449_),
    .Y(_1450_),
    .A1(_1361_),
    .A2(_1448_));
 sg13g2_nand2_1 _2017_ (.Y(_1451_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[5] ),
    .B(_1359_));
 sg13g2_o21ai_1 _2018_ (.B1(_1451_),
    .Y(_0228_),
    .A1(_1382_),
    .A2(_1450_));
 sg13g2_inv_2 _2019_ (.Y(_1452_),
    .A(_0079_));
 sg13g2_a22oi_1 _2020_ (.Y(_1453_),
    .B1(_1334_),
    .B2(_1452_),
    .A2(_1341_),
    .A1(\rsa_p[6] ));
 sg13g2_a221oi_1 _2021_ (.B2(\rsa_spi_wrapper_i.config_regs[62] ),
    .C1(net71),
    .B1(_1338_),
    .A1(\rsa_spi_wrapper_i.config_regs[14] ),
    .Y(_1454_),
    .A2(_1272_));
 sg13g2_a21oi_1 _2022_ (.A1(net71),
    .A2(_1453_),
    .Y(_1455_),
    .B1(_1454_));
 sg13g2_a22oi_1 _2023_ (.Y(_1456_),
    .B1(_1368_),
    .B2(\rsa_spi_wrapper_i.config_regs[54] ),
    .A2(_1367_),
    .A1(\rsa_const[6] ));
 sg13g2_nand2_1 _2024_ (.Y(_1457_),
    .A(\rsa_e[6] ),
    .B(_1346_));
 sg13g2_o21ai_1 _2025_ (.B1(_1457_),
    .Y(_1458_),
    .A1(_1295_),
    .A2(_1456_));
 sg13g2_nor3_1 _2026_ (.A(_1329_),
    .B(_1455_),
    .C(_1458_),
    .Y(_1459_));
 sg13g2_a21o_1 _2027_ (.A2(_1330_),
    .A1(_0078_),
    .B1(_1459_),
    .X(_1460_));
 sg13g2_nor2b_1 _2028_ (.A(net82),
    .B_N(\rsa_c[6] ),
    .Y(_1461_));
 sg13g2_o21ai_1 _2029_ (.B1(_1376_),
    .Y(_1462_),
    .A1(net86),
    .A2(_1461_));
 sg13g2_o21ai_1 _2030_ (.B1(_1462_),
    .Y(_1463_),
    .A1(_1307_),
    .A2(_1460_));
 sg13g2_nand2_1 _2031_ (.Y(_0327_),
    .A(_0077_),
    .B(net56));
 sg13g2_o21ai_1 _2032_ (.B1(_0327_),
    .Y(_0328_),
    .A1(_1361_),
    .A2(_1463_));
 sg13g2_nand2_1 _2033_ (.Y(_0329_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[6] ),
    .B(_1359_));
 sg13g2_o21ai_1 _2034_ (.B1(_0329_),
    .Y(_0229_),
    .A1(_1382_),
    .A2(_0328_));
 sg13g2_a22oi_1 _2035_ (.Y(_0330_),
    .B1(_1400_),
    .B2(\rsa_spi_wrapper_i.config_regs[63] ),
    .A2(_1390_),
    .A1(\rsa_p[7] ));
 sg13g2_buf_1 _2036_ (.A(_0082_),
    .X(_0331_));
 sg13g2_inv_1 _2037_ (.Y(_0332_),
    .A(_0331_));
 sg13g2_a221oi_1 _2038_ (.B2(\rsa_const[7] ),
    .C1(net105),
    .B1(_1403_),
    .A1(_0332_),
    .Y(_0333_),
    .A2(_1387_));
 sg13g2_a21o_1 _2039_ (.A2(_0330_),
    .A1(net105),
    .B1(_0333_),
    .X(_0334_));
 sg13g2_nand2_1 _2040_ (.Y(_0335_),
    .A(\rsa_e[7] ),
    .B(_1346_));
 sg13g2_a22oi_1 _2041_ (.Y(_0336_),
    .B1(_1300_),
    .B2(\rsa_spi_wrapper_i.config_regs[55] ),
    .A2(_1274_),
    .A1(\rsa_spi_wrapper_i.config_regs[15] ));
 sg13g2_nand3_1 _2042_ (.B(_0335_),
    .C(_0336_),
    .A(_0334_),
    .Y(_0337_));
 sg13g2_nand2_1 _2043_ (.Y(_0338_),
    .A(_0081_),
    .B(_1329_));
 sg13g2_o21ai_1 _2044_ (.B1(_0338_),
    .Y(_0339_),
    .A1(net46),
    .A2(_0337_));
 sg13g2_and2_1 _2045_ (.A(\rsa_c[7] ),
    .B(_1333_),
    .X(_0340_));
 sg13g2_o21ai_1 _2046_ (.B1(net81),
    .Y(_0341_),
    .A1(_1412_),
    .A2(_0340_));
 sg13g2_o21ai_1 _2047_ (.B1(_0341_),
    .Y(_0342_),
    .A1(net81),
    .A2(_0339_));
 sg13g2_nand2_1 _2048_ (.Y(_0343_),
    .A(_0080_),
    .B(_1357_));
 sg13g2_o21ai_1 _2049_ (.B1(_0343_),
    .Y(_0344_),
    .A1(net56),
    .A2(_0342_));
 sg13g2_nand2_1 _2050_ (.Y(_0345_),
    .A(\rsa_spi_wrapper_i.spi_miso ),
    .B(_1359_));
 sg13g2_o21ai_1 _2051_ (.B1(_0345_),
    .Y(_0230_),
    .A1(_1382_),
    .A2(_0344_));
 sg13g2_xnor2_1 _2052_ (.Y(_0346_),
    .A(_1167_),
    .B(_1318_));
 sg13g2_a21oi_1 _2053_ (.A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .A2(_1352_),
    .Y(_0231_),
    .B1(_0346_));
 sg13g2_nand2_1 _2054_ (.Y(_0347_),
    .A(_1167_),
    .B(_1318_));
 sg13g2_xnor2_1 _2055_ (.Y(_0232_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .B(_0347_));
 sg13g2_nand3_1 _2056_ (.B(_1167_),
    .C(_1318_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .Y(_0348_));
 sg13g2_xnor2_1 _2057_ (.Y(_0233_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .B(_0348_));
 sg13g2_nand3_1 _2058_ (.B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .C(_1319_),
    .A(_1167_),
    .Y(_0349_));
 sg13g2_nor2_1 _2059_ (.A(_1167_),
    .B(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .Y(_0350_));
 sg13g2_a21oi_1 _2060_ (.A1(net88),
    .A2(_0350_),
    .Y(_0351_),
    .B1(_1350_));
 sg13g2_and4_1 _2061_ (.A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .B(_1167_),
    .C(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ),
    .D(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ),
    .X(_0352_));
 sg13g2_o21ai_1 _2062_ (.B1(_1318_),
    .Y(_0353_),
    .A1(_1168_),
    .A2(_0352_));
 sg13g2_o21ai_1 _2063_ (.B1(_0353_),
    .Y(_0354_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ),
    .A2(_0351_));
 sg13g2_a21oi_1 _2064_ (.A1(_1350_),
    .A2(_0349_),
    .Y(_0234_),
    .B1(_0354_));
 sg13g2_buf_1 _2065_ (.A(\rsa_unit_i.rsa_control_fsm.load_exp ),
    .X(_0355_));
 sg13g2_nor4_1 _2066_ (.A(net109),
    .B(net110),
    .C(_1229_),
    .D(net96),
    .Y(_0356_));
 sg13g2_or4_1 _2067_ (.A(net110),
    .B(_1172_),
    .C(_1229_),
    .D(\rsa_unit_i.rsa_control_fsm.state[11] ),
    .X(_0357_));
 sg13g2_buf_1 _2068_ (.A(_0357_),
    .X(_0358_));
 sg13g2_or3_1 _2069_ (.A(net109),
    .B(\rsa_unit_i.rsa_control_fsm.state[8] ),
    .C(\rsa_unit_i.rsa_control_fsm.state[2] ),
    .X(_0359_));
 sg13g2_buf_1 _2070_ (.A(_0359_),
    .X(_0360_));
 sg13g2_nor2_1 _2071_ (.A(_0358_),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_buf_1 _2072_ (.A(_0361_),
    .X(_0362_));
 sg13g2_buf_1 _2073_ (.A(net55),
    .X(_0363_));
 sg13g2_nor3_2 _2074_ (.A(\rsa_unit_i.rsa_control_fsm.state[3] ),
    .B(net96),
    .C(\rsa_unit_i.rsa_control_fsm.state[6] ),
    .Y(_0364_));
 sg13g2_nand2_1 _2075_ (.Y(_0365_),
    .A(_0363_),
    .B(_0364_));
 sg13g2_nand2_1 _2076_ (.Y(_0366_),
    .A(net65),
    .B(_0365_));
 sg13g2_or2_1 _2077_ (.X(_0367_),
    .B(_0366_),
    .A(_0356_));
 sg13g2_buf_1 _2078_ (.A(_0367_),
    .X(_0368_));
 sg13g2_buf_1 _2079_ (.A(net29),
    .X(_0369_));
 sg13g2_nor2_1 _2080_ (.A(net109),
    .B(\rsa_unit_i.rsa_control_fsm.state[2] ),
    .Y(_0370_));
 sg13g2_buf_1 _2081_ (.A(_0370_),
    .X(_0371_));
 sg13g2_and2_1 _2082_ (.A(net108),
    .B(net70),
    .X(_0372_));
 sg13g2_buf_1 _2083_ (.A(_0372_),
    .X(_0373_));
 sg13g2_nor3_2 _2084_ (.A(net110),
    .B(_1172_),
    .C(_1229_),
    .Y(_0374_));
 sg13g2_nor2b_2 _2085_ (.A(\rsa_unit_i.rsa_control_fsm.state[10] ),
    .B_N(_0055_),
    .Y(_0375_));
 sg13g2_nand2_1 _2086_ (.Y(_0376_),
    .A(_0374_),
    .B(_0375_));
 sg13g2_buf_1 _2087_ (.A(_0376_),
    .X(_0377_));
 sg13g2_nor2_1 _2088_ (.A(net54),
    .B(net61),
    .Y(_0378_));
 sg13g2_buf_1 _2089_ (.A(_0378_),
    .X(_0379_));
 sg13g2_and2_1 _2090_ (.A(_0374_),
    .B(_0375_),
    .X(_0380_));
 sg13g2_buf_8 _2091_ (.A(_0380_),
    .X(_0381_));
 sg13g2_nand2b_1 _2092_ (.Y(_0382_),
    .B(_0381_),
    .A_N(\rsa_const[0] ));
 sg13g2_buf_1 _2093_ (.A(net54),
    .X(_0383_));
 sg13g2_a22oi_1 _2094_ (.Y(_0384_),
    .B1(_0382_),
    .B2(net44),
    .A2(net39),
    .A1(\rsa_unit_i.R_i[0] ));
 sg13g2_buf_1 _2095_ (.A(_0044_),
    .X(_0385_));
 sg13g2_nand2_2 _2096_ (.Y(_0386_),
    .A(_1232_),
    .B(_0371_));
 sg13g2_a21oi_1 _2097_ (.A1(\rsa_unit_i.rsa_control_fsm.exp[0] ),
    .A2(_0386_),
    .Y(_0387_),
    .B1(_0358_));
 sg13g2_nand2_1 _2098_ (.Y(_0388_),
    .A(_0364_),
    .B(_0387_));
 sg13g2_buf_1 _2099_ (.A(_0388_),
    .X(_0389_));
 sg13g2_mux2_1 _2100_ (.A0(_0384_),
    .A1(net95),
    .S(_0389_),
    .X(_0390_));
 sg13g2_a21o_1 _2101_ (.A2(_0365_),
    .A1(_0356_),
    .B1(_1186_),
    .X(_0391_));
 sg13g2_buf_1 _2102_ (.A(_0391_),
    .X(_0392_));
 sg13g2_nand2_1 _2103_ (.Y(_0393_),
    .A(\rsa_unit_i.R_i[0] ),
    .B(net33));
 sg13g2_o21ai_1 _2104_ (.B1(_0393_),
    .Y(_0254_),
    .A1(_0369_),
    .A2(_0390_));
 sg13g2_buf_1 _2105_ (.A(net38),
    .X(_0394_));
 sg13g2_nor2_1 _2106_ (.A(\rsa_const[1] ),
    .B(_0386_),
    .Y(_0395_));
 sg13g2_inv_1 _2107_ (.Y(_0396_),
    .A(_0027_));
 sg13g2_nor2_1 _2108_ (.A(_0396_),
    .B(net44),
    .Y(_0397_));
 sg13g2_nor3_1 _2109_ (.A(net61),
    .B(_0395_),
    .C(_0397_),
    .Y(_0398_));
 sg13g2_nand2_1 _2110_ (.Y(_0399_),
    .A(_0043_),
    .B(net36));
 sg13g2_o21ai_1 _2111_ (.B1(_0399_),
    .Y(_0400_),
    .A1(net36),
    .A2(_0398_));
 sg13g2_nand2_1 _2112_ (.Y(_0401_),
    .A(\rsa_unit_i.R_i[1] ),
    .B(net33));
 sg13g2_o21ai_1 _2113_ (.B1(_0401_),
    .Y(_0255_),
    .A1(net27),
    .A2(_0400_));
 sg13g2_nor2_1 _2114_ (.A(_0029_),
    .B(_0383_),
    .Y(_0402_));
 sg13g2_a21oi_1 _2115_ (.A1(\rsa_const[2] ),
    .A2(_0383_),
    .Y(_0403_),
    .B1(_0402_));
 sg13g2_nor2_1 _2116_ (.A(net61),
    .B(_0403_),
    .Y(_0404_));
 sg13g2_nand2_1 _2117_ (.Y(_0405_),
    .A(_0045_),
    .B(net38));
 sg13g2_o21ai_1 _2118_ (.B1(_0405_),
    .Y(_0406_),
    .A1(net36),
    .A2(_0404_));
 sg13g2_nand2_1 _2119_ (.Y(_0407_),
    .A(\rsa_unit_i.R_i[2] ),
    .B(net33));
 sg13g2_o21ai_1 _2120_ (.B1(_0407_),
    .Y(_0256_),
    .A1(net27),
    .A2(_0406_));
 sg13g2_nor2_1 _2121_ (.A(_0031_),
    .B(net54),
    .Y(_0408_));
 sg13g2_a21oi_1 _2122_ (.A1(\rsa_const[3] ),
    .A2(net44),
    .Y(_0409_),
    .B1(_0408_));
 sg13g2_nor2_1 _2123_ (.A(net61),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_nand2_1 _2124_ (.Y(_0411_),
    .A(_0046_),
    .B(net38));
 sg13g2_o21ai_1 _2125_ (.B1(_0411_),
    .Y(_0412_),
    .A1(net36),
    .A2(_0410_));
 sg13g2_nand2_1 _2126_ (.Y(_0413_),
    .A(\rsa_unit_i.R_i[3] ),
    .B(net33));
 sg13g2_o21ai_1 _2127_ (.B1(_0413_),
    .Y(_0257_),
    .A1(net27),
    .A2(_0412_));
 sg13g2_nor2_1 _2128_ (.A(_0033_),
    .B(net54),
    .Y(_0414_));
 sg13g2_a21oi_1 _2129_ (.A1(\rsa_const[4] ),
    .A2(net44),
    .Y(_0415_),
    .B1(_0414_));
 sg13g2_nor2_1 _2130_ (.A(net61),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_buf_1 _2131_ (.A(_0047_),
    .X(_0417_));
 sg13g2_nand2_1 _2132_ (.Y(_0418_),
    .A(_0417_),
    .B(net38));
 sg13g2_o21ai_1 _2133_ (.B1(_0418_),
    .Y(_0419_),
    .A1(net36),
    .A2(_0416_));
 sg13g2_nand2_1 _2134_ (.Y(_0420_),
    .A(\rsa_unit_i.R_i[4] ),
    .B(_0392_));
 sg13g2_o21ai_1 _2135_ (.B1(_0420_),
    .Y(_0258_),
    .A1(net27),
    .A2(_0419_));
 sg13g2_nor2_1 _2136_ (.A(_0035_),
    .B(net54),
    .Y(_0421_));
 sg13g2_a21oi_1 _2137_ (.A1(\rsa_const[5] ),
    .A2(net44),
    .Y(_0422_),
    .B1(_0421_));
 sg13g2_nor2_1 _2138_ (.A(net61),
    .B(_0422_),
    .Y(_0423_));
 sg13g2_nand2_1 _2139_ (.Y(_0424_),
    .A(_0048_),
    .B(net38));
 sg13g2_o21ai_1 _2140_ (.B1(_0424_),
    .Y(_0425_),
    .A1(_0394_),
    .A2(_0423_));
 sg13g2_nand2_1 _2141_ (.Y(_0426_),
    .A(\rsa_unit_i.R_i[5] ),
    .B(_0392_));
 sg13g2_o21ai_1 _2142_ (.B1(_0426_),
    .Y(_0259_),
    .A1(net27),
    .A2(_0425_));
 sg13g2_nor2_1 _2143_ (.A(_0037_),
    .B(_0373_),
    .Y(_0427_));
 sg13g2_a21oi_1 _2144_ (.A1(\rsa_const[6] ),
    .A2(net44),
    .Y(_0428_),
    .B1(_0427_));
 sg13g2_nor2_1 _2145_ (.A(_0377_),
    .B(_0428_),
    .Y(_0429_));
 sg13g2_nand2_1 _2146_ (.Y(_0430_),
    .A(_0049_),
    .B(net38));
 sg13g2_o21ai_1 _2147_ (.B1(_0430_),
    .Y(_0431_),
    .A1(_0394_),
    .A2(_0429_));
 sg13g2_nand2_1 _2148_ (.Y(_0432_),
    .A(\rsa_unit_i.R_i[6] ),
    .B(net33));
 sg13g2_o21ai_1 _2149_ (.B1(_0432_),
    .Y(_0260_),
    .A1(net27),
    .A2(_0431_));
 sg13g2_nor2_1 _2150_ (.A(_0039_),
    .B(_0373_),
    .Y(_0433_));
 sg13g2_a21oi_1 _2151_ (.A1(\rsa_const[7] ),
    .A2(net44),
    .Y(_0434_),
    .B1(_0433_));
 sg13g2_nor2_1 _2152_ (.A(_0377_),
    .B(_0434_),
    .Y(_0435_));
 sg13g2_nand2_1 _2153_ (.Y(_0436_),
    .A(_0050_),
    .B(net38));
 sg13g2_o21ai_1 _2154_ (.B1(_0436_),
    .Y(_0437_),
    .A1(net36),
    .A2(_0435_));
 sg13g2_nand2_1 _2155_ (.Y(_0438_),
    .A(\rsa_unit_i.R_i[7] ),
    .B(net33));
 sg13g2_o21ai_1 _2156_ (.B1(_0438_),
    .Y(_0261_),
    .A1(net27),
    .A2(_0437_));
 sg13g2_nor3_1 _2157_ (.A(_0041_),
    .B(net44),
    .C(net61),
    .Y(_0439_));
 sg13g2_nand2_1 _2158_ (.Y(_0440_),
    .A(_0051_),
    .B(net38));
 sg13g2_o21ai_1 _2159_ (.B1(_0440_),
    .Y(_0441_),
    .A1(net36),
    .A2(_0439_));
 sg13g2_nand2_1 _2160_ (.Y(_0442_),
    .A(\rsa_unit_i.R_i[8] ),
    .B(net33));
 sg13g2_o21ai_1 _2161_ (.B1(_0442_),
    .Y(_0262_),
    .A1(net27),
    .A2(_0441_));
 sg13g2_inv_1 _2162_ (.Y(_0443_),
    .A(_0042_));
 sg13g2_nand2_1 _2163_ (.Y(_0444_),
    .A(_0443_),
    .B(net39));
 sg13g2_nor3_1 _2164_ (.A(net29),
    .B(net36),
    .C(_0444_),
    .Y(_0445_));
 sg13g2_a21o_1 _2165_ (.A2(net33),
    .A1(\rsa_unit_i.R_i[9] ),
    .B1(_0445_),
    .X(_0263_));
 sg13g2_nor4_2 _2166_ (.A(net110),
    .B(_1172_),
    .C(_1229_),
    .Y(_0446_),
    .D(\rsa_unit_i.rsa_control_fsm.state[11] ));
 sg13g2_nor3_1 _2167_ (.A(net109),
    .B(\rsa_unit_i.rsa_control_fsm.state[8] ),
    .C(\rsa_unit_i.rsa_control_fsm.state[2] ),
    .Y(_0447_));
 sg13g2_buf_8 _2168_ (.A(_0447_),
    .X(_0448_));
 sg13g2_buf_1 _2169_ (.A(_0084_),
    .X(_0449_));
 sg13g2_inv_1 _2170_ (.Y(_0450_),
    .A(_0449_));
 sg13g2_a21oi_2 _2171_ (.B1(_0450_),
    .Y(_0451_),
    .A2(net69),
    .A1(_0446_));
 sg13g2_a21o_1 _2172_ (.A2(net45),
    .A1(_0085_),
    .B1(_0451_),
    .X(_0452_));
 sg13g2_nand2_2 _2173_ (.Y(_0453_),
    .A(_0448_),
    .B(_0364_));
 sg13g2_buf_1 _2174_ (.A(_0453_),
    .X(_0454_));
 sg13g2_mux2_1 _2175_ (.A0(_0452_),
    .A1(_0109_),
    .S(net53),
    .X(_0455_));
 sg13g2_buf_1 _2176_ (.A(_0391_),
    .X(_0456_));
 sg13g2_nand2_1 _2177_ (.Y(_0457_),
    .A(\rsa_unit_i.P_i[0] ),
    .B(net32));
 sg13g2_o21ai_1 _2178_ (.B1(_0457_),
    .Y(_0283_),
    .A1(_0369_),
    .A2(_0455_));
 sg13g2_mux2_1 _2179_ (.A0(_0087_),
    .A1(_0088_),
    .S(net45),
    .X(_0458_));
 sg13g2_mux2_1 _2180_ (.A0(_0458_),
    .A1(_0107_),
    .S(_0454_),
    .X(_0459_));
 sg13g2_buf_1 _2181_ (.A(\rsa_unit_i.P_i[1] ),
    .X(_0460_));
 sg13g2_nand2_1 _2182_ (.Y(_0461_),
    .A(net94),
    .B(net32));
 sg13g2_o21ai_1 _2183_ (.B1(_0461_),
    .Y(_0284_),
    .A1(net29),
    .A2(_0459_));
 sg13g2_inv_1 _2184_ (.Y(_0462_),
    .A(_0090_));
 sg13g2_a21oi_1 _2185_ (.A1(_0446_),
    .A2(net69),
    .Y(_0463_),
    .B1(_0462_));
 sg13g2_a21oi_1 _2186_ (.A1(_0091_),
    .A2(net45),
    .Y(_0464_),
    .B1(_0463_));
 sg13g2_nand2_1 _2187_ (.Y(_0465_),
    .A(_0110_),
    .B(_0454_));
 sg13g2_o21ai_1 _2188_ (.B1(_0465_),
    .Y(_0466_),
    .A1(net53),
    .A2(_0464_));
 sg13g2_nand2_1 _2189_ (.Y(_0467_),
    .A(\rsa_unit_i.P_i[2] ),
    .B(_0456_));
 sg13g2_o21ai_1 _2190_ (.B1(_0467_),
    .Y(_0285_),
    .A1(net29),
    .A2(_0466_));
 sg13g2_mux2_1 _2191_ (.A0(_0093_),
    .A1(_0094_),
    .S(net45),
    .X(_0468_));
 sg13g2_mux2_1 _2192_ (.A0(_0468_),
    .A1(_0112_),
    .S(net53),
    .X(_0469_));
 sg13g2_nand2_1 _2193_ (.Y(_0470_),
    .A(\rsa_unit_i.P_i[3] ),
    .B(net32));
 sg13g2_o21ai_1 _2194_ (.B1(_0470_),
    .Y(_0286_),
    .A1(net29),
    .A2(_0469_));
 sg13g2_inv_1 _2195_ (.Y(_0471_),
    .A(_0114_));
 sg13g2_nand2_2 _2196_ (.Y(_0472_),
    .A(_0446_),
    .B(net69));
 sg13g2_buf_1 _2197_ (.A(_0472_),
    .X(_0473_));
 sg13g2_and2_1 _2198_ (.A(_0096_),
    .B(net52),
    .X(_0474_));
 sg13g2_a21o_1 _2199_ (.A2(net45),
    .A1(_0097_),
    .B1(_0474_),
    .X(_0475_));
 sg13g2_nor2_1 _2200_ (.A(net53),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_a21oi_1 _2201_ (.A1(_0471_),
    .A2(net53),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_nand2_1 _2202_ (.Y(_0478_),
    .A(\rsa_unit_i.P_i[4] ),
    .B(net32));
 sg13g2_o21ai_1 _2203_ (.B1(_0478_),
    .Y(_0287_),
    .A1(net29),
    .A2(_0477_));
 sg13g2_inv_2 _2204_ (.Y(_0479_),
    .A(_0116_));
 sg13g2_inv_1 _2205_ (.Y(_0480_),
    .A(_0100_));
 sg13g2_buf_1 _2206_ (.A(_0473_),
    .X(_0481_));
 sg13g2_o21ai_1 _2207_ (.B1(_0099_),
    .Y(_0482_),
    .A1(_0358_),
    .A2(_0360_));
 sg13g2_o21ai_1 _2208_ (.B1(_0482_),
    .Y(_0483_),
    .A1(_0480_),
    .A2(net43));
 sg13g2_nor2_1 _2209_ (.A(net53),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_a21oi_1 _2210_ (.A1(_0479_),
    .A2(net53),
    .Y(_0485_),
    .B1(_0484_));
 sg13g2_nand2_1 _2211_ (.Y(_0486_),
    .A(\rsa_unit_i.P_i[5] ),
    .B(_0456_));
 sg13g2_o21ai_1 _2212_ (.B1(_0486_),
    .Y(_0288_),
    .A1(net29),
    .A2(_0485_));
 sg13g2_and2_1 _2213_ (.A(_0102_),
    .B(net52),
    .X(_0487_));
 sg13g2_a21o_1 _2214_ (.A2(net45),
    .A1(_0103_),
    .B1(_0487_),
    .X(_0488_));
 sg13g2_mux2_1 _2215_ (.A0(_0488_),
    .A1(_0020_),
    .S(_0453_),
    .X(_0489_));
 sg13g2_nand2_1 _2216_ (.Y(_0490_),
    .A(\rsa_unit_i.P_i[6] ),
    .B(net32));
 sg13g2_o21ai_1 _2217_ (.B1(_0490_),
    .Y(_0289_),
    .A1(net29),
    .A2(_0489_));
 sg13g2_and2_1 _2218_ (.A(_0105_),
    .B(net52),
    .X(_0491_));
 sg13g2_a21o_1 _2219_ (.A2(net45),
    .A1(_0106_),
    .B1(_0491_),
    .X(_0492_));
 sg13g2_mux2_1 _2220_ (.A0(_0492_),
    .A1(_0022_),
    .S(_0453_),
    .X(_0493_));
 sg13g2_nand2_1 _2221_ (.Y(_0494_),
    .A(\rsa_unit_i.P_i[7] ),
    .B(net32));
 sg13g2_o21ai_1 _2222_ (.B1(_0494_),
    .Y(_0290_),
    .A1(_0368_),
    .A2(_0493_));
 sg13g2_nand2_1 _2223_ (.Y(_0495_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[8].fa.HA1.a ),
    .B(net53));
 sg13g2_nor3_1 _2224_ (.A(_0363_),
    .B(_0367_),
    .C(_0453_),
    .Y(_0496_));
 sg13g2_o21ai_1 _2225_ (.B1(\rsa_unit_i.P_i[8] ),
    .Y(_0497_),
    .A1(net32),
    .A2(_0496_));
 sg13g2_o21ai_1 _2226_ (.B1(_0497_),
    .Y(_0291_),
    .A1(_0368_),
    .A2(_0495_));
 sg13g2_o21ai_1 _2227_ (.B1(\rsa_unit_i.P_i[9] ),
    .Y(_0498_),
    .A1(net32),
    .A2(_0496_));
 sg13g2_inv_1 _2228_ (.Y(_0292_),
    .A(_0498_));
 sg13g2_mux2_1 _2229_ (.A0(\rsa_unit_i.R_i[0] ),
    .A1(\rsa_c[0] ),
    .S(net48),
    .X(_0293_));
 sg13g2_mux2_1 _2230_ (.A0(\rsa_unit_i.R_i[1] ),
    .A1(\rsa_c[1] ),
    .S(net48),
    .X(_0294_));
 sg13g2_mux2_1 _2231_ (.A0(\rsa_unit_i.R_i[2] ),
    .A1(\rsa_c[2] ),
    .S(net48),
    .X(_0295_));
 sg13g2_mux2_1 _2232_ (.A0(\rsa_unit_i.R_i[3] ),
    .A1(\rsa_c[3] ),
    .S(net48),
    .X(_0296_));
 sg13g2_mux2_1 _2233_ (.A0(\rsa_unit_i.R_i[4] ),
    .A1(\rsa_c[4] ),
    .S(net48),
    .X(_0297_));
 sg13g2_mux2_1 _2234_ (.A0(\rsa_unit_i.R_i[5] ),
    .A1(\rsa_c[5] ),
    .S(net48),
    .X(_0298_));
 sg13g2_mux2_1 _2235_ (.A0(\rsa_unit_i.R_i[6] ),
    .A1(\rsa_c[6] ),
    .S(net48),
    .X(_0299_));
 sg13g2_mux2_1 _2236_ (.A0(\rsa_unit_i.R_i[7] ),
    .A1(\rsa_c[7] ),
    .S(net48),
    .X(_0300_));
 sg13g2_nor2_1 _2237_ (.A(net109),
    .B(net110),
    .Y(_0499_));
 sg13g2_or2_1 _2238_ (.X(_0500_),
    .B(_0499_),
    .A(_1186_));
 sg13g2_buf_1 _2239_ (.A(_0500_),
    .X(_0501_));
 sg13g2_nor3_1 _2240_ (.A(_1207_),
    .B(_1214_),
    .C(_0501_),
    .Y(_0502_));
 sg13g2_a21o_1 _2241_ (.A2(_0501_),
    .A1(_1214_),
    .B1(_0502_),
    .X(_0301_));
 sg13g2_inv_1 _2242_ (.Y(_0503_),
    .A(_0058_));
 sg13g2_nor2_1 _2243_ (.A(_1187_),
    .B(_0499_),
    .Y(_0504_));
 sg13g2_o21ai_1 _2244_ (.B1(_0504_),
    .Y(_0505_),
    .A1(_1214_),
    .A2(_0503_));
 sg13g2_nor3_1 _2245_ (.A(_0503_),
    .B(_1215_),
    .C(_0501_),
    .Y(_0506_));
 sg13g2_a21o_1 _2246_ (.A2(_0505_),
    .A1(\rsa_unit_i.rsa_control_fsm.counter_rounds[1] ),
    .B1(_0506_),
    .X(_0302_));
 sg13g2_nand4_1 _2247_ (.B(\rsa_unit_i.rsa_control_fsm.counter_rounds[1] ),
    .C(_0058_),
    .A(_1214_),
    .Y(_0507_),
    .D(_0504_));
 sg13g2_a21oi_1 _2248_ (.A1(_1214_),
    .A2(\rsa_unit_i.rsa_control_fsm.counter_rounds[1] ),
    .Y(_0508_),
    .B1(_0503_));
 sg13g2_o21ai_1 _2249_ (.B1(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ),
    .Y(_0509_),
    .A1(_0501_),
    .A2(_0508_));
 sg13g2_o21ai_1 _2250_ (.B1(_0509_),
    .Y(_0303_),
    .A1(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ),
    .A2(_0507_));
 sg13g2_nand3_1 _2251_ (.B(\rsa_unit_i.rsa_control_fsm.counter_rounds[1] ),
    .C(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ),
    .A(_1214_),
    .Y(_0510_));
 sg13g2_nor3_1 _2252_ (.A(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ),
    .B(_0501_),
    .C(_0510_),
    .Y(_0511_));
 sg13g2_a21o_1 _2253_ (.A2(_0510_),
    .A1(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ),
    .B1(_0511_),
    .X(_0512_));
 sg13g2_a22oi_1 _2254_ (.Y(_0513_),
    .B1(_0512_),
    .B2(_0058_),
    .A2(_0501_),
    .A1(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ));
 sg13g2_inv_1 _2255_ (.Y(_0304_),
    .A(_0513_));
 sg13g2_nand2_1 _2256_ (.Y(_0514_),
    .A(_0054_),
    .B(_0499_));
 sg13g2_nor4_1 _2257_ (.A(_1172_),
    .B(\rsa_unit_i.rsa_control_fsm.state[3] ),
    .C(\rsa_unit_i.rsa_control_fsm.state[8] ),
    .D(_0514_),
    .Y(_0515_));
 sg13g2_or2_1 _2258_ (.X(_0516_),
    .B(_0515_),
    .A(_1186_));
 sg13g2_buf_1 _2259_ (.A(_0516_),
    .X(_0517_));
 sg13g2_or2_1 _2260_ (.X(_0518_),
    .B(_0517_),
    .A(_0514_));
 sg13g2_nand2_1 _2261_ (.Y(_0519_),
    .A(_1176_),
    .B(_0517_));
 sg13g2_o21ai_1 _2262_ (.B1(_0519_),
    .Y(_0305_),
    .A1(_1176_),
    .A2(_0518_));
 sg13g2_nor2_1 _2263_ (.A(_1176_),
    .B(_0514_),
    .Y(_0520_));
 sg13g2_o21ai_1 _2264_ (.B1(\rsa_unit_i.rsa_control_fsm.counter_steps[1] ),
    .Y(_0521_),
    .A1(_0517_),
    .A2(_0520_));
 sg13g2_o21ai_1 _2265_ (.B1(_0521_),
    .Y(_0306_),
    .A1(_1177_),
    .A2(_0518_));
 sg13g2_nand3b_1 _2266_ (.B(\rsa_unit_i.rsa_control_fsm.counter_steps[1] ),
    .C(_1176_),
    .Y(_0522_),
    .A_N(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ));
 sg13g2_a21oi_1 _2267_ (.A1(_1176_),
    .A2(\rsa_unit_i.rsa_control_fsm.counter_steps[1] ),
    .Y(_0523_),
    .B1(_0514_));
 sg13g2_o21ai_1 _2268_ (.B1(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ),
    .Y(_0524_),
    .A1(_0517_),
    .A2(_0523_));
 sg13g2_o21ai_1 _2269_ (.B1(_0524_),
    .Y(_0307_),
    .A1(_0518_),
    .A2(_0522_));
 sg13g2_nand3_1 _2270_ (.B(\rsa_unit_i.rsa_control_fsm.counter_steps[1] ),
    .C(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ),
    .A(_1176_),
    .Y(_0525_));
 sg13g2_nor3_1 _2271_ (.A(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ),
    .B(_0517_),
    .C(_0525_),
    .Y(_0526_));
 sg13g2_a21oi_1 _2272_ (.A1(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ),
    .A2(_0525_),
    .Y(_0527_),
    .B1(_0526_));
 sg13g2_nand2_1 _2273_ (.Y(_0528_),
    .A(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ),
    .B(_0517_));
 sg13g2_o21ai_1 _2274_ (.B1(_0528_),
    .Y(_0308_),
    .A1(_0514_),
    .A2(_0527_));
 sg13g2_nor2_1 _2275_ (.A(net109),
    .B(net96),
    .Y(_0529_));
 sg13g2_a21oi_2 _2276_ (.B1(net64),
    .Y(_0530_),
    .A2(_0529_),
    .A1(net43));
 sg13g2_buf_1 _2277_ (.A(_0530_),
    .X(_0531_));
 sg13g2_buf_1 _2278_ (.A(net96),
    .X(_0532_));
 sg13g2_nor2b_1 _2279_ (.A(net80),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[1] ),
    .Y(_0533_));
 sg13g2_a22oi_1 _2280_ (.Y(_0534_),
    .B1(net43),
    .B2(_0533_),
    .A2(\rsa_e[0] ),
    .A1(net80));
 sg13g2_nor2_1 _2281_ (.A(\rsa_unit_i.rsa_control_fsm.exp[0] ),
    .B(net35),
    .Y(_0535_));
 sg13g2_a21oi_1 _2282_ (.A1(net35),
    .A2(_0534_),
    .Y(_0309_),
    .B1(_0535_));
 sg13g2_nor2b_1 _2283_ (.A(_0532_),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[2] ),
    .Y(_0536_));
 sg13g2_a22oi_1 _2284_ (.Y(_0537_),
    .B1(net43),
    .B2(_0536_),
    .A2(\rsa_e[1] ),
    .A1(net80));
 sg13g2_nor2_1 _2285_ (.A(\rsa_unit_i.rsa_control_fsm.exp[1] ),
    .B(net35),
    .Y(_0538_));
 sg13g2_a21oi_1 _2286_ (.A1(net35),
    .A2(_0537_),
    .Y(_0310_),
    .B1(_0538_));
 sg13g2_nor2b_1 _2287_ (.A(net96),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[3] ),
    .Y(_0539_));
 sg13g2_a22oi_1 _2288_ (.Y(_0540_),
    .B1(net43),
    .B2(_0539_),
    .A2(\rsa_e[2] ),
    .A1(net80));
 sg13g2_nor2_1 _2289_ (.A(\rsa_unit_i.rsa_control_fsm.exp[2] ),
    .B(_0530_),
    .Y(_0541_));
 sg13g2_a21oi_1 _2290_ (.A1(net35),
    .A2(_0540_),
    .Y(_0311_),
    .B1(_0541_));
 sg13g2_nor2b_1 _2291_ (.A(net96),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[4] ),
    .Y(_0542_));
 sg13g2_a22oi_1 _2292_ (.Y(_0543_),
    .B1(net43),
    .B2(_0542_),
    .A2(\rsa_e[3] ),
    .A1(_0532_));
 sg13g2_nor2_1 _2293_ (.A(\rsa_unit_i.rsa_control_fsm.exp[3] ),
    .B(_0530_),
    .Y(_0544_));
 sg13g2_a21oi_1 _2294_ (.A1(net35),
    .A2(_0543_),
    .Y(_0312_),
    .B1(_0544_));
 sg13g2_nor2b_1 _2295_ (.A(net96),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[5] ),
    .Y(_0545_));
 sg13g2_a22oi_1 _2296_ (.Y(_0546_),
    .B1(net43),
    .B2(_0545_),
    .A2(\rsa_e[4] ),
    .A1(net80));
 sg13g2_nor2_1 _2297_ (.A(\rsa_unit_i.rsa_control_fsm.exp[4] ),
    .B(_0530_),
    .Y(_0547_));
 sg13g2_a21oi_1 _2298_ (.A1(_0531_),
    .A2(_0546_),
    .Y(_0313_),
    .B1(_0547_));
 sg13g2_nor2b_1 _2299_ (.A(net96),
    .B_N(\rsa_unit_i.rsa_control_fsm.exp[6] ),
    .Y(_0548_));
 sg13g2_a22oi_1 _2300_ (.Y(_0549_),
    .B1(_0481_),
    .B2(_0548_),
    .A2(\rsa_e[5] ),
    .A1(net80));
 sg13g2_nor2_1 _2301_ (.A(\rsa_unit_i.rsa_control_fsm.exp[5] ),
    .B(_0530_),
    .Y(_0550_));
 sg13g2_a21oi_1 _2302_ (.A1(_0531_),
    .A2(_0549_),
    .Y(_0314_),
    .B1(_0550_));
 sg13g2_inv_1 _2303_ (.Y(_0551_),
    .A(\rsa_unit_i.rsa_control_fsm.exp[7] ));
 sg13g2_nor2_1 _2304_ (.A(_0355_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_a22oi_1 _2305_ (.Y(_0553_),
    .B1(_0481_),
    .B2(_0552_),
    .A2(\rsa_e[6] ),
    .A1(net80));
 sg13g2_nor2_1 _2306_ (.A(\rsa_unit_i.rsa_control_fsm.exp[6] ),
    .B(_0530_),
    .Y(_0554_));
 sg13g2_a21oi_1 _2307_ (.A1(net35),
    .A2(_0553_),
    .Y(_0315_),
    .B1(_0554_));
 sg13g2_nand3_1 _2308_ (.B(\rsa_e[7] ),
    .C(net65),
    .A(net80),
    .Y(_0555_));
 sg13g2_o21ai_1 _2309_ (.B1(_0555_),
    .Y(_0316_),
    .A1(_0551_),
    .A2(net35));
 sg13g2_mux2_1 _2310_ (.A0(\synchronizer_spi_clk_inst.data_sync[1] ),
    .A1(net7),
    .S(net72),
    .X(_0317_));
 sg13g2_mux2_1 _2311_ (.A0(\rsa_spi_wrapper_i.spi_clk ),
    .A1(\synchronizer_spi_clk_inst.data_sync[1] ),
    .S(net72),
    .X(_0318_));
 sg13g2_mux2_1 _2312_ (.A0(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .A1(net6),
    .S(net72),
    .X(_0319_));
 sg13g2_mux2_1 _2313_ (.A0(_1165_),
    .A1(\synchronizer_spi_cs_n_inst.data_sync[1] ),
    .S(net72),
    .X(_0320_));
 sg13g2_mux2_1 _2314_ (.A0(\synchronizer_spi_mode_cpha.data_sync[1] ),
    .A1(net5),
    .S(net87),
    .X(_0321_));
 sg13g2_mux2_1 _2315_ (.A0(cpha_sync),
    .A1(\synchronizer_spi_mode_cpha.data_sync[1] ),
    .S(net87),
    .X(_0322_));
 sg13g2_mux2_1 _2316_ (.A0(\synchronizer_spi_mode_cpol.data_sync[1] ),
    .A1(net4),
    .S(_1222_),
    .X(_0323_));
 sg13g2_mux2_1 _2317_ (.A0(cpol_sync),
    .A1(\synchronizer_spi_mode_cpol.data_sync[1] ),
    .S(_1222_),
    .X(_0324_));
 sg13g2_mux2_1 _2318_ (.A0(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .A1(net8),
    .S(net87),
    .X(_0325_));
 sg13g2_mux2_1 _2319_ (.A0(\rsa_spi_wrapper_i.spi_mosi ),
    .A1(\synchronizer_spi_mosi_inst.data_sync[1] ),
    .S(net87),
    .X(_0326_));
 sg13g2_nand2_1 _2320_ (.Y(_0556_),
    .A(_1182_),
    .B(_1175_));
 sg13g2_o21ai_1 _2321_ (.B1(_0556_),
    .Y(_0557_),
    .A1(_0118_),
    .A2(_1184_));
 sg13g2_inv_1 _2322_ (.Y(_0121_),
    .A(_0557_));
 sg13g2_buf_1 _2323_ (.A(_0366_),
    .X(_0558_));
 sg13g2_buf_1 _2324_ (.A(net31),
    .X(_0559_));
 sg13g2_nor2_1 _2325_ (.A(\rsa_unit_i.rsa_control_fsm.state[2] ),
    .B(\rsa_unit_i.rsa_control_fsm.state[6] ),
    .Y(_0560_));
 sg13g2_nand2_1 _2326_ (.Y(_0561_),
    .A(_0055_),
    .B(_0560_));
 sg13g2_buf_1 _2327_ (.A(_0561_),
    .X(_0562_));
 sg13g2_mux2_1 _2328_ (.A0(_0025_),
    .A1(_0384_),
    .S(net68),
    .X(_0563_));
 sg13g2_buf_1 _2329_ (.A(\rsa_unit_i.mmm_multiply.A_bit ),
    .X(_0564_));
 sg13g2_buf_1 _2330_ (.A(net93),
    .X(_0565_));
 sg13g2_buf_1 _2331_ (.A(net64),
    .X(_0566_));
 sg13g2_nand2_1 _2332_ (.Y(_0567_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_o21ai_1 _2333_ (.B1(_0567_),
    .Y(_0235_),
    .A1(_0559_),
    .A2(_0563_));
 sg13g2_buf_1 _2334_ (.A(net68),
    .X(_0568_));
 sg13g2_buf_1 _2335_ (.A(_0561_),
    .X(_0569_));
 sg13g2_nor2_1 _2336_ (.A(_0026_),
    .B(net67),
    .Y(_0570_));
 sg13g2_a21oi_1 _2337_ (.A1(_0398_),
    .A2(net60),
    .Y(_0571_),
    .B1(_0570_));
 sg13g2_nand2_1 _2338_ (.Y(_0572_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[1] ),
    .B(net51));
 sg13g2_o21ai_1 _2339_ (.B1(_0572_),
    .Y(_0236_),
    .A1(net28),
    .A2(_0571_));
 sg13g2_nor2_1 _2340_ (.A(_0028_),
    .B(net67),
    .Y(_0573_));
 sg13g2_a21oi_1 _2341_ (.A1(_0404_),
    .A2(net60),
    .Y(_0574_),
    .B1(_0573_));
 sg13g2_nand2_1 _2342_ (.Y(_0575_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[2] ),
    .B(net51));
 sg13g2_o21ai_1 _2343_ (.B1(_0575_),
    .Y(_0237_),
    .A1(_0559_),
    .A2(_0574_));
 sg13g2_nor2_1 _2344_ (.A(_0030_),
    .B(net67),
    .Y(_0576_));
 sg13g2_a21oi_1 _2345_ (.A1(_0410_),
    .A2(net60),
    .Y(_0577_),
    .B1(_0576_));
 sg13g2_nand2_1 _2346_ (.Y(_0578_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[3] ),
    .B(net51));
 sg13g2_o21ai_1 _2347_ (.B1(_0578_),
    .Y(_0238_),
    .A1(net28),
    .A2(_0577_));
 sg13g2_nor2_1 _2348_ (.A(_0032_),
    .B(net67),
    .Y(_0579_));
 sg13g2_a21oi_1 _2349_ (.A1(_0416_),
    .A2(net60),
    .Y(_0580_),
    .B1(_0579_));
 sg13g2_nand2_1 _2350_ (.Y(_0581_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[4] ),
    .B(net51));
 sg13g2_o21ai_1 _2351_ (.B1(_0581_),
    .Y(_0239_),
    .A1(net28),
    .A2(_0580_));
 sg13g2_nor2_1 _2352_ (.A(_0034_),
    .B(net67),
    .Y(_0582_));
 sg13g2_a21oi_1 _2353_ (.A1(_0423_),
    .A2(net60),
    .Y(_0583_),
    .B1(_0582_));
 sg13g2_nand2_1 _2354_ (.Y(_0584_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[5] ),
    .B(net51));
 sg13g2_o21ai_1 _2355_ (.B1(_0584_),
    .Y(_0240_),
    .A1(net28),
    .A2(_0583_));
 sg13g2_nor2_1 _2356_ (.A(_0036_),
    .B(net67),
    .Y(_0585_));
 sg13g2_a21oi_1 _2357_ (.A1(_0429_),
    .A2(net60),
    .Y(_0586_),
    .B1(_0585_));
 sg13g2_nand2_1 _2358_ (.Y(_0587_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[6] ),
    .B(_0566_));
 sg13g2_o21ai_1 _2359_ (.B1(_0587_),
    .Y(_0241_),
    .A1(net28),
    .A2(_0586_));
 sg13g2_nor2_1 _2360_ (.A(_0038_),
    .B(net67),
    .Y(_0588_));
 sg13g2_a21oi_1 _2361_ (.A1(_0435_),
    .A2(net60),
    .Y(_0589_),
    .B1(_0588_));
 sg13g2_nand2_1 _2362_ (.Y(_0590_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[7] ),
    .B(net51));
 sg13g2_o21ai_1 _2363_ (.B1(_0590_),
    .Y(_0242_),
    .A1(net28),
    .A2(_0589_));
 sg13g2_nor2_1 _2364_ (.A(_0040_),
    .B(net67),
    .Y(_0591_));
 sg13g2_a21oi_1 _2365_ (.A1(_0439_),
    .A2(net60),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_nand2_1 _2366_ (.Y(_0593_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[8] ),
    .B(net51));
 sg13g2_o21ai_1 _2367_ (.B1(_0593_),
    .Y(_0243_),
    .A1(net28),
    .A2(_0592_));
 sg13g2_nand3_1 _2368_ (.B(net39),
    .C(_0568_),
    .A(_0443_),
    .Y(_0594_));
 sg13g2_nand2_1 _2369_ (.Y(_0595_),
    .A(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[9] ),
    .B(net51));
 sg13g2_o21ai_1 _2370_ (.B1(_0595_),
    .Y(_0244_),
    .A1(net28),
    .A2(_0594_));
 sg13g2_or2_1 _2371_ (.X(_0596_),
    .B(_0561_),
    .A(_0366_));
 sg13g2_buf_1 _2372_ (.A(_0596_),
    .X(_0597_));
 sg13g2_buf_1 _2373_ (.A(_0597_),
    .X(_0598_));
 sg13g2_buf_1 _2374_ (.A(net26),
    .X(_0599_));
 sg13g2_nor2_1 _2375_ (.A(_1293_),
    .B(net95),
    .Y(_0600_));
 sg13g2_a21oi_1 _2376_ (.A1(net108),
    .A2(net70),
    .Y(_0601_),
    .B1(\rsa_unit_i.P_i[0] ));
 sg13g2_and2_1 _2377_ (.A(net108),
    .B(\rsa_unit_i.R_i[0] ),
    .X(_0602_));
 sg13g2_a22oi_1 _2378_ (.Y(_0603_),
    .B1(_0602_),
    .B2(net70),
    .A2(_0375_),
    .A1(_0374_));
 sg13g2_or2_1 _2379_ (.X(_0604_),
    .B(_0603_),
    .A(_0601_));
 sg13g2_buf_1 _2380_ (.A(_0604_),
    .X(_0605_));
 sg13g2_inv_1 _2381_ (.Y(_0606_),
    .A(\rsa_unit_i.P_i[0] ));
 sg13g2_nand3_1 _2382_ (.B(\rsa_spi_wrapper_i.config_regs[33] ),
    .C(net95),
    .A(_1342_),
    .Y(_0607_));
 sg13g2_nand3_1 _2383_ (.B(_1293_),
    .C(net95),
    .A(_1343_),
    .Y(_0608_));
 sg13g2_a221oi_1 _2384_ (.B2(_0608_),
    .C1(_0603_),
    .B1(_0607_),
    .A1(_0606_),
    .Y(_0609_),
    .A2(_0386_));
 sg13g2_a21o_1 _2385_ (.A2(_0605_),
    .A1(_0600_),
    .B1(_0609_),
    .X(_0610_));
 sg13g2_buf_1 _2386_ (.A(_0610_),
    .X(_0611_));
 sg13g2_nor2_2 _2387_ (.A(_0386_),
    .B(_0381_),
    .Y(_0612_));
 sg13g2_a22oi_1 _2388_ (.Y(_0613_),
    .B1(_0612_),
    .B2(_0396_),
    .A2(_0378_),
    .A1(net94));
 sg13g2_buf_1 _2389_ (.A(_0613_),
    .X(_0614_));
 sg13g2_xnor2_1 _2390_ (.Y(_0615_),
    .A(_0611_),
    .B(_0614_));
 sg13g2_inv_1 _2391_ (.Y(_0616_),
    .A(net93));
 sg13g2_nand2_2 _2392_ (.Y(_0617_),
    .A(net78),
    .B(\rsa_unit_i.mmm_multiply.adder2.fa_bit0.HA1.a ));
 sg13g2_nor2_1 _2393_ (.A(net97),
    .B(_0617_),
    .Y(_0618_));
 sg13g2_a21oi_1 _2394_ (.A1(net93),
    .A2(_0615_),
    .Y(_0619_),
    .B1(_0618_));
 sg13g2_nand2b_1 _2395_ (.Y(_0620_),
    .B(\rsa_unit_i.mmm_multiply.adder2.fa_bit0.HA1.a ),
    .A_N(_1342_));
 sg13g2_nand2_1 _2396_ (.Y(_0621_),
    .A(_1286_),
    .B(net93));
 sg13g2_o21ai_1 _2397_ (.B1(_0621_),
    .Y(_0622_),
    .A1(net93),
    .A2(_0620_));
 sg13g2_nand2b_1 _2398_ (.Y(_0623_),
    .B(_0622_),
    .A_N(net95));
 sg13g2_or4_1 _2399_ (.A(net78),
    .B(net95),
    .C(_0601_),
    .D(_0603_),
    .X(_0624_));
 sg13g2_and2_1 _2400_ (.A(_0623_),
    .B(_0624_),
    .X(_0625_));
 sg13g2_nand2_1 _2401_ (.Y(_0626_),
    .A(_0043_),
    .B(_0625_));
 sg13g2_inv_1 _2402_ (.Y(_0627_),
    .A(_0043_));
 sg13g2_nand2_1 _2403_ (.Y(_0628_),
    .A(_0623_),
    .B(_0624_));
 sg13g2_nand2_1 _2404_ (.Y(_0629_),
    .A(_0627_),
    .B(_0628_));
 sg13g2_nand2_1 _2405_ (.Y(_0630_),
    .A(_0626_),
    .B(_0629_));
 sg13g2_xnor2_1 _2406_ (.Y(_0631_),
    .A(_0619_),
    .B(_0630_));
 sg13g2_buf_1 _2407_ (.A(net64),
    .X(_0632_));
 sg13g2_nand2_1 _2408_ (.Y(_0633_),
    .A(\rsa_unit_i.mmm_multiply.adder2.fa_bit0.HA1.a ),
    .B(net50));
 sg13g2_o21ai_1 _2409_ (.B1(_0633_),
    .Y(_0245_),
    .A1(net25),
    .A2(_0631_));
 sg13g2_nor2_1 _2410_ (.A(_1386_),
    .B(_0617_),
    .Y(_0634_));
 sg13g2_inv_1 _2411_ (.Y(_0635_),
    .A(\rsa_unit_i.P_i[2] ));
 sg13g2_a21oi_1 _2412_ (.A1(net108),
    .A2(_0371_),
    .Y(_0636_),
    .B1(_0635_));
 sg13g2_a21oi_1 _2413_ (.A1(_0374_),
    .A2(_0375_),
    .Y(_0637_),
    .B1(_0029_));
 sg13g2_a22oi_1 _2414_ (.Y(_0638_),
    .B1(_0637_),
    .B2(_0372_),
    .A2(_0636_),
    .A1(_0381_));
 sg13g2_buf_1 _2415_ (.A(_0638_),
    .X(_0639_));
 sg13g2_inv_1 _2416_ (.Y(_0640_),
    .A(net42));
 sg13g2_nor2b_1 _2417_ (.A(_1342_),
    .B_N(net108),
    .Y(_0641_));
 sg13g2_nor2b_1 _2418_ (.A(_1342_),
    .B_N(\rsa_unit_i.P_i[0] ),
    .Y(_0642_));
 sg13g2_a21oi_1 _2419_ (.A1(net70),
    .A2(_0641_),
    .Y(_0643_),
    .B1(_0642_));
 sg13g2_inv_1 _2420_ (.Y(_0644_),
    .A(\rsa_unit_i.P_i[1] ));
 sg13g2_a21o_1 _2421_ (.A2(net70),
    .A1(net108),
    .B1(_0644_),
    .X(_0645_));
 sg13g2_nand4_1 _2422_ (.B(\rsa_unit_i.R_i[0] ),
    .C(_0396_),
    .A(net108),
    .Y(_0646_),
    .D(net70));
 sg13g2_mux2_1 _2423_ (.A0(_0645_),
    .A1(_0646_),
    .S(_0376_),
    .X(_0647_));
 sg13g2_o21ai_1 _2424_ (.B1(_1293_),
    .Y(_0648_),
    .A1(_0643_),
    .A2(_0647_));
 sg13g2_nor2b_1 _2425_ (.A(_1342_),
    .B_N(\rsa_unit_i.R_i[0] ),
    .Y(_0649_));
 sg13g2_a21oi_1 _2426_ (.A1(_0374_),
    .A2(_0375_),
    .Y(_0650_),
    .B1(_0027_));
 sg13g2_o21ai_1 _2427_ (.B1(net54),
    .Y(_0651_),
    .A1(_0649_),
    .A2(_0650_));
 sg13g2_a21oi_1 _2428_ (.A1(net108),
    .A2(net70),
    .Y(_0652_),
    .B1(_0644_));
 sg13g2_a21o_1 _2429_ (.A2(_0641_),
    .A1(net70),
    .B1(_0642_),
    .X(_0653_));
 sg13g2_o21ai_1 _2430_ (.B1(_0381_),
    .Y(_0654_),
    .A1(_0652_),
    .A2(_0653_));
 sg13g2_nand2_1 _2431_ (.Y(_0655_),
    .A(_0651_),
    .B(_0654_));
 sg13g2_nor2_1 _2432_ (.A(_1386_),
    .B(net78),
    .Y(_0656_));
 sg13g2_nand4_1 _2433_ (.B(_0648_),
    .C(_0655_),
    .A(_0640_),
    .Y(_0657_),
    .D(_0656_));
 sg13g2_inv_2 _2434_ (.Y(_0658_),
    .A(_1386_));
 sg13g2_nor3_1 _2435_ (.A(_0658_),
    .B(net78),
    .C(net42),
    .Y(_0659_));
 sg13g2_nand2b_1 _2436_ (.Y(_0660_),
    .B(_0659_),
    .A_N(_0648_));
 sg13g2_xor2_1 _2437_ (.B(_0605_),
    .A(net95),
    .X(_0661_));
 sg13g2_and3_1 _2438_ (.X(_0662_),
    .A(_1386_),
    .B(net93),
    .C(net42));
 sg13g2_nand4_1 _2439_ (.B(_0648_),
    .C(_0655_),
    .A(_0661_),
    .Y(_0663_),
    .D(_0662_));
 sg13g2_nand3_1 _2440_ (.B(_0660_),
    .C(_0663_),
    .A(_0657_),
    .Y(_0664_));
 sg13g2_nand3_1 _2441_ (.B(_0661_),
    .C(_0656_),
    .A(net42),
    .Y(_0665_));
 sg13g2_and2_1 _2442_ (.A(_0651_),
    .B(_0654_),
    .X(_0666_));
 sg13g2_nor2_1 _2443_ (.A(net78),
    .B(net42),
    .Y(_0667_));
 sg13g2_xnor2_1 _2444_ (.Y(_0668_),
    .A(net95),
    .B(_0605_));
 sg13g2_buf_1 _2445_ (.A(_0668_),
    .X(_0669_));
 sg13g2_a22oi_1 _2446_ (.Y(_0670_),
    .B1(_0667_),
    .B2(net34),
    .A2(_0659_),
    .A1(_0666_));
 sg13g2_o21ai_1 _2447_ (.B1(_0670_),
    .Y(_0671_),
    .A1(_0648_),
    .A2(_0665_));
 sg13g2_and4_1 _2448_ (.A(net42),
    .B(_0661_),
    .C(_0666_),
    .D(_0656_),
    .X(_0672_));
 sg13g2_nor4_2 _2449_ (.A(_0634_),
    .B(_0664_),
    .C(_0671_),
    .Y(_0673_),
    .D(_0672_));
 sg13g2_inv_1 _2450_ (.Y(_0674_),
    .A(_0045_));
 sg13g2_nand2_1 _2451_ (.Y(_0675_),
    .A(_0674_),
    .B(_0626_));
 sg13g2_a21oi_1 _2452_ (.A1(_0619_),
    .A2(_0629_),
    .Y(_0676_),
    .B1(_0675_));
 sg13g2_nand4_1 _2453_ (.B(_0611_),
    .C(_0614_),
    .A(net93),
    .Y(_0677_),
    .D(_0628_));
 sg13g2_or4_1 _2454_ (.A(net78),
    .B(_0611_),
    .C(_0614_),
    .D(_0625_),
    .X(_0678_));
 sg13g2_o21ai_1 _2455_ (.B1(_0628_),
    .Y(_0679_),
    .A1(_0627_),
    .A2(_0618_));
 sg13g2_nand4_1 _2456_ (.B(_0627_),
    .C(_0611_),
    .A(net93),
    .Y(_0680_),
    .D(_0614_));
 sg13g2_nand4_1 _2457_ (.B(_0678_),
    .C(_0679_),
    .A(_0677_),
    .Y(_0681_),
    .D(_0680_));
 sg13g2_inv_1 _2458_ (.Y(_0682_),
    .A(_0618_));
 sg13g2_nor2_1 _2459_ (.A(_0043_),
    .B(_0682_),
    .Y(_0683_));
 sg13g2_nor4_1 _2460_ (.A(net78),
    .B(_0043_),
    .C(_0611_),
    .D(_0614_),
    .Y(_0684_));
 sg13g2_nor4_2 _2461_ (.A(_0674_),
    .B(_0681_),
    .C(_0683_),
    .Y(_0685_),
    .D(_0684_));
 sg13g2_nor3_1 _2462_ (.A(_0673_),
    .B(_0676_),
    .C(_0685_),
    .Y(_0686_));
 sg13g2_o21ai_1 _2463_ (.B1(_0673_),
    .Y(_0687_),
    .A1(_0676_),
    .A2(_0685_));
 sg13g2_nand2b_1 _2464_ (.Y(_0688_),
    .B(_0687_),
    .A_N(_0686_));
 sg13g2_nand2_1 _2465_ (.Y(_0689_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[1].fa.HA1.a ),
    .B(net50));
 sg13g2_o21ai_1 _2466_ (.B1(_0689_),
    .Y(_0246_),
    .A1(net25),
    .A2(_0688_));
 sg13g2_a21o_1 _2467_ (.A2(_0629_),
    .A1(_0619_),
    .B1(_0675_),
    .X(_0690_));
 sg13g2_a21oi_1 _2468_ (.A1(_0673_),
    .A2(_0690_),
    .Y(_0691_),
    .B1(_0685_));
 sg13g2_inv_1 _2469_ (.Y(_0692_),
    .A(_0046_));
 sg13g2_nand2_1 _2470_ (.Y(_0693_),
    .A(net54),
    .B(net61));
 sg13g2_nand3_1 _2471_ (.B(_0386_),
    .C(_0381_),
    .A(\rsa_unit_i.P_i[3] ),
    .Y(_0694_));
 sg13g2_o21ai_1 _2472_ (.B1(_0694_),
    .Y(_0695_),
    .A1(_0031_),
    .A2(_0693_));
 sg13g2_nor2_1 _2473_ (.A(_0669_),
    .B(_0695_),
    .Y(_0696_));
 sg13g2_o21ai_1 _2474_ (.B1(net42),
    .Y(_0697_),
    .A1(_0643_),
    .A2(_0647_));
 sg13g2_a21oi_1 _2475_ (.A1(_1386_),
    .A2(_0639_),
    .Y(_0698_),
    .B1(_1293_));
 sg13g2_nor3_1 _2476_ (.A(net42),
    .B(_0643_),
    .C(_0647_),
    .Y(_0699_));
 sg13g2_a221oi_1 _2477_ (.B2(_0655_),
    .C1(_0699_),
    .B1(_0698_),
    .A1(_0658_),
    .Y(_0700_),
    .A2(_0697_));
 sg13g2_buf_1 _2478_ (.A(_0700_),
    .X(_0701_));
 sg13g2_mux2_1 _2479_ (.A0(_0695_),
    .A1(_0696_),
    .S(net30),
    .X(_0702_));
 sg13g2_buf_1 _2480_ (.A(_0070_),
    .X(_0703_));
 sg13g2_nor2_1 _2481_ (.A(net92),
    .B(_0616_),
    .Y(_0704_));
 sg13g2_buf_1 _2482_ (.A(net78),
    .X(_0705_));
 sg13g2_nor2_1 _2483_ (.A(_1402_),
    .B(_0705_),
    .Y(_0706_));
 sg13g2_mux2_1 _2484_ (.A0(_0696_),
    .A1(_0695_),
    .S(net30),
    .X(_0707_));
 sg13g2_nand3_1 _2485_ (.B(_0669_),
    .C(_0695_),
    .A(_0565_),
    .Y(_0708_));
 sg13g2_o21ai_1 _2486_ (.B1(_0708_),
    .Y(_0709_),
    .A1(net92),
    .A2(_0617_));
 sg13g2_a221oi_1 _2487_ (.B2(_0707_),
    .C1(_0709_),
    .B1(_0706_),
    .A1(_0702_),
    .Y(_0710_),
    .A2(_0704_));
 sg13g2_xnor2_1 _2488_ (.Y(_0711_),
    .A(_0692_),
    .B(_0710_));
 sg13g2_xnor2_1 _2489_ (.Y(_0712_),
    .A(_0691_),
    .B(_0711_));
 sg13g2_nand2_1 _2490_ (.Y(_0713_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[2].fa.HA1.a ),
    .B(net50));
 sg13g2_o21ai_1 _2491_ (.B1(_0713_),
    .Y(_0247_),
    .A1(net25),
    .A2(_0712_));
 sg13g2_nand2b_1 _2492_ (.Y(_0714_),
    .B(_0710_),
    .A_N(_0691_));
 sg13g2_inv_1 _2493_ (.Y(_0715_),
    .A(_0710_));
 sg13g2_a21o_1 _2494_ (.A2(_0715_),
    .A1(_0691_),
    .B1(_0692_),
    .X(_0716_));
 sg13g2_nand2_1 _2495_ (.Y(_0717_),
    .A(_0714_),
    .B(_0716_));
 sg13g2_nand3b_1 _2496_ (.B(net54),
    .C(_0376_),
    .Y(_0718_),
    .A_N(_0033_));
 sg13g2_nand3_1 _2497_ (.B(_0386_),
    .C(_0381_),
    .A(\rsa_unit_i.P_i[4] ),
    .Y(_0719_));
 sg13g2_nand2_2 _2498_ (.Y(_0720_),
    .A(_0718_),
    .B(_0719_));
 sg13g2_inv_1 _2499_ (.Y(_0721_),
    .A(_0031_));
 sg13g2_a22oi_1 _2500_ (.Y(_0722_),
    .B1(_0612_),
    .B2(_0721_),
    .A2(net39),
    .A1(\rsa_unit_i.P_i[3] ));
 sg13g2_a21o_1 _2501_ (.A2(net30),
    .A1(net92),
    .B1(_0722_),
    .X(_0723_));
 sg13g2_or2_1 _2502_ (.X(_0724_),
    .B(net30),
    .A(net92));
 sg13g2_and3_1 _2503_ (.X(_0725_),
    .A(_0720_),
    .B(_0723_),
    .C(_0724_));
 sg13g2_and2_1 _2504_ (.A(_0718_),
    .B(_0719_),
    .X(_0726_));
 sg13g2_nand2_1 _2505_ (.Y(_0727_),
    .A(_0661_),
    .B(_0726_));
 sg13g2_a21oi_1 _2506_ (.A1(_0723_),
    .A2(_0724_),
    .Y(_0728_),
    .B1(_0727_));
 sg13g2_buf_1 _2507_ (.A(_1419_),
    .X(_0729_));
 sg13g2_o21ai_1 _2508_ (.B1(net77),
    .Y(_0730_),
    .A1(_0725_),
    .A2(_0728_));
 sg13g2_a221oi_1 _2509_ (.B2(_0724_),
    .C1(net77),
    .B1(_0723_),
    .A1(_0718_),
    .Y(_0731_),
    .A2(_0719_));
 sg13g2_a21oi_1 _2510_ (.A1(net92),
    .A2(net30),
    .Y(_0732_),
    .B1(_0722_));
 sg13g2_nor3_1 _2511_ (.A(net77),
    .B(net34),
    .C(_0720_),
    .Y(_0733_));
 sg13g2_o21ai_1 _2512_ (.B1(_0733_),
    .Y(_0734_),
    .A1(net92),
    .A2(net30));
 sg13g2_nand2_1 _2513_ (.Y(_0735_),
    .A(net34),
    .B(_0720_));
 sg13g2_o21ai_1 _2514_ (.B1(_0735_),
    .Y(_0736_),
    .A1(_0732_),
    .A2(_0734_));
 sg13g2_nor2_1 _2515_ (.A(_0731_),
    .B(_0736_),
    .Y(_0737_));
 sg13g2_a21oi_1 _2516_ (.A1(_0730_),
    .A2(_0737_),
    .Y(_0738_),
    .B1(net66));
 sg13g2_nor2_1 _2517_ (.A(net77),
    .B(_0617_),
    .Y(_0739_));
 sg13g2_nor2_1 _2518_ (.A(_0738_),
    .B(_0739_),
    .Y(_0740_));
 sg13g2_xnor2_1 _2519_ (.Y(_0741_),
    .A(_0417_),
    .B(_0740_));
 sg13g2_xnor2_1 _2520_ (.Y(_0742_),
    .A(_0717_),
    .B(_0741_));
 sg13g2_nand2_1 _2521_ (.Y(_0743_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[3].fa.HA1.a ),
    .B(net50));
 sg13g2_o21ai_1 _2522_ (.B1(_0743_),
    .Y(_0248_),
    .A1(net25),
    .A2(_0742_));
 sg13g2_inv_1 _2523_ (.Y(_0744_),
    .A(_0048_));
 sg13g2_nor2b_1 _2524_ (.A(_0739_),
    .B_N(_0417_),
    .Y(_0745_));
 sg13g2_o21ai_1 _2525_ (.B1(net79),
    .Y(_0746_),
    .A1(_0731_),
    .A2(_0736_));
 sg13g2_nor2_1 _2526_ (.A(_1420_),
    .B(net66),
    .Y(_0747_));
 sg13g2_o21ai_1 _2527_ (.B1(_0747_),
    .Y(_0748_),
    .A1(_0725_),
    .A2(_0728_));
 sg13g2_nand3_1 _2528_ (.B(_0746_),
    .C(_0748_),
    .A(_0745_),
    .Y(_0749_));
 sg13g2_nand3_1 _2529_ (.B(_0716_),
    .C(_0749_),
    .A(_0714_),
    .Y(_0750_));
 sg13g2_nor2_1 _2530_ (.A(net66),
    .B(_0417_),
    .Y(_0751_));
 sg13g2_o21ai_1 _2531_ (.B1(_0751_),
    .Y(_0752_),
    .A1(_0731_),
    .A2(_0736_));
 sg13g2_nand2b_1 _2532_ (.Y(_0753_),
    .B(_0739_),
    .A_N(_0417_));
 sg13g2_nor3_1 _2533_ (.A(_1420_),
    .B(net66),
    .C(_0417_),
    .Y(_0754_));
 sg13g2_o21ai_1 _2534_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0725_),
    .A2(_0728_));
 sg13g2_and4_1 _2535_ (.A(_0750_),
    .B(_0752_),
    .C(_0753_),
    .D(_0755_),
    .X(_0756_));
 sg13g2_inv_1 _2536_ (.Y(_0757_),
    .A(_0035_));
 sg13g2_a22oi_1 _2537_ (.Y(_0758_),
    .B1(_0612_),
    .B2(_0757_),
    .A2(net39),
    .A1(\rsa_unit_i.P_i[5] ));
 sg13g2_buf_2 _2538_ (.A(_0758_),
    .X(_0759_));
 sg13g2_nand2_1 _2539_ (.Y(_0760_),
    .A(_1438_),
    .B(_0564_));
 sg13g2_nor2_1 _2540_ (.A(_0759_),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_nand2_1 _2541_ (.Y(_0762_),
    .A(_1437_),
    .B(_0564_));
 sg13g2_nor2_1 _2542_ (.A(_0759_),
    .B(_0762_),
    .Y(_0763_));
 sg13g2_a221oi_1 _2543_ (.B2(_1419_),
    .C1(_0722_),
    .B1(_0726_),
    .A1(_0070_),
    .Y(_0764_),
    .A2(_0701_));
 sg13g2_o21ai_1 _2544_ (.B1(_1402_),
    .Y(_0765_),
    .A1(_1420_),
    .A2(_0720_));
 sg13g2_nand2_1 _2545_ (.Y(_0766_),
    .A(_1420_),
    .B(_0720_));
 sg13g2_o21ai_1 _2546_ (.B1(_0766_),
    .Y(_0767_),
    .A1(net30),
    .A2(_0765_));
 sg13g2_nor2_1 _2547_ (.A(_0764_),
    .B(_0767_),
    .Y(_0768_));
 sg13g2_mux2_1 _2548_ (.A0(_0761_),
    .A1(_0763_),
    .S(_0768_),
    .X(_0769_));
 sg13g2_nand2_1 _2549_ (.Y(_0770_),
    .A(_0661_),
    .B(_0759_));
 sg13g2_nor4_1 _2550_ (.A(_0764_),
    .B(_0767_),
    .C(_0770_),
    .D(_0760_),
    .Y(_0771_));
 sg13g2_nor3_1 _2551_ (.A(_0768_),
    .B(_0770_),
    .C(_0762_),
    .Y(_0772_));
 sg13g2_nand3b_1 _2552_ (.B(net79),
    .C(net34),
    .Y(_0773_),
    .A_N(_0759_));
 sg13g2_o21ai_1 _2553_ (.B1(_0773_),
    .Y(_0774_),
    .A1(_1437_),
    .A2(_0617_));
 sg13g2_or4_1 _2554_ (.A(_0769_),
    .B(_0771_),
    .C(_0772_),
    .D(_0774_),
    .X(_0775_));
 sg13g2_buf_8 _2555_ (.A(_0775_),
    .X(_0776_));
 sg13g2_xnor2_1 _2556_ (.Y(_0777_),
    .A(_0756_),
    .B(_0776_));
 sg13g2_xnor2_1 _2557_ (.Y(_0778_),
    .A(_0744_),
    .B(_0777_));
 sg13g2_nand2_1 _2558_ (.Y(_0779_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[4].fa.HA1.a ),
    .B(net50));
 sg13g2_o21ai_1 _2559_ (.B1(_0779_),
    .Y(_0249_),
    .A1(net25),
    .A2(_0778_));
 sg13g2_nand3_1 _2560_ (.B(_0753_),
    .C(_0755_),
    .A(_0752_),
    .Y(_0780_));
 sg13g2_nor2_1 _2561_ (.A(_0780_),
    .B(_0776_),
    .Y(_0781_));
 sg13g2_nand4_1 _2562_ (.B(_0716_),
    .C(_0749_),
    .A(_0714_),
    .Y(_0782_),
    .D(_0776_));
 sg13g2_a21oi_1 _2563_ (.A1(_0780_),
    .A2(_0776_),
    .Y(_0783_),
    .B1(_0744_));
 sg13g2_a22oi_1 _2564_ (.Y(_0784_),
    .B1(_0782_),
    .B2(_0783_),
    .A2(_0781_),
    .A1(_0750_));
 sg13g2_nand2_1 _2565_ (.Y(_0785_),
    .A(\rsa_unit_i.P_i[6] ),
    .B(net39));
 sg13g2_o21ai_1 _2566_ (.B1(_0785_),
    .Y(_0786_),
    .A1(_0037_),
    .A2(_0693_));
 sg13g2_nand2_1 _2567_ (.Y(_0787_),
    .A(_1437_),
    .B(_0759_));
 sg13g2_o21ai_1 _2568_ (.B1(_0787_),
    .Y(_0788_),
    .A1(_0764_),
    .A2(_0767_));
 sg13g2_or2_1 _2569_ (.X(_0789_),
    .B(_0759_),
    .A(_1437_));
 sg13g2_buf_1 _2570_ (.A(_0789_),
    .X(_0790_));
 sg13g2_nor2_1 _2571_ (.A(_1452_),
    .B(net66),
    .Y(_0791_));
 sg13g2_and4_1 _2572_ (.A(_0786_),
    .B(_0788_),
    .C(_0790_),
    .D(_0791_),
    .X(_0792_));
 sg13g2_buf_1 _2573_ (.A(_0079_),
    .X(_0793_));
 sg13g2_nor4_1 _2574_ (.A(net91),
    .B(net66),
    .C(net34),
    .D(_0786_),
    .Y(_0794_));
 sg13g2_and3_1 _2575_ (.X(_0795_),
    .A(_0788_),
    .B(_0790_),
    .C(_0794_));
 sg13g2_nand3_1 _2576_ (.B(net79),
    .C(_0786_),
    .A(_1452_),
    .Y(_0796_));
 sg13g2_inv_1 _2577_ (.Y(_0797_),
    .A(_0037_));
 sg13g2_a22oi_1 _2578_ (.Y(_0798_),
    .B1(_0612_),
    .B2(_0797_),
    .A2(net39),
    .A1(\rsa_unit_i.P_i[6] ));
 sg13g2_nand3_1 _2579_ (.B(_0798_),
    .C(_0791_),
    .A(_0661_),
    .Y(_0799_));
 sg13g2_a22oi_1 _2580_ (.Y(_0800_),
    .B1(_0796_),
    .B2(_0799_),
    .A2(_0790_),
    .A1(_0788_));
 sg13g2_nand3_1 _2581_ (.B(net34),
    .C(_0786_),
    .A(net79),
    .Y(_0801_));
 sg13g2_o21ai_1 _2582_ (.B1(_0801_),
    .Y(_0802_),
    .A1(net91),
    .A2(_0617_));
 sg13g2_nor4_1 _2583_ (.A(_0792_),
    .B(_0795_),
    .C(_0800_),
    .D(_0802_),
    .Y(_0803_));
 sg13g2_and2_1 _2584_ (.A(_0049_),
    .B(_0803_),
    .X(_0804_));
 sg13g2_nor2_1 _2585_ (.A(_0049_),
    .B(_0803_),
    .Y(_0805_));
 sg13g2_or2_1 _2586_ (.X(_0806_),
    .B(_0805_),
    .A(_0804_));
 sg13g2_xor2_1 _2587_ (.B(_0806_),
    .A(_0784_),
    .X(_0807_));
 sg13g2_nand2_1 _2588_ (.Y(_0808_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[5].fa.HA1.a ),
    .B(net50));
 sg13g2_o21ai_1 _2589_ (.B1(_0808_),
    .Y(_0250_),
    .A1(net25),
    .A2(_0807_));
 sg13g2_a221oi_1 _2590_ (.B2(_0783_),
    .C1(_0804_),
    .B1(_0782_),
    .A1(_0750_),
    .Y(_0809_),
    .A2(_0781_));
 sg13g2_nor2_1 _2591_ (.A(_0805_),
    .B(_0809_),
    .Y(_0810_));
 sg13g2_nand3_1 _2592_ (.B(_0788_),
    .C(_0790_),
    .A(_0798_),
    .Y(_0811_));
 sg13g2_buf_1 _2593_ (.A(_0811_),
    .X(_0812_));
 sg13g2_a21oi_1 _2594_ (.A1(_1420_),
    .A2(_0720_),
    .Y(_0813_),
    .B1(_1438_));
 sg13g2_o21ai_1 _2595_ (.B1(_0813_),
    .Y(_0814_),
    .A1(net92),
    .A2(net30));
 sg13g2_nor2_1 _2596_ (.A(_1420_),
    .B(_0720_),
    .Y(_0815_));
 sg13g2_o21ai_1 _2597_ (.B1(_1437_),
    .Y(_0816_),
    .A1(_0759_),
    .A2(_0815_));
 sg13g2_o21ai_1 _2598_ (.B1(_0816_),
    .Y(_0817_),
    .A1(_0732_),
    .A2(_0814_));
 sg13g2_and2_1 _2599_ (.A(_0079_),
    .B(_0759_),
    .X(_0818_));
 sg13g2_nor2_1 _2600_ (.A(_1452_),
    .B(_0786_),
    .Y(_0819_));
 sg13g2_a221oi_1 _2601_ (.B2(_0768_),
    .C1(_0819_),
    .B1(_0818_),
    .A1(net91),
    .Y(_0820_),
    .A2(_0817_));
 sg13g2_nand2_1 _2602_ (.Y(_0821_),
    .A(\rsa_unit_i.P_i[7] ),
    .B(net39));
 sg13g2_o21ai_1 _2603_ (.B1(_0821_),
    .Y(_0822_),
    .A1(_0039_),
    .A2(_0693_));
 sg13g2_buf_1 _2604_ (.A(_0822_),
    .X(_0823_));
 sg13g2_nor2_1 _2605_ (.A(_0331_),
    .B(net66),
    .Y(_0824_));
 sg13g2_and4_1 _2606_ (.A(_0812_),
    .B(_0820_),
    .C(_0823_),
    .D(_0824_),
    .X(_0825_));
 sg13g2_nor2_1 _2607_ (.A(net34),
    .B(_0823_),
    .Y(_0826_));
 sg13g2_nand2_1 _2608_ (.Y(_0827_),
    .A(_0824_),
    .B(_0826_));
 sg13g2_a21oi_1 _2609_ (.A1(_0812_),
    .A2(_0820_),
    .Y(_0828_),
    .B1(_0827_));
 sg13g2_nor2_1 _2610_ (.A(_0332_),
    .B(net66),
    .Y(_0829_));
 sg13g2_nand2_1 _2611_ (.Y(_0830_),
    .A(_0823_),
    .B(_0829_));
 sg13g2_a21oi_1 _2612_ (.A1(_0812_),
    .A2(_0820_),
    .Y(_0831_),
    .B1(_0830_));
 sg13g2_and4_1 _2613_ (.A(_0812_),
    .B(_0820_),
    .C(_0826_),
    .D(_0829_),
    .X(_0832_));
 sg13g2_nor4_2 _2614_ (.A(_0825_),
    .B(_0828_),
    .C(_0831_),
    .Y(_0833_),
    .D(_0832_));
 sg13g2_nor2_1 _2615_ (.A(_0331_),
    .B(_0617_),
    .Y(_0834_));
 sg13g2_nand3_1 _2616_ (.B(net34),
    .C(_0823_),
    .A(net79),
    .Y(_0835_));
 sg13g2_nor2b_1 _2617_ (.A(_0834_),
    .B_N(_0835_),
    .Y(_0836_));
 sg13g2_and3_1 _2618_ (.X(_0837_),
    .A(_0050_),
    .B(_0833_),
    .C(_0836_));
 sg13g2_buf_8 _2619_ (.A(_0837_),
    .X(_0838_));
 sg13g2_a21oi_2 _2620_ (.B1(_0050_),
    .Y(_0839_),
    .A2(_0836_),
    .A1(_0833_));
 sg13g2_nor3_1 _2621_ (.A(_0810_),
    .B(_0838_),
    .C(_0839_),
    .Y(_0840_));
 sg13g2_o21ai_1 _2622_ (.B1(_0810_),
    .Y(_0841_),
    .A1(_0838_),
    .A2(_0839_));
 sg13g2_nand2b_1 _2623_ (.Y(_0842_),
    .B(_0841_),
    .A_N(_0840_));
 sg13g2_nand2_1 _2624_ (.Y(_0843_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[6].fa.HA1.a ),
    .B(net50));
 sg13g2_o21ai_1 _2625_ (.B1(_0843_),
    .Y(_0251_),
    .A1(net25),
    .A2(_0842_));
 sg13g2_nor3_1 _2626_ (.A(_0805_),
    .B(_0809_),
    .C(_0839_),
    .Y(_0844_));
 sg13g2_nor2_1 _2627_ (.A(_0838_),
    .B(_0844_),
    .Y(_0845_));
 sg13g2_a21oi_1 _2628_ (.A1(_0788_),
    .A2(_0790_),
    .Y(_0846_),
    .B1(_0798_));
 sg13g2_a221oi_1 _2629_ (.B2(_0332_),
    .C1(_0846_),
    .B1(_0823_),
    .A1(_1452_),
    .Y(_0847_),
    .A2(_0812_));
 sg13g2_o21ai_1 _2630_ (.B1(_0385_),
    .Y(_0848_),
    .A1(_0705_),
    .A2(_0605_));
 sg13g2_and2_1 _2631_ (.A(_0624_),
    .B(_0848_),
    .X(_0849_));
 sg13g2_o21ai_1 _2632_ (.B1(_0849_),
    .Y(_0850_),
    .A1(_0332_),
    .A2(_0823_));
 sg13g2_inv_1 _2633_ (.Y(_0851_),
    .A(_0041_));
 sg13g2_a22oi_1 _2634_ (.Y(_0852_),
    .B1(_0612_),
    .B2(_0851_),
    .A2(_0379_),
    .A1(\rsa_unit_i.P_i[8] ));
 sg13g2_o21ai_1 _2635_ (.B1(_0852_),
    .Y(_0853_),
    .A1(_0847_),
    .A2(_0850_));
 sg13g2_or3_1 _2636_ (.A(_0847_),
    .B(_0850_),
    .C(_0852_),
    .X(_0854_));
 sg13g2_and3_1 _2637_ (.X(_0855_),
    .A(net79),
    .B(_0853_),
    .C(_0854_));
 sg13g2_buf_8 _2638_ (.A(_0855_),
    .X(_0856_));
 sg13g2_xnor2_1 _2639_ (.Y(_0857_),
    .A(_0051_),
    .B(_0856_));
 sg13g2_xnor2_1 _2640_ (.Y(_0858_),
    .A(_0845_),
    .B(_0857_));
 sg13g2_nand2_1 _2641_ (.Y(_0859_),
    .A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[7].fa.HA1.a ),
    .B(net50));
 sg13g2_o21ai_1 _2642_ (.B1(_0859_),
    .Y(_0252_),
    .A1(net25),
    .A2(_0858_));
 sg13g2_and2_1 _2643_ (.A(\rsa_unit_i.mmm_multiply.adder2.gen_fa[8].fa.HA1.a ),
    .B(net64),
    .X(_0860_));
 sg13g2_nor2b_1 _2644_ (.A(_0856_),
    .B_N(_0051_),
    .Y(_0861_));
 sg13g2_nor4_1 _2645_ (.A(_0805_),
    .B(_0809_),
    .C(_0839_),
    .D(_0856_),
    .Y(_0862_));
 sg13g2_nor2b_1 _2646_ (.A(_0856_),
    .B_N(_0838_),
    .Y(_0863_));
 sg13g2_nor3_1 _2647_ (.A(_0861_),
    .B(_0862_),
    .C(_0863_),
    .Y(_0864_));
 sg13g2_o21ai_1 _2648_ (.B1(_0051_),
    .Y(_0865_),
    .A1(_0838_),
    .A2(_0844_));
 sg13g2_a22oi_1 _2649_ (.Y(_0866_),
    .B1(_0612_),
    .B2(_0443_),
    .A2(_0379_),
    .A1(\rsa_unit_i.P_i[9] ));
 sg13g2_xor2_1 _2650_ (.B(_0866_),
    .A(_0854_),
    .X(_0867_));
 sg13g2_a21oi_1 _2651_ (.A1(net79),
    .A2(_0867_),
    .Y(_0868_),
    .B1(_0597_));
 sg13g2_and3_1 _2652_ (.X(_0869_),
    .A(_0864_),
    .B(_0865_),
    .C(_0868_));
 sg13g2_nand2_1 _2653_ (.Y(_0870_),
    .A(net79),
    .B(_0867_));
 sg13g2_or2_1 _2654_ (.X(_0871_),
    .B(_0870_),
    .A(_0597_));
 sg13g2_a21oi_1 _2655_ (.A1(_0864_),
    .A2(_0865_),
    .Y(_0872_),
    .B1(_0871_));
 sg13g2_or3_1 _2656_ (.A(_0860_),
    .B(_0869_),
    .C(_0872_),
    .X(_0253_));
 sg13g2_mux2_1 _2657_ (.A0(_0083_),
    .A1(_0452_),
    .S(net68),
    .X(_0873_));
 sg13g2_buf_1 _2658_ (.A(\rsa_unit_i.mmm_square.A_bit ),
    .X(_0874_));
 sg13g2_buf_8 _2659_ (.A(_0874_),
    .X(_0875_));
 sg13g2_nand2_1 _2660_ (.Y(_0876_),
    .A(_0875_),
    .B(_0632_));
 sg13g2_o21ai_1 _2661_ (.B1(_0876_),
    .Y(_0264_),
    .A1(_0558_),
    .A2(_0873_));
 sg13g2_mux2_1 _2662_ (.A0(_0086_),
    .A1(_0458_),
    .S(net68),
    .X(_0877_));
 sg13g2_nand2_1 _2663_ (.Y(_0878_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[1] ),
    .B(_0632_));
 sg13g2_o21ai_1 _2664_ (.B1(_0878_),
    .Y(_0265_),
    .A1(net31),
    .A2(_0877_));
 sg13g2_nor2_1 _2665_ (.A(_0089_),
    .B(_0569_),
    .Y(_0879_));
 sg13g2_a21oi_1 _2666_ (.A1(_0464_),
    .A2(_0569_),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_buf_1 _2667_ (.A(net64),
    .X(_0881_));
 sg13g2_nand2_1 _2668_ (.Y(_0882_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[2] ),
    .B(net49));
 sg13g2_o21ai_1 _2669_ (.B1(_0882_),
    .Y(_0266_),
    .A1(net31),
    .A2(_0880_));
 sg13g2_mux2_1 _2670_ (.A0(_0092_),
    .A1(_0468_),
    .S(net68),
    .X(_0883_));
 sg13g2_nand2_1 _2671_ (.Y(_0884_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[3] ),
    .B(net49));
 sg13g2_o21ai_1 _2672_ (.B1(_0884_),
    .Y(_0267_),
    .A1(net31),
    .A2(_0883_));
 sg13g2_mux2_1 _2673_ (.A0(_0095_),
    .A1(_0475_),
    .S(net68),
    .X(_0885_));
 sg13g2_nand2_1 _2674_ (.Y(_0886_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[4] ),
    .B(net49));
 sg13g2_o21ai_1 _2675_ (.B1(_0886_),
    .Y(_0268_),
    .A1(net31),
    .A2(_0885_));
 sg13g2_mux2_1 _2676_ (.A0(_0098_),
    .A1(_0483_),
    .S(net68),
    .X(_0887_));
 sg13g2_nand2_1 _2677_ (.Y(_0888_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[5] ),
    .B(net49));
 sg13g2_o21ai_1 _2678_ (.B1(_0888_),
    .Y(_0269_),
    .A1(net31),
    .A2(_0887_));
 sg13g2_mux2_1 _2679_ (.A0(_0101_),
    .A1(_0488_),
    .S(net68),
    .X(_0889_));
 sg13g2_nand2_1 _2680_ (.Y(_0890_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[6] ),
    .B(net49));
 sg13g2_o21ai_1 _2681_ (.B1(_0890_),
    .Y(_0270_),
    .A1(_0558_),
    .A2(_0889_));
 sg13g2_mux2_1 _2682_ (.A0(_0104_),
    .A1(_0492_),
    .S(_0562_),
    .X(_0891_));
 sg13g2_nand2_1 _2683_ (.Y(_0892_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[7] ),
    .B(_0881_));
 sg13g2_o21ai_1 _2684_ (.B1(_0892_),
    .Y(_0271_),
    .A1(net31),
    .A2(_0891_));
 sg13g2_inv_1 _2685_ (.Y(_0893_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[9] ));
 sg13g2_nand2_1 _2686_ (.Y(_0894_),
    .A(\rsa_unit_i.P_i[8] ),
    .B(net52));
 sg13g2_mux2_1 _2687_ (.A0(_0893_),
    .A1(_0894_),
    .S(_0562_),
    .X(_0895_));
 sg13g2_nand2_1 _2688_ (.Y(_0896_),
    .A(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[8] ),
    .B(net49));
 sg13g2_o21ai_1 _2689_ (.B1(_0896_),
    .Y(_0272_),
    .A1(net31),
    .A2(_0895_));
 sg13g2_nand4_1 _2690_ (.B(net65),
    .C(net43),
    .A(\rsa_unit_i.P_i[9] ),
    .Y(_0897_),
    .D(_0568_));
 sg13g2_o21ai_1 _2691_ (.B1(_0897_),
    .Y(_0273_),
    .A1(_0893_),
    .A2(net65));
 sg13g2_inv_1 _2692_ (.Y(_0898_),
    .A(net90));
 sg13g2_buf_1 _2693_ (.A(_0108_),
    .X(_0899_));
 sg13g2_inv_1 _2694_ (.Y(_0900_),
    .A(_0899_));
 sg13g2_buf_1 _2695_ (.A(\rsa_unit_i.mmm_square.adder2.fa_bit0.HA1.a ),
    .X(_0901_));
 sg13g2_nand2_1 _2696_ (.Y(_0902_),
    .A(_1280_),
    .B(_1287_));
 sg13g2_o21ai_1 _2697_ (.B1(net97),
    .Y(_0903_),
    .A1(net89),
    .A2(_0902_));
 sg13g2_nand2b_1 _2698_ (.Y(_0904_),
    .B(net83),
    .A_N(_0899_));
 sg13g2_a22oi_1 _2699_ (.Y(_0905_),
    .B1(_0904_),
    .B2(_1281_),
    .A2(_0903_),
    .A1(_0900_));
 sg13g2_nor2b_1 _2700_ (.A(_0449_),
    .B_N(_1286_),
    .Y(_0906_));
 sg13g2_nor2_1 _2701_ (.A(net94),
    .B(_0906_),
    .Y(_0907_));
 sg13g2_nand3b_1 _2702_ (.B(net83),
    .C(net94),
    .Y(_0908_),
    .A_N(net89));
 sg13g2_a21oi_1 _2703_ (.A1(net97),
    .A2(_0908_),
    .Y(_0909_),
    .B1(_0449_));
 sg13g2_nor3_1 _2704_ (.A(net55),
    .B(_0907_),
    .C(_0909_),
    .Y(_0910_));
 sg13g2_a21oi_1 _2705_ (.A1(_0362_),
    .A2(_0905_),
    .Y(_0911_),
    .B1(_0910_));
 sg13g2_mux2_1 _2706_ (.A0(_1280_),
    .A1(net94),
    .S(_0472_),
    .X(_0912_));
 sg13g2_inv_1 _2707_ (.Y(_0913_),
    .A(net89));
 sg13g2_a21oi_1 _2708_ (.A1(net97),
    .A2(_0912_),
    .Y(_0914_),
    .B1(_0913_));
 sg13g2_nor3_1 _2709_ (.A(net75),
    .B(_0911_),
    .C(_0914_),
    .Y(_0915_));
 sg13g2_nor3_1 _2710_ (.A(_1280_),
    .B(_0899_),
    .C(net83),
    .Y(_0916_));
 sg13g2_a21oi_1 _2711_ (.A1(_1280_),
    .A2(_1287_),
    .Y(_0917_),
    .B1(_0916_));
 sg13g2_nor3_1 _2712_ (.A(_0449_),
    .B(net94),
    .C(net83),
    .Y(_0918_));
 sg13g2_a221oi_1 _2713_ (.B2(net69),
    .C1(_0918_),
    .B1(_0446_),
    .A1(_0460_),
    .Y(_0919_),
    .A2(net83));
 sg13g2_a21oi_1 _2714_ (.A1(_0362_),
    .A2(_0917_),
    .Y(_0920_),
    .B1(_0919_));
 sg13g2_nor3_1 _2715_ (.A(net97),
    .B(net75),
    .C(_0901_),
    .Y(_0921_));
 sg13g2_xnor2_1 _2716_ (.Y(_0922_),
    .A(_1280_),
    .B(_0899_));
 sg13g2_xnor2_1 _2717_ (.Y(_0923_),
    .A(_0449_),
    .B(_0460_));
 sg13g2_mux2_1 _2718_ (.A0(_0922_),
    .A1(_0923_),
    .S(_0473_),
    .X(_0924_));
 sg13g2_nand2_1 _2719_ (.Y(_0925_),
    .A(_1363_),
    .B(net89));
 sg13g2_a21oi_1 _2720_ (.A1(net90),
    .A2(_0924_),
    .Y(_0926_),
    .B1(_0925_));
 sg13g2_a21o_1 _2721_ (.A2(_0921_),
    .A1(_0920_),
    .B1(_0926_),
    .X(_0927_));
 sg13g2_nor2_1 _2722_ (.A(_0915_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_nor2_1 _2723_ (.A(_1342_),
    .B(net90),
    .Y(_0929_));
 sg13g2_and2_1 _2724_ (.A(net83),
    .B(net90),
    .X(_0930_));
 sg13g2_o21ai_1 _2725_ (.B1(net89),
    .Y(_0931_),
    .A1(_0929_),
    .A2(_0930_));
 sg13g2_nor3_1 _2726_ (.A(_0900_),
    .B(_0358_),
    .C(_0360_),
    .Y(_0932_));
 sg13g2_nor2_1 _2727_ (.A(_0451_),
    .B(_0932_),
    .Y(_0933_));
 sg13g2_nand3b_1 _2728_ (.B(_0874_),
    .C(_0933_),
    .Y(_0934_),
    .A_N(net83));
 sg13g2_a21oi_1 _2729_ (.A1(_0931_),
    .A2(_0934_),
    .Y(_0935_),
    .B1(_0109_));
 sg13g2_xor2_1 _2730_ (.B(_0935_),
    .A(_0107_),
    .X(_0936_));
 sg13g2_xnor2_1 _2731_ (.Y(_0937_),
    .A(_0928_),
    .B(_0936_));
 sg13g2_buf_1 _2732_ (.A(net89),
    .X(_0938_));
 sg13g2_nand2_1 _2733_ (.Y(_0939_),
    .A(_0938_),
    .B(_0881_));
 sg13g2_o21ai_1 _2734_ (.B1(_0939_),
    .Y(_0274_),
    .A1(_0599_),
    .A2(_0937_));
 sg13g2_nand3b_1 _2735_ (.B(_1286_),
    .C(net97),
    .Y(_0940_),
    .A_N(_0899_));
 sg13g2_a21o_1 _2736_ (.A2(_0940_),
    .A1(_1293_),
    .B1(_1281_),
    .X(_0941_));
 sg13g2_nand4_1 _2737_ (.B(_1281_),
    .C(_0900_),
    .A(_1363_),
    .Y(_0942_),
    .D(_1286_));
 sg13g2_and3_1 _2738_ (.X(_0943_),
    .A(_0111_),
    .B(_0446_),
    .C(net69));
 sg13g2_buf_8 _2739_ (.A(_0943_),
    .X(_0944_));
 sg13g2_nand3_1 _2740_ (.B(_0942_),
    .C(_0944_),
    .A(_0941_),
    .Y(_0945_));
 sg13g2_a21oi_1 _2741_ (.A1(net94),
    .A2(\rsa_spi_wrapper_i.config_regs[33] ),
    .Y(_0946_),
    .B1(_0450_));
 sg13g2_a21oi_1 _2742_ (.A1(_0463_),
    .A2(_0946_),
    .Y(_0947_),
    .B1(_0898_));
 sg13g2_o21ai_1 _2743_ (.B1(_0947_),
    .Y(_0948_),
    .A1(_0900_),
    .A2(_0945_));
 sg13g2_nand3_1 _2744_ (.B(_0938_),
    .C(_0948_),
    .A(_0658_),
    .Y(_0949_));
 sg13g2_xnor2_1 _2745_ (.Y(_0950_),
    .A(net97),
    .B(\rsa_unit_i.P_i[1] ));
 sg13g2_a22oi_1 _2746_ (.Y(_0951_),
    .B1(_0906_),
    .B2(_0950_),
    .A2(\rsa_spi_wrapper_i.config_regs[33] ),
    .A1(net94));
 sg13g2_nand3b_1 _2747_ (.B(_0090_),
    .C(net52),
    .Y(_0952_),
    .A_N(_0951_));
 sg13g2_a21oi_1 _2748_ (.A1(_1293_),
    .A2(_0940_),
    .Y(_0953_),
    .B1(_1281_));
 sg13g2_nor3_1 _2749_ (.A(_1362_),
    .B(_1280_),
    .C(_0904_),
    .Y(_0954_));
 sg13g2_o21ai_1 _2750_ (.B1(_0944_),
    .Y(_0955_),
    .A1(_0953_),
    .A2(_0954_));
 sg13g2_a21oi_1 _2751_ (.A1(_0952_),
    .A2(_0955_),
    .Y(_0956_),
    .B1(_0658_));
 sg13g2_o21ai_1 _2752_ (.B1(_0449_),
    .Y(_0957_),
    .A1(_0358_),
    .A2(_0360_));
 sg13g2_nand3_1 _2753_ (.B(_0446_),
    .C(net69),
    .A(_0899_),
    .Y(_0958_));
 sg13g2_a21oi_2 _2754_ (.B1(_0913_),
    .Y(_0959_),
    .A2(_0958_),
    .A1(_0957_));
 sg13g2_a221oi_1 _2755_ (.B2(_0958_),
    .C1(_0944_),
    .B1(_0957_),
    .A1(_0090_),
    .Y(_0960_),
    .A2(_0472_));
 sg13g2_nor4_1 _2756_ (.A(_0451_),
    .B(_0463_),
    .C(_0932_),
    .D(_0944_),
    .Y(_0961_));
 sg13g2_mux2_1 _2757_ (.A0(_0960_),
    .A1(_0961_),
    .S(_0901_),
    .X(_0962_));
 sg13g2_a21o_1 _2758_ (.A2(_0959_),
    .A1(_0956_),
    .B1(_0962_),
    .X(_0963_));
 sg13g2_nor3_1 _2759_ (.A(_0462_),
    .B(net55),
    .C(_0951_),
    .Y(_0964_));
 sg13g2_nand3_1 _2760_ (.B(_0446_),
    .C(net69),
    .A(_0111_),
    .Y(_0965_));
 sg13g2_a21oi_1 _2761_ (.A1(_0941_),
    .A2(_0942_),
    .Y(_0966_),
    .B1(_0965_));
 sg13g2_nor3_1 _2762_ (.A(net89),
    .B(_0451_),
    .C(_0932_),
    .Y(_0967_));
 sg13g2_buf_1 _2763_ (.A(_0967_),
    .X(_0968_));
 sg13g2_o21ai_1 _2764_ (.B1(_0968_),
    .Y(_0969_),
    .A1(_0964_),
    .A2(_0966_));
 sg13g2_and2_1 _2765_ (.A(_0462_),
    .B(_0951_),
    .X(_0970_));
 sg13g2_nor2_1 _2766_ (.A(_0111_),
    .B(_0472_),
    .Y(_0971_));
 sg13g2_nor2_1 _2767_ (.A(_0953_),
    .B(_0954_),
    .Y(_0972_));
 sg13g2_a221oi_1 _2768_ (.B2(_0972_),
    .C1(_0658_),
    .B1(_0971_),
    .A1(net52),
    .Y(_0973_),
    .A2(_0970_));
 sg13g2_nor3_1 _2769_ (.A(_0953_),
    .B(_0954_),
    .C(_0965_),
    .Y(_0974_));
 sg13g2_a221oi_1 _2770_ (.B2(_0950_),
    .C1(_0462_),
    .B1(_0906_),
    .A1(\rsa_unit_i.P_i[1] ),
    .Y(_0975_),
    .A2(\rsa_spi_wrapper_i.config_regs[33] ));
 sg13g2_and2_1 _2771_ (.A(net52),
    .B(_0975_),
    .X(_0976_));
 sg13g2_o21ai_1 _2772_ (.B1(_0968_),
    .Y(_0977_),
    .A1(_0974_),
    .A2(_0976_));
 sg13g2_nor2_1 _2773_ (.A(net55),
    .B(_0951_),
    .Y(_0978_));
 sg13g2_nand2_1 _2774_ (.Y(_0979_),
    .A(_0941_),
    .B(_0942_));
 sg13g2_a221oi_1 _2775_ (.B2(_0979_),
    .C1(_1386_),
    .B1(_0971_),
    .A1(_0462_),
    .Y(_0980_),
    .A2(_0978_));
 sg13g2_a22oi_1 _2776_ (.Y(_0981_),
    .B1(_0977_),
    .B2(_0980_),
    .A2(_0973_),
    .A1(_0969_));
 sg13g2_o21ai_1 _2777_ (.B1(net76),
    .Y(_0982_),
    .A1(_0963_),
    .A2(_0981_));
 sg13g2_nand2_1 _2778_ (.Y(_0983_),
    .A(_0949_),
    .B(_0982_));
 sg13g2_o21ai_1 _2779_ (.B1(_0935_),
    .Y(_0984_),
    .A1(_0915_),
    .A2(_0927_));
 sg13g2_nor3_1 _2780_ (.A(_0915_),
    .B(_0927_),
    .C(_0935_),
    .Y(_0985_));
 sg13g2_a21oi_1 _2781_ (.A1(_0107_),
    .A2(_0984_),
    .Y(_0986_),
    .B1(_0985_));
 sg13g2_xnor2_1 _2782_ (.Y(_0987_),
    .A(_0110_),
    .B(_0986_));
 sg13g2_xnor2_1 _2783_ (.Y(_0988_),
    .A(_0983_),
    .B(_0987_));
 sg13g2_nand2_1 _2784_ (.Y(_0989_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[1].fa.HA1.a ),
    .B(net49));
 sg13g2_o21ai_1 _2785_ (.B1(_0989_),
    .Y(_0275_),
    .A1(_0599_),
    .A2(_0988_));
 sg13g2_nand3_1 _2786_ (.B(_0949_),
    .C(_0982_),
    .A(_0110_),
    .Y(_0990_));
 sg13g2_inv_1 _2787_ (.Y(_0991_),
    .A(_0110_));
 sg13g2_a21o_1 _2788_ (.A2(_0983_),
    .A1(_0991_),
    .B1(_0986_),
    .X(_0992_));
 sg13g2_nand2_1 _2789_ (.Y(_0993_),
    .A(_0990_),
    .B(_0992_));
 sg13g2_nor2_1 _2790_ (.A(net92),
    .B(_0913_),
    .Y(_0994_));
 sg13g2_nand2_2 _2791_ (.Y(_0995_),
    .A(_0957_),
    .B(_0958_));
 sg13g2_mux2_1 _2792_ (.A0(_0093_),
    .A1(_0113_),
    .S(_0361_),
    .X(_0996_));
 sg13g2_buf_1 _2793_ (.A(_0996_),
    .X(_0997_));
 sg13g2_a21oi_1 _2794_ (.A1(_0472_),
    .A2(_0975_),
    .Y(_0998_),
    .B1(_1386_));
 sg13g2_nor3_1 _2795_ (.A(_0090_),
    .B(_0361_),
    .C(_0951_),
    .Y(_0999_));
 sg13g2_a221oi_1 _2796_ (.B2(_0945_),
    .C1(_0999_),
    .B1(_0998_),
    .A1(_0979_),
    .Y(_1000_),
    .A2(_0971_));
 sg13g2_buf_2 _2797_ (.A(_1000_),
    .X(_1001_));
 sg13g2_nand3_1 _2798_ (.B(net40),
    .C(_1001_),
    .A(_0995_),
    .Y(_1002_));
 sg13g2_nand2_1 _2799_ (.Y(_1003_),
    .A(net76),
    .B(_1002_));
 sg13g2_o21ai_1 _2800_ (.B1(net40),
    .Y(_1004_),
    .A1(_0959_),
    .A2(net41));
 sg13g2_mux2_1 _2801_ (.A0(_1004_),
    .A1(net40),
    .S(_1001_),
    .X(_1005_));
 sg13g2_nor2_1 _2802_ (.A(_0959_),
    .B(net41),
    .Y(_1006_));
 sg13g2_nand2b_1 _2803_ (.Y(_1007_),
    .B(_1006_),
    .A_N(net40));
 sg13g2_o21ai_1 _2804_ (.B1(_1007_),
    .Y(_1008_),
    .A1(_1402_),
    .A2(_1005_));
 sg13g2_nand2_1 _2805_ (.Y(_1009_),
    .A(net41),
    .B(net40));
 sg13g2_mux2_1 _2806_ (.A0(_0997_),
    .A1(_1009_),
    .S(_1001_),
    .X(_1010_));
 sg13g2_nor3_1 _2807_ (.A(_0703_),
    .B(net75),
    .C(_1010_),
    .Y(_1011_));
 sg13g2_a221oi_1 _2808_ (.B2(net76),
    .C1(_1011_),
    .B1(_1008_),
    .A1(_0994_),
    .Y(_1012_),
    .A2(_1003_));
 sg13g2_xnor2_1 _2809_ (.Y(_1013_),
    .A(_0112_),
    .B(_1012_));
 sg13g2_xnor2_1 _2810_ (.Y(_1014_),
    .A(_0993_),
    .B(_1013_));
 sg13g2_nand2_1 _2811_ (.Y(_1015_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[2].fa.HA1.a ),
    .B(net49));
 sg13g2_o21ai_1 _2812_ (.B1(_1015_),
    .Y(_0276_),
    .A1(_0598_),
    .A2(_1014_));
 sg13g2_nor2_1 _2813_ (.A(_0112_),
    .B(_1012_),
    .Y(_1016_));
 sg13g2_a21oi_1 _2814_ (.A1(_0990_),
    .A2(_0992_),
    .Y(_1017_),
    .B1(_1016_));
 sg13g2_a21oi_2 _2815_ (.B1(_1017_),
    .Y(_1018_),
    .A2(_1012_),
    .A1(_0112_));
 sg13g2_mux2_1 _2816_ (.A0(_0096_),
    .A1(_0115_),
    .S(net55),
    .X(_1019_));
 sg13g2_buf_8 _2817_ (.A(_1019_),
    .X(_1020_));
 sg13g2_nand2_1 _2818_ (.Y(_1021_),
    .A(net41),
    .B(net37));
 sg13g2_nand2b_1 _2819_ (.Y(_1022_),
    .B(_1402_),
    .A_N(net40));
 sg13g2_and2_1 _2820_ (.A(_0070_),
    .B(net40),
    .X(_1023_));
 sg13g2_a21o_1 _2821_ (.A2(_1022_),
    .A1(_1001_),
    .B1(_1023_),
    .X(_1024_));
 sg13g2_buf_8 _2822_ (.A(_1024_),
    .X(_1025_));
 sg13g2_xnor2_1 _2823_ (.Y(_1026_),
    .A(_1420_),
    .B(_1025_));
 sg13g2_mux2_1 _2824_ (.A0(net37),
    .A1(_1021_),
    .S(_1026_),
    .X(_1027_));
 sg13g2_nor2_1 _2825_ (.A(net74),
    .B(_0933_),
    .Y(_1028_));
 sg13g2_a21oi_1 _2826_ (.A1(_0115_),
    .A2(net55),
    .Y(_1029_),
    .B1(_0474_));
 sg13g2_a21oi_1 _2827_ (.A1(_1001_),
    .A2(_1022_),
    .Y(_1030_),
    .B1(_1023_));
 sg13g2_nand2_1 _2828_ (.Y(_1031_),
    .A(_0995_),
    .B(net37));
 sg13g2_o21ai_1 _2829_ (.B1(net90),
    .Y(_1032_),
    .A1(_1030_),
    .A2(_1031_));
 sg13g2_nor2_1 _2830_ (.A(net77),
    .B(_0913_),
    .Y(_1033_));
 sg13g2_nand4_1 _2831_ (.B(net74),
    .C(_0995_),
    .A(net77),
    .Y(_1034_),
    .D(net37));
 sg13g2_nand3_1 _2832_ (.B(_0933_),
    .C(_1029_),
    .A(net74),
    .Y(_1035_));
 sg13g2_o21ai_1 _2833_ (.B1(_1035_),
    .Y(_1036_),
    .A1(_1025_),
    .A2(_1034_));
 sg13g2_a221oi_1 _2834_ (.B2(_1033_),
    .C1(_1036_),
    .B1(_1032_),
    .A1(_1028_),
    .Y(_1037_),
    .A2(_1029_));
 sg13g2_nor2_1 _2835_ (.A(net76),
    .B(_1033_),
    .Y(_1038_));
 sg13g2_a21oi_2 _2836_ (.B1(_1038_),
    .Y(_1039_),
    .A2(_1037_),
    .A1(_1027_));
 sg13g2_xnor2_1 _2837_ (.Y(_1040_),
    .A(_0114_),
    .B(_1039_));
 sg13g2_xnor2_1 _2838_ (.Y(_1041_),
    .A(_1018_),
    .B(_1040_));
 sg13g2_nand2_1 _2839_ (.Y(_1042_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[3].fa.HA1.a ),
    .B(net59));
 sg13g2_o21ai_1 _2840_ (.B1(_1042_),
    .Y(_0277_),
    .A1(net26),
    .A2(_1041_));
 sg13g2_a21o_1 _2841_ (.A2(_1039_),
    .A1(_1018_),
    .B1(_0471_),
    .X(_1043_));
 sg13g2_o21ai_1 _2842_ (.B1(_1043_),
    .Y(_1044_),
    .A1(_1018_),
    .A2(_1039_));
 sg13g2_nor2_1 _2843_ (.A(_1029_),
    .B(_1025_),
    .Y(_1045_));
 sg13g2_nand3_1 _2844_ (.B(_0446_),
    .C(net69),
    .A(_0117_),
    .Y(_1046_));
 sg13g2_nand2_1 _2845_ (.Y(_1047_),
    .A(_0482_),
    .B(_1046_));
 sg13g2_nor2_1 _2846_ (.A(_1437_),
    .B(_1047_),
    .Y(_1048_));
 sg13g2_a21oi_1 _2847_ (.A1(_0482_),
    .A2(_1046_),
    .Y(_1049_),
    .B1(_1438_));
 sg13g2_or2_1 _2848_ (.X(_1050_),
    .B(_1049_),
    .A(_1048_));
 sg13g2_nor2_1 _2849_ (.A(_1030_),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_o21ai_1 _2850_ (.B1(net77),
    .Y(_1052_),
    .A1(_1045_),
    .A2(_1051_));
 sg13g2_o21ai_1 _2851_ (.B1(_1025_),
    .Y(_1053_),
    .A1(net77),
    .A2(net37));
 sg13g2_or2_1 _2852_ (.X(_1054_),
    .B(net41),
    .A(_0959_));
 sg13g2_nand2_1 _2853_ (.Y(_1055_),
    .A(net90),
    .B(_1054_));
 sg13g2_a221oi_1 _2854_ (.B2(_1050_),
    .C1(_1055_),
    .B1(_1053_),
    .A1(_1020_),
    .Y(_1056_),
    .A2(_1051_));
 sg13g2_nand3_1 _2855_ (.B(_1020_),
    .C(_1047_),
    .A(_0729_),
    .Y(_1057_));
 sg13g2_nand2_1 _2856_ (.Y(_1058_),
    .A(net76),
    .B(_1057_));
 sg13g2_nand4_1 _2857_ (.B(net74),
    .C(_0933_),
    .A(net90),
    .Y(_1059_),
    .D(_1047_));
 sg13g2_a21oi_1 _2858_ (.A1(_0995_),
    .A2(_1047_),
    .Y(_1060_),
    .B1(net75));
 sg13g2_or2_1 _2859_ (.X(_1061_),
    .B(_1060_),
    .A(net74));
 sg13g2_nand3_1 _2860_ (.B(net89),
    .C(_0995_),
    .A(net90),
    .Y(_1062_));
 sg13g2_nand2b_1 _2861_ (.Y(_1063_),
    .B(_1062_),
    .A_N(net41));
 sg13g2_nand4_1 _2862_ (.B(net37),
    .C(_1048_),
    .A(_0729_),
    .Y(_1064_),
    .D(_1063_));
 sg13g2_nand3_1 _2863_ (.B(_1061_),
    .C(_1064_),
    .A(_1059_),
    .Y(_1065_));
 sg13g2_a221oi_1 _2864_ (.B2(_1437_),
    .C1(_1065_),
    .B1(_1058_),
    .A1(_1052_),
    .Y(_1066_),
    .A2(_1056_));
 sg13g2_buf_1 _2865_ (.A(_1066_),
    .X(_1067_));
 sg13g2_xnor2_1 _2866_ (.Y(_1068_),
    .A(_0479_),
    .B(_1067_));
 sg13g2_xnor2_1 _2867_ (.Y(_1069_),
    .A(_1044_),
    .B(_1068_));
 sg13g2_nand2_1 _2868_ (.Y(_1070_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[4].fa.HA1.a ),
    .B(net59));
 sg13g2_o21ai_1 _2869_ (.B1(_1070_),
    .Y(_0278_),
    .A1(net26),
    .A2(_1069_));
 sg13g2_o21ai_1 _2870_ (.B1(_1039_),
    .Y(_1071_),
    .A1(_0479_),
    .A2(_1067_));
 sg13g2_o21ai_1 _2871_ (.B1(_0471_),
    .Y(_1072_),
    .A1(_0479_),
    .A2(_1067_));
 sg13g2_a221oi_1 _2872_ (.B2(_1072_),
    .C1(_1017_),
    .B1(_1071_),
    .A1(_0112_),
    .Y(_1073_),
    .A2(_1012_));
 sg13g2_nand2_1 _2873_ (.Y(_1074_),
    .A(_0479_),
    .B(_1067_));
 sg13g2_o21ai_1 _2874_ (.B1(_1074_),
    .Y(_1075_),
    .A1(_0114_),
    .A2(_1071_));
 sg13g2_nor2_1 _2875_ (.A(_1073_),
    .B(_1075_),
    .Y(_1076_));
 sg13g2_a21oi_2 _2876_ (.B1(_0487_),
    .Y(_1077_),
    .A2(net55),
    .A1(_0021_));
 sg13g2_a21o_1 _2877_ (.A2(net40),
    .A1(_0703_),
    .B1(_1049_),
    .X(_1078_));
 sg13g2_a221oi_1 _2878_ (.B2(_1001_),
    .C1(_1078_),
    .B1(_1022_),
    .A1(_1419_),
    .Y(_1079_),
    .A2(net37));
 sg13g2_nor3_1 _2879_ (.A(_1419_),
    .B(net37),
    .C(_1049_),
    .Y(_1080_));
 sg13g2_or2_1 _2880_ (.X(_1081_),
    .B(_1080_),
    .A(_1048_));
 sg13g2_nor2_2 _2881_ (.A(_1079_),
    .B(_1081_),
    .Y(_1082_));
 sg13g2_nand3_1 _2882_ (.B(_1077_),
    .C(_1082_),
    .A(net91),
    .Y(_1083_));
 sg13g2_a21o_1 _2883_ (.A2(net55),
    .A1(_0021_),
    .B1(_0487_),
    .X(_1084_));
 sg13g2_buf_1 _2884_ (.A(_1084_),
    .X(_1085_));
 sg13g2_nand3_1 _2885_ (.B(net41),
    .C(_1085_),
    .A(net91),
    .Y(_1086_));
 sg13g2_nand4_1 _2886_ (.B(net74),
    .C(_0995_),
    .A(net91),
    .Y(_1087_),
    .D(_1085_));
 sg13g2_a21o_1 _2887_ (.A2(_1087_),
    .A1(_1086_),
    .B1(_1082_),
    .X(_1088_));
 sg13g2_nor2_1 _2888_ (.A(_0995_),
    .B(_1085_),
    .Y(_1089_));
 sg13g2_a22oi_1 _2889_ (.Y(_1090_),
    .B1(_1089_),
    .B2(net74),
    .A2(_1077_),
    .A1(_1028_));
 sg13g2_nor3_1 _2890_ (.A(_1077_),
    .B(_1079_),
    .C(_1081_),
    .Y(_1091_));
 sg13g2_and2_1 _2891_ (.A(net41),
    .B(_1091_),
    .X(_1092_));
 sg13g2_nor2_1 _2892_ (.A(_1085_),
    .B(_1082_),
    .Y(_1093_));
 sg13g2_o21ai_1 _2893_ (.B1(_1452_),
    .Y(_1094_),
    .A1(_1092_),
    .A2(_1093_));
 sg13g2_nand4_1 _2894_ (.B(_1088_),
    .C(_1090_),
    .A(_1083_),
    .Y(_1095_),
    .D(_1094_));
 sg13g2_a21oi_1 _2895_ (.A1(_0995_),
    .A2(_1091_),
    .Y(_1096_),
    .B1(net75));
 sg13g2_nor3_1 _2896_ (.A(net91),
    .B(_0913_),
    .C(_1096_),
    .Y(_1097_));
 sg13g2_a21o_1 _2897_ (.A2(_1095_),
    .A1(net76),
    .B1(_1097_),
    .X(_1098_));
 sg13g2_xor2_1 _2898_ (.B(_1098_),
    .A(_0020_),
    .X(_1099_));
 sg13g2_xnor2_1 _2899_ (.Y(_1100_),
    .A(_1076_),
    .B(_1099_));
 sg13g2_nand2_1 _2900_ (.Y(_1101_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[5].fa.HA1.a ),
    .B(net59));
 sg13g2_o21ai_1 _2901_ (.B1(_1101_),
    .Y(_0279_),
    .A1(net26),
    .A2(_1100_));
 sg13g2_o21ai_1 _2902_ (.B1(_1098_),
    .Y(_1102_),
    .A1(_1073_),
    .A2(_1075_));
 sg13g2_nor3_1 _2903_ (.A(_1073_),
    .B(_1075_),
    .C(_1098_),
    .Y(_1103_));
 sg13g2_a21oi_1 _2904_ (.A1(_0020_),
    .A2(_1102_),
    .Y(_1104_),
    .B1(_1103_));
 sg13g2_a21oi_2 _2905_ (.B1(_0491_),
    .Y(_1105_),
    .A2(net45),
    .A1(_0023_));
 sg13g2_nor3_1 _2906_ (.A(_1006_),
    .B(_1093_),
    .C(_1105_),
    .Y(_1106_));
 sg13g2_a21oi_1 _2907_ (.A1(net91),
    .A2(_1085_),
    .Y(_1107_),
    .B1(_1082_));
 sg13g2_o21ai_1 _2908_ (.B1(_1105_),
    .Y(_1108_),
    .A1(_1006_),
    .A2(_1107_));
 sg13g2_nand2b_1 _2909_ (.Y(_1109_),
    .B(_1108_),
    .A_N(_1106_));
 sg13g2_or2_1 _2910_ (.X(_1110_),
    .B(_1105_),
    .A(_1082_));
 sg13g2_nand3_1 _2911_ (.B(_1077_),
    .C(_1082_),
    .A(_1054_),
    .Y(_1111_));
 sg13g2_a21oi_1 _2912_ (.A1(_1110_),
    .A2(_1111_),
    .Y(_1112_),
    .B1(_0793_));
 sg13g2_nor3_1 _2913_ (.A(_0331_),
    .B(net75),
    .C(_1112_),
    .Y(_1113_));
 sg13g2_nor2_1 _2914_ (.A(_0332_),
    .B(net75),
    .Y(_1114_));
 sg13g2_nor2_1 _2915_ (.A(_0793_),
    .B(_1091_),
    .Y(_1115_));
 sg13g2_o21ai_1 _2916_ (.B1(_1054_),
    .Y(_1116_),
    .A1(_1093_),
    .A2(_1115_));
 sg13g2_xnor2_1 _2917_ (.Y(_1117_),
    .A(_1105_),
    .B(_1116_));
 sg13g2_nand2_1 _2918_ (.Y(_1118_),
    .A(net75),
    .B(net74));
 sg13g2_nand4_1 _2919_ (.B(net76),
    .C(_1077_),
    .A(_1452_),
    .Y(_1119_),
    .D(_1105_));
 sg13g2_a21oi_1 _2920_ (.A1(_1118_),
    .A2(_1119_),
    .Y(_1120_),
    .B1(_0331_));
 sg13g2_a221oi_1 _2921_ (.B2(_1117_),
    .C1(_1120_),
    .B1(_1114_),
    .A1(_1109_),
    .Y(_1121_),
    .A2(_1113_));
 sg13g2_xor2_1 _2922_ (.B(_1121_),
    .A(_0022_),
    .X(_1122_));
 sg13g2_xnor2_1 _2923_ (.Y(_1123_),
    .A(_1104_),
    .B(_1122_));
 sg13g2_nand2_1 _2924_ (.Y(_1124_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[6].fa.HA1.a ),
    .B(net59));
 sg13g2_o21ai_1 _2925_ (.B1(_1124_),
    .Y(_0280_),
    .A1(_0598_),
    .A2(_1123_));
 sg13g2_nand2_1 _2926_ (.Y(_1125_),
    .A(_0022_),
    .B(_1121_));
 sg13g2_nor2_1 _2927_ (.A(_0022_),
    .B(_1121_),
    .Y(_1126_));
 sg13g2_a21oi_2 _2928_ (.B1(_1126_),
    .Y(_1127_),
    .A2(_1125_),
    .A1(_1104_));
 sg13g2_nand2b_1 _2929_ (.Y(_1128_),
    .B(_0331_),
    .A_N(_1105_));
 sg13g2_o21ai_1 _2930_ (.B1(_1128_),
    .Y(_1129_),
    .A1(_1093_),
    .A2(_1115_));
 sg13g2_nand2_1 _2931_ (.Y(_1130_),
    .A(_0332_),
    .B(_1105_));
 sg13g2_a21oi_1 _2932_ (.A1(_1129_),
    .A2(_1130_),
    .Y(_1131_),
    .B1(_1006_));
 sg13g2_xnor2_1 _2933_ (.Y(_1132_),
    .A(_0894_),
    .B(_1131_));
 sg13g2_nand2_1 _2934_ (.Y(_1133_),
    .A(_0875_),
    .B(_1132_));
 sg13g2_xnor2_1 _2935_ (.Y(_1134_),
    .A(_0024_),
    .B(_1133_));
 sg13g2_xnor2_1 _2936_ (.Y(_1135_),
    .A(_1127_),
    .B(_1134_));
 sg13g2_nand2_1 _2937_ (.Y(_1136_),
    .A(\rsa_unit_i.mmm_square.adder2.gen_fa[7].fa.HA1.a ),
    .B(net59));
 sg13g2_o21ai_1 _2938_ (.B1(_1136_),
    .Y(_0281_),
    .A1(net26),
    .A2(_1135_));
 sg13g2_nand2_1 _2939_ (.Y(_1137_),
    .A(_0024_),
    .B(_1133_));
 sg13g2_nand2_1 _2940_ (.Y(_1138_),
    .A(\rsa_unit_i.P_i[8] ),
    .B(_1131_));
 sg13g2_xnor2_1 _2941_ (.Y(_1139_),
    .A(\rsa_unit_i.P_i[9] ),
    .B(_1138_));
 sg13g2_nand3_1 _2942_ (.B(net52),
    .C(_1139_),
    .A(net76),
    .Y(_1140_));
 sg13g2_nand2_1 _2943_ (.Y(_1141_),
    .A(_1137_),
    .B(_1140_));
 sg13g2_or3_1 _2944_ (.A(net26),
    .B(_1127_),
    .C(_1141_),
    .X(_1142_));
 sg13g2_nor2_1 _2945_ (.A(_0024_),
    .B(_1133_),
    .Y(_1143_));
 sg13g2_nor2b_1 _2946_ (.A(net26),
    .B_N(_1140_),
    .Y(_1144_));
 sg13g2_nor3_1 _2947_ (.A(net26),
    .B(_1137_),
    .C(_1140_),
    .Y(_1145_));
 sg13g2_a21oi_1 _2948_ (.A1(_1143_),
    .A2(_1144_),
    .Y(_1146_),
    .B1(_1145_));
 sg13g2_nor3_1 _2949_ (.A(_0597_),
    .B(_1143_),
    .C(_1140_),
    .Y(_1147_));
 sg13g2_a22oi_1 _2950_ (.Y(_1148_),
    .B1(_1127_),
    .B2(_1147_),
    .A2(_1187_),
    .A1(\rsa_unit_i.mmm_square.adder2.gen_fa[8].fa.HA1.a ));
 sg13g2_nand3_1 _2951_ (.B(_1146_),
    .C(_1148_),
    .A(_1142_),
    .Y(_0282_));
 sg13g2_nand2_1 _2952_ (.Y(_0119_),
    .A(_1156_),
    .B(\rsa_en_logic_i.state[0] ));
 sg13g2_nand3_1 _2953_ (.B(net87),
    .C(_1169_),
    .A(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ),
    .Y(_1149_));
 sg13g2_inv_1 _2954_ (.Y(_1150_),
    .A(_1194_));
 sg13g2_nand2b_1 _2955_ (.Y(_1151_),
    .B(_1163_),
    .A_N(_1165_));
 sg13g2_a22oi_1 _2956_ (.Y(_1152_),
    .B1(_1151_),
    .B2(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0] ),
    .A2(_1150_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_nor3_1 _2957_ (.A(_1197_),
    .B(_1193_),
    .C(_1312_),
    .Y(_1153_));
 sg13g2_o21ai_1 _2958_ (.B1(_1311_),
    .Y(_1154_),
    .A1(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0] ),
    .A2(_1153_));
 sg13g2_and3_1 _2959_ (.X(_0120_),
    .A(_1149_),
    .B(_1152_),
    .C(_1154_));
 sg13g2_dfrbp_1 _2960_ (.CLK(clknet_leaf_20_clk),
    .RESET_B(net144),
    .D(_0121_),
    .Q_N(\rsa_unit_i.rsa_control_fsm.state[0] ),
    .Q(_0118_));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _2963__155 (.L_HI(net155));
 sg13g2_buf_1 _2963_ (.A(net155),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2964_ (.A(net156),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2965_ (.A(net157),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2966_ (.A(net158),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2967_ (.A(net152),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2968_ (.A(net153),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2969_ (.A(net154),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2970_ (.A(net159),
    .X(uio_oe[7]));
 sg13g2_buf_1 _2971_ (.A(irq),
    .X(net9));
 sg13g2_buf_1 _2972_ (.A(ui_in[4]),
    .X(net10));
 sg13g2_buf_1 _2973_ (.A(ui_in[5]),
    .X(net11));
 sg13g2_buf_1 _2974_ (.A(\rsa_spi_wrapper_i.spi_miso ),
    .X(net12));
 sg13g2_buf_1 _2975_ (.A(ui_in[4]),
    .X(net13));
 sg13g2_buf_1 _2976_ (.A(ui_in[5]),
    .X(net14));
 sg13g2_buf_1 _2977_ (.A(ui_in[6]),
    .X(net15));
 sg13g2_buf_1 _2978_ (.A(ui_in[7]),
    .X(net16));
 sg13g2_buf_1 _2979_ (.A(\rsa_spi_wrapper_i.config_regs[56] ),
    .X(net17));
 sg13g2_buf_1 _2980_ (.A(\rsa_spi_wrapper_i.config_regs[57] ),
    .X(net18));
 sg13g2_buf_1 _2981_ (.A(\rsa_spi_wrapper_i.config_regs[58] ),
    .X(net19));
 sg13g2_buf_1 _2982_ (.A(\rsa_spi_wrapper_i.config_regs[59] ),
    .X(net20));
 sg13g2_buf_1 _2983_ (.A(\rsa_spi_wrapper_i.config_regs[60] ),
    .X(net21));
 sg13g2_buf_1 _2984_ (.A(\rsa_spi_wrapper_i.config_regs[61] ),
    .X(net22));
 sg13g2_buf_1 _2985_ (.A(\rsa_spi_wrapper_i.config_regs[62] ),
    .X(net23));
 sg13g2_buf_1 _2986_ (.A(\rsa_spi_wrapper_i.config_regs[63] ),
    .X(net24));
 sg13g2_dfrbp_1 \gpio_wrapper_i.gpio_start_cmd_i.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net147),
    .D(_0122_),
    .Q_N(_1575_),
    .Q(\gpio_wrapper_i.gpio_start_cmd_i.data_dly ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.gpio_stop_cmd_i.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net147),
    .D(_0123_),
    .Q_N(_1574_),
    .Q(\gpio_wrapper_i.gpio_stop_cmd_i.data_dly ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.sync_gpio_start.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net147),
    .D(_0124_),
    .Q_N(_1573_),
    .Q(\gpio_wrapper_i.sync_gpio_start.data_sync[1] ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.sync_gpio_start.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net148),
    .D(_0125_),
    .Q_N(_1572_),
    .Q(\gpio_wrapper_i.gpio_start_cmd_i.data ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.sync_gpio_stop.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net148),
    .D(_0126_),
    .Q_N(_1571_),
    .Q(\gpio_wrapper_i.sync_gpio_stop.data_sync[1] ));
 sg13g2_dfrbp_1 \gpio_wrapper_i.sync_gpio_stop.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net147),
    .D(_0127_),
    .Q_N(_1570_),
    .Q(\gpio_wrapper_i.gpio_stop_cmd_i.data ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.irq_reg$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net149),
    .D(_0128_),
    .Q_N(_0061_),
    .Q(irq));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[0]$_DFF_PN1_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net145),
    .D(_0119_),
    .Q_N(\rsa_en_logic_i.state[0] ),
    .Q(_1591_));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net145),
    .D(_0000_),
    .Q_N(_1576_),
    .Q(\rsa_en_logic_i.state[1] ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[2]$_DFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net144),
    .D(_0001_),
    .Q_N(_1577_),
    .Q(\rsa_en_logic_i.state[2] ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[3]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net145),
    .D(_0002_),
    .Q_N(_1578_),
    .Q(\rsa_en_logic_i.state[3] ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[4]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net145),
    .D(_0003_),
    .Q_N(_1579_),
    .Q(\rsa_en_logic_i.state[4] ));
 sg13g2_dfrbp_1 \rsa_en_logic_i.state[5]$_DFF_PN0_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net144),
    .D(_0004_),
    .Q_N(_0056_),
    .Q(\rsa_en_logic_i.state[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_start_cmd_i.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net147),
    .D(_0129_),
    .Q_N(_1569_),
    .Q(\rsa_spi_wrapper_i.spi_start_cmd_i.data_dly ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net147),
    .D(_0130_),
    .Q_N(_1568_),
    .Q(\rsa_spi_wrapper_i.spi_stop_cmd_i.data_dly ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net126),
    .D(_0131_),
    .Q_N(_0059_),
    .Q(\rsa_spi_wrapper_i.config_regs[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net124),
    .D(_0132_),
    .Q_N(_0063_),
    .Q(\rsa_spi_wrapper_i.config_regs[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net120),
    .D(_0133_),
    .Q_N(_0066_),
    .Q(\rsa_spi_wrapper_i.config_regs[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net118),
    .D(_0134_),
    .Q_N(_0069_),
    .Q(\rsa_spi_wrapper_i.config_regs[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net122),
    .D(_0135_),
    .Q_N(_0072_),
    .Q(\rsa_spi_wrapper_i.config_regs[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net124),
    .D(_0136_),
    .Q_N(_0075_),
    .Q(\rsa_spi_wrapper_i.config_regs[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net124),
    .D(_0137_),
    .Q_N(_0078_),
    .Q(\rsa_spi_wrapper_i.config_regs[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[0][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net120),
    .D(_0138_),
    .Q_N(_0081_),
    .Q(\rsa_spi_wrapper_i.config_regs[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net142),
    .D(_0139_),
    .Q_N(_1567_),
    .Q(\rsa_spi_wrapper_i.config_regs[8] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net142),
    .D(_0140_),
    .Q_N(_1566_),
    .Q(\rsa_spi_wrapper_i.config_regs[9] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net122),
    .D(_0141_),
    .Q_N(_1565_),
    .Q(\rsa_spi_wrapper_i.config_regs[10] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net118),
    .D(_0142_),
    .Q_N(_1564_),
    .Q(\rsa_spi_wrapper_i.config_regs[11] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net141),
    .D(_0143_),
    .Q_N(_1563_),
    .Q(\rsa_spi_wrapper_i.config_regs[12] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net122),
    .D(_0144_),
    .Q_N(_1562_),
    .Q(\rsa_spi_wrapper_i.config_regs[13] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net141),
    .D(_0145_),
    .Q_N(_1561_),
    .Q(\rsa_spi_wrapper_i.config_regs[14] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[1][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net118),
    .D(_0146_),
    .Q_N(_1560_),
    .Q(\rsa_spi_wrapper_i.config_regs[15] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net139),
    .D(_0147_),
    .Q_N(_0108_),
    .Q(\rsa_p[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net139),
    .D(_0148_),
    .Q_N(_1559_),
    .Q(\rsa_p[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net137),
    .D(_0149_),
    .Q_N(_0111_),
    .Q(\rsa_p[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net137),
    .D(_0150_),
    .Q_N(_0113_),
    .Q(\rsa_p[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net137),
    .D(_0151_),
    .Q_N(_0115_),
    .Q(\rsa_p[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net137),
    .D(_0152_),
    .Q_N(_0117_),
    .Q(\rsa_p[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net137),
    .D(_0153_),
    .Q_N(_0021_),
    .Q(\rsa_p[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[2][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net137),
    .D(_0154_),
    .Q_N(_0023_),
    .Q(\rsa_p[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net139),
    .D(_0155_),
    .Q_N(_1558_),
    .Q(\rsa_e[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net139),
    .D(_0156_),
    .Q_N(_1557_),
    .Q(\rsa_e[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net137),
    .D(_0157_),
    .Q_N(_1556_),
    .Q(\rsa_e[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net138),
    .D(_0158_),
    .Q_N(_1555_),
    .Q(\rsa_e[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net138),
    .D(_0159_),
    .Q_N(_1554_),
    .Q(\rsa_e[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net140),
    .D(_0160_),
    .Q_N(_1553_),
    .Q(\rsa_e[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net138),
    .D(_0161_),
    .Q_N(_1552_),
    .Q(\rsa_e[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[3][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net138),
    .D(_0162_),
    .Q_N(_1551_),
    .Q(\rsa_e[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net130),
    .D(_0163_),
    .Q_N(_0060_),
    .Q(\rsa_spi_wrapper_i.config_regs[32] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net130),
    .D(_0164_),
    .Q_N(_0064_),
    .Q(\rsa_spi_wrapper_i.config_regs[33] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net118),
    .D(_0165_),
    .Q_N(_0067_),
    .Q(\rsa_spi_wrapper_i.config_regs[34] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net128),
    .D(_0166_),
    .Q_N(_0070_),
    .Q(\rsa_spi_wrapper_i.config_regs[35] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net118),
    .D(_0167_),
    .Q_N(_0073_),
    .Q(\rsa_spi_wrapper_i.config_regs[36] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net118),
    .D(_0168_),
    .Q_N(_0076_),
    .Q(\rsa_spi_wrapper_i.config_regs[37] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net116),
    .D(_0169_),
    .Q_N(_0079_),
    .Q(\rsa_spi_wrapper_i.config_regs[38] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[4][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net118),
    .D(_0170_),
    .Q_N(_0082_),
    .Q(\rsa_spi_wrapper_i.config_regs[39] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net116),
    .D(_0171_),
    .Q_N(_0085_),
    .Q(\rsa_const[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net136),
    .D(_0172_),
    .Q_N(_0088_),
    .Q(\rsa_const[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net128),
    .D(_0173_),
    .Q_N(_0091_),
    .Q(\rsa_const[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net137),
    .D(_0174_),
    .Q_N(_0094_),
    .Q(\rsa_const[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net128),
    .D(_0175_),
    .Q_N(_0097_),
    .Q(\rsa_const[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net139),
    .D(_0176_),
    .Q_N(_0100_),
    .Q(\rsa_const[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net116),
    .D(_0177_),
    .Q_N(_0103_),
    .Q(\rsa_const[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[5][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net136),
    .D(_0178_),
    .Q_N(_0106_),
    .Q(\rsa_const[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net120),
    .D(_0179_),
    .Q_N(_1550_),
    .Q(\rsa_spi_wrapper_i.config_regs[48] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net121),
    .D(_0180_),
    .Q_N(_1549_),
    .Q(\rsa_spi_wrapper_i.config_regs[49] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net119),
    .D(_0181_),
    .Q_N(_1548_),
    .Q(\rsa_spi_wrapper_i.config_regs[50] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net119),
    .D(_0182_),
    .Q_N(_1547_),
    .Q(\rsa_spi_wrapper_i.config_regs[51] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net119),
    .D(_0183_),
    .Q_N(_1546_),
    .Q(\rsa_spi_wrapper_i.config_regs[52] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net119),
    .D(_0184_),
    .Q_N(_1545_),
    .Q(\rsa_spi_wrapper_i.config_regs[53] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net121),
    .D(_0185_),
    .Q_N(_1544_),
    .Q(\rsa_spi_wrapper_i.config_regs[54] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[6][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net119),
    .D(_0186_),
    .Q_N(_1543_),
    .Q(\rsa_spi_wrapper_i.config_regs[55] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net141),
    .D(_0187_),
    .Q_N(_1542_),
    .Q(\rsa_spi_wrapper_i.config_regs[56] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net141),
    .D(_0188_),
    .Q_N(_1541_),
    .Q(\rsa_spi_wrapper_i.config_regs[57] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net141),
    .D(_0189_),
    .Q_N(_1540_),
    .Q(\rsa_spi_wrapper_i.config_regs[58] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net127),
    .D(_0190_),
    .Q_N(_1539_),
    .Q(\rsa_spi_wrapper_i.config_regs[59] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net141),
    .D(_0191_),
    .Q_N(_1538_),
    .Q(\rsa_spi_wrapper_i.config_regs[60] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0192_),
    .Q_N(_1537_),
    .Q(\rsa_spi_wrapper_i.config_regs[61] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0193_),
    .Q_N(_1536_),
    .Q(\rsa_spi_wrapper_i.config_regs[62] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.config_mem[7][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0194_),
    .Q_N(_1535_),
    .Q(\rsa_spi_wrapper_i.config_regs[63] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.addr[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net126),
    .D(_0195_),
    .Q_N(_1534_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.addr[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net127),
    .D(_0196_),
    .Q_N(_1533_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.addr[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net127),
    .D(_0197_),
    .Q_N(_0053_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.addr[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net124),
    .D(_0198_),
    .Q_N(_1532_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_addr[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net124),
    .D(_0199_),
    .Q_N(_1531_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net124),
    .D(_0200_),
    .Q_N(_1530_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net122),
    .D(_0201_),
    .Q_N(_1529_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net122),
    .D(_0202_),
    .Q_N(_1528_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net122),
    .D(_0203_),
    .Q_N(_1527_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net122),
    .D(_0204_),
    .Q_N(_1526_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net125),
    .D(_0205_),
    .Q_N(_1525_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.data[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net123),
    .D(_0206_),
    .Q_N(_1524_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.dv$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net149),
    .D(_0207_),
    .Q_N(_1523_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.reg_data_o_vld ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net124),
    .D(_0208_),
    .Q_N(_1522_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.reg_rw ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rising_edge_detector_eof.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net147),
    .D(_0209_),
    .Q_N(_1521_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_sof.data_dly ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rising_edge_detector_spi_clk.data_dly$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net148),
    .D(_0210_),
    .Q_N(_1520_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.falling_edge_detector_spi_clk.data_dly ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net125),
    .D(_0211_),
    .Q_N(_1519_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net125),
    .D(_0212_),
    .Q_N(_1518_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net124),
    .D(_0213_),
    .Q_N(_1517_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net122),
    .D(_0214_),
    .Q_N(_1516_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net123),
    .D(_0215_),
    .Q_N(_1515_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net123),
    .D(_0216_),
    .Q_N(_1514_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net123),
    .D(_0217_),
    .Q_N(_1513_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net123),
    .D(_0218_),
    .Q_N(_1512_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer[7] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net142),
    .D(_0219_),
    .Q_N(_1511_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net141),
    .D(_0220_),
    .Q_N(_1510_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net142),
    .D(_0221_),
    .Q_N(_1509_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net141),
    .D(_0222_),
    .Q_N(_1508_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.rx_buffer_counter[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0]$_DFF_PN1_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net149),
    .D(_0120_),
    .Q_N(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[0] ),
    .Q(_1592_));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net142),
    .D(_0005_),
    .Q_N(_1580_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2]$_DFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net142),
    .D(_0006_),
    .Q_N(_1581_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3]$_DFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net147),
    .D(_0007_),
    .Q_N(_1582_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4]$_DFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net149),
    .D(_0008_),
    .Q_N(_1507_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.state[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net126),
    .D(_0223_),
    .Q_N(_0062_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net126),
    .D(_0224_),
    .Q_N(_0065_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net126),
    .D(_0225_),
    .Q_N(_0068_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net126),
    .D(_0226_),
    .Q_N(_0071_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[3] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net126),
    .D(_0227_),
    .Q_N(_0074_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[4] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net126),
    .D(_0228_),
    .Q_N(_0077_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[5] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0229_),
    .Q_N(_0080_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[6] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net127),
    .D(_0230_),
    .Q_N(_1506_),
    .Q(\rsa_spi_wrapper_i.spi_miso ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net142),
    .D(_0231_),
    .Q_N(_1505_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[0] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net143),
    .D(_0232_),
    .Q_N(_1504_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[1] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net143),
    .D(_0233_),
    .Q_N(_1503_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[2] ));
 sg13g2_dfrbp_1 \rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net142),
    .D(_0234_),
    .Q_N(_1502_),
    .Q(\rsa_spi_wrapper_i.spi_wrapper_i.spi_reg_inst.tx_buffer_counter[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net116),
    .D(_0235_),
    .Q_N(_1501_),
    .Q(\rsa_unit_i.mmm_multiply.A_bit ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net112),
    .D(_0236_),
    .Q_N(_0025_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net112),
    .D(_0237_),
    .Q_N(_0026_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net112),
    .D(_0238_),
    .Q_N(_0028_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net112),
    .D(_0239_),
    .Q_N(_0030_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net113),
    .D(_0240_),
    .Q_N(_0032_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net113),
    .D(_0241_),
    .Q_N(_0034_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net113),
    .D(_0242_),
    .Q_N(_0036_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net112),
    .D(_0243_),
    .Q_N(_0038_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net112),
    .D(_0244_),
    .Q_N(_0040_),
    .Q(\rsa_unit_i.mmm_multiply.shiftreg_A_aux.A_aux[9] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net115),
    .D(_0245_),
    .Q_N(_0044_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.fa_bit0.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net112),
    .D(_0246_),
    .Q_N(_0043_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[1].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net115),
    .D(_0247_),
    .Q_N(_0045_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[2].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net115),
    .D(_0248_),
    .Q_N(_0046_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[3].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net115),
    .D(_0249_),
    .Q_N(_0047_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[4].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net115),
    .D(_0250_),
    .Q_N(_0048_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[5].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net115),
    .D(_0251_),
    .Q_N(_0049_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[6].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net115),
    .D(_0252_),
    .Q_N(_0050_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[7].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_reg_rji.reg_rji[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net116),
    .D(_0253_),
    .Q_N(_0051_),
    .Q(\rsa_unit_i.mmm_multiply.adder2.gen_fa[8].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net116),
    .D(_0254_),
    .Q_N(_1500_),
    .Q(\rsa_unit_i.R_i[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(_0255_),
    .Q_N(_0027_),
    .Q(\rsa_unit_i.R_i[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net113),
    .D(_0256_),
    .Q_N(_0029_),
    .Q(\rsa_unit_i.R_i[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net120),
    .D(_0257_),
    .Q_N(_0031_),
    .Q(\rsa_unit_i.R_i[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net114),
    .D(_0258_),
    .Q_N(_0033_),
    .Q(\rsa_unit_i.R_i[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(_0259_),
    .Q_N(_0035_),
    .Q(\rsa_unit_i.R_i[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(_0260_),
    .Q_N(_0037_),
    .Q(\rsa_unit_i.R_i[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(_0261_),
    .Q_N(_0039_),
    .Q(\rsa_unit_i.R_i[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net114),
    .D(_0262_),
    .Q_N(_0041_),
    .Q(\rsa_unit_i.R_i[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_multiply.shiftreg_result.R_i[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net112),
    .D(_0263_),
    .Q_N(_0042_),
    .Q(\rsa_unit_i.R_i[9] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0264_),
    .Q_N(_1499_),
    .Q(\rsa_unit_i.mmm_square.A_bit ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net132),
    .D(_0265_),
    .Q_N(_0083_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net132),
    .D(_0266_),
    .Q_N(_0086_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net132),
    .D(_0267_),
    .Q_N(_0089_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net132),
    .D(_0268_),
    .Q_N(_0092_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net131),
    .D(_0269_),
    .Q_N(_0095_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net135),
    .D(_0270_),
    .Q_N(_0098_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net135),
    .D(_0271_),
    .Q_N(_0101_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net131),
    .D(_0272_),
    .Q_N(_0104_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0273_),
    .Q_N(_1498_),
    .Q(\rsa_unit_i.mmm_square.shiftreg_A_aux.A_aux[9] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net130),
    .D(_0274_),
    .Q_N(_0109_),
    .Q(\rsa_unit_i.mmm_square.adder2.fa_bit0.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net134),
    .D(_0275_),
    .Q_N(_0107_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[1].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0276_),
    .Q_N(_0110_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[2].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net135),
    .D(_0277_),
    .Q_N(_0112_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[3].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0278_),
    .Q_N(_0114_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[4].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0279_),
    .Q_N(_0116_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[5].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net131),
    .D(_0280_),
    .Q_N(_0020_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[6].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net131),
    .D(_0281_),
    .Q_N(_0022_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[7].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_reg_rji.reg_rji[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net130),
    .D(_0282_),
    .Q_N(_0024_),
    .Q(\rsa_unit_i.mmm_square.adder2.gen_fa[8].fa.HA1.a ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net117),
    .D(_0283_),
    .Q_N(_0084_),
    .Q(\rsa_unit_i.P_i[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net134),
    .D(_0284_),
    .Q_N(_0087_),
    .Q(\rsa_unit_i.P_i[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0285_),
    .Q_N(_0090_),
    .Q(\rsa_unit_i.P_i[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net117),
    .D(_0286_),
    .Q_N(_0093_),
    .Q(\rsa_unit_i.P_i[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net130),
    .D(_0287_),
    .Q_N(_0096_),
    .Q(\rsa_unit_i.P_i[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net130),
    .D(_0288_),
    .Q_N(_0099_),
    .Q(\rsa_unit_i.P_i[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net116),
    .D(_0289_),
    .Q_N(_0102_),
    .Q(\rsa_unit_i.P_i[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net116),
    .D(_0290_),
    .Q_N(_0105_),
    .Q(\rsa_unit_i.P_i[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net130),
    .D(_0291_),
    .Q_N(_1497_),
    .Q(\rsa_unit_i.P_i[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.mmm_square.shiftreg_result.R_i[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net130),
    .D(_0292_),
    .Q_N(_1496_),
    .Q(\rsa_unit_i.P_i[9] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net128),
    .D(_0293_),
    .Q_N(_1495_),
    .Q(\rsa_c[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net120),
    .D(_0294_),
    .Q_N(_1494_),
    .Q(\rsa_c[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net118),
    .D(_0295_),
    .Q_N(_1493_),
    .Q(\rsa_c[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net120),
    .D(_0296_),
    .Q_N(_1492_),
    .Q(\rsa_c[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net120),
    .D(_0297_),
    .Q_N(_1491_),
    .Q(\rsa_c[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net128),
    .D(_0298_),
    .Q_N(_1490_),
    .Q(\rsa_c[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net120),
    .D(_0299_),
    .Q_N(_1489_),
    .Q(\rsa_c[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.reg_crypt.C_ex[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net128),
    .D(_0300_),
    .Q_N(_1488_),
    .Q(\rsa_c[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_rounds[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net146),
    .D(_0301_),
    .Q_N(_1487_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_rounds[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_rounds[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net145),
    .D(_0302_),
    .Q_N(_1486_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_rounds[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_rounds[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net145),
    .D(_0303_),
    .Q_N(_1485_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_rounds[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_rounds[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net146),
    .D(_0304_),
    .Q_N(_1484_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_rounds[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_steps[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net132),
    .D(_0305_),
    .Q_N(_1483_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_steps[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_steps[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net132),
    .D(_0306_),
    .Q_N(_1482_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_steps[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_steps[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net132),
    .D(_0307_),
    .Q_N(_1481_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_steps[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.counter_steps[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net132),
    .D(_0308_),
    .Q_N(_1480_),
    .Q(\rsa_unit_i.rsa_control_fsm.counter_steps[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net139),
    .D(_0309_),
    .Q_N(_1479_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[0] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net140),
    .D(_0310_),
    .Q_N(_1478_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net144),
    .D(_0311_),
    .Q_N(_1477_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net144),
    .D(_0312_),
    .Q_N(_1476_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(_0313_),
    .Q_N(_1475_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[4] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net140),
    .D(_0314_),
    .Q_N(_1474_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[5] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net139),
    .D(_0315_),
    .Q_N(_1473_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.exp[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net146),
    .D(_0316_),
    .Q_N(_1583_),
    .Q(\rsa_unit_i.rsa_control_fsm.exp[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[10]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(_0009_),
    .Q_N(_1584_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[10] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[11]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net136),
    .D(_0010_),
    .Q_N(_0055_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[11] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net133),
    .D(_0011_),
    .Q_N(_1585_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[1] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[2]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net139),
    .D(_0012_),
    .Q_N(_1586_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[2] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[3]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net133),
    .D(_0013_),
    .Q_N(_1587_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[3] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[4]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net145),
    .D(_0014_),
    .Q_N(_0058_),
    .Q(eoc_rsa));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[5]$_DFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net133),
    .D(_0015_),
    .Q_N(_1588_),
    .Q(\rsa_unit_i.rsa_control_fsm.increment_rounds ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[6]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net144),
    .D(_0016_),
    .Q_N(_1589_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[6] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[7]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net133),
    .D(_0017_),
    .Q_N(_1590_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[7] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[8]$_DFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net134),
    .D(_0018_),
    .Q_N(_0057_),
    .Q(\rsa_unit_i.rsa_control_fsm.state[8] ));
 sg13g2_dfrbp_1 \rsa_unit_i.rsa_control_fsm.state[9]$_DFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net145),
    .D(_0019_),
    .Q_N(_0054_),
    .Q(\rsa_unit_i.rsa_control_fsm.load_exp ));
 sg13g2_dfrbp_1 \synchronizer_spi_clk_inst.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net149),
    .D(_0317_),
    .Q_N(_1472_),
    .Q(\synchronizer_spi_clk_inst.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_clk_inst.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net149),
    .D(_0318_),
    .Q_N(_1471_),
    .Q(\rsa_spi_wrapper_i.spi_clk ));
 sg13g2_dfrbp_1 \synchronizer_spi_cs_n_inst.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net149),
    .D(_0319_),
    .Q_N(_1470_),
    .Q(\synchronizer_spi_cs_n_inst.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_cs_n_inst.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net149),
    .D(_0320_),
    .Q_N(_0052_),
    .Q(\rsa_spi_wrapper_i.spi_cs_n ));
 sg13g2_dfrbp_1 \synchronizer_spi_mode_cpha.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net148),
    .D(_0321_),
    .Q_N(_1469_),
    .Q(\synchronizer_spi_mode_cpha.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_mode_cpha.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net148),
    .D(_0322_),
    .Q_N(_1468_),
    .Q(cpha_sync));
 sg13g2_dfrbp_1 \synchronizer_spi_mode_cpol.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net148),
    .D(_0323_),
    .Q_N(_1467_),
    .Q(\synchronizer_spi_mode_cpol.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_mode_cpol.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net148),
    .D(_0324_),
    .Q_N(_1466_),
    .Q(cpol_sync));
 sg13g2_dfrbp_1 \synchronizer_spi_mosi_inst.gen_reclocking[0].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net143),
    .D(_0325_),
    .Q_N(_1465_),
    .Q(\synchronizer_spi_mosi_inst.data_sync[1] ));
 sg13g2_dfrbp_1 \synchronizer_spi_mosi_inst.gen_reclocking[1].reclocking_i0.data_sync$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net143),
    .D(_0326_),
    .Q_N(_1464_),
    .Q(\rsa_spi_wrapper_i.spi_mosi ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[6]),
    .X(net8));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[0]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[1]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[2]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[3]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[4]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[5]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[6]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[7]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout25 (.A(_0599_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0598_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0369_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0559_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0368_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0701_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0558_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0456_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0392_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0669_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_0531_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0394_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1020_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0389_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0379_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0997_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0968_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0639_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0481_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0383_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0363_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1330_),
    .X(net46));
 sg13g2_buf_4 fanout47 (.X(net47),
    .A(_1292_));
 sg13g2_buf_4 fanout48 (.X(net48),
    .A(_1209_));
 sg13g2_buf_2 fanout49 (.A(_0881_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0632_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0566_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0473_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0454_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0373_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0362_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1361_),
    .X(net56));
 sg13g2_buf_4 fanout57 (.X(net57),
    .A(_1319_));
 sg13g2_buf_2 fanout58 (.A(_1297_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1226_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0568_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0377_),
    .X(net61));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(_1309_));
 sg13g2_buf_2 fanout63 (.A(_1279_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1187_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1184_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0705_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0569_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0562_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0448_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0371_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1289_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_1249_));
 sg13g2_buf_2 fanout73 (.A(_1201_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0938_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0898_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0875_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0729_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0616_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0565_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0532_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1307_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1295_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1287_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1260_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1258_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1256_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1222_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1163_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_0901_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_0874_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_0793_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0703_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_0564_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0460_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0385_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0355_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1362_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1270_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_1269_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1268_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_1267_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_1266_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_1265_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_1264_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_1257_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_1255_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_1254_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1232_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1211_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1207_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_1162_),
    .X(net111));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(net114));
 sg13g2_buf_2 fanout113 (.A(net114),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(net115));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(net117));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(net117));
 sg13g2_buf_2 fanout117 (.A(net129),
    .X(net117));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(net121));
 sg13g2_buf_2 fanout119 (.A(net121),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(net121));
 sg13g2_buf_2 fanout121 (.A(net129),
    .X(net121));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(net125));
 sg13g2_buf_2 fanout123 (.A(net125),
    .X(net123));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(net125));
 sg13g2_buf_2 fanout125 (.A(net129),
    .X(net125));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(net128));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(net128));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(net129));
 sg13g2_buf_1 fanout129 (.A(net1),
    .X(net129));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(net136));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(net135));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(net134));
 sg13g2_buf_2 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(net135),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(net151),
    .X(net136));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net140));
 sg13g2_buf_2 fanout138 (.A(net140),
    .X(net138));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net140));
 sg13g2_buf_2 fanout140 (.A(net151),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net143));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net143));
 sg13g2_buf_2 fanout143 (.A(net151),
    .X(net143));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net146));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net146));
 sg13g2_buf_2 fanout146 (.A(net150),
    .X(net146));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(net150));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net150));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(net150));
 sg13g2_buf_1 fanout150 (.A(net151),
    .X(net150));
 sg13g2_buf_1 fanout151 (.A(net1),
    .X(net151));
 sg13g2_tielo _2967__152 (.L_LO(net152));
 sg13g2_tielo _2968__153 (.L_LO(net153));
 sg13g2_tielo _2969__154 (.L_LO(net154));
 sg13g2_tiehi _2964__156 (.L_HI(net156));
 sg13g2_tiehi _2965__157 (.L_HI(net157));
 sg13g2_tiehi _2966__158 (.L_HI(net158));
 sg13g2_tiehi _2970__159 (.L_HI(net159));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_leaf_29_clk));
 sg13g2_inv_2 clkload2 (.A(clknet_leaf_30_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_28_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_leaf_11_clk));
 sg13g2_inv_2 clkload5 (.A(clknet_leaf_22_clk));
 sg13g2_inv_4 clkload6 (.A(clknet_leaf_26_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_27_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_4 FILLER_0_56 ();
 sg13g2_fill_1 FILLER_0_60 ();
 sg13g2_fill_1 FILLER_0_99 ();
 sg13g2_fill_1 FILLER_0_113 ();
 sg13g2_fill_1 FILLER_0_140 ();
 sg13g2_decap_4 FILLER_0_146 ();
 sg13g2_fill_1 FILLER_0_150 ();
 sg13g2_fill_1 FILLER_0_171 ();
 sg13g2_fill_1 FILLER_0_176 ();
 sg13g2_fill_1 FILLER_0_185 ();
 sg13g2_decap_8 FILLER_0_198 ();
 sg13g2_fill_2 FILLER_0_205 ();
 sg13g2_fill_2 FILLER_0_220 ();
 sg13g2_fill_2 FILLER_0_250 ();
 sg13g2_fill_1 FILLER_0_289 ();
 sg13g2_fill_2 FILLER_0_299 ();
 sg13g2_fill_2 FILLER_0_314 ();
 sg13g2_fill_2 FILLER_0_324 ();
 sg13g2_fill_1 FILLER_0_326 ();
 sg13g2_fill_1 FILLER_0_335 ();
 sg13g2_fill_2 FILLER_0_341 ();
 sg13g2_fill_1 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_4 FILLER_0_425 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_fill_1 FILLER_1_49 ();
 sg13g2_fill_1 FILLER_1_68 ();
 sg13g2_fill_1 FILLER_1_81 ();
 sg13g2_fill_2 FILLER_1_107 ();
 sg13g2_decap_4 FILLER_1_133 ();
 sg13g2_fill_2 FILLER_1_202 ();
 sg13g2_fill_1 FILLER_1_204 ();
 sg13g2_fill_1 FILLER_1_241 ();
 sg13g2_fill_2 FILLER_1_246 ();
 sg13g2_fill_1 FILLER_1_253 ();
 sg13g2_fill_1 FILLER_1_266 ();
 sg13g2_fill_2 FILLER_1_273 ();
 sg13g2_fill_1 FILLER_1_275 ();
 sg13g2_fill_2 FILLER_1_283 ();
 sg13g2_fill_1 FILLER_1_285 ();
 sg13g2_fill_1 FILLER_1_299 ();
 sg13g2_fill_2 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_362 ();
 sg13g2_decap_8 FILLER_1_369 ();
 sg13g2_decap_8 FILLER_1_376 ();
 sg13g2_decap_8 FILLER_1_383 ();
 sg13g2_decap_8 FILLER_1_390 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_8 FILLER_1_404 ();
 sg13g2_decap_8 FILLER_1_411 ();
 sg13g2_decap_8 FILLER_1_418 ();
 sg13g2_decap_4 FILLER_1_425 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_fill_1 FILLER_2_68 ();
 sg13g2_fill_2 FILLER_2_83 ();
 sg13g2_fill_1 FILLER_2_90 ();
 sg13g2_fill_2 FILLER_2_97 ();
 sg13g2_fill_1 FILLER_2_114 ();
 sg13g2_fill_2 FILLER_2_129 ();
 sg13g2_fill_2 FILLER_2_141 ();
 sg13g2_fill_1 FILLER_2_167 ();
 sg13g2_fill_1 FILLER_2_176 ();
 sg13g2_fill_1 FILLER_2_190 ();
 sg13g2_decap_4 FILLER_2_196 ();
 sg13g2_fill_2 FILLER_2_205 ();
 sg13g2_fill_1 FILLER_2_207 ();
 sg13g2_fill_2 FILLER_2_242 ();
 sg13g2_fill_2 FILLER_2_274 ();
 sg13g2_fill_2 FILLER_2_291 ();
 sg13g2_fill_1 FILLER_2_356 ();
 sg13g2_fill_2 FILLER_2_365 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_decap_4 FILLER_3_99 ();
 sg13g2_fill_2 FILLER_3_116 ();
 sg13g2_fill_1 FILLER_3_156 ();
 sg13g2_decap_8 FILLER_3_183 ();
 sg13g2_fill_2 FILLER_3_190 ();
 sg13g2_fill_1 FILLER_3_192 ();
 sg13g2_fill_2 FILLER_3_214 ();
 sg13g2_fill_1 FILLER_3_216 ();
 sg13g2_fill_1 FILLER_3_248 ();
 sg13g2_fill_1 FILLER_3_286 ();
 sg13g2_fill_1 FILLER_3_298 ();
 sg13g2_fill_1 FILLER_3_307 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_decap_8 FILLER_3_384 ();
 sg13g2_decap_8 FILLER_3_391 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_8 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_3_412 ();
 sg13g2_decap_8 FILLER_3_419 ();
 sg13g2_decap_4 FILLER_3_426 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_4 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_125 ();
 sg13g2_fill_1 FILLER_4_132 ();
 sg13g2_decap_8 FILLER_4_188 ();
 sg13g2_fill_2 FILLER_4_199 ();
 sg13g2_fill_1 FILLER_4_209 ();
 sg13g2_fill_1 FILLER_4_215 ();
 sg13g2_fill_1 FILLER_4_220 ();
 sg13g2_fill_1 FILLER_4_249 ();
 sg13g2_fill_2 FILLER_4_306 ();
 sg13g2_fill_1 FILLER_4_313 ();
 sg13g2_fill_1 FILLER_4_319 ();
 sg13g2_fill_1 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_8 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_4_412 ();
 sg13g2_decap_8 FILLER_4_419 ();
 sg13g2_decap_4 FILLER_4_426 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_4 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_32 ();
 sg13g2_fill_2 FILLER_5_102 ();
 sg13g2_fill_1 FILLER_5_124 ();
 sg13g2_fill_1 FILLER_5_160 ();
 sg13g2_fill_1 FILLER_5_185 ();
 sg13g2_fill_1 FILLER_5_196 ();
 sg13g2_fill_2 FILLER_5_204 ();
 sg13g2_fill_1 FILLER_5_211 ();
 sg13g2_fill_2 FILLER_5_217 ();
 sg13g2_fill_1 FILLER_5_219 ();
 sg13g2_fill_1 FILLER_5_228 ();
 sg13g2_fill_2 FILLER_5_236 ();
 sg13g2_fill_1 FILLER_5_238 ();
 sg13g2_fill_1 FILLER_5_243 ();
 sg13g2_fill_2 FILLER_5_248 ();
 sg13g2_fill_1 FILLER_5_254 ();
 sg13g2_fill_1 FILLER_5_290 ();
 sg13g2_fill_2 FILLER_5_334 ();
 sg13g2_fill_1 FILLER_5_359 ();
 sg13g2_fill_2 FILLER_5_365 ();
 sg13g2_fill_1 FILLER_5_367 ();
 sg13g2_fill_2 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_409 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_fill_2 FILLER_6_28 ();
 sg13g2_fill_1 FILLER_6_30 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_fill_1 FILLER_6_42 ();
 sg13g2_fill_1 FILLER_6_65 ();
 sg13g2_fill_1 FILLER_6_87 ();
 sg13g2_fill_1 FILLER_6_107 ();
 sg13g2_fill_2 FILLER_6_166 ();
 sg13g2_fill_2 FILLER_6_178 ();
 sg13g2_fill_1 FILLER_6_185 ();
 sg13g2_fill_1 FILLER_6_190 ();
 sg13g2_fill_2 FILLER_6_196 ();
 sg13g2_fill_1 FILLER_6_198 ();
 sg13g2_fill_2 FILLER_6_203 ();
 sg13g2_fill_1 FILLER_6_284 ();
 sg13g2_fill_1 FILLER_6_327 ();
 sg13g2_fill_2 FILLER_6_353 ();
 sg13g2_decap_4 FILLER_6_381 ();
 sg13g2_fill_1 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_390 ();
 sg13g2_decap_8 FILLER_6_397 ();
 sg13g2_decap_8 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_411 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_decap_4 FILLER_6_425 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_4 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_61 ();
 sg13g2_fill_1 FILLER_7_87 ();
 sg13g2_fill_1 FILLER_7_92 ();
 sg13g2_fill_1 FILLER_7_113 ();
 sg13g2_fill_2 FILLER_7_150 ();
 sg13g2_fill_2 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_311 ();
 sg13g2_fill_2 FILLER_7_321 ();
 sg13g2_fill_1 FILLER_7_323 ();
 sg13g2_fill_1 FILLER_7_333 ();
 sg13g2_fill_1 FILLER_7_342 ();
 sg13g2_fill_1 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_409 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_fill_2 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_44 ();
 sg13g2_fill_2 FILLER_8_54 ();
 sg13g2_fill_1 FILLER_8_88 ();
 sg13g2_fill_1 FILLER_8_190 ();
 sg13g2_fill_1 FILLER_8_195 ();
 sg13g2_fill_2 FILLER_8_229 ();
 sg13g2_fill_1 FILLER_8_306 ();
 sg13g2_fill_1 FILLER_8_312 ();
 sg13g2_fill_1 FILLER_8_345 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_fill_2 FILLER_8_394 ();
 sg13g2_fill_1 FILLER_8_396 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_fill_2 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_127 ();
 sg13g2_fill_1 FILLER_9_129 ();
 sg13g2_fill_2 FILLER_9_189 ();
 sg13g2_fill_1 FILLER_9_196 ();
 sg13g2_fill_1 FILLER_9_205 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_fill_2 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_272 ();
 sg13g2_fill_1 FILLER_9_311 ();
 sg13g2_fill_2 FILLER_9_317 ();
 sg13g2_fill_1 FILLER_9_319 ();
 sg13g2_fill_1 FILLER_9_332 ();
 sg13g2_fill_2 FILLER_9_382 ();
 sg13g2_fill_1 FILLER_9_422 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_4 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_25 ();
 sg13g2_fill_2 FILLER_10_62 ();
 sg13g2_fill_1 FILLER_10_110 ();
 sg13g2_fill_2 FILLER_10_115 ();
 sg13g2_fill_1 FILLER_10_132 ();
 sg13g2_fill_1 FILLER_10_138 ();
 sg13g2_fill_1 FILLER_10_191 ();
 sg13g2_fill_1 FILLER_10_227 ();
 sg13g2_fill_2 FILLER_10_233 ();
 sg13g2_fill_1 FILLER_10_240 ();
 sg13g2_fill_1 FILLER_10_264 ();
 sg13g2_fill_2 FILLER_10_290 ();
 sg13g2_fill_1 FILLER_10_335 ();
 sg13g2_decap_4 FILLER_10_362 ();
 sg13g2_fill_2 FILLER_10_381 ();
 sg13g2_fill_2 FILLER_10_392 ();
 sg13g2_fill_2 FILLER_11_109 ();
 sg13g2_fill_2 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_204 ();
 sg13g2_fill_1 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_215 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_fill_1 FILLER_11_251 ();
 sg13g2_fill_1 FILLER_11_264 ();
 sg13g2_fill_2 FILLER_11_274 ();
 sg13g2_fill_1 FILLER_11_313 ();
 sg13g2_fill_2 FILLER_11_325 ();
 sg13g2_fill_1 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_362 ();
 sg13g2_fill_2 FILLER_11_390 ();
 sg13g2_fill_2 FILLER_11_402 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_8 ();
 sg13g2_fill_1 FILLER_12_10 ();
 sg13g2_decap_8 FILLER_12_15 ();
 sg13g2_fill_2 FILLER_12_35 ();
 sg13g2_fill_1 FILLER_12_41 ();
 sg13g2_fill_1 FILLER_12_156 ();
 sg13g2_fill_1 FILLER_12_167 ();
 sg13g2_fill_1 FILLER_12_176 ();
 sg13g2_fill_2 FILLER_12_217 ();
 sg13g2_fill_2 FILLER_12_296 ();
 sg13g2_fill_2 FILLER_12_303 ();
 sg13g2_fill_1 FILLER_12_315 ();
 sg13g2_fill_1 FILLER_12_336 ();
 sg13g2_fill_1 FILLER_12_367 ();
 sg13g2_fill_2 FILLER_12_373 ();
 sg13g2_fill_1 FILLER_12_375 ();
 sg13g2_fill_2 FILLER_12_391 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_1 FILLER_13_26 ();
 sg13g2_fill_2 FILLER_13_80 ();
 sg13g2_fill_1 FILLER_13_90 ();
 sg13g2_fill_2 FILLER_13_96 ();
 sg13g2_fill_2 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_115 ();
 sg13g2_fill_1 FILLER_13_131 ();
 sg13g2_fill_2 FILLER_13_136 ();
 sg13g2_fill_2 FILLER_13_185 ();
 sg13g2_fill_1 FILLER_13_187 ();
 sg13g2_fill_1 FILLER_13_191 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_212 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_fill_1 FILLER_13_276 ();
 sg13g2_fill_2 FILLER_13_306 ();
 sg13g2_fill_2 FILLER_13_334 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_396 ();
 sg13g2_fill_2 FILLER_13_402 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_37 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_2 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_177 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_decap_4 FILLER_14_183 ();
 sg13g2_fill_1 FILLER_14_216 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_fill_1 FILLER_14_292 ();
 sg13g2_fill_1 FILLER_14_301 ();
 sg13g2_fill_2 FILLER_14_357 ();
 sg13g2_fill_1 FILLER_14_359 ();
 sg13g2_fill_2 FILLER_14_364 ();
 sg13g2_fill_2 FILLER_14_397 ();
 sg13g2_fill_1 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_412 ();
 sg13g2_fill_2 FILLER_14_419 ();
 sg13g2_fill_1 FILLER_14_421 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_2 FILLER_15_18 ();
 sg13g2_fill_1 FILLER_15_20 ();
 sg13g2_fill_2 FILLER_15_31 ();
 sg13g2_fill_2 FILLER_15_69 ();
 sg13g2_fill_2 FILLER_15_95 ();
 sg13g2_fill_1 FILLER_15_97 ();
 sg13g2_fill_2 FILLER_15_103 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_146 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_fill_1 FILLER_15_164 ();
 sg13g2_fill_2 FILLER_15_181 ();
 sg13g2_fill_1 FILLER_15_183 ();
 sg13g2_fill_1 FILLER_15_189 ();
 sg13g2_decap_4 FILLER_15_198 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_1 FILLER_15_208 ();
 sg13g2_decap_4 FILLER_15_214 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_316 ();
 sg13g2_fill_2 FILLER_15_345 ();
 sg13g2_fill_2 FILLER_15_355 ();
 sg13g2_fill_2 FILLER_15_402 ();
 sg13g2_fill_2 FILLER_16_26 ();
 sg13g2_fill_2 FILLER_16_43 ();
 sg13g2_fill_1 FILLER_16_57 ();
 sg13g2_fill_1 FILLER_16_68 ();
 sg13g2_fill_2 FILLER_16_73 ();
 sg13g2_fill_1 FILLER_16_80 ();
 sg13g2_fill_2 FILLER_16_86 ();
 sg13g2_fill_1 FILLER_16_92 ();
 sg13g2_fill_1 FILLER_16_119 ();
 sg13g2_fill_1 FILLER_16_124 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_164 ();
 sg13g2_fill_1 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_185 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_219 ();
 sg13g2_fill_1 FILLER_16_287 ();
 sg13g2_fill_1 FILLER_16_298 ();
 sg13g2_fill_2 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_331 ();
 sg13g2_fill_1 FILLER_16_337 ();
 sg13g2_fill_1 FILLER_16_369 ();
 sg13g2_decap_4 FILLER_16_382 ();
 sg13g2_fill_1 FILLER_16_386 ();
 sg13g2_fill_2 FILLER_16_412 ();
 sg13g2_fill_1 FILLER_16_414 ();
 sg13g2_decap_8 FILLER_16_423 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_fill_2 FILLER_17_110 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_117 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_fill_1 FILLER_17_150 ();
 sg13g2_fill_1 FILLER_17_159 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_175 ();
 sg13g2_fill_2 FILLER_17_202 ();
 sg13g2_fill_2 FILLER_17_306 ();
 sg13g2_fill_2 FILLER_17_355 ();
 sg13g2_fill_2 FILLER_17_366 ();
 sg13g2_fill_1 FILLER_17_377 ();
 sg13g2_fill_2 FILLER_17_402 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_4 ();
 sg13g2_fill_2 FILLER_18_32 ();
 sg13g2_fill_1 FILLER_18_34 ();
 sg13g2_fill_1 FILLER_18_76 ();
 sg13g2_fill_1 FILLER_18_81 ();
 sg13g2_fill_1 FILLER_18_87 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_134 ();
 sg13g2_fill_2 FILLER_18_256 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_decap_4 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_328 ();
 sg13g2_fill_1 FILLER_18_336 ();
 sg13g2_fill_1 FILLER_18_346 ();
 sg13g2_fill_1 FILLER_18_358 ();
 sg13g2_fill_1 FILLER_18_364 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_1 FILLER_18_403 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_fill_2 FILLER_18_424 ();
 sg13g2_fill_1 FILLER_18_426 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_9 ();
 sg13g2_fill_1 FILLER_19_22 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_33 ();
 sg13g2_fill_2 FILLER_19_44 ();
 sg13g2_fill_1 FILLER_19_46 ();
 sg13g2_fill_2 FILLER_19_140 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_fill_1 FILLER_19_206 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_fill_2 FILLER_19_256 ();
 sg13g2_fill_2 FILLER_19_284 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_fill_2 FILLER_19_291 ();
 sg13g2_fill_1 FILLER_19_293 ();
 sg13g2_fill_2 FILLER_19_320 ();
 sg13g2_fill_1 FILLER_19_327 ();
 sg13g2_fill_1 FILLER_19_333 ();
 sg13g2_fill_1 FILLER_19_348 ();
 sg13g2_fill_1 FILLER_19_355 ();
 sg13g2_fill_2 FILLER_19_385 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_27 ();
 sg13g2_fill_1 FILLER_20_54 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_fill_2 FILLER_20_74 ();
 sg13g2_fill_2 FILLER_20_86 ();
 sg13g2_fill_1 FILLER_20_88 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_104 ();
 sg13g2_fill_1 FILLER_20_116 ();
 sg13g2_fill_2 FILLER_20_172 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_fill_1 FILLER_20_262 ();
 sg13g2_decap_4 FILLER_20_289 ();
 sg13g2_fill_2 FILLER_20_293 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_26 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_205 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_228 ();
 sg13g2_fill_2 FILLER_21_240 ();
 sg13g2_fill_1 FILLER_21_242 ();
 sg13g2_decap_4 FILLER_21_246 ();
 sg13g2_fill_1 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_decap_4 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_decap_4 FILLER_21_288 ();
 sg13g2_decap_4 FILLER_21_301 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_1 FILLER_21_323 ();
 sg13g2_decap_4 FILLER_21_328 ();
 sg13g2_fill_2 FILLER_21_332 ();
 sg13g2_fill_2 FILLER_21_343 ();
 sg13g2_fill_1 FILLER_21_390 ();
 sg13g2_fill_2 FILLER_22_8 ();
 sg13g2_fill_1 FILLER_22_10 ();
 sg13g2_decap_8 FILLER_22_34 ();
 sg13g2_fill_1 FILLER_22_41 ();
 sg13g2_decap_4 FILLER_22_78 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_fill_2 FILLER_22_137 ();
 sg13g2_fill_1 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_fill_2 FILLER_22_284 ();
 sg13g2_fill_1 FILLER_22_317 ();
 sg13g2_fill_2 FILLER_22_349 ();
 sg13g2_fill_2 FILLER_22_356 ();
 sg13g2_fill_1 FILLER_22_358 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_1 FILLER_22_365 ();
 sg13g2_fill_2 FILLER_22_384 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_fill_1 FILLER_22_392 ();
 sg13g2_fill_1 FILLER_22_403 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_13 ();
 sg13g2_fill_2 FILLER_23_53 ();
 sg13g2_fill_1 FILLER_23_55 ();
 sg13g2_fill_1 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_228 ();
 sg13g2_fill_2 FILLER_23_244 ();
 sg13g2_fill_1 FILLER_23_246 ();
 sg13g2_decap_4 FILLER_23_273 ();
 sg13g2_fill_2 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_2 ();
 sg13g2_fill_2 FILLER_24_143 ();
 sg13g2_fill_1 FILLER_24_162 ();
 sg13g2_fill_1 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_176 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_fill_1 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_fill_2 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_decap_4 FILLER_24_238 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_253 ();
 sg13g2_decap_8 FILLER_24_281 ();
 sg13g2_fill_2 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_290 ();
 sg13g2_fill_1 FILLER_24_343 ();
 sg13g2_decap_4 FILLER_24_368 ();
 sg13g2_fill_2 FILLER_24_376 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_fill_1 FILLER_25_55 ();
 sg13g2_fill_1 FILLER_25_92 ();
 sg13g2_fill_2 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_fill_1 FILLER_25_188 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_318 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_fill_1 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_179 ();
 sg13g2_fill_1 FILLER_26_190 ();
 sg13g2_fill_1 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_fill_2 FILLER_26_215 ();
 sg13g2_decap_4 FILLER_26_227 ();
 sg13g2_decap_4 FILLER_26_241 ();
 sg13g2_decap_4 FILLER_26_255 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_215 ();
 sg13g2_fill_2 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_244 ();
 sg13g2_fill_2 FILLER_27_286 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_fill_2 FILLER_27_387 ();
 sg13g2_fill_2 FILLER_27_402 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_fill_1 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_fill_1 FILLER_28_120 ();
 sg13g2_fill_2 FILLER_28_147 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_214 ();
 sg13g2_fill_1 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_401 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_1 FILLER_29_79 ();
 sg13g2_fill_2 FILLER_29_288 ();
 sg13g2_fill_1 FILLER_29_290 ();
 sg13g2_fill_1 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_367 ();
 sg13g2_fill_1 FILLER_29_402 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_1 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_119 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_fill_1 FILLER_30_160 ();
 sg13g2_fill_2 FILLER_30_166 ();
 sg13g2_fill_1 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_2 FILLER_30_197 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_decap_4 FILLER_30_236 ();
 sg13g2_fill_1 FILLER_30_240 ();
 sg13g2_decap_4 FILLER_30_261 ();
 sg13g2_fill_1 FILLER_30_265 ();
 sg13g2_decap_8 FILLER_30_274 ();
 sg13g2_decap_4 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_391 ();
 sg13g2_fill_1 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_fill_2 FILLER_31_43 ();
 sg13g2_fill_1 FILLER_31_45 ();
 sg13g2_fill_1 FILLER_31_66 ();
 sg13g2_fill_1 FILLER_31_103 ();
 sg13g2_fill_2 FILLER_31_109 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_fill_1 FILLER_31_225 ();
 sg13g2_fill_1 FILLER_31_252 ();
 sg13g2_fill_2 FILLER_31_279 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_383 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_11 ();
 sg13g2_fill_1 FILLER_32_32 ();
 sg13g2_fill_2 FILLER_32_59 ();
 sg13g2_fill_2 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_fill_1 FILLER_32_231 ();
 sg13g2_fill_2 FILLER_32_275 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_27 ();
 sg13g2_fill_2 FILLER_33_38 ();
 sg13g2_fill_2 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_2 FILLER_33_142 ();
 sg13g2_fill_1 FILLER_33_144 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_351 ();
 sg13g2_fill_2 FILLER_33_392 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_167 ();
 sg13g2_fill_1 FILLER_34_169 ();
 sg13g2_fill_2 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_fill_2 FILLER_34_236 ();
 sg13g2_fill_2 FILLER_34_262 ();
 sg13g2_fill_2 FILLER_34_415 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_2 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_37 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_114 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_157 ();
 sg13g2_fill_1 FILLER_35_162 ();
 sg13g2_fill_2 FILLER_35_194 ();
 sg13g2_fill_1 FILLER_35_196 ();
 sg13g2_fill_2 FILLER_35_223 ();
 sg13g2_fill_1 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_301 ();
 sg13g2_fill_2 FILLER_35_318 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_fill_1 FILLER_35_398 ();
 sg13g2_fill_1 FILLER_36_75 ();
 sg13g2_fill_1 FILLER_36_132 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_fill_2 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_236 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_290 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_419 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_99 ();
 sg13g2_fill_1 FILLER_37_117 ();
 sg13g2_fill_1 FILLER_37_162 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_fill_2 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_257 ();
 sg13g2_fill_2 FILLER_37_392 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_48 ();
 sg13g2_fill_2 FILLER_38_104 ();
 sg13g2_fill_1 FILLER_38_106 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_2 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_232 ();
 sg13g2_fill_1 FILLER_38_344 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_fill_2 FILLER_38_428 ();
endmodule
